`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Linear_p( // @[:@3.2]
  input  [3:0]  io_in_0, // @[:@6.4]
  input  [3:0]  io_in_3, // @[:@6.4]
  input  [3:0]  io_in_5, // @[:@6.4]
  input  [3:0]  io_in_10, // @[:@6.4]
  input  [3:0]  io_in_12, // @[:@6.4]
  input  [3:0]  io_in_13, // @[:@6.4]
  input  [3:0]  io_in_14, // @[:@6.4]
  input  [3:0]  io_in_15, // @[:@6.4]
  input  [3:0]  io_in_19, // @[:@6.4]
  input  [3:0]  io_in_21, // @[:@6.4]
  input  [3:0]  io_in_23, // @[:@6.4]
  input  [3:0]  io_in_25, // @[:@6.4]
  input  [3:0]  io_in_28, // @[:@6.4]
  input  [3:0]  io_in_29, // @[:@6.4]
  input  [3:0]  io_in_30, // @[:@6.4]
  input  [3:0]  io_in_32, // @[:@6.4]
  input  [3:0]  io_in_33, // @[:@6.4]
  input  [3:0]  io_in_34, // @[:@6.4]
  input  [3:0]  io_in_35, // @[:@6.4]
  input  [3:0]  io_in_36, // @[:@6.4]
  input  [3:0]  io_in_37, // @[:@6.4]
  input  [3:0]  io_in_38, // @[:@6.4]
  input  [3:0]  io_in_39, // @[:@6.4]
  input  [3:0]  io_in_40, // @[:@6.4]
  input  [3:0]  io_in_41, // @[:@6.4]
  input  [3:0]  io_in_42, // @[:@6.4]
  input  [3:0]  io_in_43, // @[:@6.4]
  input  [3:0]  io_in_44, // @[:@6.4]
  input  [3:0]  io_in_45, // @[:@6.4]
  input  [3:0]  io_in_46, // @[:@6.4]
  input  [3:0]  io_in_47, // @[:@6.4]
  input  [3:0]  io_in_48, // @[:@6.4]
  input  [3:0]  io_in_49, // @[:@6.4]
  input  [3:0]  io_in_50, // @[:@6.4]
  input  [3:0]  io_in_51, // @[:@6.4]
  input  [3:0]  io_in_52, // @[:@6.4]
  input  [3:0]  io_in_54, // @[:@6.4]
  input  [3:0]  io_in_56, // @[:@6.4]
  input  [3:0]  io_in_59, // @[:@6.4]
  input  [3:0]  io_in_60, // @[:@6.4]
  input  [3:0]  io_in_61, // @[:@6.4]
  input  [3:0]  io_in_62, // @[:@6.4]
  input  [3:0]  io_in_63, // @[:@6.4]
  input  [3:0]  io_in_64, // @[:@6.4]
  input  [3:0]  io_in_65, // @[:@6.4]
  input  [3:0]  io_in_66, // @[:@6.4]
  input  [3:0]  io_in_67, // @[:@6.4]
  input  [3:0]  io_in_68, // @[:@6.4]
  input  [3:0]  io_in_69, // @[:@6.4]
  input  [3:0]  io_in_70, // @[:@6.4]
  input  [3:0]  io_in_71, // @[:@6.4]
  input  [3:0]  io_in_72, // @[:@6.4]
  input  [3:0]  io_in_73, // @[:@6.4]
  input  [3:0]  io_in_74, // @[:@6.4]
  input  [3:0]  io_in_75, // @[:@6.4]
  input  [3:0]  io_in_76, // @[:@6.4]
  input  [3:0]  io_in_77, // @[:@6.4]
  input  [3:0]  io_in_78, // @[:@6.4]
  input  [3:0]  io_in_79, // @[:@6.4]
  input  [3:0]  io_in_80, // @[:@6.4]
  input  [3:0]  io_in_81, // @[:@6.4]
  input  [3:0]  io_in_82, // @[:@6.4]
  input  [3:0]  io_in_83, // @[:@6.4]
  input  [3:0]  io_in_86, // @[:@6.4]
  input  [3:0]  io_in_87, // @[:@6.4]
  input  [3:0]  io_in_88, // @[:@6.4]
  input  [3:0]  io_in_89, // @[:@6.4]
  input  [3:0]  io_in_90, // @[:@6.4]
  input  [3:0]  io_in_91, // @[:@6.4]
  input  [3:0]  io_in_92, // @[:@6.4]
  input  [3:0]  io_in_93, // @[:@6.4]
  input  [3:0]  io_in_94, // @[:@6.4]
  input  [3:0]  io_in_95, // @[:@6.4]
  input  [3:0]  io_in_96, // @[:@6.4]
  input  [3:0]  io_in_97, // @[:@6.4]
  input  [3:0]  io_in_98, // @[:@6.4]
  input  [3:0]  io_in_99, // @[:@6.4]
  input  [3:0]  io_in_100, // @[:@6.4]
  input  [3:0]  io_in_101, // @[:@6.4]
  input  [3:0]  io_in_102, // @[:@6.4]
  input  [3:0]  io_in_103, // @[:@6.4]
  input  [3:0]  io_in_104, // @[:@6.4]
  input  [3:0]  io_in_105, // @[:@6.4]
  input  [3:0]  io_in_106, // @[:@6.4]
  input  [3:0]  io_in_107, // @[:@6.4]
  input  [3:0]  io_in_108, // @[:@6.4]
  input  [3:0]  io_in_109, // @[:@6.4]
  input  [3:0]  io_in_110, // @[:@6.4]
  input  [3:0]  io_in_113, // @[:@6.4]
  input  [3:0]  io_in_114, // @[:@6.4]
  input  [3:0]  io_in_115, // @[:@6.4]
  input  [3:0]  io_in_116, // @[:@6.4]
  input  [3:0]  io_in_117, // @[:@6.4]
  input  [3:0]  io_in_118, // @[:@6.4]
  input  [3:0]  io_in_119, // @[:@6.4]
  input  [3:0]  io_in_120, // @[:@6.4]
  input  [3:0]  io_in_121, // @[:@6.4]
  input  [3:0]  io_in_122, // @[:@6.4]
  input  [3:0]  io_in_123, // @[:@6.4]
  input  [3:0]  io_in_124, // @[:@6.4]
  input  [3:0]  io_in_125, // @[:@6.4]
  input  [3:0]  io_in_126, // @[:@6.4]
  input  [3:0]  io_in_127, // @[:@6.4]
  input  [3:0]  io_in_128, // @[:@6.4]
  input  [3:0]  io_in_129, // @[:@6.4]
  input  [3:0]  io_in_130, // @[:@6.4]
  input  [3:0]  io_in_131, // @[:@6.4]
  input  [3:0]  io_in_132, // @[:@6.4]
  input  [3:0]  io_in_133, // @[:@6.4]
  input  [3:0]  io_in_134, // @[:@6.4]
  input  [3:0]  io_in_135, // @[:@6.4]
  input  [3:0]  io_in_136, // @[:@6.4]
  input  [3:0]  io_in_137, // @[:@6.4]
  input  [3:0]  io_in_138, // @[:@6.4]
  input  [3:0]  io_in_139, // @[:@6.4]
  input  [3:0]  io_in_140, // @[:@6.4]
  input  [3:0]  io_in_142, // @[:@6.4]
  input  [3:0]  io_in_143, // @[:@6.4]
  input  [3:0]  io_in_144, // @[:@6.4]
  input  [3:0]  io_in_145, // @[:@6.4]
  input  [3:0]  io_in_146, // @[:@6.4]
  input  [3:0]  io_in_147, // @[:@6.4]
  input  [3:0]  io_in_148, // @[:@6.4]
  input  [3:0]  io_in_149, // @[:@6.4]
  input  [3:0]  io_in_150, // @[:@6.4]
  input  [3:0]  io_in_151, // @[:@6.4]
  input  [3:0]  io_in_152, // @[:@6.4]
  input  [3:0]  io_in_153, // @[:@6.4]
  input  [3:0]  io_in_154, // @[:@6.4]
  input  [3:0]  io_in_155, // @[:@6.4]
  input  [3:0]  io_in_156, // @[:@6.4]
  input  [3:0]  io_in_157, // @[:@6.4]
  input  [3:0]  io_in_158, // @[:@6.4]
  input  [3:0]  io_in_159, // @[:@6.4]
  input  [3:0]  io_in_160, // @[:@6.4]
  input  [3:0]  io_in_161, // @[:@6.4]
  input  [3:0]  io_in_162, // @[:@6.4]
  input  [3:0]  io_in_163, // @[:@6.4]
  input  [3:0]  io_in_164, // @[:@6.4]
  input  [3:0]  io_in_165, // @[:@6.4]
  input  [3:0]  io_in_166, // @[:@6.4]
  input  [3:0]  io_in_167, // @[:@6.4]
  input  [3:0]  io_in_168, // @[:@6.4]
  input  [3:0]  io_in_169, // @[:@6.4]
  input  [3:0]  io_in_170, // @[:@6.4]
  input  [3:0]  io_in_171, // @[:@6.4]
  input  [3:0]  io_in_172, // @[:@6.4]
  input  [3:0]  io_in_173, // @[:@6.4]
  input  [3:0]  io_in_174, // @[:@6.4]
  input  [3:0]  io_in_175, // @[:@6.4]
  input  [3:0]  io_in_176, // @[:@6.4]
  input  [3:0]  io_in_177, // @[:@6.4]
  input  [3:0]  io_in_178, // @[:@6.4]
  input  [3:0]  io_in_179, // @[:@6.4]
  input  [3:0]  io_in_180, // @[:@6.4]
  input  [3:0]  io_in_181, // @[:@6.4]
  input  [3:0]  io_in_182, // @[:@6.4]
  input  [3:0]  io_in_183, // @[:@6.4]
  input  [3:0]  io_in_184, // @[:@6.4]
  input  [3:0]  io_in_185, // @[:@6.4]
  input  [3:0]  io_in_186, // @[:@6.4]
  input  [3:0]  io_in_187, // @[:@6.4]
  input  [3:0]  io_in_188, // @[:@6.4]
  input  [3:0]  io_in_189, // @[:@6.4]
  input  [3:0]  io_in_190, // @[:@6.4]
  input  [3:0]  io_in_191, // @[:@6.4]
  input  [3:0]  io_in_192, // @[:@6.4]
  input  [3:0]  io_in_193, // @[:@6.4]
  input  [3:0]  io_in_194, // @[:@6.4]
  input  [3:0]  io_in_195, // @[:@6.4]
  input  [3:0]  io_in_196, // @[:@6.4]
  input  [3:0]  io_in_197, // @[:@6.4]
  input  [3:0]  io_in_198, // @[:@6.4]
  input  [3:0]  io_in_199, // @[:@6.4]
  input  [3:0]  io_in_200, // @[:@6.4]
  input  [3:0]  io_in_201, // @[:@6.4]
  input  [3:0]  io_in_202, // @[:@6.4]
  input  [3:0]  io_in_203, // @[:@6.4]
  input  [3:0]  io_in_204, // @[:@6.4]
  input  [3:0]  io_in_205, // @[:@6.4]
  input  [3:0]  io_in_206, // @[:@6.4]
  input  [3:0]  io_in_207, // @[:@6.4]
  input  [3:0]  io_in_208, // @[:@6.4]
  input  [3:0]  io_in_209, // @[:@6.4]
  input  [3:0]  io_in_210, // @[:@6.4]
  input  [3:0]  io_in_211, // @[:@6.4]
  input  [3:0]  io_in_212, // @[:@6.4]
  input  [3:0]  io_in_213, // @[:@6.4]
  input  [3:0]  io_in_214, // @[:@6.4]
  input  [3:0]  io_in_215, // @[:@6.4]
  input  [3:0]  io_in_216, // @[:@6.4]
  input  [3:0]  io_in_217, // @[:@6.4]
  input  [3:0]  io_in_218, // @[:@6.4]
  input  [3:0]  io_in_219, // @[:@6.4]
  input  [3:0]  io_in_220, // @[:@6.4]
  input  [3:0]  io_in_221, // @[:@6.4]
  input  [3:0]  io_in_222, // @[:@6.4]
  input  [3:0]  io_in_223, // @[:@6.4]
  input  [3:0]  io_in_224, // @[:@6.4]
  input  [3:0]  io_in_225, // @[:@6.4]
  input  [3:0]  io_in_226, // @[:@6.4]
  input  [3:0]  io_in_227, // @[:@6.4]
  input  [3:0]  io_in_228, // @[:@6.4]
  input  [3:0]  io_in_229, // @[:@6.4]
  input  [3:0]  io_in_230, // @[:@6.4]
  input  [3:0]  io_in_231, // @[:@6.4]
  input  [3:0]  io_in_232, // @[:@6.4]
  input  [3:0]  io_in_233, // @[:@6.4]
  input  [3:0]  io_in_234, // @[:@6.4]
  input  [3:0]  io_in_235, // @[:@6.4]
  input  [3:0]  io_in_236, // @[:@6.4]
  input  [3:0]  io_in_237, // @[:@6.4]
  input  [3:0]  io_in_238, // @[:@6.4]
  input  [3:0]  io_in_239, // @[:@6.4]
  input  [3:0]  io_in_240, // @[:@6.4]
  input  [3:0]  io_in_241, // @[:@6.4]
  input  [3:0]  io_in_242, // @[:@6.4]
  input  [3:0]  io_in_243, // @[:@6.4]
  input  [3:0]  io_in_244, // @[:@6.4]
  input  [3:0]  io_in_245, // @[:@6.4]
  input  [3:0]  io_in_246, // @[:@6.4]
  input  [3:0]  io_in_247, // @[:@6.4]
  input  [3:0]  io_in_248, // @[:@6.4]
  input  [3:0]  io_in_249, // @[:@6.4]
  input  [3:0]  io_in_250, // @[:@6.4]
  input  [3:0]  io_in_251, // @[:@6.4]
  input  [3:0]  io_in_252, // @[:@6.4]
  input  [3:0]  io_in_253, // @[:@6.4]
  input  [3:0]  io_in_254, // @[:@6.4]
  input  [3:0]  io_in_255, // @[:@6.4]
  input  [3:0]  io_in_256, // @[:@6.4]
  input  [3:0]  io_in_257, // @[:@6.4]
  input  [3:0]  io_in_258, // @[:@6.4]
  input  [3:0]  io_in_259, // @[:@6.4]
  input  [3:0]  io_in_260, // @[:@6.4]
  input  [3:0]  io_in_261, // @[:@6.4]
  input  [3:0]  io_in_262, // @[:@6.4]
  input  [3:0]  io_in_263, // @[:@6.4]
  input  [3:0]  io_in_264, // @[:@6.4]
  input  [3:0]  io_in_265, // @[:@6.4]
  input  [3:0]  io_in_266, // @[:@6.4]
  input  [3:0]  io_in_267, // @[:@6.4]
  input  [3:0]  io_in_268, // @[:@6.4]
  input  [3:0]  io_in_269, // @[:@6.4]
  input  [3:0]  io_in_270, // @[:@6.4]
  input  [3:0]  io_in_271, // @[:@6.4]
  input  [3:0]  io_in_272, // @[:@6.4]
  input  [3:0]  io_in_273, // @[:@6.4]
  input  [3:0]  io_in_274, // @[:@6.4]
  input  [3:0]  io_in_275, // @[:@6.4]
  input  [3:0]  io_in_276, // @[:@6.4]
  input  [3:0]  io_in_277, // @[:@6.4]
  input  [3:0]  io_in_278, // @[:@6.4]
  input  [3:0]  io_in_279, // @[:@6.4]
  input  [3:0]  io_in_280, // @[:@6.4]
  input  [3:0]  io_in_281, // @[:@6.4]
  input  [3:0]  io_in_282, // @[:@6.4]
  input  [3:0]  io_in_283, // @[:@6.4]
  input  [3:0]  io_in_284, // @[:@6.4]
  input  [3:0]  io_in_285, // @[:@6.4]
  input  [3:0]  io_in_286, // @[:@6.4]
  input  [3:0]  io_in_287, // @[:@6.4]
  input  [3:0]  io_in_288, // @[:@6.4]
  input  [3:0]  io_in_289, // @[:@6.4]
  input  [3:0]  io_in_290, // @[:@6.4]
  input  [3:0]  io_in_291, // @[:@6.4]
  input  [3:0]  io_in_292, // @[:@6.4]
  input  [3:0]  io_in_293, // @[:@6.4]
  input  [3:0]  io_in_294, // @[:@6.4]
  input  [3:0]  io_in_295, // @[:@6.4]
  input  [3:0]  io_in_296, // @[:@6.4]
  input  [3:0]  io_in_297, // @[:@6.4]
  input  [3:0]  io_in_298, // @[:@6.4]
  input  [3:0]  io_in_299, // @[:@6.4]
  input  [3:0]  io_in_300, // @[:@6.4]
  input  [3:0]  io_in_301, // @[:@6.4]
  input  [3:0]  io_in_302, // @[:@6.4]
  input  [3:0]  io_in_303, // @[:@6.4]
  input  [3:0]  io_in_304, // @[:@6.4]
  input  [3:0]  io_in_305, // @[:@6.4]
  input  [3:0]  io_in_306, // @[:@6.4]
  input  [3:0]  io_in_307, // @[:@6.4]
  input  [3:0]  io_in_308, // @[:@6.4]
  input  [3:0]  io_in_309, // @[:@6.4]
  input  [3:0]  io_in_310, // @[:@6.4]
  input  [3:0]  io_in_311, // @[:@6.4]
  input  [3:0]  io_in_312, // @[:@6.4]
  input  [3:0]  io_in_313, // @[:@6.4]
  input  [3:0]  io_in_314, // @[:@6.4]
  input  [3:0]  io_in_315, // @[:@6.4]
  input  [3:0]  io_in_316, // @[:@6.4]
  input  [3:0]  io_in_317, // @[:@6.4]
  input  [3:0]  io_in_318, // @[:@6.4]
  input  [3:0]  io_in_319, // @[:@6.4]
  input  [3:0]  io_in_320, // @[:@6.4]
  input  [3:0]  io_in_321, // @[:@6.4]
  input  [3:0]  io_in_322, // @[:@6.4]
  input  [3:0]  io_in_323, // @[:@6.4]
  input  [3:0]  io_in_324, // @[:@6.4]
  input  [3:0]  io_in_325, // @[:@6.4]
  input  [3:0]  io_in_326, // @[:@6.4]
  input  [3:0]  io_in_327, // @[:@6.4]
  input  [3:0]  io_in_328, // @[:@6.4]
  input  [3:0]  io_in_329, // @[:@6.4]
  input  [3:0]  io_in_330, // @[:@6.4]
  input  [3:0]  io_in_331, // @[:@6.4]
  input  [3:0]  io_in_332, // @[:@6.4]
  input  [3:0]  io_in_333, // @[:@6.4]
  input  [3:0]  io_in_334, // @[:@6.4]
  input  [3:0]  io_in_335, // @[:@6.4]
  input  [3:0]  io_in_336, // @[:@6.4]
  input  [3:0]  io_in_337, // @[:@6.4]
  input  [3:0]  io_in_338, // @[:@6.4]
  input  [3:0]  io_in_339, // @[:@6.4]
  input  [3:0]  io_in_340, // @[:@6.4]
  input  [3:0]  io_in_341, // @[:@6.4]
  input  [3:0]  io_in_342, // @[:@6.4]
  input  [3:0]  io_in_343, // @[:@6.4]
  input  [3:0]  io_in_344, // @[:@6.4]
  input  [3:0]  io_in_345, // @[:@6.4]
  input  [3:0]  io_in_346, // @[:@6.4]
  input  [3:0]  io_in_347, // @[:@6.4]
  input  [3:0]  io_in_348, // @[:@6.4]
  input  [3:0]  io_in_349, // @[:@6.4]
  input  [3:0]  io_in_350, // @[:@6.4]
  input  [3:0]  io_in_351, // @[:@6.4]
  input  [3:0]  io_in_352, // @[:@6.4]
  input  [3:0]  io_in_353, // @[:@6.4]
  input  [3:0]  io_in_354, // @[:@6.4]
  input  [3:0]  io_in_355, // @[:@6.4]
  input  [3:0]  io_in_356, // @[:@6.4]
  input  [3:0]  io_in_357, // @[:@6.4]
  input  [3:0]  io_in_358, // @[:@6.4]
  input  [3:0]  io_in_359, // @[:@6.4]
  input  [3:0]  io_in_360, // @[:@6.4]
  input  [3:0]  io_in_361, // @[:@6.4]
  input  [3:0]  io_in_362, // @[:@6.4]
  input  [3:0]  io_in_363, // @[:@6.4]
  input  [3:0]  io_in_364, // @[:@6.4]
  input  [3:0]  io_in_365, // @[:@6.4]
  input  [3:0]  io_in_366, // @[:@6.4]
  input  [3:0]  io_in_367, // @[:@6.4]
  input  [3:0]  io_in_368, // @[:@6.4]
  input  [3:0]  io_in_369, // @[:@6.4]
  input  [3:0]  io_in_370, // @[:@6.4]
  input  [3:0]  io_in_371, // @[:@6.4]
  input  [3:0]  io_in_372, // @[:@6.4]
  input  [3:0]  io_in_373, // @[:@6.4]
  input  [3:0]  io_in_374, // @[:@6.4]
  input  [3:0]  io_in_375, // @[:@6.4]
  input  [3:0]  io_in_376, // @[:@6.4]
  input  [3:0]  io_in_377, // @[:@6.4]
  input  [3:0]  io_in_378, // @[:@6.4]
  input  [3:0]  io_in_379, // @[:@6.4]
  input  [3:0]  io_in_380, // @[:@6.4]
  input  [3:0]  io_in_381, // @[:@6.4]
  input  [3:0]  io_in_382, // @[:@6.4]
  input  [3:0]  io_in_383, // @[:@6.4]
  input  [3:0]  io_in_384, // @[:@6.4]
  input  [3:0]  io_in_385, // @[:@6.4]
  input  [3:0]  io_in_386, // @[:@6.4]
  input  [3:0]  io_in_387, // @[:@6.4]
  input  [3:0]  io_in_388, // @[:@6.4]
  input  [3:0]  io_in_389, // @[:@6.4]
  input  [3:0]  io_in_390, // @[:@6.4]
  input  [3:0]  io_in_391, // @[:@6.4]
  input  [3:0]  io_in_392, // @[:@6.4]
  input  [3:0]  io_in_393, // @[:@6.4]
  input  [3:0]  io_in_394, // @[:@6.4]
  input  [3:0]  io_in_395, // @[:@6.4]
  input  [3:0]  io_in_396, // @[:@6.4]
  input  [3:0]  io_in_397, // @[:@6.4]
  input  [3:0]  io_in_398, // @[:@6.4]
  input  [3:0]  io_in_399, // @[:@6.4]
  input  [3:0]  io_in_400, // @[:@6.4]
  input  [3:0]  io_in_401, // @[:@6.4]
  input  [3:0]  io_in_402, // @[:@6.4]
  input  [3:0]  io_in_403, // @[:@6.4]
  input  [3:0]  io_in_404, // @[:@6.4]
  input  [3:0]  io_in_405, // @[:@6.4]
  input  [3:0]  io_in_406, // @[:@6.4]
  input  [3:0]  io_in_407, // @[:@6.4]
  input  [3:0]  io_in_408, // @[:@6.4]
  input  [3:0]  io_in_409, // @[:@6.4]
  input  [3:0]  io_in_410, // @[:@6.4]
  input  [3:0]  io_in_411, // @[:@6.4]
  input  [3:0]  io_in_412, // @[:@6.4]
  input  [3:0]  io_in_413, // @[:@6.4]
  input  [3:0]  io_in_414, // @[:@6.4]
  input  [3:0]  io_in_415, // @[:@6.4]
  input  [3:0]  io_in_416, // @[:@6.4]
  input  [3:0]  io_in_417, // @[:@6.4]
  input  [3:0]  io_in_418, // @[:@6.4]
  input  [3:0]  io_in_419, // @[:@6.4]
  input  [3:0]  io_in_420, // @[:@6.4]
  input  [3:0]  io_in_421, // @[:@6.4]
  input  [3:0]  io_in_422, // @[:@6.4]
  input  [3:0]  io_in_423, // @[:@6.4]
  input  [3:0]  io_in_424, // @[:@6.4]
  input  [3:0]  io_in_425, // @[:@6.4]
  input  [3:0]  io_in_426, // @[:@6.4]
  input  [3:0]  io_in_427, // @[:@6.4]
  input  [3:0]  io_in_428, // @[:@6.4]
  input  [3:0]  io_in_429, // @[:@6.4]
  input  [3:0]  io_in_430, // @[:@6.4]
  input  [3:0]  io_in_431, // @[:@6.4]
  input  [3:0]  io_in_432, // @[:@6.4]
  input  [3:0]  io_in_433, // @[:@6.4]
  input  [3:0]  io_in_434, // @[:@6.4]
  input  [3:0]  io_in_435, // @[:@6.4]
  input  [3:0]  io_in_436, // @[:@6.4]
  input  [3:0]  io_in_437, // @[:@6.4]
  input  [3:0]  io_in_438, // @[:@6.4]
  input  [3:0]  io_in_439, // @[:@6.4]
  input  [3:0]  io_in_440, // @[:@6.4]
  input  [3:0]  io_in_441, // @[:@6.4]
  input  [3:0]  io_in_442, // @[:@6.4]
  input  [3:0]  io_in_443, // @[:@6.4]
  input  [3:0]  io_in_444, // @[:@6.4]
  input  [3:0]  io_in_445, // @[:@6.4]
  input  [3:0]  io_in_446, // @[:@6.4]
  input  [3:0]  io_in_447, // @[:@6.4]
  input  [3:0]  io_in_448, // @[:@6.4]
  input  [3:0]  io_in_449, // @[:@6.4]
  input  [3:0]  io_in_450, // @[:@6.4]
  input  [3:0]  io_in_451, // @[:@6.4]
  input  [3:0]  io_in_452, // @[:@6.4]
  input  [3:0]  io_in_453, // @[:@6.4]
  input  [3:0]  io_in_454, // @[:@6.4]
  input  [3:0]  io_in_455, // @[:@6.4]
  input  [3:0]  io_in_456, // @[:@6.4]
  input  [3:0]  io_in_457, // @[:@6.4]
  input  [3:0]  io_in_458, // @[:@6.4]
  input  [3:0]  io_in_459, // @[:@6.4]
  input  [3:0]  io_in_460, // @[:@6.4]
  input  [3:0]  io_in_461, // @[:@6.4]
  input  [3:0]  io_in_462, // @[:@6.4]
  input  [3:0]  io_in_463, // @[:@6.4]
  input  [3:0]  io_in_464, // @[:@6.4]
  input  [3:0]  io_in_465, // @[:@6.4]
  input  [3:0]  io_in_466, // @[:@6.4]
  input  [3:0]  io_in_467, // @[:@6.4]
  input  [3:0]  io_in_468, // @[:@6.4]
  input  [3:0]  io_in_469, // @[:@6.4]
  input  [3:0]  io_in_470, // @[:@6.4]
  input  [3:0]  io_in_471, // @[:@6.4]
  input  [3:0]  io_in_472, // @[:@6.4]
  input  [3:0]  io_in_473, // @[:@6.4]
  input  [3:0]  io_in_474, // @[:@6.4]
  input  [3:0]  io_in_475, // @[:@6.4]
  input  [3:0]  io_in_476, // @[:@6.4]
  input  [3:0]  io_in_477, // @[:@6.4]
  input  [3:0]  io_in_478, // @[:@6.4]
  input  [3:0]  io_in_479, // @[:@6.4]
  input  [3:0]  io_in_480, // @[:@6.4]
  input  [3:0]  io_in_481, // @[:@6.4]
  input  [3:0]  io_in_482, // @[:@6.4]
  input  [3:0]  io_in_483, // @[:@6.4]
  input  [3:0]  io_in_484, // @[:@6.4]
  input  [3:0]  io_in_485, // @[:@6.4]
  input  [3:0]  io_in_486, // @[:@6.4]
  input  [3:0]  io_in_487, // @[:@6.4]
  input  [3:0]  io_in_488, // @[:@6.4]
  input  [3:0]  io_in_489, // @[:@6.4]
  input  [3:0]  io_in_490, // @[:@6.4]
  input  [3:0]  io_in_491, // @[:@6.4]
  input  [3:0]  io_in_492, // @[:@6.4]
  input  [3:0]  io_in_493, // @[:@6.4]
  input  [3:0]  io_in_494, // @[:@6.4]
  input  [3:0]  io_in_495, // @[:@6.4]
  input  [3:0]  io_in_496, // @[:@6.4]
  input  [3:0]  io_in_497, // @[:@6.4]
  input  [3:0]  io_in_498, // @[:@6.4]
  input  [3:0]  io_in_499, // @[:@6.4]
  input  [3:0]  io_in_500, // @[:@6.4]
  input  [3:0]  io_in_501, // @[:@6.4]
  input  [3:0]  io_in_502, // @[:@6.4]
  input  [3:0]  io_in_503, // @[:@6.4]
  input  [3:0]  io_in_504, // @[:@6.4]
  input  [3:0]  io_in_505, // @[:@6.4]
  input  [3:0]  io_in_506, // @[:@6.4]
  input  [3:0]  io_in_507, // @[:@6.4]
  input  [3:0]  io_in_508, // @[:@6.4]
  input  [3:0]  io_in_509, // @[:@6.4]
  input  [3:0]  io_in_510, // @[:@6.4]
  input  [3:0]  io_in_511, // @[:@6.4]
  input  [3:0]  io_in_512, // @[:@6.4]
  input  [3:0]  io_in_513, // @[:@6.4]
  input  [3:0]  io_in_514, // @[:@6.4]
  input  [3:0]  io_in_515, // @[:@6.4]
  input  [3:0]  io_in_516, // @[:@6.4]
  input  [3:0]  io_in_517, // @[:@6.4]
  input  [3:0]  io_in_518, // @[:@6.4]
  input  [3:0]  io_in_519, // @[:@6.4]
  input  [3:0]  io_in_520, // @[:@6.4]
  input  [3:0]  io_in_521, // @[:@6.4]
  input  [3:0]  io_in_522, // @[:@6.4]
  input  [3:0]  io_in_523, // @[:@6.4]
  input  [3:0]  io_in_524, // @[:@6.4]
  input  [3:0]  io_in_525, // @[:@6.4]
  input  [3:0]  io_in_526, // @[:@6.4]
  input  [3:0]  io_in_527, // @[:@6.4]
  input  [3:0]  io_in_528, // @[:@6.4]
  input  [3:0]  io_in_529, // @[:@6.4]
  input  [3:0]  io_in_530, // @[:@6.4]
  input  [3:0]  io_in_531, // @[:@6.4]
  input  [3:0]  io_in_532, // @[:@6.4]
  input  [3:0]  io_in_533, // @[:@6.4]
  input  [3:0]  io_in_534, // @[:@6.4]
  input  [3:0]  io_in_535, // @[:@6.4]
  input  [3:0]  io_in_536, // @[:@6.4]
  input  [3:0]  io_in_537, // @[:@6.4]
  input  [3:0]  io_in_538, // @[:@6.4]
  input  [3:0]  io_in_539, // @[:@6.4]
  input  [3:0]  io_in_540, // @[:@6.4]
  input  [3:0]  io_in_541, // @[:@6.4]
  input  [3:0]  io_in_542, // @[:@6.4]
  input  [3:0]  io_in_543, // @[:@6.4]
  input  [3:0]  io_in_544, // @[:@6.4]
  input  [3:0]  io_in_545, // @[:@6.4]
  input  [3:0]  io_in_546, // @[:@6.4]
  input  [3:0]  io_in_547, // @[:@6.4]
  input  [3:0]  io_in_548, // @[:@6.4]
  input  [3:0]  io_in_549, // @[:@6.4]
  input  [3:0]  io_in_550, // @[:@6.4]
  input  [3:0]  io_in_551, // @[:@6.4]
  input  [3:0]  io_in_552, // @[:@6.4]
  input  [3:0]  io_in_553, // @[:@6.4]
  input  [3:0]  io_in_554, // @[:@6.4]
  input  [3:0]  io_in_555, // @[:@6.4]
  input  [3:0]  io_in_556, // @[:@6.4]
  input  [3:0]  io_in_557, // @[:@6.4]
  input  [3:0]  io_in_558, // @[:@6.4]
  input  [3:0]  io_in_559, // @[:@6.4]
  input  [3:0]  io_in_561, // @[:@6.4]
  input  [3:0]  io_in_562, // @[:@6.4]
  input  [3:0]  io_in_563, // @[:@6.4]
  input  [3:0]  io_in_564, // @[:@6.4]
  input  [3:0]  io_in_565, // @[:@6.4]
  input  [3:0]  io_in_566, // @[:@6.4]
  input  [3:0]  io_in_567, // @[:@6.4]
  input  [3:0]  io_in_568, // @[:@6.4]
  input  [3:0]  io_in_569, // @[:@6.4]
  input  [3:0]  io_in_570, // @[:@6.4]
  input  [3:0]  io_in_571, // @[:@6.4]
  input  [3:0]  io_in_572, // @[:@6.4]
  input  [3:0]  io_in_573, // @[:@6.4]
  input  [3:0]  io_in_574, // @[:@6.4]
  input  [3:0]  io_in_575, // @[:@6.4]
  input  [3:0]  io_in_576, // @[:@6.4]
  input  [3:0]  io_in_577, // @[:@6.4]
  input  [3:0]  io_in_578, // @[:@6.4]
  input  [3:0]  io_in_579, // @[:@6.4]
  input  [3:0]  io_in_580, // @[:@6.4]
  input  [3:0]  io_in_581, // @[:@6.4]
  input  [3:0]  io_in_582, // @[:@6.4]
  input  [3:0]  io_in_583, // @[:@6.4]
  input  [3:0]  io_in_584, // @[:@6.4]
  input  [3:0]  io_in_585, // @[:@6.4]
  input  [3:0]  io_in_586, // @[:@6.4]
  input  [3:0]  io_in_587, // @[:@6.4]
  input  [3:0]  io_in_588, // @[:@6.4]
  input  [3:0]  io_in_589, // @[:@6.4]
  input  [3:0]  io_in_590, // @[:@6.4]
  input  [3:0]  io_in_591, // @[:@6.4]
  input  [3:0]  io_in_592, // @[:@6.4]
  input  [3:0]  io_in_593, // @[:@6.4]
  input  [3:0]  io_in_594, // @[:@6.4]
  input  [3:0]  io_in_595, // @[:@6.4]
  input  [3:0]  io_in_596, // @[:@6.4]
  input  [3:0]  io_in_597, // @[:@6.4]
  input  [3:0]  io_in_598, // @[:@6.4]
  input  [3:0]  io_in_599, // @[:@6.4]
  input  [3:0]  io_in_600, // @[:@6.4]
  input  [3:0]  io_in_601, // @[:@6.4]
  input  [3:0]  io_in_602, // @[:@6.4]
  input  [3:0]  io_in_603, // @[:@6.4]
  input  [3:0]  io_in_604, // @[:@6.4]
  input  [3:0]  io_in_605, // @[:@6.4]
  input  [3:0]  io_in_606, // @[:@6.4]
  input  [3:0]  io_in_607, // @[:@6.4]
  input  [3:0]  io_in_608, // @[:@6.4]
  input  [3:0]  io_in_609, // @[:@6.4]
  input  [3:0]  io_in_610, // @[:@6.4]
  input  [3:0]  io_in_611, // @[:@6.4]
  input  [3:0]  io_in_612, // @[:@6.4]
  input  [3:0]  io_in_613, // @[:@6.4]
  input  [3:0]  io_in_614, // @[:@6.4]
  input  [3:0]  io_in_615, // @[:@6.4]
  input  [3:0]  io_in_616, // @[:@6.4]
  input  [3:0]  io_in_617, // @[:@6.4]
  input  [3:0]  io_in_618, // @[:@6.4]
  input  [3:0]  io_in_619, // @[:@6.4]
  input  [3:0]  io_in_620, // @[:@6.4]
  input  [3:0]  io_in_621, // @[:@6.4]
  input  [3:0]  io_in_622, // @[:@6.4]
  input  [3:0]  io_in_623, // @[:@6.4]
  input  [3:0]  io_in_624, // @[:@6.4]
  input  [3:0]  io_in_625, // @[:@6.4]
  input  [3:0]  io_in_626, // @[:@6.4]
  input  [3:0]  io_in_627, // @[:@6.4]
  input  [3:0]  io_in_628, // @[:@6.4]
  input  [3:0]  io_in_629, // @[:@6.4]
  input  [3:0]  io_in_630, // @[:@6.4]
  input  [3:0]  io_in_631, // @[:@6.4]
  input  [3:0]  io_in_632, // @[:@6.4]
  input  [3:0]  io_in_633, // @[:@6.4]
  input  [3:0]  io_in_634, // @[:@6.4]
  input  [3:0]  io_in_635, // @[:@6.4]
  input  [3:0]  io_in_636, // @[:@6.4]
  input  [3:0]  io_in_637, // @[:@6.4]
  input  [3:0]  io_in_638, // @[:@6.4]
  input  [3:0]  io_in_639, // @[:@6.4]
  input  [3:0]  io_in_640, // @[:@6.4]
  input  [3:0]  io_in_641, // @[:@6.4]
  input  [3:0]  io_in_642, // @[:@6.4]
  input  [3:0]  io_in_646, // @[:@6.4]
  input  [3:0]  io_in_647, // @[:@6.4]
  input  [3:0]  io_in_648, // @[:@6.4]
  input  [3:0]  io_in_649, // @[:@6.4]
  input  [3:0]  io_in_650, // @[:@6.4]
  input  [3:0]  io_in_651, // @[:@6.4]
  input  [3:0]  io_in_652, // @[:@6.4]
  input  [3:0]  io_in_653, // @[:@6.4]
  input  [3:0]  io_in_654, // @[:@6.4]
  input  [3:0]  io_in_655, // @[:@6.4]
  input  [3:0]  io_in_656, // @[:@6.4]
  input  [3:0]  io_in_657, // @[:@6.4]
  input  [3:0]  io_in_658, // @[:@6.4]
  input  [3:0]  io_in_659, // @[:@6.4]
  input  [3:0]  io_in_660, // @[:@6.4]
  input  [3:0]  io_in_661, // @[:@6.4]
  input  [3:0]  io_in_662, // @[:@6.4]
  input  [3:0]  io_in_663, // @[:@6.4]
  input  [3:0]  io_in_664, // @[:@6.4]
  input  [3:0]  io_in_665, // @[:@6.4]
  input  [3:0]  io_in_666, // @[:@6.4]
  input  [3:0]  io_in_667, // @[:@6.4]
  input  [3:0]  io_in_668, // @[:@6.4]
  input  [3:0]  io_in_669, // @[:@6.4]
  input  [3:0]  io_in_670, // @[:@6.4]
  input  [3:0]  io_in_673, // @[:@6.4]
  input  [3:0]  io_in_674, // @[:@6.4]
  input  [3:0]  io_in_675, // @[:@6.4]
  input  [3:0]  io_in_676, // @[:@6.4]
  input  [3:0]  io_in_677, // @[:@6.4]
  input  [3:0]  io_in_678, // @[:@6.4]
  input  [3:0]  io_in_679, // @[:@6.4]
  input  [3:0]  io_in_680, // @[:@6.4]
  input  [3:0]  io_in_681, // @[:@6.4]
  input  [3:0]  io_in_682, // @[:@6.4]
  input  [3:0]  io_in_683, // @[:@6.4]
  input  [3:0]  io_in_684, // @[:@6.4]
  input  [3:0]  io_in_685, // @[:@6.4]
  input  [3:0]  io_in_686, // @[:@6.4]
  input  [3:0]  io_in_687, // @[:@6.4]
  input  [3:0]  io_in_688, // @[:@6.4]
  input  [3:0]  io_in_689, // @[:@6.4]
  input  [3:0]  io_in_690, // @[:@6.4]
  input  [3:0]  io_in_691, // @[:@6.4]
  input  [3:0]  io_in_692, // @[:@6.4]
  input  [3:0]  io_in_693, // @[:@6.4]
  input  [3:0]  io_in_694, // @[:@6.4]
  input  [3:0]  io_in_695, // @[:@6.4]
  input  [3:0]  io_in_696, // @[:@6.4]
  input  [3:0]  io_in_697, // @[:@6.4]
  input  [3:0]  io_in_698, // @[:@6.4]
  input  [3:0]  io_in_699, // @[:@6.4]
  input  [3:0]  io_in_702, // @[:@6.4]
  input  [3:0]  io_in_703, // @[:@6.4]
  input  [3:0]  io_in_704, // @[:@6.4]
  input  [3:0]  io_in_705, // @[:@6.4]
  input  [3:0]  io_in_706, // @[:@6.4]
  input  [3:0]  io_in_707, // @[:@6.4]
  input  [3:0]  io_in_708, // @[:@6.4]
  input  [3:0]  io_in_709, // @[:@6.4]
  input  [3:0]  io_in_710, // @[:@6.4]
  input  [3:0]  io_in_711, // @[:@6.4]
  input  [3:0]  io_in_712, // @[:@6.4]
  input  [3:0]  io_in_713, // @[:@6.4]
  input  [3:0]  io_in_714, // @[:@6.4]
  input  [3:0]  io_in_715, // @[:@6.4]
  input  [3:0]  io_in_716, // @[:@6.4]
  input  [3:0]  io_in_717, // @[:@6.4]
  input  [3:0]  io_in_718, // @[:@6.4]
  input  [3:0]  io_in_719, // @[:@6.4]
  input  [3:0]  io_in_720, // @[:@6.4]
  input  [3:0]  io_in_721, // @[:@6.4]
  input  [3:0]  io_in_722, // @[:@6.4]
  input  [3:0]  io_in_723, // @[:@6.4]
  input  [3:0]  io_in_724, // @[:@6.4]
  input  [3:0]  io_in_725, // @[:@6.4]
  input  [3:0]  io_in_726, // @[:@6.4]
  input  [3:0]  io_in_728, // @[:@6.4]
  input  [3:0]  io_in_729, // @[:@6.4]
  input  [3:0]  io_in_731, // @[:@6.4]
  input  [3:0]  io_in_732, // @[:@6.4]
  input  [3:0]  io_in_733, // @[:@6.4]
  input  [3:0]  io_in_734, // @[:@6.4]
  input  [3:0]  io_in_735, // @[:@6.4]
  input  [3:0]  io_in_736, // @[:@6.4]
  input  [3:0]  io_in_737, // @[:@6.4]
  input  [3:0]  io_in_738, // @[:@6.4]
  input  [3:0]  io_in_739, // @[:@6.4]
  input  [3:0]  io_in_740, // @[:@6.4]
  input  [3:0]  io_in_741, // @[:@6.4]
  input  [3:0]  io_in_742, // @[:@6.4]
  input  [3:0]  io_in_743, // @[:@6.4]
  input  [3:0]  io_in_744, // @[:@6.4]
  input  [3:0]  io_in_745, // @[:@6.4]
  input  [3:0]  io_in_746, // @[:@6.4]
  input  [3:0]  io_in_747, // @[:@6.4]
  input  [3:0]  io_in_748, // @[:@6.4]
  input  [3:0]  io_in_749, // @[:@6.4]
  input  [3:0]  io_in_750, // @[:@6.4]
  input  [3:0]  io_in_751, // @[:@6.4]
  input  [3:0]  io_in_752, // @[:@6.4]
  input  [3:0]  io_in_753, // @[:@6.4]
  input  [3:0]  io_in_756, // @[:@6.4]
  input  [3:0]  io_in_758, // @[:@6.4]
  input  [3:0]  io_in_760, // @[:@6.4]
  input  [3:0]  io_in_761, // @[:@6.4]
  input  [3:0]  io_in_762, // @[:@6.4]
  input  [3:0]  io_in_763, // @[:@6.4]
  input  [3:0]  io_in_764, // @[:@6.4]
  input  [3:0]  io_in_765, // @[:@6.4]
  input  [3:0]  io_in_766, // @[:@6.4]
  input  [3:0]  io_in_767, // @[:@6.4]
  input  [3:0]  io_in_768, // @[:@6.4]
  input  [3:0]  io_in_769, // @[:@6.4]
  input  [3:0]  io_in_770, // @[:@6.4]
  input  [3:0]  io_in_771, // @[:@6.4]
  input  [3:0]  io_in_772, // @[:@6.4]
  input  [3:0]  io_in_773, // @[:@6.4]
  input  [3:0]  io_in_774, // @[:@6.4]
  input  [3:0]  io_in_775, // @[:@6.4]
  input  [3:0]  io_in_776, // @[:@6.4]
  input  [3:0]  io_in_777, // @[:@6.4]
  input  [3:0]  io_in_778, // @[:@6.4]
  input  [3:0]  io_in_779, // @[:@6.4]
  input  [3:0]  io_in_780, // @[:@6.4]
  output [13:0] io_out_0, // @[:@6.4]
  output [13:0] io_out_1, // @[:@6.4]
  output [13:0] io_out_2, // @[:@6.4]
  output [13:0] io_out_3, // @[:@6.4]
  output [13:0] io_out_4, // @[:@6.4]
  output [13:0] io_out_5, // @[:@6.4]
  output [13:0] io_out_6, // @[:@6.4]
  output [13:0] io_out_7, // @[:@6.4]
  output [13:0] io_out_8, // @[:@6.4]
  output [13:0] io_out_9, // @[:@6.4]
  output [13:0] io_out_10, // @[:@6.4]
  output [13:0] io_out_11, // @[:@6.4]
  output [13:0] io_out_12, // @[:@6.4]
  output [13:0] io_out_13, // @[:@6.4]
  output [13:0] io_out_14, // @[:@6.4]
  output [13:0] io_out_15 // @[:@6.4]
);
  wire [5:0] _T_54199; // @[Modules.scala 150:74:@9.4]
  wire [5:0] _T_54201; // @[Modules.scala 151:80:@10.4]
  wire [6:0] _T_54202; // @[Modules.scala 150:103:@11.4]
  wire [5:0] _T_54203; // @[Modules.scala 150:103:@12.4]
  wire [5:0] _T_54204; // @[Modules.scala 150:103:@13.4]
  wire [5:0] _T_54206; // @[Modules.scala 150:74:@15.4]
  wire [5:0] _T_54208; // @[Modules.scala 151:80:@16.4]
  wire [6:0] _T_54209; // @[Modules.scala 150:103:@17.4]
  wire [5:0] _T_54210; // @[Modules.scala 150:103:@18.4]
  wire [5:0] _T_54211; // @[Modules.scala 150:103:@19.4]
  wire [4:0] _T_54213; // @[Modules.scala 150:74:@21.4]
  wire [5:0] _T_54215; // @[Modules.scala 151:80:@22.4]
  wire [5:0] _GEN_0; // @[Modules.scala 150:103:@23.4]
  wire [6:0] _T_54216; // @[Modules.scala 150:103:@23.4]
  wire [5:0] _T_54217; // @[Modules.scala 150:103:@24.4]
  wire [5:0] _T_54218; // @[Modules.scala 150:103:@25.4]
  wire [5:0] _T_54220; // @[Modules.scala 150:74:@27.4]
  wire [5:0] _T_54222; // @[Modules.scala 151:80:@28.4]
  wire [6:0] _T_54223; // @[Modules.scala 150:103:@29.4]
  wire [5:0] _T_54224; // @[Modules.scala 150:103:@30.4]
  wire [5:0] _T_54225; // @[Modules.scala 150:103:@31.4]
  wire [5:0] _T_54227; // @[Modules.scala 150:74:@33.4]
  wire [5:0] _T_54229; // @[Modules.scala 151:80:@34.4]
  wire [6:0] _T_54230; // @[Modules.scala 150:103:@35.4]
  wire [5:0] _T_54231; // @[Modules.scala 150:103:@36.4]
  wire [5:0] _T_54232; // @[Modules.scala 150:103:@37.4]
  wire [5:0] _T_54234; // @[Modules.scala 150:74:@39.4]
  wire [5:0] _T_54236; // @[Modules.scala 151:80:@40.4]
  wire [6:0] _T_54237; // @[Modules.scala 150:103:@41.4]
  wire [5:0] _T_54238; // @[Modules.scala 150:103:@42.4]
  wire [5:0] _T_54239; // @[Modules.scala 150:103:@43.4]
  wire [5:0] _T_54241; // @[Modules.scala 150:74:@45.4]
  wire [5:0] _T_54243; // @[Modules.scala 151:80:@46.4]
  wire [6:0] _T_54244; // @[Modules.scala 150:103:@47.4]
  wire [5:0] _T_54245; // @[Modules.scala 150:103:@48.4]
  wire [5:0] _T_54246; // @[Modules.scala 150:103:@49.4]
  wire [5:0] _T_54248; // @[Modules.scala 150:74:@51.4]
  wire [5:0] _T_54250; // @[Modules.scala 151:80:@52.4]
  wire [6:0] _T_54251; // @[Modules.scala 150:103:@53.4]
  wire [5:0] _T_54252; // @[Modules.scala 150:103:@54.4]
  wire [5:0] _T_54253; // @[Modules.scala 150:103:@55.4]
  wire [5:0] _T_54255; // @[Modules.scala 150:74:@57.4]
  wire [5:0] _T_54257; // @[Modules.scala 151:80:@58.4]
  wire [6:0] _T_54258; // @[Modules.scala 150:103:@59.4]
  wire [5:0] _T_54259; // @[Modules.scala 150:103:@60.4]
  wire [5:0] _T_54260; // @[Modules.scala 150:103:@61.4]
  wire [5:0] _T_54262; // @[Modules.scala 150:74:@63.4]
  wire [5:0] _T_54264; // @[Modules.scala 151:80:@64.4]
  wire [6:0] _T_54265; // @[Modules.scala 150:103:@65.4]
  wire [5:0] _T_54266; // @[Modules.scala 150:103:@66.4]
  wire [5:0] _T_54267; // @[Modules.scala 150:103:@67.4]
  wire [5:0] _T_54269; // @[Modules.scala 150:74:@69.4]
  wire [5:0] _T_54271; // @[Modules.scala 151:80:@70.4]
  wire [6:0] _T_54272; // @[Modules.scala 150:103:@71.4]
  wire [5:0] _T_54273; // @[Modules.scala 150:103:@72.4]
  wire [5:0] _T_54274; // @[Modules.scala 150:103:@73.4]
  wire [5:0] _T_54276; // @[Modules.scala 150:74:@75.4]
  wire [5:0] _T_54278; // @[Modules.scala 151:80:@76.4]
  wire [6:0] _T_54279; // @[Modules.scala 150:103:@77.4]
  wire [5:0] _T_54280; // @[Modules.scala 150:103:@78.4]
  wire [5:0] _T_54281; // @[Modules.scala 150:103:@79.4]
  wire [5:0] _T_54283; // @[Modules.scala 150:74:@81.4]
  wire [5:0] _T_54285; // @[Modules.scala 151:80:@82.4]
  wire [6:0] _T_54286; // @[Modules.scala 150:103:@83.4]
  wire [5:0] _T_54287; // @[Modules.scala 150:103:@84.4]
  wire [5:0] _T_54288; // @[Modules.scala 150:103:@85.4]
  wire [5:0] _T_54290; // @[Modules.scala 150:74:@87.4]
  wire [5:0] _T_54292; // @[Modules.scala 151:80:@88.4]
  wire [6:0] _T_54293; // @[Modules.scala 150:103:@89.4]
  wire [5:0] _T_54294; // @[Modules.scala 150:103:@90.4]
  wire [5:0] _T_54295; // @[Modules.scala 150:103:@91.4]
  wire [5:0] _T_54297; // @[Modules.scala 150:74:@93.4]
  wire [5:0] _T_54299; // @[Modules.scala 151:80:@94.4]
  wire [6:0] _T_54300; // @[Modules.scala 150:103:@95.4]
  wire [5:0] _T_54301; // @[Modules.scala 150:103:@96.4]
  wire [5:0] _T_54302; // @[Modules.scala 150:103:@97.4]
  wire [5:0] _T_54304; // @[Modules.scala 150:74:@99.4]
  wire [5:0] _T_54306; // @[Modules.scala 151:80:@100.4]
  wire [6:0] _T_54307; // @[Modules.scala 150:103:@101.4]
  wire [5:0] _T_54308; // @[Modules.scala 150:103:@102.4]
  wire [5:0] _T_54309; // @[Modules.scala 150:103:@103.4]
  wire [5:0] _T_54311; // @[Modules.scala 150:74:@105.4]
  wire [5:0] _T_54313; // @[Modules.scala 151:80:@106.4]
  wire [6:0] _T_54314; // @[Modules.scala 150:103:@107.4]
  wire [5:0] _T_54315; // @[Modules.scala 150:103:@108.4]
  wire [5:0] _T_54316; // @[Modules.scala 150:103:@109.4]
  wire [5:0] _T_54318; // @[Modules.scala 150:74:@111.4]
  wire [5:0] _T_54320; // @[Modules.scala 151:80:@112.4]
  wire [6:0] _T_54321; // @[Modules.scala 150:103:@113.4]
  wire [5:0] _T_54322; // @[Modules.scala 150:103:@114.4]
  wire [5:0] _T_54323; // @[Modules.scala 150:103:@115.4]
  wire [5:0] _T_54325; // @[Modules.scala 150:74:@117.4]
  wire [5:0] _T_54327; // @[Modules.scala 151:80:@118.4]
  wire [6:0] _T_54328; // @[Modules.scala 150:103:@119.4]
  wire [5:0] _T_54329; // @[Modules.scala 150:103:@120.4]
  wire [5:0] _T_54330; // @[Modules.scala 150:103:@121.4]
  wire [5:0] _T_54332; // @[Modules.scala 150:74:@123.4]
  wire [5:0] _T_54334; // @[Modules.scala 151:80:@124.4]
  wire [6:0] _T_54335; // @[Modules.scala 150:103:@125.4]
  wire [5:0] _T_54336; // @[Modules.scala 150:103:@126.4]
  wire [5:0] _T_54337; // @[Modules.scala 150:103:@127.4]
  wire [5:0] _T_54339; // @[Modules.scala 150:74:@129.4]
  wire [5:0] _T_54341; // @[Modules.scala 151:80:@130.4]
  wire [6:0] _T_54342; // @[Modules.scala 150:103:@131.4]
  wire [5:0] _T_54343; // @[Modules.scala 150:103:@132.4]
  wire [5:0] _T_54344; // @[Modules.scala 150:103:@133.4]
  wire [5:0] _T_54346; // @[Modules.scala 150:74:@135.4]
  wire [5:0] _T_54348; // @[Modules.scala 151:80:@136.4]
  wire [6:0] _T_54349; // @[Modules.scala 150:103:@137.4]
  wire [5:0] _T_54350; // @[Modules.scala 150:103:@138.4]
  wire [5:0] _T_54351; // @[Modules.scala 150:103:@139.4]
  wire [5:0] _T_54353; // @[Modules.scala 150:74:@141.4]
  wire [4:0] _T_54355; // @[Modules.scala 151:80:@142.4]
  wire [5:0] _GEN_1; // @[Modules.scala 150:103:@143.4]
  wire [6:0] _T_54356; // @[Modules.scala 150:103:@143.4]
  wire [5:0] _T_54357; // @[Modules.scala 150:103:@144.4]
  wire [5:0] _T_54358; // @[Modules.scala 150:103:@145.4]
  wire [5:0] _T_54360; // @[Modules.scala 150:74:@147.4]
  wire [5:0] _T_54362; // @[Modules.scala 151:80:@148.4]
  wire [6:0] _T_54363; // @[Modules.scala 150:103:@149.4]
  wire [5:0] _T_54364; // @[Modules.scala 150:103:@150.4]
  wire [5:0] _T_54365; // @[Modules.scala 150:103:@151.4]
  wire [5:0] _T_54367; // @[Modules.scala 150:74:@153.4]
  wire [5:0] _T_54369; // @[Modules.scala 151:80:@154.4]
  wire [6:0] _T_54370; // @[Modules.scala 150:103:@155.4]
  wire [5:0] _T_54371; // @[Modules.scala 150:103:@156.4]
  wire [5:0] _T_54372; // @[Modules.scala 150:103:@157.4]
  wire [5:0] _T_54374; // @[Modules.scala 150:74:@159.4]
  wire [5:0] _T_54376; // @[Modules.scala 151:80:@160.4]
  wire [6:0] _T_54377; // @[Modules.scala 150:103:@161.4]
  wire [5:0] _T_54378; // @[Modules.scala 150:103:@162.4]
  wire [5:0] _T_54379; // @[Modules.scala 150:103:@163.4]
  wire [5:0] _T_54381; // @[Modules.scala 150:74:@165.4]
  wire [5:0] _T_54383; // @[Modules.scala 151:80:@166.4]
  wire [6:0] _T_54384; // @[Modules.scala 150:103:@167.4]
  wire [5:0] _T_54385; // @[Modules.scala 150:103:@168.4]
  wire [5:0] _T_54386; // @[Modules.scala 150:103:@169.4]
  wire [5:0] _T_54388; // @[Modules.scala 150:74:@171.4]
  wire [5:0] _T_54390; // @[Modules.scala 151:80:@172.4]
  wire [6:0] _T_54391; // @[Modules.scala 150:103:@173.4]
  wire [5:0] _T_54392; // @[Modules.scala 150:103:@174.4]
  wire [5:0] _T_54393; // @[Modules.scala 150:103:@175.4]
  wire [5:0] _T_54395; // @[Modules.scala 150:74:@177.4]
  wire [5:0] _T_54397; // @[Modules.scala 151:80:@178.4]
  wire [6:0] _T_54398; // @[Modules.scala 150:103:@179.4]
  wire [5:0] _T_54399; // @[Modules.scala 150:103:@180.4]
  wire [5:0] _T_54400; // @[Modules.scala 150:103:@181.4]
  wire [5:0] _T_54402; // @[Modules.scala 150:74:@183.4]
  wire [5:0] _T_54404; // @[Modules.scala 151:80:@184.4]
  wire [6:0] _T_54405; // @[Modules.scala 150:103:@185.4]
  wire [5:0] _T_54406; // @[Modules.scala 150:103:@186.4]
  wire [5:0] _T_54407; // @[Modules.scala 150:103:@187.4]
  wire [5:0] _T_54409; // @[Modules.scala 150:74:@189.4]
  wire [5:0] _T_54411; // @[Modules.scala 151:80:@190.4]
  wire [6:0] _T_54412; // @[Modules.scala 150:103:@191.4]
  wire [5:0] _T_54413; // @[Modules.scala 150:103:@192.4]
  wire [5:0] _T_54414; // @[Modules.scala 150:103:@193.4]
  wire [5:0] _T_54416; // @[Modules.scala 150:74:@195.4]
  wire [5:0] _T_54418; // @[Modules.scala 151:80:@196.4]
  wire [6:0] _T_54419; // @[Modules.scala 150:103:@197.4]
  wire [5:0] _T_54420; // @[Modules.scala 150:103:@198.4]
  wire [5:0] _T_54421; // @[Modules.scala 150:103:@199.4]
  wire [5:0] _T_54423; // @[Modules.scala 150:74:@201.4]
  wire [5:0] _T_54425; // @[Modules.scala 151:80:@202.4]
  wire [6:0] _T_54426; // @[Modules.scala 150:103:@203.4]
  wire [5:0] _T_54427; // @[Modules.scala 150:103:@204.4]
  wire [5:0] _T_54428; // @[Modules.scala 150:103:@205.4]
  wire [5:0] _T_54430; // @[Modules.scala 150:74:@207.4]
  wire [5:0] _T_54432; // @[Modules.scala 151:80:@208.4]
  wire [6:0] _T_54433; // @[Modules.scala 150:103:@209.4]
  wire [5:0] _T_54434; // @[Modules.scala 150:103:@210.4]
  wire [5:0] _T_54435; // @[Modules.scala 150:103:@211.4]
  wire [5:0] _T_54437; // @[Modules.scala 150:74:@213.4]
  wire [4:0] _T_54439; // @[Modules.scala 151:80:@214.4]
  wire [5:0] _GEN_2; // @[Modules.scala 150:103:@215.4]
  wire [6:0] _T_54440; // @[Modules.scala 150:103:@215.4]
  wire [5:0] _T_54441; // @[Modules.scala 150:103:@216.4]
  wire [5:0] _T_54442; // @[Modules.scala 150:103:@217.4]
  wire [5:0] _T_54444; // @[Modules.scala 150:74:@219.4]
  wire [4:0] _T_54446; // @[Modules.scala 151:80:@220.4]
  wire [5:0] _GEN_3; // @[Modules.scala 150:103:@221.4]
  wire [6:0] _T_54447; // @[Modules.scala 150:103:@221.4]
  wire [5:0] _T_54448; // @[Modules.scala 150:103:@222.4]
  wire [5:0] _T_54449; // @[Modules.scala 150:103:@223.4]
  wire [5:0] _T_54451; // @[Modules.scala 150:74:@225.4]
  wire [4:0] _T_54453; // @[Modules.scala 151:80:@226.4]
  wire [5:0] _GEN_4; // @[Modules.scala 150:103:@227.4]
  wire [6:0] _T_54454; // @[Modules.scala 150:103:@227.4]
  wire [5:0] _T_54455; // @[Modules.scala 150:103:@228.4]
  wire [5:0] _T_54456; // @[Modules.scala 150:103:@229.4]
  wire [4:0] _T_54458; // @[Modules.scala 150:74:@231.4]
  wire [5:0] _T_54460; // @[Modules.scala 151:80:@232.4]
  wire [5:0] _GEN_5; // @[Modules.scala 150:103:@233.4]
  wire [6:0] _T_54461; // @[Modules.scala 150:103:@233.4]
  wire [5:0] _T_54462; // @[Modules.scala 150:103:@234.4]
  wire [5:0] _T_54463; // @[Modules.scala 150:103:@235.4]
  wire [5:0] _T_54465; // @[Modules.scala 150:74:@237.4]
  wire [5:0] _T_54467; // @[Modules.scala 151:80:@238.4]
  wire [6:0] _T_54468; // @[Modules.scala 150:103:@239.4]
  wire [5:0] _T_54469; // @[Modules.scala 150:103:@240.4]
  wire [5:0] _T_54470; // @[Modules.scala 150:103:@241.4]
  wire [5:0] _T_54472; // @[Modules.scala 150:74:@243.4]
  wire [5:0] _T_54474; // @[Modules.scala 151:80:@244.4]
  wire [6:0] _T_54475; // @[Modules.scala 150:103:@245.4]
  wire [5:0] _T_54476; // @[Modules.scala 150:103:@246.4]
  wire [5:0] _T_54477; // @[Modules.scala 150:103:@247.4]
  wire [5:0] _T_54479; // @[Modules.scala 150:74:@249.4]
  wire [5:0] _T_54481; // @[Modules.scala 151:80:@250.4]
  wire [6:0] _T_54482; // @[Modules.scala 150:103:@251.4]
  wire [5:0] _T_54483; // @[Modules.scala 150:103:@252.4]
  wire [5:0] _T_54484; // @[Modules.scala 150:103:@253.4]
  wire [5:0] _T_54486; // @[Modules.scala 150:74:@255.4]
  wire [5:0] _T_54488; // @[Modules.scala 151:80:@256.4]
  wire [6:0] _T_54489; // @[Modules.scala 150:103:@257.4]
  wire [5:0] _T_54490; // @[Modules.scala 150:103:@258.4]
  wire [5:0] _T_54491; // @[Modules.scala 150:103:@259.4]
  wire [5:0] _T_54493; // @[Modules.scala 150:74:@261.4]
  wire [5:0] _T_54495; // @[Modules.scala 151:80:@262.4]
  wire [6:0] _T_54496; // @[Modules.scala 150:103:@263.4]
  wire [5:0] _T_54497; // @[Modules.scala 150:103:@264.4]
  wire [5:0] _T_54498; // @[Modules.scala 150:103:@265.4]
  wire [5:0] _T_54500; // @[Modules.scala 150:74:@267.4]
  wire [5:0] _T_54502; // @[Modules.scala 151:80:@268.4]
  wire [6:0] _T_54503; // @[Modules.scala 150:103:@269.4]
  wire [5:0] _T_54504; // @[Modules.scala 150:103:@270.4]
  wire [5:0] _T_54505; // @[Modules.scala 150:103:@271.4]
  wire [4:0] _T_54507; // @[Modules.scala 150:74:@273.4]
  wire [4:0] _T_54509; // @[Modules.scala 151:80:@274.4]
  wire [5:0] _T_54510; // @[Modules.scala 150:103:@275.4]
  wire [4:0] _T_54511; // @[Modules.scala 150:103:@276.4]
  wire [4:0] _T_54512; // @[Modules.scala 150:103:@277.4]
  wire [4:0] _T_54514; // @[Modules.scala 150:74:@279.4]
  wire [5:0] _T_54516; // @[Modules.scala 151:80:@280.4]
  wire [5:0] _GEN_6; // @[Modules.scala 150:103:@281.4]
  wire [6:0] _T_54517; // @[Modules.scala 150:103:@281.4]
  wire [5:0] _T_54518; // @[Modules.scala 150:103:@282.4]
  wire [5:0] _T_54519; // @[Modules.scala 150:103:@283.4]
  wire [5:0] _T_54521; // @[Modules.scala 150:74:@285.4]
  wire [4:0] _T_54523; // @[Modules.scala 151:80:@286.4]
  wire [5:0] _GEN_7; // @[Modules.scala 150:103:@287.4]
  wire [6:0] _T_54524; // @[Modules.scala 150:103:@287.4]
  wire [5:0] _T_54525; // @[Modules.scala 150:103:@288.4]
  wire [5:0] _T_54526; // @[Modules.scala 150:103:@289.4]
  wire [4:0] _T_54528; // @[Modules.scala 150:74:@291.4]
  wire [5:0] _T_54530; // @[Modules.scala 151:80:@292.4]
  wire [5:0] _GEN_8; // @[Modules.scala 150:103:@293.4]
  wire [6:0] _T_54531; // @[Modules.scala 150:103:@293.4]
  wire [5:0] _T_54532; // @[Modules.scala 150:103:@294.4]
  wire [5:0] _T_54533; // @[Modules.scala 150:103:@295.4]
  wire [5:0] _T_54535; // @[Modules.scala 150:74:@297.4]
  wire [5:0] _T_54537; // @[Modules.scala 151:80:@298.4]
  wire [6:0] _T_54538; // @[Modules.scala 150:103:@299.4]
  wire [5:0] _T_54539; // @[Modules.scala 150:103:@300.4]
  wire [5:0] _T_54540; // @[Modules.scala 150:103:@301.4]
  wire [5:0] _T_54542; // @[Modules.scala 150:74:@303.4]
  wire [4:0] _T_54544; // @[Modules.scala 151:80:@304.4]
  wire [5:0] _GEN_9; // @[Modules.scala 150:103:@305.4]
  wire [6:0] _T_54545; // @[Modules.scala 150:103:@305.4]
  wire [5:0] _T_54546; // @[Modules.scala 150:103:@306.4]
  wire [5:0] _T_54547; // @[Modules.scala 150:103:@307.4]
  wire [4:0] _T_54549; // @[Modules.scala 150:74:@309.4]
  wire [4:0] _T_54551; // @[Modules.scala 151:80:@310.4]
  wire [5:0] _T_54552; // @[Modules.scala 150:103:@311.4]
  wire [4:0] _T_54553; // @[Modules.scala 150:103:@312.4]
  wire [4:0] _T_54554; // @[Modules.scala 150:103:@313.4]
  wire [5:0] _T_54556; // @[Modules.scala 150:74:@315.4]
  wire [4:0] _T_54558; // @[Modules.scala 151:80:@316.4]
  wire [5:0] _GEN_10; // @[Modules.scala 150:103:@317.4]
  wire [6:0] _T_54559; // @[Modules.scala 150:103:@317.4]
  wire [5:0] _T_54560; // @[Modules.scala 150:103:@318.4]
  wire [5:0] _T_54561; // @[Modules.scala 150:103:@319.4]
  wire [4:0] _T_54563; // @[Modules.scala 150:74:@321.4]
  wire [4:0] _T_54565; // @[Modules.scala 151:80:@322.4]
  wire [5:0] _T_54566; // @[Modules.scala 150:103:@323.4]
  wire [4:0] _T_54567; // @[Modules.scala 150:103:@324.4]
  wire [4:0] _T_54568; // @[Modules.scala 150:103:@325.4]
  wire [4:0] _T_54570; // @[Modules.scala 150:74:@327.4]
  wire [5:0] _T_54572; // @[Modules.scala 151:80:@328.4]
  wire [5:0] _GEN_11; // @[Modules.scala 150:103:@329.4]
  wire [6:0] _T_54573; // @[Modules.scala 150:103:@329.4]
  wire [5:0] _T_54574; // @[Modules.scala 150:103:@330.4]
  wire [5:0] _T_54575; // @[Modules.scala 150:103:@331.4]
  wire [5:0] _T_54577; // @[Modules.scala 150:74:@333.4]
  wire [4:0] _T_54579; // @[Modules.scala 151:80:@334.4]
  wire [5:0] _GEN_12; // @[Modules.scala 150:103:@335.4]
  wire [6:0] _T_54580; // @[Modules.scala 150:103:@335.4]
  wire [5:0] _T_54581; // @[Modules.scala 150:103:@336.4]
  wire [5:0] _T_54582; // @[Modules.scala 150:103:@337.4]
  wire [4:0] _T_54584; // @[Modules.scala 150:74:@339.4]
  wire [5:0] _T_54586; // @[Modules.scala 151:80:@340.4]
  wire [5:0] _GEN_13; // @[Modules.scala 150:103:@341.4]
  wire [6:0] _T_54587; // @[Modules.scala 150:103:@341.4]
  wire [5:0] _T_54588; // @[Modules.scala 150:103:@342.4]
  wire [5:0] _T_54589; // @[Modules.scala 150:103:@343.4]
  wire [5:0] _T_54591; // @[Modules.scala 150:74:@345.4]
  wire [5:0] _T_54593; // @[Modules.scala 151:80:@346.4]
  wire [6:0] _T_54594; // @[Modules.scala 150:103:@347.4]
  wire [5:0] _T_54595; // @[Modules.scala 150:103:@348.4]
  wire [5:0] _T_54596; // @[Modules.scala 150:103:@349.4]
  wire [5:0] _T_54598; // @[Modules.scala 150:74:@351.4]
  wire [5:0] _T_54600; // @[Modules.scala 151:80:@352.4]
  wire [6:0] _T_54601; // @[Modules.scala 150:103:@353.4]
  wire [5:0] _T_54602; // @[Modules.scala 150:103:@354.4]
  wire [5:0] _T_54603; // @[Modules.scala 150:103:@355.4]
  wire [5:0] _T_54605; // @[Modules.scala 150:74:@357.4]
  wire [4:0] _T_54607; // @[Modules.scala 151:80:@358.4]
  wire [5:0] _GEN_14; // @[Modules.scala 150:103:@359.4]
  wire [6:0] _T_54608; // @[Modules.scala 150:103:@359.4]
  wire [5:0] _T_54609; // @[Modules.scala 150:103:@360.4]
  wire [5:0] _T_54610; // @[Modules.scala 150:103:@361.4]
  wire [4:0] _T_54612; // @[Modules.scala 150:74:@363.4]
  wire [4:0] _T_54614; // @[Modules.scala 151:80:@364.4]
  wire [5:0] _T_54615; // @[Modules.scala 150:103:@365.4]
  wire [4:0] _T_54616; // @[Modules.scala 150:103:@366.4]
  wire [4:0] _T_54617; // @[Modules.scala 150:103:@367.4]
  wire [4:0] _T_54619; // @[Modules.scala 150:74:@369.4]
  wire [4:0] _T_54621; // @[Modules.scala 151:80:@370.4]
  wire [5:0] _T_54622; // @[Modules.scala 150:103:@371.4]
  wire [4:0] _T_54623; // @[Modules.scala 150:103:@372.4]
  wire [4:0] _T_54624; // @[Modules.scala 150:103:@373.4]
  wire [4:0] _T_54626; // @[Modules.scala 150:74:@375.4]
  wire [4:0] _T_54628; // @[Modules.scala 151:80:@376.4]
  wire [5:0] _T_54629; // @[Modules.scala 150:103:@377.4]
  wire [4:0] _T_54630; // @[Modules.scala 150:103:@378.4]
  wire [4:0] _T_54631; // @[Modules.scala 150:103:@379.4]
  wire [4:0] _T_54633; // @[Modules.scala 150:74:@381.4]
  wire [4:0] _T_54635; // @[Modules.scala 151:80:@382.4]
  wire [5:0] _T_54636; // @[Modules.scala 150:103:@383.4]
  wire [4:0] _T_54637; // @[Modules.scala 150:103:@384.4]
  wire [4:0] _T_54638; // @[Modules.scala 150:103:@385.4]
  wire [4:0] _T_54640; // @[Modules.scala 150:74:@387.4]
  wire [4:0] _T_54642; // @[Modules.scala 151:80:@388.4]
  wire [5:0] _T_54643; // @[Modules.scala 150:103:@389.4]
  wire [4:0] _T_54644; // @[Modules.scala 150:103:@390.4]
  wire [4:0] _T_54645; // @[Modules.scala 150:103:@391.4]
  wire [4:0] _T_54647; // @[Modules.scala 150:74:@393.4]
  wire [4:0] _T_54649; // @[Modules.scala 151:80:@394.4]
  wire [5:0] _T_54650; // @[Modules.scala 150:103:@395.4]
  wire [4:0] _T_54651; // @[Modules.scala 150:103:@396.4]
  wire [4:0] _T_54652; // @[Modules.scala 150:103:@397.4]
  wire [5:0] _T_54654; // @[Modules.scala 150:74:@399.4]
  wire [4:0] _T_54656; // @[Modules.scala 151:80:@400.4]
  wire [5:0] _GEN_15; // @[Modules.scala 150:103:@401.4]
  wire [6:0] _T_54657; // @[Modules.scala 150:103:@401.4]
  wire [5:0] _T_54658; // @[Modules.scala 150:103:@402.4]
  wire [5:0] _T_54659; // @[Modules.scala 150:103:@403.4]
  wire [5:0] _T_54661; // @[Modules.scala 150:74:@405.4]
  wire [5:0] _T_54663; // @[Modules.scala 151:80:@406.4]
  wire [6:0] _T_54664; // @[Modules.scala 150:103:@407.4]
  wire [5:0] _T_54665; // @[Modules.scala 150:103:@408.4]
  wire [5:0] _T_54666; // @[Modules.scala 150:103:@409.4]
  wire [5:0] _T_54668; // @[Modules.scala 150:74:@411.4]
  wire [5:0] _T_54670; // @[Modules.scala 151:80:@412.4]
  wire [6:0] _T_54671; // @[Modules.scala 150:103:@413.4]
  wire [5:0] _T_54672; // @[Modules.scala 150:103:@414.4]
  wire [5:0] _T_54673; // @[Modules.scala 150:103:@415.4]
  wire [5:0] _T_54675; // @[Modules.scala 150:74:@417.4]
  wire [5:0] _T_54677; // @[Modules.scala 151:80:@418.4]
  wire [6:0] _T_54678; // @[Modules.scala 150:103:@419.4]
  wire [5:0] _T_54679; // @[Modules.scala 150:103:@420.4]
  wire [5:0] _T_54680; // @[Modules.scala 150:103:@421.4]
  wire [5:0] _T_54682; // @[Modules.scala 150:74:@423.4]
  wire [4:0] _T_54684; // @[Modules.scala 151:80:@424.4]
  wire [5:0] _GEN_16; // @[Modules.scala 150:103:@425.4]
  wire [6:0] _T_54685; // @[Modules.scala 150:103:@425.4]
  wire [5:0] _T_54686; // @[Modules.scala 150:103:@426.4]
  wire [5:0] _T_54687; // @[Modules.scala 150:103:@427.4]
  wire [5:0] _T_54689; // @[Modules.scala 150:74:@429.4]
  wire [4:0] _T_54691; // @[Modules.scala 151:80:@430.4]
  wire [5:0] _GEN_17; // @[Modules.scala 150:103:@431.4]
  wire [6:0] _T_54692; // @[Modules.scala 150:103:@431.4]
  wire [5:0] _T_54693; // @[Modules.scala 150:103:@432.4]
  wire [5:0] _T_54694; // @[Modules.scala 150:103:@433.4]
  wire [4:0] _T_54696; // @[Modules.scala 150:74:@435.4]
  wire [4:0] _T_54698; // @[Modules.scala 151:80:@436.4]
  wire [5:0] _T_54699; // @[Modules.scala 150:103:@437.4]
  wire [4:0] _T_54700; // @[Modules.scala 150:103:@438.4]
  wire [4:0] _T_54701; // @[Modules.scala 150:103:@439.4]
  wire [4:0] _T_54703; // @[Modules.scala 150:74:@441.4]
  wire [4:0] _T_54705; // @[Modules.scala 151:80:@442.4]
  wire [5:0] _T_54706; // @[Modules.scala 150:103:@443.4]
  wire [4:0] _T_54707; // @[Modules.scala 150:103:@444.4]
  wire [4:0] _T_54708; // @[Modules.scala 150:103:@445.4]
  wire [4:0] _T_54710; // @[Modules.scala 150:74:@447.4]
  wire [4:0] _T_54712; // @[Modules.scala 151:80:@448.4]
  wire [5:0] _T_54713; // @[Modules.scala 150:103:@449.4]
  wire [4:0] _T_54714; // @[Modules.scala 150:103:@450.4]
  wire [4:0] _T_54715; // @[Modules.scala 150:103:@451.4]
  wire [4:0] _T_54717; // @[Modules.scala 150:74:@453.4]
  wire [4:0] _T_54719; // @[Modules.scala 151:80:@454.4]
  wire [5:0] _T_54720; // @[Modules.scala 150:103:@455.4]
  wire [4:0] _T_54721; // @[Modules.scala 150:103:@456.4]
  wire [4:0] _T_54722; // @[Modules.scala 150:103:@457.4]
  wire [5:0] _T_54724; // @[Modules.scala 150:74:@459.4]
  wire [4:0] _T_54726; // @[Modules.scala 151:80:@460.4]
  wire [5:0] _GEN_18; // @[Modules.scala 150:103:@461.4]
  wire [6:0] _T_54727; // @[Modules.scala 150:103:@461.4]
  wire [5:0] _T_54728; // @[Modules.scala 150:103:@462.4]
  wire [5:0] _T_54729; // @[Modules.scala 150:103:@463.4]
  wire [5:0] _T_54731; // @[Modules.scala 150:74:@465.4]
  wire [5:0] _T_54733; // @[Modules.scala 151:80:@466.4]
  wire [6:0] _T_54734; // @[Modules.scala 150:103:@467.4]
  wire [5:0] _T_54735; // @[Modules.scala 150:103:@468.4]
  wire [5:0] _T_54736; // @[Modules.scala 150:103:@469.4]
  wire [5:0] _T_54738; // @[Modules.scala 150:74:@471.4]
  wire [5:0] _T_54740; // @[Modules.scala 151:80:@472.4]
  wire [6:0] _T_54741; // @[Modules.scala 150:103:@473.4]
  wire [5:0] _T_54742; // @[Modules.scala 150:103:@474.4]
  wire [5:0] _T_54743; // @[Modules.scala 150:103:@475.4]
  wire [5:0] _T_54745; // @[Modules.scala 150:74:@477.4]
  wire [5:0] _T_54747; // @[Modules.scala 151:80:@478.4]
  wire [6:0] _T_54748; // @[Modules.scala 150:103:@479.4]
  wire [5:0] _T_54749; // @[Modules.scala 150:103:@480.4]
  wire [5:0] _T_54750; // @[Modules.scala 150:103:@481.4]
  wire [5:0] _T_54752; // @[Modules.scala 150:74:@483.4]
  wire [5:0] _T_54754; // @[Modules.scala 151:80:@484.4]
  wire [6:0] _T_54755; // @[Modules.scala 150:103:@485.4]
  wire [5:0] _T_54756; // @[Modules.scala 150:103:@486.4]
  wire [5:0] _T_54757; // @[Modules.scala 150:103:@487.4]
  wire [4:0] _T_54759; // @[Modules.scala 150:74:@489.4]
  wire [5:0] _T_54761; // @[Modules.scala 151:80:@490.4]
  wire [5:0] _GEN_19; // @[Modules.scala 150:103:@491.4]
  wire [6:0] _T_54762; // @[Modules.scala 150:103:@491.4]
  wire [5:0] _T_54763; // @[Modules.scala 150:103:@492.4]
  wire [5:0] _T_54764; // @[Modules.scala 150:103:@493.4]
  wire [5:0] _T_54766; // @[Modules.scala 150:74:@495.4]
  wire [4:0] _T_54768; // @[Modules.scala 151:80:@496.4]
  wire [5:0] _GEN_20; // @[Modules.scala 150:103:@497.4]
  wire [6:0] _T_54769; // @[Modules.scala 150:103:@497.4]
  wire [5:0] _T_54770; // @[Modules.scala 150:103:@498.4]
  wire [5:0] _T_54771; // @[Modules.scala 150:103:@499.4]
  wire [4:0] _T_54773; // @[Modules.scala 150:74:@501.4]
  wire [4:0] _T_54775; // @[Modules.scala 151:80:@502.4]
  wire [5:0] _T_54776; // @[Modules.scala 150:103:@503.4]
  wire [4:0] _T_54777; // @[Modules.scala 150:103:@504.4]
  wire [4:0] _T_54778; // @[Modules.scala 150:103:@505.4]
  wire [4:0] _T_54780; // @[Modules.scala 150:74:@507.4]
  wire [4:0] _T_54782; // @[Modules.scala 151:80:@508.4]
  wire [5:0] _T_54783; // @[Modules.scala 150:103:@509.4]
  wire [4:0] _T_54784; // @[Modules.scala 150:103:@510.4]
  wire [4:0] _T_54785; // @[Modules.scala 150:103:@511.4]
  wire [4:0] _T_54787; // @[Modules.scala 150:74:@513.4]
  wire [4:0] _T_54789; // @[Modules.scala 151:80:@514.4]
  wire [5:0] _T_54790; // @[Modules.scala 150:103:@515.4]
  wire [4:0] _T_54791; // @[Modules.scala 150:103:@516.4]
  wire [4:0] _T_54792; // @[Modules.scala 150:103:@517.4]
  wire [4:0] _T_54794; // @[Modules.scala 150:74:@519.4]
  wire [4:0] _T_54796; // @[Modules.scala 151:80:@520.4]
  wire [5:0] _T_54797; // @[Modules.scala 150:103:@521.4]
  wire [4:0] _T_54798; // @[Modules.scala 150:103:@522.4]
  wire [4:0] _T_54799; // @[Modules.scala 150:103:@523.4]
  wire [4:0] _T_54801; // @[Modules.scala 150:74:@525.4]
  wire [4:0] _T_54803; // @[Modules.scala 151:80:@526.4]
  wire [5:0] _T_54804; // @[Modules.scala 150:103:@527.4]
  wire [4:0] _T_54805; // @[Modules.scala 150:103:@528.4]
  wire [4:0] _T_54806; // @[Modules.scala 150:103:@529.4]
  wire [5:0] _T_54808; // @[Modules.scala 150:74:@531.4]
  wire [4:0] _T_54810; // @[Modules.scala 151:80:@532.4]
  wire [5:0] _GEN_21; // @[Modules.scala 150:103:@533.4]
  wire [6:0] _T_54811; // @[Modules.scala 150:103:@533.4]
  wire [5:0] _T_54812; // @[Modules.scala 150:103:@534.4]
  wire [5:0] _T_54813; // @[Modules.scala 150:103:@535.4]
  wire [5:0] _T_54815; // @[Modules.scala 150:74:@537.4]
  wire [5:0] _T_54817; // @[Modules.scala 151:80:@538.4]
  wire [6:0] _T_54818; // @[Modules.scala 150:103:@539.4]
  wire [5:0] _T_54819; // @[Modules.scala 150:103:@540.4]
  wire [5:0] _T_54820; // @[Modules.scala 150:103:@541.4]
  wire [5:0] _T_54822; // @[Modules.scala 150:74:@543.4]
  wire [5:0] _T_54824; // @[Modules.scala 151:80:@544.4]
  wire [6:0] _T_54825; // @[Modules.scala 150:103:@545.4]
  wire [5:0] _T_54826; // @[Modules.scala 150:103:@546.4]
  wire [5:0] _T_54827; // @[Modules.scala 150:103:@547.4]
  wire [4:0] _T_54829; // @[Modules.scala 150:74:@549.4]
  wire [4:0] _T_54831; // @[Modules.scala 151:80:@550.4]
  wire [5:0] _T_54832; // @[Modules.scala 150:103:@551.4]
  wire [4:0] _T_54833; // @[Modules.scala 150:103:@552.4]
  wire [4:0] _T_54834; // @[Modules.scala 150:103:@553.4]
  wire [4:0] _T_54836; // @[Modules.scala 150:74:@555.4]
  wire [4:0] _T_54838; // @[Modules.scala 151:80:@556.4]
  wire [5:0] _T_54839; // @[Modules.scala 150:103:@557.4]
  wire [4:0] _T_54840; // @[Modules.scala 150:103:@558.4]
  wire [4:0] _T_54841; // @[Modules.scala 150:103:@559.4]
  wire [4:0] _T_54843; // @[Modules.scala 150:74:@561.4]
  wire [5:0] _T_54845; // @[Modules.scala 151:80:@562.4]
  wire [5:0] _GEN_22; // @[Modules.scala 150:103:@563.4]
  wire [6:0] _T_54846; // @[Modules.scala 150:103:@563.4]
  wire [5:0] _T_54847; // @[Modules.scala 150:103:@564.4]
  wire [5:0] _T_54848; // @[Modules.scala 150:103:@565.4]
  wire [5:0] _T_54850; // @[Modules.scala 150:74:@567.4]
  wire [4:0] _T_54852; // @[Modules.scala 151:80:@568.4]
  wire [5:0] _GEN_23; // @[Modules.scala 150:103:@569.4]
  wire [6:0] _T_54853; // @[Modules.scala 150:103:@569.4]
  wire [5:0] _T_54854; // @[Modules.scala 150:103:@570.4]
  wire [5:0] _T_54855; // @[Modules.scala 150:103:@571.4]
  wire [4:0] _T_54857; // @[Modules.scala 150:74:@573.4]
  wire [4:0] _T_54859; // @[Modules.scala 151:80:@574.4]
  wire [5:0] _T_54860; // @[Modules.scala 150:103:@575.4]
  wire [4:0] _T_54861; // @[Modules.scala 150:103:@576.4]
  wire [4:0] _T_54862; // @[Modules.scala 150:103:@577.4]
  wire [4:0] _T_54864; // @[Modules.scala 150:74:@579.4]
  wire [4:0] _T_54866; // @[Modules.scala 151:80:@580.4]
  wire [5:0] _T_54867; // @[Modules.scala 150:103:@581.4]
  wire [4:0] _T_54868; // @[Modules.scala 150:103:@582.4]
  wire [4:0] _T_54869; // @[Modules.scala 150:103:@583.4]
  wire [4:0] _T_54871; // @[Modules.scala 150:74:@585.4]
  wire [4:0] _T_54873; // @[Modules.scala 151:80:@586.4]
  wire [5:0] _T_54874; // @[Modules.scala 150:103:@587.4]
  wire [4:0] _T_54875; // @[Modules.scala 150:103:@588.4]
  wire [4:0] _T_54876; // @[Modules.scala 150:103:@589.4]
  wire [4:0] _T_54878; // @[Modules.scala 150:74:@591.4]
  wire [4:0] _T_54880; // @[Modules.scala 151:80:@592.4]
  wire [5:0] _T_54881; // @[Modules.scala 150:103:@593.4]
  wire [4:0] _T_54882; // @[Modules.scala 150:103:@594.4]
  wire [4:0] _T_54883; // @[Modules.scala 150:103:@595.4]
  wire [4:0] _T_54885; // @[Modules.scala 150:74:@597.4]
  wire [4:0] _T_54887; // @[Modules.scala 151:80:@598.4]
  wire [5:0] _T_54888; // @[Modules.scala 150:103:@599.4]
  wire [4:0] _T_54889; // @[Modules.scala 150:103:@600.4]
  wire [4:0] _T_54890; // @[Modules.scala 150:103:@601.4]
  wire [4:0] _T_54892; // @[Modules.scala 150:74:@603.4]
  wire [4:0] _T_54894; // @[Modules.scala 151:80:@604.4]
  wire [5:0] _T_54895; // @[Modules.scala 150:103:@605.4]
  wire [4:0] _T_54896; // @[Modules.scala 150:103:@606.4]
  wire [4:0] _T_54897; // @[Modules.scala 150:103:@607.4]
  wire [5:0] _T_54899; // @[Modules.scala 150:74:@609.4]
  wire [5:0] _T_54901; // @[Modules.scala 151:80:@610.4]
  wire [6:0] _T_54902; // @[Modules.scala 150:103:@611.4]
  wire [5:0] _T_54903; // @[Modules.scala 150:103:@612.4]
  wire [5:0] _T_54904; // @[Modules.scala 150:103:@613.4]
  wire [5:0] _T_54906; // @[Modules.scala 150:74:@615.4]
  wire [4:0] _T_54908; // @[Modules.scala 151:80:@616.4]
  wire [5:0] _GEN_24; // @[Modules.scala 150:103:@617.4]
  wire [6:0] _T_54909; // @[Modules.scala 150:103:@617.4]
  wire [5:0] _T_54910; // @[Modules.scala 150:103:@618.4]
  wire [5:0] _T_54911; // @[Modules.scala 150:103:@619.4]
  wire [4:0] _T_54913; // @[Modules.scala 150:74:@621.4]
  wire [4:0] _T_54915; // @[Modules.scala 151:80:@622.4]
  wire [5:0] _T_54916; // @[Modules.scala 150:103:@623.4]
  wire [4:0] _T_54917; // @[Modules.scala 150:103:@624.4]
  wire [4:0] _T_54918; // @[Modules.scala 150:103:@625.4]
  wire [4:0] _T_54920; // @[Modules.scala 150:74:@627.4]
  wire [4:0] _T_54922; // @[Modules.scala 151:80:@628.4]
  wire [5:0] _T_54923; // @[Modules.scala 150:103:@629.4]
  wire [4:0] _T_54924; // @[Modules.scala 150:103:@630.4]
  wire [4:0] _T_54925; // @[Modules.scala 150:103:@631.4]
  wire [4:0] _T_54927; // @[Modules.scala 150:74:@633.4]
  wire [4:0] _T_54929; // @[Modules.scala 151:80:@634.4]
  wire [5:0] _T_54930; // @[Modules.scala 150:103:@635.4]
  wire [4:0] _T_54931; // @[Modules.scala 150:103:@636.4]
  wire [4:0] _T_54932; // @[Modules.scala 150:103:@637.4]
  wire [4:0] _T_54934; // @[Modules.scala 150:74:@639.4]
  wire [4:0] _T_54936; // @[Modules.scala 151:80:@640.4]
  wire [5:0] _T_54937; // @[Modules.scala 150:103:@641.4]
  wire [4:0] _T_54938; // @[Modules.scala 150:103:@642.4]
  wire [4:0] _T_54939; // @[Modules.scala 150:103:@643.4]
  wire [4:0] _T_54941; // @[Modules.scala 150:74:@645.4]
  wire [5:0] _T_54943; // @[Modules.scala 151:80:@646.4]
  wire [5:0] _GEN_25; // @[Modules.scala 150:103:@647.4]
  wire [6:0] _T_54944; // @[Modules.scala 150:103:@647.4]
  wire [5:0] _T_54945; // @[Modules.scala 150:103:@648.4]
  wire [5:0] _T_54946; // @[Modules.scala 150:103:@649.4]
  wire [5:0] _T_54948; // @[Modules.scala 150:74:@651.4]
  wire [5:0] _T_54950; // @[Modules.scala 151:80:@652.4]
  wire [6:0] _T_54951; // @[Modules.scala 150:103:@653.4]
  wire [5:0] _T_54952; // @[Modules.scala 150:103:@654.4]
  wire [5:0] _T_54953; // @[Modules.scala 150:103:@655.4]
  wire [4:0] _T_54955; // @[Modules.scala 150:74:@657.4]
  wire [4:0] _T_54957; // @[Modules.scala 151:80:@658.4]
  wire [5:0] _T_54958; // @[Modules.scala 150:103:@659.4]
  wire [4:0] _T_54959; // @[Modules.scala 150:103:@660.4]
  wire [4:0] _T_54960; // @[Modules.scala 150:103:@661.4]
  wire [4:0] _T_54962; // @[Modules.scala 150:74:@663.4]
  wire [4:0] _T_54964; // @[Modules.scala 151:80:@664.4]
  wire [5:0] _T_54965; // @[Modules.scala 150:103:@665.4]
  wire [4:0] _T_54966; // @[Modules.scala 150:103:@666.4]
  wire [4:0] _T_54967; // @[Modules.scala 150:103:@667.4]
  wire [4:0] _T_54969; // @[Modules.scala 150:74:@669.4]
  wire [4:0] _T_54971; // @[Modules.scala 151:80:@670.4]
  wire [5:0] _T_54972; // @[Modules.scala 150:103:@671.4]
  wire [4:0] _T_54973; // @[Modules.scala 150:103:@672.4]
  wire [4:0] _T_54974; // @[Modules.scala 150:103:@673.4]
  wire [4:0] _T_54976; // @[Modules.scala 150:74:@675.4]
  wire [4:0] _T_54978; // @[Modules.scala 151:80:@676.4]
  wire [5:0] _T_54979; // @[Modules.scala 150:103:@677.4]
  wire [4:0] _T_54980; // @[Modules.scala 150:103:@678.4]
  wire [4:0] _T_54981; // @[Modules.scala 150:103:@679.4]
  wire [4:0] _T_54983; // @[Modules.scala 150:74:@681.4]
  wire [4:0] _T_54985; // @[Modules.scala 151:80:@682.4]
  wire [5:0] _T_54986; // @[Modules.scala 150:103:@683.4]
  wire [4:0] _T_54987; // @[Modules.scala 150:103:@684.4]
  wire [4:0] _T_54988; // @[Modules.scala 150:103:@685.4]
  wire [5:0] _T_54990; // @[Modules.scala 150:74:@687.4]
  wire [4:0] _T_54992; // @[Modules.scala 151:80:@688.4]
  wire [5:0] _GEN_26; // @[Modules.scala 150:103:@689.4]
  wire [6:0] _T_54993; // @[Modules.scala 150:103:@689.4]
  wire [5:0] _T_54994; // @[Modules.scala 150:103:@690.4]
  wire [5:0] _T_54995; // @[Modules.scala 150:103:@691.4]
  wire [5:0] _T_54997; // @[Modules.scala 150:74:@693.4]
  wire [4:0] _T_54999; // @[Modules.scala 151:80:@694.4]
  wire [5:0] _GEN_27; // @[Modules.scala 150:103:@695.4]
  wire [6:0] _T_55000; // @[Modules.scala 150:103:@695.4]
  wire [5:0] _T_55001; // @[Modules.scala 150:103:@696.4]
  wire [5:0] _T_55002; // @[Modules.scala 150:103:@697.4]
  wire [4:0] _T_55004; // @[Modules.scala 150:74:@699.4]
  wire [4:0] _T_55006; // @[Modules.scala 151:80:@700.4]
  wire [5:0] _T_55007; // @[Modules.scala 150:103:@701.4]
  wire [4:0] _T_55008; // @[Modules.scala 150:103:@702.4]
  wire [4:0] _T_55009; // @[Modules.scala 150:103:@703.4]
  wire [4:0] _T_55011; // @[Modules.scala 150:74:@705.4]
  wire [4:0] _T_55013; // @[Modules.scala 151:80:@706.4]
  wire [5:0] _T_55014; // @[Modules.scala 150:103:@707.4]
  wire [4:0] _T_55015; // @[Modules.scala 150:103:@708.4]
  wire [4:0] _T_55016; // @[Modules.scala 150:103:@709.4]
  wire [4:0] _T_55018; // @[Modules.scala 150:74:@711.4]
  wire [4:0] _T_55020; // @[Modules.scala 151:80:@712.4]
  wire [5:0] _T_55021; // @[Modules.scala 150:103:@713.4]
  wire [4:0] _T_55022; // @[Modules.scala 150:103:@714.4]
  wire [4:0] _T_55023; // @[Modules.scala 150:103:@715.4]
  wire [4:0] _T_55025; // @[Modules.scala 150:74:@717.4]
  wire [4:0] _T_55027; // @[Modules.scala 151:80:@718.4]
  wire [5:0] _T_55028; // @[Modules.scala 150:103:@719.4]
  wire [4:0] _T_55029; // @[Modules.scala 150:103:@720.4]
  wire [4:0] _T_55030; // @[Modules.scala 150:103:@721.4]
  wire [4:0] _T_55032; // @[Modules.scala 150:74:@723.4]
  wire [5:0] _T_55034; // @[Modules.scala 151:80:@724.4]
  wire [5:0] _GEN_28; // @[Modules.scala 150:103:@725.4]
  wire [6:0] _T_55035; // @[Modules.scala 150:103:@725.4]
  wire [5:0] _T_55036; // @[Modules.scala 150:103:@726.4]
  wire [5:0] _T_55037; // @[Modules.scala 150:103:@727.4]
  wire [4:0] _T_55039; // @[Modules.scala 150:74:@729.4]
  wire [4:0] _T_55041; // @[Modules.scala 151:80:@730.4]
  wire [5:0] _T_55042; // @[Modules.scala 150:103:@731.4]
  wire [4:0] _T_55043; // @[Modules.scala 150:103:@732.4]
  wire [4:0] _T_55044; // @[Modules.scala 150:103:@733.4]
  wire [4:0] _T_55046; // @[Modules.scala 150:74:@735.4]
  wire [4:0] _T_55048; // @[Modules.scala 151:80:@736.4]
  wire [5:0] _T_55049; // @[Modules.scala 150:103:@737.4]
  wire [4:0] _T_55050; // @[Modules.scala 150:103:@738.4]
  wire [4:0] _T_55051; // @[Modules.scala 150:103:@739.4]
  wire [4:0] _T_55053; // @[Modules.scala 150:74:@741.4]
  wire [4:0] _T_55055; // @[Modules.scala 151:80:@742.4]
  wire [5:0] _T_55056; // @[Modules.scala 150:103:@743.4]
  wire [4:0] _T_55057; // @[Modules.scala 150:103:@744.4]
  wire [4:0] _T_55058; // @[Modules.scala 150:103:@745.4]
  wire [4:0] _T_55060; // @[Modules.scala 150:74:@747.4]
  wire [4:0] _T_55062; // @[Modules.scala 151:80:@748.4]
  wire [5:0] _T_55063; // @[Modules.scala 150:103:@749.4]
  wire [4:0] _T_55064; // @[Modules.scala 150:103:@750.4]
  wire [4:0] _T_55065; // @[Modules.scala 150:103:@751.4]
  wire [4:0] _T_55067; // @[Modules.scala 150:74:@753.4]
  wire [4:0] _T_55069; // @[Modules.scala 151:80:@754.4]
  wire [5:0] _T_55070; // @[Modules.scala 150:103:@755.4]
  wire [4:0] _T_55071; // @[Modules.scala 150:103:@756.4]
  wire [4:0] _T_55072; // @[Modules.scala 150:103:@757.4]
  wire [4:0] _T_55074; // @[Modules.scala 150:74:@759.4]
  wire [5:0] _T_55076; // @[Modules.scala 151:80:@760.4]
  wire [5:0] _GEN_29; // @[Modules.scala 150:103:@761.4]
  wire [6:0] _T_55077; // @[Modules.scala 150:103:@761.4]
  wire [5:0] _T_55078; // @[Modules.scala 150:103:@762.4]
  wire [5:0] _T_55079; // @[Modules.scala 150:103:@763.4]
  wire [5:0] _T_55081; // @[Modules.scala 150:74:@765.4]
  wire [5:0] _T_55083; // @[Modules.scala 151:80:@766.4]
  wire [6:0] _T_55084; // @[Modules.scala 150:103:@767.4]
  wire [5:0] _T_55085; // @[Modules.scala 150:103:@768.4]
  wire [5:0] _T_55086; // @[Modules.scala 150:103:@769.4]
  wire [4:0] _T_55088; // @[Modules.scala 150:74:@771.4]
  wire [4:0] _T_55090; // @[Modules.scala 151:80:@772.4]
  wire [5:0] _T_55091; // @[Modules.scala 150:103:@773.4]
  wire [4:0] _T_55092; // @[Modules.scala 150:103:@774.4]
  wire [4:0] _T_55093; // @[Modules.scala 150:103:@775.4]
  wire [4:0] _T_55095; // @[Modules.scala 150:74:@777.4]
  wire [4:0] _T_55097; // @[Modules.scala 151:80:@778.4]
  wire [5:0] _T_55098; // @[Modules.scala 150:103:@779.4]
  wire [4:0] _T_55099; // @[Modules.scala 150:103:@780.4]
  wire [4:0] _T_55100; // @[Modules.scala 150:103:@781.4]
  wire [4:0] _T_55102; // @[Modules.scala 150:74:@783.4]
  wire [4:0] _T_55104; // @[Modules.scala 151:80:@784.4]
  wire [5:0] _T_55105; // @[Modules.scala 150:103:@785.4]
  wire [4:0] _T_55106; // @[Modules.scala 150:103:@786.4]
  wire [4:0] _T_55107; // @[Modules.scala 150:103:@787.4]
  wire [4:0] _T_55109; // @[Modules.scala 150:74:@789.4]
  wire [4:0] _T_55111; // @[Modules.scala 151:80:@790.4]
  wire [5:0] _T_55112; // @[Modules.scala 150:103:@791.4]
  wire [4:0] _T_55113; // @[Modules.scala 150:103:@792.4]
  wire [4:0] _T_55114; // @[Modules.scala 150:103:@793.4]
  wire [4:0] _T_55116; // @[Modules.scala 150:74:@795.4]
  wire [4:0] _T_55118; // @[Modules.scala 151:80:@796.4]
  wire [5:0] _T_55119; // @[Modules.scala 150:103:@797.4]
  wire [4:0] _T_55120; // @[Modules.scala 150:103:@798.4]
  wire [4:0] _T_55121; // @[Modules.scala 150:103:@799.4]
  wire [5:0] _T_55123; // @[Modules.scala 150:74:@801.4]
  wire [5:0] _T_55125; // @[Modules.scala 151:80:@802.4]
  wire [6:0] _T_55126; // @[Modules.scala 150:103:@803.4]
  wire [5:0] _T_55127; // @[Modules.scala 150:103:@804.4]
  wire [5:0] _T_55128; // @[Modules.scala 150:103:@805.4]
  wire [4:0] _T_55130; // @[Modules.scala 150:74:@807.4]
  wire [4:0] _T_55132; // @[Modules.scala 151:80:@808.4]
  wire [5:0] _T_55133; // @[Modules.scala 150:103:@809.4]
  wire [4:0] _T_55134; // @[Modules.scala 150:103:@810.4]
  wire [4:0] _T_55135; // @[Modules.scala 150:103:@811.4]
  wire [5:0] _T_55137; // @[Modules.scala 150:74:@813.4]
  wire [4:0] _T_55139; // @[Modules.scala 151:80:@814.4]
  wire [5:0] _GEN_30; // @[Modules.scala 150:103:@815.4]
  wire [6:0] _T_55140; // @[Modules.scala 150:103:@815.4]
  wire [5:0] _T_55141; // @[Modules.scala 150:103:@816.4]
  wire [5:0] _T_55142; // @[Modules.scala 150:103:@817.4]
  wire [4:0] _T_55144; // @[Modules.scala 150:74:@819.4]
  wire [4:0] _T_55146; // @[Modules.scala 151:80:@820.4]
  wire [5:0] _T_55147; // @[Modules.scala 150:103:@821.4]
  wire [4:0] _T_55148; // @[Modules.scala 150:103:@822.4]
  wire [4:0] _T_55149; // @[Modules.scala 150:103:@823.4]
  wire [5:0] _T_55151; // @[Modules.scala 150:74:@825.4]
  wire [4:0] _T_55153; // @[Modules.scala 151:80:@826.4]
  wire [5:0] _GEN_31; // @[Modules.scala 150:103:@827.4]
  wire [6:0] _T_55154; // @[Modules.scala 150:103:@827.4]
  wire [5:0] _T_55155; // @[Modules.scala 150:103:@828.4]
  wire [5:0] _T_55156; // @[Modules.scala 150:103:@829.4]
  wire [4:0] _T_55158; // @[Modules.scala 150:74:@831.4]
  wire [5:0] _T_55160; // @[Modules.scala 151:80:@832.4]
  wire [5:0] _GEN_32; // @[Modules.scala 150:103:@833.4]
  wire [6:0] _T_55161; // @[Modules.scala 150:103:@833.4]
  wire [5:0] _T_55162; // @[Modules.scala 150:103:@834.4]
  wire [5:0] _T_55163; // @[Modules.scala 150:103:@835.4]
  wire [5:0] _T_55165; // @[Modules.scala 150:74:@837.4]
  wire [5:0] _T_55167; // @[Modules.scala 151:80:@838.4]
  wire [6:0] _T_55168; // @[Modules.scala 150:103:@839.4]
  wire [5:0] _T_55169; // @[Modules.scala 150:103:@840.4]
  wire [5:0] _T_55170; // @[Modules.scala 150:103:@841.4]
  wire [5:0] _T_55172; // @[Modules.scala 150:74:@843.4]
  wire [5:0] _T_55174; // @[Modules.scala 151:80:@844.4]
  wire [6:0] _T_55175; // @[Modules.scala 150:103:@845.4]
  wire [5:0] _T_55176; // @[Modules.scala 150:103:@846.4]
  wire [5:0] _T_55177; // @[Modules.scala 150:103:@847.4]
  wire [4:0] _T_55179; // @[Modules.scala 150:74:@849.4]
  wire [4:0] _T_55181; // @[Modules.scala 151:80:@850.4]
  wire [5:0] _T_55182; // @[Modules.scala 150:103:@851.4]
  wire [4:0] _T_55183; // @[Modules.scala 150:103:@852.4]
  wire [4:0] _T_55184; // @[Modules.scala 150:103:@853.4]
  wire [4:0] _T_55186; // @[Modules.scala 150:74:@855.4]
  wire [4:0] _T_55188; // @[Modules.scala 151:80:@856.4]
  wire [5:0] _T_55189; // @[Modules.scala 150:103:@857.4]
  wire [4:0] _T_55190; // @[Modules.scala 150:103:@858.4]
  wire [4:0] _T_55191; // @[Modules.scala 150:103:@859.4]
  wire [4:0] _T_55193; // @[Modules.scala 150:74:@861.4]
  wire [4:0] _T_55195; // @[Modules.scala 151:80:@862.4]
  wire [5:0] _T_55196; // @[Modules.scala 150:103:@863.4]
  wire [4:0] _T_55197; // @[Modules.scala 150:103:@864.4]
  wire [4:0] _T_55198; // @[Modules.scala 150:103:@865.4]
  wire [4:0] _T_55200; // @[Modules.scala 150:74:@867.4]
  wire [4:0] _T_55202; // @[Modules.scala 151:80:@868.4]
  wire [5:0] _T_55203; // @[Modules.scala 150:103:@869.4]
  wire [4:0] _T_55204; // @[Modules.scala 150:103:@870.4]
  wire [4:0] _T_55205; // @[Modules.scala 150:103:@871.4]
  wire [4:0] _T_55207; // @[Modules.scala 150:74:@873.4]
  wire [4:0] _T_55209; // @[Modules.scala 151:80:@874.4]
  wire [5:0] _T_55210; // @[Modules.scala 150:103:@875.4]
  wire [4:0] _T_55211; // @[Modules.scala 150:103:@876.4]
  wire [4:0] _T_55212; // @[Modules.scala 150:103:@877.4]
  wire [5:0] _T_55214; // @[Modules.scala 150:74:@879.4]
  wire [4:0] _T_55216; // @[Modules.scala 151:80:@880.4]
  wire [5:0] _GEN_33; // @[Modules.scala 150:103:@881.4]
  wire [6:0] _T_55217; // @[Modules.scala 150:103:@881.4]
  wire [5:0] _T_55218; // @[Modules.scala 150:103:@882.4]
  wire [5:0] _T_55219; // @[Modules.scala 150:103:@883.4]
  wire [5:0] _T_55221; // @[Modules.scala 150:74:@885.4]
  wire [4:0] _T_55223; // @[Modules.scala 151:80:@886.4]
  wire [5:0] _GEN_34; // @[Modules.scala 150:103:@887.4]
  wire [6:0] _T_55224; // @[Modules.scala 150:103:@887.4]
  wire [5:0] _T_55225; // @[Modules.scala 150:103:@888.4]
  wire [5:0] _T_55226; // @[Modules.scala 150:103:@889.4]
  wire [4:0] _T_55228; // @[Modules.scala 150:74:@891.4]
  wire [5:0] _T_55230; // @[Modules.scala 151:80:@892.4]
  wire [5:0] _GEN_35; // @[Modules.scala 150:103:@893.4]
  wire [6:0] _T_55231; // @[Modules.scala 150:103:@893.4]
  wire [5:0] _T_55232; // @[Modules.scala 150:103:@894.4]
  wire [5:0] _T_55233; // @[Modules.scala 150:103:@895.4]
  wire [5:0] _T_55235; // @[Modules.scala 150:74:@897.4]
  wire [4:0] _T_55237; // @[Modules.scala 151:80:@898.4]
  wire [5:0] _GEN_36; // @[Modules.scala 150:103:@899.4]
  wire [6:0] _T_55238; // @[Modules.scala 150:103:@899.4]
  wire [5:0] _T_55239; // @[Modules.scala 150:103:@900.4]
  wire [5:0] _T_55240; // @[Modules.scala 150:103:@901.4]
  wire [4:0] _T_55242; // @[Modules.scala 150:74:@903.4]
  wire [5:0] _T_55244; // @[Modules.scala 151:80:@904.4]
  wire [5:0] _GEN_37; // @[Modules.scala 150:103:@905.4]
  wire [6:0] _T_55245; // @[Modules.scala 150:103:@905.4]
  wire [5:0] _T_55246; // @[Modules.scala 150:103:@906.4]
  wire [5:0] _T_55247; // @[Modules.scala 150:103:@907.4]
  wire [5:0] _T_55249; // @[Modules.scala 150:74:@909.4]
  wire [4:0] _T_55251; // @[Modules.scala 151:80:@910.4]
  wire [5:0] _GEN_38; // @[Modules.scala 150:103:@911.4]
  wire [6:0] _T_55252; // @[Modules.scala 150:103:@911.4]
  wire [5:0] _T_55253; // @[Modules.scala 150:103:@912.4]
  wire [5:0] _T_55254; // @[Modules.scala 150:103:@913.4]
  wire [5:0] _T_55256; // @[Modules.scala 150:74:@915.4]
  wire [5:0] _T_55258; // @[Modules.scala 151:80:@916.4]
  wire [6:0] _T_55259; // @[Modules.scala 150:103:@917.4]
  wire [5:0] _T_55260; // @[Modules.scala 150:103:@918.4]
  wire [5:0] _T_55261; // @[Modules.scala 150:103:@919.4]
  wire [4:0] _T_55263; // @[Modules.scala 150:74:@921.4]
  wire [4:0] _T_55265; // @[Modules.scala 151:80:@922.4]
  wire [5:0] _T_55266; // @[Modules.scala 150:103:@923.4]
  wire [4:0] _T_55267; // @[Modules.scala 150:103:@924.4]
  wire [4:0] _T_55268; // @[Modules.scala 150:103:@925.4]
  wire [4:0] _T_55270; // @[Modules.scala 150:74:@927.4]
  wire [4:0] _T_55272; // @[Modules.scala 151:80:@928.4]
  wire [5:0] _T_55273; // @[Modules.scala 150:103:@929.4]
  wire [4:0] _T_55274; // @[Modules.scala 150:103:@930.4]
  wire [4:0] _T_55275; // @[Modules.scala 150:103:@931.4]
  wire [4:0] _T_55277; // @[Modules.scala 150:74:@933.4]
  wire [4:0] _T_55279; // @[Modules.scala 151:80:@934.4]
  wire [5:0] _T_55280; // @[Modules.scala 150:103:@935.4]
  wire [4:0] _T_55281; // @[Modules.scala 150:103:@936.4]
  wire [4:0] _T_55282; // @[Modules.scala 150:103:@937.4]
  wire [4:0] _T_55284; // @[Modules.scala 150:74:@939.4]
  wire [4:0] _T_55286; // @[Modules.scala 151:80:@940.4]
  wire [5:0] _T_55287; // @[Modules.scala 150:103:@941.4]
  wire [4:0] _T_55288; // @[Modules.scala 150:103:@942.4]
  wire [4:0] _T_55289; // @[Modules.scala 150:103:@943.4]
  wire [4:0] _T_55291; // @[Modules.scala 150:74:@945.4]
  wire [5:0] _T_55293; // @[Modules.scala 151:80:@946.4]
  wire [5:0] _GEN_39; // @[Modules.scala 150:103:@947.4]
  wire [6:0] _T_55294; // @[Modules.scala 150:103:@947.4]
  wire [5:0] _T_55295; // @[Modules.scala 150:103:@948.4]
  wire [5:0] _T_55296; // @[Modules.scala 150:103:@949.4]
  wire [5:0] _T_55298; // @[Modules.scala 150:74:@951.4]
  wire [4:0] _T_55300; // @[Modules.scala 151:80:@952.4]
  wire [5:0] _GEN_40; // @[Modules.scala 150:103:@953.4]
  wire [6:0] _T_55301; // @[Modules.scala 150:103:@953.4]
  wire [5:0] _T_55302; // @[Modules.scala 150:103:@954.4]
  wire [5:0] _T_55303; // @[Modules.scala 150:103:@955.4]
  wire [4:0] _T_55305; // @[Modules.scala 150:74:@957.4]
  wire [5:0] _T_55307; // @[Modules.scala 151:80:@958.4]
  wire [5:0] _GEN_41; // @[Modules.scala 150:103:@959.4]
  wire [6:0] _T_55308; // @[Modules.scala 150:103:@959.4]
  wire [5:0] _T_55309; // @[Modules.scala 150:103:@960.4]
  wire [5:0] _T_55310; // @[Modules.scala 150:103:@961.4]
  wire [5:0] _T_55312; // @[Modules.scala 150:74:@963.4]
  wire [5:0] _T_55314; // @[Modules.scala 151:80:@964.4]
  wire [6:0] _T_55315; // @[Modules.scala 150:103:@965.4]
  wire [5:0] _T_55316; // @[Modules.scala 150:103:@966.4]
  wire [5:0] _T_55317; // @[Modules.scala 150:103:@967.4]
  wire [5:0] _T_55319; // @[Modules.scala 150:74:@969.4]
  wire [4:0] _T_55321; // @[Modules.scala 151:80:@970.4]
  wire [5:0] _GEN_42; // @[Modules.scala 150:103:@971.4]
  wire [6:0] _T_55322; // @[Modules.scala 150:103:@971.4]
  wire [5:0] _T_55323; // @[Modules.scala 150:103:@972.4]
  wire [5:0] _T_55324; // @[Modules.scala 150:103:@973.4]
  wire [5:0] _T_55326; // @[Modules.scala 150:74:@975.4]
  wire [5:0] _T_55328; // @[Modules.scala 151:80:@976.4]
  wire [6:0] _T_55329; // @[Modules.scala 150:103:@977.4]
  wire [5:0] _T_55330; // @[Modules.scala 150:103:@978.4]
  wire [5:0] _T_55331; // @[Modules.scala 150:103:@979.4]
  wire [4:0] _T_55333; // @[Modules.scala 150:74:@981.4]
  wire [5:0] _T_55335; // @[Modules.scala 151:80:@982.4]
  wire [5:0] _GEN_43; // @[Modules.scala 150:103:@983.4]
  wire [6:0] _T_55336; // @[Modules.scala 150:103:@983.4]
  wire [5:0] _T_55337; // @[Modules.scala 150:103:@984.4]
  wire [5:0] _T_55338; // @[Modules.scala 150:103:@985.4]
  wire [5:0] _T_55340; // @[Modules.scala 150:74:@987.4]
  wire [4:0] _T_55342; // @[Modules.scala 151:80:@988.4]
  wire [5:0] _GEN_44; // @[Modules.scala 150:103:@989.4]
  wire [6:0] _T_55343; // @[Modules.scala 150:103:@989.4]
  wire [5:0] _T_55344; // @[Modules.scala 150:103:@990.4]
  wire [5:0] _T_55345; // @[Modules.scala 150:103:@991.4]
  wire [4:0] _T_55347; // @[Modules.scala 150:74:@993.4]
  wire [4:0] _T_55349; // @[Modules.scala 151:80:@994.4]
  wire [5:0] _T_55350; // @[Modules.scala 150:103:@995.4]
  wire [4:0] _T_55351; // @[Modules.scala 150:103:@996.4]
  wire [4:0] _T_55352; // @[Modules.scala 150:103:@997.4]
  wire [4:0] _T_55354; // @[Modules.scala 150:74:@999.4]
  wire [4:0] _T_55356; // @[Modules.scala 151:80:@1000.4]
  wire [5:0] _T_55357; // @[Modules.scala 150:103:@1001.4]
  wire [4:0] _T_55358; // @[Modules.scala 150:103:@1002.4]
  wire [4:0] _T_55359; // @[Modules.scala 150:103:@1003.4]
  wire [4:0] _T_55361; // @[Modules.scala 150:74:@1005.4]
  wire [5:0] _T_55363; // @[Modules.scala 151:80:@1006.4]
  wire [5:0] _GEN_45; // @[Modules.scala 150:103:@1007.4]
  wire [6:0] _T_55364; // @[Modules.scala 150:103:@1007.4]
  wire [5:0] _T_55365; // @[Modules.scala 150:103:@1008.4]
  wire [5:0] _T_55366; // @[Modules.scala 150:103:@1009.4]
  wire [5:0] _T_55368; // @[Modules.scala 150:74:@1011.4]
  wire [5:0] _T_55370; // @[Modules.scala 151:80:@1012.4]
  wire [6:0] _T_55371; // @[Modules.scala 150:103:@1013.4]
  wire [5:0] _T_55372; // @[Modules.scala 150:103:@1014.4]
  wire [5:0] _T_55373; // @[Modules.scala 150:103:@1015.4]
  wire [5:0] _T_55375; // @[Modules.scala 150:74:@1017.4]
  wire [4:0] _T_55377; // @[Modules.scala 151:80:@1018.4]
  wire [5:0] _GEN_46; // @[Modules.scala 150:103:@1019.4]
  wire [6:0] _T_55378; // @[Modules.scala 150:103:@1019.4]
  wire [5:0] _T_55379; // @[Modules.scala 150:103:@1020.4]
  wire [5:0] _T_55380; // @[Modules.scala 150:103:@1021.4]
  wire [4:0] _T_55382; // @[Modules.scala 150:74:@1023.4]
  wire [5:0] _T_55384; // @[Modules.scala 151:80:@1024.4]
  wire [5:0] _GEN_47; // @[Modules.scala 150:103:@1025.4]
  wire [6:0] _T_55385; // @[Modules.scala 150:103:@1025.4]
  wire [5:0] _T_55386; // @[Modules.scala 150:103:@1026.4]
  wire [5:0] _T_55387; // @[Modules.scala 150:103:@1027.4]
  wire [5:0] _T_55389; // @[Modules.scala 150:74:@1029.4]
  wire [5:0] _T_55391; // @[Modules.scala 151:80:@1030.4]
  wire [6:0] _T_55392; // @[Modules.scala 150:103:@1031.4]
  wire [5:0] _T_55393; // @[Modules.scala 150:103:@1032.4]
  wire [5:0] _T_55394; // @[Modules.scala 150:103:@1033.4]
  wire [5:0] _T_55396; // @[Modules.scala 150:74:@1035.4]
  wire [4:0] _T_55398; // @[Modules.scala 151:80:@1036.4]
  wire [5:0] _GEN_48; // @[Modules.scala 150:103:@1037.4]
  wire [6:0] _T_55399; // @[Modules.scala 150:103:@1037.4]
  wire [5:0] _T_55400; // @[Modules.scala 150:103:@1038.4]
  wire [5:0] _T_55401; // @[Modules.scala 150:103:@1039.4]
  wire [4:0] _T_55403; // @[Modules.scala 150:74:@1041.4]
  wire [5:0] _T_55405; // @[Modules.scala 151:80:@1042.4]
  wire [5:0] _GEN_49; // @[Modules.scala 150:103:@1043.4]
  wire [6:0] _T_55406; // @[Modules.scala 150:103:@1043.4]
  wire [5:0] _T_55407; // @[Modules.scala 150:103:@1044.4]
  wire [5:0] _T_55408; // @[Modules.scala 150:103:@1045.4]
  wire [5:0] _T_55410; // @[Modules.scala 150:74:@1047.4]
  wire [5:0] _T_55412; // @[Modules.scala 151:80:@1048.4]
  wire [6:0] _T_55413; // @[Modules.scala 150:103:@1049.4]
  wire [5:0] _T_55414; // @[Modules.scala 150:103:@1050.4]
  wire [5:0] _T_55415; // @[Modules.scala 150:103:@1051.4]
  wire [4:0] _T_55417; // @[Modules.scala 150:74:@1053.4]
  wire [4:0] _T_55419; // @[Modules.scala 151:80:@1054.4]
  wire [5:0] _T_55420; // @[Modules.scala 150:103:@1055.4]
  wire [4:0] _T_55421; // @[Modules.scala 150:103:@1056.4]
  wire [4:0] _T_55422; // @[Modules.scala 150:103:@1057.4]
  wire [5:0] _T_55424; // @[Modules.scala 150:74:@1059.4]
  wire [5:0] _T_55426; // @[Modules.scala 151:80:@1060.4]
  wire [6:0] _T_55427; // @[Modules.scala 150:103:@1061.4]
  wire [5:0] _T_55428; // @[Modules.scala 150:103:@1062.4]
  wire [5:0] _T_55429; // @[Modules.scala 150:103:@1063.4]
  wire [4:0] _T_55431; // @[Modules.scala 150:74:@1065.4]
  wire [4:0] _T_55433; // @[Modules.scala 151:80:@1066.4]
  wire [5:0] _T_55434; // @[Modules.scala 150:103:@1067.4]
  wire [4:0] _T_55435; // @[Modules.scala 150:103:@1068.4]
  wire [4:0] _T_55436; // @[Modules.scala 150:103:@1069.4]
  wire [5:0] _T_55438; // @[Modules.scala 150:74:@1071.4]
  wire [5:0] _T_55440; // @[Modules.scala 151:80:@1072.4]
  wire [6:0] _T_55441; // @[Modules.scala 150:103:@1073.4]
  wire [5:0] _T_55442; // @[Modules.scala 150:103:@1074.4]
  wire [5:0] _T_55443; // @[Modules.scala 150:103:@1075.4]
  wire [5:0] _T_55445; // @[Modules.scala 150:74:@1077.4]
  wire [5:0] _T_55447; // @[Modules.scala 151:80:@1078.4]
  wire [6:0] _T_55448; // @[Modules.scala 150:103:@1079.4]
  wire [5:0] _T_55449; // @[Modules.scala 150:103:@1080.4]
  wire [5:0] _T_55450; // @[Modules.scala 150:103:@1081.4]
  wire [5:0] _T_55452; // @[Modules.scala 150:74:@1083.4]
  wire [5:0] _T_55454; // @[Modules.scala 151:80:@1084.4]
  wire [6:0] _T_55455; // @[Modules.scala 150:103:@1085.4]
  wire [5:0] _T_55456; // @[Modules.scala 150:103:@1086.4]
  wire [5:0] _T_55457; // @[Modules.scala 150:103:@1087.4]
  wire [5:0] _T_55459; // @[Modules.scala 150:74:@1089.4]
  wire [4:0] _T_55461; // @[Modules.scala 151:80:@1090.4]
  wire [5:0] _GEN_50; // @[Modules.scala 150:103:@1091.4]
  wire [6:0] _T_55462; // @[Modules.scala 150:103:@1091.4]
  wire [5:0] _T_55463; // @[Modules.scala 150:103:@1092.4]
  wire [5:0] _T_55464; // @[Modules.scala 150:103:@1093.4]
  wire [4:0] _T_55466; // @[Modules.scala 150:74:@1095.4]
  wire [5:0] _T_55468; // @[Modules.scala 151:80:@1096.4]
  wire [5:0] _GEN_51; // @[Modules.scala 150:103:@1097.4]
  wire [6:0] _T_55469; // @[Modules.scala 150:103:@1097.4]
  wire [5:0] _T_55470; // @[Modules.scala 150:103:@1098.4]
  wire [5:0] _T_55471; // @[Modules.scala 150:103:@1099.4]
  wire [5:0] _T_55473; // @[Modules.scala 150:74:@1101.4]
  wire [4:0] _T_55475; // @[Modules.scala 151:80:@1102.4]
  wire [5:0] _GEN_52; // @[Modules.scala 150:103:@1103.4]
  wire [6:0] _T_55476; // @[Modules.scala 150:103:@1103.4]
  wire [5:0] _T_55477; // @[Modules.scala 150:103:@1104.4]
  wire [5:0] _T_55478; // @[Modules.scala 150:103:@1105.4]
  wire [5:0] _T_55480; // @[Modules.scala 150:74:@1107.4]
  wire [5:0] _T_55482; // @[Modules.scala 151:80:@1108.4]
  wire [6:0] _T_55483; // @[Modules.scala 150:103:@1109.4]
  wire [5:0] _T_55484; // @[Modules.scala 150:103:@1110.4]
  wire [5:0] _T_55485; // @[Modules.scala 150:103:@1111.4]
  wire [4:0] _T_55487; // @[Modules.scala 150:74:@1113.4]
  wire [5:0] _T_55489; // @[Modules.scala 151:80:@1114.4]
  wire [5:0] _GEN_53; // @[Modules.scala 150:103:@1115.4]
  wire [6:0] _T_55490; // @[Modules.scala 150:103:@1115.4]
  wire [5:0] _T_55491; // @[Modules.scala 150:103:@1116.4]
  wire [5:0] _T_55492; // @[Modules.scala 150:103:@1117.4]
  wire [5:0] _T_55494; // @[Modules.scala 150:74:@1119.4]
  wire [5:0] _T_55496; // @[Modules.scala 151:80:@1120.4]
  wire [6:0] _T_55497; // @[Modules.scala 150:103:@1121.4]
  wire [5:0] _T_55498; // @[Modules.scala 150:103:@1122.4]
  wire [5:0] _T_55499; // @[Modules.scala 150:103:@1123.4]
  wire [5:0] _T_55501; // @[Modules.scala 150:74:@1125.4]
  wire [4:0] _T_55503; // @[Modules.scala 151:80:@1126.4]
  wire [5:0] _GEN_54; // @[Modules.scala 150:103:@1127.4]
  wire [6:0] _T_55504; // @[Modules.scala 150:103:@1127.4]
  wire [5:0] _T_55505; // @[Modules.scala 150:103:@1128.4]
  wire [5:0] _T_55506; // @[Modules.scala 150:103:@1129.4]
  wire [5:0] _T_55508; // @[Modules.scala 150:74:@1131.4]
  wire [5:0] _T_55510; // @[Modules.scala 151:80:@1132.4]
  wire [6:0] _T_55511; // @[Modules.scala 150:103:@1133.4]
  wire [5:0] _T_55512; // @[Modules.scala 150:103:@1134.4]
  wire [5:0] _T_55513; // @[Modules.scala 150:103:@1135.4]
  wire [5:0] _T_55515; // @[Modules.scala 150:74:@1137.4]
  wire [5:0] _T_55517; // @[Modules.scala 151:80:@1138.4]
  wire [6:0] _T_55518; // @[Modules.scala 150:103:@1139.4]
  wire [5:0] _T_55519; // @[Modules.scala 150:103:@1140.4]
  wire [5:0] _T_55520; // @[Modules.scala 150:103:@1141.4]
  wire [5:0] _T_55522; // @[Modules.scala 150:74:@1143.4]
  wire [5:0] _T_55524; // @[Modules.scala 151:80:@1144.4]
  wire [6:0] _T_55525; // @[Modules.scala 150:103:@1145.4]
  wire [5:0] _T_55526; // @[Modules.scala 150:103:@1146.4]
  wire [5:0] _T_55527; // @[Modules.scala 150:103:@1147.4]
  wire [4:0] _T_55529; // @[Modules.scala 150:74:@1149.4]
  wire [4:0] _T_55531; // @[Modules.scala 151:80:@1150.4]
  wire [5:0] _T_55532; // @[Modules.scala 150:103:@1151.4]
  wire [4:0] _T_55533; // @[Modules.scala 150:103:@1152.4]
  wire [4:0] _T_55534; // @[Modules.scala 150:103:@1153.4]
  wire [4:0] _T_55536; // @[Modules.scala 150:74:@1155.4]
  wire [5:0] _T_55538; // @[Modules.scala 151:80:@1156.4]
  wire [5:0] _GEN_55; // @[Modules.scala 150:103:@1157.4]
  wire [6:0] _T_55539; // @[Modules.scala 150:103:@1157.4]
  wire [5:0] _T_55540; // @[Modules.scala 150:103:@1158.4]
  wire [5:0] _T_55541; // @[Modules.scala 150:103:@1159.4]
  wire [5:0] _T_55543; // @[Modules.scala 150:74:@1161.4]
  wire [5:0] _T_55545; // @[Modules.scala 151:80:@1162.4]
  wire [6:0] _T_55546; // @[Modules.scala 150:103:@1163.4]
  wire [5:0] _T_55547; // @[Modules.scala 150:103:@1164.4]
  wire [5:0] _T_55548; // @[Modules.scala 150:103:@1165.4]
  wire [5:0] _T_55550; // @[Modules.scala 150:74:@1167.4]
  wire [5:0] _T_55552; // @[Modules.scala 151:80:@1168.4]
  wire [6:0] _T_55553; // @[Modules.scala 150:103:@1169.4]
  wire [5:0] _T_55554; // @[Modules.scala 150:103:@1170.4]
  wire [5:0] _T_55555; // @[Modules.scala 150:103:@1171.4]
  wire [5:0] _T_55557; // @[Modules.scala 150:74:@1173.4]
  wire [4:0] _T_55559; // @[Modules.scala 151:80:@1174.4]
  wire [5:0] _GEN_56; // @[Modules.scala 150:103:@1175.4]
  wire [6:0] _T_55560; // @[Modules.scala 150:103:@1175.4]
  wire [5:0] _T_55561; // @[Modules.scala 150:103:@1176.4]
  wire [5:0] _T_55562; // @[Modules.scala 150:103:@1177.4]
  wire [5:0] _T_55564; // @[Modules.scala 150:74:@1179.4]
  wire [5:0] _T_55566; // @[Modules.scala 151:80:@1180.4]
  wire [6:0] _T_55567; // @[Modules.scala 150:103:@1181.4]
  wire [5:0] _T_55568; // @[Modules.scala 150:103:@1182.4]
  wire [5:0] _T_55569; // @[Modules.scala 150:103:@1183.4]
  wire [5:0] _T_55571; // @[Modules.scala 150:74:@1185.4]
  wire [5:0] _T_55573; // @[Modules.scala 151:80:@1186.4]
  wire [6:0] _T_55574; // @[Modules.scala 150:103:@1187.4]
  wire [5:0] _T_55575; // @[Modules.scala 150:103:@1188.4]
  wire [5:0] _T_55576; // @[Modules.scala 150:103:@1189.4]
  wire [5:0] _T_55578; // @[Modules.scala 150:74:@1191.4]
  wire [4:0] _T_55580; // @[Modules.scala 151:80:@1192.4]
  wire [5:0] _GEN_57; // @[Modules.scala 150:103:@1193.4]
  wire [6:0] _T_55581; // @[Modules.scala 150:103:@1193.4]
  wire [5:0] _T_55582; // @[Modules.scala 150:103:@1194.4]
  wire [5:0] _T_55583; // @[Modules.scala 150:103:@1195.4]
  wire [4:0] _T_55585; // @[Modules.scala 150:74:@1197.4]
  wire [5:0] _T_55587; // @[Modules.scala 151:80:@1198.4]
  wire [5:0] _GEN_58; // @[Modules.scala 150:103:@1199.4]
  wire [6:0] _T_55588; // @[Modules.scala 150:103:@1199.4]
  wire [5:0] _T_55589; // @[Modules.scala 150:103:@1200.4]
  wire [5:0] _T_55590; // @[Modules.scala 150:103:@1201.4]
  wire [5:0] _T_55592; // @[Modules.scala 150:74:@1203.4]
  wire [5:0] _T_55594; // @[Modules.scala 151:80:@1204.4]
  wire [6:0] _T_55595; // @[Modules.scala 150:103:@1205.4]
  wire [5:0] _T_55596; // @[Modules.scala 150:103:@1206.4]
  wire [5:0] _T_55597; // @[Modules.scala 150:103:@1207.4]
  wire [5:0] _T_55599; // @[Modules.scala 150:74:@1209.4]
  wire [5:0] _T_55601; // @[Modules.scala 151:80:@1210.4]
  wire [6:0] _T_55602; // @[Modules.scala 150:103:@1211.4]
  wire [5:0] _T_55603; // @[Modules.scala 150:103:@1212.4]
  wire [5:0] _T_55604; // @[Modules.scala 150:103:@1213.4]
  wire [5:0] _T_55606; // @[Modules.scala 150:74:@1215.4]
  wire [4:0] _T_55608; // @[Modules.scala 151:80:@1216.4]
  wire [5:0] _GEN_59; // @[Modules.scala 150:103:@1217.4]
  wire [6:0] _T_55609; // @[Modules.scala 150:103:@1217.4]
  wire [5:0] _T_55610; // @[Modules.scala 150:103:@1218.4]
  wire [5:0] _T_55611; // @[Modules.scala 150:103:@1219.4]
  wire [4:0] _T_55613; // @[Modules.scala 150:74:@1221.4]
  wire [5:0] _T_55615; // @[Modules.scala 151:80:@1222.4]
  wire [5:0] _GEN_60; // @[Modules.scala 150:103:@1223.4]
  wire [6:0] _T_55616; // @[Modules.scala 150:103:@1223.4]
  wire [5:0] _T_55617; // @[Modules.scala 150:103:@1224.4]
  wire [5:0] _T_55618; // @[Modules.scala 150:103:@1225.4]
  wire [5:0] _T_55620; // @[Modules.scala 150:74:@1227.4]
  wire [5:0] _T_55622; // @[Modules.scala 151:80:@1228.4]
  wire [6:0] _T_55623; // @[Modules.scala 150:103:@1229.4]
  wire [5:0] _T_55624; // @[Modules.scala 150:103:@1230.4]
  wire [5:0] _T_55625; // @[Modules.scala 150:103:@1231.4]
  wire [5:0] _T_55627; // @[Modules.scala 150:74:@1233.4]
  wire [5:0] _T_55629; // @[Modules.scala 151:80:@1234.4]
  wire [6:0] _T_55630; // @[Modules.scala 150:103:@1235.4]
  wire [5:0] _T_55631; // @[Modules.scala 150:103:@1236.4]
  wire [5:0] _T_55632; // @[Modules.scala 150:103:@1237.4]
  wire [5:0] _T_55634; // @[Modules.scala 150:74:@1239.4]
  wire [5:0] _T_55636; // @[Modules.scala 151:80:@1240.4]
  wire [6:0] _T_55637; // @[Modules.scala 150:103:@1241.4]
  wire [5:0] _T_55638; // @[Modules.scala 150:103:@1242.4]
  wire [5:0] _T_55639; // @[Modules.scala 150:103:@1243.4]
  wire [5:0] _T_55641; // @[Modules.scala 150:74:@1245.4]
  wire [5:0] _T_55643; // @[Modules.scala 151:80:@1246.4]
  wire [6:0] _T_55644; // @[Modules.scala 150:103:@1247.4]
  wire [5:0] _T_55645; // @[Modules.scala 150:103:@1248.4]
  wire [5:0] _T_55646; // @[Modules.scala 150:103:@1249.4]
  wire [4:0] _T_55648; // @[Modules.scala 150:74:@1251.4]
  wire [5:0] _T_55650; // @[Modules.scala 151:80:@1252.4]
  wire [5:0] _GEN_61; // @[Modules.scala 150:103:@1253.4]
  wire [6:0] _T_55651; // @[Modules.scala 150:103:@1253.4]
  wire [5:0] _T_55652; // @[Modules.scala 150:103:@1254.4]
  wire [5:0] _T_55653; // @[Modules.scala 150:103:@1255.4]
  wire [5:0] _T_55655; // @[Modules.scala 150:74:@1257.4]
  wire [5:0] _T_55657; // @[Modules.scala 151:80:@1258.4]
  wire [6:0] _T_55658; // @[Modules.scala 150:103:@1259.4]
  wire [5:0] _T_55659; // @[Modules.scala 150:103:@1260.4]
  wire [5:0] _T_55660; // @[Modules.scala 150:103:@1261.4]
  wire [5:0] _T_55662; // @[Modules.scala 150:74:@1263.4]
  wire [5:0] _T_55664; // @[Modules.scala 151:80:@1264.4]
  wire [6:0] _T_55665; // @[Modules.scala 150:103:@1265.4]
  wire [5:0] _T_55666; // @[Modules.scala 150:103:@1266.4]
  wire [5:0] _T_55667; // @[Modules.scala 150:103:@1267.4]
  wire [5:0] _T_55669; // @[Modules.scala 150:74:@1269.4]
  wire [5:0] _T_55671; // @[Modules.scala 151:80:@1270.4]
  wire [6:0] _T_55672; // @[Modules.scala 150:103:@1271.4]
  wire [5:0] _T_55673; // @[Modules.scala 150:103:@1272.4]
  wire [5:0] _T_55674; // @[Modules.scala 150:103:@1273.4]
  wire [5:0] _T_55676; // @[Modules.scala 150:74:@1275.4]
  wire [5:0] _T_55678; // @[Modules.scala 151:80:@1276.4]
  wire [6:0] _T_55679; // @[Modules.scala 150:103:@1277.4]
  wire [5:0] _T_55680; // @[Modules.scala 150:103:@1278.4]
  wire [5:0] _T_55681; // @[Modules.scala 150:103:@1279.4]
  wire [5:0] _T_55683; // @[Modules.scala 150:74:@1281.4]
  wire [5:0] _T_55685; // @[Modules.scala 151:80:@1282.4]
  wire [6:0] _T_55686; // @[Modules.scala 150:103:@1283.4]
  wire [5:0] _T_55687; // @[Modules.scala 150:103:@1284.4]
  wire [5:0] _T_55688; // @[Modules.scala 150:103:@1285.4]
  wire [5:0] _T_55690; // @[Modules.scala 150:74:@1287.4]
  wire [5:0] _T_55692; // @[Modules.scala 151:80:@1288.4]
  wire [6:0] _T_55693; // @[Modules.scala 150:103:@1289.4]
  wire [5:0] _T_55694; // @[Modules.scala 150:103:@1290.4]
  wire [5:0] _T_55695; // @[Modules.scala 150:103:@1291.4]
  wire [5:0] _T_55697; // @[Modules.scala 150:74:@1293.4]
  wire [5:0] _T_55699; // @[Modules.scala 151:80:@1294.4]
  wire [6:0] _T_55700; // @[Modules.scala 150:103:@1295.4]
  wire [5:0] _T_55701; // @[Modules.scala 150:103:@1296.4]
  wire [5:0] _T_55702; // @[Modules.scala 150:103:@1297.4]
  wire [5:0] _T_55704; // @[Modules.scala 150:74:@1299.4]
  wire [5:0] _T_55706; // @[Modules.scala 151:80:@1300.4]
  wire [6:0] _T_55707; // @[Modules.scala 150:103:@1301.4]
  wire [5:0] _T_55708; // @[Modules.scala 150:103:@1302.4]
  wire [5:0] _T_55709; // @[Modules.scala 150:103:@1303.4]
  wire [5:0] _T_55711; // @[Modules.scala 150:74:@1305.4]
  wire [5:0] _T_55713; // @[Modules.scala 151:80:@1306.4]
  wire [6:0] _T_55714; // @[Modules.scala 150:103:@1307.4]
  wire [5:0] _T_55715; // @[Modules.scala 150:103:@1308.4]
  wire [5:0] _T_55716; // @[Modules.scala 150:103:@1309.4]
  wire [5:0] _T_55718; // @[Modules.scala 150:74:@1311.4]
  wire [5:0] _T_55720; // @[Modules.scala 151:80:@1312.4]
  wire [6:0] _T_55721; // @[Modules.scala 150:103:@1313.4]
  wire [5:0] _T_55722; // @[Modules.scala 150:103:@1314.4]
  wire [5:0] _T_55723; // @[Modules.scala 150:103:@1315.4]
  wire [4:0] _T_55725; // @[Modules.scala 150:74:@1317.4]
  wire [5:0] _T_55727; // @[Modules.scala 151:80:@1318.4]
  wire [5:0] _GEN_62; // @[Modules.scala 150:103:@1319.4]
  wire [6:0] _T_55728; // @[Modules.scala 150:103:@1319.4]
  wire [5:0] _T_55729; // @[Modules.scala 150:103:@1320.4]
  wire [5:0] _T_55730; // @[Modules.scala 150:103:@1321.4]
  wire [5:0] _T_55732; // @[Modules.scala 150:74:@1323.4]
  wire [5:0] _T_55734; // @[Modules.scala 151:80:@1324.4]
  wire [6:0] _T_55735; // @[Modules.scala 150:103:@1325.4]
  wire [5:0] _T_55736; // @[Modules.scala 150:103:@1326.4]
  wire [5:0] _T_55737; // @[Modules.scala 150:103:@1327.4]
  wire [5:0] _T_55739; // @[Modules.scala 150:74:@1329.4]
  wire [5:0] _T_55741; // @[Modules.scala 151:80:@1330.4]
  wire [6:0] _T_55742; // @[Modules.scala 150:103:@1331.4]
  wire [5:0] _T_55743; // @[Modules.scala 150:103:@1332.4]
  wire [5:0] _T_55744; // @[Modules.scala 150:103:@1333.4]
  wire [5:0] _T_55746; // @[Modules.scala 150:74:@1335.4]
  wire [5:0] _T_55748; // @[Modules.scala 151:80:@1336.4]
  wire [6:0] _T_55749; // @[Modules.scala 150:103:@1337.4]
  wire [5:0] _T_55750; // @[Modules.scala 150:103:@1338.4]
  wire [5:0] _T_55751; // @[Modules.scala 150:103:@1339.4]
  wire [5:0] _T_55753; // @[Modules.scala 150:74:@1341.4]
  wire [5:0] _T_55755; // @[Modules.scala 151:80:@1342.4]
  wire [6:0] _T_55756; // @[Modules.scala 150:103:@1343.4]
  wire [5:0] _T_55757; // @[Modules.scala 150:103:@1344.4]
  wire [5:0] _T_55758; // @[Modules.scala 150:103:@1345.4]
  wire [5:0] _T_55760; // @[Modules.scala 150:74:@1347.4]
  wire [5:0] _T_55762; // @[Modules.scala 151:80:@1348.4]
  wire [6:0] _T_55763; // @[Modules.scala 150:103:@1349.4]
  wire [5:0] _T_55764; // @[Modules.scala 150:103:@1350.4]
  wire [5:0] _T_55765; // @[Modules.scala 150:103:@1351.4]
  wire [5:0] _T_55767; // @[Modules.scala 150:74:@1353.4]
  wire [4:0] _T_55769; // @[Modules.scala 151:80:@1354.4]
  wire [5:0] _GEN_63; // @[Modules.scala 150:103:@1355.4]
  wire [6:0] _T_55770; // @[Modules.scala 150:103:@1355.4]
  wire [5:0] _T_55771; // @[Modules.scala 150:103:@1356.4]
  wire [5:0] _T_55772; // @[Modules.scala 150:103:@1357.4]
  wire [4:0] _T_55774; // @[Modules.scala 150:74:@1359.4]
  wire [5:0] _T_55776; // @[Modules.scala 151:80:@1360.4]
  wire [5:0] _GEN_64; // @[Modules.scala 150:103:@1361.4]
  wire [6:0] _T_55777; // @[Modules.scala 150:103:@1361.4]
  wire [5:0] _T_55778; // @[Modules.scala 150:103:@1362.4]
  wire [5:0] _T_55779; // @[Modules.scala 150:103:@1363.4]
  wire [5:0] _T_55781; // @[Modules.scala 150:74:@1365.4]
  wire [5:0] _T_55783; // @[Modules.scala 151:80:@1366.4]
  wire [6:0] _T_55784; // @[Modules.scala 150:103:@1367.4]
  wire [5:0] _T_55785; // @[Modules.scala 150:103:@1368.4]
  wire [5:0] _T_55786; // @[Modules.scala 150:103:@1369.4]
  wire [5:0] _T_55788; // @[Modules.scala 150:74:@1371.4]
  wire [5:0] _T_55790; // @[Modules.scala 151:80:@1372.4]
  wire [6:0] _T_55791; // @[Modules.scala 150:103:@1373.4]
  wire [5:0] _T_55792; // @[Modules.scala 150:103:@1374.4]
  wire [5:0] _T_55793; // @[Modules.scala 150:103:@1375.4]
  wire [5:0] _T_55795; // @[Modules.scala 150:74:@1377.4]
  wire [5:0] _T_55797; // @[Modules.scala 151:80:@1378.4]
  wire [6:0] _T_55798; // @[Modules.scala 150:103:@1379.4]
  wire [5:0] _T_55799; // @[Modules.scala 150:103:@1380.4]
  wire [5:0] _T_55800; // @[Modules.scala 150:103:@1381.4]
  wire [5:0] _T_55802; // @[Modules.scala 150:74:@1383.4]
  wire [5:0] _T_55804; // @[Modules.scala 151:80:@1384.4]
  wire [6:0] _T_55805; // @[Modules.scala 150:103:@1385.4]
  wire [5:0] _T_55806; // @[Modules.scala 150:103:@1386.4]
  wire [5:0] _T_55807; // @[Modules.scala 150:103:@1387.4]
  wire [5:0] _T_55809; // @[Modules.scala 150:74:@1389.4]
  wire [5:0] _T_55811; // @[Modules.scala 151:80:@1390.4]
  wire [6:0] _T_55812; // @[Modules.scala 150:103:@1391.4]
  wire [5:0] _T_55813; // @[Modules.scala 150:103:@1392.4]
  wire [5:0] _T_55814; // @[Modules.scala 150:103:@1393.4]
  wire [5:0] _T_55816; // @[Modules.scala 150:74:@1395.4]
  wire [5:0] _T_55818; // @[Modules.scala 151:80:@1396.4]
  wire [6:0] _T_55819; // @[Modules.scala 150:103:@1397.4]
  wire [5:0] _T_55820; // @[Modules.scala 150:103:@1398.4]
  wire [5:0] _T_55821; // @[Modules.scala 150:103:@1399.4]
  wire [5:0] _T_55823; // @[Modules.scala 150:74:@1401.4]
  wire [5:0] _T_55825; // @[Modules.scala 151:80:@1402.4]
  wire [6:0] _T_55826; // @[Modules.scala 150:103:@1403.4]
  wire [5:0] _T_55827; // @[Modules.scala 150:103:@1404.4]
  wire [5:0] _T_55828; // @[Modules.scala 150:103:@1405.4]
  wire [5:0] _T_55830; // @[Modules.scala 150:74:@1407.4]
  wire [5:0] _T_55832; // @[Modules.scala 151:80:@1408.4]
  wire [6:0] _T_55833; // @[Modules.scala 150:103:@1409.4]
  wire [5:0] _T_55834; // @[Modules.scala 150:103:@1410.4]
  wire [5:0] _T_55835; // @[Modules.scala 150:103:@1411.4]
  wire [4:0] _T_55837; // @[Modules.scala 150:74:@1413.4]
  wire [5:0] _T_55839; // @[Modules.scala 151:80:@1414.4]
  wire [5:0] _GEN_65; // @[Modules.scala 150:103:@1415.4]
  wire [6:0] _T_55840; // @[Modules.scala 150:103:@1415.4]
  wire [5:0] _T_55841; // @[Modules.scala 150:103:@1416.4]
  wire [5:0] _T_55842; // @[Modules.scala 150:103:@1417.4]
  wire [5:0] _T_55844; // @[Modules.scala 150:74:@1419.4]
  wire [5:0] _T_55846; // @[Modules.scala 151:80:@1420.4]
  wire [6:0] _T_55847; // @[Modules.scala 150:103:@1421.4]
  wire [5:0] _T_55848; // @[Modules.scala 150:103:@1422.4]
  wire [5:0] _T_55849; // @[Modules.scala 150:103:@1423.4]
  wire [5:0] _T_55851; // @[Modules.scala 150:74:@1425.4]
  wire [5:0] _T_55853; // @[Modules.scala 151:80:@1426.4]
  wire [6:0] _T_55854; // @[Modules.scala 150:103:@1427.4]
  wire [5:0] _T_55855; // @[Modules.scala 150:103:@1428.4]
  wire [5:0] _T_55856; // @[Modules.scala 150:103:@1429.4]
  wire [5:0] _T_55858; // @[Modules.scala 150:74:@1431.4]
  wire [5:0] _T_55860; // @[Modules.scala 151:80:@1432.4]
  wire [6:0] _T_55861; // @[Modules.scala 150:103:@1433.4]
  wire [5:0] _T_55862; // @[Modules.scala 150:103:@1434.4]
  wire [5:0] _T_55863; // @[Modules.scala 150:103:@1435.4]
  wire [5:0] _T_55865; // @[Modules.scala 150:74:@1437.4]
  wire [5:0] _T_55867; // @[Modules.scala 151:80:@1438.4]
  wire [6:0] _T_55868; // @[Modules.scala 150:103:@1439.4]
  wire [5:0] _T_55869; // @[Modules.scala 150:103:@1440.4]
  wire [5:0] _T_55870; // @[Modules.scala 150:103:@1441.4]
  wire [5:0] _T_55872; // @[Modules.scala 150:74:@1443.4]
  wire [5:0] _T_55874; // @[Modules.scala 151:80:@1444.4]
  wire [6:0] _T_55875; // @[Modules.scala 150:103:@1445.4]
  wire [5:0] _T_55876; // @[Modules.scala 150:103:@1446.4]
  wire [5:0] _T_55877; // @[Modules.scala 150:103:@1447.4]
  wire [5:0] _T_55879; // @[Modules.scala 150:74:@1449.4]
  wire [5:0] _T_55881; // @[Modules.scala 151:80:@1450.4]
  wire [6:0] _T_55882; // @[Modules.scala 150:103:@1451.4]
  wire [5:0] _T_55883; // @[Modules.scala 150:103:@1452.4]
  wire [5:0] _T_55884; // @[Modules.scala 150:103:@1453.4]
  wire [4:0] _T_55886; // @[Modules.scala 150:74:@1455.4]
  wire [5:0] _T_55888; // @[Modules.scala 151:80:@1456.4]
  wire [5:0] _GEN_66; // @[Modules.scala 150:103:@1457.4]
  wire [6:0] _T_55889; // @[Modules.scala 150:103:@1457.4]
  wire [5:0] _T_55890; // @[Modules.scala 150:103:@1458.4]
  wire [5:0] _T_55891; // @[Modules.scala 150:103:@1459.4]
  wire [4:0] _T_55893; // @[Modules.scala 150:74:@1461.4]
  wire [4:0] _T_55895; // @[Modules.scala 151:80:@1462.4]
  wire [5:0] _T_55896; // @[Modules.scala 150:103:@1463.4]
  wire [4:0] _T_55897; // @[Modules.scala 150:103:@1464.4]
  wire [4:0] _T_55898; // @[Modules.scala 150:103:@1465.4]
  wire [4:0] _T_55900; // @[Modules.scala 150:74:@1467.4]
  wire [4:0] _T_55902; // @[Modules.scala 151:80:@1468.4]
  wire [5:0] _T_55903; // @[Modules.scala 150:103:@1469.4]
  wire [4:0] _T_55904; // @[Modules.scala 150:103:@1470.4]
  wire [4:0] _T_55905; // @[Modules.scala 150:103:@1471.4]
  wire [4:0] _T_55907; // @[Modules.scala 150:74:@1473.4]
  wire [4:0] _T_55909; // @[Modules.scala 151:80:@1474.4]
  wire [5:0] _T_55910; // @[Modules.scala 150:103:@1475.4]
  wire [4:0] _T_55911; // @[Modules.scala 150:103:@1476.4]
  wire [4:0] _T_55912; // @[Modules.scala 150:103:@1477.4]
  wire [4:0] _T_55914; // @[Modules.scala 150:74:@1479.4]
  wire [4:0] _T_55916; // @[Modules.scala 151:80:@1480.4]
  wire [5:0] _T_55917; // @[Modules.scala 150:103:@1481.4]
  wire [4:0] _T_55918; // @[Modules.scala 150:103:@1482.4]
  wire [4:0] _T_55919; // @[Modules.scala 150:103:@1483.4]
  wire [5:0] _T_55921; // @[Modules.scala 150:74:@1485.4]
  wire [5:0] _T_55923; // @[Modules.scala 151:80:@1486.4]
  wire [6:0] _T_55924; // @[Modules.scala 150:103:@1487.4]
  wire [5:0] _T_55925; // @[Modules.scala 150:103:@1488.4]
  wire [5:0] _T_55926; // @[Modules.scala 150:103:@1489.4]
  wire [5:0] _T_55928; // @[Modules.scala 150:74:@1491.4]
  wire [5:0] _T_55930; // @[Modules.scala 151:80:@1492.4]
  wire [6:0] _T_55931; // @[Modules.scala 150:103:@1493.4]
  wire [5:0] _T_55932; // @[Modules.scala 150:103:@1494.4]
  wire [5:0] _T_55933; // @[Modules.scala 150:103:@1495.4]
  wire [5:0] _T_55935; // @[Modules.scala 150:74:@1497.4]
  wire [5:0] _T_55937; // @[Modules.scala 151:80:@1498.4]
  wire [6:0] _T_55938; // @[Modules.scala 150:103:@1499.4]
  wire [5:0] _T_55939; // @[Modules.scala 150:103:@1500.4]
  wire [5:0] _T_55940; // @[Modules.scala 150:103:@1501.4]
  wire [5:0] _T_55942; // @[Modules.scala 150:74:@1503.4]
  wire [5:0] _T_55944; // @[Modules.scala 151:80:@1504.4]
  wire [6:0] _T_55945; // @[Modules.scala 150:103:@1505.4]
  wire [5:0] _T_55946; // @[Modules.scala 150:103:@1506.4]
  wire [5:0] _T_55947; // @[Modules.scala 150:103:@1507.4]
  wire [5:0] _T_55949; // @[Modules.scala 150:74:@1509.4]
  wire [5:0] _T_55951; // @[Modules.scala 151:80:@1510.4]
  wire [6:0] _T_55952; // @[Modules.scala 150:103:@1511.4]
  wire [5:0] _T_55953; // @[Modules.scala 150:103:@1512.4]
  wire [5:0] _T_55954; // @[Modules.scala 150:103:@1513.4]
  wire [5:0] _T_55956; // @[Modules.scala 150:74:@1515.4]
  wire [5:0] _T_55958; // @[Modules.scala 151:80:@1516.4]
  wire [6:0] _T_55959; // @[Modules.scala 150:103:@1517.4]
  wire [5:0] _T_55960; // @[Modules.scala 150:103:@1518.4]
  wire [5:0] _T_55961; // @[Modules.scala 150:103:@1519.4]
  wire [5:0] _T_55963; // @[Modules.scala 150:74:@1521.4]
  wire [5:0] _T_55965; // @[Modules.scala 151:80:@1522.4]
  wire [6:0] _T_55966; // @[Modules.scala 150:103:@1523.4]
  wire [5:0] _T_55967; // @[Modules.scala 150:103:@1524.4]
  wire [5:0] _T_55968; // @[Modules.scala 150:103:@1525.4]
  wire [4:0] _T_55970; // @[Modules.scala 150:74:@1527.4]
  wire [4:0] _T_55972; // @[Modules.scala 151:80:@1528.4]
  wire [5:0] _T_55973; // @[Modules.scala 150:103:@1529.4]
  wire [4:0] _T_55974; // @[Modules.scala 150:103:@1530.4]
  wire [4:0] _T_55975; // @[Modules.scala 150:103:@1531.4]
  wire [4:0] _T_55977; // @[Modules.scala 150:74:@1533.4]
  wire [4:0] _T_55979; // @[Modules.scala 151:80:@1534.4]
  wire [5:0] _T_55980; // @[Modules.scala 150:103:@1535.4]
  wire [4:0] _T_55981; // @[Modules.scala 150:103:@1536.4]
  wire [4:0] _T_55982; // @[Modules.scala 150:103:@1537.4]
  wire [4:0] _T_55984; // @[Modules.scala 150:74:@1539.4]
  wire [4:0] _T_55986; // @[Modules.scala 151:80:@1540.4]
  wire [5:0] _T_55987; // @[Modules.scala 150:103:@1541.4]
  wire [4:0] _T_55988; // @[Modules.scala 150:103:@1542.4]
  wire [4:0] _T_55989; // @[Modules.scala 150:103:@1543.4]
  wire [4:0] _T_55991; // @[Modules.scala 150:74:@1545.4]
  wire [4:0] _T_55993; // @[Modules.scala 151:80:@1546.4]
  wire [5:0] _T_55994; // @[Modules.scala 150:103:@1547.4]
  wire [4:0] _T_55995; // @[Modules.scala 150:103:@1548.4]
  wire [4:0] _T_55996; // @[Modules.scala 150:103:@1549.4]
  wire [4:0] _T_55998; // @[Modules.scala 150:74:@1551.4]
  wire [4:0] _T_56000; // @[Modules.scala 151:80:@1552.4]
  wire [5:0] _T_56001; // @[Modules.scala 150:103:@1553.4]
  wire [4:0] _T_56002; // @[Modules.scala 150:103:@1554.4]
  wire [4:0] _T_56003; // @[Modules.scala 150:103:@1555.4]
  wire [4:0] _T_56005; // @[Modules.scala 150:74:@1557.4]
  wire [4:0] _T_56007; // @[Modules.scala 151:80:@1558.4]
  wire [5:0] _T_56008; // @[Modules.scala 150:103:@1559.4]
  wire [4:0] _T_56009; // @[Modules.scala 150:103:@1560.4]
  wire [4:0] _T_56010; // @[Modules.scala 150:103:@1561.4]
  wire [4:0] _T_56012; // @[Modules.scala 150:74:@1563.4]
  wire [4:0] _T_56014; // @[Modules.scala 151:80:@1564.4]
  wire [5:0] _T_56015; // @[Modules.scala 150:103:@1565.4]
  wire [4:0] _T_56016; // @[Modules.scala 150:103:@1566.4]
  wire [4:0] _T_56017; // @[Modules.scala 150:103:@1567.4]
  wire [5:0] _T_56019; // @[Modules.scala 150:74:@1569.4]
  wire [5:0] _T_56021; // @[Modules.scala 151:80:@1570.4]
  wire [6:0] _T_56022; // @[Modules.scala 150:103:@1571.4]
  wire [5:0] _T_56023; // @[Modules.scala 150:103:@1572.4]
  wire [5:0] _T_56024; // @[Modules.scala 150:103:@1573.4]
  wire [5:0] _T_56026; // @[Modules.scala 150:74:@1575.4]
  wire [4:0] _T_56028; // @[Modules.scala 151:80:@1576.4]
  wire [5:0] _GEN_67; // @[Modules.scala 150:103:@1577.4]
  wire [6:0] _T_56029; // @[Modules.scala 150:103:@1577.4]
  wire [5:0] _T_56030; // @[Modules.scala 150:103:@1578.4]
  wire [5:0] _T_56031; // @[Modules.scala 150:103:@1579.4]
  wire [5:0] _T_56033; // @[Modules.scala 150:74:@1581.4]
  wire [5:0] _T_56035; // @[Modules.scala 151:80:@1582.4]
  wire [6:0] _T_56036; // @[Modules.scala 150:103:@1583.4]
  wire [5:0] _T_56037; // @[Modules.scala 150:103:@1584.4]
  wire [5:0] _T_56038; // @[Modules.scala 150:103:@1585.4]
  wire [5:0] _T_56040; // @[Modules.scala 150:74:@1587.4]
  wire [5:0] _T_56042; // @[Modules.scala 151:80:@1588.4]
  wire [6:0] _T_56043; // @[Modules.scala 150:103:@1589.4]
  wire [5:0] _T_56044; // @[Modules.scala 150:103:@1590.4]
  wire [5:0] _T_56045; // @[Modules.scala 150:103:@1591.4]
  wire [5:0] _T_56047; // @[Modules.scala 150:74:@1593.4]
  wire [4:0] _T_56049; // @[Modules.scala 151:80:@1594.4]
  wire [5:0] _GEN_68; // @[Modules.scala 150:103:@1595.4]
  wire [6:0] _T_56050; // @[Modules.scala 150:103:@1595.4]
  wire [5:0] _T_56051; // @[Modules.scala 150:103:@1596.4]
  wire [5:0] _T_56052; // @[Modules.scala 150:103:@1597.4]
  wire [4:0] _T_56054; // @[Modules.scala 150:74:@1599.4]
  wire [4:0] _T_56056; // @[Modules.scala 151:80:@1600.4]
  wire [5:0] _T_56057; // @[Modules.scala 150:103:@1601.4]
  wire [4:0] _T_56058; // @[Modules.scala 150:103:@1602.4]
  wire [4:0] _T_56059; // @[Modules.scala 150:103:@1603.4]
  wire [4:0] _T_56061; // @[Modules.scala 150:74:@1605.4]
  wire [4:0] _T_56063; // @[Modules.scala 151:80:@1606.4]
  wire [5:0] _T_56064; // @[Modules.scala 150:103:@1607.4]
  wire [4:0] _T_56065; // @[Modules.scala 150:103:@1608.4]
  wire [4:0] _T_56066; // @[Modules.scala 150:103:@1609.4]
  wire [4:0] _T_56068; // @[Modules.scala 150:74:@1611.4]
  wire [4:0] _T_56070; // @[Modules.scala 151:80:@1612.4]
  wire [5:0] _T_56071; // @[Modules.scala 150:103:@1613.4]
  wire [4:0] _T_56072; // @[Modules.scala 150:103:@1614.4]
  wire [4:0] _T_56073; // @[Modules.scala 150:103:@1615.4]
  wire [4:0] _T_56075; // @[Modules.scala 150:74:@1617.4]
  wire [4:0] _T_56077; // @[Modules.scala 151:80:@1618.4]
  wire [5:0] _T_56078; // @[Modules.scala 150:103:@1619.4]
  wire [4:0] _T_56079; // @[Modules.scala 150:103:@1620.4]
  wire [4:0] _T_56080; // @[Modules.scala 150:103:@1621.4]
  wire [4:0] _T_56082; // @[Modules.scala 150:74:@1623.4]
  wire [4:0] _T_56084; // @[Modules.scala 151:80:@1624.4]
  wire [5:0] _T_56085; // @[Modules.scala 150:103:@1625.4]
  wire [4:0] _T_56086; // @[Modules.scala 150:103:@1626.4]
  wire [4:0] _T_56087; // @[Modules.scala 150:103:@1627.4]
  wire [4:0] _T_56089; // @[Modules.scala 150:74:@1629.4]
  wire [4:0] _T_56091; // @[Modules.scala 151:80:@1630.4]
  wire [5:0] _T_56092; // @[Modules.scala 150:103:@1631.4]
  wire [4:0] _T_56093; // @[Modules.scala 150:103:@1632.4]
  wire [4:0] _T_56094; // @[Modules.scala 150:103:@1633.4]
  wire [4:0] _T_56096; // @[Modules.scala 150:74:@1635.4]
  wire [5:0] _T_56098; // @[Modules.scala 151:80:@1636.4]
  wire [5:0] _GEN_69; // @[Modules.scala 150:103:@1637.4]
  wire [6:0] _T_56099; // @[Modules.scala 150:103:@1637.4]
  wire [5:0] _T_56100; // @[Modules.scala 150:103:@1638.4]
  wire [5:0] _T_56101; // @[Modules.scala 150:103:@1639.4]
  wire [5:0] _T_56103; // @[Modules.scala 150:74:@1641.4]
  wire [5:0] _T_56105; // @[Modules.scala 151:80:@1642.4]
  wire [6:0] _T_56106; // @[Modules.scala 150:103:@1643.4]
  wire [5:0] _T_56107; // @[Modules.scala 150:103:@1644.4]
  wire [5:0] _T_56108; // @[Modules.scala 150:103:@1645.4]
  wire [5:0] _T_56110; // @[Modules.scala 150:74:@1647.4]
  wire [5:0] _T_56112; // @[Modules.scala 151:80:@1648.4]
  wire [6:0] _T_56113; // @[Modules.scala 150:103:@1649.4]
  wire [5:0] _T_56114; // @[Modules.scala 150:103:@1650.4]
  wire [5:0] _T_56115; // @[Modules.scala 150:103:@1651.4]
  wire [5:0] _T_56117; // @[Modules.scala 150:74:@1653.4]
  wire [4:0] _T_56119; // @[Modules.scala 151:80:@1654.4]
  wire [5:0] _GEN_70; // @[Modules.scala 150:103:@1655.4]
  wire [6:0] _T_56120; // @[Modules.scala 150:103:@1655.4]
  wire [5:0] _T_56121; // @[Modules.scala 150:103:@1656.4]
  wire [5:0] _T_56122; // @[Modules.scala 150:103:@1657.4]
  wire [4:0] _T_56124; // @[Modules.scala 150:74:@1659.4]
  wire [5:0] _T_56126; // @[Modules.scala 151:80:@1660.4]
  wire [5:0] _GEN_71; // @[Modules.scala 150:103:@1661.4]
  wire [6:0] _T_56127; // @[Modules.scala 150:103:@1661.4]
  wire [5:0] _T_56128; // @[Modules.scala 150:103:@1662.4]
  wire [5:0] _T_56129; // @[Modules.scala 150:103:@1663.4]
  wire [5:0] _T_56131; // @[Modules.scala 150:74:@1665.4]
  wire [5:0] _T_56133; // @[Modules.scala 151:80:@1666.4]
  wire [6:0] _T_56134; // @[Modules.scala 150:103:@1667.4]
  wire [5:0] _T_56135; // @[Modules.scala 150:103:@1668.4]
  wire [5:0] _T_56136; // @[Modules.scala 150:103:@1669.4]
  wire [5:0] _T_56138; // @[Modules.scala 150:74:@1671.4]
  wire [5:0] _T_56140; // @[Modules.scala 151:80:@1672.4]
  wire [6:0] _T_56141; // @[Modules.scala 150:103:@1673.4]
  wire [5:0] _T_56142; // @[Modules.scala 150:103:@1674.4]
  wire [5:0] _T_56143; // @[Modules.scala 150:103:@1675.4]
  wire [4:0] _T_56145; // @[Modules.scala 150:74:@1677.4]
  wire [4:0] _T_56147; // @[Modules.scala 151:80:@1678.4]
  wire [5:0] _T_56148; // @[Modules.scala 150:103:@1679.4]
  wire [4:0] _T_56149; // @[Modules.scala 150:103:@1680.4]
  wire [4:0] _T_56150; // @[Modules.scala 150:103:@1681.4]
  wire [4:0] _T_56152; // @[Modules.scala 150:74:@1683.4]
  wire [4:0] _T_56154; // @[Modules.scala 151:80:@1684.4]
  wire [5:0] _T_56155; // @[Modules.scala 150:103:@1685.4]
  wire [4:0] _T_56156; // @[Modules.scala 150:103:@1686.4]
  wire [4:0] _T_56157; // @[Modules.scala 150:103:@1687.4]
  wire [4:0] _T_56159; // @[Modules.scala 150:74:@1689.4]
  wire [4:0] _T_56161; // @[Modules.scala 151:80:@1690.4]
  wire [5:0] _T_56162; // @[Modules.scala 150:103:@1691.4]
  wire [4:0] _T_56163; // @[Modules.scala 150:103:@1692.4]
  wire [4:0] _T_56164; // @[Modules.scala 150:103:@1693.4]
  wire [4:0] _T_56166; // @[Modules.scala 150:74:@1695.4]
  wire [4:0] _T_56168; // @[Modules.scala 151:80:@1696.4]
  wire [5:0] _T_56169; // @[Modules.scala 150:103:@1697.4]
  wire [4:0] _T_56170; // @[Modules.scala 150:103:@1698.4]
  wire [4:0] _T_56171; // @[Modules.scala 150:103:@1699.4]
  wire [4:0] _T_56173; // @[Modules.scala 150:74:@1701.4]
  wire [4:0] _T_56175; // @[Modules.scala 151:80:@1702.4]
  wire [5:0] _T_56176; // @[Modules.scala 150:103:@1703.4]
  wire [4:0] _T_56177; // @[Modules.scala 150:103:@1704.4]
  wire [4:0] _T_56178; // @[Modules.scala 150:103:@1705.4]
  wire [4:0] _T_56180; // @[Modules.scala 150:74:@1707.4]
  wire [4:0] _T_56182; // @[Modules.scala 151:80:@1708.4]
  wire [5:0] _T_56183; // @[Modules.scala 150:103:@1709.4]
  wire [4:0] _T_56184; // @[Modules.scala 150:103:@1710.4]
  wire [4:0] _T_56185; // @[Modules.scala 150:103:@1711.4]
  wire [4:0] _T_56187; // @[Modules.scala 150:74:@1713.4]
  wire [4:0] _T_56189; // @[Modules.scala 151:80:@1714.4]
  wire [5:0] _T_56190; // @[Modules.scala 150:103:@1715.4]
  wire [4:0] _T_56191; // @[Modules.scala 150:103:@1716.4]
  wire [4:0] _T_56192; // @[Modules.scala 150:103:@1717.4]
  wire [4:0] _T_56194; // @[Modules.scala 150:74:@1719.4]
  wire [5:0] _T_56196; // @[Modules.scala 151:80:@1720.4]
  wire [5:0] _GEN_72; // @[Modules.scala 150:103:@1721.4]
  wire [6:0] _T_56197; // @[Modules.scala 150:103:@1721.4]
  wire [5:0] _T_56198; // @[Modules.scala 150:103:@1722.4]
  wire [5:0] _T_56199; // @[Modules.scala 150:103:@1723.4]
  wire [5:0] _T_56201; // @[Modules.scala 150:74:@1725.4]
  wire [5:0] _T_56203; // @[Modules.scala 151:80:@1726.4]
  wire [6:0] _T_56204; // @[Modules.scala 150:103:@1727.4]
  wire [5:0] _T_56205; // @[Modules.scala 150:103:@1728.4]
  wire [5:0] _T_56206; // @[Modules.scala 150:103:@1729.4]
  wire [5:0] _T_56208; // @[Modules.scala 150:74:@1731.4]
  wire [5:0] _T_56210; // @[Modules.scala 151:80:@1732.4]
  wire [6:0] _T_56211; // @[Modules.scala 150:103:@1733.4]
  wire [5:0] _T_56212; // @[Modules.scala 150:103:@1734.4]
  wire [5:0] _T_56213; // @[Modules.scala 150:103:@1735.4]
  wire [4:0] _T_56215; // @[Modules.scala 150:74:@1737.4]
  wire [5:0] _T_56217; // @[Modules.scala 151:80:@1738.4]
  wire [5:0] _GEN_73; // @[Modules.scala 150:103:@1739.4]
  wire [6:0] _T_56218; // @[Modules.scala 150:103:@1739.4]
  wire [5:0] _T_56219; // @[Modules.scala 150:103:@1740.4]
  wire [5:0] _T_56220; // @[Modules.scala 150:103:@1741.4]
  wire [5:0] _T_56222; // @[Modules.scala 150:74:@1743.4]
  wire [4:0] _T_56224; // @[Modules.scala 151:80:@1744.4]
  wire [5:0] _GEN_74; // @[Modules.scala 150:103:@1745.4]
  wire [6:0] _T_56225; // @[Modules.scala 150:103:@1745.4]
  wire [5:0] _T_56226; // @[Modules.scala 150:103:@1746.4]
  wire [5:0] _T_56227; // @[Modules.scala 150:103:@1747.4]
  wire [4:0] _T_56229; // @[Modules.scala 150:74:@1749.4]
  wire [4:0] _T_56231; // @[Modules.scala 151:80:@1750.4]
  wire [5:0] _T_56232; // @[Modules.scala 150:103:@1751.4]
  wire [4:0] _T_56233; // @[Modules.scala 150:103:@1752.4]
  wire [4:0] _T_56234; // @[Modules.scala 150:103:@1753.4]
  wire [4:0] _T_56236; // @[Modules.scala 150:74:@1755.4]
  wire [4:0] _T_56238; // @[Modules.scala 151:80:@1756.4]
  wire [5:0] _T_56239; // @[Modules.scala 150:103:@1757.4]
  wire [4:0] _T_56240; // @[Modules.scala 150:103:@1758.4]
  wire [4:0] _T_56241; // @[Modules.scala 150:103:@1759.4]
  wire [4:0] _T_56243; // @[Modules.scala 150:74:@1761.4]
  wire [5:0] _T_56245; // @[Modules.scala 151:80:@1762.4]
  wire [5:0] _GEN_75; // @[Modules.scala 150:103:@1763.4]
  wire [6:0] _T_56246; // @[Modules.scala 150:103:@1763.4]
  wire [5:0] _T_56247; // @[Modules.scala 150:103:@1764.4]
  wire [5:0] _T_56248; // @[Modules.scala 150:103:@1765.4]
  wire [5:0] _T_56250; // @[Modules.scala 150:74:@1767.4]
  wire [5:0] _T_56252; // @[Modules.scala 151:80:@1768.4]
  wire [6:0] _T_56253; // @[Modules.scala 150:103:@1769.4]
  wire [5:0] _T_56254; // @[Modules.scala 150:103:@1770.4]
  wire [5:0] _T_56255; // @[Modules.scala 150:103:@1771.4]
  wire [4:0] _T_56257; // @[Modules.scala 150:74:@1773.4]
  wire [4:0] _T_56259; // @[Modules.scala 151:80:@1774.4]
  wire [5:0] _T_56260; // @[Modules.scala 150:103:@1775.4]
  wire [4:0] _T_56261; // @[Modules.scala 150:103:@1776.4]
  wire [4:0] _T_56262; // @[Modules.scala 150:103:@1777.4]
  wire [5:0] _T_56264; // @[Modules.scala 150:74:@1779.4]
  wire [5:0] _T_56266; // @[Modules.scala 151:80:@1780.4]
  wire [6:0] _T_56267; // @[Modules.scala 150:103:@1781.4]
  wire [5:0] _T_56268; // @[Modules.scala 150:103:@1782.4]
  wire [5:0] _T_56269; // @[Modules.scala 150:103:@1783.4]
  wire [5:0] _T_56271; // @[Modules.scala 150:74:@1785.4]
  wire [5:0] _T_56273; // @[Modules.scala 151:80:@1786.4]
  wire [6:0] _T_56274; // @[Modules.scala 150:103:@1787.4]
  wire [5:0] _T_56275; // @[Modules.scala 150:103:@1788.4]
  wire [5:0] _T_56276; // @[Modules.scala 150:103:@1789.4]
  wire [5:0] _T_56278; // @[Modules.scala 150:74:@1791.4]
  wire [5:0] _T_56280; // @[Modules.scala 151:80:@1792.4]
  wire [6:0] _T_56281; // @[Modules.scala 150:103:@1793.4]
  wire [5:0] _T_56282; // @[Modules.scala 150:103:@1794.4]
  wire [5:0] _T_56283; // @[Modules.scala 150:103:@1795.4]
  wire [5:0] _T_56285; // @[Modules.scala 150:74:@1797.4]
  wire [5:0] _T_56287; // @[Modules.scala 151:80:@1798.4]
  wire [6:0] _T_56288; // @[Modules.scala 150:103:@1799.4]
  wire [5:0] _T_56289; // @[Modules.scala 150:103:@1800.4]
  wire [5:0] _T_56290; // @[Modules.scala 150:103:@1801.4]
  wire [4:0] _T_56292; // @[Modules.scala 150:74:@1803.4]
  wire [4:0] _T_56294; // @[Modules.scala 151:80:@1804.4]
  wire [5:0] _T_56295; // @[Modules.scala 150:103:@1805.4]
  wire [4:0] _T_56296; // @[Modules.scala 150:103:@1806.4]
  wire [4:0] _T_56297; // @[Modules.scala 150:103:@1807.4]
  wire [5:0] _T_56299; // @[Modules.scala 150:74:@1809.4]
  wire [5:0] _T_56301; // @[Modules.scala 151:80:@1810.4]
  wire [6:0] _T_56302; // @[Modules.scala 150:103:@1811.4]
  wire [5:0] _T_56303; // @[Modules.scala 150:103:@1812.4]
  wire [5:0] _T_56304; // @[Modules.scala 150:103:@1813.4]
  wire [5:0] _T_56306; // @[Modules.scala 153:80:@1815.4]
  wire [13:0] buffer_0_0; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56307; // @[Modules.scala 160:64:@1817.4]
  wire [13:0] _T_56308; // @[Modules.scala 160:64:@1818.4]
  wire [13:0] buffer_0_302; // @[Modules.scala 160:64:@1819.4]
  wire [13:0] buffer_0_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56310; // @[Modules.scala 160:64:@1821.4]
  wire [13:0] _T_56311; // @[Modules.scala 160:64:@1822.4]
  wire [13:0] buffer_0_303; // @[Modules.scala 160:64:@1823.4]
  wire [13:0] buffer_0_4; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_5; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56313; // @[Modules.scala 160:64:@1825.4]
  wire [13:0] _T_56314; // @[Modules.scala 160:64:@1826.4]
  wire [13:0] buffer_0_304; // @[Modules.scala 160:64:@1827.4]
  wire [13:0] buffer_0_6; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_7; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56316; // @[Modules.scala 160:64:@1829.4]
  wire [13:0] _T_56317; // @[Modules.scala 160:64:@1830.4]
  wire [13:0] buffer_0_305; // @[Modules.scala 160:64:@1831.4]
  wire [13:0] buffer_0_8; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56319; // @[Modules.scala 160:64:@1833.4]
  wire [13:0] _T_56320; // @[Modules.scala 160:64:@1834.4]
  wire [13:0] buffer_0_306; // @[Modules.scala 160:64:@1835.4]
  wire [13:0] buffer_0_10; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56322; // @[Modules.scala 160:64:@1837.4]
  wire [13:0] _T_56323; // @[Modules.scala 160:64:@1838.4]
  wire [13:0] buffer_0_307; // @[Modules.scala 160:64:@1839.4]
  wire [13:0] buffer_0_12; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56325; // @[Modules.scala 160:64:@1841.4]
  wire [13:0] _T_56326; // @[Modules.scala 160:64:@1842.4]
  wire [13:0] buffer_0_308; // @[Modules.scala 160:64:@1843.4]
  wire [13:0] buffer_0_14; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_15; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56328; // @[Modules.scala 160:64:@1845.4]
  wire [13:0] _T_56329; // @[Modules.scala 160:64:@1846.4]
  wire [13:0] buffer_0_309; // @[Modules.scala 160:64:@1847.4]
  wire [13:0] buffer_0_16; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_17; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56331; // @[Modules.scala 160:64:@1849.4]
  wire [13:0] _T_56332; // @[Modules.scala 160:64:@1850.4]
  wire [13:0] buffer_0_310; // @[Modules.scala 160:64:@1851.4]
  wire [13:0] buffer_0_18; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_19; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56334; // @[Modules.scala 160:64:@1853.4]
  wire [13:0] _T_56335; // @[Modules.scala 160:64:@1854.4]
  wire [13:0] buffer_0_311; // @[Modules.scala 160:64:@1855.4]
  wire [13:0] buffer_0_20; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56337; // @[Modules.scala 160:64:@1857.4]
  wire [13:0] _T_56338; // @[Modules.scala 160:64:@1858.4]
  wire [13:0] buffer_0_312; // @[Modules.scala 160:64:@1859.4]
  wire [13:0] buffer_0_22; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_23; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56340; // @[Modules.scala 160:64:@1861.4]
  wire [13:0] _T_56341; // @[Modules.scala 160:64:@1862.4]
  wire [13:0] buffer_0_313; // @[Modules.scala 160:64:@1863.4]
  wire [13:0] buffer_0_24; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_25; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56343; // @[Modules.scala 160:64:@1865.4]
  wire [13:0] _T_56344; // @[Modules.scala 160:64:@1866.4]
  wire [13:0] buffer_0_314; // @[Modules.scala 160:64:@1867.4]
  wire [13:0] buffer_0_26; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56346; // @[Modules.scala 160:64:@1869.4]
  wire [13:0] _T_56347; // @[Modules.scala 160:64:@1870.4]
  wire [13:0] buffer_0_315; // @[Modules.scala 160:64:@1871.4]
  wire [13:0] buffer_0_28; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_29; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56349; // @[Modules.scala 160:64:@1873.4]
  wire [13:0] _T_56350; // @[Modules.scala 160:64:@1874.4]
  wire [13:0] buffer_0_316; // @[Modules.scala 160:64:@1875.4]
  wire [13:0] buffer_0_30; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_31; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56352; // @[Modules.scala 160:64:@1877.4]
  wire [13:0] _T_56353; // @[Modules.scala 160:64:@1878.4]
  wire [13:0] buffer_0_317; // @[Modules.scala 160:64:@1879.4]
  wire [13:0] buffer_0_32; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56355; // @[Modules.scala 160:64:@1881.4]
  wire [13:0] _T_56356; // @[Modules.scala 160:64:@1882.4]
  wire [13:0] buffer_0_318; // @[Modules.scala 160:64:@1883.4]
  wire [13:0] buffer_0_34; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56358; // @[Modules.scala 160:64:@1885.4]
  wire [13:0] _T_56359; // @[Modules.scala 160:64:@1886.4]
  wire [13:0] buffer_0_319; // @[Modules.scala 160:64:@1887.4]
  wire [13:0] buffer_0_36; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_37; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56361; // @[Modules.scala 160:64:@1889.4]
  wire [13:0] _T_56362; // @[Modules.scala 160:64:@1890.4]
  wire [13:0] buffer_0_320; // @[Modules.scala 160:64:@1891.4]
  wire [13:0] buffer_0_38; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_39; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56364; // @[Modules.scala 160:64:@1893.4]
  wire [13:0] _T_56365; // @[Modules.scala 160:64:@1894.4]
  wire [13:0] buffer_0_321; // @[Modules.scala 160:64:@1895.4]
  wire [13:0] buffer_0_40; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56367; // @[Modules.scala 160:64:@1897.4]
  wire [13:0] _T_56368; // @[Modules.scala 160:64:@1898.4]
  wire [13:0] buffer_0_322; // @[Modules.scala 160:64:@1899.4]
  wire [13:0] buffer_0_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56370; // @[Modules.scala 160:64:@1901.4]
  wire [13:0] _T_56371; // @[Modules.scala 160:64:@1902.4]
  wire [13:0] buffer_0_323; // @[Modules.scala 160:64:@1903.4]
  wire [13:0] buffer_0_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56373; // @[Modules.scala 160:64:@1905.4]
  wire [13:0] _T_56374; // @[Modules.scala 160:64:@1906.4]
  wire [13:0] buffer_0_324; // @[Modules.scala 160:64:@1907.4]
  wire [13:0] buffer_0_46; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_47; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56376; // @[Modules.scala 160:64:@1909.4]
  wire [13:0] _T_56377; // @[Modules.scala 160:64:@1910.4]
  wire [13:0] buffer_0_325; // @[Modules.scala 160:64:@1911.4]
  wire [13:0] buffer_0_48; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56379; // @[Modules.scala 160:64:@1913.4]
  wire [13:0] _T_56380; // @[Modules.scala 160:64:@1914.4]
  wire [13:0] buffer_0_326; // @[Modules.scala 160:64:@1915.4]
  wire [13:0] buffer_0_50; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56382; // @[Modules.scala 160:64:@1917.4]
  wire [13:0] _T_56383; // @[Modules.scala 160:64:@1918.4]
  wire [13:0] buffer_0_327; // @[Modules.scala 160:64:@1919.4]
  wire [13:0] buffer_0_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56385; // @[Modules.scala 160:64:@1921.4]
  wire [13:0] _T_56386; // @[Modules.scala 160:64:@1922.4]
  wire [13:0] buffer_0_328; // @[Modules.scala 160:64:@1923.4]
  wire [13:0] buffer_0_54; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56388; // @[Modules.scala 160:64:@1925.4]
  wire [13:0] _T_56389; // @[Modules.scala 160:64:@1926.4]
  wire [13:0] buffer_0_329; // @[Modules.scala 160:64:@1927.4]
  wire [13:0] buffer_0_56; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56391; // @[Modules.scala 160:64:@1929.4]
  wire [13:0] _T_56392; // @[Modules.scala 160:64:@1930.4]
  wire [13:0] buffer_0_330; // @[Modules.scala 160:64:@1931.4]
  wire [13:0] buffer_0_58; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56394; // @[Modules.scala 160:64:@1933.4]
  wire [13:0] _T_56395; // @[Modules.scala 160:64:@1934.4]
  wire [13:0] buffer_0_331; // @[Modules.scala 160:64:@1935.4]
  wire [13:0] buffer_0_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56397; // @[Modules.scala 160:64:@1937.4]
  wire [13:0] _T_56398; // @[Modules.scala 160:64:@1938.4]
  wire [13:0] buffer_0_332; // @[Modules.scala 160:64:@1939.4]
  wire [13:0] buffer_0_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56400; // @[Modules.scala 160:64:@1941.4]
  wire [13:0] _T_56401; // @[Modules.scala 160:64:@1942.4]
  wire [13:0] buffer_0_333; // @[Modules.scala 160:64:@1943.4]
  wire [13:0] buffer_0_64; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_65; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56403; // @[Modules.scala 160:64:@1945.4]
  wire [13:0] _T_56404; // @[Modules.scala 160:64:@1946.4]
  wire [13:0] buffer_0_334; // @[Modules.scala 160:64:@1947.4]
  wire [13:0] buffer_0_66; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56406; // @[Modules.scala 160:64:@1949.4]
  wire [13:0] _T_56407; // @[Modules.scala 160:64:@1950.4]
  wire [13:0] buffer_0_335; // @[Modules.scala 160:64:@1951.4]
  wire [13:0] buffer_0_68; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56409; // @[Modules.scala 160:64:@1953.4]
  wire [13:0] _T_56410; // @[Modules.scala 160:64:@1954.4]
  wire [13:0] buffer_0_336; // @[Modules.scala 160:64:@1955.4]
  wire [13:0] buffer_0_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56412; // @[Modules.scala 160:64:@1957.4]
  wire [13:0] _T_56413; // @[Modules.scala 160:64:@1958.4]
  wire [13:0] buffer_0_337; // @[Modules.scala 160:64:@1959.4]
  wire [13:0] buffer_0_72; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56415; // @[Modules.scala 160:64:@1961.4]
  wire [13:0] _T_56416; // @[Modules.scala 160:64:@1962.4]
  wire [13:0] buffer_0_338; // @[Modules.scala 160:64:@1963.4]
  wire [13:0] buffer_0_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56418; // @[Modules.scala 160:64:@1965.4]
  wire [13:0] _T_56419; // @[Modules.scala 160:64:@1966.4]
  wire [13:0] buffer_0_339; // @[Modules.scala 160:64:@1967.4]
  wire [13:0] buffer_0_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56421; // @[Modules.scala 160:64:@1969.4]
  wire [13:0] _T_56422; // @[Modules.scala 160:64:@1970.4]
  wire [13:0] buffer_0_340; // @[Modules.scala 160:64:@1971.4]
  wire [13:0] buffer_0_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56424; // @[Modules.scala 160:64:@1973.4]
  wire [13:0] _T_56425; // @[Modules.scala 160:64:@1974.4]
  wire [13:0] buffer_0_341; // @[Modules.scala 160:64:@1975.4]
  wire [13:0] buffer_0_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56427; // @[Modules.scala 160:64:@1977.4]
  wire [13:0] _T_56428; // @[Modules.scala 160:64:@1978.4]
  wire [13:0] buffer_0_342; // @[Modules.scala 160:64:@1979.4]
  wire [13:0] buffer_0_82; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_83; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56430; // @[Modules.scala 160:64:@1981.4]
  wire [13:0] _T_56431; // @[Modules.scala 160:64:@1982.4]
  wire [13:0] buffer_0_343; // @[Modules.scala 160:64:@1983.4]
  wire [13:0] buffer_0_84; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56433; // @[Modules.scala 160:64:@1985.4]
  wire [13:0] _T_56434; // @[Modules.scala 160:64:@1986.4]
  wire [13:0] buffer_0_344; // @[Modules.scala 160:64:@1987.4]
  wire [13:0] buffer_0_86; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_87; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56436; // @[Modules.scala 160:64:@1989.4]
  wire [13:0] _T_56437; // @[Modules.scala 160:64:@1990.4]
  wire [13:0] buffer_0_345; // @[Modules.scala 160:64:@1991.4]
  wire [13:0] buffer_0_88; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_89; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56439; // @[Modules.scala 160:64:@1993.4]
  wire [13:0] _T_56440; // @[Modules.scala 160:64:@1994.4]
  wire [13:0] buffer_0_346; // @[Modules.scala 160:64:@1995.4]
  wire [13:0] buffer_0_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56442; // @[Modules.scala 160:64:@1997.4]
  wire [13:0] _T_56443; // @[Modules.scala 160:64:@1998.4]
  wire [13:0] buffer_0_347; // @[Modules.scala 160:64:@1999.4]
  wire [13:0] buffer_0_92; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56445; // @[Modules.scala 160:64:@2001.4]
  wire [13:0] _T_56446; // @[Modules.scala 160:64:@2002.4]
  wire [13:0] buffer_0_348; // @[Modules.scala 160:64:@2003.4]
  wire [13:0] buffer_0_94; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56448; // @[Modules.scala 160:64:@2005.4]
  wire [13:0] _T_56449; // @[Modules.scala 160:64:@2006.4]
  wire [13:0] buffer_0_349; // @[Modules.scala 160:64:@2007.4]
  wire [13:0] buffer_0_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56451; // @[Modules.scala 160:64:@2009.4]
  wire [13:0] _T_56452; // @[Modules.scala 160:64:@2010.4]
  wire [13:0] buffer_0_350; // @[Modules.scala 160:64:@2011.4]
  wire [13:0] buffer_0_98; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_99; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56454; // @[Modules.scala 160:64:@2013.4]
  wire [13:0] _T_56455; // @[Modules.scala 160:64:@2014.4]
  wire [13:0] buffer_0_351; // @[Modules.scala 160:64:@2015.4]
  wire [13:0] buffer_0_100; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_101; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56457; // @[Modules.scala 160:64:@2017.4]
  wire [13:0] _T_56458; // @[Modules.scala 160:64:@2018.4]
  wire [13:0] buffer_0_352; // @[Modules.scala 160:64:@2019.4]
  wire [13:0] buffer_0_102; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_103; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56460; // @[Modules.scala 160:64:@2021.4]
  wire [13:0] _T_56461; // @[Modules.scala 160:64:@2022.4]
  wire [13:0] buffer_0_353; // @[Modules.scala 160:64:@2023.4]
  wire [13:0] buffer_0_104; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56463; // @[Modules.scala 160:64:@2025.4]
  wire [13:0] _T_56464; // @[Modules.scala 160:64:@2026.4]
  wire [13:0] buffer_0_354; // @[Modules.scala 160:64:@2027.4]
  wire [13:0] buffer_0_106; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56466; // @[Modules.scala 160:64:@2029.4]
  wire [13:0] _T_56467; // @[Modules.scala 160:64:@2030.4]
  wire [13:0] buffer_0_355; // @[Modules.scala 160:64:@2031.4]
  wire [13:0] buffer_0_108; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_109; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56469; // @[Modules.scala 160:64:@2033.4]
  wire [13:0] _T_56470; // @[Modules.scala 160:64:@2034.4]
  wire [13:0] buffer_0_356; // @[Modules.scala 160:64:@2035.4]
  wire [13:0] buffer_0_110; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56472; // @[Modules.scala 160:64:@2037.4]
  wire [13:0] _T_56473; // @[Modules.scala 160:64:@2038.4]
  wire [13:0] buffer_0_357; // @[Modules.scala 160:64:@2039.4]
  wire [13:0] buffer_0_112; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56475; // @[Modules.scala 160:64:@2041.4]
  wire [13:0] _T_56476; // @[Modules.scala 160:64:@2042.4]
  wire [13:0] buffer_0_358; // @[Modules.scala 160:64:@2043.4]
  wire [13:0] buffer_0_114; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56478; // @[Modules.scala 160:64:@2045.4]
  wire [13:0] _T_56479; // @[Modules.scala 160:64:@2046.4]
  wire [13:0] buffer_0_359; // @[Modules.scala 160:64:@2047.4]
  wire [13:0] buffer_0_116; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56481; // @[Modules.scala 160:64:@2049.4]
  wire [13:0] _T_56482; // @[Modules.scala 160:64:@2050.4]
  wire [13:0] buffer_0_360; // @[Modules.scala 160:64:@2051.4]
  wire [13:0] buffer_0_118; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_119; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56484; // @[Modules.scala 160:64:@2053.4]
  wire [13:0] _T_56485; // @[Modules.scala 160:64:@2054.4]
  wire [13:0] buffer_0_361; // @[Modules.scala 160:64:@2055.4]
  wire [13:0] buffer_0_120; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56487; // @[Modules.scala 160:64:@2057.4]
  wire [13:0] _T_56488; // @[Modules.scala 160:64:@2058.4]
  wire [13:0] buffer_0_362; // @[Modules.scala 160:64:@2059.4]
  wire [13:0] buffer_0_122; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56490; // @[Modules.scala 160:64:@2061.4]
  wire [13:0] _T_56491; // @[Modules.scala 160:64:@2062.4]
  wire [13:0] buffer_0_363; // @[Modules.scala 160:64:@2063.4]
  wire [13:0] buffer_0_124; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56493; // @[Modules.scala 160:64:@2065.4]
  wire [13:0] _T_56494; // @[Modules.scala 160:64:@2066.4]
  wire [13:0] buffer_0_364; // @[Modules.scala 160:64:@2067.4]
  wire [13:0] buffer_0_126; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_127; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56496; // @[Modules.scala 160:64:@2069.4]
  wire [13:0] _T_56497; // @[Modules.scala 160:64:@2070.4]
  wire [13:0] buffer_0_365; // @[Modules.scala 160:64:@2071.4]
  wire [13:0] buffer_0_128; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_129; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56499; // @[Modules.scala 160:64:@2073.4]
  wire [13:0] _T_56500; // @[Modules.scala 160:64:@2074.4]
  wire [13:0] buffer_0_366; // @[Modules.scala 160:64:@2075.4]
  wire [13:0] buffer_0_130; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56502; // @[Modules.scala 160:64:@2077.4]
  wire [13:0] _T_56503; // @[Modules.scala 160:64:@2078.4]
  wire [13:0] buffer_0_367; // @[Modules.scala 160:64:@2079.4]
  wire [13:0] buffer_0_132; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56505; // @[Modules.scala 160:64:@2081.4]
  wire [13:0] _T_56506; // @[Modules.scala 160:64:@2082.4]
  wire [13:0] buffer_0_368; // @[Modules.scala 160:64:@2083.4]
  wire [13:0] buffer_0_134; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56508; // @[Modules.scala 160:64:@2085.4]
  wire [13:0] _T_56509; // @[Modules.scala 160:64:@2086.4]
  wire [13:0] buffer_0_369; // @[Modules.scala 160:64:@2087.4]
  wire [13:0] buffer_0_136; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56511; // @[Modules.scala 160:64:@2089.4]
  wire [13:0] _T_56512; // @[Modules.scala 160:64:@2090.4]
  wire [13:0] buffer_0_370; // @[Modules.scala 160:64:@2091.4]
  wire [13:0] buffer_0_138; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_139; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56514; // @[Modules.scala 160:64:@2093.4]
  wire [13:0] _T_56515; // @[Modules.scala 160:64:@2094.4]
  wire [13:0] buffer_0_371; // @[Modules.scala 160:64:@2095.4]
  wire [13:0] buffer_0_140; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56517; // @[Modules.scala 160:64:@2097.4]
  wire [13:0] _T_56518; // @[Modules.scala 160:64:@2098.4]
  wire [13:0] buffer_0_372; // @[Modules.scala 160:64:@2099.4]
  wire [13:0] buffer_0_142; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_143; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56520; // @[Modules.scala 160:64:@2101.4]
  wire [13:0] _T_56521; // @[Modules.scala 160:64:@2102.4]
  wire [13:0] buffer_0_373; // @[Modules.scala 160:64:@2103.4]
  wire [13:0] buffer_0_144; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56523; // @[Modules.scala 160:64:@2105.4]
  wire [13:0] _T_56524; // @[Modules.scala 160:64:@2106.4]
  wire [13:0] buffer_0_374; // @[Modules.scala 160:64:@2107.4]
  wire [13:0] buffer_0_146; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56526; // @[Modules.scala 160:64:@2109.4]
  wire [13:0] _T_56527; // @[Modules.scala 160:64:@2110.4]
  wire [13:0] buffer_0_375; // @[Modules.scala 160:64:@2111.4]
  wire [13:0] buffer_0_148; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56529; // @[Modules.scala 160:64:@2113.4]
  wire [13:0] _T_56530; // @[Modules.scala 160:64:@2114.4]
  wire [13:0] buffer_0_376; // @[Modules.scala 160:64:@2115.4]
  wire [13:0] buffer_0_150; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56532; // @[Modules.scala 160:64:@2117.4]
  wire [13:0] _T_56533; // @[Modules.scala 160:64:@2118.4]
  wire [13:0] buffer_0_377; // @[Modules.scala 160:64:@2119.4]
  wire [13:0] buffer_0_152; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56535; // @[Modules.scala 160:64:@2121.4]
  wire [13:0] _T_56536; // @[Modules.scala 160:64:@2122.4]
  wire [13:0] buffer_0_378; // @[Modules.scala 160:64:@2123.4]
  wire [13:0] buffer_0_154; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56538; // @[Modules.scala 160:64:@2125.4]
  wire [13:0] _T_56539; // @[Modules.scala 160:64:@2126.4]
  wire [13:0] buffer_0_379; // @[Modules.scala 160:64:@2127.4]
  wire [13:0] buffer_0_156; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56541; // @[Modules.scala 160:64:@2129.4]
  wire [13:0] _T_56542; // @[Modules.scala 160:64:@2130.4]
  wire [13:0] buffer_0_380; // @[Modules.scala 160:64:@2131.4]
  wire [13:0] buffer_0_158; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56544; // @[Modules.scala 160:64:@2133.4]
  wire [13:0] _T_56545; // @[Modules.scala 160:64:@2134.4]
  wire [13:0] buffer_0_381; // @[Modules.scala 160:64:@2135.4]
  wire [13:0] buffer_0_160; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56547; // @[Modules.scala 160:64:@2137.4]
  wire [13:0] _T_56548; // @[Modules.scala 160:64:@2138.4]
  wire [13:0] buffer_0_382; // @[Modules.scala 160:64:@2139.4]
  wire [13:0] buffer_0_162; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_163; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56550; // @[Modules.scala 160:64:@2141.4]
  wire [13:0] _T_56551; // @[Modules.scala 160:64:@2142.4]
  wire [13:0] buffer_0_383; // @[Modules.scala 160:64:@2143.4]
  wire [13:0] buffer_0_164; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56553; // @[Modules.scala 160:64:@2145.4]
  wire [13:0] _T_56554; // @[Modules.scala 160:64:@2146.4]
  wire [13:0] buffer_0_384; // @[Modules.scala 160:64:@2147.4]
  wire [13:0] buffer_0_166; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56556; // @[Modules.scala 160:64:@2149.4]
  wire [13:0] _T_56557; // @[Modules.scala 160:64:@2150.4]
  wire [13:0] buffer_0_385; // @[Modules.scala 160:64:@2151.4]
  wire [13:0] buffer_0_168; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56559; // @[Modules.scala 160:64:@2153.4]
  wire [13:0] _T_56560; // @[Modules.scala 160:64:@2154.4]
  wire [13:0] buffer_0_386; // @[Modules.scala 160:64:@2155.4]
  wire [13:0] buffer_0_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56562; // @[Modules.scala 160:64:@2157.4]
  wire [13:0] _T_56563; // @[Modules.scala 160:64:@2158.4]
  wire [13:0] buffer_0_387; // @[Modules.scala 160:64:@2159.4]
  wire [13:0] buffer_0_172; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_173; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56565; // @[Modules.scala 160:64:@2161.4]
  wire [13:0] _T_56566; // @[Modules.scala 160:64:@2162.4]
  wire [13:0] buffer_0_388; // @[Modules.scala 160:64:@2163.4]
  wire [13:0] buffer_0_174; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56568; // @[Modules.scala 160:64:@2165.4]
  wire [13:0] _T_56569; // @[Modules.scala 160:64:@2166.4]
  wire [13:0] buffer_0_389; // @[Modules.scala 160:64:@2167.4]
  wire [13:0] buffer_0_176; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56571; // @[Modules.scala 160:64:@2169.4]
  wire [13:0] _T_56572; // @[Modules.scala 160:64:@2170.4]
  wire [13:0] buffer_0_390; // @[Modules.scala 160:64:@2171.4]
  wire [13:0] buffer_0_178; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_179; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56574; // @[Modules.scala 160:64:@2173.4]
  wire [13:0] _T_56575; // @[Modules.scala 160:64:@2174.4]
  wire [13:0] buffer_0_391; // @[Modules.scala 160:64:@2175.4]
  wire [13:0] buffer_0_180; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56577; // @[Modules.scala 160:64:@2177.4]
  wire [13:0] _T_56578; // @[Modules.scala 160:64:@2178.4]
  wire [13:0] buffer_0_392; // @[Modules.scala 160:64:@2179.4]
  wire [13:0] buffer_0_182; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56580; // @[Modules.scala 160:64:@2181.4]
  wire [13:0] _T_56581; // @[Modules.scala 160:64:@2182.4]
  wire [13:0] buffer_0_393; // @[Modules.scala 160:64:@2183.4]
  wire [13:0] buffer_0_184; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56583; // @[Modules.scala 160:64:@2185.4]
  wire [13:0] _T_56584; // @[Modules.scala 160:64:@2186.4]
  wire [13:0] buffer_0_394; // @[Modules.scala 160:64:@2187.4]
  wire [13:0] buffer_0_186; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_187; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56586; // @[Modules.scala 160:64:@2189.4]
  wire [13:0] _T_56587; // @[Modules.scala 160:64:@2190.4]
  wire [13:0] buffer_0_395; // @[Modules.scala 160:64:@2191.4]
  wire [13:0] buffer_0_188; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56589; // @[Modules.scala 160:64:@2193.4]
  wire [13:0] _T_56590; // @[Modules.scala 160:64:@2194.4]
  wire [13:0] buffer_0_396; // @[Modules.scala 160:64:@2195.4]
  wire [13:0] buffer_0_190; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56592; // @[Modules.scala 160:64:@2197.4]
  wire [13:0] _T_56593; // @[Modules.scala 160:64:@2198.4]
  wire [13:0] buffer_0_397; // @[Modules.scala 160:64:@2199.4]
  wire [13:0] buffer_0_192; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56595; // @[Modules.scala 160:64:@2201.4]
  wire [13:0] _T_56596; // @[Modules.scala 160:64:@2202.4]
  wire [13:0] buffer_0_398; // @[Modules.scala 160:64:@2203.4]
  wire [13:0] buffer_0_194; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56598; // @[Modules.scala 160:64:@2205.4]
  wire [13:0] _T_56599; // @[Modules.scala 160:64:@2206.4]
  wire [13:0] buffer_0_399; // @[Modules.scala 160:64:@2207.4]
  wire [13:0] buffer_0_196; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56601; // @[Modules.scala 160:64:@2209.4]
  wire [13:0] _T_56602; // @[Modules.scala 160:64:@2210.4]
  wire [13:0] buffer_0_400; // @[Modules.scala 160:64:@2211.4]
  wire [13:0] buffer_0_198; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56604; // @[Modules.scala 160:64:@2213.4]
  wire [13:0] _T_56605; // @[Modules.scala 160:64:@2214.4]
  wire [13:0] buffer_0_401; // @[Modules.scala 160:64:@2215.4]
  wire [13:0] buffer_0_200; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56607; // @[Modules.scala 160:64:@2217.4]
  wire [13:0] _T_56608; // @[Modules.scala 160:64:@2218.4]
  wire [13:0] buffer_0_402; // @[Modules.scala 160:64:@2219.4]
  wire [13:0] buffer_0_202; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56610; // @[Modules.scala 160:64:@2221.4]
  wire [13:0] _T_56611; // @[Modules.scala 160:64:@2222.4]
  wire [13:0] buffer_0_403; // @[Modules.scala 160:64:@2223.4]
  wire [13:0] buffer_0_204; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56613; // @[Modules.scala 160:64:@2225.4]
  wire [13:0] _T_56614; // @[Modules.scala 160:64:@2226.4]
  wire [13:0] buffer_0_404; // @[Modules.scala 160:64:@2227.4]
  wire [13:0] buffer_0_206; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56616; // @[Modules.scala 160:64:@2229.4]
  wire [13:0] _T_56617; // @[Modules.scala 160:64:@2230.4]
  wire [13:0] buffer_0_405; // @[Modules.scala 160:64:@2231.4]
  wire [13:0] buffer_0_208; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_209; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56619; // @[Modules.scala 160:64:@2233.4]
  wire [13:0] _T_56620; // @[Modules.scala 160:64:@2234.4]
  wire [13:0] buffer_0_406; // @[Modules.scala 160:64:@2235.4]
  wire [13:0] buffer_0_210; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56622; // @[Modules.scala 160:64:@2237.4]
  wire [13:0] _T_56623; // @[Modules.scala 160:64:@2238.4]
  wire [13:0] buffer_0_407; // @[Modules.scala 160:64:@2239.4]
  wire [13:0] buffer_0_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56625; // @[Modules.scala 160:64:@2241.4]
  wire [13:0] _T_56626; // @[Modules.scala 160:64:@2242.4]
  wire [13:0] buffer_0_408; // @[Modules.scala 160:64:@2243.4]
  wire [13:0] buffer_0_214; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56628; // @[Modules.scala 160:64:@2245.4]
  wire [13:0] _T_56629; // @[Modules.scala 160:64:@2246.4]
  wire [13:0] buffer_0_409; // @[Modules.scala 160:64:@2247.4]
  wire [13:0] buffer_0_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56631; // @[Modules.scala 160:64:@2249.4]
  wire [13:0] _T_56632; // @[Modules.scala 160:64:@2250.4]
  wire [13:0] buffer_0_410; // @[Modules.scala 160:64:@2251.4]
  wire [13:0] buffer_0_218; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56634; // @[Modules.scala 160:64:@2253.4]
  wire [13:0] _T_56635; // @[Modules.scala 160:64:@2254.4]
  wire [13:0] buffer_0_411; // @[Modules.scala 160:64:@2255.4]
  wire [13:0] buffer_0_220; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_221; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56637; // @[Modules.scala 160:64:@2257.4]
  wire [13:0] _T_56638; // @[Modules.scala 160:64:@2258.4]
  wire [13:0] buffer_0_412; // @[Modules.scala 160:64:@2259.4]
  wire [13:0] buffer_0_222; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56640; // @[Modules.scala 160:64:@2261.4]
  wire [13:0] _T_56641; // @[Modules.scala 160:64:@2262.4]
  wire [13:0] buffer_0_413; // @[Modules.scala 160:64:@2263.4]
  wire [13:0] buffer_0_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56643; // @[Modules.scala 160:64:@2265.4]
  wire [13:0] _T_56644; // @[Modules.scala 160:64:@2266.4]
  wire [13:0] buffer_0_414; // @[Modules.scala 160:64:@2267.4]
  wire [13:0] buffer_0_226; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56646; // @[Modules.scala 160:64:@2269.4]
  wire [13:0] _T_56647; // @[Modules.scala 160:64:@2270.4]
  wire [13:0] buffer_0_415; // @[Modules.scala 160:64:@2271.4]
  wire [13:0] buffer_0_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56649; // @[Modules.scala 160:64:@2273.4]
  wire [13:0] _T_56650; // @[Modules.scala 160:64:@2274.4]
  wire [13:0] buffer_0_416; // @[Modules.scala 160:64:@2275.4]
  wire [13:0] buffer_0_230; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56652; // @[Modules.scala 160:64:@2277.4]
  wire [13:0] _T_56653; // @[Modules.scala 160:64:@2278.4]
  wire [13:0] buffer_0_417; // @[Modules.scala 160:64:@2279.4]
  wire [13:0] buffer_0_232; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56655; // @[Modules.scala 160:64:@2281.4]
  wire [13:0] _T_56656; // @[Modules.scala 160:64:@2282.4]
  wire [13:0] buffer_0_418; // @[Modules.scala 160:64:@2283.4]
  wire [13:0] buffer_0_234; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56658; // @[Modules.scala 160:64:@2285.4]
  wire [13:0] _T_56659; // @[Modules.scala 160:64:@2286.4]
  wire [13:0] buffer_0_419; // @[Modules.scala 160:64:@2287.4]
  wire [13:0] buffer_0_236; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56661; // @[Modules.scala 160:64:@2289.4]
  wire [13:0] _T_56662; // @[Modules.scala 160:64:@2290.4]
  wire [13:0] buffer_0_420; // @[Modules.scala 160:64:@2291.4]
  wire [13:0] buffer_0_238; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56664; // @[Modules.scala 160:64:@2293.4]
  wire [13:0] _T_56665; // @[Modules.scala 160:64:@2294.4]
  wire [13:0] buffer_0_421; // @[Modules.scala 160:64:@2295.4]
  wire [13:0] buffer_0_240; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56667; // @[Modules.scala 160:64:@2297.4]
  wire [13:0] _T_56668; // @[Modules.scala 160:64:@2298.4]
  wire [13:0] buffer_0_422; // @[Modules.scala 160:64:@2299.4]
  wire [13:0] buffer_0_242; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56670; // @[Modules.scala 160:64:@2301.4]
  wire [13:0] _T_56671; // @[Modules.scala 160:64:@2302.4]
  wire [13:0] buffer_0_423; // @[Modules.scala 160:64:@2303.4]
  wire [13:0] buffer_0_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56673; // @[Modules.scala 160:64:@2305.4]
  wire [13:0] _T_56674; // @[Modules.scala 160:64:@2306.4]
  wire [13:0] buffer_0_424; // @[Modules.scala 160:64:@2307.4]
  wire [13:0] buffer_0_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56676; // @[Modules.scala 160:64:@2309.4]
  wire [13:0] _T_56677; // @[Modules.scala 160:64:@2310.4]
  wire [13:0] buffer_0_425; // @[Modules.scala 160:64:@2311.4]
  wire [13:0] buffer_0_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56679; // @[Modules.scala 160:64:@2313.4]
  wire [13:0] _T_56680; // @[Modules.scala 160:64:@2314.4]
  wire [13:0] buffer_0_426; // @[Modules.scala 160:64:@2315.4]
  wire [13:0] buffer_0_250; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56682; // @[Modules.scala 160:64:@2317.4]
  wire [13:0] _T_56683; // @[Modules.scala 160:64:@2318.4]
  wire [13:0] buffer_0_427; // @[Modules.scala 160:64:@2319.4]
  wire [13:0] buffer_0_252; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56685; // @[Modules.scala 160:64:@2321.4]
  wire [13:0] _T_56686; // @[Modules.scala 160:64:@2322.4]
  wire [13:0] buffer_0_428; // @[Modules.scala 160:64:@2323.4]
  wire [13:0] buffer_0_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56688; // @[Modules.scala 160:64:@2325.4]
  wire [13:0] _T_56689; // @[Modules.scala 160:64:@2326.4]
  wire [13:0] buffer_0_429; // @[Modules.scala 160:64:@2327.4]
  wire [13:0] buffer_0_256; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56691; // @[Modules.scala 160:64:@2329.4]
  wire [13:0] _T_56692; // @[Modules.scala 160:64:@2330.4]
  wire [13:0] buffer_0_430; // @[Modules.scala 160:64:@2331.4]
  wire [13:0] buffer_0_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56694; // @[Modules.scala 160:64:@2333.4]
  wire [13:0] _T_56695; // @[Modules.scala 160:64:@2334.4]
  wire [13:0] buffer_0_431; // @[Modules.scala 160:64:@2335.4]
  wire [13:0] buffer_0_260; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_261; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56697; // @[Modules.scala 160:64:@2337.4]
  wire [13:0] _T_56698; // @[Modules.scala 160:64:@2338.4]
  wire [13:0] buffer_0_432; // @[Modules.scala 160:64:@2339.4]
  wire [13:0] buffer_0_262; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56700; // @[Modules.scala 160:64:@2341.4]
  wire [13:0] _T_56701; // @[Modules.scala 160:64:@2342.4]
  wire [13:0] buffer_0_433; // @[Modules.scala 160:64:@2343.4]
  wire [13:0] buffer_0_264; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56703; // @[Modules.scala 160:64:@2345.4]
  wire [13:0] _T_56704; // @[Modules.scala 160:64:@2346.4]
  wire [13:0] buffer_0_434; // @[Modules.scala 160:64:@2347.4]
  wire [13:0] buffer_0_266; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_267; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56706; // @[Modules.scala 160:64:@2349.4]
  wire [13:0] _T_56707; // @[Modules.scala 160:64:@2350.4]
  wire [13:0] buffer_0_435; // @[Modules.scala 160:64:@2351.4]
  wire [13:0] buffer_0_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56709; // @[Modules.scala 160:64:@2353.4]
  wire [13:0] _T_56710; // @[Modules.scala 160:64:@2354.4]
  wire [13:0] buffer_0_436; // @[Modules.scala 160:64:@2355.4]
  wire [13:0] buffer_0_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56712; // @[Modules.scala 160:64:@2357.4]
  wire [13:0] _T_56713; // @[Modules.scala 160:64:@2358.4]
  wire [13:0] buffer_0_437; // @[Modules.scala 160:64:@2359.4]
  wire [13:0] buffer_0_272; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56715; // @[Modules.scala 160:64:@2361.4]
  wire [13:0] _T_56716; // @[Modules.scala 160:64:@2362.4]
  wire [13:0] buffer_0_438; // @[Modules.scala 160:64:@2363.4]
  wire [13:0] buffer_0_274; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_275; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56718; // @[Modules.scala 160:64:@2365.4]
  wire [13:0] _T_56719; // @[Modules.scala 160:64:@2366.4]
  wire [13:0] buffer_0_439; // @[Modules.scala 160:64:@2367.4]
  wire [13:0] buffer_0_276; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_277; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56721; // @[Modules.scala 160:64:@2369.4]
  wire [13:0] _T_56722; // @[Modules.scala 160:64:@2370.4]
  wire [13:0] buffer_0_440; // @[Modules.scala 160:64:@2371.4]
  wire [13:0] buffer_0_278; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56724; // @[Modules.scala 160:64:@2373.4]
  wire [13:0] _T_56725; // @[Modules.scala 160:64:@2374.4]
  wire [13:0] buffer_0_441; // @[Modules.scala 160:64:@2375.4]
  wire [13:0] buffer_0_280; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56727; // @[Modules.scala 160:64:@2377.4]
  wire [13:0] _T_56728; // @[Modules.scala 160:64:@2378.4]
  wire [13:0] buffer_0_442; // @[Modules.scala 160:64:@2379.4]
  wire [13:0] buffer_0_282; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56730; // @[Modules.scala 160:64:@2381.4]
  wire [13:0] _T_56731; // @[Modules.scala 160:64:@2382.4]
  wire [13:0] buffer_0_443; // @[Modules.scala 160:64:@2383.4]
  wire [13:0] buffer_0_284; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_285; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56733; // @[Modules.scala 160:64:@2385.4]
  wire [13:0] _T_56734; // @[Modules.scala 160:64:@2386.4]
  wire [13:0] buffer_0_444; // @[Modules.scala 160:64:@2387.4]
  wire [13:0] buffer_0_286; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_287; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56736; // @[Modules.scala 160:64:@2389.4]
  wire [13:0] _T_56737; // @[Modules.scala 160:64:@2390.4]
  wire [13:0] buffer_0_445; // @[Modules.scala 160:64:@2391.4]
  wire [13:0] buffer_0_288; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56739; // @[Modules.scala 160:64:@2393.4]
  wire [13:0] _T_56740; // @[Modules.scala 160:64:@2394.4]
  wire [13:0] buffer_0_446; // @[Modules.scala 160:64:@2395.4]
  wire [13:0] buffer_0_290; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56742; // @[Modules.scala 160:64:@2397.4]
  wire [13:0] _T_56743; // @[Modules.scala 160:64:@2398.4]
  wire [13:0] buffer_0_447; // @[Modules.scala 160:64:@2399.4]
  wire [13:0] buffer_0_292; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56745; // @[Modules.scala 160:64:@2401.4]
  wire [13:0] _T_56746; // @[Modules.scala 160:64:@2402.4]
  wire [13:0] buffer_0_448; // @[Modules.scala 160:64:@2403.4]
  wire [13:0] buffer_0_294; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56748; // @[Modules.scala 160:64:@2405.4]
  wire [13:0] _T_56749; // @[Modules.scala 160:64:@2406.4]
  wire [13:0] buffer_0_449; // @[Modules.scala 160:64:@2407.4]
  wire [13:0] buffer_0_296; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_297; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56751; // @[Modules.scala 160:64:@2409.4]
  wire [13:0] _T_56752; // @[Modules.scala 160:64:@2410.4]
  wire [13:0] buffer_0_450; // @[Modules.scala 160:64:@2411.4]
  wire [13:0] buffer_0_298; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56754; // @[Modules.scala 160:64:@2413.4]
  wire [13:0] _T_56755; // @[Modules.scala 160:64:@2414.4]
  wire [13:0] buffer_0_451; // @[Modules.scala 160:64:@2415.4]
  wire [13:0] buffer_0_300; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_0_301; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_56757; // @[Modules.scala 160:64:@2417.4]
  wire [13:0] _T_56758; // @[Modules.scala 160:64:@2418.4]
  wire [13:0] buffer_0_452; // @[Modules.scala 160:64:@2419.4]
  wire [14:0] _T_56760; // @[Modules.scala 166:64:@2421.4]
  wire [13:0] _T_56761; // @[Modules.scala 166:64:@2422.4]
  wire [13:0] buffer_0_453; // @[Modules.scala 166:64:@2423.4]
  wire [14:0] _T_56763; // @[Modules.scala 166:64:@2425.4]
  wire [13:0] _T_56764; // @[Modules.scala 166:64:@2426.4]
  wire [13:0] buffer_0_454; // @[Modules.scala 166:64:@2427.4]
  wire [14:0] _T_56766; // @[Modules.scala 166:64:@2429.4]
  wire [13:0] _T_56767; // @[Modules.scala 166:64:@2430.4]
  wire [13:0] buffer_0_455; // @[Modules.scala 166:64:@2431.4]
  wire [14:0] _T_56769; // @[Modules.scala 166:64:@2433.4]
  wire [13:0] _T_56770; // @[Modules.scala 166:64:@2434.4]
  wire [13:0] buffer_0_456; // @[Modules.scala 166:64:@2435.4]
  wire [14:0] _T_56772; // @[Modules.scala 166:64:@2437.4]
  wire [13:0] _T_56773; // @[Modules.scala 166:64:@2438.4]
  wire [13:0] buffer_0_457; // @[Modules.scala 166:64:@2439.4]
  wire [14:0] _T_56775; // @[Modules.scala 166:64:@2441.4]
  wire [13:0] _T_56776; // @[Modules.scala 166:64:@2442.4]
  wire [13:0] buffer_0_458; // @[Modules.scala 166:64:@2443.4]
  wire [14:0] _T_56778; // @[Modules.scala 166:64:@2445.4]
  wire [13:0] _T_56779; // @[Modules.scala 166:64:@2446.4]
  wire [13:0] buffer_0_459; // @[Modules.scala 166:64:@2447.4]
  wire [14:0] _T_56781; // @[Modules.scala 166:64:@2449.4]
  wire [13:0] _T_56782; // @[Modules.scala 166:64:@2450.4]
  wire [13:0] buffer_0_460; // @[Modules.scala 166:64:@2451.4]
  wire [14:0] _T_56784; // @[Modules.scala 166:64:@2453.4]
  wire [13:0] _T_56785; // @[Modules.scala 166:64:@2454.4]
  wire [13:0] buffer_0_461; // @[Modules.scala 166:64:@2455.4]
  wire [14:0] _T_56787; // @[Modules.scala 166:64:@2457.4]
  wire [13:0] _T_56788; // @[Modules.scala 166:64:@2458.4]
  wire [13:0] buffer_0_462; // @[Modules.scala 166:64:@2459.4]
  wire [14:0] _T_56790; // @[Modules.scala 166:64:@2461.4]
  wire [13:0] _T_56791; // @[Modules.scala 166:64:@2462.4]
  wire [13:0] buffer_0_463; // @[Modules.scala 166:64:@2463.4]
  wire [14:0] _T_56793; // @[Modules.scala 166:64:@2465.4]
  wire [13:0] _T_56794; // @[Modules.scala 166:64:@2466.4]
  wire [13:0] buffer_0_464; // @[Modules.scala 166:64:@2467.4]
  wire [14:0] _T_56796; // @[Modules.scala 166:64:@2469.4]
  wire [13:0] _T_56797; // @[Modules.scala 166:64:@2470.4]
  wire [13:0] buffer_0_465; // @[Modules.scala 166:64:@2471.4]
  wire [14:0] _T_56799; // @[Modules.scala 166:64:@2473.4]
  wire [13:0] _T_56800; // @[Modules.scala 166:64:@2474.4]
  wire [13:0] buffer_0_466; // @[Modules.scala 166:64:@2475.4]
  wire [14:0] _T_56802; // @[Modules.scala 166:64:@2477.4]
  wire [13:0] _T_56803; // @[Modules.scala 166:64:@2478.4]
  wire [13:0] buffer_0_467; // @[Modules.scala 166:64:@2479.4]
  wire [14:0] _T_56805; // @[Modules.scala 166:64:@2481.4]
  wire [13:0] _T_56806; // @[Modules.scala 166:64:@2482.4]
  wire [13:0] buffer_0_468; // @[Modules.scala 166:64:@2483.4]
  wire [14:0] _T_56808; // @[Modules.scala 166:64:@2485.4]
  wire [13:0] _T_56809; // @[Modules.scala 166:64:@2486.4]
  wire [13:0] buffer_0_469; // @[Modules.scala 166:64:@2487.4]
  wire [14:0] _T_56811; // @[Modules.scala 166:64:@2489.4]
  wire [13:0] _T_56812; // @[Modules.scala 166:64:@2490.4]
  wire [13:0] buffer_0_470; // @[Modules.scala 166:64:@2491.4]
  wire [14:0] _T_56814; // @[Modules.scala 166:64:@2493.4]
  wire [13:0] _T_56815; // @[Modules.scala 166:64:@2494.4]
  wire [13:0] buffer_0_471; // @[Modules.scala 166:64:@2495.4]
  wire [14:0] _T_56817; // @[Modules.scala 166:64:@2497.4]
  wire [13:0] _T_56818; // @[Modules.scala 166:64:@2498.4]
  wire [13:0] buffer_0_472; // @[Modules.scala 166:64:@2499.4]
  wire [14:0] _T_56820; // @[Modules.scala 166:64:@2501.4]
  wire [13:0] _T_56821; // @[Modules.scala 166:64:@2502.4]
  wire [13:0] buffer_0_473; // @[Modules.scala 166:64:@2503.4]
  wire [14:0] _T_56823; // @[Modules.scala 166:64:@2505.4]
  wire [13:0] _T_56824; // @[Modules.scala 166:64:@2506.4]
  wire [13:0] buffer_0_474; // @[Modules.scala 166:64:@2507.4]
  wire [14:0] _T_56826; // @[Modules.scala 166:64:@2509.4]
  wire [13:0] _T_56827; // @[Modules.scala 166:64:@2510.4]
  wire [13:0] buffer_0_475; // @[Modules.scala 166:64:@2511.4]
  wire [14:0] _T_56829; // @[Modules.scala 166:64:@2513.4]
  wire [13:0] _T_56830; // @[Modules.scala 166:64:@2514.4]
  wire [13:0] buffer_0_476; // @[Modules.scala 166:64:@2515.4]
  wire [14:0] _T_56832; // @[Modules.scala 166:64:@2517.4]
  wire [13:0] _T_56833; // @[Modules.scala 166:64:@2518.4]
  wire [13:0] buffer_0_477; // @[Modules.scala 166:64:@2519.4]
  wire [14:0] _T_56835; // @[Modules.scala 166:64:@2521.4]
  wire [13:0] _T_56836; // @[Modules.scala 166:64:@2522.4]
  wire [13:0] buffer_0_478; // @[Modules.scala 166:64:@2523.4]
  wire [14:0] _T_56838; // @[Modules.scala 166:64:@2525.4]
  wire [13:0] _T_56839; // @[Modules.scala 166:64:@2526.4]
  wire [13:0] buffer_0_479; // @[Modules.scala 166:64:@2527.4]
  wire [14:0] _T_56841; // @[Modules.scala 166:64:@2529.4]
  wire [13:0] _T_56842; // @[Modules.scala 166:64:@2530.4]
  wire [13:0] buffer_0_480; // @[Modules.scala 166:64:@2531.4]
  wire [14:0] _T_56844; // @[Modules.scala 166:64:@2533.4]
  wire [13:0] _T_56845; // @[Modules.scala 166:64:@2534.4]
  wire [13:0] buffer_0_481; // @[Modules.scala 166:64:@2535.4]
  wire [14:0] _T_56847; // @[Modules.scala 166:64:@2537.4]
  wire [13:0] _T_56848; // @[Modules.scala 166:64:@2538.4]
  wire [13:0] buffer_0_482; // @[Modules.scala 166:64:@2539.4]
  wire [14:0] _T_56850; // @[Modules.scala 166:64:@2541.4]
  wire [13:0] _T_56851; // @[Modules.scala 166:64:@2542.4]
  wire [13:0] buffer_0_483; // @[Modules.scala 166:64:@2543.4]
  wire [14:0] _T_56853; // @[Modules.scala 166:64:@2545.4]
  wire [13:0] _T_56854; // @[Modules.scala 166:64:@2546.4]
  wire [13:0] buffer_0_484; // @[Modules.scala 166:64:@2547.4]
  wire [14:0] _T_56856; // @[Modules.scala 166:64:@2549.4]
  wire [13:0] _T_56857; // @[Modules.scala 166:64:@2550.4]
  wire [13:0] buffer_0_485; // @[Modules.scala 166:64:@2551.4]
  wire [14:0] _T_56859; // @[Modules.scala 166:64:@2553.4]
  wire [13:0] _T_56860; // @[Modules.scala 166:64:@2554.4]
  wire [13:0] buffer_0_486; // @[Modules.scala 166:64:@2555.4]
  wire [14:0] _T_56862; // @[Modules.scala 166:64:@2557.4]
  wire [13:0] _T_56863; // @[Modules.scala 166:64:@2558.4]
  wire [13:0] buffer_0_487; // @[Modules.scala 166:64:@2559.4]
  wire [14:0] _T_56865; // @[Modules.scala 166:64:@2561.4]
  wire [13:0] _T_56866; // @[Modules.scala 166:64:@2562.4]
  wire [13:0] buffer_0_488; // @[Modules.scala 166:64:@2563.4]
  wire [14:0] _T_56868; // @[Modules.scala 166:64:@2565.4]
  wire [13:0] _T_56869; // @[Modules.scala 166:64:@2566.4]
  wire [13:0] buffer_0_489; // @[Modules.scala 166:64:@2567.4]
  wire [14:0] _T_56871; // @[Modules.scala 166:64:@2569.4]
  wire [13:0] _T_56872; // @[Modules.scala 166:64:@2570.4]
  wire [13:0] buffer_0_490; // @[Modules.scala 166:64:@2571.4]
  wire [14:0] _T_56874; // @[Modules.scala 166:64:@2573.4]
  wire [13:0] _T_56875; // @[Modules.scala 166:64:@2574.4]
  wire [13:0] buffer_0_491; // @[Modules.scala 166:64:@2575.4]
  wire [14:0] _T_56877; // @[Modules.scala 166:64:@2577.4]
  wire [13:0] _T_56878; // @[Modules.scala 166:64:@2578.4]
  wire [13:0] buffer_0_492; // @[Modules.scala 166:64:@2579.4]
  wire [14:0] _T_56880; // @[Modules.scala 166:64:@2581.4]
  wire [13:0] _T_56881; // @[Modules.scala 166:64:@2582.4]
  wire [13:0] buffer_0_493; // @[Modules.scala 166:64:@2583.4]
  wire [14:0] _T_56883; // @[Modules.scala 166:64:@2585.4]
  wire [13:0] _T_56884; // @[Modules.scala 166:64:@2586.4]
  wire [13:0] buffer_0_494; // @[Modules.scala 166:64:@2587.4]
  wire [14:0] _T_56886; // @[Modules.scala 166:64:@2589.4]
  wire [13:0] _T_56887; // @[Modules.scala 166:64:@2590.4]
  wire [13:0] buffer_0_495; // @[Modules.scala 166:64:@2591.4]
  wire [14:0] _T_56889; // @[Modules.scala 166:64:@2593.4]
  wire [13:0] _T_56890; // @[Modules.scala 166:64:@2594.4]
  wire [13:0] buffer_0_496; // @[Modules.scala 166:64:@2595.4]
  wire [14:0] _T_56892; // @[Modules.scala 166:64:@2597.4]
  wire [13:0] _T_56893; // @[Modules.scala 166:64:@2598.4]
  wire [13:0] buffer_0_497; // @[Modules.scala 166:64:@2599.4]
  wire [14:0] _T_56895; // @[Modules.scala 166:64:@2601.4]
  wire [13:0] _T_56896; // @[Modules.scala 166:64:@2602.4]
  wire [13:0] buffer_0_498; // @[Modules.scala 166:64:@2603.4]
  wire [14:0] _T_56898; // @[Modules.scala 166:64:@2605.4]
  wire [13:0] _T_56899; // @[Modules.scala 166:64:@2606.4]
  wire [13:0] buffer_0_499; // @[Modules.scala 166:64:@2607.4]
  wire [14:0] _T_56901; // @[Modules.scala 166:64:@2609.4]
  wire [13:0] _T_56902; // @[Modules.scala 166:64:@2610.4]
  wire [13:0] buffer_0_500; // @[Modules.scala 166:64:@2611.4]
  wire [14:0] _T_56904; // @[Modules.scala 166:64:@2613.4]
  wire [13:0] _T_56905; // @[Modules.scala 166:64:@2614.4]
  wire [13:0] buffer_0_501; // @[Modules.scala 166:64:@2615.4]
  wire [14:0] _T_56907; // @[Modules.scala 166:64:@2617.4]
  wire [13:0] _T_56908; // @[Modules.scala 166:64:@2618.4]
  wire [13:0] buffer_0_502; // @[Modules.scala 166:64:@2619.4]
  wire [14:0] _T_56910; // @[Modules.scala 166:64:@2621.4]
  wire [13:0] _T_56911; // @[Modules.scala 166:64:@2622.4]
  wire [13:0] buffer_0_503; // @[Modules.scala 166:64:@2623.4]
  wire [14:0] _T_56913; // @[Modules.scala 166:64:@2625.4]
  wire [13:0] _T_56914; // @[Modules.scala 166:64:@2626.4]
  wire [13:0] buffer_0_504; // @[Modules.scala 166:64:@2627.4]
  wire [14:0] _T_56916; // @[Modules.scala 166:64:@2629.4]
  wire [13:0] _T_56917; // @[Modules.scala 166:64:@2630.4]
  wire [13:0] buffer_0_505; // @[Modules.scala 166:64:@2631.4]
  wire [14:0] _T_56919; // @[Modules.scala 166:64:@2633.4]
  wire [13:0] _T_56920; // @[Modules.scala 166:64:@2634.4]
  wire [13:0] buffer_0_506; // @[Modules.scala 166:64:@2635.4]
  wire [14:0] _T_56922; // @[Modules.scala 166:64:@2637.4]
  wire [13:0] _T_56923; // @[Modules.scala 166:64:@2638.4]
  wire [13:0] buffer_0_507; // @[Modules.scala 166:64:@2639.4]
  wire [14:0] _T_56925; // @[Modules.scala 166:64:@2641.4]
  wire [13:0] _T_56926; // @[Modules.scala 166:64:@2642.4]
  wire [13:0] buffer_0_508; // @[Modules.scala 166:64:@2643.4]
  wire [14:0] _T_56928; // @[Modules.scala 166:64:@2645.4]
  wire [13:0] _T_56929; // @[Modules.scala 166:64:@2646.4]
  wire [13:0] buffer_0_509; // @[Modules.scala 166:64:@2647.4]
  wire [14:0] _T_56931; // @[Modules.scala 166:64:@2649.4]
  wire [13:0] _T_56932; // @[Modules.scala 166:64:@2650.4]
  wire [13:0] buffer_0_510; // @[Modules.scala 166:64:@2651.4]
  wire [14:0] _T_56934; // @[Modules.scala 166:64:@2653.4]
  wire [13:0] _T_56935; // @[Modules.scala 166:64:@2654.4]
  wire [13:0] buffer_0_511; // @[Modules.scala 166:64:@2655.4]
  wire [14:0] _T_56937; // @[Modules.scala 166:64:@2657.4]
  wire [13:0] _T_56938; // @[Modules.scala 166:64:@2658.4]
  wire [13:0] buffer_0_512; // @[Modules.scala 166:64:@2659.4]
  wire [14:0] _T_56940; // @[Modules.scala 166:64:@2661.4]
  wire [13:0] _T_56941; // @[Modules.scala 166:64:@2662.4]
  wire [13:0] buffer_0_513; // @[Modules.scala 166:64:@2663.4]
  wire [14:0] _T_56943; // @[Modules.scala 166:64:@2665.4]
  wire [13:0] _T_56944; // @[Modules.scala 166:64:@2666.4]
  wire [13:0] buffer_0_514; // @[Modules.scala 166:64:@2667.4]
  wire [14:0] _T_56946; // @[Modules.scala 166:64:@2669.4]
  wire [13:0] _T_56947; // @[Modules.scala 166:64:@2670.4]
  wire [13:0] buffer_0_515; // @[Modules.scala 166:64:@2671.4]
  wire [14:0] _T_56949; // @[Modules.scala 166:64:@2673.4]
  wire [13:0] _T_56950; // @[Modules.scala 166:64:@2674.4]
  wire [13:0] buffer_0_516; // @[Modules.scala 166:64:@2675.4]
  wire [14:0] _T_56952; // @[Modules.scala 166:64:@2677.4]
  wire [13:0] _T_56953; // @[Modules.scala 166:64:@2678.4]
  wire [13:0] buffer_0_517; // @[Modules.scala 166:64:@2679.4]
  wire [14:0] _T_56955; // @[Modules.scala 166:64:@2681.4]
  wire [13:0] _T_56956; // @[Modules.scala 166:64:@2682.4]
  wire [13:0] buffer_0_518; // @[Modules.scala 166:64:@2683.4]
  wire [14:0] _T_56958; // @[Modules.scala 166:64:@2685.4]
  wire [13:0] _T_56959; // @[Modules.scala 166:64:@2686.4]
  wire [13:0] buffer_0_519; // @[Modules.scala 166:64:@2687.4]
  wire [14:0] _T_56961; // @[Modules.scala 166:64:@2689.4]
  wire [13:0] _T_56962; // @[Modules.scala 166:64:@2690.4]
  wire [13:0] buffer_0_520; // @[Modules.scala 166:64:@2691.4]
  wire [14:0] _T_56964; // @[Modules.scala 166:64:@2693.4]
  wire [13:0] _T_56965; // @[Modules.scala 166:64:@2694.4]
  wire [13:0] buffer_0_521; // @[Modules.scala 166:64:@2695.4]
  wire [14:0] _T_56967; // @[Modules.scala 166:64:@2697.4]
  wire [13:0] _T_56968; // @[Modules.scala 166:64:@2698.4]
  wire [13:0] buffer_0_522; // @[Modules.scala 166:64:@2699.4]
  wire [14:0] _T_56970; // @[Modules.scala 166:64:@2701.4]
  wire [13:0] _T_56971; // @[Modules.scala 166:64:@2702.4]
  wire [13:0] buffer_0_523; // @[Modules.scala 166:64:@2703.4]
  wire [14:0] _T_56973; // @[Modules.scala 166:64:@2705.4]
  wire [13:0] _T_56974; // @[Modules.scala 166:64:@2706.4]
  wire [13:0] buffer_0_524; // @[Modules.scala 166:64:@2707.4]
  wire [14:0] _T_56976; // @[Modules.scala 166:64:@2709.4]
  wire [13:0] _T_56977; // @[Modules.scala 166:64:@2710.4]
  wire [13:0] buffer_0_525; // @[Modules.scala 166:64:@2711.4]
  wire [14:0] _T_56979; // @[Modules.scala 166:64:@2713.4]
  wire [13:0] _T_56980; // @[Modules.scala 166:64:@2714.4]
  wire [13:0] buffer_0_526; // @[Modules.scala 166:64:@2715.4]
  wire [14:0] _T_56982; // @[Modules.scala 166:64:@2717.4]
  wire [13:0] _T_56983; // @[Modules.scala 166:64:@2718.4]
  wire [13:0] buffer_0_527; // @[Modules.scala 166:64:@2719.4]
  wire [14:0] _T_56985; // @[Modules.scala 166:64:@2721.4]
  wire [13:0] _T_56986; // @[Modules.scala 166:64:@2722.4]
  wire [13:0] buffer_0_528; // @[Modules.scala 166:64:@2723.4]
  wire [14:0] _T_56988; // @[Modules.scala 166:64:@2725.4]
  wire [13:0] _T_56989; // @[Modules.scala 166:64:@2726.4]
  wire [13:0] buffer_0_529; // @[Modules.scala 166:64:@2727.4]
  wire [14:0] _T_56991; // @[Modules.scala 166:64:@2729.4]
  wire [13:0] _T_56992; // @[Modules.scala 166:64:@2730.4]
  wire [13:0] buffer_0_530; // @[Modules.scala 166:64:@2731.4]
  wire [14:0] _T_56994; // @[Modules.scala 166:64:@2733.4]
  wire [13:0] _T_56995; // @[Modules.scala 166:64:@2734.4]
  wire [13:0] buffer_0_531; // @[Modules.scala 166:64:@2735.4]
  wire [14:0] _T_56997; // @[Modules.scala 166:64:@2737.4]
  wire [13:0] _T_56998; // @[Modules.scala 166:64:@2738.4]
  wire [13:0] buffer_0_532; // @[Modules.scala 166:64:@2739.4]
  wire [14:0] _T_57000; // @[Modules.scala 166:64:@2741.4]
  wire [13:0] _T_57001; // @[Modules.scala 166:64:@2742.4]
  wire [13:0] buffer_0_533; // @[Modules.scala 166:64:@2743.4]
  wire [14:0] _T_57003; // @[Modules.scala 166:64:@2745.4]
  wire [13:0] _T_57004; // @[Modules.scala 166:64:@2746.4]
  wire [13:0] buffer_0_534; // @[Modules.scala 166:64:@2747.4]
  wire [14:0] _T_57006; // @[Modules.scala 166:64:@2749.4]
  wire [13:0] _T_57007; // @[Modules.scala 166:64:@2750.4]
  wire [13:0] buffer_0_535; // @[Modules.scala 166:64:@2751.4]
  wire [14:0] _T_57009; // @[Modules.scala 166:64:@2753.4]
  wire [13:0] _T_57010; // @[Modules.scala 166:64:@2754.4]
  wire [13:0] buffer_0_536; // @[Modules.scala 166:64:@2755.4]
  wire [14:0] _T_57012; // @[Modules.scala 166:64:@2757.4]
  wire [13:0] _T_57013; // @[Modules.scala 166:64:@2758.4]
  wire [13:0] buffer_0_537; // @[Modules.scala 166:64:@2759.4]
  wire [14:0] _T_57015; // @[Modules.scala 166:64:@2761.4]
  wire [13:0] _T_57016; // @[Modules.scala 166:64:@2762.4]
  wire [13:0] buffer_0_538; // @[Modules.scala 166:64:@2763.4]
  wire [14:0] _T_57018; // @[Modules.scala 166:64:@2765.4]
  wire [13:0] _T_57019; // @[Modules.scala 166:64:@2766.4]
  wire [13:0] buffer_0_539; // @[Modules.scala 166:64:@2767.4]
  wire [14:0] _T_57021; // @[Modules.scala 166:64:@2769.4]
  wire [13:0] _T_57022; // @[Modules.scala 166:64:@2770.4]
  wire [13:0] buffer_0_540; // @[Modules.scala 166:64:@2771.4]
  wire [14:0] _T_57024; // @[Modules.scala 166:64:@2773.4]
  wire [13:0] _T_57025; // @[Modules.scala 166:64:@2774.4]
  wire [13:0] buffer_0_541; // @[Modules.scala 166:64:@2775.4]
  wire [14:0] _T_57027; // @[Modules.scala 166:64:@2777.4]
  wire [13:0] _T_57028; // @[Modules.scala 166:64:@2778.4]
  wire [13:0] buffer_0_542; // @[Modules.scala 166:64:@2779.4]
  wire [14:0] _T_57030; // @[Modules.scala 166:64:@2781.4]
  wire [13:0] _T_57031; // @[Modules.scala 166:64:@2782.4]
  wire [13:0] buffer_0_543; // @[Modules.scala 166:64:@2783.4]
  wire [14:0] _T_57033; // @[Modules.scala 166:64:@2785.4]
  wire [13:0] _T_57034; // @[Modules.scala 166:64:@2786.4]
  wire [13:0] buffer_0_544; // @[Modules.scala 166:64:@2787.4]
  wire [14:0] _T_57036; // @[Modules.scala 166:64:@2789.4]
  wire [13:0] _T_57037; // @[Modules.scala 166:64:@2790.4]
  wire [13:0] buffer_0_545; // @[Modules.scala 166:64:@2791.4]
  wire [14:0] _T_57039; // @[Modules.scala 166:64:@2793.4]
  wire [13:0] _T_57040; // @[Modules.scala 166:64:@2794.4]
  wire [13:0] buffer_0_546; // @[Modules.scala 166:64:@2795.4]
  wire [14:0] _T_57042; // @[Modules.scala 166:64:@2797.4]
  wire [13:0] _T_57043; // @[Modules.scala 166:64:@2798.4]
  wire [13:0] buffer_0_547; // @[Modules.scala 166:64:@2799.4]
  wire [14:0] _T_57045; // @[Modules.scala 166:64:@2801.4]
  wire [13:0] _T_57046; // @[Modules.scala 166:64:@2802.4]
  wire [13:0] buffer_0_548; // @[Modules.scala 166:64:@2803.4]
  wire [14:0] _T_57048; // @[Modules.scala 166:64:@2805.4]
  wire [13:0] _T_57049; // @[Modules.scala 166:64:@2806.4]
  wire [13:0] buffer_0_549; // @[Modules.scala 166:64:@2807.4]
  wire [14:0] _T_57051; // @[Modules.scala 166:64:@2809.4]
  wire [13:0] _T_57052; // @[Modules.scala 166:64:@2810.4]
  wire [13:0] buffer_0_550; // @[Modules.scala 166:64:@2811.4]
  wire [14:0] _T_57054; // @[Modules.scala 166:64:@2813.4]
  wire [13:0] _T_57055; // @[Modules.scala 166:64:@2814.4]
  wire [13:0] buffer_0_551; // @[Modules.scala 166:64:@2815.4]
  wire [14:0] _T_57057; // @[Modules.scala 166:64:@2817.4]
  wire [13:0] _T_57058; // @[Modules.scala 166:64:@2818.4]
  wire [13:0] buffer_0_552; // @[Modules.scala 166:64:@2819.4]
  wire [14:0] _T_57060; // @[Modules.scala 166:64:@2821.4]
  wire [13:0] _T_57061; // @[Modules.scala 166:64:@2822.4]
  wire [13:0] buffer_0_553; // @[Modules.scala 166:64:@2823.4]
  wire [14:0] _T_57063; // @[Modules.scala 166:64:@2825.4]
  wire [13:0] _T_57064; // @[Modules.scala 166:64:@2826.4]
  wire [13:0] buffer_0_554; // @[Modules.scala 166:64:@2827.4]
  wire [14:0] _T_57066; // @[Modules.scala 166:64:@2829.4]
  wire [13:0] _T_57067; // @[Modules.scala 166:64:@2830.4]
  wire [13:0] buffer_0_555; // @[Modules.scala 166:64:@2831.4]
  wire [14:0] _T_57069; // @[Modules.scala 166:64:@2833.4]
  wire [13:0] _T_57070; // @[Modules.scala 166:64:@2834.4]
  wire [13:0] buffer_0_556; // @[Modules.scala 166:64:@2835.4]
  wire [14:0] _T_57072; // @[Modules.scala 166:64:@2837.4]
  wire [13:0] _T_57073; // @[Modules.scala 166:64:@2838.4]
  wire [13:0] buffer_0_557; // @[Modules.scala 166:64:@2839.4]
  wire [14:0] _T_57075; // @[Modules.scala 166:64:@2841.4]
  wire [13:0] _T_57076; // @[Modules.scala 166:64:@2842.4]
  wire [13:0] buffer_0_558; // @[Modules.scala 166:64:@2843.4]
  wire [14:0] _T_57078; // @[Modules.scala 166:64:@2845.4]
  wire [13:0] _T_57079; // @[Modules.scala 166:64:@2846.4]
  wire [13:0] buffer_0_559; // @[Modules.scala 166:64:@2847.4]
  wire [14:0] _T_57081; // @[Modules.scala 166:64:@2849.4]
  wire [13:0] _T_57082; // @[Modules.scala 166:64:@2850.4]
  wire [13:0] buffer_0_560; // @[Modules.scala 166:64:@2851.4]
  wire [14:0] _T_57084; // @[Modules.scala 166:64:@2853.4]
  wire [13:0] _T_57085; // @[Modules.scala 166:64:@2854.4]
  wire [13:0] buffer_0_561; // @[Modules.scala 166:64:@2855.4]
  wire [14:0] _T_57087; // @[Modules.scala 166:64:@2857.4]
  wire [13:0] _T_57088; // @[Modules.scala 166:64:@2858.4]
  wire [13:0] buffer_0_562; // @[Modules.scala 166:64:@2859.4]
  wire [14:0] _T_57090; // @[Modules.scala 166:64:@2861.4]
  wire [13:0] _T_57091; // @[Modules.scala 166:64:@2862.4]
  wire [13:0] buffer_0_563; // @[Modules.scala 166:64:@2863.4]
  wire [14:0] _T_57093; // @[Modules.scala 166:64:@2865.4]
  wire [13:0] _T_57094; // @[Modules.scala 166:64:@2866.4]
  wire [13:0] buffer_0_564; // @[Modules.scala 166:64:@2867.4]
  wire [14:0] _T_57096; // @[Modules.scala 172:66:@2869.4]
  wire [13:0] _T_57097; // @[Modules.scala 172:66:@2870.4]
  wire [13:0] buffer_0_565; // @[Modules.scala 172:66:@2871.4]
  wire [14:0] _T_57099; // @[Modules.scala 160:64:@2873.4]
  wire [13:0] _T_57100; // @[Modules.scala 160:64:@2874.4]
  wire [13:0] buffer_0_566; // @[Modules.scala 160:64:@2875.4]
  wire [14:0] _T_57102; // @[Modules.scala 160:64:@2877.4]
  wire [13:0] _T_57103; // @[Modules.scala 160:64:@2878.4]
  wire [13:0] buffer_0_567; // @[Modules.scala 160:64:@2879.4]
  wire [14:0] _T_57105; // @[Modules.scala 160:64:@2881.4]
  wire [13:0] _T_57106; // @[Modules.scala 160:64:@2882.4]
  wire [13:0] buffer_0_568; // @[Modules.scala 160:64:@2883.4]
  wire [14:0] _T_57108; // @[Modules.scala 160:64:@2885.4]
  wire [13:0] _T_57109; // @[Modules.scala 160:64:@2886.4]
  wire [13:0] buffer_0_569; // @[Modules.scala 160:64:@2887.4]
  wire [14:0] _T_57111; // @[Modules.scala 160:64:@2889.4]
  wire [13:0] _T_57112; // @[Modules.scala 160:64:@2890.4]
  wire [13:0] buffer_0_570; // @[Modules.scala 160:64:@2891.4]
  wire [14:0] _T_57114; // @[Modules.scala 160:64:@2893.4]
  wire [13:0] _T_57115; // @[Modules.scala 160:64:@2894.4]
  wire [13:0] buffer_0_571; // @[Modules.scala 160:64:@2895.4]
  wire [14:0] _T_57117; // @[Modules.scala 160:64:@2897.4]
  wire [13:0] _T_57118; // @[Modules.scala 160:64:@2898.4]
  wire [13:0] buffer_0_572; // @[Modules.scala 160:64:@2899.4]
  wire [14:0] _T_57120; // @[Modules.scala 160:64:@2901.4]
  wire [13:0] _T_57121; // @[Modules.scala 160:64:@2902.4]
  wire [13:0] buffer_0_573; // @[Modules.scala 160:64:@2903.4]
  wire [14:0] _T_57123; // @[Modules.scala 160:64:@2905.4]
  wire [13:0] _T_57124; // @[Modules.scala 160:64:@2906.4]
  wire [13:0] buffer_0_574; // @[Modules.scala 160:64:@2907.4]
  wire [14:0] _T_57126; // @[Modules.scala 160:64:@2909.4]
  wire [13:0] _T_57127; // @[Modules.scala 160:64:@2910.4]
  wire [13:0] buffer_0_575; // @[Modules.scala 160:64:@2911.4]
  wire [14:0] _T_57129; // @[Modules.scala 160:64:@2913.4]
  wire [13:0] _T_57130; // @[Modules.scala 160:64:@2914.4]
  wire [13:0] buffer_0_576; // @[Modules.scala 160:64:@2915.4]
  wire [14:0] _T_57132; // @[Modules.scala 160:64:@2917.4]
  wire [13:0] _T_57133; // @[Modules.scala 160:64:@2918.4]
  wire [13:0] buffer_0_577; // @[Modules.scala 160:64:@2919.4]
  wire [14:0] _T_57135; // @[Modules.scala 160:64:@2921.4]
  wire [13:0] _T_57136; // @[Modules.scala 160:64:@2922.4]
  wire [13:0] buffer_0_578; // @[Modules.scala 160:64:@2923.4]
  wire [14:0] _T_57138; // @[Modules.scala 160:64:@2925.4]
  wire [13:0] _T_57139; // @[Modules.scala 160:64:@2926.4]
  wire [13:0] buffer_0_579; // @[Modules.scala 160:64:@2927.4]
  wire [14:0] _T_57141; // @[Modules.scala 160:64:@2929.4]
  wire [13:0] _T_57142; // @[Modules.scala 160:64:@2930.4]
  wire [13:0] buffer_0_580; // @[Modules.scala 160:64:@2931.4]
  wire [14:0] _T_57144; // @[Modules.scala 160:64:@2933.4]
  wire [13:0] _T_57145; // @[Modules.scala 160:64:@2934.4]
  wire [13:0] buffer_0_581; // @[Modules.scala 160:64:@2935.4]
  wire [14:0] _T_57147; // @[Modules.scala 160:64:@2937.4]
  wire [13:0] _T_57148; // @[Modules.scala 160:64:@2938.4]
  wire [13:0] buffer_0_582; // @[Modules.scala 160:64:@2939.4]
  wire [14:0] _T_57150; // @[Modules.scala 160:64:@2941.4]
  wire [13:0] _T_57151; // @[Modules.scala 160:64:@2942.4]
  wire [13:0] buffer_0_583; // @[Modules.scala 160:64:@2943.4]
  wire [14:0] _T_57153; // @[Modules.scala 160:64:@2945.4]
  wire [13:0] _T_57154; // @[Modules.scala 160:64:@2946.4]
  wire [13:0] buffer_0_584; // @[Modules.scala 160:64:@2947.4]
  wire [14:0] _T_57156; // @[Modules.scala 166:64:@2949.4]
  wire [13:0] _T_57157; // @[Modules.scala 166:64:@2950.4]
  wire [13:0] buffer_0_585; // @[Modules.scala 166:64:@2951.4]
  wire [14:0] _T_57159; // @[Modules.scala 166:64:@2953.4]
  wire [13:0] _T_57160; // @[Modules.scala 166:64:@2954.4]
  wire [13:0] buffer_0_586; // @[Modules.scala 166:64:@2955.4]
  wire [14:0] _T_57162; // @[Modules.scala 166:64:@2957.4]
  wire [13:0] _T_57163; // @[Modules.scala 166:64:@2958.4]
  wire [13:0] buffer_0_587; // @[Modules.scala 166:64:@2959.4]
  wire [14:0] _T_57165; // @[Modules.scala 166:64:@2961.4]
  wire [13:0] _T_57166; // @[Modules.scala 166:64:@2962.4]
  wire [13:0] buffer_0_588; // @[Modules.scala 166:64:@2963.4]
  wire [14:0] _T_57168; // @[Modules.scala 166:64:@2965.4]
  wire [13:0] _T_57169; // @[Modules.scala 166:64:@2966.4]
  wire [13:0] buffer_0_589; // @[Modules.scala 166:64:@2967.4]
  wire [14:0] _T_57171; // @[Modules.scala 166:64:@2969.4]
  wire [13:0] _T_57172; // @[Modules.scala 166:64:@2970.4]
  wire [13:0] buffer_0_590; // @[Modules.scala 166:64:@2971.4]
  wire [14:0] _T_57174; // @[Modules.scala 166:64:@2973.4]
  wire [13:0] _T_57175; // @[Modules.scala 166:64:@2974.4]
  wire [13:0] buffer_0_591; // @[Modules.scala 166:64:@2975.4]
  wire [14:0] _T_57177; // @[Modules.scala 166:64:@2977.4]
  wire [13:0] _T_57178; // @[Modules.scala 166:64:@2978.4]
  wire [13:0] buffer_0_592; // @[Modules.scala 166:64:@2979.4]
  wire [14:0] _T_57180; // @[Modules.scala 166:64:@2981.4]
  wire [13:0] _T_57181; // @[Modules.scala 166:64:@2982.4]
  wire [13:0] buffer_0_593; // @[Modules.scala 166:64:@2983.4]
  wire [14:0] _T_57183; // @[Modules.scala 166:64:@2985.4]
  wire [13:0] _T_57184; // @[Modules.scala 166:64:@2986.4]
  wire [13:0] buffer_0_594; // @[Modules.scala 166:64:@2987.4]
  wire [14:0] _T_57186; // @[Modules.scala 166:64:@2989.4]
  wire [13:0] _T_57187; // @[Modules.scala 166:64:@2990.4]
  wire [13:0] buffer_0_595; // @[Modules.scala 166:64:@2991.4]
  wire [14:0] _T_57189; // @[Modules.scala 166:64:@2993.4]
  wire [13:0] _T_57190; // @[Modules.scala 166:64:@2994.4]
  wire [13:0] buffer_0_596; // @[Modules.scala 166:64:@2995.4]
  wire [14:0] _T_57192; // @[Modules.scala 166:64:@2997.4]
  wire [13:0] _T_57193; // @[Modules.scala 166:64:@2998.4]
  wire [13:0] buffer_0_597; // @[Modules.scala 166:64:@2999.4]
  wire [14:0] _T_57195; // @[Modules.scala 172:66:@3001.4]
  wire [13:0] _T_57196; // @[Modules.scala 172:66:@3002.4]
  wire [13:0] buffer_0_598; // @[Modules.scala 172:66:@3003.4]
  wire [14:0] _T_57198; // @[Modules.scala 166:64:@3005.4]
  wire [13:0] _T_57199; // @[Modules.scala 166:64:@3006.4]
  wire [13:0] buffer_0_599; // @[Modules.scala 166:64:@3007.4]
  wire [14:0] _T_57201; // @[Modules.scala 166:64:@3009.4]
  wire [13:0] _T_57202; // @[Modules.scala 166:64:@3010.4]
  wire [13:0] buffer_0_600; // @[Modules.scala 166:64:@3011.4]
  wire [14:0] _T_57204; // @[Modules.scala 160:64:@3013.4]
  wire [13:0] _T_57205; // @[Modules.scala 160:64:@3014.4]
  wire [13:0] buffer_0_601; // @[Modules.scala 160:64:@3015.4]
  wire [14:0] _T_57207; // @[Modules.scala 172:66:@3017.4]
  wire [13:0] _T_57208; // @[Modules.scala 172:66:@3018.4]
  wire [13:0] buffer_0_602; // @[Modules.scala 172:66:@3019.4]
  wire [5:0] _T_57225; // @[Modules.scala 143:74:@3214.4]
  wire [4:0] _T_57227; // @[Modules.scala 144:80:@3215.4]
  wire [5:0] _GEN_76; // @[Modules.scala 143:103:@3216.4]
  wire [6:0] _T_57228; // @[Modules.scala 143:103:@3216.4]
  wire [5:0] _T_57229; // @[Modules.scala 143:103:@3217.4]
  wire [5:0] _T_57230; // @[Modules.scala 143:103:@3218.4]
  wire [5:0] _T_57232; // @[Modules.scala 143:74:@3220.4]
  wire [5:0] _T_57234; // @[Modules.scala 144:80:@3221.4]
  wire [6:0] _T_57235; // @[Modules.scala 143:103:@3222.4]
  wire [5:0] _T_57236; // @[Modules.scala 143:103:@3223.4]
  wire [5:0] _T_57237; // @[Modules.scala 143:103:@3224.4]
  wire [4:0] _T_57239; // @[Modules.scala 143:74:@3226.4]
  wire [4:0] _T_57241; // @[Modules.scala 144:80:@3227.4]
  wire [5:0] _T_57242; // @[Modules.scala 143:103:@3228.4]
  wire [4:0] _T_57243; // @[Modules.scala 143:103:@3229.4]
  wire [4:0] _T_57244; // @[Modules.scala 143:103:@3230.4]
  wire [4:0] _T_57248; // @[Modules.scala 144:80:@3233.4]
  wire [5:0] _GEN_77; // @[Modules.scala 143:103:@3234.4]
  wire [6:0] _T_57249; // @[Modules.scala 143:103:@3234.4]
  wire [5:0] _T_57250; // @[Modules.scala 143:103:@3235.4]
  wire [5:0] _T_57251; // @[Modules.scala 143:103:@3236.4]
  wire [4:0] _T_57253; // @[Modules.scala 143:74:@3238.4]
  wire [4:0] _T_57255; // @[Modules.scala 144:80:@3239.4]
  wire [5:0] _T_57256; // @[Modules.scala 143:103:@3240.4]
  wire [4:0] _T_57257; // @[Modules.scala 143:103:@3241.4]
  wire [4:0] _T_57258; // @[Modules.scala 143:103:@3242.4]
  wire [4:0] _T_57260; // @[Modules.scala 143:74:@3244.4]
  wire [4:0] _T_57262; // @[Modules.scala 144:80:@3245.4]
  wire [5:0] _T_57263; // @[Modules.scala 143:103:@3246.4]
  wire [4:0] _T_57264; // @[Modules.scala 143:103:@3247.4]
  wire [4:0] _T_57265; // @[Modules.scala 143:103:@3248.4]
  wire [4:0] _T_57267; // @[Modules.scala 143:74:@3250.4]
  wire [5:0] _GEN_78; // @[Modules.scala 143:103:@3252.4]
  wire [6:0] _T_57270; // @[Modules.scala 143:103:@3252.4]
  wire [5:0] _T_57271; // @[Modules.scala 143:103:@3253.4]
  wire [5:0] _T_57272; // @[Modules.scala 143:103:@3254.4]
  wire [4:0] _T_57274; // @[Modules.scala 143:74:@3256.4]
  wire [4:0] _T_57276; // @[Modules.scala 144:80:@3257.4]
  wire [5:0] _T_57277; // @[Modules.scala 143:103:@3258.4]
  wire [4:0] _T_57278; // @[Modules.scala 143:103:@3259.4]
  wire [4:0] _T_57279; // @[Modules.scala 143:103:@3260.4]
  wire [4:0] _T_57281; // @[Modules.scala 143:74:@3262.4]
  wire [5:0] _GEN_79; // @[Modules.scala 143:103:@3264.4]
  wire [6:0] _T_57284; // @[Modules.scala 143:103:@3264.4]
  wire [5:0] _T_57285; // @[Modules.scala 143:103:@3265.4]
  wire [5:0] _T_57286; // @[Modules.scala 143:103:@3266.4]
  wire [4:0] _T_57288; // @[Modules.scala 143:74:@3268.4]
  wire [5:0] _GEN_80; // @[Modules.scala 143:103:@3270.4]
  wire [6:0] _T_57291; // @[Modules.scala 143:103:@3270.4]
  wire [5:0] _T_57292; // @[Modules.scala 143:103:@3271.4]
  wire [5:0] _T_57293; // @[Modules.scala 143:103:@3272.4]
  wire [4:0] _T_57297; // @[Modules.scala 144:80:@3275.4]
  wire [5:0] _GEN_81; // @[Modules.scala 143:103:@3276.4]
  wire [6:0] _T_57298; // @[Modules.scala 143:103:@3276.4]
  wire [5:0] _T_57299; // @[Modules.scala 143:103:@3277.4]
  wire [5:0] _T_57300; // @[Modules.scala 143:103:@3278.4]
  wire [4:0] _T_57302; // @[Modules.scala 143:74:@3280.4]
  wire [4:0] _T_57304; // @[Modules.scala 144:80:@3281.4]
  wire [5:0] _T_57305; // @[Modules.scala 143:103:@3282.4]
  wire [4:0] _T_57306; // @[Modules.scala 143:103:@3283.4]
  wire [4:0] _T_57307; // @[Modules.scala 143:103:@3284.4]
  wire [4:0] _T_57309; // @[Modules.scala 143:74:@3286.4]
  wire [4:0] _T_57311; // @[Modules.scala 144:80:@3287.4]
  wire [5:0] _T_57312; // @[Modules.scala 143:103:@3288.4]
  wire [4:0] _T_57313; // @[Modules.scala 143:103:@3289.4]
  wire [4:0] _T_57314; // @[Modules.scala 143:103:@3290.4]
  wire [4:0] _T_57316; // @[Modules.scala 143:74:@3292.4]
  wire [4:0] _T_57318; // @[Modules.scala 144:80:@3293.4]
  wire [5:0] _T_57319; // @[Modules.scala 143:103:@3294.4]
  wire [4:0] _T_57320; // @[Modules.scala 143:103:@3295.4]
  wire [4:0] _T_57321; // @[Modules.scala 143:103:@3296.4]
  wire [4:0] _T_57323; // @[Modules.scala 143:74:@3298.4]
  wire [4:0] _T_57325; // @[Modules.scala 144:80:@3299.4]
  wire [5:0] _T_57326; // @[Modules.scala 143:103:@3300.4]
  wire [4:0] _T_57327; // @[Modules.scala 143:103:@3301.4]
  wire [4:0] _T_57328; // @[Modules.scala 143:103:@3302.4]
  wire [4:0] _T_57330; // @[Modules.scala 143:74:@3304.4]
  wire [4:0] _T_57332; // @[Modules.scala 144:80:@3305.4]
  wire [5:0] _T_57333; // @[Modules.scala 143:103:@3306.4]
  wire [4:0] _T_57334; // @[Modules.scala 143:103:@3307.4]
  wire [4:0] _T_57335; // @[Modules.scala 143:103:@3308.4]
  wire [4:0] _T_57337; // @[Modules.scala 143:74:@3310.4]
  wire [4:0] _T_57339; // @[Modules.scala 144:80:@3311.4]
  wire [5:0] _T_57340; // @[Modules.scala 143:103:@3312.4]
  wire [4:0] _T_57341; // @[Modules.scala 143:103:@3313.4]
  wire [4:0] _T_57342; // @[Modules.scala 143:103:@3314.4]
  wire [6:0] _T_57347; // @[Modules.scala 143:103:@3318.4]
  wire [5:0] _T_57348; // @[Modules.scala 143:103:@3319.4]
  wire [5:0] _T_57349; // @[Modules.scala 143:103:@3320.4]
  wire [6:0] _T_57354; // @[Modules.scala 143:103:@3324.4]
  wire [5:0] _T_57355; // @[Modules.scala 143:103:@3325.4]
  wire [5:0] _T_57356; // @[Modules.scala 143:103:@3326.4]
  wire [6:0] _T_57361; // @[Modules.scala 143:103:@3330.4]
  wire [5:0] _T_57362; // @[Modules.scala 143:103:@3331.4]
  wire [5:0] _T_57363; // @[Modules.scala 143:103:@3332.4]
  wire [6:0] _T_57368; // @[Modules.scala 143:103:@3336.4]
  wire [5:0] _T_57369; // @[Modules.scala 143:103:@3337.4]
  wire [5:0] _T_57370; // @[Modules.scala 143:103:@3338.4]
  wire [6:0] _T_57375; // @[Modules.scala 143:103:@3342.4]
  wire [5:0] _T_57376; // @[Modules.scala 143:103:@3343.4]
  wire [5:0] _T_57377; // @[Modules.scala 143:103:@3344.4]
  wire [4:0] _T_57379; // @[Modules.scala 143:74:@3346.4]
  wire [4:0] _T_57381; // @[Modules.scala 144:80:@3347.4]
  wire [5:0] _T_57382; // @[Modules.scala 143:103:@3348.4]
  wire [4:0] _T_57383; // @[Modules.scala 143:103:@3349.4]
  wire [4:0] _T_57384; // @[Modules.scala 143:103:@3350.4]
  wire [4:0] _T_57386; // @[Modules.scala 143:74:@3352.4]
  wire [4:0] _T_57388; // @[Modules.scala 144:80:@3353.4]
  wire [5:0] _T_57389; // @[Modules.scala 143:103:@3354.4]
  wire [4:0] _T_57390; // @[Modules.scala 143:103:@3355.4]
  wire [4:0] _T_57391; // @[Modules.scala 143:103:@3356.4]
  wire [4:0] _T_57393; // @[Modules.scala 143:74:@3358.4]
  wire [4:0] _T_57395; // @[Modules.scala 144:80:@3359.4]
  wire [5:0] _T_57396; // @[Modules.scala 143:103:@3360.4]
  wire [4:0] _T_57397; // @[Modules.scala 143:103:@3361.4]
  wire [4:0] _T_57398; // @[Modules.scala 143:103:@3362.4]
  wire [4:0] _T_57400; // @[Modules.scala 143:74:@3364.4]
  wire [4:0] _T_57402; // @[Modules.scala 144:80:@3365.4]
  wire [5:0] _T_57403; // @[Modules.scala 143:103:@3366.4]
  wire [4:0] _T_57404; // @[Modules.scala 143:103:@3367.4]
  wire [4:0] _T_57405; // @[Modules.scala 143:103:@3368.4]
  wire [4:0] _T_57409; // @[Modules.scala 144:80:@3371.4]
  wire [5:0] _GEN_83; // @[Modules.scala 143:103:@3372.4]
  wire [6:0] _T_57410; // @[Modules.scala 143:103:@3372.4]
  wire [5:0] _T_57411; // @[Modules.scala 143:103:@3373.4]
  wire [5:0] _T_57412; // @[Modules.scala 143:103:@3374.4]
  wire [4:0] _T_57414; // @[Modules.scala 143:74:@3376.4]
  wire [4:0] _T_57416; // @[Modules.scala 144:80:@3377.4]
  wire [5:0] _T_57417; // @[Modules.scala 143:103:@3378.4]
  wire [4:0] _T_57418; // @[Modules.scala 143:103:@3379.4]
  wire [4:0] _T_57419; // @[Modules.scala 143:103:@3380.4]
  wire [4:0] _T_57421; // @[Modules.scala 143:74:@3382.4]
  wire [4:0] _T_57423; // @[Modules.scala 144:80:@3383.4]
  wire [5:0] _T_57424; // @[Modules.scala 143:103:@3384.4]
  wire [4:0] _T_57425; // @[Modules.scala 143:103:@3385.4]
  wire [4:0] _T_57426; // @[Modules.scala 143:103:@3386.4]
  wire [4:0] _T_57428; // @[Modules.scala 143:74:@3388.4]
  wire [4:0] _T_57430; // @[Modules.scala 144:80:@3389.4]
  wire [5:0] _T_57431; // @[Modules.scala 143:103:@3390.4]
  wire [4:0] _T_57432; // @[Modules.scala 143:103:@3391.4]
  wire [4:0] _T_57433; // @[Modules.scala 143:103:@3392.4]
  wire [4:0] _T_57435; // @[Modules.scala 143:74:@3394.4]
  wire [5:0] _GEN_84; // @[Modules.scala 143:103:@3396.4]
  wire [6:0] _T_57438; // @[Modules.scala 143:103:@3396.4]
  wire [5:0] _T_57439; // @[Modules.scala 143:103:@3397.4]
  wire [5:0] _T_57440; // @[Modules.scala 143:103:@3398.4]
  wire [5:0] _T_57442; // @[Modules.scala 143:74:@3400.4]
  wire [6:0] _T_57445; // @[Modules.scala 143:103:@3402.4]
  wire [5:0] _T_57446; // @[Modules.scala 143:103:@3403.4]
  wire [5:0] _T_57447; // @[Modules.scala 143:103:@3404.4]
  wire [5:0] _T_57449; // @[Modules.scala 143:74:@3406.4]
  wire [5:0] _T_57451; // @[Modules.scala 144:80:@3407.4]
  wire [6:0] _T_57452; // @[Modules.scala 143:103:@3408.4]
  wire [5:0] _T_57453; // @[Modules.scala 143:103:@3409.4]
  wire [5:0] _T_57454; // @[Modules.scala 143:103:@3410.4]
  wire [5:0] _T_57456; // @[Modules.scala 143:74:@3412.4]
  wire [5:0] _T_57458; // @[Modules.scala 144:80:@3413.4]
  wire [6:0] _T_57459; // @[Modules.scala 143:103:@3414.4]
  wire [5:0] _T_57460; // @[Modules.scala 143:103:@3415.4]
  wire [5:0] _T_57461; // @[Modules.scala 143:103:@3416.4]
  wire [6:0] _T_57466; // @[Modules.scala 143:103:@3420.4]
  wire [5:0] _T_57467; // @[Modules.scala 143:103:@3421.4]
  wire [5:0] _T_57468; // @[Modules.scala 143:103:@3422.4]
  wire [6:0] _T_57473; // @[Modules.scala 143:103:@3426.4]
  wire [5:0] _T_57474; // @[Modules.scala 143:103:@3427.4]
  wire [5:0] _T_57475; // @[Modules.scala 143:103:@3428.4]
  wire [6:0] _T_57480; // @[Modules.scala 143:103:@3432.4]
  wire [5:0] _T_57481; // @[Modules.scala 143:103:@3433.4]
  wire [5:0] _T_57482; // @[Modules.scala 143:103:@3434.4]
  wire [4:0] _T_57486; // @[Modules.scala 144:80:@3437.4]
  wire [5:0] _GEN_85; // @[Modules.scala 143:103:@3438.4]
  wire [6:0] _T_57487; // @[Modules.scala 143:103:@3438.4]
  wire [5:0] _T_57488; // @[Modules.scala 143:103:@3439.4]
  wire [5:0] _T_57489; // @[Modules.scala 143:103:@3440.4]
  wire [5:0] _T_57498; // @[Modules.scala 143:74:@3448.4]
  wire [6:0] _T_57501; // @[Modules.scala 143:103:@3450.4]
  wire [5:0] _T_57502; // @[Modules.scala 143:103:@3451.4]
  wire [5:0] _T_57503; // @[Modules.scala 143:103:@3452.4]
  wire [5:0] _T_57507; // @[Modules.scala 144:80:@3455.4]
  wire [6:0] _T_57508; // @[Modules.scala 143:103:@3456.4]
  wire [5:0] _T_57509; // @[Modules.scala 143:103:@3457.4]
  wire [5:0] _T_57510; // @[Modules.scala 143:103:@3458.4]
  wire [5:0] _T_57512; // @[Modules.scala 143:74:@3460.4]
  wire [5:0] _T_57514; // @[Modules.scala 144:80:@3461.4]
  wire [6:0] _T_57515; // @[Modules.scala 143:103:@3462.4]
  wire [5:0] _T_57516; // @[Modules.scala 143:103:@3463.4]
  wire [5:0] _T_57517; // @[Modules.scala 143:103:@3464.4]
  wire [4:0] _T_57521; // @[Modules.scala 144:80:@3467.4]
  wire [5:0] _GEN_86; // @[Modules.scala 143:103:@3468.4]
  wire [6:0] _T_57522; // @[Modules.scala 143:103:@3468.4]
  wire [5:0] _T_57523; // @[Modules.scala 143:103:@3469.4]
  wire [5:0] _T_57524; // @[Modules.scala 143:103:@3470.4]
  wire [5:0] _T_57526; // @[Modules.scala 143:74:@3472.4]
  wire [6:0] _T_57529; // @[Modules.scala 143:103:@3474.4]
  wire [5:0] _T_57530; // @[Modules.scala 143:103:@3475.4]
  wire [5:0] _T_57531; // @[Modules.scala 143:103:@3476.4]
  wire [5:0] _T_57533; // @[Modules.scala 143:74:@3478.4]
  wire [5:0] _T_57535; // @[Modules.scala 144:80:@3479.4]
  wire [6:0] _T_57536; // @[Modules.scala 143:103:@3480.4]
  wire [5:0] _T_57537; // @[Modules.scala 143:103:@3481.4]
  wire [5:0] _T_57538; // @[Modules.scala 143:103:@3482.4]
  wire [5:0] _T_57540; // @[Modules.scala 143:74:@3484.4]
  wire [5:0] _T_57542; // @[Modules.scala 144:80:@3485.4]
  wire [6:0] _T_57543; // @[Modules.scala 143:103:@3486.4]
  wire [5:0] _T_57544; // @[Modules.scala 143:103:@3487.4]
  wire [5:0] _T_57545; // @[Modules.scala 143:103:@3488.4]
  wire [5:0] _T_57556; // @[Modules.scala 144:80:@3497.4]
  wire [6:0] _T_57557; // @[Modules.scala 143:103:@3498.4]
  wire [5:0] _T_57558; // @[Modules.scala 143:103:@3499.4]
  wire [5:0] _T_57559; // @[Modules.scala 143:103:@3500.4]
  wire [4:0] _T_57561; // @[Modules.scala 143:74:@3502.4]
  wire [4:0] _T_57563; // @[Modules.scala 144:80:@3503.4]
  wire [5:0] _T_57564; // @[Modules.scala 143:103:@3504.4]
  wire [4:0] _T_57565; // @[Modules.scala 143:103:@3505.4]
  wire [4:0] _T_57566; // @[Modules.scala 143:103:@3506.4]
  wire [5:0] _T_57571; // @[Modules.scala 143:103:@3510.4]
  wire [4:0] _T_57572; // @[Modules.scala 143:103:@3511.4]
  wire [4:0] _T_57573; // @[Modules.scala 143:103:@3512.4]
  wire [4:0] _T_57575; // @[Modules.scala 143:74:@3514.4]
  wire [5:0] _GEN_87; // @[Modules.scala 143:103:@3516.4]
  wire [6:0] _T_57578; // @[Modules.scala 143:103:@3516.4]
  wire [5:0] _T_57579; // @[Modules.scala 143:103:@3517.4]
  wire [5:0] _T_57580; // @[Modules.scala 143:103:@3518.4]
  wire [5:0] _T_57585; // @[Modules.scala 143:103:@3522.4]
  wire [4:0] _T_57586; // @[Modules.scala 143:103:@3523.4]
  wire [4:0] _T_57587; // @[Modules.scala 143:103:@3524.4]
  wire [5:0] _T_57592; // @[Modules.scala 143:103:@3528.4]
  wire [4:0] _T_57593; // @[Modules.scala 143:103:@3529.4]
  wire [4:0] _T_57594; // @[Modules.scala 143:103:@3530.4]
  wire [4:0] _T_57596; // @[Modules.scala 143:74:@3532.4]
  wire [5:0] _GEN_88; // @[Modules.scala 143:103:@3534.4]
  wire [6:0] _T_57599; // @[Modules.scala 143:103:@3534.4]
  wire [5:0] _T_57600; // @[Modules.scala 143:103:@3535.4]
  wire [5:0] _T_57601; // @[Modules.scala 143:103:@3536.4]
  wire [4:0] _T_57619; // @[Modules.scala 144:80:@3551.4]
  wire [5:0] _GEN_90; // @[Modules.scala 143:103:@3552.4]
  wire [6:0] _T_57620; // @[Modules.scala 143:103:@3552.4]
  wire [5:0] _T_57621; // @[Modules.scala 143:103:@3553.4]
  wire [5:0] _T_57622; // @[Modules.scala 143:103:@3554.4]
  wire [5:0] _T_57626; // @[Modules.scala 144:80:@3557.4]
  wire [6:0] _T_57627; // @[Modules.scala 143:103:@3558.4]
  wire [5:0] _T_57628; // @[Modules.scala 143:103:@3559.4]
  wire [5:0] _T_57629; // @[Modules.scala 143:103:@3560.4]
  wire [5:0] _T_57631; // @[Modules.scala 143:74:@3562.4]
  wire [5:0] _T_57633; // @[Modules.scala 144:80:@3563.4]
  wire [6:0] _T_57634; // @[Modules.scala 143:103:@3564.4]
  wire [5:0] _T_57635; // @[Modules.scala 143:103:@3565.4]
  wire [5:0] _T_57636; // @[Modules.scala 143:103:@3566.4]
  wire [5:0] _T_57638; // @[Modules.scala 143:74:@3568.4]
  wire [5:0] _T_57640; // @[Modules.scala 144:80:@3569.4]
  wire [6:0] _T_57641; // @[Modules.scala 143:103:@3570.4]
  wire [5:0] _T_57642; // @[Modules.scala 143:103:@3571.4]
  wire [5:0] _T_57643; // @[Modules.scala 143:103:@3572.4]
  wire [5:0] _T_57645; // @[Modules.scala 143:74:@3574.4]
  wire [5:0] _GEN_92; // @[Modules.scala 143:103:@3576.4]
  wire [6:0] _T_57648; // @[Modules.scala 143:103:@3576.4]
  wire [5:0] _T_57649; // @[Modules.scala 143:103:@3577.4]
  wire [5:0] _T_57650; // @[Modules.scala 143:103:@3578.4]
  wire [5:0] _T_57655; // @[Modules.scala 143:103:@3582.4]
  wire [4:0] _T_57656; // @[Modules.scala 143:103:@3583.4]
  wire [4:0] _T_57657; // @[Modules.scala 143:103:@3584.4]
  wire [5:0] _T_57662; // @[Modules.scala 143:103:@3588.4]
  wire [4:0] _T_57663; // @[Modules.scala 143:103:@3589.4]
  wire [4:0] _T_57664; // @[Modules.scala 143:103:@3590.4]
  wire [5:0] _T_57669; // @[Modules.scala 143:103:@3594.4]
  wire [4:0] _T_57670; // @[Modules.scala 143:103:@3595.4]
  wire [4:0] _T_57671; // @[Modules.scala 143:103:@3596.4]
  wire [5:0] _T_57675; // @[Modules.scala 144:80:@3599.4]
  wire [5:0] _GEN_93; // @[Modules.scala 143:103:@3600.4]
  wire [6:0] _T_57676; // @[Modules.scala 143:103:@3600.4]
  wire [5:0] _T_57677; // @[Modules.scala 143:103:@3601.4]
  wire [5:0] _T_57678; // @[Modules.scala 143:103:@3602.4]
  wire [4:0] _T_57701; // @[Modules.scala 143:74:@3622.4]
  wire [5:0] _T_57704; // @[Modules.scala 143:103:@3624.4]
  wire [4:0] _T_57705; // @[Modules.scala 143:103:@3625.4]
  wire [4:0] _T_57706; // @[Modules.scala 143:103:@3626.4]
  wire [5:0] _T_57708; // @[Modules.scala 143:74:@3628.4]
  wire [5:0] _T_57710; // @[Modules.scala 144:80:@3629.4]
  wire [6:0] _T_57711; // @[Modules.scala 143:103:@3630.4]
  wire [5:0] _T_57712; // @[Modules.scala 143:103:@3631.4]
  wire [5:0] _T_57713; // @[Modules.scala 143:103:@3632.4]
  wire [5:0] _T_57715; // @[Modules.scala 143:74:@3634.4]
  wire [5:0] _T_57717; // @[Modules.scala 144:80:@3635.4]
  wire [6:0] _T_57718; // @[Modules.scala 143:103:@3636.4]
  wire [5:0] _T_57719; // @[Modules.scala 143:103:@3637.4]
  wire [5:0] _T_57720; // @[Modules.scala 143:103:@3638.4]
  wire [5:0] _T_57722; // @[Modules.scala 143:74:@3640.4]
  wire [5:0] _T_57724; // @[Modules.scala 144:80:@3641.4]
  wire [6:0] _T_57725; // @[Modules.scala 143:103:@3642.4]
  wire [5:0] _T_57726; // @[Modules.scala 143:103:@3643.4]
  wire [5:0] _T_57727; // @[Modules.scala 143:103:@3644.4]
  wire [5:0] _T_57729; // @[Modules.scala 143:74:@3646.4]
  wire [5:0] _GEN_94; // @[Modules.scala 143:103:@3648.4]
  wire [6:0] _T_57732; // @[Modules.scala 143:103:@3648.4]
  wire [5:0] _T_57733; // @[Modules.scala 143:103:@3649.4]
  wire [5:0] _T_57734; // @[Modules.scala 143:103:@3650.4]
  wire [5:0] _T_57736; // @[Modules.scala 143:74:@3652.4]
  wire [5:0] _T_57738; // @[Modules.scala 144:80:@3653.4]
  wire [6:0] _T_57739; // @[Modules.scala 143:103:@3654.4]
  wire [5:0] _T_57740; // @[Modules.scala 143:103:@3655.4]
  wire [5:0] _T_57741; // @[Modules.scala 143:103:@3656.4]
  wire [4:0] _T_57757; // @[Modules.scala 143:74:@3670.4]
  wire [4:0] _T_57759; // @[Modules.scala 144:80:@3671.4]
  wire [5:0] _T_57760; // @[Modules.scala 143:103:@3672.4]
  wire [4:0] _T_57761; // @[Modules.scala 143:103:@3673.4]
  wire [4:0] _T_57762; // @[Modules.scala 143:103:@3674.4]
  wire [5:0] _T_57764; // @[Modules.scala 143:74:@3676.4]
  wire [6:0] _T_57767; // @[Modules.scala 143:103:@3678.4]
  wire [5:0] _T_57768; // @[Modules.scala 143:103:@3679.4]
  wire [5:0] _T_57769; // @[Modules.scala 143:103:@3680.4]
  wire [6:0] _T_57774; // @[Modules.scala 143:103:@3684.4]
  wire [5:0] _T_57775; // @[Modules.scala 143:103:@3685.4]
  wire [5:0] _T_57776; // @[Modules.scala 143:103:@3686.4]
  wire [6:0] _T_57781; // @[Modules.scala 143:103:@3690.4]
  wire [5:0] _T_57782; // @[Modules.scala 143:103:@3691.4]
  wire [5:0] _T_57783; // @[Modules.scala 143:103:@3692.4]
  wire [4:0] _T_57787; // @[Modules.scala 144:80:@3695.4]
  wire [5:0] _GEN_95; // @[Modules.scala 143:103:@3696.4]
  wire [6:0] _T_57788; // @[Modules.scala 143:103:@3696.4]
  wire [5:0] _T_57789; // @[Modules.scala 143:103:@3697.4]
  wire [5:0] _T_57790; // @[Modules.scala 143:103:@3698.4]
  wire [4:0] _T_57794; // @[Modules.scala 144:80:@3701.4]
  wire [5:0] _T_57795; // @[Modules.scala 143:103:@3702.4]
  wire [4:0] _T_57796; // @[Modules.scala 143:103:@3703.4]
  wire [4:0] _T_57797; // @[Modules.scala 143:103:@3704.4]
  wire [5:0] _T_57799; // @[Modules.scala 143:74:@3706.4]
  wire [6:0] _T_57802; // @[Modules.scala 143:103:@3708.4]
  wire [5:0] _T_57803; // @[Modules.scala 143:103:@3709.4]
  wire [5:0] _T_57804; // @[Modules.scala 143:103:@3710.4]
  wire [5:0] _T_57806; // @[Modules.scala 143:74:@3712.4]
  wire [5:0] _T_57808; // @[Modules.scala 144:80:@3713.4]
  wire [6:0] _T_57809; // @[Modules.scala 143:103:@3714.4]
  wire [5:0] _T_57810; // @[Modules.scala 143:103:@3715.4]
  wire [5:0] _T_57811; // @[Modules.scala 143:103:@3716.4]
  wire [5:0] _T_57813; // @[Modules.scala 143:74:@3718.4]
  wire [5:0] _T_57815; // @[Modules.scala 144:80:@3719.4]
  wire [6:0] _T_57816; // @[Modules.scala 143:103:@3720.4]
  wire [5:0] _T_57817; // @[Modules.scala 143:103:@3721.4]
  wire [5:0] _T_57818; // @[Modules.scala 143:103:@3722.4]
  wire [4:0] _T_57848; // @[Modules.scala 143:74:@3748.4]
  wire [5:0] _T_57850; // @[Modules.scala 144:80:@3749.4]
  wire [5:0] _GEN_96; // @[Modules.scala 143:103:@3750.4]
  wire [6:0] _T_57851; // @[Modules.scala 143:103:@3750.4]
  wire [5:0] _T_57852; // @[Modules.scala 143:103:@3751.4]
  wire [5:0] _T_57853; // @[Modules.scala 143:103:@3752.4]
  wire [5:0] _T_57857; // @[Modules.scala 144:80:@3755.4]
  wire [6:0] _T_57858; // @[Modules.scala 143:103:@3756.4]
  wire [5:0] _T_57859; // @[Modules.scala 143:103:@3757.4]
  wire [5:0] _T_57860; // @[Modules.scala 143:103:@3758.4]
  wire [5:0] _T_57864; // @[Modules.scala 144:80:@3761.4]
  wire [6:0] _T_57865; // @[Modules.scala 143:103:@3762.4]
  wire [5:0] _T_57866; // @[Modules.scala 143:103:@3763.4]
  wire [5:0] _T_57867; // @[Modules.scala 143:103:@3764.4]
  wire [4:0] _T_57869; // @[Modules.scala 143:74:@3766.4]
  wire [5:0] _T_57872; // @[Modules.scala 143:103:@3768.4]
  wire [4:0] _T_57873; // @[Modules.scala 143:103:@3769.4]
  wire [4:0] _T_57874; // @[Modules.scala 143:103:@3770.4]
  wire [6:0] _T_57886; // @[Modules.scala 143:103:@3780.4]
  wire [5:0] _T_57887; // @[Modules.scala 143:103:@3781.4]
  wire [5:0] _T_57888; // @[Modules.scala 143:103:@3782.4]
  wire [5:0] _T_57890; // @[Modules.scala 143:74:@3784.4]
  wire [5:0] _T_57892; // @[Modules.scala 144:80:@3785.4]
  wire [6:0] _T_57893; // @[Modules.scala 143:103:@3786.4]
  wire [5:0] _T_57894; // @[Modules.scala 143:103:@3787.4]
  wire [5:0] _T_57895; // @[Modules.scala 143:103:@3788.4]
  wire [5:0] _T_57897; // @[Modules.scala 143:74:@3790.4]
  wire [5:0] _T_57899; // @[Modules.scala 144:80:@3791.4]
  wire [6:0] _T_57900; // @[Modules.scala 143:103:@3792.4]
  wire [5:0] _T_57901; // @[Modules.scala 143:103:@3793.4]
  wire [5:0] _T_57902; // @[Modules.scala 143:103:@3794.4]
  wire [5:0] _T_57904; // @[Modules.scala 143:74:@3796.4]
  wire [5:0] _GEN_97; // @[Modules.scala 143:103:@3798.4]
  wire [6:0] _T_57907; // @[Modules.scala 143:103:@3798.4]
  wire [5:0] _T_57908; // @[Modules.scala 143:103:@3799.4]
  wire [5:0] _T_57909; // @[Modules.scala 143:103:@3800.4]
  wire [5:0] _T_57927; // @[Modules.scala 144:80:@3815.4]
  wire [5:0] _GEN_98; // @[Modules.scala 143:103:@3816.4]
  wire [6:0] _T_57928; // @[Modules.scala 143:103:@3816.4]
  wire [5:0] _T_57929; // @[Modules.scala 143:103:@3817.4]
  wire [5:0] _T_57930; // @[Modules.scala 143:103:@3818.4]
  wire [5:0] _T_57941; // @[Modules.scala 144:80:@3827.4]
  wire [6:0] _T_57942; // @[Modules.scala 143:103:@3828.4]
  wire [5:0] _T_57943; // @[Modules.scala 143:103:@3829.4]
  wire [5:0] _T_57944; // @[Modules.scala 143:103:@3830.4]
  wire [5:0] _T_57949; // @[Modules.scala 143:103:@3834.4]
  wire [4:0] _T_57950; // @[Modules.scala 143:103:@3835.4]
  wire [4:0] _T_57951; // @[Modules.scala 143:103:@3836.4]
  wire [5:0] _T_57956; // @[Modules.scala 143:103:@3840.4]
  wire [4:0] _T_57957; // @[Modules.scala 143:103:@3841.4]
  wire [4:0] _T_57958; // @[Modules.scala 143:103:@3842.4]
  wire [5:0] _T_57962; // @[Modules.scala 144:80:@3845.4]
  wire [5:0] _GEN_99; // @[Modules.scala 143:103:@3846.4]
  wire [6:0] _T_57963; // @[Modules.scala 143:103:@3846.4]
  wire [5:0] _T_57964; // @[Modules.scala 143:103:@3847.4]
  wire [5:0] _T_57965; // @[Modules.scala 143:103:@3848.4]
  wire [6:0] _T_57970; // @[Modules.scala 143:103:@3852.4]
  wire [5:0] _T_57971; // @[Modules.scala 143:103:@3853.4]
  wire [5:0] _T_57972; // @[Modules.scala 143:103:@3854.4]
  wire [5:0] _T_57976; // @[Modules.scala 144:80:@3857.4]
  wire [6:0] _T_57977; // @[Modules.scala 143:103:@3858.4]
  wire [5:0] _T_57978; // @[Modules.scala 143:103:@3859.4]
  wire [5:0] _T_57979; // @[Modules.scala 143:103:@3860.4]
  wire [5:0] _T_57981; // @[Modules.scala 143:74:@3862.4]
  wire [5:0] _T_57983; // @[Modules.scala 144:80:@3863.4]
  wire [6:0] _T_57984; // @[Modules.scala 143:103:@3864.4]
  wire [5:0] _T_57985; // @[Modules.scala 143:103:@3865.4]
  wire [5:0] _T_57986; // @[Modules.scala 143:103:@3866.4]
  wire [5:0] _T_57988; // @[Modules.scala 143:74:@3868.4]
  wire [5:0] _T_57990; // @[Modules.scala 144:80:@3869.4]
  wire [6:0] _T_57991; // @[Modules.scala 143:103:@3870.4]
  wire [5:0] _T_57992; // @[Modules.scala 143:103:@3871.4]
  wire [5:0] _T_57993; // @[Modules.scala 143:103:@3872.4]
  wire [5:0] _T_57998; // @[Modules.scala 143:103:@3876.4]
  wire [4:0] _T_57999; // @[Modules.scala 143:103:@3877.4]
  wire [4:0] _T_58000; // @[Modules.scala 143:103:@3878.4]
  wire [5:0] _T_58005; // @[Modules.scala 143:103:@3882.4]
  wire [4:0] _T_58006; // @[Modules.scala 143:103:@3883.4]
  wire [4:0] _T_58007; // @[Modules.scala 143:103:@3884.4]
  wire [5:0] _T_58009; // @[Modules.scala 143:74:@3886.4]
  wire [5:0] _T_58011; // @[Modules.scala 144:80:@3887.4]
  wire [6:0] _T_58012; // @[Modules.scala 143:103:@3888.4]
  wire [5:0] _T_58013; // @[Modules.scala 143:103:@3889.4]
  wire [5:0] _T_58014; // @[Modules.scala 143:103:@3890.4]
  wire [5:0] _T_58018; // @[Modules.scala 144:80:@3893.4]
  wire [6:0] _T_58019; // @[Modules.scala 143:103:@3894.4]
  wire [5:0] _T_58020; // @[Modules.scala 143:103:@3895.4]
  wire [5:0] _T_58021; // @[Modules.scala 143:103:@3896.4]
  wire [5:0] _T_58025; // @[Modules.scala 144:80:@3899.4]
  wire [6:0] _T_58026; // @[Modules.scala 143:103:@3900.4]
  wire [5:0] _T_58027; // @[Modules.scala 143:103:@3901.4]
  wire [5:0] _T_58028; // @[Modules.scala 143:103:@3902.4]
  wire [5:0] _T_58032; // @[Modules.scala 144:80:@3905.4]
  wire [5:0] _GEN_100; // @[Modules.scala 143:103:@3906.4]
  wire [6:0] _T_58033; // @[Modules.scala 143:103:@3906.4]
  wire [5:0] _T_58034; // @[Modules.scala 143:103:@3907.4]
  wire [5:0] _T_58035; // @[Modules.scala 143:103:@3908.4]
  wire [5:0] _T_58040; // @[Modules.scala 143:103:@3912.4]
  wire [4:0] _T_58041; // @[Modules.scala 143:103:@3913.4]
  wire [4:0] _T_58042; // @[Modules.scala 143:103:@3914.4]
  wire [5:0] _T_58047; // @[Modules.scala 143:103:@3918.4]
  wire [4:0] _T_58048; // @[Modules.scala 143:103:@3919.4]
  wire [4:0] _T_58049; // @[Modules.scala 143:103:@3920.4]
  wire [5:0] _T_58053; // @[Modules.scala 144:80:@3923.4]
  wire [5:0] _GEN_101; // @[Modules.scala 143:103:@3924.4]
  wire [6:0] _T_58054; // @[Modules.scala 143:103:@3924.4]
  wire [5:0] _T_58055; // @[Modules.scala 143:103:@3925.4]
  wire [5:0] _T_58056; // @[Modules.scala 143:103:@3926.4]
  wire [5:0] _T_58058; // @[Modules.scala 143:74:@3928.4]
  wire [6:0] _T_58061; // @[Modules.scala 143:103:@3930.4]
  wire [5:0] _T_58062; // @[Modules.scala 143:103:@3931.4]
  wire [5:0] _T_58063; // @[Modules.scala 143:103:@3932.4]
  wire [5:0] _T_58065; // @[Modules.scala 143:74:@3934.4]
  wire [5:0] _T_58067; // @[Modules.scala 144:80:@3935.4]
  wire [6:0] _T_58068; // @[Modules.scala 143:103:@3936.4]
  wire [5:0] _T_58069; // @[Modules.scala 143:103:@3937.4]
  wire [5:0] _T_58070; // @[Modules.scala 143:103:@3938.4]
  wire [5:0] _T_58072; // @[Modules.scala 143:74:@3940.4]
  wire [5:0] _T_58074; // @[Modules.scala 144:80:@3941.4]
  wire [6:0] _T_58075; // @[Modules.scala 143:103:@3942.4]
  wire [5:0] _T_58076; // @[Modules.scala 143:103:@3943.4]
  wire [5:0] _T_58077; // @[Modules.scala 143:103:@3944.4]
  wire [5:0] _T_58079; // @[Modules.scala 143:74:@3946.4]
  wire [5:0] _T_58081; // @[Modules.scala 144:80:@3947.4]
  wire [6:0] _T_58082; // @[Modules.scala 143:103:@3948.4]
  wire [5:0] _T_58083; // @[Modules.scala 143:103:@3949.4]
  wire [5:0] _T_58084; // @[Modules.scala 143:103:@3950.4]
  wire [5:0] _T_58089; // @[Modules.scala 143:103:@3954.4]
  wire [4:0] _T_58090; // @[Modules.scala 143:103:@3955.4]
  wire [4:0] _T_58091; // @[Modules.scala 143:103:@3956.4]
  wire [4:0] _T_58095; // @[Modules.scala 144:80:@3959.4]
  wire [5:0] _T_58096; // @[Modules.scala 143:103:@3960.4]
  wire [4:0] _T_58097; // @[Modules.scala 143:103:@3961.4]
  wire [4:0] _T_58098; // @[Modules.scala 143:103:@3962.4]
  wire [5:0] _T_58100; // @[Modules.scala 143:74:@3964.4]
  wire [5:0] _T_58102; // @[Modules.scala 144:80:@3965.4]
  wire [6:0] _T_58103; // @[Modules.scala 143:103:@3966.4]
  wire [5:0] _T_58104; // @[Modules.scala 143:103:@3967.4]
  wire [5:0] _T_58105; // @[Modules.scala 143:103:@3968.4]
  wire [4:0] _T_58107; // @[Modules.scala 143:74:@3970.4]
  wire [4:0] _T_58109; // @[Modules.scala 144:80:@3971.4]
  wire [5:0] _T_58110; // @[Modules.scala 143:103:@3972.4]
  wire [4:0] _T_58111; // @[Modules.scala 143:103:@3973.4]
  wire [4:0] _T_58112; // @[Modules.scala 143:103:@3974.4]
  wire [5:0] _T_58116; // @[Modules.scala 144:80:@3977.4]
  wire [6:0] _T_58117; // @[Modules.scala 143:103:@3978.4]
  wire [5:0] _T_58118; // @[Modules.scala 143:103:@3979.4]
  wire [5:0] _T_58119; // @[Modules.scala 143:103:@3980.4]
  wire [5:0] _T_58121; // @[Modules.scala 143:74:@3982.4]
  wire [5:0] _GEN_102; // @[Modules.scala 143:103:@3984.4]
  wire [6:0] _T_58124; // @[Modules.scala 143:103:@3984.4]
  wire [5:0] _T_58125; // @[Modules.scala 143:103:@3985.4]
  wire [5:0] _T_58126; // @[Modules.scala 143:103:@3986.4]
  wire [5:0] _T_58131; // @[Modules.scala 143:103:@3990.4]
  wire [4:0] _T_58132; // @[Modules.scala 143:103:@3991.4]
  wire [4:0] _T_58133; // @[Modules.scala 143:103:@3992.4]
  wire [5:0] _T_58138; // @[Modules.scala 143:103:@3996.4]
  wire [4:0] _T_58139; // @[Modules.scala 143:103:@3997.4]
  wire [4:0] _T_58140; // @[Modules.scala 143:103:@3998.4]
  wire [5:0] _T_58142; // @[Modules.scala 143:74:@4000.4]
  wire [6:0] _T_58145; // @[Modules.scala 143:103:@4002.4]
  wire [5:0] _T_58146; // @[Modules.scala 143:103:@4003.4]
  wire [5:0] _T_58147; // @[Modules.scala 143:103:@4004.4]
  wire [5:0] _T_58151; // @[Modules.scala 144:80:@4007.4]
  wire [6:0] _T_58152; // @[Modules.scala 143:103:@4008.4]
  wire [5:0] _T_58153; // @[Modules.scala 143:103:@4009.4]
  wire [5:0] _T_58154; // @[Modules.scala 143:103:@4010.4]
  wire [5:0] _T_58156; // @[Modules.scala 143:74:@4012.4]
  wire [5:0] _T_58158; // @[Modules.scala 144:80:@4013.4]
  wire [6:0] _T_58159; // @[Modules.scala 143:103:@4014.4]
  wire [5:0] _T_58160; // @[Modules.scala 143:103:@4015.4]
  wire [5:0] _T_58161; // @[Modules.scala 143:103:@4016.4]
  wire [5:0] _T_58163; // @[Modules.scala 143:74:@4018.4]
  wire [6:0] _T_58166; // @[Modules.scala 143:103:@4020.4]
  wire [5:0] _T_58167; // @[Modules.scala 143:103:@4021.4]
  wire [5:0] _T_58168; // @[Modules.scala 143:103:@4022.4]
  wire [5:0] _T_58170; // @[Modules.scala 143:74:@4024.4]
  wire [4:0] _T_58172; // @[Modules.scala 144:80:@4025.4]
  wire [5:0] _GEN_103; // @[Modules.scala 143:103:@4026.4]
  wire [6:0] _T_58173; // @[Modules.scala 143:103:@4026.4]
  wire [5:0] _T_58174; // @[Modules.scala 143:103:@4027.4]
  wire [5:0] _T_58175; // @[Modules.scala 143:103:@4028.4]
  wire [5:0] _T_58177; // @[Modules.scala 143:74:@4030.4]
  wire [6:0] _T_58180; // @[Modules.scala 143:103:@4032.4]
  wire [5:0] _T_58181; // @[Modules.scala 143:103:@4033.4]
  wire [5:0] _T_58182; // @[Modules.scala 143:103:@4034.4]
  wire [6:0] _T_58187; // @[Modules.scala 143:103:@4038.4]
  wire [5:0] _T_58188; // @[Modules.scala 143:103:@4039.4]
  wire [5:0] _T_58189; // @[Modules.scala 143:103:@4040.4]
  wire [4:0] _T_58191; // @[Modules.scala 143:74:@4042.4]
  wire [4:0] _T_58193; // @[Modules.scala 144:80:@4043.4]
  wire [5:0] _T_58194; // @[Modules.scala 143:103:@4044.4]
  wire [4:0] _T_58195; // @[Modules.scala 143:103:@4045.4]
  wire [4:0] _T_58196; // @[Modules.scala 143:103:@4046.4]
  wire [5:0] _T_58200; // @[Modules.scala 144:80:@4049.4]
  wire [6:0] _T_58201; // @[Modules.scala 143:103:@4050.4]
  wire [5:0] _T_58202; // @[Modules.scala 143:103:@4051.4]
  wire [5:0] _T_58203; // @[Modules.scala 143:103:@4052.4]
  wire [5:0] _T_58205; // @[Modules.scala 143:74:@4054.4]
  wire [5:0] _T_58207; // @[Modules.scala 144:80:@4055.4]
  wire [6:0] _T_58208; // @[Modules.scala 143:103:@4056.4]
  wire [5:0] _T_58209; // @[Modules.scala 143:103:@4057.4]
  wire [5:0] _T_58210; // @[Modules.scala 143:103:@4058.4]
  wire [5:0] _T_58212; // @[Modules.scala 143:74:@4060.4]
  wire [5:0] _GEN_105; // @[Modules.scala 143:103:@4062.4]
  wire [6:0] _T_58215; // @[Modules.scala 143:103:@4062.4]
  wire [5:0] _T_58216; // @[Modules.scala 143:103:@4063.4]
  wire [5:0] _T_58217; // @[Modules.scala 143:103:@4064.4]
  wire [5:0] _T_58222; // @[Modules.scala 143:103:@4068.4]
  wire [4:0] _T_58223; // @[Modules.scala 143:103:@4069.4]
  wire [4:0] _T_58224; // @[Modules.scala 143:103:@4070.4]
  wire [5:0] _T_58226; // @[Modules.scala 143:74:@4072.4]
  wire [6:0] _T_58229; // @[Modules.scala 143:103:@4074.4]
  wire [5:0] _T_58230; // @[Modules.scala 143:103:@4075.4]
  wire [5:0] _T_58231; // @[Modules.scala 143:103:@4076.4]
  wire [5:0] _T_58233; // @[Modules.scala 143:74:@4078.4]
  wire [5:0] _T_58235; // @[Modules.scala 144:80:@4079.4]
  wire [6:0] _T_58236; // @[Modules.scala 143:103:@4080.4]
  wire [5:0] _T_58237; // @[Modules.scala 143:103:@4081.4]
  wire [5:0] _T_58238; // @[Modules.scala 143:103:@4082.4]
  wire [5:0] _T_58240; // @[Modules.scala 143:74:@4084.4]
  wire [6:0] _T_58243; // @[Modules.scala 143:103:@4086.4]
  wire [5:0] _T_58244; // @[Modules.scala 143:103:@4087.4]
  wire [5:0] _T_58245; // @[Modules.scala 143:103:@4088.4]
  wire [5:0] _T_58247; // @[Modules.scala 143:74:@4090.4]
  wire [5:0] _T_58249; // @[Modules.scala 144:80:@4091.4]
  wire [6:0] _T_58250; // @[Modules.scala 143:103:@4092.4]
  wire [5:0] _T_58251; // @[Modules.scala 143:103:@4093.4]
  wire [5:0] _T_58252; // @[Modules.scala 143:103:@4094.4]
  wire [4:0] _T_58254; // @[Modules.scala 143:74:@4096.4]
  wire [5:0] _T_58257; // @[Modules.scala 143:103:@4098.4]
  wire [4:0] _T_58258; // @[Modules.scala 143:103:@4099.4]
  wire [4:0] _T_58259; // @[Modules.scala 143:103:@4100.4]
  wire [4:0] _T_58261; // @[Modules.scala 143:74:@4102.4]
  wire [4:0] _T_58263; // @[Modules.scala 144:80:@4103.4]
  wire [5:0] _T_58264; // @[Modules.scala 143:103:@4104.4]
  wire [4:0] _T_58265; // @[Modules.scala 143:103:@4105.4]
  wire [4:0] _T_58266; // @[Modules.scala 143:103:@4106.4]
  wire [5:0] _T_58268; // @[Modules.scala 143:74:@4108.4]
  wire [5:0] _T_58270; // @[Modules.scala 144:80:@4109.4]
  wire [6:0] _T_58271; // @[Modules.scala 143:103:@4110.4]
  wire [5:0] _T_58272; // @[Modules.scala 143:103:@4111.4]
  wire [5:0] _T_58273; // @[Modules.scala 143:103:@4112.4]
  wire [4:0] _T_58277; // @[Modules.scala 144:80:@4115.4]
  wire [5:0] _GEN_106; // @[Modules.scala 143:103:@4116.4]
  wire [6:0] _T_58278; // @[Modules.scala 143:103:@4116.4]
  wire [5:0] _T_58279; // @[Modules.scala 143:103:@4117.4]
  wire [5:0] _T_58280; // @[Modules.scala 143:103:@4118.4]
  wire [5:0] _T_58282; // @[Modules.scala 143:74:@4120.4]
  wire [6:0] _T_58285; // @[Modules.scala 143:103:@4122.4]
  wire [5:0] _T_58286; // @[Modules.scala 143:103:@4123.4]
  wire [5:0] _T_58287; // @[Modules.scala 143:103:@4124.4]
  wire [5:0] _T_58289; // @[Modules.scala 143:74:@4126.4]
  wire [5:0] _T_58291; // @[Modules.scala 144:80:@4127.4]
  wire [6:0] _T_58292; // @[Modules.scala 143:103:@4128.4]
  wire [5:0] _T_58293; // @[Modules.scala 143:103:@4129.4]
  wire [5:0] _T_58294; // @[Modules.scala 143:103:@4130.4]
  wire [5:0] _T_58296; // @[Modules.scala 143:74:@4132.4]
  wire [5:0] _GEN_107; // @[Modules.scala 143:103:@4134.4]
  wire [6:0] _T_58299; // @[Modules.scala 143:103:@4134.4]
  wire [5:0] _T_58300; // @[Modules.scala 143:103:@4135.4]
  wire [5:0] _T_58301; // @[Modules.scala 143:103:@4136.4]
  wire [5:0] _T_58306; // @[Modules.scala 143:103:@4140.4]
  wire [4:0] _T_58307; // @[Modules.scala 143:103:@4141.4]
  wire [4:0] _T_58308; // @[Modules.scala 143:103:@4142.4]
  wire [5:0] _T_58310; // @[Modules.scala 143:74:@4144.4]
  wire [6:0] _T_58313; // @[Modules.scala 143:103:@4146.4]
  wire [5:0] _T_58314; // @[Modules.scala 143:103:@4147.4]
  wire [5:0] _T_58315; // @[Modules.scala 143:103:@4148.4]
  wire [4:0] _T_58326; // @[Modules.scala 144:80:@4157.4]
  wire [5:0] _T_58327; // @[Modules.scala 143:103:@4158.4]
  wire [4:0] _T_58328; // @[Modules.scala 143:103:@4159.4]
  wire [4:0] _T_58329; // @[Modules.scala 143:103:@4160.4]
  wire [4:0] _T_58331; // @[Modules.scala 143:74:@4162.4]
  wire [4:0] _T_58333; // @[Modules.scala 144:80:@4163.4]
  wire [5:0] _T_58334; // @[Modules.scala 143:103:@4164.4]
  wire [4:0] _T_58335; // @[Modules.scala 143:103:@4165.4]
  wire [4:0] _T_58336; // @[Modules.scala 143:103:@4166.4]
  wire [4:0] _T_58338; // @[Modules.scala 143:74:@4168.4]
  wire [4:0] _T_58340; // @[Modules.scala 144:80:@4169.4]
  wire [5:0] _T_58341; // @[Modules.scala 143:103:@4170.4]
  wire [4:0] _T_58342; // @[Modules.scala 143:103:@4171.4]
  wire [4:0] _T_58343; // @[Modules.scala 143:103:@4172.4]
  wire [4:0] _T_58347; // @[Modules.scala 144:80:@4175.4]
  wire [5:0] _T_58348; // @[Modules.scala 143:103:@4176.4]
  wire [4:0] _T_58349; // @[Modules.scala 143:103:@4177.4]
  wire [4:0] _T_58350; // @[Modules.scala 143:103:@4178.4]
  wire [4:0] _T_58352; // @[Modules.scala 143:74:@4180.4]
  wire [5:0] _T_58355; // @[Modules.scala 143:103:@4182.4]
  wire [4:0] _T_58356; // @[Modules.scala 143:103:@4183.4]
  wire [4:0] _T_58357; // @[Modules.scala 143:103:@4184.4]
  wire [5:0] _T_58361; // @[Modules.scala 144:80:@4187.4]
  wire [6:0] _T_58362; // @[Modules.scala 143:103:@4188.4]
  wire [5:0] _T_58363; // @[Modules.scala 143:103:@4189.4]
  wire [5:0] _T_58364; // @[Modules.scala 143:103:@4190.4]
  wire [4:0] _T_58375; // @[Modules.scala 144:80:@4199.4]
  wire [5:0] _T_58376; // @[Modules.scala 143:103:@4200.4]
  wire [4:0] _T_58377; // @[Modules.scala 143:103:@4201.4]
  wire [4:0] _T_58378; // @[Modules.scala 143:103:@4202.4]
  wire [4:0] _T_58382; // @[Modules.scala 144:80:@4205.4]
  wire [5:0] _T_58383; // @[Modules.scala 143:103:@4206.4]
  wire [4:0] _T_58384; // @[Modules.scala 143:103:@4207.4]
  wire [4:0] _T_58385; // @[Modules.scala 143:103:@4208.4]
  wire [4:0] _T_58387; // @[Modules.scala 143:74:@4210.4]
  wire [5:0] _GEN_109; // @[Modules.scala 143:103:@4212.4]
  wire [6:0] _T_58390; // @[Modules.scala 143:103:@4212.4]
  wire [5:0] _T_58391; // @[Modules.scala 143:103:@4213.4]
  wire [5:0] _T_58392; // @[Modules.scala 143:103:@4214.4]
  wire [6:0] _T_58397; // @[Modules.scala 143:103:@4218.4]
  wire [5:0] _T_58398; // @[Modules.scala 143:103:@4219.4]
  wire [5:0] _T_58399; // @[Modules.scala 143:103:@4220.4]
  wire [4:0] _T_58401; // @[Modules.scala 143:74:@4222.4]
  wire [5:0] _T_58403; // @[Modules.scala 144:80:@4223.4]
  wire [5:0] _GEN_111; // @[Modules.scala 143:103:@4224.4]
  wire [6:0] _T_58404; // @[Modules.scala 143:103:@4224.4]
  wire [5:0] _T_58405; // @[Modules.scala 143:103:@4225.4]
  wire [5:0] _T_58406; // @[Modules.scala 143:103:@4226.4]
  wire [4:0] _T_58410; // @[Modules.scala 144:80:@4229.4]
  wire [5:0] _T_58411; // @[Modules.scala 143:103:@4230.4]
  wire [4:0] _T_58412; // @[Modules.scala 143:103:@4231.4]
  wire [4:0] _T_58413; // @[Modules.scala 143:103:@4232.4]
  wire [4:0] _T_58415; // @[Modules.scala 143:74:@4234.4]
  wire [4:0] _T_58417; // @[Modules.scala 144:80:@4235.4]
  wire [5:0] _T_58418; // @[Modules.scala 143:103:@4236.4]
  wire [4:0] _T_58419; // @[Modules.scala 143:103:@4237.4]
  wire [4:0] _T_58420; // @[Modules.scala 143:103:@4238.4]
  wire [5:0] _T_58424; // @[Modules.scala 144:80:@4241.4]
  wire [6:0] _T_58425; // @[Modules.scala 143:103:@4242.4]
  wire [5:0] _T_58426; // @[Modules.scala 143:103:@4243.4]
  wire [5:0] _T_58427; // @[Modules.scala 143:103:@4244.4]
  wire [5:0] _GEN_112; // @[Modules.scala 143:103:@4248.4]
  wire [6:0] _T_58432; // @[Modules.scala 143:103:@4248.4]
  wire [5:0] _T_58433; // @[Modules.scala 143:103:@4249.4]
  wire [5:0] _T_58434; // @[Modules.scala 143:103:@4250.4]
  wire [5:0] _T_58438; // @[Modules.scala 144:80:@4253.4]
  wire [6:0] _T_58439; // @[Modules.scala 143:103:@4254.4]
  wire [5:0] _T_58440; // @[Modules.scala 143:103:@4255.4]
  wire [5:0] _T_58441; // @[Modules.scala 143:103:@4256.4]
  wire [4:0] _T_58445; // @[Modules.scala 144:80:@4259.4]
  wire [5:0] _T_58446; // @[Modules.scala 143:103:@4260.4]
  wire [4:0] _T_58447; // @[Modules.scala 143:103:@4261.4]
  wire [4:0] _T_58448; // @[Modules.scala 143:103:@4262.4]
  wire [4:0] _T_58450; // @[Modules.scala 143:74:@4264.4]
  wire [4:0] _T_58452; // @[Modules.scala 144:80:@4265.4]
  wire [5:0] _T_58453; // @[Modules.scala 143:103:@4266.4]
  wire [4:0] _T_58454; // @[Modules.scala 143:103:@4267.4]
  wire [4:0] _T_58455; // @[Modules.scala 143:103:@4268.4]
  wire [4:0] _T_58457; // @[Modules.scala 143:74:@4270.4]
  wire [4:0] _T_58459; // @[Modules.scala 144:80:@4271.4]
  wire [5:0] _T_58460; // @[Modules.scala 143:103:@4272.4]
  wire [4:0] _T_58461; // @[Modules.scala 143:103:@4273.4]
  wire [4:0] _T_58462; // @[Modules.scala 143:103:@4274.4]
  wire [4:0] _T_58464; // @[Modules.scala 143:74:@4276.4]
  wire [4:0] _T_58466; // @[Modules.scala 144:80:@4277.4]
  wire [5:0] _T_58467; // @[Modules.scala 143:103:@4278.4]
  wire [4:0] _T_58468; // @[Modules.scala 143:103:@4279.4]
  wire [4:0] _T_58469; // @[Modules.scala 143:103:@4280.4]
  wire [4:0] _T_58471; // @[Modules.scala 143:74:@4282.4]
  wire [4:0] _T_58473; // @[Modules.scala 144:80:@4283.4]
  wire [5:0] _T_58474; // @[Modules.scala 143:103:@4284.4]
  wire [4:0] _T_58475; // @[Modules.scala 143:103:@4285.4]
  wire [4:0] _T_58476; // @[Modules.scala 143:103:@4286.4]
  wire [5:0] _T_58478; // @[Modules.scala 143:74:@4288.4]
  wire [5:0] _T_58480; // @[Modules.scala 144:80:@4289.4]
  wire [6:0] _T_58481; // @[Modules.scala 143:103:@4290.4]
  wire [5:0] _T_58482; // @[Modules.scala 143:103:@4291.4]
  wire [5:0] _T_58483; // @[Modules.scala 143:103:@4292.4]
  wire [5:0] _T_58485; // @[Modules.scala 143:74:@4294.4]
  wire [6:0] _T_58488; // @[Modules.scala 143:103:@4296.4]
  wire [5:0] _T_58489; // @[Modules.scala 143:103:@4297.4]
  wire [5:0] _T_58490; // @[Modules.scala 143:103:@4298.4]
  wire [4:0] _T_58492; // @[Modules.scala 143:74:@4300.4]
  wire [4:0] _T_58494; // @[Modules.scala 144:80:@4301.4]
  wire [5:0] _T_58495; // @[Modules.scala 143:103:@4302.4]
  wire [4:0] _T_58496; // @[Modules.scala 143:103:@4303.4]
  wire [4:0] _T_58497; // @[Modules.scala 143:103:@4304.4]
  wire [5:0] _T_58501; // @[Modules.scala 144:80:@4307.4]
  wire [6:0] _T_58502; // @[Modules.scala 143:103:@4308.4]
  wire [5:0] _T_58503; // @[Modules.scala 143:103:@4309.4]
  wire [5:0] _T_58504; // @[Modules.scala 143:103:@4310.4]
  wire [4:0] _T_58520; // @[Modules.scala 143:74:@4324.4]
  wire [4:0] _T_58522; // @[Modules.scala 144:80:@4325.4]
  wire [5:0] _T_58523; // @[Modules.scala 143:103:@4326.4]
  wire [4:0] _T_58524; // @[Modules.scala 143:103:@4327.4]
  wire [4:0] _T_58525; // @[Modules.scala 143:103:@4328.4]
  wire [4:0] _T_58527; // @[Modules.scala 143:74:@4330.4]
  wire [4:0] _T_58529; // @[Modules.scala 144:80:@4331.4]
  wire [5:0] _T_58530; // @[Modules.scala 143:103:@4332.4]
  wire [4:0] _T_58531; // @[Modules.scala 143:103:@4333.4]
  wire [4:0] _T_58532; // @[Modules.scala 143:103:@4334.4]
  wire [4:0] _T_58536; // @[Modules.scala 144:80:@4337.4]
  wire [5:0] _T_58537; // @[Modules.scala 143:103:@4338.4]
  wire [4:0] _T_58538; // @[Modules.scala 143:103:@4339.4]
  wire [4:0] _T_58539; // @[Modules.scala 143:103:@4340.4]
  wire [4:0] _T_58541; // @[Modules.scala 143:74:@4342.4]
  wire [4:0] _T_58543; // @[Modules.scala 144:80:@4343.4]
  wire [5:0] _T_58544; // @[Modules.scala 143:103:@4344.4]
  wire [4:0] _T_58545; // @[Modules.scala 143:103:@4345.4]
  wire [4:0] _T_58546; // @[Modules.scala 143:103:@4346.4]
  wire [4:0] _T_58548; // @[Modules.scala 143:74:@4348.4]
  wire [4:0] _T_58550; // @[Modules.scala 144:80:@4349.4]
  wire [5:0] _T_58551; // @[Modules.scala 143:103:@4350.4]
  wire [4:0] _T_58552; // @[Modules.scala 143:103:@4351.4]
  wire [4:0] _T_58553; // @[Modules.scala 143:103:@4352.4]
  wire [5:0] _T_58557; // @[Modules.scala 144:80:@4355.4]
  wire [5:0] _GEN_115; // @[Modules.scala 143:103:@4356.4]
  wire [6:0] _T_58558; // @[Modules.scala 143:103:@4356.4]
  wire [5:0] _T_58559; // @[Modules.scala 143:103:@4357.4]
  wire [5:0] _T_58560; // @[Modules.scala 143:103:@4358.4]
  wire [4:0] _T_58562; // @[Modules.scala 143:74:@4360.4]
  wire [4:0] _T_58564; // @[Modules.scala 144:80:@4361.4]
  wire [5:0] _T_58565; // @[Modules.scala 143:103:@4362.4]
  wire [4:0] _T_58566; // @[Modules.scala 143:103:@4363.4]
  wire [4:0] _T_58567; // @[Modules.scala 143:103:@4364.4]
  wire [5:0] _T_58569; // @[Modules.scala 143:74:@4366.4]
  wire [4:0] _T_58571; // @[Modules.scala 144:80:@4367.4]
  wire [5:0] _GEN_116; // @[Modules.scala 143:103:@4368.4]
  wire [6:0] _T_58572; // @[Modules.scala 143:103:@4368.4]
  wire [5:0] _T_58573; // @[Modules.scala 143:103:@4369.4]
  wire [5:0] _T_58574; // @[Modules.scala 143:103:@4370.4]
  wire [4:0] _T_58576; // @[Modules.scala 143:74:@4372.4]
  wire [4:0] _T_58578; // @[Modules.scala 144:80:@4373.4]
  wire [5:0] _T_58579; // @[Modules.scala 143:103:@4374.4]
  wire [4:0] _T_58580; // @[Modules.scala 143:103:@4375.4]
  wire [4:0] _T_58581; // @[Modules.scala 143:103:@4376.4]
  wire [6:0] _T_58586; // @[Modules.scala 143:103:@4380.4]
  wire [5:0] _T_58587; // @[Modules.scala 143:103:@4381.4]
  wire [5:0] _T_58588; // @[Modules.scala 143:103:@4382.4]
  wire [5:0] _T_58590; // @[Modules.scala 143:74:@4384.4]
  wire [6:0] _T_58593; // @[Modules.scala 143:103:@4386.4]
  wire [5:0] _T_58594; // @[Modules.scala 143:103:@4387.4]
  wire [5:0] _T_58595; // @[Modules.scala 143:103:@4388.4]
  wire [4:0] _T_58599; // @[Modules.scala 144:80:@4391.4]
  wire [5:0] _GEN_117; // @[Modules.scala 143:103:@4392.4]
  wire [6:0] _T_58600; // @[Modules.scala 143:103:@4392.4]
  wire [5:0] _T_58601; // @[Modules.scala 143:103:@4393.4]
  wire [5:0] _T_58602; // @[Modules.scala 143:103:@4394.4]
  wire [4:0] _T_58606; // @[Modules.scala 144:80:@4397.4]
  wire [5:0] _T_58607; // @[Modules.scala 143:103:@4398.4]
  wire [4:0] _T_58608; // @[Modules.scala 143:103:@4399.4]
  wire [4:0] _T_58609; // @[Modules.scala 143:103:@4400.4]
  wire [4:0] _T_58613; // @[Modules.scala 144:80:@4403.4]
  wire [5:0] _T_58614; // @[Modules.scala 143:103:@4404.4]
  wire [4:0] _T_58615; // @[Modules.scala 143:103:@4405.4]
  wire [4:0] _T_58616; // @[Modules.scala 143:103:@4406.4]
  wire [4:0] _T_58618; // @[Modules.scala 143:74:@4408.4]
  wire [4:0] _T_58620; // @[Modules.scala 144:80:@4409.4]
  wire [5:0] _T_58621; // @[Modules.scala 143:103:@4410.4]
  wire [4:0] _T_58622; // @[Modules.scala 143:103:@4411.4]
  wire [4:0] _T_58623; // @[Modules.scala 143:103:@4412.4]
  wire [4:0] _T_58625; // @[Modules.scala 143:74:@4414.4]
  wire [4:0] _T_58627; // @[Modules.scala 144:80:@4415.4]
  wire [5:0] _T_58628; // @[Modules.scala 143:103:@4416.4]
  wire [4:0] _T_58629; // @[Modules.scala 143:103:@4417.4]
  wire [4:0] _T_58630; // @[Modules.scala 143:103:@4418.4]
  wire [5:0] _T_58632; // @[Modules.scala 143:74:@4420.4]
  wire [6:0] _T_58635; // @[Modules.scala 143:103:@4422.4]
  wire [5:0] _T_58636; // @[Modules.scala 143:103:@4423.4]
  wire [5:0] _T_58637; // @[Modules.scala 143:103:@4424.4]
  wire [4:0] _T_58639; // @[Modules.scala 143:74:@4426.4]
  wire [4:0] _T_58641; // @[Modules.scala 144:80:@4427.4]
  wire [5:0] _T_58642; // @[Modules.scala 143:103:@4428.4]
  wire [4:0] _T_58643; // @[Modules.scala 143:103:@4429.4]
  wire [4:0] _T_58644; // @[Modules.scala 143:103:@4430.4]
  wire [4:0] _T_58646; // @[Modules.scala 143:74:@4432.4]
  wire [4:0] _T_58648; // @[Modules.scala 144:80:@4433.4]
  wire [5:0] _T_58649; // @[Modules.scala 143:103:@4434.4]
  wire [4:0] _T_58650; // @[Modules.scala 143:103:@4435.4]
  wire [4:0] _T_58651; // @[Modules.scala 143:103:@4436.4]
  wire [5:0] _T_58655; // @[Modules.scala 144:80:@4439.4]
  wire [6:0] _T_58656; // @[Modules.scala 143:103:@4440.4]
  wire [5:0] _T_58657; // @[Modules.scala 143:103:@4441.4]
  wire [5:0] _T_58658; // @[Modules.scala 143:103:@4442.4]
  wire [4:0] _T_58660; // @[Modules.scala 143:74:@4444.4]
  wire [5:0] _GEN_119; // @[Modules.scala 143:103:@4446.4]
  wire [6:0] _T_58663; // @[Modules.scala 143:103:@4446.4]
  wire [5:0] _T_58664; // @[Modules.scala 143:103:@4447.4]
  wire [5:0] _T_58665; // @[Modules.scala 143:103:@4448.4]
  wire [6:0] _T_58670; // @[Modules.scala 143:103:@4452.4]
  wire [5:0] _T_58671; // @[Modules.scala 143:103:@4453.4]
  wire [5:0] _T_58672; // @[Modules.scala 143:103:@4454.4]
  wire [4:0] _T_58674; // @[Modules.scala 143:74:@4456.4]
  wire [4:0] _T_58676; // @[Modules.scala 144:80:@4457.4]
  wire [5:0] _T_58677; // @[Modules.scala 143:103:@4458.4]
  wire [4:0] _T_58678; // @[Modules.scala 143:103:@4459.4]
  wire [4:0] _T_58679; // @[Modules.scala 143:103:@4460.4]
  wire [4:0] _T_58681; // @[Modules.scala 143:74:@4462.4]
  wire [4:0] _T_58683; // @[Modules.scala 144:80:@4463.4]
  wire [5:0] _T_58684; // @[Modules.scala 143:103:@4464.4]
  wire [4:0] _T_58685; // @[Modules.scala 143:103:@4465.4]
  wire [4:0] _T_58686; // @[Modules.scala 143:103:@4466.4]
  wire [4:0] _T_58688; // @[Modules.scala 143:74:@4468.4]
  wire [4:0] _T_58690; // @[Modules.scala 144:80:@4469.4]
  wire [5:0] _T_58691; // @[Modules.scala 143:103:@4470.4]
  wire [4:0] _T_58692; // @[Modules.scala 143:103:@4471.4]
  wire [4:0] _T_58693; // @[Modules.scala 143:103:@4472.4]
  wire [4:0] _T_58695; // @[Modules.scala 143:74:@4474.4]
  wire [4:0] _T_58697; // @[Modules.scala 144:80:@4475.4]
  wire [5:0] _T_58698; // @[Modules.scala 143:103:@4476.4]
  wire [4:0] _T_58699; // @[Modules.scala 143:103:@4477.4]
  wire [4:0] _T_58700; // @[Modules.scala 143:103:@4478.4]
  wire [4:0] _T_58704; // @[Modules.scala 144:80:@4481.4]
  wire [5:0] _GEN_120; // @[Modules.scala 143:103:@4482.4]
  wire [6:0] _T_58705; // @[Modules.scala 143:103:@4482.4]
  wire [5:0] _T_58706; // @[Modules.scala 143:103:@4483.4]
  wire [5:0] _T_58707; // @[Modules.scala 143:103:@4484.4]
  wire [4:0] _T_58709; // @[Modules.scala 143:74:@4486.4]
  wire [4:0] _T_58711; // @[Modules.scala 144:80:@4487.4]
  wire [5:0] _T_58712; // @[Modules.scala 143:103:@4488.4]
  wire [4:0] _T_58713; // @[Modules.scala 143:103:@4489.4]
  wire [4:0] _T_58714; // @[Modules.scala 143:103:@4490.4]
  wire [4:0] _T_58718; // @[Modules.scala 144:80:@4493.4]
  wire [5:0] _GEN_121; // @[Modules.scala 143:103:@4494.4]
  wire [6:0] _T_58719; // @[Modules.scala 143:103:@4494.4]
  wire [5:0] _T_58720; // @[Modules.scala 143:103:@4495.4]
  wire [5:0] _T_58721; // @[Modules.scala 143:103:@4496.4]
  wire [4:0] _T_58723; // @[Modules.scala 143:74:@4498.4]
  wire [4:0] _T_58725; // @[Modules.scala 144:80:@4499.4]
  wire [5:0] _T_58726; // @[Modules.scala 143:103:@4500.4]
  wire [4:0] _T_58727; // @[Modules.scala 143:103:@4501.4]
  wire [4:0] _T_58728; // @[Modules.scala 143:103:@4502.4]
  wire [4:0] _T_58730; // @[Modules.scala 143:74:@4504.4]
  wire [4:0] _T_58732; // @[Modules.scala 144:80:@4505.4]
  wire [5:0] _T_58733; // @[Modules.scala 143:103:@4506.4]
  wire [4:0] _T_58734; // @[Modules.scala 143:103:@4507.4]
  wire [4:0] _T_58735; // @[Modules.scala 143:103:@4508.4]
  wire [4:0] _T_58737; // @[Modules.scala 143:74:@4510.4]
  wire [5:0] _T_58740; // @[Modules.scala 143:103:@4512.4]
  wire [4:0] _T_58741; // @[Modules.scala 143:103:@4513.4]
  wire [4:0] _T_58742; // @[Modules.scala 143:103:@4514.4]
  wire [6:0] _T_58747; // @[Modules.scala 143:103:@4518.4]
  wire [5:0] _T_58748; // @[Modules.scala 143:103:@4519.4]
  wire [5:0] _T_58749; // @[Modules.scala 143:103:@4520.4]
  wire [4:0] _T_58753; // @[Modules.scala 144:80:@4523.4]
  wire [5:0] _GEN_122; // @[Modules.scala 143:103:@4524.4]
  wire [6:0] _T_58754; // @[Modules.scala 143:103:@4524.4]
  wire [5:0] _T_58755; // @[Modules.scala 143:103:@4525.4]
  wire [5:0] _T_58756; // @[Modules.scala 143:103:@4526.4]
  wire [4:0] _T_58758; // @[Modules.scala 143:74:@4528.4]
  wire [4:0] _T_58760; // @[Modules.scala 144:80:@4529.4]
  wire [5:0] _T_58761; // @[Modules.scala 143:103:@4530.4]
  wire [4:0] _T_58762; // @[Modules.scala 143:103:@4531.4]
  wire [4:0] _T_58763; // @[Modules.scala 143:103:@4532.4]
  wire [4:0] _T_58765; // @[Modules.scala 143:74:@4534.4]
  wire [4:0] _T_58767; // @[Modules.scala 144:80:@4535.4]
  wire [5:0] _T_58768; // @[Modules.scala 143:103:@4536.4]
  wire [4:0] _T_58769; // @[Modules.scala 143:103:@4537.4]
  wire [4:0] _T_58770; // @[Modules.scala 143:103:@4538.4]
  wire [4:0] _T_58774; // @[Modules.scala 144:80:@4541.4]
  wire [5:0] _GEN_123; // @[Modules.scala 143:103:@4542.4]
  wire [6:0] _T_58775; // @[Modules.scala 143:103:@4542.4]
  wire [5:0] _T_58776; // @[Modules.scala 143:103:@4543.4]
  wire [5:0] _T_58777; // @[Modules.scala 143:103:@4544.4]
  wire [4:0] _T_58779; // @[Modules.scala 143:74:@4546.4]
  wire [4:0] _T_58781; // @[Modules.scala 144:80:@4547.4]
  wire [5:0] _T_58782; // @[Modules.scala 143:103:@4548.4]
  wire [4:0] _T_58783; // @[Modules.scala 143:103:@4549.4]
  wire [4:0] _T_58784; // @[Modules.scala 143:103:@4550.4]
  wire [5:0] _T_58786; // @[Modules.scala 143:74:@4552.4]
  wire [5:0] _T_58788; // @[Modules.scala 144:80:@4553.4]
  wire [6:0] _T_58789; // @[Modules.scala 143:103:@4554.4]
  wire [5:0] _T_58790; // @[Modules.scala 143:103:@4555.4]
  wire [5:0] _T_58791; // @[Modules.scala 143:103:@4556.4]
  wire [4:0] _T_58793; // @[Modules.scala 143:74:@4558.4]
  wire [5:0] _T_58796; // @[Modules.scala 143:103:@4560.4]
  wire [4:0] _T_58797; // @[Modules.scala 143:103:@4561.4]
  wire [4:0] _T_58798; // @[Modules.scala 143:103:@4562.4]
  wire [4:0] _T_58800; // @[Modules.scala 143:74:@4564.4]
  wire [4:0] _T_58802; // @[Modules.scala 144:80:@4565.4]
  wire [5:0] _T_58803; // @[Modules.scala 143:103:@4566.4]
  wire [4:0] _T_58804; // @[Modules.scala 143:103:@4567.4]
  wire [4:0] _T_58805; // @[Modules.scala 143:103:@4568.4]
  wire [4:0] _T_58807; // @[Modules.scala 143:74:@4570.4]
  wire [5:0] _T_58809; // @[Modules.scala 144:80:@4571.4]
  wire [5:0] _GEN_124; // @[Modules.scala 143:103:@4572.4]
  wire [6:0] _T_58810; // @[Modules.scala 143:103:@4572.4]
  wire [5:0] _T_58811; // @[Modules.scala 143:103:@4573.4]
  wire [5:0] _T_58812; // @[Modules.scala 143:103:@4574.4]
  wire [4:0] _T_58814; // @[Modules.scala 143:74:@4576.4]
  wire [4:0] _T_58816; // @[Modules.scala 144:80:@4577.4]
  wire [5:0] _T_58817; // @[Modules.scala 143:103:@4578.4]
  wire [4:0] _T_58818; // @[Modules.scala 143:103:@4579.4]
  wire [4:0] _T_58819; // @[Modules.scala 143:103:@4580.4]
  wire [4:0] _T_58837; // @[Modules.scala 144:80:@4595.4]
  wire [5:0] _GEN_125; // @[Modules.scala 143:103:@4596.4]
  wire [6:0] _T_58838; // @[Modules.scala 143:103:@4596.4]
  wire [5:0] _T_58839; // @[Modules.scala 143:103:@4597.4]
  wire [5:0] _T_58840; // @[Modules.scala 143:103:@4598.4]
  wire [4:0] _T_58844; // @[Modules.scala 144:80:@4601.4]
  wire [5:0] _GEN_126; // @[Modules.scala 143:103:@4602.4]
  wire [6:0] _T_58845; // @[Modules.scala 143:103:@4602.4]
  wire [5:0] _T_58846; // @[Modules.scala 143:103:@4603.4]
  wire [5:0] _T_58847; // @[Modules.scala 143:103:@4604.4]
  wire [4:0] _T_58849; // @[Modules.scala 143:74:@4606.4]
  wire [4:0] _T_58851; // @[Modules.scala 144:80:@4607.4]
  wire [5:0] _T_58852; // @[Modules.scala 143:103:@4608.4]
  wire [4:0] _T_58853; // @[Modules.scala 143:103:@4609.4]
  wire [4:0] _T_58854; // @[Modules.scala 143:103:@4610.4]
  wire [4:0] _T_58856; // @[Modules.scala 143:74:@4612.4]
  wire [5:0] _T_58858; // @[Modules.scala 144:80:@4613.4]
  wire [5:0] _GEN_127; // @[Modules.scala 143:103:@4614.4]
  wire [6:0] _T_58859; // @[Modules.scala 143:103:@4614.4]
  wire [5:0] _T_58860; // @[Modules.scala 143:103:@4615.4]
  wire [5:0] _T_58861; // @[Modules.scala 143:103:@4616.4]
  wire [4:0] _T_58865; // @[Modules.scala 144:80:@4619.4]
  wire [5:0] _T_58866; // @[Modules.scala 143:103:@4620.4]
  wire [4:0] _T_58867; // @[Modules.scala 143:103:@4621.4]
  wire [4:0] _T_58868; // @[Modules.scala 143:103:@4622.4]
  wire [4:0] _T_58870; // @[Modules.scala 143:74:@4624.4]
  wire [4:0] _T_58872; // @[Modules.scala 144:80:@4625.4]
  wire [5:0] _T_58873; // @[Modules.scala 143:103:@4626.4]
  wire [4:0] _T_58874; // @[Modules.scala 143:103:@4627.4]
  wire [4:0] _T_58875; // @[Modules.scala 143:103:@4628.4]
  wire [4:0] _T_58877; // @[Modules.scala 143:74:@4630.4]
  wire [4:0] _T_58879; // @[Modules.scala 144:80:@4631.4]
  wire [5:0] _T_58880; // @[Modules.scala 143:103:@4632.4]
  wire [4:0] _T_58881; // @[Modules.scala 143:103:@4633.4]
  wire [4:0] _T_58882; // @[Modules.scala 143:103:@4634.4]
  wire [4:0] _T_58886; // @[Modules.scala 144:80:@4637.4]
  wire [5:0] _GEN_128; // @[Modules.scala 143:103:@4638.4]
  wire [6:0] _T_58887; // @[Modules.scala 143:103:@4638.4]
  wire [5:0] _T_58888; // @[Modules.scala 143:103:@4639.4]
  wire [5:0] _T_58889; // @[Modules.scala 143:103:@4640.4]
  wire [4:0] _T_58891; // @[Modules.scala 143:74:@4642.4]
  wire [5:0] _GEN_129; // @[Modules.scala 143:103:@4644.4]
  wire [6:0] _T_58894; // @[Modules.scala 143:103:@4644.4]
  wire [5:0] _T_58895; // @[Modules.scala 143:103:@4645.4]
  wire [5:0] _T_58896; // @[Modules.scala 143:103:@4646.4]
  wire [5:0] _T_58912; // @[Modules.scala 143:74:@4660.4]
  wire [6:0] _T_58915; // @[Modules.scala 143:103:@4662.4]
  wire [5:0] _T_58916; // @[Modules.scala 143:103:@4663.4]
  wire [5:0] _T_58917; // @[Modules.scala 143:103:@4664.4]
  wire [5:0] _T_58919; // @[Modules.scala 143:74:@4666.4]
  wire [5:0] _GEN_130; // @[Modules.scala 143:103:@4668.4]
  wire [6:0] _T_58922; // @[Modules.scala 143:103:@4668.4]
  wire [5:0] _T_58923; // @[Modules.scala 143:103:@4669.4]
  wire [5:0] _T_58924; // @[Modules.scala 143:103:@4670.4]
  wire [5:0] _T_58929; // @[Modules.scala 143:103:@4674.4]
  wire [4:0] _T_58930; // @[Modules.scala 143:103:@4675.4]
  wire [4:0] _T_58931; // @[Modules.scala 143:103:@4676.4]
  wire [5:0] _T_58933; // @[Modules.scala 143:74:@4678.4]
  wire [5:0] _GEN_131; // @[Modules.scala 143:103:@4680.4]
  wire [6:0] _T_58936; // @[Modules.scala 143:103:@4680.4]
  wire [5:0] _T_58937; // @[Modules.scala 143:103:@4681.4]
  wire [5:0] _T_58938; // @[Modules.scala 143:103:@4682.4]
  wire [4:0] _T_58940; // @[Modules.scala 143:74:@4684.4]
  wire [4:0] _T_58942; // @[Modules.scala 144:80:@4685.4]
  wire [5:0] _T_58943; // @[Modules.scala 143:103:@4686.4]
  wire [4:0] _T_58944; // @[Modules.scala 143:103:@4687.4]
  wire [4:0] _T_58945; // @[Modules.scala 143:103:@4688.4]
  wire [4:0] _T_58947; // @[Modules.scala 143:74:@4690.4]
  wire [4:0] _T_58949; // @[Modules.scala 144:80:@4691.4]
  wire [5:0] _T_58950; // @[Modules.scala 143:103:@4692.4]
  wire [4:0] _T_58951; // @[Modules.scala 143:103:@4693.4]
  wire [4:0] _T_58952; // @[Modules.scala 143:103:@4694.4]
  wire [4:0] _T_58954; // @[Modules.scala 143:74:@4696.4]
  wire [5:0] _GEN_132; // @[Modules.scala 143:103:@4698.4]
  wire [6:0] _T_58957; // @[Modules.scala 143:103:@4698.4]
  wire [5:0] _T_58958; // @[Modules.scala 143:103:@4699.4]
  wire [5:0] _T_58959; // @[Modules.scala 143:103:@4700.4]
  wire [6:0] _T_58964; // @[Modules.scala 143:103:@4704.4]
  wire [5:0] _T_58965; // @[Modules.scala 143:103:@4705.4]
  wire [5:0] _T_58966; // @[Modules.scala 143:103:@4706.4]
  wire [5:0] _T_58982; // @[Modules.scala 143:74:@4720.4]
  wire [5:0] _T_58984; // @[Modules.scala 144:80:@4721.4]
  wire [6:0] _T_58985; // @[Modules.scala 143:103:@4722.4]
  wire [5:0] _T_58986; // @[Modules.scala 143:103:@4723.4]
  wire [5:0] _T_58987; // @[Modules.scala 143:103:@4724.4]
  wire [5:0] _T_58992; // @[Modules.scala 143:103:@4728.4]
  wire [4:0] _T_58993; // @[Modules.scala 143:103:@4729.4]
  wire [4:0] _T_58994; // @[Modules.scala 143:103:@4730.4]
  wire [5:0] _T_58999; // @[Modules.scala 143:103:@4734.4]
  wire [4:0] _T_59000; // @[Modules.scala 143:103:@4735.4]
  wire [4:0] _T_59001; // @[Modules.scala 143:103:@4736.4]
  wire [5:0] _T_59003; // @[Modules.scala 143:74:@4738.4]
  wire [5:0] _T_59005; // @[Modules.scala 144:80:@4739.4]
  wire [6:0] _T_59006; // @[Modules.scala 143:103:@4740.4]
  wire [5:0] _T_59007; // @[Modules.scala 143:103:@4741.4]
  wire [5:0] _T_59008; // @[Modules.scala 143:103:@4742.4]
  wire [4:0] _T_59017; // @[Modules.scala 143:74:@4750.4]
  wire [4:0] _T_59019; // @[Modules.scala 144:80:@4751.4]
  wire [5:0] _T_59020; // @[Modules.scala 143:103:@4752.4]
  wire [4:0] _T_59021; // @[Modules.scala 143:103:@4753.4]
  wire [4:0] _T_59022; // @[Modules.scala 143:103:@4754.4]
  wire [4:0] _T_59024; // @[Modules.scala 143:74:@4756.4]
  wire [5:0] _GEN_133; // @[Modules.scala 143:103:@4758.4]
  wire [6:0] _T_59027; // @[Modules.scala 143:103:@4758.4]
  wire [5:0] _T_59028; // @[Modules.scala 143:103:@4759.4]
  wire [5:0] _T_59029; // @[Modules.scala 143:103:@4760.4]
  wire [5:0] _T_59033; // @[Modules.scala 144:80:@4763.4]
  wire [6:0] _T_59034; // @[Modules.scala 143:103:@4764.4]
  wire [5:0] _T_59035; // @[Modules.scala 143:103:@4765.4]
  wire [5:0] _T_59036; // @[Modules.scala 143:103:@4766.4]
  wire [5:0] _T_59054; // @[Modules.scala 144:80:@4781.4]
  wire [6:0] _T_59055; // @[Modules.scala 143:103:@4782.4]
  wire [5:0] _T_59056; // @[Modules.scala 143:103:@4783.4]
  wire [5:0] _T_59057; // @[Modules.scala 143:103:@4784.4]
  wire [5:0] _T_59059; // @[Modules.scala 143:74:@4786.4]
  wire [5:0] _T_59061; // @[Modules.scala 144:80:@4787.4]
  wire [6:0] _T_59062; // @[Modules.scala 143:103:@4788.4]
  wire [5:0] _T_59063; // @[Modules.scala 143:103:@4789.4]
  wire [5:0] _T_59064; // @[Modules.scala 143:103:@4790.4]
  wire [4:0] _T_59066; // @[Modules.scala 143:74:@4792.4]
  wire [5:0] _T_59069; // @[Modules.scala 143:103:@4794.4]
  wire [4:0] _T_59070; // @[Modules.scala 143:103:@4795.4]
  wire [4:0] _T_59071; // @[Modules.scala 143:103:@4796.4]
  wire [5:0] _T_59075; // @[Modules.scala 144:80:@4799.4]
  wire [5:0] _GEN_134; // @[Modules.scala 143:103:@4800.4]
  wire [6:0] _T_59076; // @[Modules.scala 143:103:@4800.4]
  wire [5:0] _T_59077; // @[Modules.scala 143:103:@4801.4]
  wire [5:0] _T_59078; // @[Modules.scala 143:103:@4802.4]
  wire [5:0] _T_59080; // @[Modules.scala 143:74:@4804.4]
  wire [5:0] _T_59082; // @[Modules.scala 144:80:@4805.4]
  wire [6:0] _T_59083; // @[Modules.scala 143:103:@4806.4]
  wire [5:0] _T_59084; // @[Modules.scala 143:103:@4807.4]
  wire [5:0] _T_59085; // @[Modules.scala 143:103:@4808.4]
  wire [5:0] _T_59087; // @[Modules.scala 143:74:@4810.4]
  wire [5:0] _T_59089; // @[Modules.scala 144:80:@4811.4]
  wire [6:0] _T_59090; // @[Modules.scala 143:103:@4812.4]
  wire [5:0] _T_59091; // @[Modules.scala 143:103:@4813.4]
  wire [5:0] _T_59092; // @[Modules.scala 143:103:@4814.4]
  wire [5:0] _T_59094; // @[Modules.scala 143:74:@4816.4]
  wire [5:0] _GEN_135; // @[Modules.scala 143:103:@4818.4]
  wire [6:0] _T_59097; // @[Modules.scala 143:103:@4818.4]
  wire [5:0] _T_59098; // @[Modules.scala 143:103:@4819.4]
  wire [5:0] _T_59099; // @[Modules.scala 143:103:@4820.4]
  wire [5:0] _T_59104; // @[Modules.scala 143:103:@4824.4]
  wire [4:0] _T_59105; // @[Modules.scala 143:103:@4825.4]
  wire [4:0] _T_59106; // @[Modules.scala 143:103:@4826.4]
  wire [4:0] _T_59108; // @[Modules.scala 143:74:@4828.4]
  wire [5:0] _GEN_136; // @[Modules.scala 143:103:@4830.4]
  wire [6:0] _T_59111; // @[Modules.scala 143:103:@4830.4]
  wire [5:0] _T_59112; // @[Modules.scala 143:103:@4831.4]
  wire [5:0] _T_59113; // @[Modules.scala 143:103:@4832.4]
  wire [4:0] _T_59115; // @[Modules.scala 143:74:@4834.4]
  wire [5:0] _GEN_137; // @[Modules.scala 143:103:@4836.4]
  wire [6:0] _T_59118; // @[Modules.scala 143:103:@4836.4]
  wire [5:0] _T_59119; // @[Modules.scala 143:103:@4837.4]
  wire [5:0] _T_59120; // @[Modules.scala 143:103:@4838.4]
  wire [4:0] _T_59122; // @[Modules.scala 143:74:@4840.4]
  wire [5:0] _T_59124; // @[Modules.scala 144:80:@4841.4]
  wire [5:0] _GEN_138; // @[Modules.scala 143:103:@4842.4]
  wire [6:0] _T_59125; // @[Modules.scala 143:103:@4842.4]
  wire [5:0] _T_59126; // @[Modules.scala 143:103:@4843.4]
  wire [5:0] _T_59127; // @[Modules.scala 143:103:@4844.4]
  wire [5:0] _T_59129; // @[Modules.scala 143:74:@4846.4]
  wire [5:0] _T_59131; // @[Modules.scala 144:80:@4847.4]
  wire [6:0] _T_59132; // @[Modules.scala 143:103:@4848.4]
  wire [5:0] _T_59133; // @[Modules.scala 143:103:@4849.4]
  wire [5:0] _T_59134; // @[Modules.scala 143:103:@4850.4]
  wire [6:0] _T_59139; // @[Modules.scala 143:103:@4854.4]
  wire [5:0] _T_59140; // @[Modules.scala 143:103:@4855.4]
  wire [5:0] _T_59141; // @[Modules.scala 143:103:@4856.4]
  wire [6:0] _T_59146; // @[Modules.scala 143:103:@4860.4]
  wire [5:0] _T_59147; // @[Modules.scala 143:103:@4861.4]
  wire [5:0] _T_59148; // @[Modules.scala 143:103:@4862.4]
  wire [5:0] _T_59152; // @[Modules.scala 144:80:@4865.4]
  wire [6:0] _T_59153; // @[Modules.scala 143:103:@4866.4]
  wire [5:0] _T_59154; // @[Modules.scala 143:103:@4867.4]
  wire [5:0] _T_59155; // @[Modules.scala 143:103:@4868.4]
  wire [5:0] _T_59157; // @[Modules.scala 143:74:@4870.4]
  wire [5:0] _T_59159; // @[Modules.scala 144:80:@4871.4]
  wire [6:0] _T_59160; // @[Modules.scala 143:103:@4872.4]
  wire [5:0] _T_59161; // @[Modules.scala 143:103:@4873.4]
  wire [5:0] _T_59162; // @[Modules.scala 143:103:@4874.4]
  wire [5:0] _T_59164; // @[Modules.scala 143:74:@4876.4]
  wire [5:0] _T_59166; // @[Modules.scala 144:80:@4877.4]
  wire [6:0] _T_59167; // @[Modules.scala 143:103:@4878.4]
  wire [5:0] _T_59168; // @[Modules.scala 143:103:@4879.4]
  wire [5:0] _T_59169; // @[Modules.scala 143:103:@4880.4]
  wire [5:0] _T_59171; // @[Modules.scala 143:74:@4882.4]
  wire [5:0] _T_59173; // @[Modules.scala 144:80:@4883.4]
  wire [6:0] _T_59174; // @[Modules.scala 143:103:@4884.4]
  wire [5:0] _T_59175; // @[Modules.scala 143:103:@4885.4]
  wire [5:0] _T_59176; // @[Modules.scala 143:103:@4886.4]
  wire [5:0] _T_59178; // @[Modules.scala 143:74:@4888.4]
  wire [5:0] _T_59180; // @[Modules.scala 144:80:@4889.4]
  wire [6:0] _T_59181; // @[Modules.scala 143:103:@4890.4]
  wire [5:0] _T_59182; // @[Modules.scala 143:103:@4891.4]
  wire [5:0] _T_59183; // @[Modules.scala 143:103:@4892.4]
  wire [5:0] _T_59185; // @[Modules.scala 143:74:@4894.4]
  wire [5:0] _GEN_139; // @[Modules.scala 143:103:@4896.4]
  wire [6:0] _T_59188; // @[Modules.scala 143:103:@4896.4]
  wire [5:0] _T_59189; // @[Modules.scala 143:103:@4897.4]
  wire [5:0] _T_59190; // @[Modules.scala 143:103:@4898.4]
  wire [4:0] _T_59194; // @[Modules.scala 144:80:@4901.4]
  wire [5:0] _T_59195; // @[Modules.scala 143:103:@4902.4]
  wire [4:0] _T_59196; // @[Modules.scala 143:103:@4903.4]
  wire [4:0] _T_59197; // @[Modules.scala 143:103:@4904.4]
  wire [4:0] _T_59199; // @[Modules.scala 143:74:@4906.4]
  wire [5:0] _T_59201; // @[Modules.scala 144:80:@4907.4]
  wire [5:0] _GEN_140; // @[Modules.scala 143:103:@4908.4]
  wire [6:0] _T_59202; // @[Modules.scala 143:103:@4908.4]
  wire [5:0] _T_59203; // @[Modules.scala 143:103:@4909.4]
  wire [5:0] _T_59204; // @[Modules.scala 143:103:@4910.4]
  wire [5:0] _T_59206; // @[Modules.scala 143:74:@4912.4]
  wire [6:0] _T_59209; // @[Modules.scala 143:103:@4914.4]
  wire [5:0] _T_59210; // @[Modules.scala 143:103:@4915.4]
  wire [5:0] _T_59211; // @[Modules.scala 143:103:@4916.4]
  wire [5:0] _T_59227; // @[Modules.scala 143:74:@4930.4]
  wire [5:0] _T_59229; // @[Modules.scala 144:80:@4931.4]
  wire [6:0] _T_59230; // @[Modules.scala 143:103:@4932.4]
  wire [5:0] _T_59231; // @[Modules.scala 143:103:@4933.4]
  wire [5:0] _T_59232; // @[Modules.scala 143:103:@4934.4]
  wire [5:0] _T_59234; // @[Modules.scala 143:74:@4936.4]
  wire [6:0] _T_59237; // @[Modules.scala 143:103:@4938.4]
  wire [5:0] _T_59238; // @[Modules.scala 143:103:@4939.4]
  wire [5:0] _T_59239; // @[Modules.scala 143:103:@4940.4]
  wire [5:0] _T_59243; // @[Modules.scala 144:80:@4943.4]
  wire [6:0] _T_59244; // @[Modules.scala 143:103:@4944.4]
  wire [5:0] _T_59245; // @[Modules.scala 143:103:@4945.4]
  wire [5:0] _T_59246; // @[Modules.scala 143:103:@4946.4]
  wire [5:0] _T_59248; // @[Modules.scala 143:74:@4948.4]
  wire [5:0] _T_59250; // @[Modules.scala 144:80:@4949.4]
  wire [6:0] _T_59251; // @[Modules.scala 143:103:@4950.4]
  wire [5:0] _T_59252; // @[Modules.scala 143:103:@4951.4]
  wire [5:0] _T_59253; // @[Modules.scala 143:103:@4952.4]
  wire [5:0] _T_59255; // @[Modules.scala 143:74:@4954.4]
  wire [6:0] _T_59258; // @[Modules.scala 143:103:@4956.4]
  wire [5:0] _T_59259; // @[Modules.scala 143:103:@4957.4]
  wire [5:0] _T_59260; // @[Modules.scala 143:103:@4958.4]
  wire [5:0] _T_59264; // @[Modules.scala 144:80:@4961.4]
  wire [6:0] _T_59265; // @[Modules.scala 143:103:@4962.4]
  wire [5:0] _T_59266; // @[Modules.scala 143:103:@4963.4]
  wire [5:0] _T_59267; // @[Modules.scala 143:103:@4964.4]
  wire [4:0] _T_59269; // @[Modules.scala 143:74:@4966.4]
  wire [5:0] _GEN_142; // @[Modules.scala 143:103:@4968.4]
  wire [6:0] _T_59272; // @[Modules.scala 143:103:@4968.4]
  wire [5:0] _T_59273; // @[Modules.scala 143:103:@4969.4]
  wire [5:0] _T_59274; // @[Modules.scala 143:103:@4970.4]
  wire [5:0] _T_59276; // @[Modules.scala 143:74:@4972.4]
  wire [5:0] _T_59278; // @[Modules.scala 144:80:@4973.4]
  wire [6:0] _T_59279; // @[Modules.scala 143:103:@4974.4]
  wire [5:0] _T_59280; // @[Modules.scala 143:103:@4975.4]
  wire [5:0] _T_59281; // @[Modules.scala 143:103:@4976.4]
  wire [4:0] _T_59290; // @[Modules.scala 143:74:@4984.4]
  wire [4:0] _T_59292; // @[Modules.scala 144:80:@4985.4]
  wire [5:0] _T_59293; // @[Modules.scala 143:103:@4986.4]
  wire [4:0] _T_59294; // @[Modules.scala 143:103:@4987.4]
  wire [4:0] _T_59295; // @[Modules.scala 143:103:@4988.4]
  wire [6:0] _T_59300; // @[Modules.scala 143:103:@4992.4]
  wire [5:0] _T_59301; // @[Modules.scala 143:103:@4993.4]
  wire [5:0] _T_59302; // @[Modules.scala 143:103:@4994.4]
  wire [6:0] _T_59307; // @[Modules.scala 143:103:@4998.4]
  wire [5:0] _T_59308; // @[Modules.scala 143:103:@4999.4]
  wire [5:0] _T_59309; // @[Modules.scala 143:103:@5000.4]
  wire [5:0] _T_59313; // @[Modules.scala 144:80:@5003.4]
  wire [6:0] _T_59314; // @[Modules.scala 143:103:@5004.4]
  wire [5:0] _T_59315; // @[Modules.scala 143:103:@5005.4]
  wire [5:0] _T_59316; // @[Modules.scala 143:103:@5006.4]
  wire [5:0] _T_59318; // @[Modules.scala 143:74:@5008.4]
  wire [5:0] _T_59320; // @[Modules.scala 144:80:@5009.4]
  wire [6:0] _T_59321; // @[Modules.scala 143:103:@5010.4]
  wire [5:0] _T_59322; // @[Modules.scala 143:103:@5011.4]
  wire [5:0] _T_59323; // @[Modules.scala 143:103:@5012.4]
  wire [4:0] _T_59327; // @[Modules.scala 144:80:@5015.4]
  wire [5:0] _GEN_143; // @[Modules.scala 143:103:@5016.4]
  wire [6:0] _T_59328; // @[Modules.scala 143:103:@5016.4]
  wire [5:0] _T_59329; // @[Modules.scala 143:103:@5017.4]
  wire [5:0] _T_59330; // @[Modules.scala 143:103:@5018.4]
  wire [4:0] _T_59332; // @[Modules.scala 143:74:@5020.4]
  wire [4:0] _T_59334; // @[Modules.scala 144:80:@5021.4]
  wire [5:0] _T_59335; // @[Modules.scala 143:103:@5022.4]
  wire [4:0] _T_59336; // @[Modules.scala 143:103:@5023.4]
  wire [4:0] _T_59337; // @[Modules.scala 143:103:@5024.4]
  wire [13:0] buffer_1_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59341; // @[Modules.scala 160:64:@5030.4]
  wire [13:0] _T_59342; // @[Modules.scala 160:64:@5031.4]
  wire [13:0] buffer_1_305; // @[Modules.scala 160:64:@5032.4]
  wire [13:0] buffer_1_4; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_5; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59344; // @[Modules.scala 160:64:@5034.4]
  wire [13:0] _T_59345; // @[Modules.scala 160:64:@5035.4]
  wire [13:0] buffer_1_306; // @[Modules.scala 160:64:@5036.4]
  wire [13:0] buffer_1_6; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_7; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59347; // @[Modules.scala 160:64:@5038.4]
  wire [13:0] _T_59348; // @[Modules.scala 160:64:@5039.4]
  wire [13:0] buffer_1_307; // @[Modules.scala 160:64:@5040.4]
  wire [13:0] buffer_1_8; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59350; // @[Modules.scala 160:64:@5042.4]
  wire [13:0] _T_59351; // @[Modules.scala 160:64:@5043.4]
  wire [13:0] buffer_1_308; // @[Modules.scala 160:64:@5044.4]
  wire [13:0] buffer_1_10; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59353; // @[Modules.scala 160:64:@5046.4]
  wire [13:0] _T_59354; // @[Modules.scala 160:64:@5047.4]
  wire [13:0] buffer_1_309; // @[Modules.scala 160:64:@5048.4]
  wire [13:0] buffer_1_12; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59356; // @[Modules.scala 160:64:@5050.4]
  wire [13:0] _T_59357; // @[Modules.scala 160:64:@5051.4]
  wire [13:0] buffer_1_310; // @[Modules.scala 160:64:@5052.4]
  wire [13:0] buffer_1_14; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_15; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59359; // @[Modules.scala 160:64:@5054.4]
  wire [13:0] _T_59360; // @[Modules.scala 160:64:@5055.4]
  wire [13:0] buffer_1_311; // @[Modules.scala 160:64:@5056.4]
  wire [13:0] buffer_1_16; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_17; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59362; // @[Modules.scala 160:64:@5058.4]
  wire [13:0] _T_59363; // @[Modules.scala 160:64:@5059.4]
  wire [13:0] buffer_1_312; // @[Modules.scala 160:64:@5060.4]
  wire [13:0] buffer_1_18; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_19; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59365; // @[Modules.scala 160:64:@5062.4]
  wire [13:0] _T_59366; // @[Modules.scala 160:64:@5063.4]
  wire [13:0] buffer_1_313; // @[Modules.scala 160:64:@5064.4]
  wire [13:0] buffer_1_20; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59368; // @[Modules.scala 160:64:@5066.4]
  wire [13:0] _T_59369; // @[Modules.scala 160:64:@5067.4]
  wire [13:0] buffer_1_314; // @[Modules.scala 160:64:@5068.4]
  wire [13:0] buffer_1_22; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_23; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59371; // @[Modules.scala 160:64:@5070.4]
  wire [13:0] _T_59372; // @[Modules.scala 160:64:@5071.4]
  wire [13:0] buffer_1_315; // @[Modules.scala 160:64:@5072.4]
  wire [13:0] buffer_1_24; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_25; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59374; // @[Modules.scala 160:64:@5074.4]
  wire [13:0] _T_59375; // @[Modules.scala 160:64:@5075.4]
  wire [13:0] buffer_1_316; // @[Modules.scala 160:64:@5076.4]
  wire [13:0] buffer_1_26; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59377; // @[Modules.scala 160:64:@5078.4]
  wire [13:0] _T_59378; // @[Modules.scala 160:64:@5079.4]
  wire [13:0] buffer_1_317; // @[Modules.scala 160:64:@5080.4]
  wire [13:0] buffer_1_28; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_29; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59380; // @[Modules.scala 160:64:@5082.4]
  wire [13:0] _T_59381; // @[Modules.scala 160:64:@5083.4]
  wire [13:0] buffer_1_318; // @[Modules.scala 160:64:@5084.4]
  wire [13:0] buffer_1_30; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_31; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59383; // @[Modules.scala 160:64:@5086.4]
  wire [13:0] _T_59384; // @[Modules.scala 160:64:@5087.4]
  wire [13:0] buffer_1_319; // @[Modules.scala 160:64:@5088.4]
  wire [13:0] buffer_1_32; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59386; // @[Modules.scala 160:64:@5090.4]
  wire [13:0] _T_59387; // @[Modules.scala 160:64:@5091.4]
  wire [13:0] buffer_1_320; // @[Modules.scala 160:64:@5092.4]
  wire [13:0] buffer_1_34; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59389; // @[Modules.scala 160:64:@5094.4]
  wire [13:0] _T_59390; // @[Modules.scala 160:64:@5095.4]
  wire [13:0] buffer_1_321; // @[Modules.scala 160:64:@5096.4]
  wire [13:0] buffer_1_36; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_37; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59392; // @[Modules.scala 160:64:@5098.4]
  wire [13:0] _T_59393; // @[Modules.scala 160:64:@5099.4]
  wire [13:0] buffer_1_322; // @[Modules.scala 160:64:@5100.4]
  wire [13:0] buffer_1_38; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_39; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59395; // @[Modules.scala 160:64:@5102.4]
  wire [13:0] _T_59396; // @[Modules.scala 160:64:@5103.4]
  wire [13:0] buffer_1_323; // @[Modules.scala 160:64:@5104.4]
  wire [13:0] buffer_1_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59398; // @[Modules.scala 160:64:@5106.4]
  wire [13:0] _T_59399; // @[Modules.scala 160:64:@5107.4]
  wire [13:0] buffer_1_324; // @[Modules.scala 160:64:@5108.4]
  wire [13:0] buffer_1_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59401; // @[Modules.scala 160:64:@5110.4]
  wire [13:0] _T_59402; // @[Modules.scala 160:64:@5111.4]
  wire [13:0] buffer_1_325; // @[Modules.scala 160:64:@5112.4]
  wire [13:0] buffer_1_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59404; // @[Modules.scala 160:64:@5114.4]
  wire [13:0] _T_59405; // @[Modules.scala 160:64:@5115.4]
  wire [13:0] buffer_1_326; // @[Modules.scala 160:64:@5116.4]
  wire [13:0] buffer_1_46; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_47; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59407; // @[Modules.scala 160:64:@5118.4]
  wire [13:0] _T_59408; // @[Modules.scala 160:64:@5119.4]
  wire [13:0] buffer_1_327; // @[Modules.scala 160:64:@5120.4]
  wire [13:0] buffer_1_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59410; // @[Modules.scala 160:64:@5122.4]
  wire [13:0] _T_59411; // @[Modules.scala 160:64:@5123.4]
  wire [13:0] buffer_1_328; // @[Modules.scala 160:64:@5124.4]
  wire [13:0] buffer_1_50; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59413; // @[Modules.scala 160:64:@5126.4]
  wire [13:0] _T_59414; // @[Modules.scala 160:64:@5127.4]
  wire [13:0] buffer_1_329; // @[Modules.scala 160:64:@5128.4]
  wire [13:0] buffer_1_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59416; // @[Modules.scala 160:64:@5130.4]
  wire [13:0] _T_59417; // @[Modules.scala 160:64:@5131.4]
  wire [13:0] buffer_1_330; // @[Modules.scala 160:64:@5132.4]
  wire [13:0] buffer_1_54; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59419; // @[Modules.scala 160:64:@5134.4]
  wire [13:0] _T_59420; // @[Modules.scala 160:64:@5135.4]
  wire [13:0] buffer_1_331; // @[Modules.scala 160:64:@5136.4]
  wire [14:0] _T_59422; // @[Modules.scala 160:64:@5138.4]
  wire [13:0] _T_59423; // @[Modules.scala 160:64:@5139.4]
  wire [13:0] buffer_1_332; // @[Modules.scala 160:64:@5140.4]
  wire [13:0] buffer_1_58; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59425; // @[Modules.scala 160:64:@5142.4]
  wire [13:0] _T_59426; // @[Modules.scala 160:64:@5143.4]
  wire [13:0] buffer_1_333; // @[Modules.scala 160:64:@5144.4]
  wire [13:0] buffer_1_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59428; // @[Modules.scala 160:64:@5146.4]
  wire [13:0] _T_59429; // @[Modules.scala 160:64:@5147.4]
  wire [13:0] buffer_1_334; // @[Modules.scala 160:64:@5148.4]
  wire [13:0] buffer_1_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59431; // @[Modules.scala 160:64:@5150.4]
  wire [13:0] _T_59432; // @[Modules.scala 160:64:@5151.4]
  wire [13:0] buffer_1_335; // @[Modules.scala 160:64:@5152.4]
  wire [13:0] buffer_1_64; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_65; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59434; // @[Modules.scala 160:64:@5154.4]
  wire [13:0] _T_59435; // @[Modules.scala 160:64:@5155.4]
  wire [13:0] buffer_1_336; // @[Modules.scala 160:64:@5156.4]
  wire [13:0] buffer_1_66; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59437; // @[Modules.scala 160:64:@5158.4]
  wire [13:0] _T_59438; // @[Modules.scala 160:64:@5159.4]
  wire [13:0] buffer_1_337; // @[Modules.scala 160:64:@5160.4]
  wire [14:0] _T_59440; // @[Modules.scala 160:64:@5162.4]
  wire [13:0] _T_59441; // @[Modules.scala 160:64:@5163.4]
  wire [13:0] buffer_1_338; // @[Modules.scala 160:64:@5164.4]
  wire [13:0] buffer_1_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59443; // @[Modules.scala 160:64:@5166.4]
  wire [13:0] _T_59444; // @[Modules.scala 160:64:@5167.4]
  wire [13:0] buffer_1_339; // @[Modules.scala 160:64:@5168.4]
  wire [13:0] buffer_1_72; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59446; // @[Modules.scala 160:64:@5170.4]
  wire [13:0] _T_59447; // @[Modules.scala 160:64:@5171.4]
  wire [13:0] buffer_1_340; // @[Modules.scala 160:64:@5172.4]
  wire [13:0] buffer_1_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59449; // @[Modules.scala 160:64:@5174.4]
  wire [13:0] _T_59450; // @[Modules.scala 160:64:@5175.4]
  wire [13:0] buffer_1_341; // @[Modules.scala 160:64:@5176.4]
  wire [14:0] _T_59452; // @[Modules.scala 160:64:@5178.4]
  wire [13:0] _T_59453; // @[Modules.scala 160:64:@5179.4]
  wire [13:0] buffer_1_342; // @[Modules.scala 160:64:@5180.4]
  wire [13:0] buffer_1_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59455; // @[Modules.scala 160:64:@5182.4]
  wire [13:0] _T_59456; // @[Modules.scala 160:64:@5183.4]
  wire [13:0] buffer_1_343; // @[Modules.scala 160:64:@5184.4]
  wire [13:0] buffer_1_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59458; // @[Modules.scala 160:64:@5186.4]
  wire [13:0] _T_59459; // @[Modules.scala 160:64:@5187.4]
  wire [13:0] buffer_1_344; // @[Modules.scala 160:64:@5188.4]
  wire [13:0] buffer_1_82; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_83; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59461; // @[Modules.scala 160:64:@5190.4]
  wire [13:0] _T_59462; // @[Modules.scala 160:64:@5191.4]
  wire [13:0] buffer_1_345; // @[Modules.scala 160:64:@5192.4]
  wire [13:0] buffer_1_84; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59464; // @[Modules.scala 160:64:@5194.4]
  wire [13:0] _T_59465; // @[Modules.scala 160:64:@5195.4]
  wire [13:0] buffer_1_346; // @[Modules.scala 160:64:@5196.4]
  wire [13:0] buffer_1_86; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59467; // @[Modules.scala 160:64:@5198.4]
  wire [13:0] _T_59468; // @[Modules.scala 160:64:@5199.4]
  wire [13:0] buffer_1_347; // @[Modules.scala 160:64:@5200.4]
  wire [13:0] buffer_1_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59473; // @[Modules.scala 160:64:@5206.4]
  wire [13:0] _T_59474; // @[Modules.scala 160:64:@5207.4]
  wire [13:0] buffer_1_349; // @[Modules.scala 160:64:@5208.4]
  wire [13:0] buffer_1_92; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59476; // @[Modules.scala 160:64:@5210.4]
  wire [13:0] _T_59477; // @[Modules.scala 160:64:@5211.4]
  wire [13:0] buffer_1_350; // @[Modules.scala 160:64:@5212.4]
  wire [13:0] buffer_1_94; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59479; // @[Modules.scala 160:64:@5214.4]
  wire [13:0] _T_59480; // @[Modules.scala 160:64:@5215.4]
  wire [13:0] buffer_1_351; // @[Modules.scala 160:64:@5216.4]
  wire [13:0] buffer_1_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59482; // @[Modules.scala 160:64:@5218.4]
  wire [13:0] _T_59483; // @[Modules.scala 160:64:@5219.4]
  wire [13:0] buffer_1_352; // @[Modules.scala 160:64:@5220.4]
  wire [13:0] buffer_1_98; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_99; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59485; // @[Modules.scala 160:64:@5222.4]
  wire [13:0] _T_59486; // @[Modules.scala 160:64:@5223.4]
  wire [13:0] buffer_1_353; // @[Modules.scala 160:64:@5224.4]
  wire [14:0] _T_59488; // @[Modules.scala 160:64:@5226.4]
  wire [13:0] _T_59489; // @[Modules.scala 160:64:@5227.4]
  wire [13:0] buffer_1_354; // @[Modules.scala 160:64:@5228.4]
  wire [13:0] buffer_1_102; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59491; // @[Modules.scala 160:64:@5230.4]
  wire [13:0] _T_59492; // @[Modules.scala 160:64:@5231.4]
  wire [13:0] buffer_1_355; // @[Modules.scala 160:64:@5232.4]
  wire [13:0] buffer_1_104; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59494; // @[Modules.scala 160:64:@5234.4]
  wire [13:0] _T_59495; // @[Modules.scala 160:64:@5235.4]
  wire [13:0] buffer_1_356; // @[Modules.scala 160:64:@5236.4]
  wire [13:0] buffer_1_106; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59497; // @[Modules.scala 160:64:@5238.4]
  wire [13:0] _T_59498; // @[Modules.scala 160:64:@5239.4]
  wire [13:0] buffer_1_357; // @[Modules.scala 160:64:@5240.4]
  wire [13:0] buffer_1_108; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_109; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59500; // @[Modules.scala 160:64:@5242.4]
  wire [13:0] _T_59501; // @[Modules.scala 160:64:@5243.4]
  wire [13:0] buffer_1_358; // @[Modules.scala 160:64:@5244.4]
  wire [13:0] buffer_1_110; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59503; // @[Modules.scala 160:64:@5246.4]
  wire [13:0] _T_59504; // @[Modules.scala 160:64:@5247.4]
  wire [13:0] buffer_1_359; // @[Modules.scala 160:64:@5248.4]
  wire [13:0] buffer_1_112; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59506; // @[Modules.scala 160:64:@5250.4]
  wire [13:0] _T_59507; // @[Modules.scala 160:64:@5251.4]
  wire [13:0] buffer_1_360; // @[Modules.scala 160:64:@5252.4]
  wire [13:0] buffer_1_114; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59509; // @[Modules.scala 160:64:@5254.4]
  wire [13:0] _T_59510; // @[Modules.scala 160:64:@5255.4]
  wire [13:0] buffer_1_361; // @[Modules.scala 160:64:@5256.4]
  wire [13:0] buffer_1_116; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59512; // @[Modules.scala 160:64:@5258.4]
  wire [13:0] _T_59513; // @[Modules.scala 160:64:@5259.4]
  wire [13:0] buffer_1_362; // @[Modules.scala 160:64:@5260.4]
  wire [13:0] buffer_1_118; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_119; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59515; // @[Modules.scala 160:64:@5262.4]
  wire [13:0] _T_59516; // @[Modules.scala 160:64:@5263.4]
  wire [13:0] buffer_1_363; // @[Modules.scala 160:64:@5264.4]
  wire [13:0] buffer_1_120; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59518; // @[Modules.scala 160:64:@5266.4]
  wire [13:0] _T_59519; // @[Modules.scala 160:64:@5267.4]
  wire [13:0] buffer_1_364; // @[Modules.scala 160:64:@5268.4]
  wire [13:0] buffer_1_122; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59521; // @[Modules.scala 160:64:@5270.4]
  wire [13:0] _T_59522; // @[Modules.scala 160:64:@5271.4]
  wire [13:0] buffer_1_365; // @[Modules.scala 160:64:@5272.4]
  wire [13:0] buffer_1_124; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59524; // @[Modules.scala 160:64:@5274.4]
  wire [13:0] _T_59525; // @[Modules.scala 160:64:@5275.4]
  wire [13:0] buffer_1_366; // @[Modules.scala 160:64:@5276.4]
  wire [13:0] buffer_1_126; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_127; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59527; // @[Modules.scala 160:64:@5278.4]
  wire [13:0] _T_59528; // @[Modules.scala 160:64:@5279.4]
  wire [13:0] buffer_1_367; // @[Modules.scala 160:64:@5280.4]
  wire [13:0] buffer_1_128; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_129; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59530; // @[Modules.scala 160:64:@5282.4]
  wire [13:0] _T_59531; // @[Modules.scala 160:64:@5283.4]
  wire [13:0] buffer_1_368; // @[Modules.scala 160:64:@5284.4]
  wire [13:0] buffer_1_130; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59533; // @[Modules.scala 160:64:@5286.4]
  wire [13:0] _T_59534; // @[Modules.scala 160:64:@5287.4]
  wire [13:0] buffer_1_369; // @[Modules.scala 160:64:@5288.4]
  wire [13:0] buffer_1_132; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59536; // @[Modules.scala 160:64:@5290.4]
  wire [13:0] _T_59537; // @[Modules.scala 160:64:@5291.4]
  wire [13:0] buffer_1_370; // @[Modules.scala 160:64:@5292.4]
  wire [13:0] buffer_1_134; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59539; // @[Modules.scala 160:64:@5294.4]
  wire [13:0] _T_59540; // @[Modules.scala 160:64:@5295.4]
  wire [13:0] buffer_1_371; // @[Modules.scala 160:64:@5296.4]
  wire [13:0] buffer_1_136; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59542; // @[Modules.scala 160:64:@5298.4]
  wire [13:0] _T_59543; // @[Modules.scala 160:64:@5299.4]
  wire [13:0] buffer_1_372; // @[Modules.scala 160:64:@5300.4]
  wire [13:0] buffer_1_138; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_139; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59545; // @[Modules.scala 160:64:@5302.4]
  wire [13:0] _T_59546; // @[Modules.scala 160:64:@5303.4]
  wire [13:0] buffer_1_373; // @[Modules.scala 160:64:@5304.4]
  wire [13:0] buffer_1_140; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59548; // @[Modules.scala 160:64:@5306.4]
  wire [13:0] _T_59549; // @[Modules.scala 160:64:@5307.4]
  wire [13:0] buffer_1_374; // @[Modules.scala 160:64:@5308.4]
  wire [13:0] buffer_1_142; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_143; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59551; // @[Modules.scala 160:64:@5310.4]
  wire [13:0] _T_59552; // @[Modules.scala 160:64:@5311.4]
  wire [13:0] buffer_1_375; // @[Modules.scala 160:64:@5312.4]
  wire [13:0] buffer_1_144; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59554; // @[Modules.scala 160:64:@5314.4]
  wire [13:0] _T_59555; // @[Modules.scala 160:64:@5315.4]
  wire [13:0] buffer_1_376; // @[Modules.scala 160:64:@5316.4]
  wire [13:0] buffer_1_146; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59557; // @[Modules.scala 160:64:@5318.4]
  wire [13:0] _T_59558; // @[Modules.scala 160:64:@5319.4]
  wire [13:0] buffer_1_377; // @[Modules.scala 160:64:@5320.4]
  wire [13:0] buffer_1_148; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59560; // @[Modules.scala 160:64:@5322.4]
  wire [13:0] _T_59561; // @[Modules.scala 160:64:@5323.4]
  wire [13:0] buffer_1_378; // @[Modules.scala 160:64:@5324.4]
  wire [13:0] buffer_1_150; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59563; // @[Modules.scala 160:64:@5326.4]
  wire [13:0] _T_59564; // @[Modules.scala 160:64:@5327.4]
  wire [13:0] buffer_1_379; // @[Modules.scala 160:64:@5328.4]
  wire [13:0] buffer_1_152; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59566; // @[Modules.scala 160:64:@5330.4]
  wire [13:0] _T_59567; // @[Modules.scala 160:64:@5331.4]
  wire [13:0] buffer_1_380; // @[Modules.scala 160:64:@5332.4]
  wire [13:0] buffer_1_154; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59569; // @[Modules.scala 160:64:@5334.4]
  wire [13:0] _T_59570; // @[Modules.scala 160:64:@5335.4]
  wire [13:0] buffer_1_381; // @[Modules.scala 160:64:@5336.4]
  wire [13:0] buffer_1_156; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59572; // @[Modules.scala 160:64:@5338.4]
  wire [13:0] _T_59573; // @[Modules.scala 160:64:@5339.4]
  wire [13:0] buffer_1_382; // @[Modules.scala 160:64:@5340.4]
  wire [13:0] buffer_1_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59575; // @[Modules.scala 160:64:@5342.4]
  wire [13:0] _T_59576; // @[Modules.scala 160:64:@5343.4]
  wire [13:0] buffer_1_383; // @[Modules.scala 160:64:@5344.4]
  wire [13:0] buffer_1_160; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59578; // @[Modules.scala 160:64:@5346.4]
  wire [13:0] _T_59579; // @[Modules.scala 160:64:@5347.4]
  wire [13:0] buffer_1_384; // @[Modules.scala 160:64:@5348.4]
  wire [13:0] buffer_1_162; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_163; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59581; // @[Modules.scala 160:64:@5350.4]
  wire [13:0] _T_59582; // @[Modules.scala 160:64:@5351.4]
  wire [13:0] buffer_1_385; // @[Modules.scala 160:64:@5352.4]
  wire [13:0] buffer_1_164; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59584; // @[Modules.scala 160:64:@5354.4]
  wire [13:0] _T_59585; // @[Modules.scala 160:64:@5355.4]
  wire [13:0] buffer_1_386; // @[Modules.scala 160:64:@5356.4]
  wire [13:0] buffer_1_166; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59587; // @[Modules.scala 160:64:@5358.4]
  wire [13:0] _T_59588; // @[Modules.scala 160:64:@5359.4]
  wire [13:0] buffer_1_387; // @[Modules.scala 160:64:@5360.4]
  wire [13:0] buffer_1_168; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59590; // @[Modules.scala 160:64:@5362.4]
  wire [13:0] _T_59591; // @[Modules.scala 160:64:@5363.4]
  wire [13:0] buffer_1_388; // @[Modules.scala 160:64:@5364.4]
  wire [13:0] buffer_1_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59593; // @[Modules.scala 160:64:@5366.4]
  wire [13:0] _T_59594; // @[Modules.scala 160:64:@5367.4]
  wire [13:0] buffer_1_389; // @[Modules.scala 160:64:@5368.4]
  wire [13:0] buffer_1_172; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_173; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59596; // @[Modules.scala 160:64:@5370.4]
  wire [13:0] _T_59597; // @[Modules.scala 160:64:@5371.4]
  wire [13:0] buffer_1_390; // @[Modules.scala 160:64:@5372.4]
  wire [13:0] buffer_1_174; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59599; // @[Modules.scala 160:64:@5374.4]
  wire [13:0] _T_59600; // @[Modules.scala 160:64:@5375.4]
  wire [13:0] buffer_1_391; // @[Modules.scala 160:64:@5376.4]
  wire [13:0] buffer_1_176; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59602; // @[Modules.scala 160:64:@5378.4]
  wire [13:0] _T_59603; // @[Modules.scala 160:64:@5379.4]
  wire [13:0] buffer_1_392; // @[Modules.scala 160:64:@5380.4]
  wire [13:0] buffer_1_178; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_179; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59605; // @[Modules.scala 160:64:@5382.4]
  wire [13:0] _T_59606; // @[Modules.scala 160:64:@5383.4]
  wire [13:0] buffer_1_393; // @[Modules.scala 160:64:@5384.4]
  wire [13:0] buffer_1_180; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59608; // @[Modules.scala 160:64:@5386.4]
  wire [13:0] _T_59609; // @[Modules.scala 160:64:@5387.4]
  wire [13:0] buffer_1_394; // @[Modules.scala 160:64:@5388.4]
  wire [13:0] buffer_1_182; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59611; // @[Modules.scala 160:64:@5390.4]
  wire [13:0] _T_59612; // @[Modules.scala 160:64:@5391.4]
  wire [13:0] buffer_1_395; // @[Modules.scala 160:64:@5392.4]
  wire [13:0] buffer_1_184; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59614; // @[Modules.scala 160:64:@5394.4]
  wire [13:0] _T_59615; // @[Modules.scala 160:64:@5395.4]
  wire [13:0] buffer_1_396; // @[Modules.scala 160:64:@5396.4]
  wire [13:0] buffer_1_187; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59617; // @[Modules.scala 160:64:@5398.4]
  wire [13:0] _T_59618; // @[Modules.scala 160:64:@5399.4]
  wire [13:0] buffer_1_397; // @[Modules.scala 160:64:@5400.4]
  wire [13:0] buffer_1_188; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59620; // @[Modules.scala 160:64:@5402.4]
  wire [13:0] _T_59621; // @[Modules.scala 160:64:@5403.4]
  wire [13:0] buffer_1_398; // @[Modules.scala 160:64:@5404.4]
  wire [13:0] buffer_1_190; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59623; // @[Modules.scala 160:64:@5406.4]
  wire [13:0] _T_59624; // @[Modules.scala 160:64:@5407.4]
  wire [13:0] buffer_1_399; // @[Modules.scala 160:64:@5408.4]
  wire [13:0] buffer_1_192; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59626; // @[Modules.scala 160:64:@5410.4]
  wire [13:0] _T_59627; // @[Modules.scala 160:64:@5411.4]
  wire [13:0] buffer_1_400; // @[Modules.scala 160:64:@5412.4]
  wire [13:0] buffer_1_194; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59629; // @[Modules.scala 160:64:@5414.4]
  wire [13:0] _T_59630; // @[Modules.scala 160:64:@5415.4]
  wire [13:0] buffer_1_401; // @[Modules.scala 160:64:@5416.4]
  wire [13:0] buffer_1_196; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59632; // @[Modules.scala 160:64:@5418.4]
  wire [13:0] _T_59633; // @[Modules.scala 160:64:@5419.4]
  wire [13:0] buffer_1_402; // @[Modules.scala 160:64:@5420.4]
  wire [13:0] buffer_1_198; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59635; // @[Modules.scala 160:64:@5422.4]
  wire [13:0] _T_59636; // @[Modules.scala 160:64:@5423.4]
  wire [13:0] buffer_1_403; // @[Modules.scala 160:64:@5424.4]
  wire [13:0] buffer_1_200; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59638; // @[Modules.scala 160:64:@5426.4]
  wire [13:0] _T_59639; // @[Modules.scala 160:64:@5427.4]
  wire [13:0] buffer_1_404; // @[Modules.scala 160:64:@5428.4]
  wire [13:0] buffer_1_202; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59641; // @[Modules.scala 160:64:@5430.4]
  wire [13:0] _T_59642; // @[Modules.scala 160:64:@5431.4]
  wire [13:0] buffer_1_405; // @[Modules.scala 160:64:@5432.4]
  wire [13:0] buffer_1_204; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59644; // @[Modules.scala 160:64:@5434.4]
  wire [13:0] _T_59645; // @[Modules.scala 160:64:@5435.4]
  wire [13:0] buffer_1_406; // @[Modules.scala 160:64:@5436.4]
  wire [13:0] buffer_1_206; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59647; // @[Modules.scala 160:64:@5438.4]
  wire [13:0] _T_59648; // @[Modules.scala 160:64:@5439.4]
  wire [13:0] buffer_1_407; // @[Modules.scala 160:64:@5440.4]
  wire [13:0] buffer_1_208; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_209; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59650; // @[Modules.scala 160:64:@5442.4]
  wire [13:0] _T_59651; // @[Modules.scala 160:64:@5443.4]
  wire [13:0] buffer_1_408; // @[Modules.scala 160:64:@5444.4]
  wire [13:0] buffer_1_210; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59653; // @[Modules.scala 160:64:@5446.4]
  wire [13:0] _T_59654; // @[Modules.scala 160:64:@5447.4]
  wire [13:0] buffer_1_409; // @[Modules.scala 160:64:@5448.4]
  wire [13:0] buffer_1_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59656; // @[Modules.scala 160:64:@5450.4]
  wire [13:0] _T_59657; // @[Modules.scala 160:64:@5451.4]
  wire [13:0] buffer_1_410; // @[Modules.scala 160:64:@5452.4]
  wire [13:0] buffer_1_214; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59659; // @[Modules.scala 160:64:@5454.4]
  wire [13:0] _T_59660; // @[Modules.scala 160:64:@5455.4]
  wire [13:0] buffer_1_411; // @[Modules.scala 160:64:@5456.4]
  wire [13:0] buffer_1_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59662; // @[Modules.scala 160:64:@5458.4]
  wire [13:0] _T_59663; // @[Modules.scala 160:64:@5459.4]
  wire [13:0] buffer_1_412; // @[Modules.scala 160:64:@5460.4]
  wire [13:0] buffer_1_218; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59665; // @[Modules.scala 160:64:@5462.4]
  wire [13:0] _T_59666; // @[Modules.scala 160:64:@5463.4]
  wire [13:0] buffer_1_413; // @[Modules.scala 160:64:@5464.4]
  wire [13:0] buffer_1_220; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_221; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59668; // @[Modules.scala 160:64:@5466.4]
  wire [13:0] _T_59669; // @[Modules.scala 160:64:@5467.4]
  wire [13:0] buffer_1_414; // @[Modules.scala 160:64:@5468.4]
  wire [13:0] buffer_1_222; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59671; // @[Modules.scala 160:64:@5470.4]
  wire [13:0] _T_59672; // @[Modules.scala 160:64:@5471.4]
  wire [13:0] buffer_1_415; // @[Modules.scala 160:64:@5472.4]
  wire [13:0] buffer_1_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59674; // @[Modules.scala 160:64:@5474.4]
  wire [13:0] _T_59675; // @[Modules.scala 160:64:@5475.4]
  wire [13:0] buffer_1_416; // @[Modules.scala 160:64:@5476.4]
  wire [13:0] buffer_1_226; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59677; // @[Modules.scala 160:64:@5478.4]
  wire [13:0] _T_59678; // @[Modules.scala 160:64:@5479.4]
  wire [13:0] buffer_1_417; // @[Modules.scala 160:64:@5480.4]
  wire [13:0] buffer_1_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59680; // @[Modules.scala 160:64:@5482.4]
  wire [13:0] _T_59681; // @[Modules.scala 160:64:@5483.4]
  wire [13:0] buffer_1_418; // @[Modules.scala 160:64:@5484.4]
  wire [13:0] buffer_1_232; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59686; // @[Modules.scala 160:64:@5490.4]
  wire [13:0] _T_59687; // @[Modules.scala 160:64:@5491.4]
  wire [13:0] buffer_1_420; // @[Modules.scala 160:64:@5492.4]
  wire [13:0] buffer_1_234; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59689; // @[Modules.scala 160:64:@5494.4]
  wire [13:0] _T_59690; // @[Modules.scala 160:64:@5495.4]
  wire [13:0] buffer_1_421; // @[Modules.scala 160:64:@5496.4]
  wire [13:0] buffer_1_236; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59692; // @[Modules.scala 160:64:@5498.4]
  wire [13:0] _T_59693; // @[Modules.scala 160:64:@5499.4]
  wire [13:0] buffer_1_422; // @[Modules.scala 160:64:@5500.4]
  wire [13:0] buffer_1_238; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59695; // @[Modules.scala 160:64:@5502.4]
  wire [13:0] _T_59696; // @[Modules.scala 160:64:@5503.4]
  wire [13:0] buffer_1_423; // @[Modules.scala 160:64:@5504.4]
  wire [13:0] buffer_1_240; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59698; // @[Modules.scala 160:64:@5506.4]
  wire [13:0] _T_59699; // @[Modules.scala 160:64:@5507.4]
  wire [13:0] buffer_1_424; // @[Modules.scala 160:64:@5508.4]
  wire [13:0] buffer_1_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59701; // @[Modules.scala 160:64:@5510.4]
  wire [13:0] _T_59702; // @[Modules.scala 160:64:@5511.4]
  wire [13:0] buffer_1_425; // @[Modules.scala 160:64:@5512.4]
  wire [13:0] buffer_1_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59704; // @[Modules.scala 160:64:@5514.4]
  wire [13:0] _T_59705; // @[Modules.scala 160:64:@5515.4]
  wire [13:0] buffer_1_426; // @[Modules.scala 160:64:@5516.4]
  wire [13:0] buffer_1_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59707; // @[Modules.scala 160:64:@5518.4]
  wire [13:0] _T_59708; // @[Modules.scala 160:64:@5519.4]
  wire [13:0] buffer_1_427; // @[Modules.scala 160:64:@5520.4]
  wire [13:0] buffer_1_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59710; // @[Modules.scala 160:64:@5522.4]
  wire [13:0] _T_59711; // @[Modules.scala 160:64:@5523.4]
  wire [13:0] buffer_1_428; // @[Modules.scala 160:64:@5524.4]
  wire [13:0] buffer_1_250; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59713; // @[Modules.scala 160:64:@5526.4]
  wire [13:0] _T_59714; // @[Modules.scala 160:64:@5527.4]
  wire [13:0] buffer_1_429; // @[Modules.scala 160:64:@5528.4]
  wire [13:0] buffer_1_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59716; // @[Modules.scala 160:64:@5530.4]
  wire [13:0] _T_59717; // @[Modules.scala 160:64:@5531.4]
  wire [13:0] buffer_1_430; // @[Modules.scala 160:64:@5532.4]
  wire [13:0] buffer_1_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59719; // @[Modules.scala 160:64:@5534.4]
  wire [13:0] _T_59720; // @[Modules.scala 160:64:@5535.4]
  wire [13:0] buffer_1_431; // @[Modules.scala 160:64:@5536.4]
  wire [13:0] buffer_1_256; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59722; // @[Modules.scala 160:64:@5538.4]
  wire [13:0] _T_59723; // @[Modules.scala 160:64:@5539.4]
  wire [13:0] buffer_1_432; // @[Modules.scala 160:64:@5540.4]
  wire [13:0] buffer_1_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59725; // @[Modules.scala 160:64:@5542.4]
  wire [13:0] _T_59726; // @[Modules.scala 160:64:@5543.4]
  wire [13:0] buffer_1_433; // @[Modules.scala 160:64:@5544.4]
  wire [13:0] buffer_1_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59728; // @[Modules.scala 160:64:@5546.4]
  wire [13:0] _T_59729; // @[Modules.scala 160:64:@5547.4]
  wire [13:0] buffer_1_434; // @[Modules.scala 160:64:@5548.4]
  wire [13:0] buffer_1_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59731; // @[Modules.scala 160:64:@5550.4]
  wire [13:0] _T_59732; // @[Modules.scala 160:64:@5551.4]
  wire [13:0] buffer_1_435; // @[Modules.scala 160:64:@5552.4]
  wire [13:0] buffer_1_264; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59734; // @[Modules.scala 160:64:@5554.4]
  wire [13:0] _T_59735; // @[Modules.scala 160:64:@5555.4]
  wire [13:0] buffer_1_436; // @[Modules.scala 160:64:@5556.4]
  wire [13:0] buffer_1_266; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_267; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59737; // @[Modules.scala 160:64:@5558.4]
  wire [13:0] _T_59738; // @[Modules.scala 160:64:@5559.4]
  wire [13:0] buffer_1_437; // @[Modules.scala 160:64:@5560.4]
  wire [13:0] buffer_1_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59740; // @[Modules.scala 160:64:@5562.4]
  wire [13:0] _T_59741; // @[Modules.scala 160:64:@5563.4]
  wire [13:0] buffer_1_438; // @[Modules.scala 160:64:@5564.4]
  wire [13:0] buffer_1_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59743; // @[Modules.scala 160:64:@5566.4]
  wire [13:0] _T_59744; // @[Modules.scala 160:64:@5567.4]
  wire [13:0] buffer_1_439; // @[Modules.scala 160:64:@5568.4]
  wire [13:0] buffer_1_272; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59746; // @[Modules.scala 160:64:@5570.4]
  wire [13:0] _T_59747; // @[Modules.scala 160:64:@5571.4]
  wire [13:0] buffer_1_440; // @[Modules.scala 160:64:@5572.4]
  wire [13:0] buffer_1_274; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_275; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59749; // @[Modules.scala 160:64:@5574.4]
  wire [13:0] _T_59750; // @[Modules.scala 160:64:@5575.4]
  wire [13:0] buffer_1_441; // @[Modules.scala 160:64:@5576.4]
  wire [13:0] buffer_1_276; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_277; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59752; // @[Modules.scala 160:64:@5578.4]
  wire [13:0] _T_59753; // @[Modules.scala 160:64:@5579.4]
  wire [13:0] buffer_1_442; // @[Modules.scala 160:64:@5580.4]
  wire [13:0] buffer_1_278; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59755; // @[Modules.scala 160:64:@5582.4]
  wire [13:0] _T_59756; // @[Modules.scala 160:64:@5583.4]
  wire [13:0] buffer_1_443; // @[Modules.scala 160:64:@5584.4]
  wire [13:0] buffer_1_280; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59758; // @[Modules.scala 160:64:@5586.4]
  wire [13:0] _T_59759; // @[Modules.scala 160:64:@5587.4]
  wire [13:0] buffer_1_444; // @[Modules.scala 160:64:@5588.4]
  wire [13:0] buffer_1_282; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59761; // @[Modules.scala 160:64:@5590.4]
  wire [13:0] _T_59762; // @[Modules.scala 160:64:@5591.4]
  wire [13:0] buffer_1_445; // @[Modules.scala 160:64:@5592.4]
  wire [13:0] buffer_1_284; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_285; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59764; // @[Modules.scala 160:64:@5594.4]
  wire [13:0] _T_59765; // @[Modules.scala 160:64:@5595.4]
  wire [13:0] buffer_1_446; // @[Modules.scala 160:64:@5596.4]
  wire [13:0] buffer_1_288; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59770; // @[Modules.scala 160:64:@5602.4]
  wire [13:0] _T_59771; // @[Modules.scala 160:64:@5603.4]
  wire [13:0] buffer_1_448; // @[Modules.scala 160:64:@5604.4]
  wire [13:0] buffer_1_290; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59773; // @[Modules.scala 160:64:@5606.4]
  wire [13:0] _T_59774; // @[Modules.scala 160:64:@5607.4]
  wire [13:0] buffer_1_449; // @[Modules.scala 160:64:@5608.4]
  wire [13:0] buffer_1_292; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59776; // @[Modules.scala 160:64:@5610.4]
  wire [13:0] _T_59777; // @[Modules.scala 160:64:@5611.4]
  wire [13:0] buffer_1_450; // @[Modules.scala 160:64:@5612.4]
  wire [13:0] buffer_1_294; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59779; // @[Modules.scala 160:64:@5614.4]
  wire [13:0] _T_59780; // @[Modules.scala 160:64:@5615.4]
  wire [13:0] buffer_1_451; // @[Modules.scala 160:64:@5616.4]
  wire [13:0] buffer_1_297; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59782; // @[Modules.scala 160:64:@5618.4]
  wire [13:0] _T_59783; // @[Modules.scala 160:64:@5619.4]
  wire [13:0] buffer_1_452; // @[Modules.scala 160:64:@5620.4]
  wire [13:0] buffer_1_298; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59785; // @[Modules.scala 160:64:@5622.4]
  wire [13:0] _T_59786; // @[Modules.scala 160:64:@5623.4]
  wire [13:0] buffer_1_453; // @[Modules.scala 160:64:@5624.4]
  wire [13:0] buffer_1_300; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_301; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59788; // @[Modules.scala 160:64:@5626.4]
  wire [13:0] _T_59789; // @[Modules.scala 160:64:@5627.4]
  wire [13:0] buffer_1_454; // @[Modules.scala 160:64:@5628.4]
  wire [13:0] buffer_1_302; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_1_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_59791; // @[Modules.scala 160:64:@5630.4]
  wire [13:0] _T_59792; // @[Modules.scala 160:64:@5631.4]
  wire [13:0] buffer_1_455; // @[Modules.scala 160:64:@5632.4]
  wire [14:0] _T_59794; // @[Modules.scala 160:64:@5634.4]
  wire [13:0] _T_59795; // @[Modules.scala 160:64:@5635.4]
  wire [13:0] buffer_1_456; // @[Modules.scala 160:64:@5636.4]
  wire [14:0] _T_59797; // @[Modules.scala 160:64:@5638.4]
  wire [13:0] _T_59798; // @[Modules.scala 160:64:@5639.4]
  wire [13:0] buffer_1_457; // @[Modules.scala 160:64:@5640.4]
  wire [14:0] _T_59800; // @[Modules.scala 160:64:@5642.4]
  wire [13:0] _T_59801; // @[Modules.scala 160:64:@5643.4]
  wire [13:0] buffer_1_458; // @[Modules.scala 160:64:@5644.4]
  wire [14:0] _T_59803; // @[Modules.scala 160:64:@5646.4]
  wire [13:0] _T_59804; // @[Modules.scala 160:64:@5647.4]
  wire [13:0] buffer_1_459; // @[Modules.scala 160:64:@5648.4]
  wire [14:0] _T_59806; // @[Modules.scala 160:64:@5650.4]
  wire [13:0] _T_59807; // @[Modules.scala 160:64:@5651.4]
  wire [13:0] buffer_1_460; // @[Modules.scala 160:64:@5652.4]
  wire [14:0] _T_59809; // @[Modules.scala 160:64:@5654.4]
  wire [13:0] _T_59810; // @[Modules.scala 160:64:@5655.4]
  wire [13:0] buffer_1_461; // @[Modules.scala 160:64:@5656.4]
  wire [14:0] _T_59812; // @[Modules.scala 160:64:@5658.4]
  wire [13:0] _T_59813; // @[Modules.scala 160:64:@5659.4]
  wire [13:0] buffer_1_462; // @[Modules.scala 160:64:@5660.4]
  wire [14:0] _T_59815; // @[Modules.scala 160:64:@5662.4]
  wire [13:0] _T_59816; // @[Modules.scala 160:64:@5663.4]
  wire [13:0] buffer_1_463; // @[Modules.scala 160:64:@5664.4]
  wire [14:0] _T_59818; // @[Modules.scala 160:64:@5666.4]
  wire [13:0] _T_59819; // @[Modules.scala 160:64:@5667.4]
  wire [13:0] buffer_1_464; // @[Modules.scala 160:64:@5668.4]
  wire [14:0] _T_59821; // @[Modules.scala 160:64:@5670.4]
  wire [13:0] _T_59822; // @[Modules.scala 160:64:@5671.4]
  wire [13:0] buffer_1_465; // @[Modules.scala 160:64:@5672.4]
  wire [14:0] _T_59824; // @[Modules.scala 160:64:@5674.4]
  wire [13:0] _T_59825; // @[Modules.scala 160:64:@5675.4]
  wire [13:0] buffer_1_466; // @[Modules.scala 160:64:@5676.4]
  wire [14:0] _T_59827; // @[Modules.scala 160:64:@5678.4]
  wire [13:0] _T_59828; // @[Modules.scala 160:64:@5679.4]
  wire [13:0] buffer_1_467; // @[Modules.scala 160:64:@5680.4]
  wire [14:0] _T_59830; // @[Modules.scala 160:64:@5682.4]
  wire [13:0] _T_59831; // @[Modules.scala 160:64:@5683.4]
  wire [13:0] buffer_1_468; // @[Modules.scala 160:64:@5684.4]
  wire [14:0] _T_59833; // @[Modules.scala 160:64:@5686.4]
  wire [13:0] _T_59834; // @[Modules.scala 160:64:@5687.4]
  wire [13:0] buffer_1_469; // @[Modules.scala 160:64:@5688.4]
  wire [14:0] _T_59836; // @[Modules.scala 160:64:@5690.4]
  wire [13:0] _T_59837; // @[Modules.scala 160:64:@5691.4]
  wire [13:0] buffer_1_470; // @[Modules.scala 160:64:@5692.4]
  wire [14:0] _T_59839; // @[Modules.scala 160:64:@5694.4]
  wire [13:0] _T_59840; // @[Modules.scala 160:64:@5695.4]
  wire [13:0] buffer_1_471; // @[Modules.scala 160:64:@5696.4]
  wire [14:0] _T_59842; // @[Modules.scala 160:64:@5698.4]
  wire [13:0] _T_59843; // @[Modules.scala 160:64:@5699.4]
  wire [13:0] buffer_1_472; // @[Modules.scala 160:64:@5700.4]
  wire [14:0] _T_59845; // @[Modules.scala 160:64:@5702.4]
  wire [13:0] _T_59846; // @[Modules.scala 160:64:@5703.4]
  wire [13:0] buffer_1_473; // @[Modules.scala 160:64:@5704.4]
  wire [14:0] _T_59848; // @[Modules.scala 160:64:@5706.4]
  wire [13:0] _T_59849; // @[Modules.scala 160:64:@5707.4]
  wire [13:0] buffer_1_474; // @[Modules.scala 160:64:@5708.4]
  wire [14:0] _T_59851; // @[Modules.scala 160:64:@5710.4]
  wire [13:0] _T_59852; // @[Modules.scala 160:64:@5711.4]
  wire [13:0] buffer_1_475; // @[Modules.scala 160:64:@5712.4]
  wire [14:0] _T_59854; // @[Modules.scala 160:64:@5714.4]
  wire [13:0] _T_59855; // @[Modules.scala 160:64:@5715.4]
  wire [13:0] buffer_1_476; // @[Modules.scala 160:64:@5716.4]
  wire [14:0] _T_59857; // @[Modules.scala 160:64:@5718.4]
  wire [13:0] _T_59858; // @[Modules.scala 160:64:@5719.4]
  wire [13:0] buffer_1_477; // @[Modules.scala 160:64:@5720.4]
  wire [14:0] _T_59860; // @[Modules.scala 160:64:@5722.4]
  wire [13:0] _T_59861; // @[Modules.scala 160:64:@5723.4]
  wire [13:0] buffer_1_478; // @[Modules.scala 160:64:@5724.4]
  wire [14:0] _T_59863; // @[Modules.scala 160:64:@5726.4]
  wire [13:0] _T_59864; // @[Modules.scala 160:64:@5727.4]
  wire [13:0] buffer_1_479; // @[Modules.scala 160:64:@5728.4]
  wire [14:0] _T_59866; // @[Modules.scala 160:64:@5730.4]
  wire [13:0] _T_59867; // @[Modules.scala 160:64:@5731.4]
  wire [13:0] buffer_1_480; // @[Modules.scala 160:64:@5732.4]
  wire [14:0] _T_59869; // @[Modules.scala 160:64:@5734.4]
  wire [13:0] _T_59870; // @[Modules.scala 160:64:@5735.4]
  wire [13:0] buffer_1_481; // @[Modules.scala 160:64:@5736.4]
  wire [14:0] _T_59872; // @[Modules.scala 160:64:@5738.4]
  wire [13:0] _T_59873; // @[Modules.scala 160:64:@5739.4]
  wire [13:0] buffer_1_482; // @[Modules.scala 160:64:@5740.4]
  wire [14:0] _T_59875; // @[Modules.scala 160:64:@5742.4]
  wire [13:0] _T_59876; // @[Modules.scala 160:64:@5743.4]
  wire [13:0] buffer_1_483; // @[Modules.scala 160:64:@5744.4]
  wire [14:0] _T_59878; // @[Modules.scala 160:64:@5746.4]
  wire [13:0] _T_59879; // @[Modules.scala 160:64:@5747.4]
  wire [13:0] buffer_1_484; // @[Modules.scala 160:64:@5748.4]
  wire [14:0] _T_59881; // @[Modules.scala 160:64:@5750.4]
  wire [13:0] _T_59882; // @[Modules.scala 160:64:@5751.4]
  wire [13:0] buffer_1_485; // @[Modules.scala 160:64:@5752.4]
  wire [14:0] _T_59884; // @[Modules.scala 160:64:@5754.4]
  wire [13:0] _T_59885; // @[Modules.scala 160:64:@5755.4]
  wire [13:0] buffer_1_486; // @[Modules.scala 160:64:@5756.4]
  wire [14:0] _T_59887; // @[Modules.scala 160:64:@5758.4]
  wire [13:0] _T_59888; // @[Modules.scala 160:64:@5759.4]
  wire [13:0] buffer_1_487; // @[Modules.scala 160:64:@5760.4]
  wire [14:0] _T_59890; // @[Modules.scala 160:64:@5762.4]
  wire [13:0] _T_59891; // @[Modules.scala 160:64:@5763.4]
  wire [13:0] buffer_1_488; // @[Modules.scala 160:64:@5764.4]
  wire [14:0] _T_59893; // @[Modules.scala 160:64:@5766.4]
  wire [13:0] _T_59894; // @[Modules.scala 160:64:@5767.4]
  wire [13:0] buffer_1_489; // @[Modules.scala 160:64:@5768.4]
  wire [14:0] _T_59896; // @[Modules.scala 160:64:@5770.4]
  wire [13:0] _T_59897; // @[Modules.scala 160:64:@5771.4]
  wire [13:0] buffer_1_490; // @[Modules.scala 160:64:@5772.4]
  wire [14:0] _T_59899; // @[Modules.scala 160:64:@5774.4]
  wire [13:0] _T_59900; // @[Modules.scala 160:64:@5775.4]
  wire [13:0] buffer_1_491; // @[Modules.scala 160:64:@5776.4]
  wire [14:0] _T_59902; // @[Modules.scala 160:64:@5778.4]
  wire [13:0] _T_59903; // @[Modules.scala 160:64:@5779.4]
  wire [13:0] buffer_1_492; // @[Modules.scala 160:64:@5780.4]
  wire [14:0] _T_59905; // @[Modules.scala 160:64:@5782.4]
  wire [13:0] _T_59906; // @[Modules.scala 160:64:@5783.4]
  wire [13:0] buffer_1_493; // @[Modules.scala 160:64:@5784.4]
  wire [14:0] _T_59908; // @[Modules.scala 160:64:@5786.4]
  wire [13:0] _T_59909; // @[Modules.scala 160:64:@5787.4]
  wire [13:0] buffer_1_494; // @[Modules.scala 160:64:@5788.4]
  wire [14:0] _T_59911; // @[Modules.scala 160:64:@5790.4]
  wire [13:0] _T_59912; // @[Modules.scala 160:64:@5791.4]
  wire [13:0] buffer_1_495; // @[Modules.scala 160:64:@5792.4]
  wire [14:0] _T_59914; // @[Modules.scala 160:64:@5794.4]
  wire [13:0] _T_59915; // @[Modules.scala 160:64:@5795.4]
  wire [13:0] buffer_1_496; // @[Modules.scala 160:64:@5796.4]
  wire [14:0] _T_59917; // @[Modules.scala 160:64:@5798.4]
  wire [13:0] _T_59918; // @[Modules.scala 160:64:@5799.4]
  wire [13:0] buffer_1_497; // @[Modules.scala 160:64:@5800.4]
  wire [14:0] _T_59920; // @[Modules.scala 160:64:@5802.4]
  wire [13:0] _T_59921; // @[Modules.scala 160:64:@5803.4]
  wire [13:0] buffer_1_498; // @[Modules.scala 160:64:@5804.4]
  wire [14:0] _T_59923; // @[Modules.scala 160:64:@5806.4]
  wire [13:0] _T_59924; // @[Modules.scala 160:64:@5807.4]
  wire [13:0] buffer_1_499; // @[Modules.scala 160:64:@5808.4]
  wire [14:0] _T_59926; // @[Modules.scala 160:64:@5810.4]
  wire [13:0] _T_59927; // @[Modules.scala 160:64:@5811.4]
  wire [13:0] buffer_1_500; // @[Modules.scala 160:64:@5812.4]
  wire [14:0] _T_59929; // @[Modules.scala 160:64:@5814.4]
  wire [13:0] _T_59930; // @[Modules.scala 160:64:@5815.4]
  wire [13:0] buffer_1_501; // @[Modules.scala 160:64:@5816.4]
  wire [14:0] _T_59932; // @[Modules.scala 160:64:@5818.4]
  wire [13:0] _T_59933; // @[Modules.scala 160:64:@5819.4]
  wire [13:0] buffer_1_502; // @[Modules.scala 160:64:@5820.4]
  wire [14:0] _T_59935; // @[Modules.scala 160:64:@5822.4]
  wire [13:0] _T_59936; // @[Modules.scala 160:64:@5823.4]
  wire [13:0] buffer_1_503; // @[Modules.scala 160:64:@5824.4]
  wire [14:0] _T_59938; // @[Modules.scala 160:64:@5826.4]
  wire [13:0] _T_59939; // @[Modules.scala 160:64:@5827.4]
  wire [13:0] buffer_1_504; // @[Modules.scala 160:64:@5828.4]
  wire [14:0] _T_59941; // @[Modules.scala 160:64:@5830.4]
  wire [13:0] _T_59942; // @[Modules.scala 160:64:@5831.4]
  wire [13:0] buffer_1_505; // @[Modules.scala 160:64:@5832.4]
  wire [14:0] _T_59944; // @[Modules.scala 160:64:@5834.4]
  wire [13:0] _T_59945; // @[Modules.scala 160:64:@5835.4]
  wire [13:0] buffer_1_506; // @[Modules.scala 160:64:@5836.4]
  wire [14:0] _T_59947; // @[Modules.scala 160:64:@5838.4]
  wire [13:0] _T_59948; // @[Modules.scala 160:64:@5839.4]
  wire [13:0] buffer_1_507; // @[Modules.scala 160:64:@5840.4]
  wire [14:0] _T_59950; // @[Modules.scala 160:64:@5842.4]
  wire [13:0] _T_59951; // @[Modules.scala 160:64:@5843.4]
  wire [13:0] buffer_1_508; // @[Modules.scala 160:64:@5844.4]
  wire [14:0] _T_59953; // @[Modules.scala 160:64:@5846.4]
  wire [13:0] _T_59954; // @[Modules.scala 160:64:@5847.4]
  wire [13:0] buffer_1_509; // @[Modules.scala 160:64:@5848.4]
  wire [14:0] _T_59956; // @[Modules.scala 160:64:@5850.4]
  wire [13:0] _T_59957; // @[Modules.scala 160:64:@5851.4]
  wire [13:0] buffer_1_510; // @[Modules.scala 160:64:@5852.4]
  wire [14:0] _T_59959; // @[Modules.scala 160:64:@5854.4]
  wire [13:0] _T_59960; // @[Modules.scala 160:64:@5855.4]
  wire [13:0] buffer_1_511; // @[Modules.scala 160:64:@5856.4]
  wire [14:0] _T_59962; // @[Modules.scala 160:64:@5858.4]
  wire [13:0] _T_59963; // @[Modules.scala 160:64:@5859.4]
  wire [13:0] buffer_1_512; // @[Modules.scala 160:64:@5860.4]
  wire [14:0] _T_59965; // @[Modules.scala 160:64:@5862.4]
  wire [13:0] _T_59966; // @[Modules.scala 160:64:@5863.4]
  wire [13:0] buffer_1_513; // @[Modules.scala 160:64:@5864.4]
  wire [14:0] _T_59968; // @[Modules.scala 160:64:@5866.4]
  wire [13:0] _T_59969; // @[Modules.scala 160:64:@5867.4]
  wire [13:0] buffer_1_514; // @[Modules.scala 160:64:@5868.4]
  wire [14:0] _T_59971; // @[Modules.scala 160:64:@5870.4]
  wire [13:0] _T_59972; // @[Modules.scala 160:64:@5871.4]
  wire [13:0] buffer_1_515; // @[Modules.scala 160:64:@5872.4]
  wire [14:0] _T_59974; // @[Modules.scala 160:64:@5874.4]
  wire [13:0] _T_59975; // @[Modules.scala 160:64:@5875.4]
  wire [13:0] buffer_1_516; // @[Modules.scala 160:64:@5876.4]
  wire [14:0] _T_59977; // @[Modules.scala 160:64:@5878.4]
  wire [13:0] _T_59978; // @[Modules.scala 160:64:@5879.4]
  wire [13:0] buffer_1_517; // @[Modules.scala 160:64:@5880.4]
  wire [14:0] _T_59980; // @[Modules.scala 160:64:@5882.4]
  wire [13:0] _T_59981; // @[Modules.scala 160:64:@5883.4]
  wire [13:0] buffer_1_518; // @[Modules.scala 160:64:@5884.4]
  wire [14:0] _T_59983; // @[Modules.scala 160:64:@5886.4]
  wire [13:0] _T_59984; // @[Modules.scala 160:64:@5887.4]
  wire [13:0] buffer_1_519; // @[Modules.scala 160:64:@5888.4]
  wire [14:0] _T_59986; // @[Modules.scala 160:64:@5890.4]
  wire [13:0] _T_59987; // @[Modules.scala 160:64:@5891.4]
  wire [13:0] buffer_1_520; // @[Modules.scala 160:64:@5892.4]
  wire [14:0] _T_59989; // @[Modules.scala 160:64:@5894.4]
  wire [13:0] _T_59990; // @[Modules.scala 160:64:@5895.4]
  wire [13:0] buffer_1_521; // @[Modules.scala 160:64:@5896.4]
  wire [14:0] _T_59992; // @[Modules.scala 160:64:@5898.4]
  wire [13:0] _T_59993; // @[Modules.scala 160:64:@5899.4]
  wire [13:0] buffer_1_522; // @[Modules.scala 160:64:@5900.4]
  wire [14:0] _T_59995; // @[Modules.scala 160:64:@5902.4]
  wire [13:0] _T_59996; // @[Modules.scala 160:64:@5903.4]
  wire [13:0] buffer_1_523; // @[Modules.scala 160:64:@5904.4]
  wire [14:0] _T_59998; // @[Modules.scala 160:64:@5906.4]
  wire [13:0] _T_59999; // @[Modules.scala 160:64:@5907.4]
  wire [13:0] buffer_1_524; // @[Modules.scala 160:64:@5908.4]
  wire [14:0] _T_60001; // @[Modules.scala 160:64:@5910.4]
  wire [13:0] _T_60002; // @[Modules.scala 160:64:@5911.4]
  wire [13:0] buffer_1_525; // @[Modules.scala 160:64:@5912.4]
  wire [14:0] _T_60004; // @[Modules.scala 160:64:@5914.4]
  wire [13:0] _T_60005; // @[Modules.scala 160:64:@5915.4]
  wire [13:0] buffer_1_526; // @[Modules.scala 160:64:@5916.4]
  wire [14:0] _T_60007; // @[Modules.scala 160:64:@5918.4]
  wire [13:0] _T_60008; // @[Modules.scala 160:64:@5919.4]
  wire [13:0] buffer_1_527; // @[Modules.scala 160:64:@5920.4]
  wire [14:0] _T_60010; // @[Modules.scala 160:64:@5922.4]
  wire [13:0] _T_60011; // @[Modules.scala 160:64:@5923.4]
  wire [13:0] buffer_1_528; // @[Modules.scala 160:64:@5924.4]
  wire [14:0] _T_60013; // @[Modules.scala 160:64:@5926.4]
  wire [13:0] _T_60014; // @[Modules.scala 160:64:@5927.4]
  wire [13:0] buffer_1_529; // @[Modules.scala 160:64:@5928.4]
  wire [14:0] _T_60016; // @[Modules.scala 160:64:@5930.4]
  wire [13:0] _T_60017; // @[Modules.scala 160:64:@5931.4]
  wire [13:0] buffer_1_530; // @[Modules.scala 160:64:@5932.4]
  wire [14:0] _T_60019; // @[Modules.scala 160:64:@5934.4]
  wire [13:0] _T_60020; // @[Modules.scala 160:64:@5935.4]
  wire [13:0] buffer_1_531; // @[Modules.scala 160:64:@5936.4]
  wire [14:0] _T_60022; // @[Modules.scala 160:64:@5938.4]
  wire [13:0] _T_60023; // @[Modules.scala 160:64:@5939.4]
  wire [13:0] buffer_1_532; // @[Modules.scala 160:64:@5940.4]
  wire [14:0] _T_60025; // @[Modules.scala 160:64:@5942.4]
  wire [13:0] _T_60026; // @[Modules.scala 160:64:@5943.4]
  wire [13:0] buffer_1_533; // @[Modules.scala 160:64:@5944.4]
  wire [14:0] _T_60028; // @[Modules.scala 160:64:@5946.4]
  wire [13:0] _T_60029; // @[Modules.scala 160:64:@5947.4]
  wire [13:0] buffer_1_534; // @[Modules.scala 160:64:@5948.4]
  wire [14:0] _T_60031; // @[Modules.scala 160:64:@5950.4]
  wire [13:0] _T_60032; // @[Modules.scala 160:64:@5951.4]
  wire [13:0] buffer_1_535; // @[Modules.scala 160:64:@5952.4]
  wire [14:0] _T_60034; // @[Modules.scala 160:64:@5954.4]
  wire [13:0] _T_60035; // @[Modules.scala 160:64:@5955.4]
  wire [13:0] buffer_1_536; // @[Modules.scala 160:64:@5956.4]
  wire [14:0] _T_60037; // @[Modules.scala 160:64:@5958.4]
  wire [13:0] _T_60038; // @[Modules.scala 160:64:@5959.4]
  wire [13:0] buffer_1_537; // @[Modules.scala 160:64:@5960.4]
  wire [14:0] _T_60040; // @[Modules.scala 160:64:@5962.4]
  wire [13:0] _T_60041; // @[Modules.scala 160:64:@5963.4]
  wire [13:0] buffer_1_538; // @[Modules.scala 160:64:@5964.4]
  wire [14:0] _T_60043; // @[Modules.scala 160:64:@5966.4]
  wire [13:0] _T_60044; // @[Modules.scala 160:64:@5967.4]
  wire [13:0] buffer_1_539; // @[Modules.scala 160:64:@5968.4]
  wire [14:0] _T_60046; // @[Modules.scala 160:64:@5970.4]
  wire [13:0] _T_60047; // @[Modules.scala 160:64:@5971.4]
  wire [13:0] buffer_1_540; // @[Modules.scala 160:64:@5972.4]
  wire [14:0] _T_60049; // @[Modules.scala 160:64:@5974.4]
  wire [13:0] _T_60050; // @[Modules.scala 160:64:@5975.4]
  wire [13:0] buffer_1_541; // @[Modules.scala 160:64:@5976.4]
  wire [14:0] _T_60052; // @[Modules.scala 160:64:@5978.4]
  wire [13:0] _T_60053; // @[Modules.scala 160:64:@5979.4]
  wire [13:0] buffer_1_542; // @[Modules.scala 160:64:@5980.4]
  wire [14:0] _T_60055; // @[Modules.scala 160:64:@5982.4]
  wire [13:0] _T_60056; // @[Modules.scala 160:64:@5983.4]
  wire [13:0] buffer_1_543; // @[Modules.scala 160:64:@5984.4]
  wire [14:0] _T_60058; // @[Modules.scala 160:64:@5986.4]
  wire [13:0] _T_60059; // @[Modules.scala 160:64:@5987.4]
  wire [13:0] buffer_1_544; // @[Modules.scala 160:64:@5988.4]
  wire [14:0] _T_60061; // @[Modules.scala 160:64:@5990.4]
  wire [13:0] _T_60062; // @[Modules.scala 160:64:@5991.4]
  wire [13:0] buffer_1_545; // @[Modules.scala 160:64:@5992.4]
  wire [14:0] _T_60064; // @[Modules.scala 160:64:@5994.4]
  wire [13:0] _T_60065; // @[Modules.scala 160:64:@5995.4]
  wire [13:0] buffer_1_546; // @[Modules.scala 160:64:@5996.4]
  wire [14:0] _T_60067; // @[Modules.scala 160:64:@5998.4]
  wire [13:0] _T_60068; // @[Modules.scala 160:64:@5999.4]
  wire [13:0] buffer_1_547; // @[Modules.scala 160:64:@6000.4]
  wire [14:0] _T_60070; // @[Modules.scala 160:64:@6002.4]
  wire [13:0] _T_60071; // @[Modules.scala 160:64:@6003.4]
  wire [13:0] buffer_1_548; // @[Modules.scala 160:64:@6004.4]
  wire [14:0] _T_60073; // @[Modules.scala 160:64:@6006.4]
  wire [13:0] _T_60074; // @[Modules.scala 160:64:@6007.4]
  wire [13:0] buffer_1_549; // @[Modules.scala 160:64:@6008.4]
  wire [14:0] _T_60076; // @[Modules.scala 160:64:@6010.4]
  wire [13:0] _T_60077; // @[Modules.scala 160:64:@6011.4]
  wire [13:0] buffer_1_550; // @[Modules.scala 160:64:@6012.4]
  wire [14:0] _T_60079; // @[Modules.scala 160:64:@6014.4]
  wire [13:0] _T_60080; // @[Modules.scala 160:64:@6015.4]
  wire [13:0] buffer_1_551; // @[Modules.scala 160:64:@6016.4]
  wire [14:0] _T_60082; // @[Modules.scala 160:64:@6018.4]
  wire [13:0] _T_60083; // @[Modules.scala 160:64:@6019.4]
  wire [13:0] buffer_1_552; // @[Modules.scala 160:64:@6020.4]
  wire [14:0] _T_60085; // @[Modules.scala 160:64:@6022.4]
  wire [13:0] _T_60086; // @[Modules.scala 160:64:@6023.4]
  wire [13:0] buffer_1_553; // @[Modules.scala 160:64:@6024.4]
  wire [14:0] _T_60088; // @[Modules.scala 160:64:@6026.4]
  wire [13:0] _T_60089; // @[Modules.scala 160:64:@6027.4]
  wire [13:0] buffer_1_554; // @[Modules.scala 160:64:@6028.4]
  wire [14:0] _T_60091; // @[Modules.scala 160:64:@6030.4]
  wire [13:0] _T_60092; // @[Modules.scala 160:64:@6031.4]
  wire [13:0] buffer_1_555; // @[Modules.scala 160:64:@6032.4]
  wire [14:0] _T_60094; // @[Modules.scala 160:64:@6034.4]
  wire [13:0] _T_60095; // @[Modules.scala 160:64:@6035.4]
  wire [13:0] buffer_1_556; // @[Modules.scala 160:64:@6036.4]
  wire [14:0] _T_60097; // @[Modules.scala 160:64:@6038.4]
  wire [13:0] _T_60098; // @[Modules.scala 160:64:@6039.4]
  wire [13:0] buffer_1_557; // @[Modules.scala 160:64:@6040.4]
  wire [14:0] _T_60100; // @[Modules.scala 160:64:@6042.4]
  wire [13:0] _T_60101; // @[Modules.scala 160:64:@6043.4]
  wire [13:0] buffer_1_558; // @[Modules.scala 160:64:@6044.4]
  wire [14:0] _T_60103; // @[Modules.scala 160:64:@6046.4]
  wire [13:0] _T_60104; // @[Modules.scala 160:64:@6047.4]
  wire [13:0] buffer_1_559; // @[Modules.scala 160:64:@6048.4]
  wire [14:0] _T_60106; // @[Modules.scala 160:64:@6050.4]
  wire [13:0] _T_60107; // @[Modules.scala 160:64:@6051.4]
  wire [13:0] buffer_1_560; // @[Modules.scala 160:64:@6052.4]
  wire [14:0] _T_60109; // @[Modules.scala 160:64:@6054.4]
  wire [13:0] _T_60110; // @[Modules.scala 160:64:@6055.4]
  wire [13:0] buffer_1_561; // @[Modules.scala 160:64:@6056.4]
  wire [14:0] _T_60112; // @[Modules.scala 160:64:@6058.4]
  wire [13:0] _T_60113; // @[Modules.scala 160:64:@6059.4]
  wire [13:0] buffer_1_562; // @[Modules.scala 160:64:@6060.4]
  wire [14:0] _T_60115; // @[Modules.scala 160:64:@6062.4]
  wire [13:0] _T_60116; // @[Modules.scala 160:64:@6063.4]
  wire [13:0] buffer_1_563; // @[Modules.scala 160:64:@6064.4]
  wire [14:0] _T_60118; // @[Modules.scala 160:64:@6066.4]
  wire [13:0] _T_60119; // @[Modules.scala 160:64:@6067.4]
  wire [13:0] buffer_1_564; // @[Modules.scala 160:64:@6068.4]
  wire [14:0] _T_60121; // @[Modules.scala 160:64:@6070.4]
  wire [13:0] _T_60122; // @[Modules.scala 160:64:@6071.4]
  wire [13:0] buffer_1_565; // @[Modules.scala 160:64:@6072.4]
  wire [14:0] _T_60124; // @[Modules.scala 160:64:@6074.4]
  wire [13:0] _T_60125; // @[Modules.scala 160:64:@6075.4]
  wire [13:0] buffer_1_566; // @[Modules.scala 160:64:@6076.4]
  wire [14:0] _T_60127; // @[Modules.scala 160:64:@6078.4]
  wire [13:0] _T_60128; // @[Modules.scala 160:64:@6079.4]
  wire [13:0] buffer_1_567; // @[Modules.scala 160:64:@6080.4]
  wire [14:0] _T_60130; // @[Modules.scala 160:64:@6082.4]
  wire [13:0] _T_60131; // @[Modules.scala 160:64:@6083.4]
  wire [13:0] buffer_1_568; // @[Modules.scala 160:64:@6084.4]
  wire [14:0] _T_60133; // @[Modules.scala 160:64:@6086.4]
  wire [13:0] _T_60134; // @[Modules.scala 160:64:@6087.4]
  wire [13:0] buffer_1_569; // @[Modules.scala 160:64:@6088.4]
  wire [14:0] _T_60136; // @[Modules.scala 160:64:@6090.4]
  wire [13:0] _T_60137; // @[Modules.scala 160:64:@6091.4]
  wire [13:0] buffer_1_570; // @[Modules.scala 160:64:@6092.4]
  wire [14:0] _T_60139; // @[Modules.scala 160:64:@6094.4]
  wire [13:0] _T_60140; // @[Modules.scala 160:64:@6095.4]
  wire [13:0] buffer_1_571; // @[Modules.scala 160:64:@6096.4]
  wire [14:0] _T_60142; // @[Modules.scala 160:64:@6098.4]
  wire [13:0] _T_60143; // @[Modules.scala 160:64:@6099.4]
  wire [13:0] buffer_1_572; // @[Modules.scala 160:64:@6100.4]
  wire [14:0] _T_60145; // @[Modules.scala 160:64:@6102.4]
  wire [13:0] _T_60146; // @[Modules.scala 160:64:@6103.4]
  wire [13:0] buffer_1_573; // @[Modules.scala 160:64:@6104.4]
  wire [14:0] _T_60148; // @[Modules.scala 160:64:@6106.4]
  wire [13:0] _T_60149; // @[Modules.scala 160:64:@6107.4]
  wire [13:0] buffer_1_574; // @[Modules.scala 160:64:@6108.4]
  wire [14:0] _T_60151; // @[Modules.scala 160:64:@6110.4]
  wire [13:0] _T_60152; // @[Modules.scala 160:64:@6111.4]
  wire [13:0] buffer_1_575; // @[Modules.scala 160:64:@6112.4]
  wire [14:0] _T_60154; // @[Modules.scala 160:64:@6114.4]
  wire [13:0] _T_60155; // @[Modules.scala 160:64:@6115.4]
  wire [13:0] buffer_1_576; // @[Modules.scala 160:64:@6116.4]
  wire [14:0] _T_60157; // @[Modules.scala 160:64:@6118.4]
  wire [13:0] _T_60158; // @[Modules.scala 160:64:@6119.4]
  wire [13:0] buffer_1_577; // @[Modules.scala 160:64:@6120.4]
  wire [14:0] _T_60160; // @[Modules.scala 160:64:@6122.4]
  wire [13:0] _T_60161; // @[Modules.scala 160:64:@6123.4]
  wire [13:0] buffer_1_578; // @[Modules.scala 160:64:@6124.4]
  wire [14:0] _T_60163; // @[Modules.scala 160:64:@6126.4]
  wire [13:0] _T_60164; // @[Modules.scala 160:64:@6127.4]
  wire [13:0] buffer_1_579; // @[Modules.scala 160:64:@6128.4]
  wire [14:0] _T_60166; // @[Modules.scala 160:64:@6130.4]
  wire [13:0] _T_60167; // @[Modules.scala 160:64:@6131.4]
  wire [13:0] buffer_1_580; // @[Modules.scala 160:64:@6132.4]
  wire [14:0] _T_60169; // @[Modules.scala 160:64:@6134.4]
  wire [13:0] _T_60170; // @[Modules.scala 160:64:@6135.4]
  wire [13:0] buffer_1_581; // @[Modules.scala 160:64:@6136.4]
  wire [14:0] _T_60172; // @[Modules.scala 160:64:@6138.4]
  wire [13:0] _T_60173; // @[Modules.scala 160:64:@6139.4]
  wire [13:0] buffer_1_582; // @[Modules.scala 160:64:@6140.4]
  wire [14:0] _T_60175; // @[Modules.scala 160:64:@6142.4]
  wire [13:0] _T_60176; // @[Modules.scala 160:64:@6143.4]
  wire [13:0] buffer_1_583; // @[Modules.scala 160:64:@6144.4]
  wire [14:0] _T_60178; // @[Modules.scala 160:64:@6146.4]
  wire [13:0] _T_60179; // @[Modules.scala 160:64:@6147.4]
  wire [13:0] buffer_1_584; // @[Modules.scala 160:64:@6148.4]
  wire [14:0] _T_60181; // @[Modules.scala 160:64:@6150.4]
  wire [13:0] _T_60182; // @[Modules.scala 160:64:@6151.4]
  wire [13:0] buffer_1_585; // @[Modules.scala 160:64:@6152.4]
  wire [14:0] _T_60184; // @[Modules.scala 160:64:@6154.4]
  wire [13:0] _T_60185; // @[Modules.scala 160:64:@6155.4]
  wire [13:0] buffer_1_586; // @[Modules.scala 160:64:@6156.4]
  wire [14:0] _T_60187; // @[Modules.scala 160:64:@6158.4]
  wire [13:0] _T_60188; // @[Modules.scala 160:64:@6159.4]
  wire [13:0] buffer_1_587; // @[Modules.scala 160:64:@6160.4]
  wire [14:0] _T_60190; // @[Modules.scala 160:64:@6162.4]
  wire [13:0] _T_60191; // @[Modules.scala 160:64:@6163.4]
  wire [13:0] buffer_1_588; // @[Modules.scala 160:64:@6164.4]
  wire [14:0] _T_60193; // @[Modules.scala 166:64:@6166.4]
  wire [13:0] _T_60194; // @[Modules.scala 166:64:@6167.4]
  wire [13:0] buffer_1_589; // @[Modules.scala 166:64:@6168.4]
  wire [14:0] _T_60196; // @[Modules.scala 166:64:@6170.4]
  wire [13:0] _T_60197; // @[Modules.scala 166:64:@6171.4]
  wire [13:0] buffer_1_590; // @[Modules.scala 166:64:@6172.4]
  wire [14:0] _T_60199; // @[Modules.scala 166:64:@6174.4]
  wire [13:0] _T_60200; // @[Modules.scala 166:64:@6175.4]
  wire [13:0] buffer_1_591; // @[Modules.scala 166:64:@6176.4]
  wire [14:0] _T_60202; // @[Modules.scala 166:64:@6178.4]
  wire [13:0] _T_60203; // @[Modules.scala 166:64:@6179.4]
  wire [13:0] buffer_1_592; // @[Modules.scala 166:64:@6180.4]
  wire [14:0] _T_60205; // @[Modules.scala 166:64:@6182.4]
  wire [13:0] _T_60206; // @[Modules.scala 166:64:@6183.4]
  wire [13:0] buffer_1_593; // @[Modules.scala 166:64:@6184.4]
  wire [14:0] _T_60208; // @[Modules.scala 166:64:@6186.4]
  wire [13:0] _T_60209; // @[Modules.scala 166:64:@6187.4]
  wire [13:0] buffer_1_594; // @[Modules.scala 166:64:@6188.4]
  wire [14:0] _T_60211; // @[Modules.scala 166:64:@6190.4]
  wire [13:0] _T_60212; // @[Modules.scala 166:64:@6191.4]
  wire [13:0] buffer_1_595; // @[Modules.scala 166:64:@6192.4]
  wire [14:0] _T_60214; // @[Modules.scala 166:64:@6194.4]
  wire [13:0] _T_60215; // @[Modules.scala 166:64:@6195.4]
  wire [13:0] buffer_1_596; // @[Modules.scala 166:64:@6196.4]
  wire [14:0] _T_60217; // @[Modules.scala 166:64:@6198.4]
  wire [13:0] _T_60218; // @[Modules.scala 166:64:@6199.4]
  wire [13:0] buffer_1_597; // @[Modules.scala 166:64:@6200.4]
  wire [14:0] _T_60220; // @[Modules.scala 166:64:@6202.4]
  wire [13:0] _T_60221; // @[Modules.scala 166:64:@6203.4]
  wire [13:0] buffer_1_598; // @[Modules.scala 166:64:@6204.4]
  wire [14:0] _T_60223; // @[Modules.scala 166:64:@6206.4]
  wire [13:0] _T_60224; // @[Modules.scala 166:64:@6207.4]
  wire [13:0] buffer_1_599; // @[Modules.scala 166:64:@6208.4]
  wire [14:0] _T_60226; // @[Modules.scala 166:64:@6210.4]
  wire [13:0] _T_60227; // @[Modules.scala 166:64:@6211.4]
  wire [13:0] buffer_1_600; // @[Modules.scala 166:64:@6212.4]
  wire [14:0] _T_60229; // @[Modules.scala 166:64:@6214.4]
  wire [13:0] _T_60230; // @[Modules.scala 166:64:@6215.4]
  wire [13:0] buffer_1_601; // @[Modules.scala 166:64:@6216.4]
  wire [14:0] _T_60232; // @[Modules.scala 172:66:@6218.4]
  wire [13:0] _T_60233; // @[Modules.scala 172:66:@6219.4]
  wire [13:0] buffer_1_602; // @[Modules.scala 172:66:@6220.4]
  wire [14:0] _T_60235; // @[Modules.scala 166:64:@6222.4]
  wire [13:0] _T_60236; // @[Modules.scala 166:64:@6223.4]
  wire [13:0] buffer_1_603; // @[Modules.scala 166:64:@6224.4]
  wire [14:0] _T_60238; // @[Modules.scala 166:64:@6226.4]
  wire [13:0] _T_60239; // @[Modules.scala 166:64:@6227.4]
  wire [13:0] buffer_1_604; // @[Modules.scala 166:64:@6228.4]
  wire [14:0] _T_60241; // @[Modules.scala 160:64:@6230.4]
  wire [13:0] _T_60242; // @[Modules.scala 160:64:@6231.4]
  wire [13:0] buffer_1_605; // @[Modules.scala 160:64:@6232.4]
  wire [14:0] _T_60244; // @[Modules.scala 172:66:@6234.4]
  wire [13:0] _T_60245; // @[Modules.scala 172:66:@6235.4]
  wire [13:0] buffer_1_606; // @[Modules.scala 172:66:@6236.4]
  wire [4:0] _T_60248; // @[Modules.scala 143:74:@6415.4]
  wire [4:0] _T_60250; // @[Modules.scala 144:80:@6416.4]
  wire [5:0] _T_60251; // @[Modules.scala 143:103:@6417.4]
  wire [4:0] _T_60252; // @[Modules.scala 143:103:@6418.4]
  wire [4:0] _T_60253; // @[Modules.scala 143:103:@6419.4]
  wire [4:0] _T_60255; // @[Modules.scala 143:74:@6421.4]
  wire [4:0] _T_60257; // @[Modules.scala 144:80:@6422.4]
  wire [5:0] _T_60258; // @[Modules.scala 143:103:@6423.4]
  wire [4:0] _T_60259; // @[Modules.scala 143:103:@6424.4]
  wire [4:0] _T_60260; // @[Modules.scala 143:103:@6425.4]
  wire [4:0] _T_60264; // @[Modules.scala 144:80:@6428.4]
  wire [5:0] _T_60265; // @[Modules.scala 143:103:@6429.4]
  wire [4:0] _T_60266; // @[Modules.scala 143:103:@6430.4]
  wire [4:0] _T_60267; // @[Modules.scala 143:103:@6431.4]
  wire [4:0] _T_60269; // @[Modules.scala 143:74:@6433.4]
  wire [4:0] _T_60271; // @[Modules.scala 144:80:@6434.4]
  wire [5:0] _T_60272; // @[Modules.scala 143:103:@6435.4]
  wire [4:0] _T_60273; // @[Modules.scala 143:103:@6436.4]
  wire [4:0] _T_60274; // @[Modules.scala 143:103:@6437.4]
  wire [6:0] _T_60279; // @[Modules.scala 143:103:@6441.4]
  wire [5:0] _T_60280; // @[Modules.scala 143:103:@6442.4]
  wire [5:0] _T_60281; // @[Modules.scala 143:103:@6443.4]
  wire [6:0] _T_60286; // @[Modules.scala 143:103:@6447.4]
  wire [5:0] _T_60287; // @[Modules.scala 143:103:@6448.4]
  wire [5:0] _T_60288; // @[Modules.scala 143:103:@6449.4]
  wire [5:0] _T_60293; // @[Modules.scala 143:103:@6453.4]
  wire [4:0] _T_60294; // @[Modules.scala 143:103:@6454.4]
  wire [4:0] _T_60295; // @[Modules.scala 143:103:@6455.4]
  wire [4:0] _T_60299; // @[Modules.scala 144:80:@6458.4]
  wire [5:0] _GEN_144; // @[Modules.scala 143:103:@6459.4]
  wire [6:0] _T_60300; // @[Modules.scala 143:103:@6459.4]
  wire [5:0] _T_60301; // @[Modules.scala 143:103:@6460.4]
  wire [5:0] _T_60302; // @[Modules.scala 143:103:@6461.4]
  wire [5:0] _T_60307; // @[Modules.scala 143:103:@6465.4]
  wire [4:0] _T_60308; // @[Modules.scala 143:103:@6466.4]
  wire [4:0] _T_60309; // @[Modules.scala 143:103:@6467.4]
  wire [4:0] _T_60327; // @[Modules.scala 144:80:@6482.4]
  wire [5:0] _T_60328; // @[Modules.scala 143:103:@6483.4]
  wire [4:0] _T_60329; // @[Modules.scala 143:103:@6484.4]
  wire [4:0] _T_60330; // @[Modules.scala 143:103:@6485.4]
  wire [4:0] _T_60332; // @[Modules.scala 143:74:@6487.4]
  wire [4:0] _T_60334; // @[Modules.scala 144:80:@6488.4]
  wire [5:0] _T_60335; // @[Modules.scala 143:103:@6489.4]
  wire [4:0] _T_60336; // @[Modules.scala 143:103:@6490.4]
  wire [4:0] _T_60337; // @[Modules.scala 143:103:@6491.4]
  wire [5:0] _T_60342; // @[Modules.scala 143:103:@6495.4]
  wire [4:0] _T_60343; // @[Modules.scala 143:103:@6496.4]
  wire [4:0] _T_60344; // @[Modules.scala 143:103:@6497.4]
  wire [5:0] _T_60349; // @[Modules.scala 143:103:@6501.4]
  wire [4:0] _T_60350; // @[Modules.scala 143:103:@6502.4]
  wire [4:0] _T_60351; // @[Modules.scala 143:103:@6503.4]
  wire [5:0] _T_60356; // @[Modules.scala 143:103:@6507.4]
  wire [4:0] _T_60357; // @[Modules.scala 143:103:@6508.4]
  wire [4:0] _T_60358; // @[Modules.scala 143:103:@6509.4]
  wire [5:0] _T_60363; // @[Modules.scala 143:103:@6513.4]
  wire [4:0] _T_60364; // @[Modules.scala 143:103:@6514.4]
  wire [4:0] _T_60365; // @[Modules.scala 143:103:@6515.4]
  wire [5:0] _GEN_145; // @[Modules.scala 143:103:@6519.4]
  wire [6:0] _T_60370; // @[Modules.scala 143:103:@6519.4]
  wire [5:0] _T_60371; // @[Modules.scala 143:103:@6520.4]
  wire [5:0] _T_60372; // @[Modules.scala 143:103:@6521.4]
  wire [4:0] _T_60402; // @[Modules.scala 143:74:@6547.4]
  wire [4:0] _T_60404; // @[Modules.scala 144:80:@6548.4]
  wire [5:0] _T_60405; // @[Modules.scala 143:103:@6549.4]
  wire [4:0] _T_60406; // @[Modules.scala 143:103:@6550.4]
  wire [4:0] _T_60407; // @[Modules.scala 143:103:@6551.4]
  wire [6:0] _T_60412; // @[Modules.scala 143:103:@6555.4]
  wire [5:0] _T_60413; // @[Modules.scala 143:103:@6556.4]
  wire [5:0] _T_60414; // @[Modules.scala 143:103:@6557.4]
  wire [5:0] _GEN_147; // @[Modules.scala 143:103:@6561.4]
  wire [6:0] _T_60419; // @[Modules.scala 143:103:@6561.4]
  wire [5:0] _T_60420; // @[Modules.scala 143:103:@6562.4]
  wire [5:0] _T_60421; // @[Modules.scala 143:103:@6563.4]
  wire [4:0] _T_60430; // @[Modules.scala 143:74:@6571.4]
  wire [5:0] _GEN_148; // @[Modules.scala 143:103:@6573.4]
  wire [6:0] _T_60433; // @[Modules.scala 143:103:@6573.4]
  wire [5:0] _T_60434; // @[Modules.scala 143:103:@6574.4]
  wire [5:0] _T_60435; // @[Modules.scala 143:103:@6575.4]
  wire [6:0] _T_60440; // @[Modules.scala 143:103:@6579.4]
  wire [5:0] _T_60441; // @[Modules.scala 143:103:@6580.4]
  wire [5:0] _T_60442; // @[Modules.scala 143:103:@6581.4]
  wire [6:0] _T_60447; // @[Modules.scala 143:103:@6585.4]
  wire [5:0] _T_60448; // @[Modules.scala 143:103:@6586.4]
  wire [5:0] _T_60449; // @[Modules.scala 143:103:@6587.4]
  wire [6:0] _T_60454; // @[Modules.scala 143:103:@6591.4]
  wire [5:0] _T_60455; // @[Modules.scala 143:103:@6592.4]
  wire [5:0] _T_60456; // @[Modules.scala 143:103:@6593.4]
  wire [6:0] _T_60461; // @[Modules.scala 143:103:@6597.4]
  wire [5:0] _T_60462; // @[Modules.scala 143:103:@6598.4]
  wire [5:0] _T_60463; // @[Modules.scala 143:103:@6599.4]
  wire [6:0] _T_60468; // @[Modules.scala 143:103:@6603.4]
  wire [5:0] _T_60469; // @[Modules.scala 143:103:@6604.4]
  wire [5:0] _T_60470; // @[Modules.scala 143:103:@6605.4]
  wire [4:0] _T_60474; // @[Modules.scala 144:80:@6608.4]
  wire [5:0] _T_60475; // @[Modules.scala 143:103:@6609.4]
  wire [4:0] _T_60476; // @[Modules.scala 143:103:@6610.4]
  wire [4:0] _T_60477; // @[Modules.scala 143:103:@6611.4]
  wire [6:0] _T_60482; // @[Modules.scala 143:103:@6615.4]
  wire [5:0] _T_60483; // @[Modules.scala 143:103:@6616.4]
  wire [5:0] _T_60484; // @[Modules.scala 143:103:@6617.4]
  wire [5:0] _T_60488; // @[Modules.scala 144:80:@6620.4]
  wire [6:0] _T_60489; // @[Modules.scala 143:103:@6621.4]
  wire [5:0] _T_60490; // @[Modules.scala 143:103:@6622.4]
  wire [5:0] _T_60491; // @[Modules.scala 143:103:@6623.4]
  wire [4:0] _T_60495; // @[Modules.scala 144:80:@6626.4]
  wire [5:0] _GEN_150; // @[Modules.scala 143:103:@6627.4]
  wire [6:0] _T_60496; // @[Modules.scala 143:103:@6627.4]
  wire [5:0] _T_60497; // @[Modules.scala 143:103:@6628.4]
  wire [5:0] _T_60498; // @[Modules.scala 143:103:@6629.4]
  wire [4:0] _T_60500; // @[Modules.scala 143:74:@6631.4]
  wire [4:0] _T_60502; // @[Modules.scala 144:80:@6632.4]
  wire [5:0] _T_60503; // @[Modules.scala 143:103:@6633.4]
  wire [4:0] _T_60504; // @[Modules.scala 143:103:@6634.4]
  wire [4:0] _T_60505; // @[Modules.scala 143:103:@6635.4]
  wire [4:0] _T_60507; // @[Modules.scala 143:74:@6637.4]
  wire [4:0] _T_60509; // @[Modules.scala 144:80:@6638.4]
  wire [5:0] _T_60510; // @[Modules.scala 143:103:@6639.4]
  wire [4:0] _T_60511; // @[Modules.scala 143:103:@6640.4]
  wire [4:0] _T_60512; // @[Modules.scala 143:103:@6641.4]
  wire [4:0] _T_60514; // @[Modules.scala 143:74:@6643.4]
  wire [5:0] _GEN_151; // @[Modules.scala 143:103:@6645.4]
  wire [6:0] _T_60517; // @[Modules.scala 143:103:@6645.4]
  wire [5:0] _T_60518; // @[Modules.scala 143:103:@6646.4]
  wire [5:0] _T_60519; // @[Modules.scala 143:103:@6647.4]
  wire [4:0] _T_60544; // @[Modules.scala 144:80:@6668.4]
  wire [5:0] _GEN_152; // @[Modules.scala 143:103:@6669.4]
  wire [6:0] _T_60545; // @[Modules.scala 143:103:@6669.4]
  wire [5:0] _T_60546; // @[Modules.scala 143:103:@6670.4]
  wire [5:0] _T_60547; // @[Modules.scala 143:103:@6671.4]
  wire [5:0] _T_60549; // @[Modules.scala 143:74:@6673.4]
  wire [4:0] _T_60551; // @[Modules.scala 144:80:@6674.4]
  wire [5:0] _GEN_153; // @[Modules.scala 143:103:@6675.4]
  wire [6:0] _T_60552; // @[Modules.scala 143:103:@6675.4]
  wire [5:0] _T_60553; // @[Modules.scala 143:103:@6676.4]
  wire [5:0] _T_60554; // @[Modules.scala 143:103:@6677.4]
  wire [4:0] _T_60556; // @[Modules.scala 143:74:@6679.4]
  wire [5:0] _GEN_154; // @[Modules.scala 143:103:@6681.4]
  wire [6:0] _T_60559; // @[Modules.scala 143:103:@6681.4]
  wire [5:0] _T_60560; // @[Modules.scala 143:103:@6682.4]
  wire [5:0] _T_60561; // @[Modules.scala 143:103:@6683.4]
  wire [4:0] _T_60563; // @[Modules.scala 143:74:@6685.4]
  wire [5:0] _T_60566; // @[Modules.scala 143:103:@6687.4]
  wire [4:0] _T_60567; // @[Modules.scala 143:103:@6688.4]
  wire [4:0] _T_60568; // @[Modules.scala 143:103:@6689.4]
  wire [6:0] _T_60573; // @[Modules.scala 143:103:@6693.4]
  wire [5:0] _T_60574; // @[Modules.scala 143:103:@6694.4]
  wire [5:0] _T_60575; // @[Modules.scala 143:103:@6695.4]
  wire [4:0] _T_60577; // @[Modules.scala 143:74:@6697.4]
  wire [4:0] _T_60579; // @[Modules.scala 144:80:@6698.4]
  wire [5:0] _T_60580; // @[Modules.scala 143:103:@6699.4]
  wire [4:0] _T_60581; // @[Modules.scala 143:103:@6700.4]
  wire [4:0] _T_60582; // @[Modules.scala 143:103:@6701.4]
  wire [4:0] _T_60584; // @[Modules.scala 143:74:@6703.4]
  wire [4:0] _T_60586; // @[Modules.scala 144:80:@6704.4]
  wire [5:0] _T_60587; // @[Modules.scala 143:103:@6705.4]
  wire [4:0] _T_60588; // @[Modules.scala 143:103:@6706.4]
  wire [4:0] _T_60589; // @[Modules.scala 143:103:@6707.4]
  wire [5:0] _T_60605; // @[Modules.scala 143:74:@6721.4]
  wire [4:0] _T_60607; // @[Modules.scala 144:80:@6722.4]
  wire [5:0] _GEN_155; // @[Modules.scala 143:103:@6723.4]
  wire [6:0] _T_60608; // @[Modules.scala 143:103:@6723.4]
  wire [5:0] _T_60609; // @[Modules.scala 143:103:@6724.4]
  wire [5:0] _T_60610; // @[Modules.scala 143:103:@6725.4]
  wire [5:0] _T_60614; // @[Modules.scala 144:80:@6728.4]
  wire [6:0] _T_60615; // @[Modules.scala 143:103:@6729.4]
  wire [5:0] _T_60616; // @[Modules.scala 143:103:@6730.4]
  wire [5:0] _T_60617; // @[Modules.scala 143:103:@6731.4]
  wire [5:0] _T_60619; // @[Modules.scala 143:74:@6733.4]
  wire [6:0] _T_60622; // @[Modules.scala 143:103:@6735.4]
  wire [5:0] _T_60623; // @[Modules.scala 143:103:@6736.4]
  wire [5:0] _T_60624; // @[Modules.scala 143:103:@6737.4]
  wire [5:0] _T_60628; // @[Modules.scala 144:80:@6740.4]
  wire [6:0] _T_60629; // @[Modules.scala 143:103:@6741.4]
  wire [5:0] _T_60630; // @[Modules.scala 143:103:@6742.4]
  wire [5:0] _T_60631; // @[Modules.scala 143:103:@6743.4]
  wire [5:0] _T_60633; // @[Modules.scala 143:74:@6745.4]
  wire [4:0] _T_60635; // @[Modules.scala 144:80:@6746.4]
  wire [5:0] _GEN_159; // @[Modules.scala 143:103:@6747.4]
  wire [6:0] _T_60636; // @[Modules.scala 143:103:@6747.4]
  wire [5:0] _T_60637; // @[Modules.scala 143:103:@6748.4]
  wire [5:0] _T_60638; // @[Modules.scala 143:103:@6749.4]
  wire [4:0] _T_60642; // @[Modules.scala 144:80:@6752.4]
  wire [5:0] _GEN_160; // @[Modules.scala 143:103:@6753.4]
  wire [6:0] _T_60643; // @[Modules.scala 143:103:@6753.4]
  wire [5:0] _T_60644; // @[Modules.scala 143:103:@6754.4]
  wire [5:0] _T_60645; // @[Modules.scala 143:103:@6755.4]
  wire [4:0] _T_60647; // @[Modules.scala 143:74:@6757.4]
  wire [5:0] _GEN_161; // @[Modules.scala 143:103:@6759.4]
  wire [6:0] _T_60650; // @[Modules.scala 143:103:@6759.4]
  wire [5:0] _T_60651; // @[Modules.scala 143:103:@6760.4]
  wire [5:0] _T_60652; // @[Modules.scala 143:103:@6761.4]
  wire [4:0] _T_60656; // @[Modules.scala 144:80:@6764.4]
  wire [5:0] _T_60657; // @[Modules.scala 143:103:@6765.4]
  wire [4:0] _T_60658; // @[Modules.scala 143:103:@6766.4]
  wire [4:0] _T_60659; // @[Modules.scala 143:103:@6767.4]
  wire [4:0] _T_60668; // @[Modules.scala 143:74:@6775.4]
  wire [5:0] _T_60671; // @[Modules.scala 143:103:@6777.4]
  wire [4:0] _T_60672; // @[Modules.scala 143:103:@6778.4]
  wire [4:0] _T_60673; // @[Modules.scala 143:103:@6779.4]
  wire [5:0] _T_60678; // @[Modules.scala 143:103:@6783.4]
  wire [4:0] _T_60679; // @[Modules.scala 143:103:@6784.4]
  wire [4:0] _T_60680; // @[Modules.scala 143:103:@6785.4]
  wire [4:0] _T_60689; // @[Modules.scala 143:74:@6793.4]
  wire [4:0] _T_60691; // @[Modules.scala 144:80:@6794.4]
  wire [5:0] _T_60692; // @[Modules.scala 143:103:@6795.4]
  wire [4:0] _T_60693; // @[Modules.scala 143:103:@6796.4]
  wire [4:0] _T_60694; // @[Modules.scala 143:103:@6797.4]
  wire [5:0] _T_60698; // @[Modules.scala 144:80:@6800.4]
  wire [5:0] _GEN_162; // @[Modules.scala 143:103:@6801.4]
  wire [6:0] _T_60699; // @[Modules.scala 143:103:@6801.4]
  wire [5:0] _T_60700; // @[Modules.scala 143:103:@6802.4]
  wire [5:0] _T_60701; // @[Modules.scala 143:103:@6803.4]
  wire [4:0] _T_60717; // @[Modules.scala 143:74:@6817.4]
  wire [4:0] _T_60719; // @[Modules.scala 144:80:@6818.4]
  wire [5:0] _T_60720; // @[Modules.scala 143:103:@6819.4]
  wire [4:0] _T_60721; // @[Modules.scala 143:103:@6820.4]
  wire [4:0] _T_60722; // @[Modules.scala 143:103:@6821.4]
  wire [4:0] _T_60724; // @[Modules.scala 143:74:@6823.4]
  wire [4:0] _T_60726; // @[Modules.scala 144:80:@6824.4]
  wire [5:0] _T_60727; // @[Modules.scala 143:103:@6825.4]
  wire [4:0] _T_60728; // @[Modules.scala 143:103:@6826.4]
  wire [4:0] _T_60729; // @[Modules.scala 143:103:@6827.4]
  wire [4:0] _T_60733; // @[Modules.scala 144:80:@6830.4]
  wire [5:0] _GEN_164; // @[Modules.scala 143:103:@6831.4]
  wire [6:0] _T_60734; // @[Modules.scala 143:103:@6831.4]
  wire [5:0] _T_60735; // @[Modules.scala 143:103:@6832.4]
  wire [5:0] _T_60736; // @[Modules.scala 143:103:@6833.4]
  wire [4:0] _T_60740; // @[Modules.scala 144:80:@6836.4]
  wire [5:0] _T_60741; // @[Modules.scala 143:103:@6837.4]
  wire [4:0] _T_60742; // @[Modules.scala 143:103:@6838.4]
  wire [4:0] _T_60743; // @[Modules.scala 143:103:@6839.4]
  wire [4:0] _T_60745; // @[Modules.scala 143:74:@6841.4]
  wire [4:0] _T_60747; // @[Modules.scala 144:80:@6842.4]
  wire [5:0] _T_60748; // @[Modules.scala 143:103:@6843.4]
  wire [4:0] _T_60749; // @[Modules.scala 143:103:@6844.4]
  wire [4:0] _T_60750; // @[Modules.scala 143:103:@6845.4]
  wire [4:0] _T_60752; // @[Modules.scala 143:74:@6847.4]
  wire [4:0] _T_60754; // @[Modules.scala 144:80:@6848.4]
  wire [5:0] _T_60755; // @[Modules.scala 143:103:@6849.4]
  wire [4:0] _T_60756; // @[Modules.scala 143:103:@6850.4]
  wire [4:0] _T_60757; // @[Modules.scala 143:103:@6851.4]
  wire [4:0] _T_60759; // @[Modules.scala 143:74:@6853.4]
  wire [5:0] _T_60762; // @[Modules.scala 143:103:@6855.4]
  wire [4:0] _T_60763; // @[Modules.scala 143:103:@6856.4]
  wire [4:0] _T_60764; // @[Modules.scala 143:103:@6857.4]
  wire [4:0] _T_60773; // @[Modules.scala 143:74:@6865.4]
  wire [5:0] _T_60776; // @[Modules.scala 143:103:@6867.4]
  wire [4:0] _T_60777; // @[Modules.scala 143:103:@6868.4]
  wire [4:0] _T_60778; // @[Modules.scala 143:103:@6869.4]
  wire [5:0] _T_60783; // @[Modules.scala 143:103:@6873.4]
  wire [4:0] _T_60784; // @[Modules.scala 143:103:@6874.4]
  wire [4:0] _T_60785; // @[Modules.scala 143:103:@6875.4]
  wire [4:0] _T_60808; // @[Modules.scala 143:74:@6895.4]
  wire [4:0] _T_60810; // @[Modules.scala 144:80:@6896.4]
  wire [5:0] _T_60811; // @[Modules.scala 143:103:@6897.4]
  wire [4:0] _T_60812; // @[Modules.scala 143:103:@6898.4]
  wire [4:0] _T_60813; // @[Modules.scala 143:103:@6899.4]
  wire [4:0] _T_60815; // @[Modules.scala 143:74:@6901.4]
  wire [4:0] _T_60817; // @[Modules.scala 144:80:@6902.4]
  wire [5:0] _T_60818; // @[Modules.scala 143:103:@6903.4]
  wire [4:0] _T_60819; // @[Modules.scala 143:103:@6904.4]
  wire [4:0] _T_60820; // @[Modules.scala 143:103:@6905.4]
  wire [4:0] _T_60822; // @[Modules.scala 143:74:@6907.4]
  wire [5:0] _T_60825; // @[Modules.scala 143:103:@6909.4]
  wire [4:0] _T_60826; // @[Modules.scala 143:103:@6910.4]
  wire [4:0] _T_60827; // @[Modules.scala 143:103:@6911.4]
  wire [4:0] _T_60829; // @[Modules.scala 143:74:@6913.4]
  wire [4:0] _T_60831; // @[Modules.scala 144:80:@6914.4]
  wire [5:0] _T_60832; // @[Modules.scala 143:103:@6915.4]
  wire [4:0] _T_60833; // @[Modules.scala 143:103:@6916.4]
  wire [4:0] _T_60834; // @[Modules.scala 143:103:@6917.4]
  wire [4:0] _T_60838; // @[Modules.scala 144:80:@6920.4]
  wire [5:0] _GEN_165; // @[Modules.scala 143:103:@6921.4]
  wire [6:0] _T_60839; // @[Modules.scala 143:103:@6921.4]
  wire [5:0] _T_60840; // @[Modules.scala 143:103:@6922.4]
  wire [5:0] _T_60841; // @[Modules.scala 143:103:@6923.4]
  wire [4:0] _T_60843; // @[Modules.scala 143:74:@6925.4]
  wire [4:0] _T_60845; // @[Modules.scala 144:80:@6926.4]
  wire [5:0] _T_60846; // @[Modules.scala 143:103:@6927.4]
  wire [4:0] _T_60847; // @[Modules.scala 143:103:@6928.4]
  wire [4:0] _T_60848; // @[Modules.scala 143:103:@6929.4]
  wire [4:0] _T_60850; // @[Modules.scala 143:74:@6931.4]
  wire [5:0] _T_60853; // @[Modules.scala 143:103:@6933.4]
  wire [4:0] _T_60854; // @[Modules.scala 143:103:@6934.4]
  wire [4:0] _T_60855; // @[Modules.scala 143:103:@6935.4]
  wire [5:0] _T_60860; // @[Modules.scala 143:103:@6939.4]
  wire [4:0] _T_60861; // @[Modules.scala 143:103:@6940.4]
  wire [4:0] _T_60862; // @[Modules.scala 143:103:@6941.4]
  wire [5:0] _T_60867; // @[Modules.scala 143:103:@6945.4]
  wire [4:0] _T_60868; // @[Modules.scala 143:103:@6946.4]
  wire [4:0] _T_60869; // @[Modules.scala 143:103:@6947.4]
  wire [5:0] _T_60874; // @[Modules.scala 143:103:@6951.4]
  wire [4:0] _T_60875; // @[Modules.scala 143:103:@6952.4]
  wire [4:0] _T_60876; // @[Modules.scala 143:103:@6953.4]
  wire [5:0] _T_60881; // @[Modules.scala 143:103:@6957.4]
  wire [4:0] _T_60882; // @[Modules.scala 143:103:@6958.4]
  wire [4:0] _T_60883; // @[Modules.scala 143:103:@6959.4]
  wire [5:0] _T_60888; // @[Modules.scala 143:103:@6963.4]
  wire [4:0] _T_60889; // @[Modules.scala 143:103:@6964.4]
  wire [4:0] _T_60890; // @[Modules.scala 143:103:@6965.4]
  wire [6:0] _T_60895; // @[Modules.scala 143:103:@6969.4]
  wire [5:0] _T_60896; // @[Modules.scala 143:103:@6970.4]
  wire [5:0] _T_60897; // @[Modules.scala 143:103:@6971.4]
  wire [4:0] _T_60899; // @[Modules.scala 143:74:@6973.4]
  wire [4:0] _T_60901; // @[Modules.scala 144:80:@6974.4]
  wire [5:0] _T_60902; // @[Modules.scala 143:103:@6975.4]
  wire [4:0] _T_60903; // @[Modules.scala 143:103:@6976.4]
  wire [4:0] _T_60904; // @[Modules.scala 143:103:@6977.4]
  wire [4:0] _T_60906; // @[Modules.scala 143:74:@6979.4]
  wire [4:0] _T_60908; // @[Modules.scala 144:80:@6980.4]
  wire [5:0] _T_60909; // @[Modules.scala 143:103:@6981.4]
  wire [4:0] _T_60910; // @[Modules.scala 143:103:@6982.4]
  wire [4:0] _T_60911; // @[Modules.scala 143:103:@6983.4]
  wire [4:0] _T_60913; // @[Modules.scala 143:74:@6985.4]
  wire [5:0] _T_60916; // @[Modules.scala 143:103:@6987.4]
  wire [4:0] _T_60917; // @[Modules.scala 143:103:@6988.4]
  wire [4:0] _T_60918; // @[Modules.scala 143:103:@6989.4]
  wire [4:0] _T_60920; // @[Modules.scala 143:74:@6991.4]
  wire [5:0] _T_60922; // @[Modules.scala 144:80:@6992.4]
  wire [5:0] _GEN_167; // @[Modules.scala 143:103:@6993.4]
  wire [6:0] _T_60923; // @[Modules.scala 143:103:@6993.4]
  wire [5:0] _T_60924; // @[Modules.scala 143:103:@6994.4]
  wire [5:0] _T_60925; // @[Modules.scala 143:103:@6995.4]
  wire [5:0] _T_60930; // @[Modules.scala 143:103:@6999.4]
  wire [4:0] _T_60931; // @[Modules.scala 143:103:@7000.4]
  wire [4:0] _T_60932; // @[Modules.scala 143:103:@7001.4]
  wire [4:0] _T_60934; // @[Modules.scala 143:74:@7003.4]
  wire [4:0] _T_60936; // @[Modules.scala 144:80:@7004.4]
  wire [5:0] _T_60937; // @[Modules.scala 143:103:@7005.4]
  wire [4:0] _T_60938; // @[Modules.scala 143:103:@7006.4]
  wire [4:0] _T_60939; // @[Modules.scala 143:103:@7007.4]
  wire [5:0] _T_60944; // @[Modules.scala 143:103:@7011.4]
  wire [4:0] _T_60945; // @[Modules.scala 143:103:@7012.4]
  wire [4:0] _T_60946; // @[Modules.scala 143:103:@7013.4]
  wire [4:0] _T_60983; // @[Modules.scala 143:74:@7045.4]
  wire [4:0] _T_60985; // @[Modules.scala 144:80:@7046.4]
  wire [5:0] _T_60986; // @[Modules.scala 143:103:@7047.4]
  wire [4:0] _T_60987; // @[Modules.scala 143:103:@7048.4]
  wire [4:0] _T_60988; // @[Modules.scala 143:103:@7049.4]
  wire [5:0] _T_60993; // @[Modules.scala 143:103:@7053.4]
  wire [4:0] _T_60994; // @[Modules.scala 143:103:@7054.4]
  wire [4:0] _T_60995; // @[Modules.scala 143:103:@7055.4]
  wire [5:0] _T_61000; // @[Modules.scala 143:103:@7059.4]
  wire [4:0] _T_61001; // @[Modules.scala 143:103:@7060.4]
  wire [4:0] _T_61002; // @[Modules.scala 143:103:@7061.4]
  wire [5:0] _T_61004; // @[Modules.scala 143:74:@7063.4]
  wire [5:0] _T_61006; // @[Modules.scala 144:80:@7064.4]
  wire [6:0] _T_61007; // @[Modules.scala 143:103:@7065.4]
  wire [5:0] _T_61008; // @[Modules.scala 143:103:@7066.4]
  wire [5:0] _T_61009; // @[Modules.scala 143:103:@7067.4]
  wire [4:0] _T_61013; // @[Modules.scala 144:80:@7070.4]
  wire [5:0] _T_61014; // @[Modules.scala 143:103:@7071.4]
  wire [4:0] _T_61015; // @[Modules.scala 143:103:@7072.4]
  wire [4:0] _T_61016; // @[Modules.scala 143:103:@7073.4]
  wire [4:0] _T_61018; // @[Modules.scala 143:74:@7075.4]
  wire [4:0] _T_61020; // @[Modules.scala 144:80:@7076.4]
  wire [5:0] _T_61021; // @[Modules.scala 143:103:@7077.4]
  wire [4:0] _T_61022; // @[Modules.scala 143:103:@7078.4]
  wire [4:0] _T_61023; // @[Modules.scala 143:103:@7079.4]
  wire [4:0] _T_61025; // @[Modules.scala 143:74:@7081.4]
  wire [5:0] _T_61028; // @[Modules.scala 143:103:@7083.4]
  wire [4:0] _T_61029; // @[Modules.scala 143:103:@7084.4]
  wire [4:0] _T_61030; // @[Modules.scala 143:103:@7085.4]
  wire [5:0] _T_61035; // @[Modules.scala 143:103:@7089.4]
  wire [4:0] _T_61036; // @[Modules.scala 143:103:@7090.4]
  wire [4:0] _T_61037; // @[Modules.scala 143:103:@7091.4]
  wire [5:0] _T_61042; // @[Modules.scala 143:103:@7095.4]
  wire [4:0] _T_61043; // @[Modules.scala 143:103:@7096.4]
  wire [4:0] _T_61044; // @[Modules.scala 143:103:@7097.4]
  wire [4:0] _T_61062; // @[Modules.scala 144:80:@7112.4]
  wire [5:0] _GEN_168; // @[Modules.scala 143:103:@7113.4]
  wire [6:0] _T_61063; // @[Modules.scala 143:103:@7113.4]
  wire [5:0] _T_61064; // @[Modules.scala 143:103:@7114.4]
  wire [5:0] _T_61065; // @[Modules.scala 143:103:@7115.4]
  wire [4:0] _T_61069; // @[Modules.scala 144:80:@7118.4]
  wire [5:0] _T_61070; // @[Modules.scala 143:103:@7119.4]
  wire [4:0] _T_61071; // @[Modules.scala 143:103:@7120.4]
  wire [4:0] _T_61072; // @[Modules.scala 143:103:@7121.4]
  wire [5:0] _T_61077; // @[Modules.scala 143:103:@7125.4]
  wire [4:0] _T_61078; // @[Modules.scala 143:103:@7126.4]
  wire [4:0] _T_61079; // @[Modules.scala 143:103:@7127.4]
  wire [5:0] _T_61081; // @[Modules.scala 143:74:@7129.4]
  wire [5:0] _T_61083; // @[Modules.scala 144:80:@7130.4]
  wire [6:0] _T_61084; // @[Modules.scala 143:103:@7131.4]
  wire [5:0] _T_61085; // @[Modules.scala 143:103:@7132.4]
  wire [5:0] _T_61086; // @[Modules.scala 143:103:@7133.4]
  wire [5:0] _T_61088; // @[Modules.scala 143:74:@7135.4]
  wire [5:0] _T_61090; // @[Modules.scala 144:80:@7136.4]
  wire [6:0] _T_61091; // @[Modules.scala 143:103:@7137.4]
  wire [5:0] _T_61092; // @[Modules.scala 143:103:@7138.4]
  wire [5:0] _T_61093; // @[Modules.scala 143:103:@7139.4]
  wire [5:0] _T_61095; // @[Modules.scala 143:74:@7141.4]
  wire [5:0] _T_61097; // @[Modules.scala 144:80:@7142.4]
  wire [6:0] _T_61098; // @[Modules.scala 143:103:@7143.4]
  wire [5:0] _T_61099; // @[Modules.scala 143:103:@7144.4]
  wire [5:0] _T_61100; // @[Modules.scala 143:103:@7145.4]
  wire [4:0] _T_61104; // @[Modules.scala 144:80:@7148.4]
  wire [5:0] _T_61105; // @[Modules.scala 143:103:@7149.4]
  wire [4:0] _T_61106; // @[Modules.scala 143:103:@7150.4]
  wire [4:0] _T_61107; // @[Modules.scala 143:103:@7151.4]
  wire [4:0] _T_61109; // @[Modules.scala 143:74:@7153.4]
  wire [5:0] _GEN_169; // @[Modules.scala 143:103:@7155.4]
  wire [6:0] _T_61112; // @[Modules.scala 143:103:@7155.4]
  wire [5:0] _T_61113; // @[Modules.scala 143:103:@7156.4]
  wire [5:0] _T_61114; // @[Modules.scala 143:103:@7157.4]
  wire [6:0] _T_61119; // @[Modules.scala 143:103:@7161.4]
  wire [5:0] _T_61120; // @[Modules.scala 143:103:@7162.4]
  wire [5:0] _T_61121; // @[Modules.scala 143:103:@7163.4]
  wire [5:0] _GEN_170; // @[Modules.scala 143:103:@7185.4]
  wire [6:0] _T_61147; // @[Modules.scala 143:103:@7185.4]
  wire [5:0] _T_61148; // @[Modules.scala 143:103:@7186.4]
  wire [5:0] _T_61149; // @[Modules.scala 143:103:@7187.4]
  wire [4:0] _T_61153; // @[Modules.scala 144:80:@7190.4]
  wire [5:0] _T_61154; // @[Modules.scala 143:103:@7191.4]
  wire [4:0] _T_61155; // @[Modules.scala 143:103:@7192.4]
  wire [4:0] _T_61156; // @[Modules.scala 143:103:@7193.4]
  wire [5:0] _T_61160; // @[Modules.scala 144:80:@7196.4]
  wire [5:0] _GEN_171; // @[Modules.scala 143:103:@7197.4]
  wire [6:0] _T_61161; // @[Modules.scala 143:103:@7197.4]
  wire [5:0] _T_61162; // @[Modules.scala 143:103:@7198.4]
  wire [5:0] _T_61163; // @[Modules.scala 143:103:@7199.4]
  wire [5:0] _T_61165; // @[Modules.scala 143:74:@7201.4]
  wire [5:0] _T_61167; // @[Modules.scala 144:80:@7202.4]
  wire [6:0] _T_61168; // @[Modules.scala 143:103:@7203.4]
  wire [5:0] _T_61169; // @[Modules.scala 143:103:@7204.4]
  wire [5:0] _T_61170; // @[Modules.scala 143:103:@7205.4]
  wire [5:0] _T_61172; // @[Modules.scala 143:74:@7207.4]
  wire [5:0] _T_61174; // @[Modules.scala 144:80:@7208.4]
  wire [6:0] _T_61175; // @[Modules.scala 143:103:@7209.4]
  wire [5:0] _T_61176; // @[Modules.scala 143:103:@7210.4]
  wire [5:0] _T_61177; // @[Modules.scala 143:103:@7211.4]
  wire [5:0] _T_61179; // @[Modules.scala 143:74:@7213.4]
  wire [5:0] _T_61181; // @[Modules.scala 144:80:@7214.4]
  wire [6:0] _T_61182; // @[Modules.scala 143:103:@7215.4]
  wire [5:0] _T_61183; // @[Modules.scala 143:103:@7216.4]
  wire [5:0] _T_61184; // @[Modules.scala 143:103:@7217.4]
  wire [4:0] _T_61188; // @[Modules.scala 144:80:@7220.4]
  wire [5:0] _GEN_172; // @[Modules.scala 143:103:@7221.4]
  wire [6:0] _T_61189; // @[Modules.scala 143:103:@7221.4]
  wire [5:0] _T_61190; // @[Modules.scala 143:103:@7222.4]
  wire [5:0] _T_61191; // @[Modules.scala 143:103:@7223.4]
  wire [6:0] _T_61210; // @[Modules.scala 143:103:@7239.4]
  wire [5:0] _T_61211; // @[Modules.scala 143:103:@7240.4]
  wire [5:0] _T_61212; // @[Modules.scala 143:103:@7241.4]
  wire [5:0] _T_61214; // @[Modules.scala 143:74:@7243.4]
  wire [5:0] _T_61216; // @[Modules.scala 144:80:@7244.4]
  wire [6:0] _T_61217; // @[Modules.scala 143:103:@7245.4]
  wire [5:0] _T_61218; // @[Modules.scala 143:103:@7246.4]
  wire [5:0] _T_61219; // @[Modules.scala 143:103:@7247.4]
  wire [5:0] _T_61224; // @[Modules.scala 143:103:@7251.4]
  wire [4:0] _T_61225; // @[Modules.scala 143:103:@7252.4]
  wire [4:0] _T_61226; // @[Modules.scala 143:103:@7253.4]
  wire [4:0] _T_61230; // @[Modules.scala 144:80:@7256.4]
  wire [5:0] _T_61231; // @[Modules.scala 143:103:@7257.4]
  wire [4:0] _T_61232; // @[Modules.scala 143:103:@7258.4]
  wire [4:0] _T_61233; // @[Modules.scala 143:103:@7259.4]
  wire [4:0] _T_61235; // @[Modules.scala 143:74:@7261.4]
  wire [5:0] _GEN_173; // @[Modules.scala 143:103:@7263.4]
  wire [6:0] _T_61238; // @[Modules.scala 143:103:@7263.4]
  wire [5:0] _T_61239; // @[Modules.scala 143:103:@7264.4]
  wire [5:0] _T_61240; // @[Modules.scala 143:103:@7265.4]
  wire [4:0] _T_61244; // @[Modules.scala 144:80:@7268.4]
  wire [5:0] _T_61245; // @[Modules.scala 143:103:@7269.4]
  wire [4:0] _T_61246; // @[Modules.scala 143:103:@7270.4]
  wire [4:0] _T_61247; // @[Modules.scala 143:103:@7271.4]
  wire [5:0] _GEN_174; // @[Modules.scala 143:103:@7275.4]
  wire [6:0] _T_61252; // @[Modules.scala 143:103:@7275.4]
  wire [5:0] _T_61253; // @[Modules.scala 143:103:@7276.4]
  wire [5:0] _T_61254; // @[Modules.scala 143:103:@7277.4]
  wire [5:0] _T_61258; // @[Modules.scala 144:80:@7280.4]
  wire [6:0] _T_61259; // @[Modules.scala 143:103:@7281.4]
  wire [5:0] _T_61260; // @[Modules.scala 143:103:@7282.4]
  wire [5:0] _T_61261; // @[Modules.scala 143:103:@7283.4]
  wire [5:0] _T_61265; // @[Modules.scala 144:80:@7286.4]
  wire [6:0] _T_61266; // @[Modules.scala 143:103:@7287.4]
  wire [5:0] _T_61267; // @[Modules.scala 143:103:@7288.4]
  wire [5:0] _T_61268; // @[Modules.scala 143:103:@7289.4]
  wire [5:0] _T_61270; // @[Modules.scala 143:74:@7291.4]
  wire [5:0] _T_61272; // @[Modules.scala 144:80:@7292.4]
  wire [6:0] _T_61273; // @[Modules.scala 143:103:@7293.4]
  wire [5:0] _T_61274; // @[Modules.scala 143:103:@7294.4]
  wire [5:0] _T_61275; // @[Modules.scala 143:103:@7295.4]
  wire [5:0] _T_61277; // @[Modules.scala 143:74:@7297.4]
  wire [6:0] _T_61280; // @[Modules.scala 143:103:@7299.4]
  wire [5:0] _T_61281; // @[Modules.scala 143:103:@7300.4]
  wire [5:0] _T_61282; // @[Modules.scala 143:103:@7301.4]
  wire [4:0] _T_61284; // @[Modules.scala 143:74:@7303.4]
  wire [5:0] _GEN_175; // @[Modules.scala 143:103:@7305.4]
  wire [6:0] _T_61287; // @[Modules.scala 143:103:@7305.4]
  wire [5:0] _T_61288; // @[Modules.scala 143:103:@7306.4]
  wire [5:0] _T_61289; // @[Modules.scala 143:103:@7307.4]
  wire [6:0] _T_61294; // @[Modules.scala 143:103:@7311.4]
  wire [5:0] _T_61295; // @[Modules.scala 143:103:@7312.4]
  wire [5:0] _T_61296; // @[Modules.scala 143:103:@7313.4]
  wire [6:0] _T_61301; // @[Modules.scala 143:103:@7317.4]
  wire [5:0] _T_61302; // @[Modules.scala 143:103:@7318.4]
  wire [5:0] _T_61303; // @[Modules.scala 143:103:@7319.4]
  wire [5:0] _T_61305; // @[Modules.scala 143:74:@7321.4]
  wire [5:0] _T_61307; // @[Modules.scala 144:80:@7322.4]
  wire [6:0] _T_61308; // @[Modules.scala 143:103:@7323.4]
  wire [5:0] _T_61309; // @[Modules.scala 143:103:@7324.4]
  wire [5:0] _T_61310; // @[Modules.scala 143:103:@7325.4]
  wire [6:0] _T_61315; // @[Modules.scala 143:103:@7329.4]
  wire [5:0] _T_61316; // @[Modules.scala 143:103:@7330.4]
  wire [5:0] _T_61317; // @[Modules.scala 143:103:@7331.4]
  wire [5:0] _T_61322; // @[Modules.scala 143:103:@7335.4]
  wire [4:0] _T_61323; // @[Modules.scala 143:103:@7336.4]
  wire [4:0] _T_61324; // @[Modules.scala 143:103:@7337.4]
  wire [4:0] _T_61326; // @[Modules.scala 143:74:@7339.4]
  wire [5:0] _GEN_176; // @[Modules.scala 143:103:@7341.4]
  wire [6:0] _T_61329; // @[Modules.scala 143:103:@7341.4]
  wire [5:0] _T_61330; // @[Modules.scala 143:103:@7342.4]
  wire [5:0] _T_61331; // @[Modules.scala 143:103:@7343.4]
  wire [6:0] _T_61336; // @[Modules.scala 143:103:@7347.4]
  wire [5:0] _T_61337; // @[Modules.scala 143:103:@7348.4]
  wire [5:0] _T_61338; // @[Modules.scala 143:103:@7349.4]
  wire [6:0] _T_61343; // @[Modules.scala 143:103:@7353.4]
  wire [5:0] _T_61344; // @[Modules.scala 143:103:@7354.4]
  wire [5:0] _T_61345; // @[Modules.scala 143:103:@7355.4]
  wire [5:0] _T_61349; // @[Modules.scala 144:80:@7358.4]
  wire [6:0] _T_61350; // @[Modules.scala 143:103:@7359.4]
  wire [5:0] _T_61351; // @[Modules.scala 143:103:@7360.4]
  wire [5:0] _T_61352; // @[Modules.scala 143:103:@7361.4]
  wire [5:0] _T_61354; // @[Modules.scala 143:74:@7363.4]
  wire [6:0] _T_61357; // @[Modules.scala 143:103:@7365.4]
  wire [5:0] _T_61358; // @[Modules.scala 143:103:@7366.4]
  wire [5:0] _T_61359; // @[Modules.scala 143:103:@7367.4]
  wire [5:0] _T_61361; // @[Modules.scala 143:74:@7369.4]
  wire [5:0] _T_61363; // @[Modules.scala 144:80:@7370.4]
  wire [6:0] _T_61364; // @[Modules.scala 143:103:@7371.4]
  wire [5:0] _T_61365; // @[Modules.scala 143:103:@7372.4]
  wire [5:0] _T_61366; // @[Modules.scala 143:103:@7373.4]
  wire [5:0] _T_61368; // @[Modules.scala 143:74:@7375.4]
  wire [5:0] _T_61370; // @[Modules.scala 144:80:@7376.4]
  wire [6:0] _T_61371; // @[Modules.scala 143:103:@7377.4]
  wire [5:0] _T_61372; // @[Modules.scala 143:103:@7378.4]
  wire [5:0] _T_61373; // @[Modules.scala 143:103:@7379.4]
  wire [6:0] _T_61378; // @[Modules.scala 143:103:@7383.4]
  wire [5:0] _T_61379; // @[Modules.scala 143:103:@7384.4]
  wire [5:0] _T_61380; // @[Modules.scala 143:103:@7385.4]
  wire [5:0] _T_61382; // @[Modules.scala 143:74:@7387.4]
  wire [5:0] _T_61384; // @[Modules.scala 144:80:@7388.4]
  wire [6:0] _T_61385; // @[Modules.scala 143:103:@7389.4]
  wire [5:0] _T_61386; // @[Modules.scala 143:103:@7390.4]
  wire [5:0] _T_61387; // @[Modules.scala 143:103:@7391.4]
  wire [5:0] _T_61391; // @[Modules.scala 144:80:@7394.4]
  wire [6:0] _T_61392; // @[Modules.scala 143:103:@7395.4]
  wire [5:0] _T_61393; // @[Modules.scala 143:103:@7396.4]
  wire [5:0] _T_61394; // @[Modules.scala 143:103:@7397.4]
  wire [5:0] _T_61398; // @[Modules.scala 144:80:@7400.4]
  wire [6:0] _T_61399; // @[Modules.scala 143:103:@7401.4]
  wire [5:0] _T_61400; // @[Modules.scala 143:103:@7402.4]
  wire [5:0] _T_61401; // @[Modules.scala 143:103:@7403.4]
  wire [5:0] _T_61403; // @[Modules.scala 143:74:@7405.4]
  wire [6:0] _T_61406; // @[Modules.scala 143:103:@7407.4]
  wire [5:0] _T_61407; // @[Modules.scala 143:103:@7408.4]
  wire [5:0] _T_61408; // @[Modules.scala 143:103:@7409.4]
  wire [4:0] _T_61412; // @[Modules.scala 144:80:@7412.4]
  wire [5:0] _T_61413; // @[Modules.scala 143:103:@7413.4]
  wire [4:0] _T_61414; // @[Modules.scala 143:103:@7414.4]
  wire [4:0] _T_61415; // @[Modules.scala 143:103:@7415.4]
  wire [5:0] _T_61419; // @[Modules.scala 144:80:@7418.4]
  wire [6:0] _T_61420; // @[Modules.scala 143:103:@7419.4]
  wire [5:0] _T_61421; // @[Modules.scala 143:103:@7420.4]
  wire [5:0] _T_61422; // @[Modules.scala 143:103:@7421.4]
  wire [6:0] _T_61427; // @[Modules.scala 143:103:@7425.4]
  wire [5:0] _T_61428; // @[Modules.scala 143:103:@7426.4]
  wire [5:0] _T_61429; // @[Modules.scala 143:103:@7427.4]
  wire [5:0] _T_61431; // @[Modules.scala 143:74:@7429.4]
  wire [5:0] _T_61433; // @[Modules.scala 144:80:@7430.4]
  wire [6:0] _T_61434; // @[Modules.scala 143:103:@7431.4]
  wire [5:0] _T_61435; // @[Modules.scala 143:103:@7432.4]
  wire [5:0] _T_61436; // @[Modules.scala 143:103:@7433.4]
  wire [5:0] _T_61438; // @[Modules.scala 143:74:@7435.4]
  wire [5:0] _T_61440; // @[Modules.scala 144:80:@7436.4]
  wire [6:0] _T_61441; // @[Modules.scala 143:103:@7437.4]
  wire [5:0] _T_61442; // @[Modules.scala 143:103:@7438.4]
  wire [5:0] _T_61443; // @[Modules.scala 143:103:@7439.4]
  wire [5:0] _T_61445; // @[Modules.scala 143:74:@7441.4]
  wire [5:0] _T_61447; // @[Modules.scala 144:80:@7442.4]
  wire [6:0] _T_61448; // @[Modules.scala 143:103:@7443.4]
  wire [5:0] _T_61449; // @[Modules.scala 143:103:@7444.4]
  wire [5:0] _T_61450; // @[Modules.scala 143:103:@7445.4]
  wire [4:0] _T_61454; // @[Modules.scala 144:80:@7448.4]
  wire [5:0] _GEN_177; // @[Modules.scala 143:103:@7449.4]
  wire [6:0] _T_61455; // @[Modules.scala 143:103:@7449.4]
  wire [5:0] _T_61456; // @[Modules.scala 143:103:@7450.4]
  wire [5:0] _T_61457; // @[Modules.scala 143:103:@7451.4]
  wire [6:0] _T_61462; // @[Modules.scala 143:103:@7455.4]
  wire [5:0] _T_61463; // @[Modules.scala 143:103:@7456.4]
  wire [5:0] _T_61464; // @[Modules.scala 143:103:@7457.4]
  wire [5:0] _T_61466; // @[Modules.scala 143:74:@7459.4]
  wire [5:0] _T_61468; // @[Modules.scala 144:80:@7460.4]
  wire [6:0] _T_61469; // @[Modules.scala 143:103:@7461.4]
  wire [5:0] _T_61470; // @[Modules.scala 143:103:@7462.4]
  wire [5:0] _T_61471; // @[Modules.scala 143:103:@7463.4]
  wire [4:0] _T_61473; // @[Modules.scala 143:74:@7465.4]
  wire [4:0] _T_61475; // @[Modules.scala 144:80:@7466.4]
  wire [5:0] _T_61476; // @[Modules.scala 143:103:@7467.4]
  wire [4:0] _T_61477; // @[Modules.scala 143:103:@7468.4]
  wire [4:0] _T_61478; // @[Modules.scala 143:103:@7469.4]
  wire [6:0] _T_61483; // @[Modules.scala 143:103:@7473.4]
  wire [5:0] _T_61484; // @[Modules.scala 143:103:@7474.4]
  wire [5:0] _T_61485; // @[Modules.scala 143:103:@7475.4]
  wire [5:0] _T_61489; // @[Modules.scala 144:80:@7478.4]
  wire [6:0] _T_61490; // @[Modules.scala 143:103:@7479.4]
  wire [5:0] _T_61491; // @[Modules.scala 143:103:@7480.4]
  wire [5:0] _T_61492; // @[Modules.scala 143:103:@7481.4]
  wire [4:0] _T_61496; // @[Modules.scala 144:80:@7484.4]
  wire [5:0] _T_61497; // @[Modules.scala 143:103:@7485.4]
  wire [4:0] _T_61498; // @[Modules.scala 143:103:@7486.4]
  wire [4:0] _T_61499; // @[Modules.scala 143:103:@7487.4]
  wire [5:0] _T_61503; // @[Modules.scala 144:80:@7490.4]
  wire [5:0] _GEN_179; // @[Modules.scala 143:103:@7491.4]
  wire [6:0] _T_61504; // @[Modules.scala 143:103:@7491.4]
  wire [5:0] _T_61505; // @[Modules.scala 143:103:@7492.4]
  wire [5:0] _T_61506; // @[Modules.scala 143:103:@7493.4]
  wire [4:0] _T_61510; // @[Modules.scala 144:80:@7496.4]
  wire [5:0] _GEN_180; // @[Modules.scala 143:103:@7497.4]
  wire [6:0] _T_61511; // @[Modules.scala 143:103:@7497.4]
  wire [5:0] _T_61512; // @[Modules.scala 143:103:@7498.4]
  wire [5:0] _T_61513; // @[Modules.scala 143:103:@7499.4]
  wire [5:0] _T_61522; // @[Modules.scala 143:74:@7507.4]
  wire [6:0] _T_61525; // @[Modules.scala 143:103:@7509.4]
  wire [5:0] _T_61526; // @[Modules.scala 143:103:@7510.4]
  wire [5:0] _T_61527; // @[Modules.scala 143:103:@7511.4]
  wire [5:0] _GEN_181; // @[Modules.scala 143:103:@7515.4]
  wire [6:0] _T_61532; // @[Modules.scala 143:103:@7515.4]
  wire [5:0] _T_61533; // @[Modules.scala 143:103:@7516.4]
  wire [5:0] _T_61534; // @[Modules.scala 143:103:@7517.4]
  wire [4:0] _T_61536; // @[Modules.scala 143:74:@7519.4]
  wire [5:0] _GEN_182; // @[Modules.scala 143:103:@7521.4]
  wire [6:0] _T_61539; // @[Modules.scala 143:103:@7521.4]
  wire [5:0] _T_61540; // @[Modules.scala 143:103:@7522.4]
  wire [5:0] _T_61541; // @[Modules.scala 143:103:@7523.4]
  wire [5:0] _T_61545; // @[Modules.scala 144:80:@7526.4]
  wire [6:0] _T_61546; // @[Modules.scala 143:103:@7527.4]
  wire [5:0] _T_61547; // @[Modules.scala 143:103:@7528.4]
  wire [5:0] _T_61548; // @[Modules.scala 143:103:@7529.4]
  wire [4:0] _T_61552; // @[Modules.scala 144:80:@7532.4]
  wire [5:0] _GEN_183; // @[Modules.scala 143:103:@7533.4]
  wire [6:0] _T_61553; // @[Modules.scala 143:103:@7533.4]
  wire [5:0] _T_61554; // @[Modules.scala 143:103:@7534.4]
  wire [5:0] _T_61555; // @[Modules.scala 143:103:@7535.4]
  wire [5:0] _T_61557; // @[Modules.scala 143:74:@7537.4]
  wire [6:0] _T_61560; // @[Modules.scala 143:103:@7539.4]
  wire [5:0] _T_61561; // @[Modules.scala 143:103:@7540.4]
  wire [5:0] _T_61562; // @[Modules.scala 143:103:@7541.4]
  wire [4:0] _T_61564; // @[Modules.scala 143:74:@7543.4]
  wire [5:0] _T_61567; // @[Modules.scala 143:103:@7545.4]
  wire [4:0] _T_61568; // @[Modules.scala 143:103:@7546.4]
  wire [4:0] _T_61569; // @[Modules.scala 143:103:@7547.4]
  wire [4:0] _T_61573; // @[Modules.scala 144:80:@7550.4]
  wire [5:0] _T_61574; // @[Modules.scala 143:103:@7551.4]
  wire [4:0] _T_61575; // @[Modules.scala 143:103:@7552.4]
  wire [4:0] _T_61576; // @[Modules.scala 143:103:@7553.4]
  wire [4:0] _T_61578; // @[Modules.scala 143:74:@7555.4]
  wire [5:0] _T_61580; // @[Modules.scala 144:80:@7556.4]
  wire [5:0] _GEN_184; // @[Modules.scala 143:103:@7557.4]
  wire [6:0] _T_61581; // @[Modules.scala 143:103:@7557.4]
  wire [5:0] _T_61582; // @[Modules.scala 143:103:@7558.4]
  wire [5:0] _T_61583; // @[Modules.scala 143:103:@7559.4]
  wire [4:0] _T_61585; // @[Modules.scala 143:74:@7561.4]
  wire [4:0] _T_61587; // @[Modules.scala 144:80:@7562.4]
  wire [5:0] _T_61588; // @[Modules.scala 143:103:@7563.4]
  wire [4:0] _T_61589; // @[Modules.scala 143:103:@7564.4]
  wire [4:0] _T_61590; // @[Modules.scala 143:103:@7565.4]
  wire [4:0] _T_61592; // @[Modules.scala 143:74:@7567.4]
  wire [5:0] _T_61595; // @[Modules.scala 143:103:@7569.4]
  wire [4:0] _T_61596; // @[Modules.scala 143:103:@7570.4]
  wire [4:0] _T_61597; // @[Modules.scala 143:103:@7571.4]
  wire [5:0] _T_61601; // @[Modules.scala 144:80:@7574.4]
  wire [5:0] _GEN_185; // @[Modules.scala 143:103:@7575.4]
  wire [6:0] _T_61602; // @[Modules.scala 143:103:@7575.4]
  wire [5:0] _T_61603; // @[Modules.scala 143:103:@7576.4]
  wire [5:0] _T_61604; // @[Modules.scala 143:103:@7577.4]
  wire [5:0] _T_61606; // @[Modules.scala 143:74:@7579.4]
  wire [6:0] _T_61609; // @[Modules.scala 143:103:@7581.4]
  wire [5:0] _T_61610; // @[Modules.scala 143:103:@7582.4]
  wire [5:0] _T_61611; // @[Modules.scala 143:103:@7583.4]
  wire [6:0] _T_61616; // @[Modules.scala 143:103:@7587.4]
  wire [5:0] _T_61617; // @[Modules.scala 143:103:@7588.4]
  wire [5:0] _T_61618; // @[Modules.scala 143:103:@7589.4]
  wire [5:0] _T_61622; // @[Modules.scala 144:80:@7592.4]
  wire [6:0] _T_61623; // @[Modules.scala 143:103:@7593.4]
  wire [5:0] _T_61624; // @[Modules.scala 143:103:@7594.4]
  wire [5:0] _T_61625; // @[Modules.scala 143:103:@7595.4]
  wire [4:0] _T_61629; // @[Modules.scala 144:80:@7598.4]
  wire [5:0] _GEN_186; // @[Modules.scala 143:103:@7599.4]
  wire [6:0] _T_61630; // @[Modules.scala 143:103:@7599.4]
  wire [5:0] _T_61631; // @[Modules.scala 143:103:@7600.4]
  wire [5:0] _T_61632; // @[Modules.scala 143:103:@7601.4]
  wire [5:0] _T_61637; // @[Modules.scala 143:103:@7605.4]
  wire [4:0] _T_61638; // @[Modules.scala 143:103:@7606.4]
  wire [4:0] _T_61639; // @[Modules.scala 143:103:@7607.4]
  wire [4:0] _T_61643; // @[Modules.scala 144:80:@7610.4]
  wire [5:0] _T_61644; // @[Modules.scala 143:103:@7611.4]
  wire [4:0] _T_61645; // @[Modules.scala 143:103:@7612.4]
  wire [4:0] _T_61646; // @[Modules.scala 143:103:@7613.4]
  wire [6:0] _T_61651; // @[Modules.scala 143:103:@7617.4]
  wire [5:0] _T_61652; // @[Modules.scala 143:103:@7618.4]
  wire [5:0] _T_61653; // @[Modules.scala 143:103:@7619.4]
  wire [4:0] _T_61657; // @[Modules.scala 144:80:@7622.4]
  wire [5:0] _GEN_188; // @[Modules.scala 143:103:@7623.4]
  wire [6:0] _T_61658; // @[Modules.scala 143:103:@7623.4]
  wire [5:0] _T_61659; // @[Modules.scala 143:103:@7624.4]
  wire [5:0] _T_61660; // @[Modules.scala 143:103:@7625.4]
  wire [4:0] _T_61662; // @[Modules.scala 143:74:@7627.4]
  wire [5:0] _T_61665; // @[Modules.scala 143:103:@7629.4]
  wire [4:0] _T_61666; // @[Modules.scala 143:103:@7630.4]
  wire [4:0] _T_61667; // @[Modules.scala 143:103:@7631.4]
  wire [5:0] _T_61676; // @[Modules.scala 143:74:@7639.4]
  wire [6:0] _T_61679; // @[Modules.scala 143:103:@7641.4]
  wire [5:0] _T_61680; // @[Modules.scala 143:103:@7642.4]
  wire [5:0] _T_61681; // @[Modules.scala 143:103:@7643.4]
  wire [4:0] _T_61699; // @[Modules.scala 144:80:@7658.4]
  wire [5:0] _GEN_189; // @[Modules.scala 143:103:@7659.4]
  wire [6:0] _T_61700; // @[Modules.scala 143:103:@7659.4]
  wire [5:0] _T_61701; // @[Modules.scala 143:103:@7660.4]
  wire [5:0] _T_61702; // @[Modules.scala 143:103:@7661.4]
  wire [4:0] _T_61706; // @[Modules.scala 144:80:@7664.4]
  wire [5:0] _GEN_190; // @[Modules.scala 143:103:@7665.4]
  wire [6:0] _T_61707; // @[Modules.scala 143:103:@7665.4]
  wire [5:0] _T_61708; // @[Modules.scala 143:103:@7666.4]
  wire [5:0] _T_61709; // @[Modules.scala 143:103:@7667.4]
  wire [4:0] _T_61725; // @[Modules.scala 143:74:@7681.4]
  wire [5:0] _GEN_191; // @[Modules.scala 143:103:@7683.4]
  wire [6:0] _T_61728; // @[Modules.scala 143:103:@7683.4]
  wire [5:0] _T_61729; // @[Modules.scala 143:103:@7684.4]
  wire [5:0] _T_61730; // @[Modules.scala 143:103:@7685.4]
  wire [6:0] _T_61735; // @[Modules.scala 143:103:@7689.4]
  wire [5:0] _T_61736; // @[Modules.scala 143:103:@7690.4]
  wire [5:0] _T_61737; // @[Modules.scala 143:103:@7691.4]
  wire [4:0] _T_61739; // @[Modules.scala 143:74:@7693.4]
  wire [4:0] _T_61741; // @[Modules.scala 144:80:@7694.4]
  wire [5:0] _T_61742; // @[Modules.scala 143:103:@7695.4]
  wire [4:0] _T_61743; // @[Modules.scala 143:103:@7696.4]
  wire [4:0] _T_61744; // @[Modules.scala 143:103:@7697.4]
  wire [4:0] _T_61753; // @[Modules.scala 143:74:@7705.4]
  wire [5:0] _T_61756; // @[Modules.scala 143:103:@7707.4]
  wire [4:0] _T_61757; // @[Modules.scala 143:103:@7708.4]
  wire [4:0] _T_61758; // @[Modules.scala 143:103:@7709.4]
  wire [5:0] _GEN_192; // @[Modules.scala 143:103:@7713.4]
  wire [6:0] _T_61763; // @[Modules.scala 143:103:@7713.4]
  wire [5:0] _T_61764; // @[Modules.scala 143:103:@7714.4]
  wire [5:0] _T_61765; // @[Modules.scala 143:103:@7715.4]
  wire [5:0] _GEN_193; // @[Modules.scala 143:103:@7719.4]
  wire [6:0] _T_61770; // @[Modules.scala 143:103:@7719.4]
  wire [5:0] _T_61771; // @[Modules.scala 143:103:@7720.4]
  wire [5:0] _T_61772; // @[Modules.scala 143:103:@7721.4]
  wire [4:0] _T_61774; // @[Modules.scala 143:74:@7723.4]
  wire [5:0] _GEN_194; // @[Modules.scala 143:103:@7725.4]
  wire [6:0] _T_61777; // @[Modules.scala 143:103:@7725.4]
  wire [5:0] _T_61778; // @[Modules.scala 143:103:@7726.4]
  wire [5:0] _T_61779; // @[Modules.scala 143:103:@7727.4]
  wire [5:0] _GEN_195; // @[Modules.scala 143:103:@7731.4]
  wire [6:0] _T_61784; // @[Modules.scala 143:103:@7731.4]
  wire [5:0] _T_61785; // @[Modules.scala 143:103:@7732.4]
  wire [5:0] _T_61786; // @[Modules.scala 143:103:@7733.4]
  wire [5:0] _T_61809; // @[Modules.scala 143:74:@7753.4]
  wire [6:0] _T_61812; // @[Modules.scala 143:103:@7755.4]
  wire [5:0] _T_61813; // @[Modules.scala 143:103:@7756.4]
  wire [5:0] _T_61814; // @[Modules.scala 143:103:@7757.4]
  wire [4:0] _T_61816; // @[Modules.scala 143:74:@7759.4]
  wire [4:0] _T_61818; // @[Modules.scala 144:80:@7760.4]
  wire [5:0] _T_61819; // @[Modules.scala 143:103:@7761.4]
  wire [4:0] _T_61820; // @[Modules.scala 143:103:@7762.4]
  wire [4:0] _T_61821; // @[Modules.scala 143:103:@7763.4]
  wire [5:0] _T_61826; // @[Modules.scala 143:103:@7767.4]
  wire [4:0] _T_61827; // @[Modules.scala 143:103:@7768.4]
  wire [4:0] _T_61828; // @[Modules.scala 143:103:@7769.4]
  wire [4:0] _T_61830; // @[Modules.scala 143:74:@7771.4]
  wire [4:0] _T_61832; // @[Modules.scala 144:80:@7772.4]
  wire [5:0] _T_61833; // @[Modules.scala 143:103:@7773.4]
  wire [4:0] _T_61834; // @[Modules.scala 143:103:@7774.4]
  wire [4:0] _T_61835; // @[Modules.scala 143:103:@7775.4]
  wire [4:0] _T_61837; // @[Modules.scala 143:74:@7777.4]
  wire [4:0] _T_61839; // @[Modules.scala 144:80:@7778.4]
  wire [5:0] _T_61840; // @[Modules.scala 143:103:@7779.4]
  wire [4:0] _T_61841; // @[Modules.scala 143:103:@7780.4]
  wire [4:0] _T_61842; // @[Modules.scala 143:103:@7781.4]
  wire [5:0] _T_61846; // @[Modules.scala 144:80:@7784.4]
  wire [6:0] _T_61847; // @[Modules.scala 143:103:@7785.4]
  wire [5:0] _T_61848; // @[Modules.scala 143:103:@7786.4]
  wire [5:0] _T_61849; // @[Modules.scala 143:103:@7787.4]
  wire [5:0] _T_61851; // @[Modules.scala 143:74:@7789.4]
  wire [5:0] _GEN_196; // @[Modules.scala 143:103:@7791.4]
  wire [6:0] _T_61854; // @[Modules.scala 143:103:@7791.4]
  wire [5:0] _T_61855; // @[Modules.scala 143:103:@7792.4]
  wire [5:0] _T_61856; // @[Modules.scala 143:103:@7793.4]
  wire [4:0] _T_61858; // @[Modules.scala 143:74:@7795.4]
  wire [5:0] _T_61861; // @[Modules.scala 143:103:@7797.4]
  wire [4:0] _T_61862; // @[Modules.scala 143:103:@7798.4]
  wire [4:0] _T_61863; // @[Modules.scala 143:103:@7799.4]
  wire [5:0] _T_61868; // @[Modules.scala 143:103:@7803.4]
  wire [4:0] _T_61869; // @[Modules.scala 143:103:@7804.4]
  wire [4:0] _T_61870; // @[Modules.scala 143:103:@7805.4]
  wire [5:0] _GEN_197; // @[Modules.scala 143:103:@7809.4]
  wire [6:0] _T_61875; // @[Modules.scala 143:103:@7809.4]
  wire [5:0] _T_61876; // @[Modules.scala 143:103:@7810.4]
  wire [5:0] _T_61877; // @[Modules.scala 143:103:@7811.4]
  wire [4:0] _T_61879; // @[Modules.scala 143:74:@7813.4]
  wire [5:0] _GEN_198; // @[Modules.scala 143:103:@7815.4]
  wire [6:0] _T_61882; // @[Modules.scala 143:103:@7815.4]
  wire [5:0] _T_61883; // @[Modules.scala 143:103:@7816.4]
  wire [5:0] _T_61884; // @[Modules.scala 143:103:@7817.4]
  wire [6:0] _T_61889; // @[Modules.scala 143:103:@7821.4]
  wire [5:0] _T_61890; // @[Modules.scala 143:103:@7822.4]
  wire [5:0] _T_61891; // @[Modules.scala 143:103:@7823.4]
  wire [4:0] _T_61895; // @[Modules.scala 144:80:@7826.4]
  wire [5:0] _GEN_199; // @[Modules.scala 143:103:@7827.4]
  wire [6:0] _T_61896; // @[Modules.scala 143:103:@7827.4]
  wire [5:0] _T_61897; // @[Modules.scala 143:103:@7828.4]
  wire [5:0] _T_61898; // @[Modules.scala 143:103:@7829.4]
  wire [4:0] _T_61900; // @[Modules.scala 143:74:@7831.4]
  wire [4:0] _T_61902; // @[Modules.scala 144:80:@7832.4]
  wire [5:0] _T_61903; // @[Modules.scala 143:103:@7833.4]
  wire [4:0] _T_61904; // @[Modules.scala 143:103:@7834.4]
  wire [4:0] _T_61905; // @[Modules.scala 143:103:@7835.4]
  wire [4:0] _T_61907; // @[Modules.scala 143:74:@7837.4]
  wire [5:0] _T_61910; // @[Modules.scala 143:103:@7839.4]
  wire [4:0] _T_61911; // @[Modules.scala 143:103:@7840.4]
  wire [4:0] _T_61912; // @[Modules.scala 143:103:@7841.4]
  wire [4:0] _T_61914; // @[Modules.scala 143:74:@7843.4]
  wire [4:0] _T_61916; // @[Modules.scala 144:80:@7844.4]
  wire [5:0] _T_61917; // @[Modules.scala 143:103:@7845.4]
  wire [4:0] _T_61918; // @[Modules.scala 143:103:@7846.4]
  wire [4:0] _T_61919; // @[Modules.scala 143:103:@7847.4]
  wire [4:0] _T_61921; // @[Modules.scala 143:74:@7849.4]
  wire [5:0] _T_61923; // @[Modules.scala 144:80:@7850.4]
  wire [5:0] _GEN_200; // @[Modules.scala 143:103:@7851.4]
  wire [6:0] _T_61924; // @[Modules.scala 143:103:@7851.4]
  wire [5:0] _T_61925; // @[Modules.scala 143:103:@7852.4]
  wire [5:0] _T_61926; // @[Modules.scala 143:103:@7853.4]
  wire [6:0] _T_61931; // @[Modules.scala 143:103:@7857.4]
  wire [5:0] _T_61932; // @[Modules.scala 143:103:@7858.4]
  wire [5:0] _T_61933; // @[Modules.scala 143:103:@7859.4]
  wire [5:0] _T_61937; // @[Modules.scala 144:80:@7862.4]
  wire [6:0] _T_61938; // @[Modules.scala 143:103:@7863.4]
  wire [5:0] _T_61939; // @[Modules.scala 143:103:@7864.4]
  wire [5:0] _T_61940; // @[Modules.scala 143:103:@7865.4]
  wire [4:0] _T_61944; // @[Modules.scala 144:80:@7868.4]
  wire [5:0] _T_61945; // @[Modules.scala 143:103:@7869.4]
  wire [4:0] _T_61946; // @[Modules.scala 143:103:@7870.4]
  wire [4:0] _T_61947; // @[Modules.scala 143:103:@7871.4]
  wire [5:0] _GEN_201; // @[Modules.scala 143:103:@7881.4]
  wire [6:0] _T_61959; // @[Modules.scala 143:103:@7881.4]
  wire [5:0] _T_61960; // @[Modules.scala 143:103:@7882.4]
  wire [5:0] _T_61961; // @[Modules.scala 143:103:@7883.4]
  wire [5:0] _GEN_202; // @[Modules.scala 143:103:@7887.4]
  wire [6:0] _T_61966; // @[Modules.scala 143:103:@7887.4]
  wire [5:0] _T_61967; // @[Modules.scala 143:103:@7888.4]
  wire [5:0] _T_61968; // @[Modules.scala 143:103:@7889.4]
  wire [6:0] _T_61973; // @[Modules.scala 143:103:@7893.4]
  wire [5:0] _T_61974; // @[Modules.scala 143:103:@7894.4]
  wire [5:0] _T_61975; // @[Modules.scala 143:103:@7895.4]
  wire [4:0] _T_61979; // @[Modules.scala 144:80:@7898.4]
  wire [5:0] _GEN_203; // @[Modules.scala 143:103:@7899.4]
  wire [6:0] _T_61980; // @[Modules.scala 143:103:@7899.4]
  wire [5:0] _T_61981; // @[Modules.scala 143:103:@7900.4]
  wire [5:0] _T_61982; // @[Modules.scala 143:103:@7901.4]
  wire [4:0] _T_61984; // @[Modules.scala 143:74:@7903.4]
  wire [4:0] _T_61986; // @[Modules.scala 144:80:@7904.4]
  wire [5:0] _T_61987; // @[Modules.scala 143:103:@7905.4]
  wire [4:0] _T_61988; // @[Modules.scala 143:103:@7906.4]
  wire [4:0] _T_61989; // @[Modules.scala 143:103:@7907.4]
  wire [4:0] _T_61991; // @[Modules.scala 143:74:@7909.4]
  wire [5:0] _T_61994; // @[Modules.scala 143:103:@7911.4]
  wire [4:0] _T_61995; // @[Modules.scala 143:103:@7912.4]
  wire [4:0] _T_61996; // @[Modules.scala 143:103:@7913.4]
  wire [4:0] _T_61998; // @[Modules.scala 143:74:@7915.4]
  wire [4:0] _T_62000; // @[Modules.scala 144:80:@7916.4]
  wire [5:0] _T_62001; // @[Modules.scala 143:103:@7917.4]
  wire [4:0] _T_62002; // @[Modules.scala 143:103:@7918.4]
  wire [4:0] _T_62003; // @[Modules.scala 143:103:@7919.4]
  wire [4:0] _T_62005; // @[Modules.scala 143:74:@7921.4]
  wire [5:0] _T_62008; // @[Modules.scala 143:103:@7923.4]
  wire [4:0] _T_62009; // @[Modules.scala 143:103:@7924.4]
  wire [4:0] _T_62010; // @[Modules.scala 143:103:@7925.4]
  wire [5:0] _T_62015; // @[Modules.scala 143:103:@7929.4]
  wire [4:0] _T_62016; // @[Modules.scala 143:103:@7930.4]
  wire [4:0] _T_62017; // @[Modules.scala 143:103:@7931.4]
  wire [5:0] _T_62022; // @[Modules.scala 143:103:@7935.4]
  wire [4:0] _T_62023; // @[Modules.scala 143:103:@7936.4]
  wire [4:0] _T_62024; // @[Modules.scala 143:103:@7937.4]
  wire [5:0] _T_62026; // @[Modules.scala 143:74:@7939.4]
  wire [6:0] _T_62029; // @[Modules.scala 143:103:@7941.4]
  wire [5:0] _T_62030; // @[Modules.scala 143:103:@7942.4]
  wire [5:0] _T_62031; // @[Modules.scala 143:103:@7943.4]
  wire [6:0] _T_62036; // @[Modules.scala 143:103:@7947.4]
  wire [5:0] _T_62037; // @[Modules.scala 143:103:@7948.4]
  wire [5:0] _T_62038; // @[Modules.scala 143:103:@7949.4]
  wire [4:0] _T_62049; // @[Modules.scala 144:80:@7958.4]
  wire [5:0] _GEN_205; // @[Modules.scala 143:103:@7959.4]
  wire [6:0] _T_62050; // @[Modules.scala 143:103:@7959.4]
  wire [5:0] _T_62051; // @[Modules.scala 143:103:@7960.4]
  wire [5:0] _T_62052; // @[Modules.scala 143:103:@7961.4]
  wire [4:0] _T_62054; // @[Modules.scala 143:74:@7963.4]
  wire [4:0] _T_62056; // @[Modules.scala 144:80:@7964.4]
  wire [5:0] _T_62057; // @[Modules.scala 143:103:@7965.4]
  wire [4:0] _T_62058; // @[Modules.scala 143:103:@7966.4]
  wire [4:0] _T_62059; // @[Modules.scala 143:103:@7967.4]
  wire [4:0] _T_62061; // @[Modules.scala 143:74:@7969.4]
  wire [4:0] _T_62063; // @[Modules.scala 144:80:@7970.4]
  wire [5:0] _T_62064; // @[Modules.scala 143:103:@7971.4]
  wire [4:0] _T_62065; // @[Modules.scala 143:103:@7972.4]
  wire [4:0] _T_62066; // @[Modules.scala 143:103:@7973.4]
  wire [5:0] _T_62103; // @[Modules.scala 143:74:@8005.4]
  wire [6:0] _T_62106; // @[Modules.scala 143:103:@8007.4]
  wire [5:0] _T_62107; // @[Modules.scala 143:103:@8008.4]
  wire [5:0] _T_62108; // @[Modules.scala 143:103:@8009.4]
  wire [5:0] _T_62110; // @[Modules.scala 143:74:@8011.4]
  wire [5:0] _T_62112; // @[Modules.scala 144:80:@8012.4]
  wire [6:0] _T_62113; // @[Modules.scala 143:103:@8013.4]
  wire [5:0] _T_62114; // @[Modules.scala 143:103:@8014.4]
  wire [5:0] _T_62115; // @[Modules.scala 143:103:@8015.4]
  wire [4:0] _T_62126; // @[Modules.scala 144:80:@8024.4]
  wire [5:0] _T_62127; // @[Modules.scala 143:103:@8025.4]
  wire [4:0] _T_62128; // @[Modules.scala 143:103:@8026.4]
  wire [4:0] _T_62129; // @[Modules.scala 143:103:@8027.4]
  wire [4:0] _T_62138; // @[Modules.scala 143:74:@8035.4]
  wire [4:0] _T_62140; // @[Modules.scala 144:80:@8036.4]
  wire [5:0] _T_62141; // @[Modules.scala 143:103:@8037.4]
  wire [4:0] _T_62142; // @[Modules.scala 143:103:@8038.4]
  wire [4:0] _T_62143; // @[Modules.scala 143:103:@8039.4]
  wire [4:0] _T_62145; // @[Modules.scala 143:74:@8041.4]
  wire [4:0] _T_62147; // @[Modules.scala 144:80:@8042.4]
  wire [5:0] _T_62148; // @[Modules.scala 143:103:@8043.4]
  wire [4:0] _T_62149; // @[Modules.scala 143:103:@8044.4]
  wire [4:0] _T_62150; // @[Modules.scala 143:103:@8045.4]
  wire [6:0] _T_62155; // @[Modules.scala 143:103:@8049.4]
  wire [5:0] _T_62156; // @[Modules.scala 143:103:@8050.4]
  wire [5:0] _T_62157; // @[Modules.scala 143:103:@8051.4]
  wire [5:0] _T_62159; // @[Modules.scala 143:74:@8053.4]
  wire [5:0] _GEN_206; // @[Modules.scala 143:103:@8055.4]
  wire [6:0] _T_62162; // @[Modules.scala 143:103:@8055.4]
  wire [5:0] _T_62163; // @[Modules.scala 143:103:@8056.4]
  wire [5:0] _T_62164; // @[Modules.scala 143:103:@8057.4]
  wire [6:0] _T_62183; // @[Modules.scala 143:103:@8073.4]
  wire [5:0] _T_62184; // @[Modules.scala 143:103:@8074.4]
  wire [5:0] _T_62185; // @[Modules.scala 143:103:@8075.4]
  wire [5:0] _T_62187; // @[Modules.scala 143:74:@8077.4]
  wire [5:0] _T_62189; // @[Modules.scala 144:80:@8078.4]
  wire [6:0] _T_62190; // @[Modules.scala 143:103:@8079.4]
  wire [5:0] _T_62191; // @[Modules.scala 143:103:@8080.4]
  wire [5:0] _T_62192; // @[Modules.scala 143:103:@8081.4]
  wire [5:0] _T_62194; // @[Modules.scala 143:74:@8083.4]
  wire [6:0] _T_62197; // @[Modules.scala 143:103:@8085.4]
  wire [5:0] _T_62198; // @[Modules.scala 143:103:@8086.4]
  wire [5:0] _T_62199; // @[Modules.scala 143:103:@8087.4]
  wire [4:0] _T_62203; // @[Modules.scala 144:80:@8090.4]
  wire [5:0] _GEN_208; // @[Modules.scala 143:103:@8091.4]
  wire [6:0] _T_62204; // @[Modules.scala 143:103:@8091.4]
  wire [5:0] _T_62205; // @[Modules.scala 143:103:@8092.4]
  wire [5:0] _T_62206; // @[Modules.scala 143:103:@8093.4]
  wire [4:0] _T_62210; // @[Modules.scala 144:80:@8096.4]
  wire [5:0] _T_62211; // @[Modules.scala 143:103:@8097.4]
  wire [4:0] _T_62212; // @[Modules.scala 143:103:@8098.4]
  wire [4:0] _T_62213; // @[Modules.scala 143:103:@8099.4]
  wire [4:0] _T_62215; // @[Modules.scala 143:74:@8101.4]
  wire [5:0] _GEN_209; // @[Modules.scala 143:103:@8103.4]
  wire [6:0] _T_62218; // @[Modules.scala 143:103:@8103.4]
  wire [5:0] _T_62219; // @[Modules.scala 143:103:@8104.4]
  wire [5:0] _T_62220; // @[Modules.scala 143:103:@8105.4]
  wire [6:0] _T_62225; // @[Modules.scala 143:103:@8109.4]
  wire [5:0] _T_62226; // @[Modules.scala 143:103:@8110.4]
  wire [5:0] _T_62227; // @[Modules.scala 143:103:@8111.4]
  wire [4:0] _T_62231; // @[Modules.scala 144:80:@8114.4]
  wire [5:0] _GEN_211; // @[Modules.scala 143:103:@8115.4]
  wire [6:0] _T_62232; // @[Modules.scala 143:103:@8115.4]
  wire [5:0] _T_62233; // @[Modules.scala 143:103:@8116.4]
  wire [5:0] _T_62234; // @[Modules.scala 143:103:@8117.4]
  wire [5:0] _T_62239; // @[Modules.scala 143:103:@8121.4]
  wire [4:0] _T_62240; // @[Modules.scala 143:103:@8122.4]
  wire [4:0] _T_62241; // @[Modules.scala 143:103:@8123.4]
  wire [5:0] _T_62246; // @[Modules.scala 143:103:@8127.4]
  wire [4:0] _T_62247; // @[Modules.scala 143:103:@8128.4]
  wire [4:0] _T_62248; // @[Modules.scala 143:103:@8129.4]
  wire [5:0] _GEN_212; // @[Modules.scala 143:103:@8133.4]
  wire [6:0] _T_62253; // @[Modules.scala 143:103:@8133.4]
  wire [5:0] _T_62254; // @[Modules.scala 143:103:@8134.4]
  wire [5:0] _T_62255; // @[Modules.scala 143:103:@8135.4]
  wire [5:0] _GEN_213; // @[Modules.scala 143:103:@8139.4]
  wire [6:0] _T_62260; // @[Modules.scala 143:103:@8139.4]
  wire [5:0] _T_62261; // @[Modules.scala 143:103:@8140.4]
  wire [5:0] _T_62262; // @[Modules.scala 143:103:@8141.4]
  wire [5:0] _T_62273; // @[Modules.scala 144:80:@8150.4]
  wire [5:0] _GEN_214; // @[Modules.scala 143:103:@8151.4]
  wire [6:0] _T_62274; // @[Modules.scala 143:103:@8151.4]
  wire [5:0] _T_62275; // @[Modules.scala 143:103:@8152.4]
  wire [5:0] _T_62276; // @[Modules.scala 143:103:@8153.4]
  wire [5:0] _T_62278; // @[Modules.scala 143:74:@8155.4]
  wire [5:0] _T_62280; // @[Modules.scala 144:80:@8156.4]
  wire [6:0] _T_62281; // @[Modules.scala 143:103:@8157.4]
  wire [5:0] _T_62282; // @[Modules.scala 143:103:@8158.4]
  wire [5:0] _T_62283; // @[Modules.scala 143:103:@8159.4]
  wire [5:0] _T_62285; // @[Modules.scala 143:74:@8161.4]
  wire [6:0] _T_62288; // @[Modules.scala 143:103:@8163.4]
  wire [5:0] _T_62289; // @[Modules.scala 143:103:@8164.4]
  wire [5:0] _T_62290; // @[Modules.scala 143:103:@8165.4]
  wire [4:0] _T_62294; // @[Modules.scala 144:80:@8168.4]
  wire [5:0] _GEN_215; // @[Modules.scala 143:103:@8169.4]
  wire [6:0] _T_62295; // @[Modules.scala 143:103:@8169.4]
  wire [5:0] _T_62296; // @[Modules.scala 143:103:@8170.4]
  wire [5:0] _T_62297; // @[Modules.scala 143:103:@8171.4]
  wire [4:0] _T_62299; // @[Modules.scala 143:74:@8173.4]
  wire [4:0] _T_62301; // @[Modules.scala 144:80:@8174.4]
  wire [5:0] _T_62302; // @[Modules.scala 143:103:@8175.4]
  wire [4:0] _T_62303; // @[Modules.scala 143:103:@8176.4]
  wire [4:0] _T_62304; // @[Modules.scala 143:103:@8177.4]
  wire [4:0] _T_62306; // @[Modules.scala 143:74:@8179.4]
  wire [4:0] _T_62308; // @[Modules.scala 144:80:@8180.4]
  wire [5:0] _T_62309; // @[Modules.scala 143:103:@8181.4]
  wire [4:0] _T_62310; // @[Modules.scala 143:103:@8182.4]
  wire [4:0] _T_62311; // @[Modules.scala 143:103:@8183.4]
  wire [4:0] _T_62313; // @[Modules.scala 143:74:@8185.4]
  wire [5:0] _T_62316; // @[Modules.scala 143:103:@8187.4]
  wire [4:0] _T_62317; // @[Modules.scala 143:103:@8188.4]
  wire [4:0] _T_62318; // @[Modules.scala 143:103:@8189.4]
  wire [4:0] _T_62320; // @[Modules.scala 143:74:@8191.4]
  wire [4:0] _T_62322; // @[Modules.scala 144:80:@8192.4]
  wire [5:0] _T_62323; // @[Modules.scala 143:103:@8193.4]
  wire [4:0] _T_62324; // @[Modules.scala 143:103:@8194.4]
  wire [4:0] _T_62325; // @[Modules.scala 143:103:@8195.4]
  wire [4:0] _T_62327; // @[Modules.scala 143:74:@8197.4]
  wire [5:0] _T_62330; // @[Modules.scala 143:103:@8199.4]
  wire [4:0] _T_62331; // @[Modules.scala 143:103:@8200.4]
  wire [4:0] _T_62332; // @[Modules.scala 143:103:@8201.4]
  wire [5:0] _GEN_216; // @[Modules.scala 143:103:@8205.4]
  wire [6:0] _T_62337; // @[Modules.scala 143:103:@8205.4]
  wire [5:0] _T_62338; // @[Modules.scala 143:103:@8206.4]
  wire [5:0] _T_62339; // @[Modules.scala 143:103:@8207.4]
  wire [5:0] _T_62344; // @[Modules.scala 143:103:@8211.4]
  wire [4:0] _T_62345; // @[Modules.scala 143:103:@8212.4]
  wire [4:0] _T_62346; // @[Modules.scala 143:103:@8213.4]
  wire [4:0] _T_62348; // @[Modules.scala 143:74:@8215.4]
  wire [4:0] _T_62350; // @[Modules.scala 144:80:@8216.4]
  wire [5:0] _T_62351; // @[Modules.scala 143:103:@8217.4]
  wire [4:0] _T_62352; // @[Modules.scala 143:103:@8218.4]
  wire [4:0] _T_62353; // @[Modules.scala 143:103:@8219.4]
  wire [4:0] _T_62362; // @[Modules.scala 143:74:@8227.4]
  wire [5:0] _T_62365; // @[Modules.scala 143:103:@8229.4]
  wire [4:0] _T_62366; // @[Modules.scala 143:103:@8230.4]
  wire [4:0] _T_62367; // @[Modules.scala 143:103:@8231.4]
  wire [4:0] _T_62371; // @[Modules.scala 144:80:@8234.4]
  wire [5:0] _T_62372; // @[Modules.scala 143:103:@8235.4]
  wire [4:0] _T_62373; // @[Modules.scala 143:103:@8236.4]
  wire [4:0] _T_62374; // @[Modules.scala 143:103:@8237.4]
  wire [4:0] _T_62376; // @[Modules.scala 143:74:@8239.4]
  wire [5:0] _T_62379; // @[Modules.scala 143:103:@8241.4]
  wire [4:0] _T_62380; // @[Modules.scala 143:103:@8242.4]
  wire [4:0] _T_62381; // @[Modules.scala 143:103:@8243.4]
  wire [4:0] _T_62385; // @[Modules.scala 144:80:@8246.4]
  wire [5:0] _T_62386; // @[Modules.scala 143:103:@8247.4]
  wire [4:0] _T_62387; // @[Modules.scala 143:103:@8248.4]
  wire [4:0] _T_62388; // @[Modules.scala 143:103:@8249.4]
  wire [4:0] _T_62390; // @[Modules.scala 143:74:@8251.4]
  wire [4:0] _T_62392; // @[Modules.scala 144:80:@8252.4]
  wire [5:0] _T_62393; // @[Modules.scala 143:103:@8253.4]
  wire [4:0] _T_62394; // @[Modules.scala 143:103:@8254.4]
  wire [4:0] _T_62395; // @[Modules.scala 143:103:@8255.4]
  wire [4:0] _T_62397; // @[Modules.scala 143:74:@8257.4]
  wire [4:0] _T_62399; // @[Modules.scala 144:80:@8258.4]
  wire [5:0] _T_62400; // @[Modules.scala 143:103:@8259.4]
  wire [4:0] _T_62401; // @[Modules.scala 143:103:@8260.4]
  wire [4:0] _T_62402; // @[Modules.scala 143:103:@8261.4]
  wire [4:0] _T_62404; // @[Modules.scala 143:74:@8263.4]
  wire [5:0] _GEN_217; // @[Modules.scala 143:103:@8265.4]
  wire [6:0] _T_62407; // @[Modules.scala 143:103:@8265.4]
  wire [5:0] _T_62408; // @[Modules.scala 143:103:@8266.4]
  wire [5:0] _T_62409; // @[Modules.scala 143:103:@8267.4]
  wire [6:0] _T_62414; // @[Modules.scala 143:103:@8271.4]
  wire [5:0] _T_62415; // @[Modules.scala 143:103:@8272.4]
  wire [5:0] _T_62416; // @[Modules.scala 143:103:@8273.4]
  wire [13:0] buffer_2_0; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62417; // @[Modules.scala 160:64:@8275.4]
  wire [13:0] _T_62418; // @[Modules.scala 160:64:@8276.4]
  wire [13:0] buffer_2_310; // @[Modules.scala 160:64:@8277.4]
  wire [13:0] buffer_2_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62420; // @[Modules.scala 160:64:@8279.4]
  wire [13:0] _T_62421; // @[Modules.scala 160:64:@8280.4]
  wire [13:0] buffer_2_311; // @[Modules.scala 160:64:@8281.4]
  wire [13:0] buffer_2_4; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_5; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62423; // @[Modules.scala 160:64:@8283.4]
  wire [13:0] _T_62424; // @[Modules.scala 160:64:@8284.4]
  wire [13:0] buffer_2_312; // @[Modules.scala 160:64:@8285.4]
  wire [13:0] buffer_2_6; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_7; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62426; // @[Modules.scala 160:64:@8287.4]
  wire [13:0] _T_62427; // @[Modules.scala 160:64:@8288.4]
  wire [13:0] buffer_2_313; // @[Modules.scala 160:64:@8289.4]
  wire [13:0] buffer_2_8; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62429; // @[Modules.scala 160:64:@8291.4]
  wire [13:0] _T_62430; // @[Modules.scala 160:64:@8292.4]
  wire [13:0] buffer_2_314; // @[Modules.scala 160:64:@8293.4]
  wire [13:0] buffer_2_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62432; // @[Modules.scala 160:64:@8295.4]
  wire [13:0] _T_62433; // @[Modules.scala 160:64:@8296.4]
  wire [13:0] buffer_2_315; // @[Modules.scala 160:64:@8297.4]
  wire [13:0] buffer_2_12; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62435; // @[Modules.scala 160:64:@8299.4]
  wire [13:0] _T_62436; // @[Modules.scala 160:64:@8300.4]
  wire [13:0] buffer_2_316; // @[Modules.scala 160:64:@8301.4]
  wire [13:0] buffer_2_14; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_15; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62438; // @[Modules.scala 160:64:@8303.4]
  wire [13:0] _T_62439; // @[Modules.scala 160:64:@8304.4]
  wire [13:0] buffer_2_317; // @[Modules.scala 160:64:@8305.4]
  wire [13:0] buffer_2_16; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_17; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62441; // @[Modules.scala 160:64:@8307.4]
  wire [13:0] _T_62442; // @[Modules.scala 160:64:@8308.4]
  wire [13:0] buffer_2_318; // @[Modules.scala 160:64:@8309.4]
  wire [14:0] _T_62444; // @[Modules.scala 160:64:@8311.4]
  wire [13:0] _T_62445; // @[Modules.scala 160:64:@8312.4]
  wire [13:0] buffer_2_319; // @[Modules.scala 160:64:@8313.4]
  wire [14:0] _T_62447; // @[Modules.scala 160:64:@8315.4]
  wire [13:0] _T_62448; // @[Modules.scala 160:64:@8316.4]
  wire [13:0] buffer_2_320; // @[Modules.scala 160:64:@8317.4]
  wire [13:0] buffer_2_22; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_23; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62450; // @[Modules.scala 160:64:@8319.4]
  wire [13:0] _T_62451; // @[Modules.scala 160:64:@8320.4]
  wire [13:0] buffer_2_321; // @[Modules.scala 160:64:@8321.4]
  wire [13:0] buffer_2_24; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62453; // @[Modules.scala 160:64:@8323.4]
  wire [13:0] _T_62454; // @[Modules.scala 160:64:@8324.4]
  wire [13:0] buffer_2_322; // @[Modules.scala 160:64:@8325.4]
  wire [13:0] buffer_2_26; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62456; // @[Modules.scala 160:64:@8327.4]
  wire [13:0] _T_62457; // @[Modules.scala 160:64:@8328.4]
  wire [13:0] buffer_2_323; // @[Modules.scala 160:64:@8329.4]
  wire [13:0] buffer_2_28; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_29; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62459; // @[Modules.scala 160:64:@8331.4]
  wire [13:0] _T_62460; // @[Modules.scala 160:64:@8332.4]
  wire [13:0] buffer_2_324; // @[Modules.scala 160:64:@8333.4]
  wire [13:0] buffer_2_30; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_31; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62462; // @[Modules.scala 160:64:@8335.4]
  wire [13:0] _T_62463; // @[Modules.scala 160:64:@8336.4]
  wire [13:0] buffer_2_325; // @[Modules.scala 160:64:@8337.4]
  wire [13:0] buffer_2_32; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62465; // @[Modules.scala 160:64:@8339.4]
  wire [13:0] _T_62466; // @[Modules.scala 160:64:@8340.4]
  wire [13:0] buffer_2_326; // @[Modules.scala 160:64:@8341.4]
  wire [13:0] buffer_2_34; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62468; // @[Modules.scala 160:64:@8343.4]
  wire [13:0] _T_62469; // @[Modules.scala 160:64:@8344.4]
  wire [13:0] buffer_2_327; // @[Modules.scala 160:64:@8345.4]
  wire [13:0] buffer_2_36; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_37; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62471; // @[Modules.scala 160:64:@8347.4]
  wire [13:0] _T_62472; // @[Modules.scala 160:64:@8348.4]
  wire [13:0] buffer_2_328; // @[Modules.scala 160:64:@8349.4]
  wire [13:0] buffer_2_38; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62474; // @[Modules.scala 160:64:@8351.4]
  wire [13:0] _T_62475; // @[Modules.scala 160:64:@8352.4]
  wire [13:0] buffer_2_329; // @[Modules.scala 160:64:@8353.4]
  wire [14:0] _T_62477; // @[Modules.scala 160:64:@8355.4]
  wire [13:0] _T_62478; // @[Modules.scala 160:64:@8356.4]
  wire [13:0] buffer_2_330; // @[Modules.scala 160:64:@8357.4]
  wire [13:0] buffer_2_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62480; // @[Modules.scala 160:64:@8359.4]
  wire [13:0] _T_62481; // @[Modules.scala 160:64:@8360.4]
  wire [13:0] buffer_2_331; // @[Modules.scala 160:64:@8361.4]
  wire [13:0] buffer_2_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62483; // @[Modules.scala 160:64:@8363.4]
  wire [13:0] _T_62484; // @[Modules.scala 160:64:@8364.4]
  wire [13:0] buffer_2_332; // @[Modules.scala 160:64:@8365.4]
  wire [13:0] buffer_2_46; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_47; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62486; // @[Modules.scala 160:64:@8367.4]
  wire [13:0] _T_62487; // @[Modules.scala 160:64:@8368.4]
  wire [13:0] buffer_2_333; // @[Modules.scala 160:64:@8369.4]
  wire [13:0] buffer_2_48; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62489; // @[Modules.scala 160:64:@8371.4]
  wire [13:0] _T_62490; // @[Modules.scala 160:64:@8372.4]
  wire [13:0] buffer_2_334; // @[Modules.scala 160:64:@8373.4]
  wire [13:0] buffer_2_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62492; // @[Modules.scala 160:64:@8375.4]
  wire [13:0] _T_62493; // @[Modules.scala 160:64:@8376.4]
  wire [13:0] buffer_2_335; // @[Modules.scala 160:64:@8377.4]
  wire [13:0] buffer_2_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62495; // @[Modules.scala 160:64:@8379.4]
  wire [13:0] _T_62496; // @[Modules.scala 160:64:@8380.4]
  wire [13:0] buffer_2_336; // @[Modules.scala 160:64:@8381.4]
  wire [13:0] buffer_2_54; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62498; // @[Modules.scala 160:64:@8383.4]
  wire [13:0] _T_62499; // @[Modules.scala 160:64:@8384.4]
  wire [13:0] buffer_2_337; // @[Modules.scala 160:64:@8385.4]
  wire [13:0] buffer_2_56; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62501; // @[Modules.scala 160:64:@8387.4]
  wire [13:0] _T_62502; // @[Modules.scala 160:64:@8388.4]
  wire [13:0] buffer_2_338; // @[Modules.scala 160:64:@8389.4]
  wire [13:0] buffer_2_58; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62504; // @[Modules.scala 160:64:@8391.4]
  wire [13:0] _T_62505; // @[Modules.scala 160:64:@8392.4]
  wire [13:0] buffer_2_339; // @[Modules.scala 160:64:@8393.4]
  wire [13:0] buffer_2_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62507; // @[Modules.scala 160:64:@8395.4]
  wire [13:0] _T_62508; // @[Modules.scala 160:64:@8396.4]
  wire [13:0] buffer_2_340; // @[Modules.scala 160:64:@8397.4]
  wire [13:0] buffer_2_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62510; // @[Modules.scala 160:64:@8399.4]
  wire [13:0] _T_62511; // @[Modules.scala 160:64:@8400.4]
  wire [13:0] buffer_2_341; // @[Modules.scala 160:64:@8401.4]
  wire [13:0] buffer_2_64; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62513; // @[Modules.scala 160:64:@8403.4]
  wire [13:0] _T_62514; // @[Modules.scala 160:64:@8404.4]
  wire [13:0] buffer_2_342; // @[Modules.scala 160:64:@8405.4]
  wire [13:0] buffer_2_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62516; // @[Modules.scala 160:64:@8407.4]
  wire [13:0] _T_62517; // @[Modules.scala 160:64:@8408.4]
  wire [13:0] buffer_2_343; // @[Modules.scala 160:64:@8409.4]
  wire [13:0] buffer_2_68; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62519; // @[Modules.scala 160:64:@8411.4]
  wire [13:0] _T_62520; // @[Modules.scala 160:64:@8412.4]
  wire [13:0] buffer_2_344; // @[Modules.scala 160:64:@8413.4]
  wire [13:0] buffer_2_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62522; // @[Modules.scala 160:64:@8415.4]
  wire [13:0] _T_62523; // @[Modules.scala 160:64:@8416.4]
  wire [13:0] buffer_2_345; // @[Modules.scala 160:64:@8417.4]
  wire [13:0] buffer_2_72; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62525; // @[Modules.scala 160:64:@8419.4]
  wire [13:0] _T_62526; // @[Modules.scala 160:64:@8420.4]
  wire [13:0] buffer_2_346; // @[Modules.scala 160:64:@8421.4]
  wire [13:0] buffer_2_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62528; // @[Modules.scala 160:64:@8423.4]
  wire [13:0] _T_62529; // @[Modules.scala 160:64:@8424.4]
  wire [13:0] buffer_2_347; // @[Modules.scala 160:64:@8425.4]
  wire [13:0] buffer_2_76; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62531; // @[Modules.scala 160:64:@8427.4]
  wire [13:0] _T_62532; // @[Modules.scala 160:64:@8428.4]
  wire [13:0] buffer_2_348; // @[Modules.scala 160:64:@8429.4]
  wire [13:0] buffer_2_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62537; // @[Modules.scala 160:64:@8435.4]
  wire [13:0] _T_62538; // @[Modules.scala 160:64:@8436.4]
  wire [13:0] buffer_2_350; // @[Modules.scala 160:64:@8437.4]
  wire [13:0] buffer_2_82; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_83; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62540; // @[Modules.scala 160:64:@8439.4]
  wire [13:0] _T_62541; // @[Modules.scala 160:64:@8440.4]
  wire [13:0] buffer_2_351; // @[Modules.scala 160:64:@8441.4]
  wire [13:0] buffer_2_84; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62543; // @[Modules.scala 160:64:@8443.4]
  wire [13:0] _T_62544; // @[Modules.scala 160:64:@8444.4]
  wire [13:0] buffer_2_352; // @[Modules.scala 160:64:@8445.4]
  wire [13:0] buffer_2_86; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_87; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62546; // @[Modules.scala 160:64:@8447.4]
  wire [13:0] _T_62547; // @[Modules.scala 160:64:@8448.4]
  wire [13:0] buffer_2_353; // @[Modules.scala 160:64:@8449.4]
  wire [13:0] buffer_2_88; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_89; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62549; // @[Modules.scala 160:64:@8451.4]
  wire [13:0] _T_62550; // @[Modules.scala 160:64:@8452.4]
  wire [13:0] buffer_2_354; // @[Modules.scala 160:64:@8453.4]
  wire [13:0] buffer_2_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62552; // @[Modules.scala 160:64:@8455.4]
  wire [13:0] _T_62553; // @[Modules.scala 160:64:@8456.4]
  wire [13:0] buffer_2_355; // @[Modules.scala 160:64:@8457.4]
  wire [13:0] buffer_2_92; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62555; // @[Modules.scala 160:64:@8459.4]
  wire [13:0] _T_62556; // @[Modules.scala 160:64:@8460.4]
  wire [13:0] buffer_2_356; // @[Modules.scala 160:64:@8461.4]
  wire [13:0] buffer_2_94; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62558; // @[Modules.scala 160:64:@8463.4]
  wire [13:0] _T_62559; // @[Modules.scala 160:64:@8464.4]
  wire [13:0] buffer_2_357; // @[Modules.scala 160:64:@8465.4]
  wire [13:0] buffer_2_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62561; // @[Modules.scala 160:64:@8467.4]
  wire [13:0] _T_62562; // @[Modules.scala 160:64:@8468.4]
  wire [13:0] buffer_2_358; // @[Modules.scala 160:64:@8469.4]
  wire [13:0] buffer_2_98; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_99; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62564; // @[Modules.scala 160:64:@8471.4]
  wire [13:0] _T_62565; // @[Modules.scala 160:64:@8472.4]
  wire [13:0] buffer_2_359; // @[Modules.scala 160:64:@8473.4]
  wire [14:0] _T_62567; // @[Modules.scala 160:64:@8475.4]
  wire [13:0] _T_62568; // @[Modules.scala 160:64:@8476.4]
  wire [13:0] buffer_2_360; // @[Modules.scala 160:64:@8477.4]
  wire [13:0] buffer_2_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62573; // @[Modules.scala 160:64:@8483.4]
  wire [13:0] _T_62574; // @[Modules.scala 160:64:@8484.4]
  wire [13:0] buffer_2_362; // @[Modules.scala 160:64:@8485.4]
  wire [13:0] buffer_2_106; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62576; // @[Modules.scala 160:64:@8487.4]
  wire [13:0] _T_62577; // @[Modules.scala 160:64:@8488.4]
  wire [13:0] buffer_2_363; // @[Modules.scala 160:64:@8489.4]
  wire [13:0] buffer_2_108; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_109; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62579; // @[Modules.scala 160:64:@8491.4]
  wire [13:0] _T_62580; // @[Modules.scala 160:64:@8492.4]
  wire [13:0] buffer_2_364; // @[Modules.scala 160:64:@8493.4]
  wire [13:0] buffer_2_110; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62582; // @[Modules.scala 160:64:@8495.4]
  wire [13:0] _T_62583; // @[Modules.scala 160:64:@8496.4]
  wire [13:0] buffer_2_365; // @[Modules.scala 160:64:@8497.4]
  wire [13:0] buffer_2_112; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62585; // @[Modules.scala 160:64:@8499.4]
  wire [13:0] _T_62586; // @[Modules.scala 160:64:@8500.4]
  wire [13:0] buffer_2_366; // @[Modules.scala 160:64:@8501.4]
  wire [13:0] buffer_2_116; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62591; // @[Modules.scala 160:64:@8507.4]
  wire [13:0] _T_62592; // @[Modules.scala 160:64:@8508.4]
  wire [13:0] buffer_2_368; // @[Modules.scala 160:64:@8509.4]
  wire [13:0] buffer_2_118; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_119; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62594; // @[Modules.scala 160:64:@8511.4]
  wire [13:0] _T_62595; // @[Modules.scala 160:64:@8512.4]
  wire [13:0] buffer_2_369; // @[Modules.scala 160:64:@8513.4]
  wire [13:0] buffer_2_120; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62597; // @[Modules.scala 160:64:@8515.4]
  wire [13:0] _T_62598; // @[Modules.scala 160:64:@8516.4]
  wire [13:0] buffer_2_370; // @[Modules.scala 160:64:@8517.4]
  wire [13:0] buffer_2_122; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62600; // @[Modules.scala 160:64:@8519.4]
  wire [13:0] _T_62601; // @[Modules.scala 160:64:@8520.4]
  wire [13:0] buffer_2_371; // @[Modules.scala 160:64:@8521.4]
  wire [13:0] buffer_2_124; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62603; // @[Modules.scala 160:64:@8523.4]
  wire [13:0] _T_62604; // @[Modules.scala 160:64:@8524.4]
  wire [13:0] buffer_2_372; // @[Modules.scala 160:64:@8525.4]
  wire [14:0] _T_62606; // @[Modules.scala 160:64:@8527.4]
  wire [13:0] _T_62607; // @[Modules.scala 160:64:@8528.4]
  wire [13:0] buffer_2_373; // @[Modules.scala 160:64:@8529.4]
  wire [13:0] buffer_2_128; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_129; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62609; // @[Modules.scala 160:64:@8531.4]
  wire [13:0] _T_62610; // @[Modules.scala 160:64:@8532.4]
  wire [13:0] buffer_2_374; // @[Modules.scala 160:64:@8533.4]
  wire [13:0] buffer_2_130; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62612; // @[Modules.scala 160:64:@8535.4]
  wire [13:0] _T_62613; // @[Modules.scala 160:64:@8536.4]
  wire [13:0] buffer_2_375; // @[Modules.scala 160:64:@8537.4]
  wire [13:0] buffer_2_132; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62615; // @[Modules.scala 160:64:@8539.4]
  wire [13:0] _T_62616; // @[Modules.scala 160:64:@8540.4]
  wire [13:0] buffer_2_376; // @[Modules.scala 160:64:@8541.4]
  wire [13:0] buffer_2_134; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62618; // @[Modules.scala 160:64:@8543.4]
  wire [13:0] _T_62619; // @[Modules.scala 160:64:@8544.4]
  wire [13:0] buffer_2_377; // @[Modules.scala 160:64:@8545.4]
  wire [13:0] buffer_2_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62621; // @[Modules.scala 160:64:@8547.4]
  wire [13:0] _T_62622; // @[Modules.scala 160:64:@8548.4]
  wire [13:0] buffer_2_378; // @[Modules.scala 160:64:@8549.4]
  wire [13:0] buffer_2_138; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_139; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62624; // @[Modules.scala 160:64:@8551.4]
  wire [13:0] _T_62625; // @[Modules.scala 160:64:@8552.4]
  wire [13:0] buffer_2_379; // @[Modules.scala 160:64:@8553.4]
  wire [13:0] buffer_2_140; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62627; // @[Modules.scala 160:64:@8555.4]
  wire [13:0] _T_62628; // @[Modules.scala 160:64:@8556.4]
  wire [13:0] buffer_2_380; // @[Modules.scala 160:64:@8557.4]
  wire [13:0] buffer_2_142; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_143; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62630; // @[Modules.scala 160:64:@8559.4]
  wire [13:0] _T_62631; // @[Modules.scala 160:64:@8560.4]
  wire [13:0] buffer_2_381; // @[Modules.scala 160:64:@8561.4]
  wire [13:0] buffer_2_144; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62633; // @[Modules.scala 160:64:@8563.4]
  wire [13:0] _T_62634; // @[Modules.scala 160:64:@8564.4]
  wire [13:0] buffer_2_382; // @[Modules.scala 160:64:@8565.4]
  wire [13:0] buffer_2_146; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62636; // @[Modules.scala 160:64:@8567.4]
  wire [13:0] _T_62637; // @[Modules.scala 160:64:@8568.4]
  wire [13:0] buffer_2_383; // @[Modules.scala 160:64:@8569.4]
  wire [13:0] buffer_2_148; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62639; // @[Modules.scala 160:64:@8571.4]
  wire [13:0] _T_62640; // @[Modules.scala 160:64:@8572.4]
  wire [13:0] buffer_2_384; // @[Modules.scala 160:64:@8573.4]
  wire [13:0] buffer_2_150; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62642; // @[Modules.scala 160:64:@8575.4]
  wire [13:0] _T_62643; // @[Modules.scala 160:64:@8576.4]
  wire [13:0] buffer_2_385; // @[Modules.scala 160:64:@8577.4]
  wire [13:0] buffer_2_152; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62645; // @[Modules.scala 160:64:@8579.4]
  wire [13:0] _T_62646; // @[Modules.scala 160:64:@8580.4]
  wire [13:0] buffer_2_386; // @[Modules.scala 160:64:@8581.4]
  wire [13:0] buffer_2_154; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62648; // @[Modules.scala 160:64:@8583.4]
  wire [13:0] _T_62649; // @[Modules.scala 160:64:@8584.4]
  wire [13:0] buffer_2_387; // @[Modules.scala 160:64:@8585.4]
  wire [13:0] buffer_2_156; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62651; // @[Modules.scala 160:64:@8587.4]
  wire [13:0] _T_62652; // @[Modules.scala 160:64:@8588.4]
  wire [13:0] buffer_2_388; // @[Modules.scala 160:64:@8589.4]
  wire [13:0] buffer_2_158; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62654; // @[Modules.scala 160:64:@8591.4]
  wire [13:0] _T_62655; // @[Modules.scala 160:64:@8592.4]
  wire [13:0] buffer_2_389; // @[Modules.scala 160:64:@8593.4]
  wire [13:0] buffer_2_160; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62657; // @[Modules.scala 160:64:@8595.4]
  wire [13:0] _T_62658; // @[Modules.scala 160:64:@8596.4]
  wire [13:0] buffer_2_390; // @[Modules.scala 160:64:@8597.4]
  wire [13:0] buffer_2_162; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_163; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62660; // @[Modules.scala 160:64:@8599.4]
  wire [13:0] _T_62661; // @[Modules.scala 160:64:@8600.4]
  wire [13:0] buffer_2_391; // @[Modules.scala 160:64:@8601.4]
  wire [13:0] buffer_2_164; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62663; // @[Modules.scala 160:64:@8603.4]
  wire [13:0] _T_62664; // @[Modules.scala 160:64:@8604.4]
  wire [13:0] buffer_2_392; // @[Modules.scala 160:64:@8605.4]
  wire [13:0] buffer_2_166; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62666; // @[Modules.scala 160:64:@8607.4]
  wire [13:0] _T_62667; // @[Modules.scala 160:64:@8608.4]
  wire [13:0] buffer_2_393; // @[Modules.scala 160:64:@8609.4]
  wire [13:0] buffer_2_168; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62669; // @[Modules.scala 160:64:@8611.4]
  wire [13:0] _T_62670; // @[Modules.scala 160:64:@8612.4]
  wire [13:0] buffer_2_394; // @[Modules.scala 160:64:@8613.4]
  wire [13:0] buffer_2_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62672; // @[Modules.scala 160:64:@8615.4]
  wire [13:0] _T_62673; // @[Modules.scala 160:64:@8616.4]
  wire [13:0] buffer_2_395; // @[Modules.scala 160:64:@8617.4]
  wire [13:0] buffer_2_172; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_173; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62675; // @[Modules.scala 160:64:@8619.4]
  wire [13:0] _T_62676; // @[Modules.scala 160:64:@8620.4]
  wire [13:0] buffer_2_396; // @[Modules.scala 160:64:@8621.4]
  wire [13:0] buffer_2_174; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62678; // @[Modules.scala 160:64:@8623.4]
  wire [13:0] _T_62679; // @[Modules.scala 160:64:@8624.4]
  wire [13:0] buffer_2_397; // @[Modules.scala 160:64:@8625.4]
  wire [13:0] buffer_2_176; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62681; // @[Modules.scala 160:64:@8627.4]
  wire [13:0] _T_62682; // @[Modules.scala 160:64:@8628.4]
  wire [13:0] buffer_2_398; // @[Modules.scala 160:64:@8629.4]
  wire [13:0] buffer_2_178; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_179; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62684; // @[Modules.scala 160:64:@8631.4]
  wire [13:0] _T_62685; // @[Modules.scala 160:64:@8632.4]
  wire [13:0] buffer_2_399; // @[Modules.scala 160:64:@8633.4]
  wire [13:0] buffer_2_180; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62687; // @[Modules.scala 160:64:@8635.4]
  wire [13:0] _T_62688; // @[Modules.scala 160:64:@8636.4]
  wire [13:0] buffer_2_400; // @[Modules.scala 160:64:@8637.4]
  wire [13:0] buffer_2_182; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62690; // @[Modules.scala 160:64:@8639.4]
  wire [13:0] _T_62691; // @[Modules.scala 160:64:@8640.4]
  wire [13:0] buffer_2_401; // @[Modules.scala 160:64:@8641.4]
  wire [13:0] buffer_2_184; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62693; // @[Modules.scala 160:64:@8643.4]
  wire [13:0] _T_62694; // @[Modules.scala 160:64:@8644.4]
  wire [13:0] buffer_2_402; // @[Modules.scala 160:64:@8645.4]
  wire [13:0] buffer_2_186; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_187; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62696; // @[Modules.scala 160:64:@8647.4]
  wire [13:0] _T_62697; // @[Modules.scala 160:64:@8648.4]
  wire [13:0] buffer_2_403; // @[Modules.scala 160:64:@8649.4]
  wire [13:0] buffer_2_188; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62699; // @[Modules.scala 160:64:@8651.4]
  wire [13:0] _T_62700; // @[Modules.scala 160:64:@8652.4]
  wire [13:0] buffer_2_404; // @[Modules.scala 160:64:@8653.4]
  wire [13:0] buffer_2_190; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62702; // @[Modules.scala 160:64:@8655.4]
  wire [13:0] _T_62703; // @[Modules.scala 160:64:@8656.4]
  wire [13:0] buffer_2_405; // @[Modules.scala 160:64:@8657.4]
  wire [13:0] buffer_2_192; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62705; // @[Modules.scala 160:64:@8659.4]
  wire [13:0] _T_62706; // @[Modules.scala 160:64:@8660.4]
  wire [13:0] buffer_2_406; // @[Modules.scala 160:64:@8661.4]
  wire [13:0] buffer_2_194; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62708; // @[Modules.scala 160:64:@8663.4]
  wire [13:0] _T_62709; // @[Modules.scala 160:64:@8664.4]
  wire [13:0] buffer_2_407; // @[Modules.scala 160:64:@8665.4]
  wire [13:0] buffer_2_196; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62711; // @[Modules.scala 160:64:@8667.4]
  wire [13:0] _T_62712; // @[Modules.scala 160:64:@8668.4]
  wire [13:0] buffer_2_408; // @[Modules.scala 160:64:@8669.4]
  wire [13:0] buffer_2_198; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62714; // @[Modules.scala 160:64:@8671.4]
  wire [13:0] _T_62715; // @[Modules.scala 160:64:@8672.4]
  wire [13:0] buffer_2_409; // @[Modules.scala 160:64:@8673.4]
  wire [13:0] buffer_2_200; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62717; // @[Modules.scala 160:64:@8675.4]
  wire [13:0] _T_62718; // @[Modules.scala 160:64:@8676.4]
  wire [13:0] buffer_2_410; // @[Modules.scala 160:64:@8677.4]
  wire [13:0] buffer_2_202; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62720; // @[Modules.scala 160:64:@8679.4]
  wire [13:0] _T_62721; // @[Modules.scala 160:64:@8680.4]
  wire [13:0] buffer_2_411; // @[Modules.scala 160:64:@8681.4]
  wire [13:0] buffer_2_204; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62723; // @[Modules.scala 160:64:@8683.4]
  wire [13:0] _T_62724; // @[Modules.scala 160:64:@8684.4]
  wire [13:0] buffer_2_412; // @[Modules.scala 160:64:@8685.4]
  wire [13:0] buffer_2_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62726; // @[Modules.scala 160:64:@8687.4]
  wire [13:0] _T_62727; // @[Modules.scala 160:64:@8688.4]
  wire [13:0] buffer_2_413; // @[Modules.scala 160:64:@8689.4]
  wire [13:0] buffer_2_208; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62729; // @[Modules.scala 160:64:@8691.4]
  wire [13:0] _T_62730; // @[Modules.scala 160:64:@8692.4]
  wire [13:0] buffer_2_414; // @[Modules.scala 160:64:@8693.4]
  wire [13:0] buffer_2_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62732; // @[Modules.scala 160:64:@8695.4]
  wire [13:0] _T_62733; // @[Modules.scala 160:64:@8696.4]
  wire [13:0] buffer_2_415; // @[Modules.scala 160:64:@8697.4]
  wire [13:0] buffer_2_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62735; // @[Modules.scala 160:64:@8699.4]
  wire [13:0] _T_62736; // @[Modules.scala 160:64:@8700.4]
  wire [13:0] buffer_2_416; // @[Modules.scala 160:64:@8701.4]
  wire [13:0] buffer_2_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62738; // @[Modules.scala 160:64:@8703.4]
  wire [13:0] _T_62739; // @[Modules.scala 160:64:@8704.4]
  wire [13:0] buffer_2_417; // @[Modules.scala 160:64:@8705.4]
  wire [13:0] buffer_2_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62741; // @[Modules.scala 160:64:@8707.4]
  wire [13:0] _T_62742; // @[Modules.scala 160:64:@8708.4]
  wire [13:0] buffer_2_418; // @[Modules.scala 160:64:@8709.4]
  wire [13:0] buffer_2_218; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62744; // @[Modules.scala 160:64:@8711.4]
  wire [13:0] _T_62745; // @[Modules.scala 160:64:@8712.4]
  wire [13:0] buffer_2_419; // @[Modules.scala 160:64:@8713.4]
  wire [13:0] buffer_2_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62750; // @[Modules.scala 160:64:@8719.4]
  wire [13:0] _T_62751; // @[Modules.scala 160:64:@8720.4]
  wire [13:0] buffer_2_421; // @[Modules.scala 160:64:@8721.4]
  wire [13:0] buffer_2_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62753; // @[Modules.scala 160:64:@8723.4]
  wire [13:0] _T_62754; // @[Modules.scala 160:64:@8724.4]
  wire [13:0] buffer_2_422; // @[Modules.scala 160:64:@8725.4]
  wire [13:0] buffer_2_226; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62756; // @[Modules.scala 160:64:@8727.4]
  wire [13:0] _T_62757; // @[Modules.scala 160:64:@8728.4]
  wire [13:0] buffer_2_423; // @[Modules.scala 160:64:@8729.4]
  wire [13:0] buffer_2_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62759; // @[Modules.scala 160:64:@8731.4]
  wire [13:0] _T_62760; // @[Modules.scala 160:64:@8732.4]
  wire [13:0] buffer_2_424; // @[Modules.scala 160:64:@8733.4]
  wire [13:0] buffer_2_230; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62762; // @[Modules.scala 160:64:@8735.4]
  wire [13:0] _T_62763; // @[Modules.scala 160:64:@8736.4]
  wire [13:0] buffer_2_425; // @[Modules.scala 160:64:@8737.4]
  wire [13:0] buffer_2_232; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62765; // @[Modules.scala 160:64:@8739.4]
  wire [13:0] _T_62766; // @[Modules.scala 160:64:@8740.4]
  wire [13:0] buffer_2_426; // @[Modules.scala 160:64:@8741.4]
  wire [13:0] buffer_2_234; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62768; // @[Modules.scala 160:64:@8743.4]
  wire [13:0] _T_62769; // @[Modules.scala 160:64:@8744.4]
  wire [13:0] buffer_2_427; // @[Modules.scala 160:64:@8745.4]
  wire [13:0] buffer_2_236; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62771; // @[Modules.scala 160:64:@8747.4]
  wire [13:0] _T_62772; // @[Modules.scala 160:64:@8748.4]
  wire [13:0] buffer_2_428; // @[Modules.scala 160:64:@8749.4]
  wire [13:0] buffer_2_238; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62774; // @[Modules.scala 160:64:@8751.4]
  wire [13:0] _T_62775; // @[Modules.scala 160:64:@8752.4]
  wire [13:0] buffer_2_429; // @[Modules.scala 160:64:@8753.4]
  wire [13:0] buffer_2_240; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62777; // @[Modules.scala 160:64:@8755.4]
  wire [13:0] _T_62778; // @[Modules.scala 160:64:@8756.4]
  wire [13:0] buffer_2_430; // @[Modules.scala 160:64:@8757.4]
  wire [13:0] buffer_2_242; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62780; // @[Modules.scala 160:64:@8759.4]
  wire [13:0] _T_62781; // @[Modules.scala 160:64:@8760.4]
  wire [13:0] buffer_2_431; // @[Modules.scala 160:64:@8761.4]
  wire [13:0] buffer_2_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62783; // @[Modules.scala 160:64:@8763.4]
  wire [13:0] _T_62784; // @[Modules.scala 160:64:@8764.4]
  wire [13:0] buffer_2_432; // @[Modules.scala 160:64:@8765.4]
  wire [13:0] buffer_2_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62786; // @[Modules.scala 160:64:@8767.4]
  wire [13:0] _T_62787; // @[Modules.scala 160:64:@8768.4]
  wire [13:0] buffer_2_433; // @[Modules.scala 160:64:@8769.4]
  wire [13:0] buffer_2_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62789; // @[Modules.scala 160:64:@8771.4]
  wire [13:0] _T_62790; // @[Modules.scala 160:64:@8772.4]
  wire [13:0] buffer_2_434; // @[Modules.scala 160:64:@8773.4]
  wire [13:0] buffer_2_250; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62792; // @[Modules.scala 160:64:@8775.4]
  wire [13:0] _T_62793; // @[Modules.scala 160:64:@8776.4]
  wire [13:0] buffer_2_435; // @[Modules.scala 160:64:@8777.4]
  wire [13:0] buffer_2_252; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62795; // @[Modules.scala 160:64:@8779.4]
  wire [13:0] _T_62796; // @[Modules.scala 160:64:@8780.4]
  wire [13:0] buffer_2_436; // @[Modules.scala 160:64:@8781.4]
  wire [13:0] buffer_2_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62798; // @[Modules.scala 160:64:@8783.4]
  wire [13:0] _T_62799; // @[Modules.scala 160:64:@8784.4]
  wire [13:0] buffer_2_437; // @[Modules.scala 160:64:@8785.4]
  wire [13:0] buffer_2_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62801; // @[Modules.scala 160:64:@8787.4]
  wire [13:0] _T_62802; // @[Modules.scala 160:64:@8788.4]
  wire [13:0] buffer_2_438; // @[Modules.scala 160:64:@8789.4]
  wire [13:0] buffer_2_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62804; // @[Modules.scala 160:64:@8791.4]
  wire [13:0] _T_62805; // @[Modules.scala 160:64:@8792.4]
  wire [13:0] buffer_2_439; // @[Modules.scala 160:64:@8793.4]
  wire [14:0] _T_62807; // @[Modules.scala 160:64:@8795.4]
  wire [13:0] _T_62808; // @[Modules.scala 160:64:@8796.4]
  wire [13:0] buffer_2_440; // @[Modules.scala 160:64:@8797.4]
  wire [14:0] _T_62810; // @[Modules.scala 160:64:@8799.4]
  wire [13:0] _T_62811; // @[Modules.scala 160:64:@8800.4]
  wire [13:0] buffer_2_441; // @[Modules.scala 160:64:@8801.4]
  wire [13:0] buffer_2_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62813; // @[Modules.scala 160:64:@8803.4]
  wire [13:0] _T_62814; // @[Modules.scala 160:64:@8804.4]
  wire [13:0] buffer_2_442; // @[Modules.scala 160:64:@8805.4]
  wire [13:0] buffer_2_266; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62816; // @[Modules.scala 160:64:@8807.4]
  wire [13:0] _T_62817; // @[Modules.scala 160:64:@8808.4]
  wire [13:0] buffer_2_443; // @[Modules.scala 160:64:@8809.4]
  wire [13:0] buffer_2_268; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62819; // @[Modules.scala 160:64:@8811.4]
  wire [13:0] _T_62820; // @[Modules.scala 160:64:@8812.4]
  wire [13:0] buffer_2_444; // @[Modules.scala 160:64:@8813.4]
  wire [13:0] buffer_2_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62822; // @[Modules.scala 160:64:@8815.4]
  wire [13:0] _T_62823; // @[Modules.scala 160:64:@8816.4]
  wire [13:0] buffer_2_445; // @[Modules.scala 160:64:@8817.4]
  wire [13:0] buffer_2_272; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62825; // @[Modules.scala 160:64:@8819.4]
  wire [13:0] _T_62826; // @[Modules.scala 160:64:@8820.4]
  wire [13:0] buffer_2_446; // @[Modules.scala 160:64:@8821.4]
  wire [14:0] _T_62828; // @[Modules.scala 160:64:@8823.4]
  wire [13:0] _T_62829; // @[Modules.scala 160:64:@8824.4]
  wire [13:0] buffer_2_447; // @[Modules.scala 160:64:@8825.4]
  wire [13:0] buffer_2_276; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_277; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62831; // @[Modules.scala 160:64:@8827.4]
  wire [13:0] _T_62832; // @[Modules.scala 160:64:@8828.4]
  wire [13:0] buffer_2_448; // @[Modules.scala 160:64:@8829.4]
  wire [13:0] buffer_2_278; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62834; // @[Modules.scala 160:64:@8831.4]
  wire [13:0] _T_62835; // @[Modules.scala 160:64:@8832.4]
  wire [13:0] buffer_2_449; // @[Modules.scala 160:64:@8833.4]
  wire [13:0] buffer_2_280; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62837; // @[Modules.scala 160:64:@8835.4]
  wire [13:0] _T_62838; // @[Modules.scala 160:64:@8836.4]
  wire [13:0] buffer_2_450; // @[Modules.scala 160:64:@8837.4]
  wire [13:0] buffer_2_282; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62840; // @[Modules.scala 160:64:@8839.4]
  wire [13:0] _T_62841; // @[Modules.scala 160:64:@8840.4]
  wire [13:0] buffer_2_451; // @[Modules.scala 160:64:@8841.4]
  wire [13:0] buffer_2_284; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_285; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62843; // @[Modules.scala 160:64:@8843.4]
  wire [13:0] _T_62844; // @[Modules.scala 160:64:@8844.4]
  wire [13:0] buffer_2_452; // @[Modules.scala 160:64:@8845.4]
  wire [13:0] buffer_2_286; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_287; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62846; // @[Modules.scala 160:64:@8847.4]
  wire [13:0] _T_62847; // @[Modules.scala 160:64:@8848.4]
  wire [13:0] buffer_2_453; // @[Modules.scala 160:64:@8849.4]
  wire [13:0] buffer_2_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62849; // @[Modules.scala 160:64:@8851.4]
  wire [13:0] _T_62850; // @[Modules.scala 160:64:@8852.4]
  wire [13:0] buffer_2_454; // @[Modules.scala 160:64:@8853.4]
  wire [13:0] buffer_2_290; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62852; // @[Modules.scala 160:64:@8855.4]
  wire [13:0] _T_62853; // @[Modules.scala 160:64:@8856.4]
  wire [13:0] buffer_2_455; // @[Modules.scala 160:64:@8857.4]
  wire [13:0] buffer_2_292; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62855; // @[Modules.scala 160:64:@8859.4]
  wire [13:0] _T_62856; // @[Modules.scala 160:64:@8860.4]
  wire [13:0] buffer_2_456; // @[Modules.scala 160:64:@8861.4]
  wire [13:0] buffer_2_294; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62858; // @[Modules.scala 160:64:@8863.4]
  wire [13:0] _T_62859; // @[Modules.scala 160:64:@8864.4]
  wire [13:0] buffer_2_457; // @[Modules.scala 160:64:@8865.4]
  wire [13:0] buffer_2_296; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_297; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62861; // @[Modules.scala 160:64:@8867.4]
  wire [13:0] _T_62862; // @[Modules.scala 160:64:@8868.4]
  wire [13:0] buffer_2_458; // @[Modules.scala 160:64:@8869.4]
  wire [13:0] buffer_2_298; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62864; // @[Modules.scala 160:64:@8871.4]
  wire [13:0] _T_62865; // @[Modules.scala 160:64:@8872.4]
  wire [13:0] buffer_2_459; // @[Modules.scala 160:64:@8873.4]
  wire [13:0] buffer_2_300; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62867; // @[Modules.scala 160:64:@8875.4]
  wire [13:0] _T_62868; // @[Modules.scala 160:64:@8876.4]
  wire [13:0] buffer_2_460; // @[Modules.scala 160:64:@8877.4]
  wire [13:0] buffer_2_302; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62870; // @[Modules.scala 160:64:@8879.4]
  wire [13:0] _T_62871; // @[Modules.scala 160:64:@8880.4]
  wire [13:0] buffer_2_461; // @[Modules.scala 160:64:@8881.4]
  wire [13:0] buffer_2_304; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_305; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62873; // @[Modules.scala 160:64:@8883.4]
  wire [13:0] _T_62874; // @[Modules.scala 160:64:@8884.4]
  wire [13:0] buffer_2_462; // @[Modules.scala 160:64:@8885.4]
  wire [13:0] buffer_2_306; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_307; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62876; // @[Modules.scala 160:64:@8887.4]
  wire [13:0] _T_62877; // @[Modules.scala 160:64:@8888.4]
  wire [13:0] buffer_2_463; // @[Modules.scala 160:64:@8889.4]
  wire [13:0] buffer_2_308; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_2_309; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_62879; // @[Modules.scala 160:64:@8891.4]
  wire [13:0] _T_62880; // @[Modules.scala 160:64:@8892.4]
  wire [13:0] buffer_2_464; // @[Modules.scala 160:64:@8893.4]
  wire [14:0] _T_62882; // @[Modules.scala 166:64:@8895.4]
  wire [13:0] _T_62883; // @[Modules.scala 166:64:@8896.4]
  wire [13:0] buffer_2_465; // @[Modules.scala 166:64:@8897.4]
  wire [14:0] _T_62885; // @[Modules.scala 166:64:@8899.4]
  wire [13:0] _T_62886; // @[Modules.scala 166:64:@8900.4]
  wire [13:0] buffer_2_466; // @[Modules.scala 166:64:@8901.4]
  wire [14:0] _T_62888; // @[Modules.scala 166:64:@8903.4]
  wire [13:0] _T_62889; // @[Modules.scala 166:64:@8904.4]
  wire [13:0] buffer_2_467; // @[Modules.scala 166:64:@8905.4]
  wire [14:0] _T_62891; // @[Modules.scala 166:64:@8907.4]
  wire [13:0] _T_62892; // @[Modules.scala 166:64:@8908.4]
  wire [13:0] buffer_2_468; // @[Modules.scala 166:64:@8909.4]
  wire [14:0] _T_62894; // @[Modules.scala 166:64:@8911.4]
  wire [13:0] _T_62895; // @[Modules.scala 166:64:@8912.4]
  wire [13:0] buffer_2_469; // @[Modules.scala 166:64:@8913.4]
  wire [14:0] _T_62897; // @[Modules.scala 166:64:@8915.4]
  wire [13:0] _T_62898; // @[Modules.scala 166:64:@8916.4]
  wire [13:0] buffer_2_470; // @[Modules.scala 166:64:@8917.4]
  wire [14:0] _T_62900; // @[Modules.scala 166:64:@8919.4]
  wire [13:0] _T_62901; // @[Modules.scala 166:64:@8920.4]
  wire [13:0] buffer_2_471; // @[Modules.scala 166:64:@8921.4]
  wire [14:0] _T_62903; // @[Modules.scala 166:64:@8923.4]
  wire [13:0] _T_62904; // @[Modules.scala 166:64:@8924.4]
  wire [13:0] buffer_2_472; // @[Modules.scala 166:64:@8925.4]
  wire [14:0] _T_62906; // @[Modules.scala 166:64:@8927.4]
  wire [13:0] _T_62907; // @[Modules.scala 166:64:@8928.4]
  wire [13:0] buffer_2_473; // @[Modules.scala 166:64:@8929.4]
  wire [14:0] _T_62909; // @[Modules.scala 166:64:@8931.4]
  wire [13:0] _T_62910; // @[Modules.scala 166:64:@8932.4]
  wire [13:0] buffer_2_474; // @[Modules.scala 166:64:@8933.4]
  wire [14:0] _T_62912; // @[Modules.scala 166:64:@8935.4]
  wire [13:0] _T_62913; // @[Modules.scala 166:64:@8936.4]
  wire [13:0] buffer_2_475; // @[Modules.scala 166:64:@8937.4]
  wire [14:0] _T_62915; // @[Modules.scala 166:64:@8939.4]
  wire [13:0] _T_62916; // @[Modules.scala 166:64:@8940.4]
  wire [13:0] buffer_2_476; // @[Modules.scala 166:64:@8941.4]
  wire [14:0] _T_62918; // @[Modules.scala 166:64:@8943.4]
  wire [13:0] _T_62919; // @[Modules.scala 166:64:@8944.4]
  wire [13:0] buffer_2_477; // @[Modules.scala 166:64:@8945.4]
  wire [14:0] _T_62921; // @[Modules.scala 166:64:@8947.4]
  wire [13:0] _T_62922; // @[Modules.scala 166:64:@8948.4]
  wire [13:0] buffer_2_478; // @[Modules.scala 166:64:@8949.4]
  wire [14:0] _T_62924; // @[Modules.scala 166:64:@8951.4]
  wire [13:0] _T_62925; // @[Modules.scala 166:64:@8952.4]
  wire [13:0] buffer_2_479; // @[Modules.scala 166:64:@8953.4]
  wire [14:0] _T_62927; // @[Modules.scala 166:64:@8955.4]
  wire [13:0] _T_62928; // @[Modules.scala 166:64:@8956.4]
  wire [13:0] buffer_2_480; // @[Modules.scala 166:64:@8957.4]
  wire [14:0] _T_62930; // @[Modules.scala 166:64:@8959.4]
  wire [13:0] _T_62931; // @[Modules.scala 166:64:@8960.4]
  wire [13:0] buffer_2_481; // @[Modules.scala 166:64:@8961.4]
  wire [14:0] _T_62933; // @[Modules.scala 166:64:@8963.4]
  wire [13:0] _T_62934; // @[Modules.scala 166:64:@8964.4]
  wire [13:0] buffer_2_482; // @[Modules.scala 166:64:@8965.4]
  wire [14:0] _T_62936; // @[Modules.scala 166:64:@8967.4]
  wire [13:0] _T_62937; // @[Modules.scala 166:64:@8968.4]
  wire [13:0] buffer_2_483; // @[Modules.scala 166:64:@8969.4]
  wire [14:0] _T_62939; // @[Modules.scala 166:64:@8971.4]
  wire [13:0] _T_62940; // @[Modules.scala 166:64:@8972.4]
  wire [13:0] buffer_2_484; // @[Modules.scala 166:64:@8973.4]
  wire [14:0] _T_62942; // @[Modules.scala 166:64:@8975.4]
  wire [13:0] _T_62943; // @[Modules.scala 166:64:@8976.4]
  wire [13:0] buffer_2_485; // @[Modules.scala 166:64:@8977.4]
  wire [14:0] _T_62945; // @[Modules.scala 166:64:@8979.4]
  wire [13:0] _T_62946; // @[Modules.scala 166:64:@8980.4]
  wire [13:0] buffer_2_486; // @[Modules.scala 166:64:@8981.4]
  wire [14:0] _T_62948; // @[Modules.scala 166:64:@8983.4]
  wire [13:0] _T_62949; // @[Modules.scala 166:64:@8984.4]
  wire [13:0] buffer_2_487; // @[Modules.scala 166:64:@8985.4]
  wire [14:0] _T_62951; // @[Modules.scala 166:64:@8987.4]
  wire [13:0] _T_62952; // @[Modules.scala 166:64:@8988.4]
  wire [13:0] buffer_2_488; // @[Modules.scala 166:64:@8989.4]
  wire [14:0] _T_62954; // @[Modules.scala 166:64:@8991.4]
  wire [13:0] _T_62955; // @[Modules.scala 166:64:@8992.4]
  wire [13:0] buffer_2_489; // @[Modules.scala 166:64:@8993.4]
  wire [14:0] _T_62957; // @[Modules.scala 166:64:@8995.4]
  wire [13:0] _T_62958; // @[Modules.scala 166:64:@8996.4]
  wire [13:0] buffer_2_490; // @[Modules.scala 166:64:@8997.4]
  wire [14:0] _T_62960; // @[Modules.scala 166:64:@8999.4]
  wire [13:0] _T_62961; // @[Modules.scala 166:64:@9000.4]
  wire [13:0] buffer_2_491; // @[Modules.scala 166:64:@9001.4]
  wire [14:0] _T_62963; // @[Modules.scala 166:64:@9003.4]
  wire [13:0] _T_62964; // @[Modules.scala 166:64:@9004.4]
  wire [13:0] buffer_2_492; // @[Modules.scala 166:64:@9005.4]
  wire [14:0] _T_62966; // @[Modules.scala 166:64:@9007.4]
  wire [13:0] _T_62967; // @[Modules.scala 166:64:@9008.4]
  wire [13:0] buffer_2_493; // @[Modules.scala 166:64:@9009.4]
  wire [14:0] _T_62969; // @[Modules.scala 166:64:@9011.4]
  wire [13:0] _T_62970; // @[Modules.scala 166:64:@9012.4]
  wire [13:0] buffer_2_494; // @[Modules.scala 166:64:@9013.4]
  wire [14:0] _T_62972; // @[Modules.scala 166:64:@9015.4]
  wire [13:0] _T_62973; // @[Modules.scala 166:64:@9016.4]
  wire [13:0] buffer_2_495; // @[Modules.scala 166:64:@9017.4]
  wire [14:0] _T_62975; // @[Modules.scala 166:64:@9019.4]
  wire [13:0] _T_62976; // @[Modules.scala 166:64:@9020.4]
  wire [13:0] buffer_2_496; // @[Modules.scala 166:64:@9021.4]
  wire [14:0] _T_62978; // @[Modules.scala 166:64:@9023.4]
  wire [13:0] _T_62979; // @[Modules.scala 166:64:@9024.4]
  wire [13:0] buffer_2_497; // @[Modules.scala 166:64:@9025.4]
  wire [14:0] _T_62981; // @[Modules.scala 166:64:@9027.4]
  wire [13:0] _T_62982; // @[Modules.scala 166:64:@9028.4]
  wire [13:0] buffer_2_498; // @[Modules.scala 166:64:@9029.4]
  wire [14:0] _T_62984; // @[Modules.scala 166:64:@9031.4]
  wire [13:0] _T_62985; // @[Modules.scala 166:64:@9032.4]
  wire [13:0] buffer_2_499; // @[Modules.scala 166:64:@9033.4]
  wire [14:0] _T_62987; // @[Modules.scala 166:64:@9035.4]
  wire [13:0] _T_62988; // @[Modules.scala 166:64:@9036.4]
  wire [13:0] buffer_2_500; // @[Modules.scala 166:64:@9037.4]
  wire [14:0] _T_62990; // @[Modules.scala 166:64:@9039.4]
  wire [13:0] _T_62991; // @[Modules.scala 166:64:@9040.4]
  wire [13:0] buffer_2_501; // @[Modules.scala 166:64:@9041.4]
  wire [14:0] _T_62993; // @[Modules.scala 166:64:@9043.4]
  wire [13:0] _T_62994; // @[Modules.scala 166:64:@9044.4]
  wire [13:0] buffer_2_502; // @[Modules.scala 166:64:@9045.4]
  wire [14:0] _T_62996; // @[Modules.scala 166:64:@9047.4]
  wire [13:0] _T_62997; // @[Modules.scala 166:64:@9048.4]
  wire [13:0] buffer_2_503; // @[Modules.scala 166:64:@9049.4]
  wire [14:0] _T_62999; // @[Modules.scala 166:64:@9051.4]
  wire [13:0] _T_63000; // @[Modules.scala 166:64:@9052.4]
  wire [13:0] buffer_2_504; // @[Modules.scala 166:64:@9053.4]
  wire [14:0] _T_63002; // @[Modules.scala 166:64:@9055.4]
  wire [13:0] _T_63003; // @[Modules.scala 166:64:@9056.4]
  wire [13:0] buffer_2_505; // @[Modules.scala 166:64:@9057.4]
  wire [14:0] _T_63005; // @[Modules.scala 166:64:@9059.4]
  wire [13:0] _T_63006; // @[Modules.scala 166:64:@9060.4]
  wire [13:0] buffer_2_506; // @[Modules.scala 166:64:@9061.4]
  wire [14:0] _T_63008; // @[Modules.scala 166:64:@9063.4]
  wire [13:0] _T_63009; // @[Modules.scala 166:64:@9064.4]
  wire [13:0] buffer_2_507; // @[Modules.scala 166:64:@9065.4]
  wire [14:0] _T_63011; // @[Modules.scala 166:64:@9067.4]
  wire [13:0] _T_63012; // @[Modules.scala 166:64:@9068.4]
  wire [13:0] buffer_2_508; // @[Modules.scala 166:64:@9069.4]
  wire [14:0] _T_63014; // @[Modules.scala 166:64:@9071.4]
  wire [13:0] _T_63015; // @[Modules.scala 166:64:@9072.4]
  wire [13:0] buffer_2_509; // @[Modules.scala 166:64:@9073.4]
  wire [14:0] _T_63017; // @[Modules.scala 166:64:@9075.4]
  wire [13:0] _T_63018; // @[Modules.scala 166:64:@9076.4]
  wire [13:0] buffer_2_510; // @[Modules.scala 166:64:@9077.4]
  wire [14:0] _T_63020; // @[Modules.scala 166:64:@9079.4]
  wire [13:0] _T_63021; // @[Modules.scala 166:64:@9080.4]
  wire [13:0] buffer_2_511; // @[Modules.scala 166:64:@9081.4]
  wire [14:0] _T_63023; // @[Modules.scala 166:64:@9083.4]
  wire [13:0] _T_63024; // @[Modules.scala 166:64:@9084.4]
  wire [13:0] buffer_2_512; // @[Modules.scala 166:64:@9085.4]
  wire [14:0] _T_63026; // @[Modules.scala 166:64:@9087.4]
  wire [13:0] _T_63027; // @[Modules.scala 166:64:@9088.4]
  wire [13:0] buffer_2_513; // @[Modules.scala 166:64:@9089.4]
  wire [14:0] _T_63029; // @[Modules.scala 166:64:@9091.4]
  wire [13:0] _T_63030; // @[Modules.scala 166:64:@9092.4]
  wire [13:0] buffer_2_514; // @[Modules.scala 166:64:@9093.4]
  wire [14:0] _T_63032; // @[Modules.scala 166:64:@9095.4]
  wire [13:0] _T_63033; // @[Modules.scala 166:64:@9096.4]
  wire [13:0] buffer_2_515; // @[Modules.scala 166:64:@9097.4]
  wire [14:0] _T_63035; // @[Modules.scala 166:64:@9099.4]
  wire [13:0] _T_63036; // @[Modules.scala 166:64:@9100.4]
  wire [13:0] buffer_2_516; // @[Modules.scala 166:64:@9101.4]
  wire [14:0] _T_63038; // @[Modules.scala 166:64:@9103.4]
  wire [13:0] _T_63039; // @[Modules.scala 166:64:@9104.4]
  wire [13:0] buffer_2_517; // @[Modules.scala 166:64:@9105.4]
  wire [14:0] _T_63041; // @[Modules.scala 166:64:@9107.4]
  wire [13:0] _T_63042; // @[Modules.scala 166:64:@9108.4]
  wire [13:0] buffer_2_518; // @[Modules.scala 166:64:@9109.4]
  wire [14:0] _T_63044; // @[Modules.scala 166:64:@9111.4]
  wire [13:0] _T_63045; // @[Modules.scala 166:64:@9112.4]
  wire [13:0] buffer_2_519; // @[Modules.scala 166:64:@9113.4]
  wire [14:0] _T_63047; // @[Modules.scala 166:64:@9115.4]
  wire [13:0] _T_63048; // @[Modules.scala 166:64:@9116.4]
  wire [13:0] buffer_2_520; // @[Modules.scala 166:64:@9117.4]
  wire [14:0] _T_63050; // @[Modules.scala 166:64:@9119.4]
  wire [13:0] _T_63051; // @[Modules.scala 166:64:@9120.4]
  wire [13:0] buffer_2_521; // @[Modules.scala 166:64:@9121.4]
  wire [14:0] _T_63053; // @[Modules.scala 166:64:@9123.4]
  wire [13:0] _T_63054; // @[Modules.scala 166:64:@9124.4]
  wire [13:0] buffer_2_522; // @[Modules.scala 166:64:@9125.4]
  wire [14:0] _T_63056; // @[Modules.scala 166:64:@9127.4]
  wire [13:0] _T_63057; // @[Modules.scala 166:64:@9128.4]
  wire [13:0] buffer_2_523; // @[Modules.scala 166:64:@9129.4]
  wire [14:0] _T_63059; // @[Modules.scala 166:64:@9131.4]
  wire [13:0] _T_63060; // @[Modules.scala 166:64:@9132.4]
  wire [13:0] buffer_2_524; // @[Modules.scala 166:64:@9133.4]
  wire [14:0] _T_63062; // @[Modules.scala 166:64:@9135.4]
  wire [13:0] _T_63063; // @[Modules.scala 166:64:@9136.4]
  wire [13:0] buffer_2_525; // @[Modules.scala 166:64:@9137.4]
  wire [14:0] _T_63065; // @[Modules.scala 166:64:@9139.4]
  wire [13:0] _T_63066; // @[Modules.scala 166:64:@9140.4]
  wire [13:0] buffer_2_526; // @[Modules.scala 166:64:@9141.4]
  wire [14:0] _T_63068; // @[Modules.scala 166:64:@9143.4]
  wire [13:0] _T_63069; // @[Modules.scala 166:64:@9144.4]
  wire [13:0] buffer_2_527; // @[Modules.scala 166:64:@9145.4]
  wire [14:0] _T_63071; // @[Modules.scala 166:64:@9147.4]
  wire [13:0] _T_63072; // @[Modules.scala 166:64:@9148.4]
  wire [13:0] buffer_2_528; // @[Modules.scala 166:64:@9149.4]
  wire [14:0] _T_63074; // @[Modules.scala 166:64:@9151.4]
  wire [13:0] _T_63075; // @[Modules.scala 166:64:@9152.4]
  wire [13:0] buffer_2_529; // @[Modules.scala 166:64:@9153.4]
  wire [14:0] _T_63077; // @[Modules.scala 166:64:@9155.4]
  wire [13:0] _T_63078; // @[Modules.scala 166:64:@9156.4]
  wire [13:0] buffer_2_530; // @[Modules.scala 166:64:@9157.4]
  wire [14:0] _T_63080; // @[Modules.scala 166:64:@9159.4]
  wire [13:0] _T_63081; // @[Modules.scala 166:64:@9160.4]
  wire [13:0] buffer_2_531; // @[Modules.scala 166:64:@9161.4]
  wire [14:0] _T_63083; // @[Modules.scala 166:64:@9163.4]
  wire [13:0] _T_63084; // @[Modules.scala 166:64:@9164.4]
  wire [13:0] buffer_2_532; // @[Modules.scala 166:64:@9165.4]
  wire [14:0] _T_63086; // @[Modules.scala 166:64:@9167.4]
  wire [13:0] _T_63087; // @[Modules.scala 166:64:@9168.4]
  wire [13:0] buffer_2_533; // @[Modules.scala 166:64:@9169.4]
  wire [14:0] _T_63089; // @[Modules.scala 166:64:@9171.4]
  wire [13:0] _T_63090; // @[Modules.scala 166:64:@9172.4]
  wire [13:0] buffer_2_534; // @[Modules.scala 166:64:@9173.4]
  wire [14:0] _T_63092; // @[Modules.scala 166:64:@9175.4]
  wire [13:0] _T_63093; // @[Modules.scala 166:64:@9176.4]
  wire [13:0] buffer_2_535; // @[Modules.scala 166:64:@9177.4]
  wire [14:0] _T_63095; // @[Modules.scala 166:64:@9179.4]
  wire [13:0] _T_63096; // @[Modules.scala 166:64:@9180.4]
  wire [13:0] buffer_2_536; // @[Modules.scala 166:64:@9181.4]
  wire [14:0] _T_63098; // @[Modules.scala 166:64:@9183.4]
  wire [13:0] _T_63099; // @[Modules.scala 166:64:@9184.4]
  wire [13:0] buffer_2_537; // @[Modules.scala 166:64:@9185.4]
  wire [14:0] _T_63101; // @[Modules.scala 166:64:@9187.4]
  wire [13:0] _T_63102; // @[Modules.scala 166:64:@9188.4]
  wire [13:0] buffer_2_538; // @[Modules.scala 166:64:@9189.4]
  wire [14:0] _T_63104; // @[Modules.scala 166:64:@9191.4]
  wire [13:0] _T_63105; // @[Modules.scala 166:64:@9192.4]
  wire [13:0] buffer_2_539; // @[Modules.scala 166:64:@9193.4]
  wire [14:0] _T_63107; // @[Modules.scala 166:64:@9195.4]
  wire [13:0] _T_63108; // @[Modules.scala 166:64:@9196.4]
  wire [13:0] buffer_2_540; // @[Modules.scala 166:64:@9197.4]
  wire [14:0] _T_63110; // @[Modules.scala 166:64:@9199.4]
  wire [13:0] _T_63111; // @[Modules.scala 166:64:@9200.4]
  wire [13:0] buffer_2_541; // @[Modules.scala 166:64:@9201.4]
  wire [14:0] _T_63113; // @[Modules.scala 166:64:@9203.4]
  wire [13:0] _T_63114; // @[Modules.scala 166:64:@9204.4]
  wire [13:0] buffer_2_542; // @[Modules.scala 166:64:@9205.4]
  wire [14:0] _T_63116; // @[Modules.scala 166:64:@9207.4]
  wire [13:0] _T_63117; // @[Modules.scala 166:64:@9208.4]
  wire [13:0] buffer_2_543; // @[Modules.scala 166:64:@9209.4]
  wire [14:0] _T_63119; // @[Modules.scala 166:64:@9211.4]
  wire [13:0] _T_63120; // @[Modules.scala 166:64:@9212.4]
  wire [13:0] buffer_2_544; // @[Modules.scala 166:64:@9213.4]
  wire [14:0] _T_63122; // @[Modules.scala 166:64:@9215.4]
  wire [13:0] _T_63123; // @[Modules.scala 166:64:@9216.4]
  wire [13:0] buffer_2_545; // @[Modules.scala 166:64:@9217.4]
  wire [14:0] _T_63125; // @[Modules.scala 166:64:@9219.4]
  wire [13:0] _T_63126; // @[Modules.scala 166:64:@9220.4]
  wire [13:0] buffer_2_546; // @[Modules.scala 166:64:@9221.4]
  wire [14:0] _T_63128; // @[Modules.scala 166:64:@9223.4]
  wire [13:0] _T_63129; // @[Modules.scala 166:64:@9224.4]
  wire [13:0] buffer_2_547; // @[Modules.scala 166:64:@9225.4]
  wire [14:0] _T_63131; // @[Modules.scala 166:64:@9227.4]
  wire [13:0] _T_63132; // @[Modules.scala 166:64:@9228.4]
  wire [13:0] buffer_2_548; // @[Modules.scala 166:64:@9229.4]
  wire [14:0] _T_63134; // @[Modules.scala 166:64:@9231.4]
  wire [13:0] _T_63135; // @[Modules.scala 166:64:@9232.4]
  wire [13:0] buffer_2_549; // @[Modules.scala 166:64:@9233.4]
  wire [14:0] _T_63137; // @[Modules.scala 166:64:@9235.4]
  wire [13:0] _T_63138; // @[Modules.scala 166:64:@9236.4]
  wire [13:0] buffer_2_550; // @[Modules.scala 166:64:@9237.4]
  wire [14:0] _T_63140; // @[Modules.scala 166:64:@9239.4]
  wire [13:0] _T_63141; // @[Modules.scala 166:64:@9240.4]
  wire [13:0] buffer_2_551; // @[Modules.scala 166:64:@9241.4]
  wire [14:0] _T_63143; // @[Modules.scala 166:64:@9243.4]
  wire [13:0] _T_63144; // @[Modules.scala 166:64:@9244.4]
  wire [13:0] buffer_2_552; // @[Modules.scala 166:64:@9245.4]
  wire [14:0] _T_63146; // @[Modules.scala 166:64:@9247.4]
  wire [13:0] _T_63147; // @[Modules.scala 166:64:@9248.4]
  wire [13:0] buffer_2_553; // @[Modules.scala 166:64:@9249.4]
  wire [14:0] _T_63149; // @[Modules.scala 166:64:@9251.4]
  wire [13:0] _T_63150; // @[Modules.scala 166:64:@9252.4]
  wire [13:0] buffer_2_554; // @[Modules.scala 166:64:@9253.4]
  wire [14:0] _T_63152; // @[Modules.scala 166:64:@9255.4]
  wire [13:0] _T_63153; // @[Modules.scala 166:64:@9256.4]
  wire [13:0] buffer_2_555; // @[Modules.scala 166:64:@9257.4]
  wire [14:0] _T_63155; // @[Modules.scala 166:64:@9259.4]
  wire [13:0] _T_63156; // @[Modules.scala 166:64:@9260.4]
  wire [13:0] buffer_2_556; // @[Modules.scala 166:64:@9261.4]
  wire [14:0] _T_63158; // @[Modules.scala 166:64:@9263.4]
  wire [13:0] _T_63159; // @[Modules.scala 166:64:@9264.4]
  wire [13:0] buffer_2_557; // @[Modules.scala 166:64:@9265.4]
  wire [14:0] _T_63161; // @[Modules.scala 166:64:@9267.4]
  wire [13:0] _T_63162; // @[Modules.scala 166:64:@9268.4]
  wire [13:0] buffer_2_558; // @[Modules.scala 166:64:@9269.4]
  wire [14:0] _T_63164; // @[Modules.scala 166:64:@9271.4]
  wire [13:0] _T_63165; // @[Modules.scala 166:64:@9272.4]
  wire [13:0] buffer_2_559; // @[Modules.scala 166:64:@9273.4]
  wire [14:0] _T_63167; // @[Modules.scala 166:64:@9275.4]
  wire [13:0] _T_63168; // @[Modules.scala 166:64:@9276.4]
  wire [13:0] buffer_2_560; // @[Modules.scala 166:64:@9277.4]
  wire [14:0] _T_63170; // @[Modules.scala 166:64:@9279.4]
  wire [13:0] _T_63171; // @[Modules.scala 166:64:@9280.4]
  wire [13:0] buffer_2_561; // @[Modules.scala 166:64:@9281.4]
  wire [14:0] _T_63173; // @[Modules.scala 166:64:@9283.4]
  wire [13:0] _T_63174; // @[Modules.scala 166:64:@9284.4]
  wire [13:0] buffer_2_562; // @[Modules.scala 166:64:@9285.4]
  wire [14:0] _T_63176; // @[Modules.scala 166:64:@9287.4]
  wire [13:0] _T_63177; // @[Modules.scala 166:64:@9288.4]
  wire [13:0] buffer_2_563; // @[Modules.scala 166:64:@9289.4]
  wire [14:0] _T_63179; // @[Modules.scala 166:64:@9291.4]
  wire [13:0] _T_63180; // @[Modules.scala 166:64:@9292.4]
  wire [13:0] buffer_2_564; // @[Modules.scala 166:64:@9293.4]
  wire [14:0] _T_63182; // @[Modules.scala 166:64:@9295.4]
  wire [13:0] _T_63183; // @[Modules.scala 166:64:@9296.4]
  wire [13:0] buffer_2_565; // @[Modules.scala 166:64:@9297.4]
  wire [14:0] _T_63185; // @[Modules.scala 166:64:@9299.4]
  wire [13:0] _T_63186; // @[Modules.scala 166:64:@9300.4]
  wire [13:0] buffer_2_566; // @[Modules.scala 166:64:@9301.4]
  wire [14:0] _T_63188; // @[Modules.scala 166:64:@9303.4]
  wire [13:0] _T_63189; // @[Modules.scala 166:64:@9304.4]
  wire [13:0] buffer_2_567; // @[Modules.scala 166:64:@9305.4]
  wire [14:0] _T_63191; // @[Modules.scala 166:64:@9307.4]
  wire [13:0] _T_63192; // @[Modules.scala 166:64:@9308.4]
  wire [13:0] buffer_2_568; // @[Modules.scala 166:64:@9309.4]
  wire [14:0] _T_63194; // @[Modules.scala 166:64:@9311.4]
  wire [13:0] _T_63195; // @[Modules.scala 166:64:@9312.4]
  wire [13:0] buffer_2_569; // @[Modules.scala 166:64:@9313.4]
  wire [14:0] _T_63197; // @[Modules.scala 166:64:@9315.4]
  wire [13:0] _T_63198; // @[Modules.scala 166:64:@9316.4]
  wire [13:0] buffer_2_570; // @[Modules.scala 166:64:@9317.4]
  wire [14:0] _T_63200; // @[Modules.scala 166:64:@9319.4]
  wire [13:0] _T_63201; // @[Modules.scala 166:64:@9320.4]
  wire [13:0] buffer_2_571; // @[Modules.scala 166:64:@9321.4]
  wire [14:0] _T_63203; // @[Modules.scala 166:64:@9323.4]
  wire [13:0] _T_63204; // @[Modules.scala 166:64:@9324.4]
  wire [13:0] buffer_2_572; // @[Modules.scala 166:64:@9325.4]
  wire [14:0] _T_63206; // @[Modules.scala 166:64:@9327.4]
  wire [13:0] _T_63207; // @[Modules.scala 166:64:@9328.4]
  wire [13:0] buffer_2_573; // @[Modules.scala 166:64:@9329.4]
  wire [14:0] _T_63209; // @[Modules.scala 166:64:@9331.4]
  wire [13:0] _T_63210; // @[Modules.scala 166:64:@9332.4]
  wire [13:0] buffer_2_574; // @[Modules.scala 166:64:@9333.4]
  wire [14:0] _T_63212; // @[Modules.scala 166:64:@9335.4]
  wire [13:0] _T_63213; // @[Modules.scala 166:64:@9336.4]
  wire [13:0] buffer_2_575; // @[Modules.scala 166:64:@9337.4]
  wire [14:0] _T_63215; // @[Modules.scala 166:64:@9339.4]
  wire [13:0] _T_63216; // @[Modules.scala 166:64:@9340.4]
  wire [13:0] buffer_2_576; // @[Modules.scala 166:64:@9341.4]
  wire [14:0] _T_63218; // @[Modules.scala 166:64:@9343.4]
  wire [13:0] _T_63219; // @[Modules.scala 166:64:@9344.4]
  wire [13:0] buffer_2_577; // @[Modules.scala 166:64:@9345.4]
  wire [14:0] _T_63221; // @[Modules.scala 166:64:@9347.4]
  wire [13:0] _T_63222; // @[Modules.scala 166:64:@9348.4]
  wire [13:0] buffer_2_578; // @[Modules.scala 166:64:@9349.4]
  wire [14:0] _T_63224; // @[Modules.scala 166:64:@9351.4]
  wire [13:0] _T_63225; // @[Modules.scala 166:64:@9352.4]
  wire [13:0] buffer_2_579; // @[Modules.scala 166:64:@9353.4]
  wire [14:0] _T_63227; // @[Modules.scala 172:66:@9355.4]
  wire [13:0] _T_63228; // @[Modules.scala 172:66:@9356.4]
  wire [13:0] buffer_2_580; // @[Modules.scala 172:66:@9357.4]
  wire [14:0] _T_63230; // @[Modules.scala 166:64:@9359.4]
  wire [13:0] _T_63231; // @[Modules.scala 166:64:@9360.4]
  wire [13:0] buffer_2_581; // @[Modules.scala 166:64:@9361.4]
  wire [14:0] _T_63233; // @[Modules.scala 166:64:@9363.4]
  wire [13:0] _T_63234; // @[Modules.scala 166:64:@9364.4]
  wire [13:0] buffer_2_582; // @[Modules.scala 166:64:@9365.4]
  wire [14:0] _T_63236; // @[Modules.scala 166:64:@9367.4]
  wire [13:0] _T_63237; // @[Modules.scala 166:64:@9368.4]
  wire [13:0] buffer_2_583; // @[Modules.scala 166:64:@9369.4]
  wire [14:0] _T_63239; // @[Modules.scala 166:64:@9371.4]
  wire [13:0] _T_63240; // @[Modules.scala 166:64:@9372.4]
  wire [13:0] buffer_2_584; // @[Modules.scala 166:64:@9373.4]
  wire [14:0] _T_63242; // @[Modules.scala 166:64:@9375.4]
  wire [13:0] _T_63243; // @[Modules.scala 166:64:@9376.4]
  wire [13:0] buffer_2_585; // @[Modules.scala 166:64:@9377.4]
  wire [14:0] _T_63245; // @[Modules.scala 166:64:@9379.4]
  wire [13:0] _T_63246; // @[Modules.scala 166:64:@9380.4]
  wire [13:0] buffer_2_586; // @[Modules.scala 166:64:@9381.4]
  wire [14:0] _T_63248; // @[Modules.scala 166:64:@9383.4]
  wire [13:0] _T_63249; // @[Modules.scala 166:64:@9384.4]
  wire [13:0] buffer_2_587; // @[Modules.scala 166:64:@9385.4]
  wire [14:0] _T_63251; // @[Modules.scala 166:64:@9387.4]
  wire [13:0] _T_63252; // @[Modules.scala 166:64:@9388.4]
  wire [13:0] buffer_2_588; // @[Modules.scala 166:64:@9389.4]
  wire [14:0] _T_63254; // @[Modules.scala 166:64:@9391.4]
  wire [13:0] _T_63255; // @[Modules.scala 166:64:@9392.4]
  wire [13:0] buffer_2_589; // @[Modules.scala 166:64:@9393.4]
  wire [14:0] _T_63257; // @[Modules.scala 166:64:@9395.4]
  wire [13:0] _T_63258; // @[Modules.scala 166:64:@9396.4]
  wire [13:0] buffer_2_590; // @[Modules.scala 166:64:@9397.4]
  wire [14:0] _T_63260; // @[Modules.scala 166:64:@9399.4]
  wire [13:0] _T_63261; // @[Modules.scala 166:64:@9400.4]
  wire [13:0] buffer_2_591; // @[Modules.scala 166:64:@9401.4]
  wire [14:0] _T_63263; // @[Modules.scala 166:64:@9403.4]
  wire [13:0] _T_63264; // @[Modules.scala 166:64:@9404.4]
  wire [13:0] buffer_2_592; // @[Modules.scala 166:64:@9405.4]
  wire [14:0] _T_63266; // @[Modules.scala 166:64:@9407.4]
  wire [13:0] _T_63267; // @[Modules.scala 166:64:@9408.4]
  wire [13:0] buffer_2_593; // @[Modules.scala 166:64:@9409.4]
  wire [14:0] _T_63269; // @[Modules.scala 166:64:@9411.4]
  wire [13:0] _T_63270; // @[Modules.scala 166:64:@9412.4]
  wire [13:0] buffer_2_594; // @[Modules.scala 166:64:@9413.4]
  wire [14:0] _T_63272; // @[Modules.scala 166:64:@9415.4]
  wire [13:0] _T_63273; // @[Modules.scala 166:64:@9416.4]
  wire [13:0] buffer_2_595; // @[Modules.scala 166:64:@9417.4]
  wire [14:0] _T_63275; // @[Modules.scala 166:64:@9419.4]
  wire [13:0] _T_63276; // @[Modules.scala 166:64:@9420.4]
  wire [13:0] buffer_2_596; // @[Modules.scala 166:64:@9421.4]
  wire [14:0] _T_63278; // @[Modules.scala 166:64:@9423.4]
  wire [13:0] _T_63279; // @[Modules.scala 166:64:@9424.4]
  wire [13:0] buffer_2_597; // @[Modules.scala 166:64:@9425.4]
  wire [14:0] _T_63281; // @[Modules.scala 166:64:@9427.4]
  wire [13:0] _T_63282; // @[Modules.scala 166:64:@9428.4]
  wire [13:0] buffer_2_598; // @[Modules.scala 166:64:@9429.4]
  wire [14:0] _T_63284; // @[Modules.scala 166:64:@9431.4]
  wire [13:0] _T_63285; // @[Modules.scala 166:64:@9432.4]
  wire [13:0] buffer_2_599; // @[Modules.scala 166:64:@9433.4]
  wire [14:0] _T_63287; // @[Modules.scala 166:64:@9435.4]
  wire [13:0] _T_63288; // @[Modules.scala 166:64:@9436.4]
  wire [13:0] buffer_2_600; // @[Modules.scala 166:64:@9437.4]
  wire [14:0] _T_63290; // @[Modules.scala 166:64:@9439.4]
  wire [13:0] _T_63291; // @[Modules.scala 166:64:@9440.4]
  wire [13:0] buffer_2_601; // @[Modules.scala 166:64:@9441.4]
  wire [14:0] _T_63293; // @[Modules.scala 166:64:@9443.4]
  wire [13:0] _T_63294; // @[Modules.scala 166:64:@9444.4]
  wire [13:0] buffer_2_602; // @[Modules.scala 166:64:@9445.4]
  wire [14:0] _T_63296; // @[Modules.scala 166:64:@9447.4]
  wire [13:0] _T_63297; // @[Modules.scala 166:64:@9448.4]
  wire [13:0] buffer_2_603; // @[Modules.scala 166:64:@9449.4]
  wire [14:0] _T_63299; // @[Modules.scala 166:64:@9451.4]
  wire [13:0] _T_63300; // @[Modules.scala 166:64:@9452.4]
  wire [13:0] buffer_2_604; // @[Modules.scala 166:64:@9453.4]
  wire [14:0] _T_63302; // @[Modules.scala 166:64:@9455.4]
  wire [13:0] _T_63303; // @[Modules.scala 166:64:@9456.4]
  wire [13:0] buffer_2_605; // @[Modules.scala 166:64:@9457.4]
  wire [14:0] _T_63305; // @[Modules.scala 166:64:@9459.4]
  wire [13:0] _T_63306; // @[Modules.scala 166:64:@9460.4]
  wire [13:0] buffer_2_606; // @[Modules.scala 166:64:@9461.4]
  wire [14:0] _T_63308; // @[Modules.scala 166:64:@9463.4]
  wire [13:0] _T_63309; // @[Modules.scala 166:64:@9464.4]
  wire [13:0] buffer_2_607; // @[Modules.scala 166:64:@9465.4]
  wire [14:0] _T_63311; // @[Modules.scala 166:64:@9467.4]
  wire [13:0] _T_63312; // @[Modules.scala 166:64:@9468.4]
  wire [13:0] buffer_2_608; // @[Modules.scala 166:64:@9469.4]
  wire [14:0] _T_63314; // @[Modules.scala 172:66:@9471.4]
  wire [13:0] _T_63315; // @[Modules.scala 172:66:@9472.4]
  wire [13:0] buffer_2_609; // @[Modules.scala 172:66:@9473.4]
  wire [14:0] _T_63317; // @[Modules.scala 160:64:@9475.4]
  wire [13:0] _T_63318; // @[Modules.scala 160:64:@9476.4]
  wire [13:0] buffer_2_610; // @[Modules.scala 160:64:@9477.4]
  wire [14:0] _T_63320; // @[Modules.scala 160:64:@9479.4]
  wire [13:0] _T_63321; // @[Modules.scala 160:64:@9480.4]
  wire [13:0] buffer_2_611; // @[Modules.scala 160:64:@9481.4]
  wire [14:0] _T_63323; // @[Modules.scala 160:64:@9483.4]
  wire [13:0] _T_63324; // @[Modules.scala 160:64:@9484.4]
  wire [13:0] buffer_2_612; // @[Modules.scala 160:64:@9485.4]
  wire [14:0] _T_63326; // @[Modules.scala 160:64:@9487.4]
  wire [13:0] _T_63327; // @[Modules.scala 160:64:@9488.4]
  wire [13:0] buffer_2_613; // @[Modules.scala 160:64:@9489.4]
  wire [14:0] _T_63329; // @[Modules.scala 160:64:@9491.4]
  wire [13:0] _T_63330; // @[Modules.scala 160:64:@9492.4]
  wire [13:0] buffer_2_614; // @[Modules.scala 160:64:@9493.4]
  wire [14:0] _T_63332; // @[Modules.scala 166:64:@9495.4]
  wire [13:0] _T_63333; // @[Modules.scala 166:64:@9496.4]
  wire [13:0] buffer_2_615; // @[Modules.scala 166:64:@9497.4]
  wire [14:0] _T_63335; // @[Modules.scala 166:64:@9499.4]
  wire [13:0] _T_63336; // @[Modules.scala 166:64:@9500.4]
  wire [13:0] buffer_2_616; // @[Modules.scala 166:64:@9501.4]
  wire [14:0] _T_63338; // @[Modules.scala 160:64:@9503.4]
  wire [13:0] _T_63339; // @[Modules.scala 160:64:@9504.4]
  wire [13:0] buffer_2_617; // @[Modules.scala 160:64:@9505.4]
  wire [14:0] _T_63341; // @[Modules.scala 172:66:@9507.4]
  wire [13:0] _T_63342; // @[Modules.scala 172:66:@9508.4]
  wire [13:0] buffer_2_618; // @[Modules.scala 172:66:@9509.4]
  wire [6:0] _T_63362; // @[Modules.scala 150:103:@9690.4]
  wire [5:0] _T_63363; // @[Modules.scala 150:103:@9691.4]
  wire [5:0] _T_63364; // @[Modules.scala 150:103:@9692.4]
  wire [4:0] _T_63375; // @[Modules.scala 151:80:@9701.4]
  wire [5:0] _T_63376; // @[Modules.scala 150:103:@9702.4]
  wire [4:0] _T_63377; // @[Modules.scala 150:103:@9703.4]
  wire [4:0] _T_63378; // @[Modules.scala 150:103:@9704.4]
  wire [5:0] _GEN_218; // @[Modules.scala 150:103:@9714.4]
  wire [6:0] _T_63390; // @[Modules.scala 150:103:@9714.4]
  wire [5:0] _T_63391; // @[Modules.scala 150:103:@9715.4]
  wire [5:0] _T_63392; // @[Modules.scala 150:103:@9716.4]
  wire [5:0] _T_63397; // @[Modules.scala 150:103:@9720.4]
  wire [4:0] _T_63398; // @[Modules.scala 150:103:@9721.4]
  wire [4:0] _T_63399; // @[Modules.scala 150:103:@9722.4]
  wire [4:0] _T_63403; // @[Modules.scala 151:80:@9725.4]
  wire [5:0] _T_63404; // @[Modules.scala 150:103:@9726.4]
  wire [4:0] _T_63405; // @[Modules.scala 150:103:@9727.4]
  wire [4:0] _T_63406; // @[Modules.scala 150:103:@9728.4]
  wire [4:0] _T_63408; // @[Modules.scala 150:74:@9730.4]
  wire [5:0] _T_63411; // @[Modules.scala 150:103:@9732.4]
  wire [4:0] _T_63412; // @[Modules.scala 150:103:@9733.4]
  wire [4:0] _T_63413; // @[Modules.scala 150:103:@9734.4]
  wire [6:0] _T_63418; // @[Modules.scala 150:103:@9738.4]
  wire [5:0] _T_63419; // @[Modules.scala 150:103:@9739.4]
  wire [5:0] _T_63420; // @[Modules.scala 150:103:@9740.4]
  wire [4:0] _T_63422; // @[Modules.scala 150:74:@9742.4]
  wire [5:0] _T_63425; // @[Modules.scala 150:103:@9744.4]
  wire [4:0] _T_63426; // @[Modules.scala 150:103:@9745.4]
  wire [4:0] _T_63427; // @[Modules.scala 150:103:@9746.4]
  wire [5:0] _T_63429; // @[Modules.scala 150:74:@9748.4]
  wire [6:0] _T_63432; // @[Modules.scala 150:103:@9750.4]
  wire [5:0] _T_63433; // @[Modules.scala 150:103:@9751.4]
  wire [5:0] _T_63434; // @[Modules.scala 150:103:@9752.4]
  wire [5:0] _GEN_220; // @[Modules.scala 150:103:@9756.4]
  wire [6:0] _T_63439; // @[Modules.scala 150:103:@9756.4]
  wire [5:0] _T_63440; // @[Modules.scala 150:103:@9757.4]
  wire [5:0] _T_63441; // @[Modules.scala 150:103:@9758.4]
  wire [5:0] _T_63467; // @[Modules.scala 150:103:@9780.4]
  wire [4:0] _T_63468; // @[Modules.scala 150:103:@9781.4]
  wire [4:0] _T_63469; // @[Modules.scala 150:103:@9782.4]
  wire [5:0] _GEN_221; // @[Modules.scala 150:103:@9786.4]
  wire [6:0] _T_63474; // @[Modules.scala 150:103:@9786.4]
  wire [5:0] _T_63475; // @[Modules.scala 150:103:@9787.4]
  wire [5:0] _T_63476; // @[Modules.scala 150:103:@9788.4]
  wire [4:0] _T_63485; // @[Modules.scala 150:74:@9796.4]
  wire [4:0] _T_63487; // @[Modules.scala 151:80:@9797.4]
  wire [5:0] _T_63488; // @[Modules.scala 150:103:@9798.4]
  wire [4:0] _T_63489; // @[Modules.scala 150:103:@9799.4]
  wire [4:0] _T_63490; // @[Modules.scala 150:103:@9800.4]
  wire [4:0] _T_63492; // @[Modules.scala 150:74:@9802.4]
  wire [5:0] _T_63495; // @[Modules.scala 150:103:@9804.4]
  wire [4:0] _T_63496; // @[Modules.scala 150:103:@9805.4]
  wire [4:0] _T_63497; // @[Modules.scala 150:103:@9806.4]
  wire [4:0] _T_63499; // @[Modules.scala 150:74:@9808.4]
  wire [5:0] _T_63502; // @[Modules.scala 150:103:@9810.4]
  wire [4:0] _T_63503; // @[Modules.scala 150:103:@9811.4]
  wire [4:0] _T_63504; // @[Modules.scala 150:103:@9812.4]
  wire [5:0] _T_63509; // @[Modules.scala 150:103:@9816.4]
  wire [4:0] _T_63510; // @[Modules.scala 150:103:@9817.4]
  wire [4:0] _T_63511; // @[Modules.scala 150:103:@9818.4]
  wire [5:0] _T_63516; // @[Modules.scala 150:103:@9822.4]
  wire [4:0] _T_63517; // @[Modules.scala 150:103:@9823.4]
  wire [4:0] _T_63518; // @[Modules.scala 150:103:@9824.4]
  wire [5:0] _T_63523; // @[Modules.scala 150:103:@9828.4]
  wire [4:0] _T_63524; // @[Modules.scala 150:103:@9829.4]
  wire [4:0] _T_63525; // @[Modules.scala 150:103:@9830.4]
  wire [5:0] _T_63530; // @[Modules.scala 150:103:@9834.4]
  wire [4:0] _T_63531; // @[Modules.scala 150:103:@9835.4]
  wire [4:0] _T_63532; // @[Modules.scala 150:103:@9836.4]
  wire [5:0] _T_63537; // @[Modules.scala 150:103:@9840.4]
  wire [4:0] _T_63538; // @[Modules.scala 150:103:@9841.4]
  wire [4:0] _T_63539; // @[Modules.scala 150:103:@9842.4]
  wire [4:0] _T_63541; // @[Modules.scala 150:74:@9844.4]
  wire [4:0] _T_63543; // @[Modules.scala 151:80:@9845.4]
  wire [5:0] _T_63544; // @[Modules.scala 150:103:@9846.4]
  wire [4:0] _T_63545; // @[Modules.scala 150:103:@9847.4]
  wire [4:0] _T_63546; // @[Modules.scala 150:103:@9848.4]
  wire [5:0] _T_63551; // @[Modules.scala 150:103:@9852.4]
  wire [4:0] _T_63552; // @[Modules.scala 150:103:@9853.4]
  wire [4:0] _T_63553; // @[Modules.scala 150:103:@9854.4]
  wire [5:0] _T_63558; // @[Modules.scala 150:103:@9858.4]
  wire [4:0] _T_63559; // @[Modules.scala 150:103:@9859.4]
  wire [4:0] _T_63560; // @[Modules.scala 150:103:@9860.4]
  wire [5:0] _GEN_222; // @[Modules.scala 150:103:@9864.4]
  wire [6:0] _T_63565; // @[Modules.scala 150:103:@9864.4]
  wire [5:0] _T_63566; // @[Modules.scala 150:103:@9865.4]
  wire [5:0] _T_63567; // @[Modules.scala 150:103:@9866.4]
  wire [4:0] _T_63571; // @[Modules.scala 151:80:@9869.4]
  wire [5:0] _T_63572; // @[Modules.scala 150:103:@9870.4]
  wire [4:0] _T_63573; // @[Modules.scala 150:103:@9871.4]
  wire [4:0] _T_63574; // @[Modules.scala 150:103:@9872.4]
  wire [4:0] _T_63585; // @[Modules.scala 151:80:@9881.4]
  wire [5:0] _T_63586; // @[Modules.scala 150:103:@9882.4]
  wire [4:0] _T_63587; // @[Modules.scala 150:103:@9883.4]
  wire [4:0] _T_63588; // @[Modules.scala 150:103:@9884.4]
  wire [4:0] _T_63590; // @[Modules.scala 150:74:@9886.4]
  wire [5:0] _T_63593; // @[Modules.scala 150:103:@9888.4]
  wire [4:0] _T_63594; // @[Modules.scala 150:103:@9889.4]
  wire [4:0] _T_63595; // @[Modules.scala 150:103:@9890.4]
  wire [4:0] _T_63599; // @[Modules.scala 151:80:@9893.4]
  wire [5:0] _T_63600; // @[Modules.scala 150:103:@9894.4]
  wire [4:0] _T_63601; // @[Modules.scala 150:103:@9895.4]
  wire [4:0] _T_63602; // @[Modules.scala 150:103:@9896.4]
  wire [4:0] _T_63604; // @[Modules.scala 150:74:@9898.4]
  wire [4:0] _T_63606; // @[Modules.scala 151:80:@9899.4]
  wire [5:0] _T_63607; // @[Modules.scala 150:103:@9900.4]
  wire [4:0] _T_63608; // @[Modules.scala 150:103:@9901.4]
  wire [4:0] _T_63609; // @[Modules.scala 150:103:@9902.4]
  wire [5:0] _T_63614; // @[Modules.scala 150:103:@9906.4]
  wire [4:0] _T_63615; // @[Modules.scala 150:103:@9907.4]
  wire [4:0] _T_63616; // @[Modules.scala 150:103:@9908.4]
  wire [5:0] _T_63621; // @[Modules.scala 150:103:@9912.4]
  wire [4:0] _T_63622; // @[Modules.scala 150:103:@9913.4]
  wire [4:0] _T_63623; // @[Modules.scala 150:103:@9914.4]
  wire [5:0] _GEN_223; // @[Modules.scala 150:103:@9918.4]
  wire [6:0] _T_63628; // @[Modules.scala 150:103:@9918.4]
  wire [5:0] _T_63629; // @[Modules.scala 150:103:@9919.4]
  wire [5:0] _T_63630; // @[Modules.scala 150:103:@9920.4]
  wire [6:0] _T_63635; // @[Modules.scala 150:103:@9924.4]
  wire [5:0] _T_63636; // @[Modules.scala 150:103:@9925.4]
  wire [5:0] _T_63637; // @[Modules.scala 150:103:@9926.4]
  wire [6:0] _T_63649; // @[Modules.scala 150:103:@9936.4]
  wire [5:0] _T_63650; // @[Modules.scala 150:103:@9937.4]
  wire [5:0] _T_63651; // @[Modules.scala 150:103:@9938.4]
  wire [6:0] _T_63656; // @[Modules.scala 150:103:@9942.4]
  wire [5:0] _T_63657; // @[Modules.scala 150:103:@9943.4]
  wire [5:0] _T_63658; // @[Modules.scala 150:103:@9944.4]
  wire [6:0] _T_63663; // @[Modules.scala 150:103:@9948.4]
  wire [5:0] _T_63664; // @[Modules.scala 150:103:@9949.4]
  wire [5:0] _T_63665; // @[Modules.scala 150:103:@9950.4]
  wire [4:0] _T_63669; // @[Modules.scala 151:80:@9953.4]
  wire [5:0] _T_63670; // @[Modules.scala 150:103:@9954.4]
  wire [4:0] _T_63671; // @[Modules.scala 150:103:@9955.4]
  wire [4:0] _T_63672; // @[Modules.scala 150:103:@9956.4]
  wire [4:0] _T_63683; // @[Modules.scala 151:80:@9965.4]
  wire [5:0] _T_63684; // @[Modules.scala 150:103:@9966.4]
  wire [4:0] _T_63685; // @[Modules.scala 150:103:@9967.4]
  wire [4:0] _T_63686; // @[Modules.scala 150:103:@9968.4]
  wire [4:0] _T_63688; // @[Modules.scala 150:74:@9970.4]
  wire [5:0] _T_63691; // @[Modules.scala 150:103:@9972.4]
  wire [4:0] _T_63692; // @[Modules.scala 150:103:@9973.4]
  wire [4:0] _T_63693; // @[Modules.scala 150:103:@9974.4]
  wire [5:0] _T_63698; // @[Modules.scala 150:103:@9978.4]
  wire [4:0] _T_63699; // @[Modules.scala 150:103:@9979.4]
  wire [4:0] _T_63700; // @[Modules.scala 150:103:@9980.4]
  wire [5:0] _T_63704; // @[Modules.scala 151:80:@9983.4]
  wire [5:0] _GEN_224; // @[Modules.scala 150:103:@9984.4]
  wire [6:0] _T_63705; // @[Modules.scala 150:103:@9984.4]
  wire [5:0] _T_63706; // @[Modules.scala 150:103:@9985.4]
  wire [5:0] _T_63707; // @[Modules.scala 150:103:@9986.4]
  wire [5:0] _T_63712; // @[Modules.scala 150:103:@9990.4]
  wire [4:0] _T_63713; // @[Modules.scala 150:103:@9991.4]
  wire [4:0] _T_63714; // @[Modules.scala 150:103:@9992.4]
  wire [5:0] _T_63719; // @[Modules.scala 150:103:@9996.4]
  wire [4:0] _T_63720; // @[Modules.scala 150:103:@9997.4]
  wire [4:0] _T_63721; // @[Modules.scala 150:103:@9998.4]
  wire [5:0] _T_63723; // @[Modules.scala 150:74:@10000.4]
  wire [6:0] _T_63726; // @[Modules.scala 150:103:@10002.4]
  wire [5:0] _T_63727; // @[Modules.scala 150:103:@10003.4]
  wire [5:0] _T_63728; // @[Modules.scala 150:103:@10004.4]
  wire [5:0] _T_63730; // @[Modules.scala 150:74:@10006.4]
  wire [6:0] _T_63733; // @[Modules.scala 150:103:@10008.4]
  wire [5:0] _T_63734; // @[Modules.scala 150:103:@10009.4]
  wire [5:0] _T_63735; // @[Modules.scala 150:103:@10010.4]
  wire [5:0] _T_63739; // @[Modules.scala 151:80:@10013.4]
  wire [6:0] _T_63740; // @[Modules.scala 150:103:@10014.4]
  wire [5:0] _T_63741; // @[Modules.scala 150:103:@10015.4]
  wire [5:0] _T_63742; // @[Modules.scala 150:103:@10016.4]
  wire [4:0] _T_63746; // @[Modules.scala 151:80:@10019.4]
  wire [5:0] _GEN_225; // @[Modules.scala 150:103:@10020.4]
  wire [6:0] _T_63747; // @[Modules.scala 150:103:@10020.4]
  wire [5:0] _T_63748; // @[Modules.scala 150:103:@10021.4]
  wire [5:0] _T_63749; // @[Modules.scala 150:103:@10022.4]
  wire [6:0] _T_63754; // @[Modules.scala 150:103:@10026.4]
  wire [5:0] _T_63755; // @[Modules.scala 150:103:@10027.4]
  wire [5:0] _T_63756; // @[Modules.scala 150:103:@10028.4]
  wire [4:0] _T_63760; // @[Modules.scala 151:80:@10031.4]
  wire [5:0] _T_63761; // @[Modules.scala 150:103:@10032.4]
  wire [4:0] _T_63762; // @[Modules.scala 150:103:@10033.4]
  wire [4:0] _T_63763; // @[Modules.scala 150:103:@10034.4]
  wire [5:0] _T_63768; // @[Modules.scala 150:103:@10038.4]
  wire [4:0] _T_63769; // @[Modules.scala 150:103:@10039.4]
  wire [4:0] _T_63770; // @[Modules.scala 150:103:@10040.4]
  wire [4:0] _T_63772; // @[Modules.scala 150:74:@10042.4]
  wire [4:0] _T_63774; // @[Modules.scala 151:80:@10043.4]
  wire [5:0] _T_63775; // @[Modules.scala 150:103:@10044.4]
  wire [4:0] _T_63776; // @[Modules.scala 150:103:@10045.4]
  wire [4:0] _T_63777; // @[Modules.scala 150:103:@10046.4]
  wire [5:0] _T_63782; // @[Modules.scala 150:103:@10050.4]
  wire [4:0] _T_63783; // @[Modules.scala 150:103:@10051.4]
  wire [4:0] _T_63784; // @[Modules.scala 150:103:@10052.4]
  wire [5:0] _GEN_227; // @[Modules.scala 150:103:@10056.4]
  wire [6:0] _T_63789; // @[Modules.scala 150:103:@10056.4]
  wire [5:0] _T_63790; // @[Modules.scala 150:103:@10057.4]
  wire [5:0] _T_63791; // @[Modules.scala 150:103:@10058.4]
  wire [5:0] _T_63796; // @[Modules.scala 150:103:@10062.4]
  wire [4:0] _T_63797; // @[Modules.scala 150:103:@10063.4]
  wire [4:0] _T_63798; // @[Modules.scala 150:103:@10064.4]
  wire [5:0] _T_63810; // @[Modules.scala 150:103:@10074.4]
  wire [4:0] _T_63811; // @[Modules.scala 150:103:@10075.4]
  wire [4:0] _T_63812; // @[Modules.scala 150:103:@10076.4]
  wire [5:0] _T_63814; // @[Modules.scala 150:74:@10078.4]
  wire [6:0] _T_63817; // @[Modules.scala 150:103:@10080.4]
  wire [5:0] _T_63818; // @[Modules.scala 150:103:@10081.4]
  wire [5:0] _T_63819; // @[Modules.scala 150:103:@10082.4]
  wire [5:0] _T_63821; // @[Modules.scala 150:74:@10084.4]
  wire [5:0] _T_63823; // @[Modules.scala 151:80:@10085.4]
  wire [6:0] _T_63824; // @[Modules.scala 150:103:@10086.4]
  wire [5:0] _T_63825; // @[Modules.scala 150:103:@10087.4]
  wire [5:0] _T_63826; // @[Modules.scala 150:103:@10088.4]
  wire [4:0] _T_63828; // @[Modules.scala 150:74:@10090.4]
  wire [5:0] _GEN_228; // @[Modules.scala 150:103:@10092.4]
  wire [6:0] _T_63831; // @[Modules.scala 150:103:@10092.4]
  wire [5:0] _T_63832; // @[Modules.scala 150:103:@10093.4]
  wire [5:0] _T_63833; // @[Modules.scala 150:103:@10094.4]
  wire [4:0] _T_63835; // @[Modules.scala 150:74:@10096.4]
  wire [5:0] _T_63838; // @[Modules.scala 150:103:@10098.4]
  wire [4:0] _T_63839; // @[Modules.scala 150:103:@10099.4]
  wire [4:0] _T_63840; // @[Modules.scala 150:103:@10100.4]
  wire [5:0] _T_63845; // @[Modules.scala 150:103:@10104.4]
  wire [4:0] _T_63846; // @[Modules.scala 150:103:@10105.4]
  wire [4:0] _T_63847; // @[Modules.scala 150:103:@10106.4]
  wire [5:0] _T_63852; // @[Modules.scala 150:103:@10110.4]
  wire [4:0] _T_63853; // @[Modules.scala 150:103:@10111.4]
  wire [4:0] _T_63854; // @[Modules.scala 150:103:@10112.4]
  wire [5:0] _T_63859; // @[Modules.scala 150:103:@10116.4]
  wire [4:0] _T_63860; // @[Modules.scala 150:103:@10117.4]
  wire [4:0] _T_63861; // @[Modules.scala 150:103:@10118.4]
  wire [5:0] _T_63866; // @[Modules.scala 150:103:@10122.4]
  wire [4:0] _T_63867; // @[Modules.scala 150:103:@10123.4]
  wire [4:0] _T_63868; // @[Modules.scala 150:103:@10124.4]
  wire [5:0] _GEN_229; // @[Modules.scala 150:103:@10128.4]
  wire [6:0] _T_63873; // @[Modules.scala 150:103:@10128.4]
  wire [5:0] _T_63874; // @[Modules.scala 150:103:@10129.4]
  wire [5:0] _T_63875; // @[Modules.scala 150:103:@10130.4]
  wire [6:0] _T_63880; // @[Modules.scala 150:103:@10134.4]
  wire [5:0] _T_63881; // @[Modules.scala 150:103:@10135.4]
  wire [5:0] _T_63882; // @[Modules.scala 150:103:@10136.4]
  wire [5:0] _T_63884; // @[Modules.scala 150:74:@10138.4]
  wire [5:0] _GEN_230; // @[Modules.scala 150:103:@10140.4]
  wire [6:0] _T_63887; // @[Modules.scala 150:103:@10140.4]
  wire [5:0] _T_63888; // @[Modules.scala 150:103:@10141.4]
  wire [5:0] _T_63889; // @[Modules.scala 150:103:@10142.4]
  wire [5:0] _T_63893; // @[Modules.scala 151:80:@10145.4]
  wire [5:0] _GEN_231; // @[Modules.scala 150:103:@10146.4]
  wire [6:0] _T_63894; // @[Modules.scala 150:103:@10146.4]
  wire [5:0] _T_63895; // @[Modules.scala 150:103:@10147.4]
  wire [5:0] _T_63896; // @[Modules.scala 150:103:@10148.4]
  wire [5:0] _T_63898; // @[Modules.scala 150:74:@10150.4]
  wire [5:0] _T_63900; // @[Modules.scala 151:80:@10151.4]
  wire [6:0] _T_63901; // @[Modules.scala 150:103:@10152.4]
  wire [5:0] _T_63902; // @[Modules.scala 150:103:@10153.4]
  wire [5:0] _T_63903; // @[Modules.scala 150:103:@10154.4]
  wire [5:0] _T_63905; // @[Modules.scala 150:74:@10156.4]
  wire [5:0] _T_63907; // @[Modules.scala 151:80:@10157.4]
  wire [6:0] _T_63908; // @[Modules.scala 150:103:@10158.4]
  wire [5:0] _T_63909; // @[Modules.scala 150:103:@10159.4]
  wire [5:0] _T_63910; // @[Modules.scala 150:103:@10160.4]
  wire [5:0] _T_63915; // @[Modules.scala 150:103:@10164.4]
  wire [4:0] _T_63916; // @[Modules.scala 150:103:@10165.4]
  wire [4:0] _T_63917; // @[Modules.scala 150:103:@10166.4]
  wire [5:0] _T_63943; // @[Modules.scala 150:103:@10188.4]
  wire [4:0] _T_63944; // @[Modules.scala 150:103:@10189.4]
  wire [4:0] _T_63945; // @[Modules.scala 150:103:@10190.4]
  wire [5:0] _T_63950; // @[Modules.scala 150:103:@10194.4]
  wire [4:0] _T_63951; // @[Modules.scala 150:103:@10195.4]
  wire [4:0] _T_63952; // @[Modules.scala 150:103:@10196.4]
  wire [5:0] _T_63968; // @[Modules.scala 150:74:@10210.4]
  wire [5:0] _T_63970; // @[Modules.scala 151:80:@10211.4]
  wire [6:0] _T_63971; // @[Modules.scala 150:103:@10212.4]
  wire [5:0] _T_63972; // @[Modules.scala 150:103:@10213.4]
  wire [5:0] _T_63973; // @[Modules.scala 150:103:@10214.4]
  wire [5:0] _T_63975; // @[Modules.scala 150:74:@10216.4]
  wire [5:0] _T_63977; // @[Modules.scala 151:80:@10217.4]
  wire [6:0] _T_63978; // @[Modules.scala 150:103:@10218.4]
  wire [5:0] _T_63979; // @[Modules.scala 150:103:@10219.4]
  wire [5:0] _T_63980; // @[Modules.scala 150:103:@10220.4]
  wire [5:0] _T_63982; // @[Modules.scala 150:74:@10222.4]
  wire [5:0] _T_63984; // @[Modules.scala 151:80:@10223.4]
  wire [6:0] _T_63985; // @[Modules.scala 150:103:@10224.4]
  wire [5:0] _T_63986; // @[Modules.scala 150:103:@10225.4]
  wire [5:0] _T_63987; // @[Modules.scala 150:103:@10226.4]
  wire [5:0] _T_63989; // @[Modules.scala 150:74:@10228.4]
  wire [6:0] _T_63992; // @[Modules.scala 150:103:@10230.4]
  wire [5:0] _T_63993; // @[Modules.scala 150:103:@10231.4]
  wire [5:0] _T_63994; // @[Modules.scala 150:103:@10232.4]
  wire [4:0] _T_63996; // @[Modules.scala 150:74:@10234.4]
  wire [5:0] _T_63999; // @[Modules.scala 150:103:@10236.4]
  wire [4:0] _T_64000; // @[Modules.scala 150:103:@10237.4]
  wire [4:0] _T_64001; // @[Modules.scala 150:103:@10238.4]
  wire [5:0] _T_64006; // @[Modules.scala 150:103:@10242.4]
  wire [4:0] _T_64007; // @[Modules.scala 150:103:@10243.4]
  wire [4:0] _T_64008; // @[Modules.scala 150:103:@10244.4]
  wire [5:0] _T_64013; // @[Modules.scala 150:103:@10248.4]
  wire [4:0] _T_64014; // @[Modules.scala 150:103:@10249.4]
  wire [4:0] _T_64015; // @[Modules.scala 150:103:@10250.4]
  wire [5:0] _T_64019; // @[Modules.scala 151:80:@10253.4]
  wire [6:0] _T_64020; // @[Modules.scala 150:103:@10254.4]
  wire [5:0] _T_64021; // @[Modules.scala 150:103:@10255.4]
  wire [5:0] _T_64022; // @[Modules.scala 150:103:@10256.4]
  wire [5:0] _T_64026; // @[Modules.scala 151:80:@10259.4]
  wire [6:0] _T_64027; // @[Modules.scala 150:103:@10260.4]
  wire [5:0] _T_64028; // @[Modules.scala 150:103:@10261.4]
  wire [5:0] _T_64029; // @[Modules.scala 150:103:@10262.4]
  wire [5:0] _T_64034; // @[Modules.scala 150:103:@10266.4]
  wire [4:0] _T_64035; // @[Modules.scala 150:103:@10267.4]
  wire [4:0] _T_64036; // @[Modules.scala 150:103:@10268.4]
  wire [5:0] _T_64041; // @[Modules.scala 150:103:@10272.4]
  wire [4:0] _T_64042; // @[Modules.scala 150:103:@10273.4]
  wire [4:0] _T_64043; // @[Modules.scala 150:103:@10274.4]
  wire [5:0] _T_64061; // @[Modules.scala 151:80:@10289.4]
  wire [5:0] _GEN_233; // @[Modules.scala 150:103:@10290.4]
  wire [6:0] _T_64062; // @[Modules.scala 150:103:@10290.4]
  wire [5:0] _T_64063; // @[Modules.scala 150:103:@10291.4]
  wire [5:0] _T_64064; // @[Modules.scala 150:103:@10292.4]
  wire [5:0] _T_64066; // @[Modules.scala 150:74:@10294.4]
  wire [5:0] _T_64068; // @[Modules.scala 151:80:@10295.4]
  wire [6:0] _T_64069; // @[Modules.scala 150:103:@10296.4]
  wire [5:0] _T_64070; // @[Modules.scala 150:103:@10297.4]
  wire [5:0] _T_64071; // @[Modules.scala 150:103:@10298.4]
  wire [5:0] _T_64073; // @[Modules.scala 150:74:@10300.4]
  wire [5:0] _T_64075; // @[Modules.scala 151:80:@10301.4]
  wire [6:0] _T_64076; // @[Modules.scala 150:103:@10302.4]
  wire [5:0] _T_64077; // @[Modules.scala 150:103:@10303.4]
  wire [5:0] _T_64078; // @[Modules.scala 150:103:@10304.4]
  wire [5:0] _GEN_234; // @[Modules.scala 150:103:@10314.4]
  wire [6:0] _T_64090; // @[Modules.scala 150:103:@10314.4]
  wire [5:0] _T_64091; // @[Modules.scala 150:103:@10315.4]
  wire [5:0] _T_64092; // @[Modules.scala 150:103:@10316.4]
  wire [5:0] _T_64097; // @[Modules.scala 150:103:@10320.4]
  wire [4:0] _T_64098; // @[Modules.scala 150:103:@10321.4]
  wire [4:0] _T_64099; // @[Modules.scala 150:103:@10322.4]
  wire [5:0] _T_64103; // @[Modules.scala 151:80:@10325.4]
  wire [5:0] _GEN_235; // @[Modules.scala 150:103:@10326.4]
  wire [6:0] _T_64104; // @[Modules.scala 150:103:@10326.4]
  wire [5:0] _T_64105; // @[Modules.scala 150:103:@10327.4]
  wire [5:0] _T_64106; // @[Modules.scala 150:103:@10328.4]
  wire [5:0] _T_64108; // @[Modules.scala 150:74:@10330.4]
  wire [6:0] _T_64111; // @[Modules.scala 150:103:@10332.4]
  wire [5:0] _T_64112; // @[Modules.scala 150:103:@10333.4]
  wire [5:0] _T_64113; // @[Modules.scala 150:103:@10334.4]
  wire [5:0] _T_64115; // @[Modules.scala 150:74:@10336.4]
  wire [6:0] _T_64118; // @[Modules.scala 150:103:@10338.4]
  wire [5:0] _T_64119; // @[Modules.scala 150:103:@10339.4]
  wire [5:0] _T_64120; // @[Modules.scala 150:103:@10340.4]
  wire [5:0] _T_64122; // @[Modules.scala 150:74:@10342.4]
  wire [5:0] _T_64124; // @[Modules.scala 151:80:@10343.4]
  wire [6:0] _T_64125; // @[Modules.scala 150:103:@10344.4]
  wire [5:0] _T_64126; // @[Modules.scala 150:103:@10345.4]
  wire [5:0] _T_64127; // @[Modules.scala 150:103:@10346.4]
  wire [5:0] _T_64132; // @[Modules.scala 150:103:@10350.4]
  wire [4:0] _T_64133; // @[Modules.scala 150:103:@10351.4]
  wire [4:0] _T_64134; // @[Modules.scala 150:103:@10352.4]
  wire [5:0] _T_64139; // @[Modules.scala 150:103:@10356.4]
  wire [4:0] _T_64140; // @[Modules.scala 150:103:@10357.4]
  wire [4:0] _T_64141; // @[Modules.scala 150:103:@10358.4]
  wire [5:0] _T_64164; // @[Modules.scala 150:74:@10378.4]
  wire [5:0] _T_64166; // @[Modules.scala 151:80:@10379.4]
  wire [6:0] _T_64167; // @[Modules.scala 150:103:@10380.4]
  wire [5:0] _T_64168; // @[Modules.scala 150:103:@10381.4]
  wire [5:0] _T_64169; // @[Modules.scala 150:103:@10382.4]
  wire [5:0] _T_64171; // @[Modules.scala 150:74:@10384.4]
  wire [4:0] _T_64173; // @[Modules.scala 151:80:@10385.4]
  wire [5:0] _GEN_236; // @[Modules.scala 150:103:@10386.4]
  wire [6:0] _T_64174; // @[Modules.scala 150:103:@10386.4]
  wire [5:0] _T_64175; // @[Modules.scala 150:103:@10387.4]
  wire [5:0] _T_64176; // @[Modules.scala 150:103:@10388.4]
  wire [5:0] _T_64181; // @[Modules.scala 150:103:@10392.4]
  wire [4:0] _T_64182; // @[Modules.scala 150:103:@10393.4]
  wire [4:0] _T_64183; // @[Modules.scala 150:103:@10394.4]
  wire [5:0] _T_64194; // @[Modules.scala 151:80:@10403.4]
  wire [6:0] _T_64195; // @[Modules.scala 150:103:@10404.4]
  wire [5:0] _T_64196; // @[Modules.scala 150:103:@10405.4]
  wire [5:0] _T_64197; // @[Modules.scala 150:103:@10406.4]
  wire [6:0] _T_64202; // @[Modules.scala 150:103:@10410.4]
  wire [5:0] _T_64203; // @[Modules.scala 150:103:@10411.4]
  wire [5:0] _T_64204; // @[Modules.scala 150:103:@10412.4]
  wire [6:0] _T_64209; // @[Modules.scala 150:103:@10416.4]
  wire [5:0] _T_64210; // @[Modules.scala 150:103:@10417.4]
  wire [5:0] _T_64211; // @[Modules.scala 150:103:@10418.4]
  wire [6:0] _T_64216; // @[Modules.scala 150:103:@10422.4]
  wire [5:0] _T_64217; // @[Modules.scala 150:103:@10423.4]
  wire [5:0] _T_64218; // @[Modules.scala 150:103:@10424.4]
  wire [6:0] _T_64223; // @[Modules.scala 150:103:@10428.4]
  wire [5:0] _T_64224; // @[Modules.scala 150:103:@10429.4]
  wire [5:0] _T_64225; // @[Modules.scala 150:103:@10430.4]
  wire [6:0] _T_64230; // @[Modules.scala 150:103:@10434.4]
  wire [5:0] _T_64231; // @[Modules.scala 150:103:@10435.4]
  wire [5:0] _T_64232; // @[Modules.scala 150:103:@10436.4]
  wire [5:0] _T_64262; // @[Modules.scala 150:74:@10462.4]
  wire [5:0] _T_64264; // @[Modules.scala 151:80:@10463.4]
  wire [6:0] _T_64265; // @[Modules.scala 150:103:@10464.4]
  wire [5:0] _T_64266; // @[Modules.scala 150:103:@10465.4]
  wire [5:0] _T_64267; // @[Modules.scala 150:103:@10466.4]
  wire [6:0] _T_64272; // @[Modules.scala 150:103:@10470.4]
  wire [5:0] _T_64273; // @[Modules.scala 150:103:@10471.4]
  wire [5:0] _T_64274; // @[Modules.scala 150:103:@10472.4]
  wire [5:0] _GEN_239; // @[Modules.scala 150:103:@10482.4]
  wire [6:0] _T_64286; // @[Modules.scala 150:103:@10482.4]
  wire [5:0] _T_64287; // @[Modules.scala 150:103:@10483.4]
  wire [5:0] _T_64288; // @[Modules.scala 150:103:@10484.4]
  wire [6:0] _T_64293; // @[Modules.scala 150:103:@10488.4]
  wire [5:0] _T_64294; // @[Modules.scala 150:103:@10489.4]
  wire [5:0] _T_64295; // @[Modules.scala 150:103:@10490.4]
  wire [4:0] _T_64334; // @[Modules.scala 151:80:@10523.4]
  wire [5:0] _T_64335; // @[Modules.scala 150:103:@10524.4]
  wire [4:0] _T_64336; // @[Modules.scala 150:103:@10525.4]
  wire [4:0] _T_64337; // @[Modules.scala 150:103:@10526.4]
  wire [5:0] _T_64342; // @[Modules.scala 150:103:@10530.4]
  wire [4:0] _T_64343; // @[Modules.scala 150:103:@10531.4]
  wire [4:0] _T_64344; // @[Modules.scala 150:103:@10532.4]
  wire [5:0] _T_64349; // @[Modules.scala 150:103:@10536.4]
  wire [4:0] _T_64350; // @[Modules.scala 150:103:@10537.4]
  wire [4:0] _T_64351; // @[Modules.scala 150:103:@10538.4]
  wire [5:0] _T_64355; // @[Modules.scala 151:80:@10541.4]
  wire [6:0] _T_64356; // @[Modules.scala 150:103:@10542.4]
  wire [5:0] _T_64357; // @[Modules.scala 150:103:@10543.4]
  wire [5:0] _T_64358; // @[Modules.scala 150:103:@10544.4]
  wire [5:0] _GEN_240; // @[Modules.scala 150:103:@10548.4]
  wire [6:0] _T_64363; // @[Modules.scala 150:103:@10548.4]
  wire [5:0] _T_64364; // @[Modules.scala 150:103:@10549.4]
  wire [5:0] _T_64365; // @[Modules.scala 150:103:@10550.4]
  wire [6:0] _T_64377; // @[Modules.scala 150:103:@10560.4]
  wire [5:0] _T_64378; // @[Modules.scala 150:103:@10561.4]
  wire [5:0] _T_64379; // @[Modules.scala 150:103:@10562.4]
  wire [6:0] _T_64412; // @[Modules.scala 150:103:@10590.4]
  wire [5:0] _T_64413; // @[Modules.scala 150:103:@10591.4]
  wire [5:0] _T_64414; // @[Modules.scala 150:103:@10592.4]
  wire [6:0] _T_64433; // @[Modules.scala 150:103:@10608.4]
  wire [5:0] _T_64434; // @[Modules.scala 150:103:@10609.4]
  wire [5:0] _T_64435; // @[Modules.scala 150:103:@10610.4]
  wire [5:0] _T_64440; // @[Modules.scala 150:103:@10614.4]
  wire [4:0] _T_64441; // @[Modules.scala 150:103:@10615.4]
  wire [4:0] _T_64442; // @[Modules.scala 150:103:@10616.4]
  wire [5:0] _T_64447; // @[Modules.scala 150:103:@10620.4]
  wire [4:0] _T_64448; // @[Modules.scala 150:103:@10621.4]
  wire [4:0] _T_64449; // @[Modules.scala 150:103:@10622.4]
  wire [6:0] _T_64454; // @[Modules.scala 150:103:@10626.4]
  wire [5:0] _T_64455; // @[Modules.scala 150:103:@10627.4]
  wire [5:0] _T_64456; // @[Modules.scala 150:103:@10628.4]
  wire [4:0] _T_64458; // @[Modules.scala 150:74:@10630.4]
  wire [5:0] _GEN_242; // @[Modules.scala 150:103:@10632.4]
  wire [6:0] _T_64461; // @[Modules.scala 150:103:@10632.4]
  wire [5:0] _T_64462; // @[Modules.scala 150:103:@10633.4]
  wire [5:0] _T_64463; // @[Modules.scala 150:103:@10634.4]
  wire [6:0] _T_64489; // @[Modules.scala 150:103:@10656.4]
  wire [5:0] _T_64490; // @[Modules.scala 150:103:@10657.4]
  wire [5:0] _T_64491; // @[Modules.scala 150:103:@10658.4]
  wire [6:0] _T_64496; // @[Modules.scala 150:103:@10662.4]
  wire [5:0] _T_64497; // @[Modules.scala 150:103:@10663.4]
  wire [5:0] _T_64498; // @[Modules.scala 150:103:@10664.4]
  wire [5:0] _GEN_243; // @[Modules.scala 150:103:@10674.4]
  wire [6:0] _T_64510; // @[Modules.scala 150:103:@10674.4]
  wire [5:0] _T_64511; // @[Modules.scala 150:103:@10675.4]
  wire [5:0] _T_64512; // @[Modules.scala 150:103:@10676.4]
  wire [6:0] _T_64531; // @[Modules.scala 150:103:@10692.4]
  wire [5:0] _T_64532; // @[Modules.scala 150:103:@10693.4]
  wire [5:0] _T_64533; // @[Modules.scala 150:103:@10694.4]
  wire [5:0] _GEN_245; // @[Modules.scala 150:103:@10704.4]
  wire [6:0] _T_64545; // @[Modules.scala 150:103:@10704.4]
  wire [5:0] _T_64546; // @[Modules.scala 150:103:@10705.4]
  wire [5:0] _T_64547; // @[Modules.scala 150:103:@10706.4]
  wire [5:0] _T_64549; // @[Modules.scala 150:74:@10708.4]
  wire [6:0] _T_64552; // @[Modules.scala 150:103:@10710.4]
  wire [5:0] _T_64553; // @[Modules.scala 150:103:@10711.4]
  wire [5:0] _T_64554; // @[Modules.scala 150:103:@10712.4]
  wire [5:0] _T_64573; // @[Modules.scala 150:103:@10728.4]
  wire [4:0] _T_64574; // @[Modules.scala 150:103:@10729.4]
  wire [4:0] _T_64575; // @[Modules.scala 150:103:@10730.4]
  wire [4:0] _T_64579; // @[Modules.scala 151:80:@10733.4]
  wire [5:0] _T_64580; // @[Modules.scala 150:103:@10734.4]
  wire [4:0] _T_64581; // @[Modules.scala 150:103:@10735.4]
  wire [4:0] _T_64582; // @[Modules.scala 150:103:@10736.4]
  wire [5:0] _T_64587; // @[Modules.scala 150:103:@10740.4]
  wire [4:0] _T_64588; // @[Modules.scala 150:103:@10741.4]
  wire [4:0] _T_64589; // @[Modules.scala 150:103:@10742.4]
  wire [5:0] _T_64608; // @[Modules.scala 150:103:@10758.4]
  wire [4:0] _T_64609; // @[Modules.scala 150:103:@10759.4]
  wire [4:0] _T_64610; // @[Modules.scala 150:103:@10760.4]
  wire [4:0] _T_64614; // @[Modules.scala 151:80:@10763.4]
  wire [5:0] _T_64615; // @[Modules.scala 150:103:@10764.4]
  wire [4:0] _T_64616; // @[Modules.scala 150:103:@10765.4]
  wire [4:0] _T_64617; // @[Modules.scala 150:103:@10766.4]
  wire [5:0] _T_64622; // @[Modules.scala 150:103:@10770.4]
  wire [4:0] _T_64623; // @[Modules.scala 150:103:@10771.4]
  wire [4:0] _T_64624; // @[Modules.scala 150:103:@10772.4]
  wire [5:0] _T_64635; // @[Modules.scala 151:80:@10781.4]
  wire [5:0] _GEN_247; // @[Modules.scala 150:103:@10782.4]
  wire [6:0] _T_64636; // @[Modules.scala 150:103:@10782.4]
  wire [5:0] _T_64637; // @[Modules.scala 150:103:@10783.4]
  wire [5:0] _T_64638; // @[Modules.scala 150:103:@10784.4]
  wire [6:0] _T_64643; // @[Modules.scala 150:103:@10788.4]
  wire [5:0] _T_64644; // @[Modules.scala 150:103:@10789.4]
  wire [5:0] _T_64645; // @[Modules.scala 150:103:@10790.4]
  wire [5:0] _T_64649; // @[Modules.scala 151:80:@10793.4]
  wire [6:0] _T_64650; // @[Modules.scala 150:103:@10794.4]
  wire [5:0] _T_64651; // @[Modules.scala 150:103:@10795.4]
  wire [5:0] _T_64652; // @[Modules.scala 150:103:@10796.4]
  wire [5:0] _T_64671; // @[Modules.scala 150:103:@10812.4]
  wire [4:0] _T_64672; // @[Modules.scala 150:103:@10813.4]
  wire [4:0] _T_64673; // @[Modules.scala 150:103:@10814.4]
  wire [4:0] _T_64675; // @[Modules.scala 150:74:@10816.4]
  wire [4:0] _T_64677; // @[Modules.scala 151:80:@10817.4]
  wire [5:0] _T_64678; // @[Modules.scala 150:103:@10818.4]
  wire [4:0] _T_64679; // @[Modules.scala 150:103:@10819.4]
  wire [4:0] _T_64680; // @[Modules.scala 150:103:@10820.4]
  wire [5:0] _T_64699; // @[Modules.scala 150:103:@10836.4]
  wire [4:0] _T_64700; // @[Modules.scala 150:103:@10837.4]
  wire [4:0] _T_64701; // @[Modules.scala 150:103:@10838.4]
  wire [5:0] _GEN_249; // @[Modules.scala 150:103:@10842.4]
  wire [6:0] _T_64706; // @[Modules.scala 150:103:@10842.4]
  wire [5:0] _T_64707; // @[Modules.scala 150:103:@10843.4]
  wire [5:0] _T_64708; // @[Modules.scala 150:103:@10844.4]
  wire [5:0] _T_64713; // @[Modules.scala 150:103:@10848.4]
  wire [4:0] _T_64714; // @[Modules.scala 150:103:@10849.4]
  wire [4:0] _T_64715; // @[Modules.scala 150:103:@10850.4]
  wire [5:0] _T_64720; // @[Modules.scala 150:103:@10854.4]
  wire [4:0] _T_64721; // @[Modules.scala 150:103:@10855.4]
  wire [4:0] _T_64722; // @[Modules.scala 150:103:@10856.4]
  wire [5:0] _T_64726; // @[Modules.scala 151:80:@10859.4]
  wire [6:0] _T_64727; // @[Modules.scala 150:103:@10860.4]
  wire [5:0] _T_64728; // @[Modules.scala 150:103:@10861.4]
  wire [5:0] _T_64729; // @[Modules.scala 150:103:@10862.4]
  wire [6:0] _T_64748; // @[Modules.scala 150:103:@10878.4]
  wire [5:0] _T_64749; // @[Modules.scala 150:103:@10879.4]
  wire [5:0] _T_64750; // @[Modules.scala 150:103:@10880.4]
  wire [4:0] _T_64754; // @[Modules.scala 151:80:@10883.4]
  wire [5:0] _T_64755; // @[Modules.scala 150:103:@10884.4]
  wire [4:0] _T_64756; // @[Modules.scala 150:103:@10885.4]
  wire [4:0] _T_64757; // @[Modules.scala 150:103:@10886.4]
  wire [4:0] _T_64768; // @[Modules.scala 151:80:@10895.4]
  wire [5:0] _T_64769; // @[Modules.scala 150:103:@10896.4]
  wire [4:0] _T_64770; // @[Modules.scala 150:103:@10897.4]
  wire [4:0] _T_64771; // @[Modules.scala 150:103:@10898.4]
  wire [5:0] _GEN_251; // @[Modules.scala 150:103:@10902.4]
  wire [6:0] _T_64776; // @[Modules.scala 150:103:@10902.4]
  wire [5:0] _T_64777; // @[Modules.scala 150:103:@10903.4]
  wire [5:0] _T_64778; // @[Modules.scala 150:103:@10904.4]
  wire [4:0] _T_64782; // @[Modules.scala 151:80:@10907.4]
  wire [5:0] _GEN_252; // @[Modules.scala 150:103:@10908.4]
  wire [6:0] _T_64783; // @[Modules.scala 150:103:@10908.4]
  wire [5:0] _T_64784; // @[Modules.scala 150:103:@10909.4]
  wire [5:0] _T_64785; // @[Modules.scala 150:103:@10910.4]
  wire [5:0] _T_64790; // @[Modules.scala 150:103:@10914.4]
  wire [4:0] _T_64791; // @[Modules.scala 150:103:@10915.4]
  wire [4:0] _T_64792; // @[Modules.scala 150:103:@10916.4]
  wire [5:0] _T_64796; // @[Modules.scala 151:80:@10919.4]
  wire [6:0] _T_64797; // @[Modules.scala 150:103:@10920.4]
  wire [5:0] _T_64798; // @[Modules.scala 150:103:@10921.4]
  wire [5:0] _T_64799; // @[Modules.scala 150:103:@10922.4]
  wire [5:0] _GEN_254; // @[Modules.scala 150:103:@10926.4]
  wire [6:0] _T_64804; // @[Modules.scala 150:103:@10926.4]
  wire [5:0] _T_64805; // @[Modules.scala 150:103:@10927.4]
  wire [5:0] _T_64806; // @[Modules.scala 150:103:@10928.4]
  wire [6:0] _T_64825; // @[Modules.scala 150:103:@10944.4]
  wire [5:0] _T_64826; // @[Modules.scala 150:103:@10945.4]
  wire [5:0] _T_64827; // @[Modules.scala 150:103:@10946.4]
  wire [4:0] _T_64829; // @[Modules.scala 150:74:@10948.4]
  wire [4:0] _T_64831; // @[Modules.scala 151:80:@10949.4]
  wire [5:0] _T_64832; // @[Modules.scala 150:103:@10950.4]
  wire [4:0] _T_64833; // @[Modules.scala 150:103:@10951.4]
  wire [4:0] _T_64834; // @[Modules.scala 150:103:@10952.4]
  wire [4:0] _T_64838; // @[Modules.scala 151:80:@10955.4]
  wire [5:0] _GEN_256; // @[Modules.scala 150:103:@10956.4]
  wire [6:0] _T_64839; // @[Modules.scala 150:103:@10956.4]
  wire [5:0] _T_64840; // @[Modules.scala 150:103:@10957.4]
  wire [5:0] _T_64841; // @[Modules.scala 150:103:@10958.4]
  wire [5:0] _T_64846; // @[Modules.scala 150:103:@10962.4]
  wire [4:0] _T_64847; // @[Modules.scala 150:103:@10963.4]
  wire [4:0] _T_64848; // @[Modules.scala 150:103:@10964.4]
  wire [5:0] _T_64853; // @[Modules.scala 150:103:@10968.4]
  wire [4:0] _T_64854; // @[Modules.scala 150:103:@10969.4]
  wire [4:0] _T_64855; // @[Modules.scala 150:103:@10970.4]
  wire [5:0] _GEN_257; // @[Modules.scala 150:103:@10974.4]
  wire [6:0] _T_64860; // @[Modules.scala 150:103:@10974.4]
  wire [5:0] _T_64861; // @[Modules.scala 150:103:@10975.4]
  wire [5:0] _T_64862; // @[Modules.scala 150:103:@10976.4]
  wire [6:0] _T_64867; // @[Modules.scala 150:103:@10980.4]
  wire [5:0] _T_64868; // @[Modules.scala 150:103:@10981.4]
  wire [5:0] _T_64869; // @[Modules.scala 150:103:@10982.4]
  wire [4:0] _T_64871; // @[Modules.scala 150:74:@10984.4]
  wire [5:0] _T_64874; // @[Modules.scala 150:103:@10986.4]
  wire [4:0] _T_64875; // @[Modules.scala 150:103:@10987.4]
  wire [4:0] _T_64876; // @[Modules.scala 150:103:@10988.4]
  wire [5:0] _T_64881; // @[Modules.scala 150:103:@10992.4]
  wire [4:0] _T_64882; // @[Modules.scala 150:103:@10993.4]
  wire [4:0] _T_64883; // @[Modules.scala 150:103:@10994.4]
  wire [5:0] _T_64888; // @[Modules.scala 150:103:@10998.4]
  wire [4:0] _T_64889; // @[Modules.scala 150:103:@10999.4]
  wire [4:0] _T_64890; // @[Modules.scala 150:103:@11000.4]
  wire [4:0] _T_64906; // @[Modules.scala 150:74:@11014.4]
  wire [5:0] _T_64909; // @[Modules.scala 150:103:@11016.4]
  wire [4:0] _T_64910; // @[Modules.scala 150:103:@11017.4]
  wire [4:0] _T_64911; // @[Modules.scala 150:103:@11018.4]
  wire [4:0] _T_64920; // @[Modules.scala 150:74:@11026.4]
  wire [5:0] _GEN_259; // @[Modules.scala 150:103:@11028.4]
  wire [6:0] _T_64923; // @[Modules.scala 150:103:@11028.4]
  wire [5:0] _T_64924; // @[Modules.scala 150:103:@11029.4]
  wire [5:0] _T_64925; // @[Modules.scala 150:103:@11030.4]
  wire [5:0] _T_64930; // @[Modules.scala 150:103:@11034.4]
  wire [4:0] _T_64931; // @[Modules.scala 150:103:@11035.4]
  wire [4:0] _T_64932; // @[Modules.scala 150:103:@11036.4]
  wire [5:0] _GEN_260; // @[Modules.scala 150:103:@11040.4]
  wire [6:0] _T_64937; // @[Modules.scala 150:103:@11040.4]
  wire [5:0] _T_64938; // @[Modules.scala 150:103:@11041.4]
  wire [5:0] _T_64939; // @[Modules.scala 150:103:@11042.4]
  wire [5:0] _T_64943; // @[Modules.scala 151:80:@11045.4]
  wire [5:0] _GEN_261; // @[Modules.scala 150:103:@11046.4]
  wire [6:0] _T_64944; // @[Modules.scala 150:103:@11046.4]
  wire [5:0] _T_64945; // @[Modules.scala 150:103:@11047.4]
  wire [5:0] _T_64946; // @[Modules.scala 150:103:@11048.4]
  wire [4:0] _T_64948; // @[Modules.scala 150:74:@11050.4]
  wire [4:0] _T_64950; // @[Modules.scala 151:80:@11051.4]
  wire [5:0] _T_64951; // @[Modules.scala 150:103:@11052.4]
  wire [4:0] _T_64952; // @[Modules.scala 150:103:@11053.4]
  wire [4:0] _T_64953; // @[Modules.scala 150:103:@11054.4]
  wire [5:0] _T_64969; // @[Modules.scala 150:74:@11068.4]
  wire [5:0] _GEN_262; // @[Modules.scala 150:103:@11070.4]
  wire [6:0] _T_64972; // @[Modules.scala 150:103:@11070.4]
  wire [5:0] _T_64973; // @[Modules.scala 150:103:@11071.4]
  wire [5:0] _T_64974; // @[Modules.scala 150:103:@11072.4]
  wire [5:0] _T_64979; // @[Modules.scala 150:103:@11076.4]
  wire [4:0] _T_64980; // @[Modules.scala 150:103:@11077.4]
  wire [4:0] _T_64981; // @[Modules.scala 150:103:@11078.4]
  wire [4:0] _T_64985; // @[Modules.scala 151:80:@11081.4]
  wire [5:0] _T_64986; // @[Modules.scala 150:103:@11082.4]
  wire [4:0] _T_64987; // @[Modules.scala 150:103:@11083.4]
  wire [4:0] _T_64988; // @[Modules.scala 150:103:@11084.4]
  wire [5:0] _T_65004; // @[Modules.scala 150:74:@11098.4]
  wire [6:0] _T_65007; // @[Modules.scala 150:103:@11100.4]
  wire [5:0] _T_65008; // @[Modules.scala 150:103:@11101.4]
  wire [5:0] _T_65009; // @[Modules.scala 150:103:@11102.4]
  wire [5:0] _T_65028; // @[Modules.scala 150:103:@11118.4]
  wire [4:0] _T_65029; // @[Modules.scala 150:103:@11119.4]
  wire [4:0] _T_65030; // @[Modules.scala 150:103:@11120.4]
  wire [5:0] _T_65035; // @[Modules.scala 150:103:@11124.4]
  wire [4:0] _T_65036; // @[Modules.scala 150:103:@11125.4]
  wire [4:0] _T_65037; // @[Modules.scala 150:103:@11126.4]
  wire [4:0] _T_65048; // @[Modules.scala 151:80:@11135.4]
  wire [5:0] _GEN_265; // @[Modules.scala 150:103:@11136.4]
  wire [6:0] _T_65049; // @[Modules.scala 150:103:@11136.4]
  wire [5:0] _T_65050; // @[Modules.scala 150:103:@11137.4]
  wire [5:0] _T_65051; // @[Modules.scala 150:103:@11138.4]
  wire [5:0] _T_65056; // @[Modules.scala 150:103:@11142.4]
  wire [4:0] _T_65057; // @[Modules.scala 150:103:@11143.4]
  wire [4:0] _T_65058; // @[Modules.scala 150:103:@11144.4]
  wire [6:0] _T_65063; // @[Modules.scala 150:103:@11148.4]
  wire [5:0] _T_65064; // @[Modules.scala 150:103:@11149.4]
  wire [5:0] _T_65065; // @[Modules.scala 150:103:@11150.4]
  wire [4:0] _T_65074; // @[Modules.scala 150:74:@11158.4]
  wire [5:0] _GEN_267; // @[Modules.scala 150:103:@11160.4]
  wire [6:0] _T_65077; // @[Modules.scala 150:103:@11160.4]
  wire [5:0] _T_65078; // @[Modules.scala 150:103:@11161.4]
  wire [5:0] _T_65079; // @[Modules.scala 150:103:@11162.4]
  wire [4:0] _T_65083; // @[Modules.scala 151:80:@11165.4]
  wire [5:0] _GEN_268; // @[Modules.scala 150:103:@11166.4]
  wire [6:0] _T_65084; // @[Modules.scala 150:103:@11166.4]
  wire [5:0] _T_65085; // @[Modules.scala 150:103:@11167.4]
  wire [5:0] _T_65086; // @[Modules.scala 150:103:@11168.4]
  wire [5:0] _T_65091; // @[Modules.scala 150:103:@11172.4]
  wire [4:0] _T_65092; // @[Modules.scala 150:103:@11173.4]
  wire [4:0] _T_65093; // @[Modules.scala 150:103:@11174.4]
  wire [5:0] _T_65098; // @[Modules.scala 150:103:@11178.4]
  wire [4:0] _T_65099; // @[Modules.scala 150:103:@11179.4]
  wire [4:0] _T_65100; // @[Modules.scala 150:103:@11180.4]
  wire [5:0] _T_65105; // @[Modules.scala 150:103:@11184.4]
  wire [4:0] _T_65106; // @[Modules.scala 150:103:@11185.4]
  wire [4:0] _T_65107; // @[Modules.scala 150:103:@11186.4]
  wire [5:0] _T_65112; // @[Modules.scala 150:103:@11190.4]
  wire [4:0] _T_65113; // @[Modules.scala 150:103:@11191.4]
  wire [4:0] _T_65114; // @[Modules.scala 150:103:@11192.4]
  wire [5:0] _T_65125; // @[Modules.scala 151:80:@11201.4]
  wire [5:0] _GEN_269; // @[Modules.scala 150:103:@11202.4]
  wire [6:0] _T_65126; // @[Modules.scala 150:103:@11202.4]
  wire [5:0] _T_65127; // @[Modules.scala 150:103:@11203.4]
  wire [5:0] _T_65128; // @[Modules.scala 150:103:@11204.4]
  wire [5:0] _T_65130; // @[Modules.scala 150:74:@11206.4]
  wire [6:0] _T_65133; // @[Modules.scala 150:103:@11208.4]
  wire [5:0] _T_65134; // @[Modules.scala 150:103:@11209.4]
  wire [5:0] _T_65135; // @[Modules.scala 150:103:@11210.4]
  wire [6:0] _T_65140; // @[Modules.scala 150:103:@11214.4]
  wire [5:0] _T_65141; // @[Modules.scala 150:103:@11215.4]
  wire [5:0] _T_65142; // @[Modules.scala 150:103:@11216.4]
  wire [5:0] _GEN_270; // @[Modules.scala 150:103:@11220.4]
  wire [6:0] _T_65147; // @[Modules.scala 150:103:@11220.4]
  wire [5:0] _T_65148; // @[Modules.scala 150:103:@11221.4]
  wire [5:0] _T_65149; // @[Modules.scala 150:103:@11222.4]
  wire [5:0] _GEN_271; // @[Modules.scala 150:103:@11226.4]
  wire [6:0] _T_65154; // @[Modules.scala 150:103:@11226.4]
  wire [5:0] _T_65155; // @[Modules.scala 150:103:@11227.4]
  wire [5:0] _T_65156; // @[Modules.scala 150:103:@11228.4]
  wire [4:0] _T_65160; // @[Modules.scala 151:80:@11231.4]
  wire [5:0] _T_65161; // @[Modules.scala 150:103:@11232.4]
  wire [4:0] _T_65162; // @[Modules.scala 150:103:@11233.4]
  wire [4:0] _T_65163; // @[Modules.scala 150:103:@11234.4]
  wire [4:0] _T_65165; // @[Modules.scala 150:74:@11236.4]
  wire [5:0] _T_65168; // @[Modules.scala 150:103:@11238.4]
  wire [4:0] _T_65169; // @[Modules.scala 150:103:@11239.4]
  wire [4:0] _T_65170; // @[Modules.scala 150:103:@11240.4]
  wire [5:0] _T_65188; // @[Modules.scala 151:80:@11255.4]
  wire [6:0] _T_65189; // @[Modules.scala 150:103:@11256.4]
  wire [5:0] _T_65190; // @[Modules.scala 150:103:@11257.4]
  wire [5:0] _T_65191; // @[Modules.scala 150:103:@11258.4]
  wire [5:0] _T_65193; // @[Modules.scala 150:74:@11260.4]
  wire [5:0] _T_65195; // @[Modules.scala 151:80:@11261.4]
  wire [6:0] _T_65196; // @[Modules.scala 150:103:@11262.4]
  wire [5:0] _T_65197; // @[Modules.scala 150:103:@11263.4]
  wire [5:0] _T_65198; // @[Modules.scala 150:103:@11264.4]
  wire [5:0] _T_65200; // @[Modules.scala 150:74:@11266.4]
  wire [6:0] _T_65203; // @[Modules.scala 150:103:@11268.4]
  wire [5:0] _T_65204; // @[Modules.scala 150:103:@11269.4]
  wire [5:0] _T_65205; // @[Modules.scala 150:103:@11270.4]
  wire [5:0] _T_65221; // @[Modules.scala 150:74:@11284.4]
  wire [6:0] _T_65224; // @[Modules.scala 150:103:@11286.4]
  wire [5:0] _T_65225; // @[Modules.scala 150:103:@11287.4]
  wire [5:0] _T_65226; // @[Modules.scala 150:103:@11288.4]
  wire [4:0] _T_65230; // @[Modules.scala 151:80:@11291.4]
  wire [5:0] _T_65231; // @[Modules.scala 150:103:@11292.4]
  wire [4:0] _T_65232; // @[Modules.scala 150:103:@11293.4]
  wire [4:0] _T_65233; // @[Modules.scala 150:103:@11294.4]
  wire [5:0] _GEN_273; // @[Modules.scala 150:103:@11298.4]
  wire [6:0] _T_65238; // @[Modules.scala 150:103:@11298.4]
  wire [5:0] _T_65239; // @[Modules.scala 150:103:@11299.4]
  wire [5:0] _T_65240; // @[Modules.scala 150:103:@11300.4]
  wire [5:0] _T_65245; // @[Modules.scala 150:103:@11304.4]
  wire [4:0] _T_65246; // @[Modules.scala 150:103:@11305.4]
  wire [4:0] _T_65247; // @[Modules.scala 150:103:@11306.4]
  wire [4:0] _T_65251; // @[Modules.scala 151:80:@11309.4]
  wire [5:0] _T_65252; // @[Modules.scala 150:103:@11310.4]
  wire [4:0] _T_65253; // @[Modules.scala 150:103:@11311.4]
  wire [4:0] _T_65254; // @[Modules.scala 150:103:@11312.4]
  wire [5:0] _T_65259; // @[Modules.scala 150:103:@11316.4]
  wire [4:0] _T_65260; // @[Modules.scala 150:103:@11317.4]
  wire [4:0] _T_65261; // @[Modules.scala 150:103:@11318.4]
  wire [4:0] _T_65265; // @[Modules.scala 151:80:@11321.4]
  wire [5:0] _T_65266; // @[Modules.scala 150:103:@11322.4]
  wire [4:0] _T_65267; // @[Modules.scala 150:103:@11323.4]
  wire [4:0] _T_65268; // @[Modules.scala 150:103:@11324.4]
  wire [5:0] _T_65280; // @[Modules.scala 150:103:@11334.4]
  wire [4:0] _T_65281; // @[Modules.scala 150:103:@11335.4]
  wire [4:0] _T_65282; // @[Modules.scala 150:103:@11336.4]
  wire [5:0] _GEN_274; // @[Modules.scala 150:103:@11340.4]
  wire [6:0] _T_65287; // @[Modules.scala 150:103:@11340.4]
  wire [5:0] _T_65288; // @[Modules.scala 150:103:@11341.4]
  wire [5:0] _T_65289; // @[Modules.scala 150:103:@11342.4]
  wire [6:0] _T_65301; // @[Modules.scala 150:103:@11352.4]
  wire [5:0] _T_65302; // @[Modules.scala 150:103:@11353.4]
  wire [5:0] _T_65303; // @[Modules.scala 150:103:@11354.4]
  wire [6:0] _T_65308; // @[Modules.scala 150:103:@11358.4]
  wire [5:0] _T_65309; // @[Modules.scala 150:103:@11359.4]
  wire [5:0] _T_65310; // @[Modules.scala 150:103:@11360.4]
  wire [4:0] _T_65314; // @[Modules.scala 151:80:@11363.4]
  wire [5:0] _GEN_275; // @[Modules.scala 150:103:@11364.4]
  wire [6:0] _T_65315; // @[Modules.scala 150:103:@11364.4]
  wire [5:0] _T_65316; // @[Modules.scala 150:103:@11365.4]
  wire [5:0] _T_65317; // @[Modules.scala 150:103:@11366.4]
  wire [6:0] _T_65329; // @[Modules.scala 150:103:@11376.4]
  wire [5:0] _T_65330; // @[Modules.scala 150:103:@11377.4]
  wire [5:0] _T_65331; // @[Modules.scala 150:103:@11378.4]
  wire [5:0] _T_65336; // @[Modules.scala 150:103:@11382.4]
  wire [4:0] _T_65337; // @[Modules.scala 150:103:@11383.4]
  wire [4:0] _T_65338; // @[Modules.scala 150:103:@11384.4]
  wire [4:0] _T_65340; // @[Modules.scala 150:74:@11386.4]
  wire [4:0] _T_65342; // @[Modules.scala 151:80:@11387.4]
  wire [5:0] _T_65343; // @[Modules.scala 150:103:@11388.4]
  wire [4:0] _T_65344; // @[Modules.scala 150:103:@11389.4]
  wire [4:0] _T_65345; // @[Modules.scala 150:103:@11390.4]
  wire [4:0] _T_65347; // @[Modules.scala 150:74:@11392.4]
  wire [5:0] _T_65350; // @[Modules.scala 150:103:@11394.4]
  wire [4:0] _T_65351; // @[Modules.scala 150:103:@11395.4]
  wire [4:0] _T_65352; // @[Modules.scala 150:103:@11396.4]
  wire [4:0] _T_65354; // @[Modules.scala 150:74:@11398.4]
  wire [5:0] _T_65357; // @[Modules.scala 150:103:@11400.4]
  wire [4:0] _T_65358; // @[Modules.scala 150:103:@11401.4]
  wire [4:0] _T_65359; // @[Modules.scala 150:103:@11402.4]
  wire [5:0] _GEN_277; // @[Modules.scala 150:103:@11412.4]
  wire [6:0] _T_65371; // @[Modules.scala 150:103:@11412.4]
  wire [5:0] _T_65372; // @[Modules.scala 150:103:@11413.4]
  wire [5:0] _T_65373; // @[Modules.scala 150:103:@11414.4]
  wire [5:0] _T_65382; // @[Modules.scala 150:74:@11422.4]
  wire [5:0] _T_65384; // @[Modules.scala 151:80:@11423.4]
  wire [6:0] _T_65385; // @[Modules.scala 150:103:@11424.4]
  wire [5:0] _T_65386; // @[Modules.scala 150:103:@11425.4]
  wire [5:0] _T_65387; // @[Modules.scala 150:103:@11426.4]
  wire [5:0] _T_65392; // @[Modules.scala 150:103:@11430.4]
  wire [4:0] _T_65393; // @[Modules.scala 150:103:@11431.4]
  wire [4:0] _T_65394; // @[Modules.scala 150:103:@11432.4]
  wire [6:0] _T_65399; // @[Modules.scala 150:103:@11436.4]
  wire [5:0] _T_65400; // @[Modules.scala 150:103:@11437.4]
  wire [5:0] _T_65401; // @[Modules.scala 150:103:@11438.4]
  wire [6:0] _T_65406; // @[Modules.scala 150:103:@11442.4]
  wire [5:0] _T_65407; // @[Modules.scala 150:103:@11443.4]
  wire [5:0] _T_65408; // @[Modules.scala 150:103:@11444.4]
  wire [4:0] _T_65410; // @[Modules.scala 150:74:@11446.4]
  wire [5:0] _T_65413; // @[Modules.scala 150:103:@11448.4]
  wire [4:0] _T_65414; // @[Modules.scala 150:103:@11449.4]
  wire [4:0] _T_65415; // @[Modules.scala 150:103:@11450.4]
  wire [5:0] _T_65455; // @[Modules.scala 150:103:@11484.4]
  wire [4:0] _T_65456; // @[Modules.scala 150:103:@11485.4]
  wire [4:0] _T_65457; // @[Modules.scala 150:103:@11486.4]
  wire [5:0] _GEN_278; // @[Modules.scala 150:103:@11496.4]
  wire [6:0] _T_65469; // @[Modules.scala 150:103:@11496.4]
  wire [5:0] _T_65470; // @[Modules.scala 150:103:@11497.4]
  wire [5:0] _T_65471; // @[Modules.scala 150:103:@11498.4]
  wire [4:0] _T_65475; // @[Modules.scala 151:80:@11501.4]
  wire [5:0] _T_65476; // @[Modules.scala 150:103:@11502.4]
  wire [4:0] _T_65477; // @[Modules.scala 150:103:@11503.4]
  wire [4:0] _T_65478; // @[Modules.scala 150:103:@11504.4]
  wire [5:0] _T_65525; // @[Modules.scala 150:103:@11544.4]
  wire [4:0] _T_65526; // @[Modules.scala 150:103:@11545.4]
  wire [4:0] _T_65527; // @[Modules.scala 150:103:@11546.4]
  wire [4:0] _T_65529; // @[Modules.scala 150:74:@11548.4]
  wire [5:0] _T_65532; // @[Modules.scala 150:103:@11550.4]
  wire [4:0] _T_65533; // @[Modules.scala 150:103:@11551.4]
  wire [4:0] _T_65534; // @[Modules.scala 150:103:@11552.4]
  wire [13:0] buffer_3_2; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65540; // @[Modules.scala 160:64:@11560.4]
  wire [13:0] _T_65541; // @[Modules.scala 160:64:@11561.4]
  wire [13:0] buffer_3_315; // @[Modules.scala 160:64:@11562.4]
  wire [13:0] buffer_3_4; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65543; // @[Modules.scala 160:64:@11564.4]
  wire [13:0] _T_65544; // @[Modules.scala 160:64:@11565.4]
  wire [13:0] buffer_3_316; // @[Modules.scala 160:64:@11566.4]
  wire [13:0] buffer_3_6; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_7; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65546; // @[Modules.scala 160:64:@11568.4]
  wire [13:0] _T_65547; // @[Modules.scala 160:64:@11569.4]
  wire [13:0] buffer_3_317; // @[Modules.scala 160:64:@11570.4]
  wire [13:0] buffer_3_8; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65549; // @[Modules.scala 160:64:@11572.4]
  wire [13:0] _T_65550; // @[Modules.scala 160:64:@11573.4]
  wire [13:0] buffer_3_318; // @[Modules.scala 160:64:@11574.4]
  wire [13:0] buffer_3_10; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65552; // @[Modules.scala 160:64:@11576.4]
  wire [13:0] _T_65553; // @[Modules.scala 160:64:@11577.4]
  wire [13:0] buffer_3_319; // @[Modules.scala 160:64:@11578.4]
  wire [13:0] buffer_3_12; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65555; // @[Modules.scala 160:64:@11580.4]
  wire [13:0] _T_65556; // @[Modules.scala 160:64:@11581.4]
  wire [13:0] buffer_3_320; // @[Modules.scala 160:64:@11582.4]
  wire [13:0] buffer_3_17; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65561; // @[Modules.scala 160:64:@11588.4]
  wire [13:0] _T_65562; // @[Modules.scala 160:64:@11589.4]
  wire [13:0] buffer_3_322; // @[Modules.scala 160:64:@11590.4]
  wire [13:0] buffer_3_18; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65564; // @[Modules.scala 160:64:@11592.4]
  wire [13:0] _T_65565; // @[Modules.scala 160:64:@11593.4]
  wire [13:0] buffer_3_323; // @[Modules.scala 160:64:@11594.4]
  wire [13:0] buffer_3_20; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65567; // @[Modules.scala 160:64:@11596.4]
  wire [13:0] _T_65568; // @[Modules.scala 160:64:@11597.4]
  wire [13:0] buffer_3_324; // @[Modules.scala 160:64:@11598.4]
  wire [13:0] buffer_3_22; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_23; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65570; // @[Modules.scala 160:64:@11600.4]
  wire [13:0] _T_65571; // @[Modules.scala 160:64:@11601.4]
  wire [13:0] buffer_3_325; // @[Modules.scala 160:64:@11602.4]
  wire [13:0] buffer_3_24; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_25; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65573; // @[Modules.scala 160:64:@11604.4]
  wire [13:0] _T_65574; // @[Modules.scala 160:64:@11605.4]
  wire [13:0] buffer_3_326; // @[Modules.scala 160:64:@11606.4]
  wire [13:0] buffer_3_26; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65576; // @[Modules.scala 160:64:@11608.4]
  wire [13:0] _T_65577; // @[Modules.scala 160:64:@11609.4]
  wire [13:0] buffer_3_327; // @[Modules.scala 160:64:@11610.4]
  wire [13:0] buffer_3_28; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_29; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65579; // @[Modules.scala 160:64:@11612.4]
  wire [13:0] _T_65580; // @[Modules.scala 160:64:@11613.4]
  wire [13:0] buffer_3_328; // @[Modules.scala 160:64:@11614.4]
  wire [13:0] buffer_3_30; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_31; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65582; // @[Modules.scala 160:64:@11616.4]
  wire [13:0] _T_65583; // @[Modules.scala 160:64:@11617.4]
  wire [13:0] buffer_3_329; // @[Modules.scala 160:64:@11618.4]
  wire [13:0] buffer_3_32; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65585; // @[Modules.scala 160:64:@11620.4]
  wire [13:0] _T_65586; // @[Modules.scala 160:64:@11621.4]
  wire [13:0] buffer_3_330; // @[Modules.scala 160:64:@11622.4]
  wire [13:0] buffer_3_34; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65588; // @[Modules.scala 160:64:@11624.4]
  wire [13:0] _T_65589; // @[Modules.scala 160:64:@11625.4]
  wire [13:0] buffer_3_331; // @[Modules.scala 160:64:@11626.4]
  wire [13:0] buffer_3_36; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_37; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65591; // @[Modules.scala 160:64:@11628.4]
  wire [13:0] _T_65592; // @[Modules.scala 160:64:@11629.4]
  wire [13:0] buffer_3_332; // @[Modules.scala 160:64:@11630.4]
  wire [13:0] buffer_3_38; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_39; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65594; // @[Modules.scala 160:64:@11632.4]
  wire [13:0] _T_65595; // @[Modules.scala 160:64:@11633.4]
  wire [13:0] buffer_3_333; // @[Modules.scala 160:64:@11634.4]
  wire [13:0] buffer_3_40; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65597; // @[Modules.scala 160:64:@11636.4]
  wire [13:0] _T_65598; // @[Modules.scala 160:64:@11637.4]
  wire [13:0] buffer_3_334; // @[Modules.scala 160:64:@11638.4]
  wire [13:0] buffer_3_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65600; // @[Modules.scala 160:64:@11640.4]
  wire [13:0] _T_65601; // @[Modules.scala 160:64:@11641.4]
  wire [13:0] buffer_3_335; // @[Modules.scala 160:64:@11642.4]
  wire [13:0] buffer_3_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65603; // @[Modules.scala 160:64:@11644.4]
  wire [13:0] _T_65604; // @[Modules.scala 160:64:@11645.4]
  wire [13:0] buffer_3_336; // @[Modules.scala 160:64:@11646.4]
  wire [13:0] buffer_3_46; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65606; // @[Modules.scala 160:64:@11648.4]
  wire [13:0] _T_65607; // @[Modules.scala 160:64:@11649.4]
  wire [13:0] buffer_3_337; // @[Modules.scala 160:64:@11650.4]
  wire [13:0] buffer_3_48; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65609; // @[Modules.scala 160:64:@11652.4]
  wire [13:0] _T_65610; // @[Modules.scala 160:64:@11653.4]
  wire [13:0] buffer_3_338; // @[Modules.scala 160:64:@11654.4]
  wire [13:0] buffer_3_50; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65612; // @[Modules.scala 160:64:@11656.4]
  wire [13:0] _T_65613; // @[Modules.scala 160:64:@11657.4]
  wire [13:0] buffer_3_339; // @[Modules.scala 160:64:@11658.4]
  wire [13:0] buffer_3_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65615; // @[Modules.scala 160:64:@11660.4]
  wire [13:0] _T_65616; // @[Modules.scala 160:64:@11661.4]
  wire [13:0] buffer_3_340; // @[Modules.scala 160:64:@11662.4]
  wire [13:0] buffer_3_54; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65618; // @[Modules.scala 160:64:@11664.4]
  wire [13:0] _T_65619; // @[Modules.scala 160:64:@11665.4]
  wire [13:0] buffer_3_341; // @[Modules.scala 160:64:@11666.4]
  wire [13:0] buffer_3_56; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65621; // @[Modules.scala 160:64:@11668.4]
  wire [13:0] _T_65622; // @[Modules.scala 160:64:@11669.4]
  wire [13:0] buffer_3_342; // @[Modules.scala 160:64:@11670.4]
  wire [13:0] buffer_3_58; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65624; // @[Modules.scala 160:64:@11672.4]
  wire [13:0] _T_65625; // @[Modules.scala 160:64:@11673.4]
  wire [13:0] buffer_3_343; // @[Modules.scala 160:64:@11674.4]
  wire [13:0] buffer_3_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65627; // @[Modules.scala 160:64:@11676.4]
  wire [13:0] _T_65628; // @[Modules.scala 160:64:@11677.4]
  wire [13:0] buffer_3_344; // @[Modules.scala 160:64:@11678.4]
  wire [13:0] buffer_3_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65630; // @[Modules.scala 160:64:@11680.4]
  wire [13:0] _T_65631; // @[Modules.scala 160:64:@11681.4]
  wire [13:0] buffer_3_345; // @[Modules.scala 160:64:@11682.4]
  wire [13:0] buffer_3_64; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65633; // @[Modules.scala 160:64:@11684.4]
  wire [13:0] _T_65634; // @[Modules.scala 160:64:@11685.4]
  wire [13:0] buffer_3_346; // @[Modules.scala 160:64:@11686.4]
  wire [13:0] buffer_3_66; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65636; // @[Modules.scala 160:64:@11688.4]
  wire [13:0] _T_65637; // @[Modules.scala 160:64:@11689.4]
  wire [13:0] buffer_3_347; // @[Modules.scala 160:64:@11690.4]
  wire [13:0] buffer_3_68; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65639; // @[Modules.scala 160:64:@11692.4]
  wire [13:0] _T_65640; // @[Modules.scala 160:64:@11693.4]
  wire [13:0] buffer_3_348; // @[Modules.scala 160:64:@11694.4]
  wire [13:0] buffer_3_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65642; // @[Modules.scala 160:64:@11696.4]
  wire [13:0] _T_65643; // @[Modules.scala 160:64:@11697.4]
  wire [13:0] buffer_3_349; // @[Modules.scala 160:64:@11698.4]
  wire [13:0] buffer_3_72; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65645; // @[Modules.scala 160:64:@11700.4]
  wire [13:0] _T_65646; // @[Modules.scala 160:64:@11701.4]
  wire [13:0] buffer_3_350; // @[Modules.scala 160:64:@11702.4]
  wire [13:0] buffer_3_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65648; // @[Modules.scala 160:64:@11704.4]
  wire [13:0] _T_65649; // @[Modules.scala 160:64:@11705.4]
  wire [13:0] buffer_3_351; // @[Modules.scala 160:64:@11706.4]
  wire [13:0] buffer_3_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65651; // @[Modules.scala 160:64:@11708.4]
  wire [13:0] _T_65652; // @[Modules.scala 160:64:@11709.4]
  wire [13:0] buffer_3_352; // @[Modules.scala 160:64:@11710.4]
  wire [13:0] buffer_3_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65654; // @[Modules.scala 160:64:@11712.4]
  wire [13:0] _T_65655; // @[Modules.scala 160:64:@11713.4]
  wire [13:0] buffer_3_353; // @[Modules.scala 160:64:@11714.4]
  wire [13:0] buffer_3_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65657; // @[Modules.scala 160:64:@11716.4]
  wire [13:0] _T_65658; // @[Modules.scala 160:64:@11717.4]
  wire [13:0] buffer_3_354; // @[Modules.scala 160:64:@11718.4]
  wire [13:0] buffer_3_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65663; // @[Modules.scala 160:64:@11724.4]
  wire [13:0] _T_65664; // @[Modules.scala 160:64:@11725.4]
  wire [13:0] buffer_3_356; // @[Modules.scala 160:64:@11726.4]
  wire [13:0] buffer_3_86; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65666; // @[Modules.scala 160:64:@11728.4]
  wire [13:0] _T_65667; // @[Modules.scala 160:64:@11729.4]
  wire [13:0] buffer_3_357; // @[Modules.scala 160:64:@11730.4]
  wire [13:0] buffer_3_89; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65669; // @[Modules.scala 160:64:@11732.4]
  wire [13:0] _T_65670; // @[Modules.scala 160:64:@11733.4]
  wire [13:0] buffer_3_358; // @[Modules.scala 160:64:@11734.4]
  wire [13:0] buffer_3_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65672; // @[Modules.scala 160:64:@11736.4]
  wire [13:0] _T_65673; // @[Modules.scala 160:64:@11737.4]
  wire [13:0] buffer_3_359; // @[Modules.scala 160:64:@11738.4]
  wire [13:0] buffer_3_92; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65675; // @[Modules.scala 160:64:@11740.4]
  wire [13:0] _T_65676; // @[Modules.scala 160:64:@11741.4]
  wire [13:0] buffer_3_360; // @[Modules.scala 160:64:@11742.4]
  wire [13:0] buffer_3_94; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65678; // @[Modules.scala 160:64:@11744.4]
  wire [13:0] _T_65679; // @[Modules.scala 160:64:@11745.4]
  wire [13:0] buffer_3_361; // @[Modules.scala 160:64:@11746.4]
  wire [13:0] buffer_3_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65681; // @[Modules.scala 160:64:@11748.4]
  wire [13:0] _T_65682; // @[Modules.scala 160:64:@11749.4]
  wire [13:0] buffer_3_362; // @[Modules.scala 160:64:@11750.4]
  wire [13:0] buffer_3_98; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_99; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65684; // @[Modules.scala 160:64:@11752.4]
  wire [13:0] _T_65685; // @[Modules.scala 160:64:@11753.4]
  wire [13:0] buffer_3_363; // @[Modules.scala 160:64:@11754.4]
  wire [13:0] buffer_3_102; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_103; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65690; // @[Modules.scala 160:64:@11760.4]
  wire [13:0] _T_65691; // @[Modules.scala 160:64:@11761.4]
  wire [13:0] buffer_3_365; // @[Modules.scala 160:64:@11762.4]
  wire [13:0] buffer_3_104; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65693; // @[Modules.scala 160:64:@11764.4]
  wire [13:0] _T_65694; // @[Modules.scala 160:64:@11765.4]
  wire [13:0] buffer_3_366; // @[Modules.scala 160:64:@11766.4]
  wire [13:0] buffer_3_106; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65696; // @[Modules.scala 160:64:@11768.4]
  wire [13:0] _T_65697; // @[Modules.scala 160:64:@11769.4]
  wire [13:0] buffer_3_367; // @[Modules.scala 160:64:@11770.4]
  wire [13:0] buffer_3_108; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_109; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65699; // @[Modules.scala 160:64:@11772.4]
  wire [13:0] _T_65700; // @[Modules.scala 160:64:@11773.4]
  wire [13:0] buffer_3_368; // @[Modules.scala 160:64:@11774.4]
  wire [13:0] buffer_3_110; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65702; // @[Modules.scala 160:64:@11776.4]
  wire [13:0] _T_65703; // @[Modules.scala 160:64:@11777.4]
  wire [13:0] buffer_3_369; // @[Modules.scala 160:64:@11778.4]
  wire [13:0] buffer_3_112; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65705; // @[Modules.scala 160:64:@11780.4]
  wire [13:0] _T_65706; // @[Modules.scala 160:64:@11781.4]
  wire [13:0] buffer_3_370; // @[Modules.scala 160:64:@11782.4]
  wire [13:0] buffer_3_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65711; // @[Modules.scala 160:64:@11788.4]
  wire [13:0] _T_65712; // @[Modules.scala 160:64:@11789.4]
  wire [13:0] buffer_3_372; // @[Modules.scala 160:64:@11790.4]
  wire [13:0] buffer_3_118; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_119; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65714; // @[Modules.scala 160:64:@11792.4]
  wire [13:0] _T_65715; // @[Modules.scala 160:64:@11793.4]
  wire [13:0] buffer_3_373; // @[Modules.scala 160:64:@11794.4]
  wire [13:0] buffer_3_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65717; // @[Modules.scala 160:64:@11796.4]
  wire [13:0] _T_65718; // @[Modules.scala 160:64:@11797.4]
  wire [13:0] buffer_3_374; // @[Modules.scala 160:64:@11798.4]
  wire [13:0] buffer_3_122; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65720; // @[Modules.scala 160:64:@11800.4]
  wire [13:0] _T_65721; // @[Modules.scala 160:64:@11801.4]
  wire [13:0] buffer_3_375; // @[Modules.scala 160:64:@11802.4]
  wire [13:0] buffer_3_124; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65723; // @[Modules.scala 160:64:@11804.4]
  wire [13:0] _T_65724; // @[Modules.scala 160:64:@11805.4]
  wire [13:0] buffer_3_376; // @[Modules.scala 160:64:@11806.4]
  wire [13:0] buffer_3_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65726; // @[Modules.scala 160:64:@11808.4]
  wire [13:0] _T_65727; // @[Modules.scala 160:64:@11809.4]
  wire [13:0] buffer_3_377; // @[Modules.scala 160:64:@11810.4]
  wire [14:0] _T_65729; // @[Modules.scala 160:64:@11812.4]
  wire [13:0] _T_65730; // @[Modules.scala 160:64:@11813.4]
  wire [13:0] buffer_3_378; // @[Modules.scala 160:64:@11814.4]
  wire [13:0] buffer_3_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65732; // @[Modules.scala 160:64:@11816.4]
  wire [13:0] _T_65733; // @[Modules.scala 160:64:@11817.4]
  wire [13:0] buffer_3_379; // @[Modules.scala 160:64:@11818.4]
  wire [13:0] buffer_3_132; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65735; // @[Modules.scala 160:64:@11820.4]
  wire [13:0] _T_65736; // @[Modules.scala 160:64:@11821.4]
  wire [13:0] buffer_3_380; // @[Modules.scala 160:64:@11822.4]
  wire [13:0] buffer_3_134; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65738; // @[Modules.scala 160:64:@11824.4]
  wire [13:0] _T_65739; // @[Modules.scala 160:64:@11825.4]
  wire [13:0] buffer_3_381; // @[Modules.scala 160:64:@11826.4]
  wire [14:0] _T_65741; // @[Modules.scala 160:64:@11828.4]
  wire [13:0] _T_65742; // @[Modules.scala 160:64:@11829.4]
  wire [13:0] buffer_3_382; // @[Modules.scala 160:64:@11830.4]
  wire [14:0] _T_65744; // @[Modules.scala 160:64:@11832.4]
  wire [13:0] _T_65745; // @[Modules.scala 160:64:@11833.4]
  wire [13:0] buffer_3_383; // @[Modules.scala 160:64:@11834.4]
  wire [13:0] buffer_3_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65747; // @[Modules.scala 160:64:@11836.4]
  wire [13:0] _T_65748; // @[Modules.scala 160:64:@11837.4]
  wire [13:0] buffer_3_384; // @[Modules.scala 160:64:@11838.4]
  wire [13:0] buffer_3_142; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_143; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65750; // @[Modules.scala 160:64:@11840.4]
  wire [13:0] _T_65751; // @[Modules.scala 160:64:@11841.4]
  wire [13:0] buffer_3_385; // @[Modules.scala 160:64:@11842.4]
  wire [13:0] buffer_3_144; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65753; // @[Modules.scala 160:64:@11844.4]
  wire [13:0] _T_65754; // @[Modules.scala 160:64:@11845.4]
  wire [13:0] buffer_3_386; // @[Modules.scala 160:64:@11846.4]
  wire [13:0] buffer_3_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65756; // @[Modules.scala 160:64:@11848.4]
  wire [13:0] _T_65757; // @[Modules.scala 160:64:@11849.4]
  wire [13:0] buffer_3_387; // @[Modules.scala 160:64:@11850.4]
  wire [13:0] buffer_3_152; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65765; // @[Modules.scala 160:64:@11860.4]
  wire [13:0] _T_65766; // @[Modules.scala 160:64:@11861.4]
  wire [13:0] buffer_3_390; // @[Modules.scala 160:64:@11862.4]
  wire [13:0] buffer_3_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65768; // @[Modules.scala 160:64:@11864.4]
  wire [13:0] _T_65769; // @[Modules.scala 160:64:@11865.4]
  wire [13:0] buffer_3_391; // @[Modules.scala 160:64:@11866.4]
  wire [13:0] buffer_3_156; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65771; // @[Modules.scala 160:64:@11868.4]
  wire [13:0] _T_65772; // @[Modules.scala 160:64:@11869.4]
  wire [13:0] buffer_3_392; // @[Modules.scala 160:64:@11870.4]
  wire [13:0] buffer_3_158; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65774; // @[Modules.scala 160:64:@11872.4]
  wire [13:0] _T_65775; // @[Modules.scala 160:64:@11873.4]
  wire [13:0] buffer_3_393; // @[Modules.scala 160:64:@11874.4]
  wire [14:0] _T_65777; // @[Modules.scala 160:64:@11876.4]
  wire [13:0] _T_65778; // @[Modules.scala 160:64:@11877.4]
  wire [13:0] buffer_3_394; // @[Modules.scala 160:64:@11878.4]
  wire [13:0] buffer_3_163; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65780; // @[Modules.scala 160:64:@11880.4]
  wire [13:0] _T_65781; // @[Modules.scala 160:64:@11881.4]
  wire [13:0] buffer_3_395; // @[Modules.scala 160:64:@11882.4]
  wire [13:0] buffer_3_164; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65783; // @[Modules.scala 160:64:@11884.4]
  wire [13:0] _T_65784; // @[Modules.scala 160:64:@11885.4]
  wire [13:0] buffer_3_396; // @[Modules.scala 160:64:@11886.4]
  wire [13:0] buffer_3_166; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65786; // @[Modules.scala 160:64:@11888.4]
  wire [13:0] _T_65787; // @[Modules.scala 160:64:@11889.4]
  wire [13:0] buffer_3_397; // @[Modules.scala 160:64:@11890.4]
  wire [13:0] buffer_3_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65789; // @[Modules.scala 160:64:@11892.4]
  wire [13:0] _T_65790; // @[Modules.scala 160:64:@11893.4]
  wire [13:0] buffer_3_398; // @[Modules.scala 160:64:@11894.4]
  wire [13:0] buffer_3_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65792; // @[Modules.scala 160:64:@11896.4]
  wire [13:0] _T_65793; // @[Modules.scala 160:64:@11897.4]
  wire [13:0] buffer_3_399; // @[Modules.scala 160:64:@11898.4]
  wire [13:0] buffer_3_172; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65795; // @[Modules.scala 160:64:@11900.4]
  wire [13:0] _T_65796; // @[Modules.scala 160:64:@11901.4]
  wire [13:0] buffer_3_400; // @[Modules.scala 160:64:@11902.4]
  wire [13:0] buffer_3_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65798; // @[Modules.scala 160:64:@11904.4]
  wire [13:0] _T_65799; // @[Modules.scala 160:64:@11905.4]
  wire [13:0] buffer_3_401; // @[Modules.scala 160:64:@11906.4]
  wire [13:0] buffer_3_176; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65801; // @[Modules.scala 160:64:@11908.4]
  wire [13:0] _T_65802; // @[Modules.scala 160:64:@11909.4]
  wire [13:0] buffer_3_402; // @[Modules.scala 160:64:@11910.4]
  wire [14:0] _T_65804; // @[Modules.scala 160:64:@11912.4]
  wire [13:0] _T_65805; // @[Modules.scala 160:64:@11913.4]
  wire [13:0] buffer_3_403; // @[Modules.scala 160:64:@11914.4]
  wire [13:0] buffer_3_180; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65807; // @[Modules.scala 160:64:@11916.4]
  wire [13:0] _T_65808; // @[Modules.scala 160:64:@11917.4]
  wire [13:0] buffer_3_404; // @[Modules.scala 160:64:@11918.4]
  wire [13:0] buffer_3_182; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65810; // @[Modules.scala 160:64:@11920.4]
  wire [13:0] _T_65811; // @[Modules.scala 160:64:@11921.4]
  wire [13:0] buffer_3_405; // @[Modules.scala 160:64:@11922.4]
  wire [13:0] buffer_3_184; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65813; // @[Modules.scala 160:64:@11924.4]
  wire [13:0] _T_65814; // @[Modules.scala 160:64:@11925.4]
  wire [13:0] buffer_3_406; // @[Modules.scala 160:64:@11926.4]
  wire [13:0] buffer_3_186; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65816; // @[Modules.scala 160:64:@11928.4]
  wire [13:0] _T_65817; // @[Modules.scala 160:64:@11929.4]
  wire [13:0] buffer_3_407; // @[Modules.scala 160:64:@11930.4]
  wire [13:0] buffer_3_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65819; // @[Modules.scala 160:64:@11932.4]
  wire [13:0] _T_65820; // @[Modules.scala 160:64:@11933.4]
  wire [13:0] buffer_3_408; // @[Modules.scala 160:64:@11934.4]
  wire [13:0] buffer_3_190; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65822; // @[Modules.scala 160:64:@11936.4]
  wire [13:0] _T_65823; // @[Modules.scala 160:64:@11937.4]
  wire [13:0] buffer_3_409; // @[Modules.scala 160:64:@11938.4]
  wire [13:0] buffer_3_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65825; // @[Modules.scala 160:64:@11940.4]
  wire [13:0] _T_65826; // @[Modules.scala 160:64:@11941.4]
  wire [13:0] buffer_3_410; // @[Modules.scala 160:64:@11942.4]
  wire [13:0] buffer_3_194; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65828; // @[Modules.scala 160:64:@11944.4]
  wire [13:0] _T_65829; // @[Modules.scala 160:64:@11945.4]
  wire [13:0] buffer_3_411; // @[Modules.scala 160:64:@11946.4]
  wire [13:0] buffer_3_196; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65831; // @[Modules.scala 160:64:@11948.4]
  wire [13:0] _T_65832; // @[Modules.scala 160:64:@11949.4]
  wire [13:0] buffer_3_412; // @[Modules.scala 160:64:@11950.4]
  wire [14:0] _T_65834; // @[Modules.scala 160:64:@11952.4]
  wire [13:0] _T_65835; // @[Modules.scala 160:64:@11953.4]
  wire [13:0] buffer_3_413; // @[Modules.scala 160:64:@11954.4]
  wire [13:0] buffer_3_200; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65837; // @[Modules.scala 160:64:@11956.4]
  wire [13:0] _T_65838; // @[Modules.scala 160:64:@11957.4]
  wire [13:0] buffer_3_414; // @[Modules.scala 160:64:@11958.4]
  wire [13:0] buffer_3_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65840; // @[Modules.scala 160:64:@11960.4]
  wire [13:0] _T_65841; // @[Modules.scala 160:64:@11961.4]
  wire [13:0] buffer_3_415; // @[Modules.scala 160:64:@11962.4]
  wire [13:0] buffer_3_204; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65843; // @[Modules.scala 160:64:@11964.4]
  wire [13:0] _T_65844; // @[Modules.scala 160:64:@11965.4]
  wire [13:0] buffer_3_416; // @[Modules.scala 160:64:@11966.4]
  wire [13:0] buffer_3_206; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65846; // @[Modules.scala 160:64:@11968.4]
  wire [13:0] _T_65847; // @[Modules.scala 160:64:@11969.4]
  wire [13:0] buffer_3_417; // @[Modules.scala 160:64:@11970.4]
  wire [13:0] buffer_3_208; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65849; // @[Modules.scala 160:64:@11972.4]
  wire [13:0] _T_65850; // @[Modules.scala 160:64:@11973.4]
  wire [13:0] buffer_3_418; // @[Modules.scala 160:64:@11974.4]
  wire [13:0] buffer_3_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65852; // @[Modules.scala 160:64:@11976.4]
  wire [13:0] _T_65853; // @[Modules.scala 160:64:@11977.4]
  wire [13:0] buffer_3_419; // @[Modules.scala 160:64:@11978.4]
  wire [13:0] buffer_3_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65855; // @[Modules.scala 160:64:@11980.4]
  wire [13:0] _T_65856; // @[Modules.scala 160:64:@11981.4]
  wire [13:0] buffer_3_420; // @[Modules.scala 160:64:@11982.4]
  wire [13:0] buffer_3_214; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65858; // @[Modules.scala 160:64:@11984.4]
  wire [13:0] _T_65859; // @[Modules.scala 160:64:@11985.4]
  wire [13:0] buffer_3_421; // @[Modules.scala 160:64:@11986.4]
  wire [13:0] buffer_3_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65861; // @[Modules.scala 160:64:@11988.4]
  wire [13:0] _T_65862; // @[Modules.scala 160:64:@11989.4]
  wire [13:0] buffer_3_422; // @[Modules.scala 160:64:@11990.4]
  wire [13:0] buffer_3_218; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65864; // @[Modules.scala 160:64:@11992.4]
  wire [13:0] _T_65865; // @[Modules.scala 160:64:@11993.4]
  wire [13:0] buffer_3_423; // @[Modules.scala 160:64:@11994.4]
  wire [13:0] buffer_3_220; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65867; // @[Modules.scala 160:64:@11996.4]
  wire [13:0] _T_65868; // @[Modules.scala 160:64:@11997.4]
  wire [13:0] buffer_3_424; // @[Modules.scala 160:64:@11998.4]
  wire [13:0] buffer_3_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65870; // @[Modules.scala 160:64:@12000.4]
  wire [13:0] _T_65871; // @[Modules.scala 160:64:@12001.4]
  wire [13:0] buffer_3_425; // @[Modules.scala 160:64:@12002.4]
  wire [13:0] buffer_3_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65873; // @[Modules.scala 160:64:@12004.4]
  wire [13:0] _T_65874; // @[Modules.scala 160:64:@12005.4]
  wire [13:0] buffer_3_426; // @[Modules.scala 160:64:@12006.4]
  wire [13:0] buffer_3_226; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65876; // @[Modules.scala 160:64:@12008.4]
  wire [13:0] _T_65877; // @[Modules.scala 160:64:@12009.4]
  wire [13:0] buffer_3_427; // @[Modules.scala 160:64:@12010.4]
  wire [13:0] buffer_3_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65879; // @[Modules.scala 160:64:@12012.4]
  wire [13:0] _T_65880; // @[Modules.scala 160:64:@12013.4]
  wire [13:0] buffer_3_428; // @[Modules.scala 160:64:@12014.4]
  wire [13:0] buffer_3_232; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65885; // @[Modules.scala 160:64:@12020.4]
  wire [13:0] _T_65886; // @[Modules.scala 160:64:@12021.4]
  wire [13:0] buffer_3_430; // @[Modules.scala 160:64:@12022.4]
  wire [13:0] buffer_3_234; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65888; // @[Modules.scala 160:64:@12024.4]
  wire [13:0] _T_65889; // @[Modules.scala 160:64:@12025.4]
  wire [13:0] buffer_3_431; // @[Modules.scala 160:64:@12026.4]
  wire [13:0] buffer_3_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65891; // @[Modules.scala 160:64:@12028.4]
  wire [13:0] _T_65892; // @[Modules.scala 160:64:@12029.4]
  wire [13:0] buffer_3_432; // @[Modules.scala 160:64:@12030.4]
  wire [14:0] _T_65894; // @[Modules.scala 160:64:@12032.4]
  wire [13:0] _T_65895; // @[Modules.scala 160:64:@12033.4]
  wire [13:0] buffer_3_433; // @[Modules.scala 160:64:@12034.4]
  wire [13:0] buffer_3_240; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65897; // @[Modules.scala 160:64:@12036.4]
  wire [13:0] _T_65898; // @[Modules.scala 160:64:@12037.4]
  wire [13:0] buffer_3_434; // @[Modules.scala 160:64:@12038.4]
  wire [13:0] buffer_3_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65900; // @[Modules.scala 160:64:@12040.4]
  wire [13:0] _T_65901; // @[Modules.scala 160:64:@12041.4]
  wire [13:0] buffer_3_435; // @[Modules.scala 160:64:@12042.4]
  wire [13:0] buffer_3_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65903; // @[Modules.scala 160:64:@12044.4]
  wire [13:0] _T_65904; // @[Modules.scala 160:64:@12045.4]
  wire [13:0] buffer_3_436; // @[Modules.scala 160:64:@12046.4]
  wire [13:0] buffer_3_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65906; // @[Modules.scala 160:64:@12048.4]
  wire [13:0] _T_65907; // @[Modules.scala 160:64:@12049.4]
  wire [13:0] buffer_3_437; // @[Modules.scala 160:64:@12050.4]
  wire [13:0] buffer_3_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65909; // @[Modules.scala 160:64:@12052.4]
  wire [13:0] _T_65910; // @[Modules.scala 160:64:@12053.4]
  wire [13:0] buffer_3_438; // @[Modules.scala 160:64:@12054.4]
  wire [13:0] buffer_3_250; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65912; // @[Modules.scala 160:64:@12056.4]
  wire [13:0] _T_65913; // @[Modules.scala 160:64:@12057.4]
  wire [13:0] buffer_3_439; // @[Modules.scala 160:64:@12058.4]
  wire [13:0] buffer_3_252; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65915; // @[Modules.scala 160:64:@12060.4]
  wire [13:0] _T_65916; // @[Modules.scala 160:64:@12061.4]
  wire [13:0] buffer_3_440; // @[Modules.scala 160:64:@12062.4]
  wire [13:0] buffer_3_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65918; // @[Modules.scala 160:64:@12064.4]
  wire [13:0] _T_65919; // @[Modules.scala 160:64:@12065.4]
  wire [13:0] buffer_3_441; // @[Modules.scala 160:64:@12066.4]
  wire [13:0] buffer_3_256; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65921; // @[Modules.scala 160:64:@12068.4]
  wire [13:0] _T_65922; // @[Modules.scala 160:64:@12069.4]
  wire [13:0] buffer_3_442; // @[Modules.scala 160:64:@12070.4]
  wire [13:0] buffer_3_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65924; // @[Modules.scala 160:64:@12072.4]
  wire [13:0] _T_65925; // @[Modules.scala 160:64:@12073.4]
  wire [13:0] buffer_3_443; // @[Modules.scala 160:64:@12074.4]
  wire [13:0] buffer_3_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65927; // @[Modules.scala 160:64:@12076.4]
  wire [13:0] _T_65928; // @[Modules.scala 160:64:@12077.4]
  wire [13:0] buffer_3_444; // @[Modules.scala 160:64:@12078.4]
  wire [13:0] buffer_3_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65930; // @[Modules.scala 160:64:@12080.4]
  wire [13:0] _T_65931; // @[Modules.scala 160:64:@12081.4]
  wire [13:0] buffer_3_445; // @[Modules.scala 160:64:@12082.4]
  wire [13:0] buffer_3_264; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65933; // @[Modules.scala 160:64:@12084.4]
  wire [13:0] _T_65934; // @[Modules.scala 160:64:@12085.4]
  wire [13:0] buffer_3_446; // @[Modules.scala 160:64:@12086.4]
  wire [14:0] _T_65936; // @[Modules.scala 160:64:@12088.4]
  wire [13:0] _T_65937; // @[Modules.scala 160:64:@12089.4]
  wire [13:0] buffer_3_447; // @[Modules.scala 160:64:@12090.4]
  wire [13:0] buffer_3_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65939; // @[Modules.scala 160:64:@12092.4]
  wire [13:0] _T_65940; // @[Modules.scala 160:64:@12093.4]
  wire [13:0] buffer_3_448; // @[Modules.scala 160:64:@12094.4]
  wire [13:0] buffer_3_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65942; // @[Modules.scala 160:64:@12096.4]
  wire [13:0] _T_65943; // @[Modules.scala 160:64:@12097.4]
  wire [13:0] buffer_3_449; // @[Modules.scala 160:64:@12098.4]
  wire [13:0] buffer_3_272; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65945; // @[Modules.scala 160:64:@12100.4]
  wire [13:0] _T_65946; // @[Modules.scala 160:64:@12101.4]
  wire [13:0] buffer_3_450; // @[Modules.scala 160:64:@12102.4]
  wire [13:0] buffer_3_274; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65948; // @[Modules.scala 160:64:@12104.4]
  wire [13:0] _T_65949; // @[Modules.scala 160:64:@12105.4]
  wire [13:0] buffer_3_451; // @[Modules.scala 160:64:@12106.4]
  wire [13:0] buffer_3_276; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_277; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65951; // @[Modules.scala 160:64:@12108.4]
  wire [13:0] _T_65952; // @[Modules.scala 160:64:@12109.4]
  wire [13:0] buffer_3_452; // @[Modules.scala 160:64:@12110.4]
  wire [13:0] buffer_3_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65954; // @[Modules.scala 160:64:@12112.4]
  wire [13:0] _T_65955; // @[Modules.scala 160:64:@12113.4]
  wire [13:0] buffer_3_453; // @[Modules.scala 160:64:@12114.4]
  wire [13:0] buffer_3_280; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65957; // @[Modules.scala 160:64:@12116.4]
  wire [13:0] _T_65958; // @[Modules.scala 160:64:@12117.4]
  wire [13:0] buffer_3_454; // @[Modules.scala 160:64:@12118.4]
  wire [13:0] buffer_3_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65960; // @[Modules.scala 160:64:@12120.4]
  wire [13:0] _T_65961; // @[Modules.scala 160:64:@12121.4]
  wire [13:0] buffer_3_455; // @[Modules.scala 160:64:@12122.4]
  wire [13:0] buffer_3_284; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_285; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65963; // @[Modules.scala 160:64:@12124.4]
  wire [13:0] _T_65964; // @[Modules.scala 160:64:@12125.4]
  wire [13:0] buffer_3_456; // @[Modules.scala 160:64:@12126.4]
  wire [13:0] buffer_3_286; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_287; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65966; // @[Modules.scala 160:64:@12128.4]
  wire [13:0] _T_65967; // @[Modules.scala 160:64:@12129.4]
  wire [13:0] buffer_3_457; // @[Modules.scala 160:64:@12130.4]
  wire [13:0] buffer_3_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65969; // @[Modules.scala 160:64:@12132.4]
  wire [13:0] _T_65970; // @[Modules.scala 160:64:@12133.4]
  wire [13:0] buffer_3_458; // @[Modules.scala 160:64:@12134.4]
  wire [13:0] buffer_3_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65972; // @[Modules.scala 160:64:@12136.4]
  wire [13:0] _T_65973; // @[Modules.scala 160:64:@12137.4]
  wire [13:0] buffer_3_459; // @[Modules.scala 160:64:@12138.4]
  wire [13:0] buffer_3_292; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65975; // @[Modules.scala 160:64:@12140.4]
  wire [13:0] _T_65976; // @[Modules.scala 160:64:@12141.4]
  wire [13:0] buffer_3_460; // @[Modules.scala 160:64:@12142.4]
  wire [13:0] buffer_3_294; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65978; // @[Modules.scala 160:64:@12144.4]
  wire [13:0] _T_65979; // @[Modules.scala 160:64:@12145.4]
  wire [13:0] buffer_3_461; // @[Modules.scala 160:64:@12146.4]
  wire [14:0] _T_65981; // @[Modules.scala 160:64:@12148.4]
  wire [13:0] _T_65982; // @[Modules.scala 160:64:@12149.4]
  wire [13:0] buffer_3_462; // @[Modules.scala 160:64:@12150.4]
  wire [14:0] _T_65984; // @[Modules.scala 160:64:@12152.4]
  wire [13:0] _T_65985; // @[Modules.scala 160:64:@12153.4]
  wire [13:0] buffer_3_463; // @[Modules.scala 160:64:@12154.4]
  wire [13:0] buffer_3_301; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65987; // @[Modules.scala 160:64:@12156.4]
  wire [13:0] _T_65988; // @[Modules.scala 160:64:@12157.4]
  wire [13:0] buffer_3_464; // @[Modules.scala 160:64:@12158.4]
  wire [13:0] buffer_3_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65990; // @[Modules.scala 160:64:@12160.4]
  wire [13:0] _T_65991; // @[Modules.scala 160:64:@12161.4]
  wire [13:0] buffer_3_465; // @[Modules.scala 160:64:@12162.4]
  wire [13:0] buffer_3_304; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_65993; // @[Modules.scala 160:64:@12164.4]
  wire [13:0] _T_65994; // @[Modules.scala 160:64:@12165.4]
  wire [13:0] buffer_3_466; // @[Modules.scala 160:64:@12166.4]
  wire [14:0] _T_65996; // @[Modules.scala 160:64:@12168.4]
  wire [13:0] _T_65997; // @[Modules.scala 160:64:@12169.4]
  wire [13:0] buffer_3_467; // @[Modules.scala 160:64:@12170.4]
  wire [14:0] _T_65999; // @[Modules.scala 160:64:@12172.4]
  wire [13:0] _T_66000; // @[Modules.scala 160:64:@12173.4]
  wire [13:0] buffer_3_468; // @[Modules.scala 160:64:@12174.4]
  wire [13:0] buffer_3_311; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_66002; // @[Modules.scala 160:64:@12176.4]
  wire [13:0] _T_66003; // @[Modules.scala 160:64:@12177.4]
  wire [13:0] buffer_3_469; // @[Modules.scala 160:64:@12178.4]
  wire [13:0] buffer_3_312; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_3_313; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_66005; // @[Modules.scala 160:64:@12180.4]
  wire [13:0] _T_66006; // @[Modules.scala 160:64:@12181.4]
  wire [13:0] buffer_3_470; // @[Modules.scala 160:64:@12182.4]
  wire [14:0] _T_66008; // @[Modules.scala 166:64:@12184.4]
  wire [13:0] _T_66009; // @[Modules.scala 166:64:@12185.4]
  wire [13:0] buffer_3_471; // @[Modules.scala 166:64:@12186.4]
  wire [14:0] _T_66011; // @[Modules.scala 166:64:@12188.4]
  wire [13:0] _T_66012; // @[Modules.scala 166:64:@12189.4]
  wire [13:0] buffer_3_472; // @[Modules.scala 166:64:@12190.4]
  wire [14:0] _T_66014; // @[Modules.scala 166:64:@12192.4]
  wire [13:0] _T_66015; // @[Modules.scala 166:64:@12193.4]
  wire [13:0] buffer_3_473; // @[Modules.scala 166:64:@12194.4]
  wire [14:0] _T_66017; // @[Modules.scala 166:64:@12196.4]
  wire [13:0] _T_66018; // @[Modules.scala 166:64:@12197.4]
  wire [13:0] buffer_3_474; // @[Modules.scala 166:64:@12198.4]
  wire [14:0] _T_66020; // @[Modules.scala 166:64:@12200.4]
  wire [13:0] _T_66021; // @[Modules.scala 166:64:@12201.4]
  wire [13:0] buffer_3_475; // @[Modules.scala 166:64:@12202.4]
  wire [14:0] _T_66023; // @[Modules.scala 166:64:@12204.4]
  wire [13:0] _T_66024; // @[Modules.scala 166:64:@12205.4]
  wire [13:0] buffer_3_476; // @[Modules.scala 166:64:@12206.4]
  wire [14:0] _T_66026; // @[Modules.scala 166:64:@12208.4]
  wire [13:0] _T_66027; // @[Modules.scala 166:64:@12209.4]
  wire [13:0] buffer_3_477; // @[Modules.scala 166:64:@12210.4]
  wire [14:0] _T_66029; // @[Modules.scala 166:64:@12212.4]
  wire [13:0] _T_66030; // @[Modules.scala 166:64:@12213.4]
  wire [13:0] buffer_3_478; // @[Modules.scala 166:64:@12214.4]
  wire [14:0] _T_66032; // @[Modules.scala 166:64:@12216.4]
  wire [13:0] _T_66033; // @[Modules.scala 166:64:@12217.4]
  wire [13:0] buffer_3_479; // @[Modules.scala 166:64:@12218.4]
  wire [14:0] _T_66035; // @[Modules.scala 166:64:@12220.4]
  wire [13:0] _T_66036; // @[Modules.scala 166:64:@12221.4]
  wire [13:0] buffer_3_480; // @[Modules.scala 166:64:@12222.4]
  wire [14:0] _T_66038; // @[Modules.scala 166:64:@12224.4]
  wire [13:0] _T_66039; // @[Modules.scala 166:64:@12225.4]
  wire [13:0] buffer_3_481; // @[Modules.scala 166:64:@12226.4]
  wire [14:0] _T_66041; // @[Modules.scala 166:64:@12228.4]
  wire [13:0] _T_66042; // @[Modules.scala 166:64:@12229.4]
  wire [13:0] buffer_3_482; // @[Modules.scala 166:64:@12230.4]
  wire [14:0] _T_66044; // @[Modules.scala 166:64:@12232.4]
  wire [13:0] _T_66045; // @[Modules.scala 166:64:@12233.4]
  wire [13:0] buffer_3_483; // @[Modules.scala 166:64:@12234.4]
  wire [14:0] _T_66047; // @[Modules.scala 166:64:@12236.4]
  wire [13:0] _T_66048; // @[Modules.scala 166:64:@12237.4]
  wire [13:0] buffer_3_484; // @[Modules.scala 166:64:@12238.4]
  wire [14:0] _T_66050; // @[Modules.scala 166:64:@12240.4]
  wire [13:0] _T_66051; // @[Modules.scala 166:64:@12241.4]
  wire [13:0] buffer_3_485; // @[Modules.scala 166:64:@12242.4]
  wire [14:0] _T_66053; // @[Modules.scala 166:64:@12244.4]
  wire [13:0] _T_66054; // @[Modules.scala 166:64:@12245.4]
  wire [13:0] buffer_3_486; // @[Modules.scala 166:64:@12246.4]
  wire [14:0] _T_66056; // @[Modules.scala 166:64:@12248.4]
  wire [13:0] _T_66057; // @[Modules.scala 166:64:@12249.4]
  wire [13:0] buffer_3_487; // @[Modules.scala 166:64:@12250.4]
  wire [14:0] _T_66059; // @[Modules.scala 166:64:@12252.4]
  wire [13:0] _T_66060; // @[Modules.scala 166:64:@12253.4]
  wire [13:0] buffer_3_488; // @[Modules.scala 166:64:@12254.4]
  wire [14:0] _T_66062; // @[Modules.scala 166:64:@12256.4]
  wire [13:0] _T_66063; // @[Modules.scala 166:64:@12257.4]
  wire [13:0] buffer_3_489; // @[Modules.scala 166:64:@12258.4]
  wire [14:0] _T_66065; // @[Modules.scala 166:64:@12260.4]
  wire [13:0] _T_66066; // @[Modules.scala 166:64:@12261.4]
  wire [13:0] buffer_3_490; // @[Modules.scala 166:64:@12262.4]
  wire [14:0] _T_66068; // @[Modules.scala 166:64:@12264.4]
  wire [13:0] _T_66069; // @[Modules.scala 166:64:@12265.4]
  wire [13:0] buffer_3_491; // @[Modules.scala 166:64:@12266.4]
  wire [14:0] _T_66071; // @[Modules.scala 166:64:@12268.4]
  wire [13:0] _T_66072; // @[Modules.scala 166:64:@12269.4]
  wire [13:0] buffer_3_492; // @[Modules.scala 166:64:@12270.4]
  wire [14:0] _T_66074; // @[Modules.scala 166:64:@12272.4]
  wire [13:0] _T_66075; // @[Modules.scala 166:64:@12273.4]
  wire [13:0] buffer_3_493; // @[Modules.scala 166:64:@12274.4]
  wire [14:0] _T_66077; // @[Modules.scala 166:64:@12276.4]
  wire [13:0] _T_66078; // @[Modules.scala 166:64:@12277.4]
  wire [13:0] buffer_3_494; // @[Modules.scala 166:64:@12278.4]
  wire [14:0] _T_66080; // @[Modules.scala 166:64:@12280.4]
  wire [13:0] _T_66081; // @[Modules.scala 166:64:@12281.4]
  wire [13:0] buffer_3_495; // @[Modules.scala 166:64:@12282.4]
  wire [14:0] _T_66083; // @[Modules.scala 166:64:@12284.4]
  wire [13:0] _T_66084; // @[Modules.scala 166:64:@12285.4]
  wire [13:0] buffer_3_496; // @[Modules.scala 166:64:@12286.4]
  wire [14:0] _T_66086; // @[Modules.scala 166:64:@12288.4]
  wire [13:0] _T_66087; // @[Modules.scala 166:64:@12289.4]
  wire [13:0] buffer_3_497; // @[Modules.scala 166:64:@12290.4]
  wire [14:0] _T_66089; // @[Modules.scala 166:64:@12292.4]
  wire [13:0] _T_66090; // @[Modules.scala 166:64:@12293.4]
  wire [13:0] buffer_3_498; // @[Modules.scala 166:64:@12294.4]
  wire [14:0] _T_66092; // @[Modules.scala 166:64:@12296.4]
  wire [13:0] _T_66093; // @[Modules.scala 166:64:@12297.4]
  wire [13:0] buffer_3_499; // @[Modules.scala 166:64:@12298.4]
  wire [14:0] _T_66095; // @[Modules.scala 166:64:@12300.4]
  wire [13:0] _T_66096; // @[Modules.scala 166:64:@12301.4]
  wire [13:0] buffer_3_500; // @[Modules.scala 166:64:@12302.4]
  wire [14:0] _T_66098; // @[Modules.scala 166:64:@12304.4]
  wire [13:0] _T_66099; // @[Modules.scala 166:64:@12305.4]
  wire [13:0] buffer_3_501; // @[Modules.scala 166:64:@12306.4]
  wire [14:0] _T_66101; // @[Modules.scala 166:64:@12308.4]
  wire [13:0] _T_66102; // @[Modules.scala 166:64:@12309.4]
  wire [13:0] buffer_3_502; // @[Modules.scala 166:64:@12310.4]
  wire [14:0] _T_66104; // @[Modules.scala 166:64:@12312.4]
  wire [13:0] _T_66105; // @[Modules.scala 166:64:@12313.4]
  wire [13:0] buffer_3_503; // @[Modules.scala 166:64:@12314.4]
  wire [14:0] _T_66107; // @[Modules.scala 166:64:@12316.4]
  wire [13:0] _T_66108; // @[Modules.scala 166:64:@12317.4]
  wire [13:0] buffer_3_504; // @[Modules.scala 166:64:@12318.4]
  wire [14:0] _T_66110; // @[Modules.scala 166:64:@12320.4]
  wire [13:0] _T_66111; // @[Modules.scala 166:64:@12321.4]
  wire [13:0] buffer_3_505; // @[Modules.scala 166:64:@12322.4]
  wire [14:0] _T_66113; // @[Modules.scala 166:64:@12324.4]
  wire [13:0] _T_66114; // @[Modules.scala 166:64:@12325.4]
  wire [13:0] buffer_3_506; // @[Modules.scala 166:64:@12326.4]
  wire [14:0] _T_66116; // @[Modules.scala 166:64:@12328.4]
  wire [13:0] _T_66117; // @[Modules.scala 166:64:@12329.4]
  wire [13:0] buffer_3_507; // @[Modules.scala 166:64:@12330.4]
  wire [14:0] _T_66122; // @[Modules.scala 166:64:@12336.4]
  wire [13:0] _T_66123; // @[Modules.scala 166:64:@12337.4]
  wire [13:0] buffer_3_509; // @[Modules.scala 166:64:@12338.4]
  wire [14:0] _T_66125; // @[Modules.scala 166:64:@12340.4]
  wire [13:0] _T_66126; // @[Modules.scala 166:64:@12341.4]
  wire [13:0] buffer_3_510; // @[Modules.scala 166:64:@12342.4]
  wire [14:0] _T_66128; // @[Modules.scala 166:64:@12344.4]
  wire [13:0] _T_66129; // @[Modules.scala 166:64:@12345.4]
  wire [13:0] buffer_3_511; // @[Modules.scala 166:64:@12346.4]
  wire [14:0] _T_66131; // @[Modules.scala 166:64:@12348.4]
  wire [13:0] _T_66132; // @[Modules.scala 166:64:@12349.4]
  wire [13:0] buffer_3_512; // @[Modules.scala 166:64:@12350.4]
  wire [14:0] _T_66134; // @[Modules.scala 166:64:@12352.4]
  wire [13:0] _T_66135; // @[Modules.scala 166:64:@12353.4]
  wire [13:0] buffer_3_513; // @[Modules.scala 166:64:@12354.4]
  wire [14:0] _T_66137; // @[Modules.scala 166:64:@12356.4]
  wire [13:0] _T_66138; // @[Modules.scala 166:64:@12357.4]
  wire [13:0] buffer_3_514; // @[Modules.scala 166:64:@12358.4]
  wire [14:0] _T_66140; // @[Modules.scala 166:64:@12360.4]
  wire [13:0] _T_66141; // @[Modules.scala 166:64:@12361.4]
  wire [13:0] buffer_3_515; // @[Modules.scala 166:64:@12362.4]
  wire [14:0] _T_66143; // @[Modules.scala 166:64:@12364.4]
  wire [13:0] _T_66144; // @[Modules.scala 166:64:@12365.4]
  wire [13:0] buffer_3_516; // @[Modules.scala 166:64:@12366.4]
  wire [14:0] _T_66146; // @[Modules.scala 166:64:@12368.4]
  wire [13:0] _T_66147; // @[Modules.scala 166:64:@12369.4]
  wire [13:0] buffer_3_517; // @[Modules.scala 166:64:@12370.4]
  wire [14:0] _T_66149; // @[Modules.scala 166:64:@12372.4]
  wire [13:0] _T_66150; // @[Modules.scala 166:64:@12373.4]
  wire [13:0] buffer_3_518; // @[Modules.scala 166:64:@12374.4]
  wire [14:0] _T_66152; // @[Modules.scala 166:64:@12376.4]
  wire [13:0] _T_66153; // @[Modules.scala 166:64:@12377.4]
  wire [13:0] buffer_3_519; // @[Modules.scala 166:64:@12378.4]
  wire [14:0] _T_66155; // @[Modules.scala 166:64:@12380.4]
  wire [13:0] _T_66156; // @[Modules.scala 166:64:@12381.4]
  wire [13:0] buffer_3_520; // @[Modules.scala 166:64:@12382.4]
  wire [14:0] _T_66158; // @[Modules.scala 166:64:@12384.4]
  wire [13:0] _T_66159; // @[Modules.scala 166:64:@12385.4]
  wire [13:0] buffer_3_521; // @[Modules.scala 166:64:@12386.4]
  wire [14:0] _T_66161; // @[Modules.scala 166:64:@12388.4]
  wire [13:0] _T_66162; // @[Modules.scala 166:64:@12389.4]
  wire [13:0] buffer_3_522; // @[Modules.scala 166:64:@12390.4]
  wire [14:0] _T_66164; // @[Modules.scala 166:64:@12392.4]
  wire [13:0] _T_66165; // @[Modules.scala 166:64:@12393.4]
  wire [13:0] buffer_3_523; // @[Modules.scala 166:64:@12394.4]
  wire [14:0] _T_66167; // @[Modules.scala 166:64:@12396.4]
  wire [13:0] _T_66168; // @[Modules.scala 166:64:@12397.4]
  wire [13:0] buffer_3_524; // @[Modules.scala 166:64:@12398.4]
  wire [14:0] _T_66170; // @[Modules.scala 166:64:@12400.4]
  wire [13:0] _T_66171; // @[Modules.scala 166:64:@12401.4]
  wire [13:0] buffer_3_525; // @[Modules.scala 166:64:@12402.4]
  wire [14:0] _T_66173; // @[Modules.scala 166:64:@12404.4]
  wire [13:0] _T_66174; // @[Modules.scala 166:64:@12405.4]
  wire [13:0] buffer_3_526; // @[Modules.scala 166:64:@12406.4]
  wire [14:0] _T_66176; // @[Modules.scala 166:64:@12408.4]
  wire [13:0] _T_66177; // @[Modules.scala 166:64:@12409.4]
  wire [13:0] buffer_3_527; // @[Modules.scala 166:64:@12410.4]
  wire [14:0] _T_66179; // @[Modules.scala 166:64:@12412.4]
  wire [13:0] _T_66180; // @[Modules.scala 166:64:@12413.4]
  wire [13:0] buffer_3_528; // @[Modules.scala 166:64:@12414.4]
  wire [14:0] _T_66182; // @[Modules.scala 166:64:@12416.4]
  wire [13:0] _T_66183; // @[Modules.scala 166:64:@12417.4]
  wire [13:0] buffer_3_529; // @[Modules.scala 166:64:@12418.4]
  wire [14:0] _T_66185; // @[Modules.scala 166:64:@12420.4]
  wire [13:0] _T_66186; // @[Modules.scala 166:64:@12421.4]
  wire [13:0] buffer_3_530; // @[Modules.scala 166:64:@12422.4]
  wire [14:0] _T_66188; // @[Modules.scala 166:64:@12424.4]
  wire [13:0] _T_66189; // @[Modules.scala 166:64:@12425.4]
  wire [13:0] buffer_3_531; // @[Modules.scala 166:64:@12426.4]
  wire [14:0] _T_66191; // @[Modules.scala 166:64:@12428.4]
  wire [13:0] _T_66192; // @[Modules.scala 166:64:@12429.4]
  wire [13:0] buffer_3_532; // @[Modules.scala 166:64:@12430.4]
  wire [14:0] _T_66194; // @[Modules.scala 166:64:@12432.4]
  wire [13:0] _T_66195; // @[Modules.scala 166:64:@12433.4]
  wire [13:0] buffer_3_533; // @[Modules.scala 166:64:@12434.4]
  wire [14:0] _T_66197; // @[Modules.scala 166:64:@12436.4]
  wire [13:0] _T_66198; // @[Modules.scala 166:64:@12437.4]
  wire [13:0] buffer_3_534; // @[Modules.scala 166:64:@12438.4]
  wire [14:0] _T_66200; // @[Modules.scala 166:64:@12440.4]
  wire [13:0] _T_66201; // @[Modules.scala 166:64:@12441.4]
  wire [13:0] buffer_3_535; // @[Modules.scala 166:64:@12442.4]
  wire [14:0] _T_66203; // @[Modules.scala 166:64:@12444.4]
  wire [13:0] _T_66204; // @[Modules.scala 166:64:@12445.4]
  wire [13:0] buffer_3_536; // @[Modules.scala 166:64:@12446.4]
  wire [14:0] _T_66206; // @[Modules.scala 166:64:@12448.4]
  wire [13:0] _T_66207; // @[Modules.scala 166:64:@12449.4]
  wire [13:0] buffer_3_537; // @[Modules.scala 166:64:@12450.4]
  wire [14:0] _T_66209; // @[Modules.scala 166:64:@12452.4]
  wire [13:0] _T_66210; // @[Modules.scala 166:64:@12453.4]
  wire [13:0] buffer_3_538; // @[Modules.scala 166:64:@12454.4]
  wire [14:0] _T_66212; // @[Modules.scala 166:64:@12456.4]
  wire [13:0] _T_66213; // @[Modules.scala 166:64:@12457.4]
  wire [13:0] buffer_3_539; // @[Modules.scala 166:64:@12458.4]
  wire [14:0] _T_66215; // @[Modules.scala 166:64:@12460.4]
  wire [13:0] _T_66216; // @[Modules.scala 166:64:@12461.4]
  wire [13:0] buffer_3_540; // @[Modules.scala 166:64:@12462.4]
  wire [14:0] _T_66218; // @[Modules.scala 166:64:@12464.4]
  wire [13:0] _T_66219; // @[Modules.scala 166:64:@12465.4]
  wire [13:0] buffer_3_541; // @[Modules.scala 166:64:@12466.4]
  wire [14:0] _T_66221; // @[Modules.scala 166:64:@12468.4]
  wire [13:0] _T_66222; // @[Modules.scala 166:64:@12469.4]
  wire [13:0] buffer_3_542; // @[Modules.scala 166:64:@12470.4]
  wire [14:0] _T_66224; // @[Modules.scala 166:64:@12472.4]
  wire [13:0] _T_66225; // @[Modules.scala 166:64:@12473.4]
  wire [13:0] buffer_3_543; // @[Modules.scala 166:64:@12474.4]
  wire [14:0] _T_66227; // @[Modules.scala 166:64:@12476.4]
  wire [13:0] _T_66228; // @[Modules.scala 166:64:@12477.4]
  wire [13:0] buffer_3_544; // @[Modules.scala 166:64:@12478.4]
  wire [14:0] _T_66230; // @[Modules.scala 166:64:@12480.4]
  wire [13:0] _T_66231; // @[Modules.scala 166:64:@12481.4]
  wire [13:0] buffer_3_545; // @[Modules.scala 166:64:@12482.4]
  wire [14:0] _T_66233; // @[Modules.scala 166:64:@12484.4]
  wire [13:0] _T_66234; // @[Modules.scala 166:64:@12485.4]
  wire [13:0] buffer_3_546; // @[Modules.scala 166:64:@12486.4]
  wire [14:0] _T_66236; // @[Modules.scala 166:64:@12488.4]
  wire [13:0] _T_66237; // @[Modules.scala 166:64:@12489.4]
  wire [13:0] buffer_3_547; // @[Modules.scala 166:64:@12490.4]
  wire [14:0] _T_66239; // @[Modules.scala 166:64:@12492.4]
  wire [13:0] _T_66240; // @[Modules.scala 166:64:@12493.4]
  wire [13:0] buffer_3_548; // @[Modules.scala 166:64:@12494.4]
  wire [14:0] _T_66242; // @[Modules.scala 160:64:@12496.4]
  wire [13:0] _T_66243; // @[Modules.scala 160:64:@12497.4]
  wire [13:0] buffer_3_549; // @[Modules.scala 160:64:@12498.4]
  wire [14:0] _T_66245; // @[Modules.scala 160:64:@12500.4]
  wire [13:0] _T_66246; // @[Modules.scala 160:64:@12501.4]
  wire [13:0] buffer_3_550; // @[Modules.scala 160:64:@12502.4]
  wire [14:0] _T_66248; // @[Modules.scala 160:64:@12504.4]
  wire [13:0] _T_66249; // @[Modules.scala 160:64:@12505.4]
  wire [13:0] buffer_3_551; // @[Modules.scala 160:64:@12506.4]
  wire [14:0] _T_66251; // @[Modules.scala 160:64:@12508.4]
  wire [13:0] _T_66252; // @[Modules.scala 160:64:@12509.4]
  wire [13:0] buffer_3_552; // @[Modules.scala 160:64:@12510.4]
  wire [14:0] _T_66254; // @[Modules.scala 160:64:@12512.4]
  wire [13:0] _T_66255; // @[Modules.scala 160:64:@12513.4]
  wire [13:0] buffer_3_553; // @[Modules.scala 160:64:@12514.4]
  wire [14:0] _T_66257; // @[Modules.scala 160:64:@12516.4]
  wire [13:0] _T_66258; // @[Modules.scala 160:64:@12517.4]
  wire [13:0] buffer_3_554; // @[Modules.scala 160:64:@12518.4]
  wire [14:0] _T_66260; // @[Modules.scala 160:64:@12520.4]
  wire [13:0] _T_66261; // @[Modules.scala 160:64:@12521.4]
  wire [13:0] buffer_3_555; // @[Modules.scala 160:64:@12522.4]
  wire [14:0] _T_66263; // @[Modules.scala 160:64:@12524.4]
  wire [13:0] _T_66264; // @[Modules.scala 160:64:@12525.4]
  wire [13:0] buffer_3_556; // @[Modules.scala 160:64:@12526.4]
  wire [14:0] _T_66266; // @[Modules.scala 160:64:@12528.4]
  wire [13:0] _T_66267; // @[Modules.scala 160:64:@12529.4]
  wire [13:0] buffer_3_557; // @[Modules.scala 160:64:@12530.4]
  wire [14:0] _T_66269; // @[Modules.scala 160:64:@12532.4]
  wire [13:0] _T_66270; // @[Modules.scala 160:64:@12533.4]
  wire [13:0] buffer_3_558; // @[Modules.scala 160:64:@12534.4]
  wire [14:0] _T_66272; // @[Modules.scala 160:64:@12536.4]
  wire [13:0] _T_66273; // @[Modules.scala 160:64:@12537.4]
  wire [13:0] buffer_3_559; // @[Modules.scala 160:64:@12538.4]
  wire [14:0] _T_66275; // @[Modules.scala 160:64:@12540.4]
  wire [13:0] _T_66276; // @[Modules.scala 160:64:@12541.4]
  wire [13:0] buffer_3_560; // @[Modules.scala 160:64:@12542.4]
  wire [14:0] _T_66278; // @[Modules.scala 160:64:@12544.4]
  wire [13:0] _T_66279; // @[Modules.scala 160:64:@12545.4]
  wire [13:0] buffer_3_561; // @[Modules.scala 160:64:@12546.4]
  wire [14:0] _T_66281; // @[Modules.scala 160:64:@12548.4]
  wire [13:0] _T_66282; // @[Modules.scala 160:64:@12549.4]
  wire [13:0] buffer_3_562; // @[Modules.scala 160:64:@12550.4]
  wire [14:0] _T_66284; // @[Modules.scala 160:64:@12552.4]
  wire [13:0] _T_66285; // @[Modules.scala 160:64:@12553.4]
  wire [13:0] buffer_3_563; // @[Modules.scala 160:64:@12554.4]
  wire [14:0] _T_66287; // @[Modules.scala 160:64:@12556.4]
  wire [13:0] _T_66288; // @[Modules.scala 160:64:@12557.4]
  wire [13:0] buffer_3_564; // @[Modules.scala 160:64:@12558.4]
  wire [14:0] _T_66290; // @[Modules.scala 160:64:@12560.4]
  wire [13:0] _T_66291; // @[Modules.scala 160:64:@12561.4]
  wire [13:0] buffer_3_565; // @[Modules.scala 160:64:@12562.4]
  wire [14:0] _T_66293; // @[Modules.scala 160:64:@12564.4]
  wire [13:0] _T_66294; // @[Modules.scala 160:64:@12565.4]
  wire [13:0] buffer_3_566; // @[Modules.scala 160:64:@12566.4]
  wire [14:0] _T_66296; // @[Modules.scala 160:64:@12568.4]
  wire [13:0] _T_66297; // @[Modules.scala 160:64:@12569.4]
  wire [13:0] buffer_3_567; // @[Modules.scala 160:64:@12570.4]
  wire [14:0] _T_66299; // @[Modules.scala 160:64:@12572.4]
  wire [13:0] _T_66300; // @[Modules.scala 160:64:@12573.4]
  wire [13:0] buffer_3_568; // @[Modules.scala 160:64:@12574.4]
  wire [14:0] _T_66302; // @[Modules.scala 160:64:@12576.4]
  wire [13:0] _T_66303; // @[Modules.scala 160:64:@12577.4]
  wire [13:0] buffer_3_569; // @[Modules.scala 160:64:@12578.4]
  wire [14:0] _T_66305; // @[Modules.scala 160:64:@12580.4]
  wire [13:0] _T_66306; // @[Modules.scala 160:64:@12581.4]
  wire [13:0] buffer_3_570; // @[Modules.scala 160:64:@12582.4]
  wire [14:0] _T_66308; // @[Modules.scala 160:64:@12584.4]
  wire [13:0] _T_66309; // @[Modules.scala 160:64:@12585.4]
  wire [13:0] buffer_3_571; // @[Modules.scala 160:64:@12586.4]
  wire [14:0] _T_66311; // @[Modules.scala 160:64:@12588.4]
  wire [13:0] _T_66312; // @[Modules.scala 160:64:@12589.4]
  wire [13:0] buffer_3_572; // @[Modules.scala 160:64:@12590.4]
  wire [14:0] _T_66314; // @[Modules.scala 160:64:@12592.4]
  wire [13:0] _T_66315; // @[Modules.scala 160:64:@12593.4]
  wire [13:0] buffer_3_573; // @[Modules.scala 160:64:@12594.4]
  wire [14:0] _T_66317; // @[Modules.scala 160:64:@12596.4]
  wire [13:0] _T_66318; // @[Modules.scala 160:64:@12597.4]
  wire [13:0] buffer_3_574; // @[Modules.scala 160:64:@12598.4]
  wire [14:0] _T_66320; // @[Modules.scala 160:64:@12600.4]
  wire [13:0] _T_66321; // @[Modules.scala 160:64:@12601.4]
  wire [13:0] buffer_3_575; // @[Modules.scala 160:64:@12602.4]
  wire [14:0] _T_66323; // @[Modules.scala 160:64:@12604.4]
  wire [13:0] _T_66324; // @[Modules.scala 160:64:@12605.4]
  wire [13:0] buffer_3_576; // @[Modules.scala 160:64:@12606.4]
  wire [14:0] _T_66326; // @[Modules.scala 160:64:@12608.4]
  wire [13:0] _T_66327; // @[Modules.scala 160:64:@12609.4]
  wire [13:0] buffer_3_577; // @[Modules.scala 160:64:@12610.4]
  wire [14:0] _T_66329; // @[Modules.scala 160:64:@12612.4]
  wire [13:0] _T_66330; // @[Modules.scala 160:64:@12613.4]
  wire [13:0] buffer_3_578; // @[Modules.scala 160:64:@12614.4]
  wire [14:0] _T_66332; // @[Modules.scala 160:64:@12616.4]
  wire [13:0] _T_66333; // @[Modules.scala 160:64:@12617.4]
  wire [13:0] buffer_3_579; // @[Modules.scala 160:64:@12618.4]
  wire [14:0] _T_66335; // @[Modules.scala 160:64:@12620.4]
  wire [13:0] _T_66336; // @[Modules.scala 160:64:@12621.4]
  wire [13:0] buffer_3_580; // @[Modules.scala 160:64:@12622.4]
  wire [14:0] _T_66338; // @[Modules.scala 160:64:@12624.4]
  wire [13:0] _T_66339; // @[Modules.scala 160:64:@12625.4]
  wire [13:0] buffer_3_581; // @[Modules.scala 160:64:@12626.4]
  wire [14:0] _T_66341; // @[Modules.scala 160:64:@12628.4]
  wire [13:0] _T_66342; // @[Modules.scala 160:64:@12629.4]
  wire [13:0] buffer_3_582; // @[Modules.scala 160:64:@12630.4]
  wire [14:0] _T_66344; // @[Modules.scala 160:64:@12632.4]
  wire [13:0] _T_66345; // @[Modules.scala 160:64:@12633.4]
  wire [13:0] buffer_3_583; // @[Modules.scala 160:64:@12634.4]
  wire [14:0] _T_66347; // @[Modules.scala 160:64:@12636.4]
  wire [13:0] _T_66348; // @[Modules.scala 160:64:@12637.4]
  wire [13:0] buffer_3_584; // @[Modules.scala 160:64:@12638.4]
  wire [14:0] _T_66350; // @[Modules.scala 160:64:@12640.4]
  wire [13:0] _T_66351; // @[Modules.scala 160:64:@12641.4]
  wire [13:0] buffer_3_585; // @[Modules.scala 160:64:@12642.4]
  wire [14:0] _T_66353; // @[Modules.scala 160:64:@12644.4]
  wire [13:0] _T_66354; // @[Modules.scala 160:64:@12645.4]
  wire [13:0] buffer_3_586; // @[Modules.scala 160:64:@12646.4]
  wire [14:0] _T_66356; // @[Modules.scala 160:64:@12648.4]
  wire [13:0] _T_66357; // @[Modules.scala 160:64:@12649.4]
  wire [13:0] buffer_3_587; // @[Modules.scala 160:64:@12650.4]
  wire [14:0] _T_66359; // @[Modules.scala 166:64:@12652.4]
  wire [13:0] _T_66360; // @[Modules.scala 166:64:@12653.4]
  wire [13:0] buffer_3_588; // @[Modules.scala 166:64:@12654.4]
  wire [14:0] _T_66362; // @[Modules.scala 166:64:@12656.4]
  wire [13:0] _T_66363; // @[Modules.scala 166:64:@12657.4]
  wire [13:0] buffer_3_589; // @[Modules.scala 166:64:@12658.4]
  wire [14:0] _T_66365; // @[Modules.scala 166:64:@12660.4]
  wire [13:0] _T_66366; // @[Modules.scala 166:64:@12661.4]
  wire [13:0] buffer_3_590; // @[Modules.scala 166:64:@12662.4]
  wire [14:0] _T_66368; // @[Modules.scala 166:64:@12664.4]
  wire [13:0] _T_66369; // @[Modules.scala 166:64:@12665.4]
  wire [13:0] buffer_3_591; // @[Modules.scala 166:64:@12666.4]
  wire [14:0] _T_66371; // @[Modules.scala 166:64:@12668.4]
  wire [13:0] _T_66372; // @[Modules.scala 166:64:@12669.4]
  wire [13:0] buffer_3_592; // @[Modules.scala 166:64:@12670.4]
  wire [14:0] _T_66374; // @[Modules.scala 166:64:@12672.4]
  wire [13:0] _T_66375; // @[Modules.scala 166:64:@12673.4]
  wire [13:0] buffer_3_593; // @[Modules.scala 166:64:@12674.4]
  wire [14:0] _T_66377; // @[Modules.scala 166:64:@12676.4]
  wire [13:0] _T_66378; // @[Modules.scala 166:64:@12677.4]
  wire [13:0] buffer_3_594; // @[Modules.scala 166:64:@12678.4]
  wire [14:0] _T_66380; // @[Modules.scala 166:64:@12680.4]
  wire [13:0] _T_66381; // @[Modules.scala 166:64:@12681.4]
  wire [13:0] buffer_3_595; // @[Modules.scala 166:64:@12682.4]
  wire [14:0] _T_66383; // @[Modules.scala 166:64:@12684.4]
  wire [13:0] _T_66384; // @[Modules.scala 166:64:@12685.4]
  wire [13:0] buffer_3_596; // @[Modules.scala 166:64:@12686.4]
  wire [14:0] _T_66386; // @[Modules.scala 166:64:@12688.4]
  wire [13:0] _T_66387; // @[Modules.scala 166:64:@12689.4]
  wire [13:0] buffer_3_597; // @[Modules.scala 166:64:@12690.4]
  wire [14:0] _T_66389; // @[Modules.scala 166:64:@12692.4]
  wire [13:0] _T_66390; // @[Modules.scala 166:64:@12693.4]
  wire [13:0] buffer_3_598; // @[Modules.scala 166:64:@12694.4]
  wire [14:0] _T_66392; // @[Modules.scala 166:64:@12696.4]
  wire [13:0] _T_66393; // @[Modules.scala 166:64:@12697.4]
  wire [13:0] buffer_3_599; // @[Modules.scala 166:64:@12698.4]
  wire [14:0] _T_66395; // @[Modules.scala 166:64:@12700.4]
  wire [13:0] _T_66396; // @[Modules.scala 166:64:@12701.4]
  wire [13:0] buffer_3_600; // @[Modules.scala 166:64:@12702.4]
  wire [14:0] _T_66398; // @[Modules.scala 166:64:@12704.4]
  wire [13:0] _T_66399; // @[Modules.scala 166:64:@12705.4]
  wire [13:0] buffer_3_601; // @[Modules.scala 166:64:@12706.4]
  wire [14:0] _T_66401; // @[Modules.scala 166:64:@12708.4]
  wire [13:0] _T_66402; // @[Modules.scala 166:64:@12709.4]
  wire [13:0] buffer_3_602; // @[Modules.scala 166:64:@12710.4]
  wire [14:0] _T_66404; // @[Modules.scala 166:64:@12712.4]
  wire [13:0] _T_66405; // @[Modules.scala 166:64:@12713.4]
  wire [13:0] buffer_3_603; // @[Modules.scala 166:64:@12714.4]
  wire [14:0] _T_66407; // @[Modules.scala 166:64:@12716.4]
  wire [13:0] _T_66408; // @[Modules.scala 166:64:@12717.4]
  wire [13:0] buffer_3_604; // @[Modules.scala 166:64:@12718.4]
  wire [14:0] _T_66410; // @[Modules.scala 166:64:@12720.4]
  wire [13:0] _T_66411; // @[Modules.scala 166:64:@12721.4]
  wire [13:0] buffer_3_605; // @[Modules.scala 166:64:@12722.4]
  wire [14:0] _T_66413; // @[Modules.scala 166:64:@12724.4]
  wire [13:0] _T_66414; // @[Modules.scala 166:64:@12725.4]
  wire [13:0] buffer_3_606; // @[Modules.scala 166:64:@12726.4]
  wire [14:0] _T_66416; // @[Modules.scala 172:66:@12728.4]
  wire [13:0] _T_66417; // @[Modules.scala 172:66:@12729.4]
  wire [13:0] buffer_3_607; // @[Modules.scala 172:66:@12730.4]
  wire [14:0] _T_66419; // @[Modules.scala 160:64:@12732.4]
  wire [13:0] _T_66420; // @[Modules.scala 160:64:@12733.4]
  wire [13:0] buffer_3_608; // @[Modules.scala 160:64:@12734.4]
  wire [14:0] _T_66422; // @[Modules.scala 160:64:@12736.4]
  wire [13:0] _T_66423; // @[Modules.scala 160:64:@12737.4]
  wire [13:0] buffer_3_609; // @[Modules.scala 160:64:@12738.4]
  wire [14:0] _T_66425; // @[Modules.scala 160:64:@12740.4]
  wire [13:0] _T_66426; // @[Modules.scala 160:64:@12741.4]
  wire [13:0] buffer_3_610; // @[Modules.scala 160:64:@12742.4]
  wire [14:0] _T_66428; // @[Modules.scala 160:64:@12744.4]
  wire [13:0] _T_66429; // @[Modules.scala 160:64:@12745.4]
  wire [13:0] buffer_3_611; // @[Modules.scala 160:64:@12746.4]
  wire [14:0] _T_66431; // @[Modules.scala 160:64:@12748.4]
  wire [13:0] _T_66432; // @[Modules.scala 160:64:@12749.4]
  wire [13:0] buffer_3_612; // @[Modules.scala 160:64:@12750.4]
  wire [14:0] _T_66434; // @[Modules.scala 160:64:@12752.4]
  wire [13:0] _T_66435; // @[Modules.scala 160:64:@12753.4]
  wire [13:0] buffer_3_613; // @[Modules.scala 160:64:@12754.4]
  wire [14:0] _T_66437; // @[Modules.scala 160:64:@12756.4]
  wire [13:0] _T_66438; // @[Modules.scala 160:64:@12757.4]
  wire [13:0] buffer_3_614; // @[Modules.scala 160:64:@12758.4]
  wire [14:0] _T_66440; // @[Modules.scala 160:64:@12760.4]
  wire [13:0] _T_66441; // @[Modules.scala 160:64:@12761.4]
  wire [13:0] buffer_3_615; // @[Modules.scala 160:64:@12762.4]
  wire [14:0] _T_66443; // @[Modules.scala 160:64:@12764.4]
  wire [13:0] _T_66444; // @[Modules.scala 160:64:@12765.4]
  wire [13:0] buffer_3_616; // @[Modules.scala 160:64:@12766.4]
  wire [14:0] _T_66446; // @[Modules.scala 160:64:@12768.4]
  wire [13:0] _T_66447; // @[Modules.scala 160:64:@12769.4]
  wire [13:0] buffer_3_617; // @[Modules.scala 160:64:@12770.4]
  wire [14:0] _T_66449; // @[Modules.scala 160:64:@12772.4]
  wire [13:0] _T_66450; // @[Modules.scala 160:64:@12773.4]
  wire [13:0] buffer_3_618; // @[Modules.scala 160:64:@12774.4]
  wire [14:0] _T_66452; // @[Modules.scala 160:64:@12776.4]
  wire [13:0] _T_66453; // @[Modules.scala 160:64:@12777.4]
  wire [13:0] buffer_3_619; // @[Modules.scala 160:64:@12778.4]
  wire [14:0] _T_66455; // @[Modules.scala 160:64:@12780.4]
  wire [13:0] _T_66456; // @[Modules.scala 160:64:@12781.4]
  wire [13:0] buffer_3_620; // @[Modules.scala 160:64:@12782.4]
  wire [14:0] _T_66458; // @[Modules.scala 160:64:@12784.4]
  wire [13:0] _T_66459; // @[Modules.scala 160:64:@12785.4]
  wire [13:0] buffer_3_621; // @[Modules.scala 160:64:@12786.4]
  wire [14:0] _T_66461; // @[Modules.scala 160:64:@12788.4]
  wire [13:0] _T_66462; // @[Modules.scala 160:64:@12789.4]
  wire [13:0] buffer_3_622; // @[Modules.scala 160:64:@12790.4]
  wire [14:0] _T_66464; // @[Modules.scala 166:64:@12792.4]
  wire [13:0] _T_66465; // @[Modules.scala 166:64:@12793.4]
  wire [13:0] buffer_3_623; // @[Modules.scala 166:64:@12794.4]
  wire [14:0] _T_66467; // @[Modules.scala 166:64:@12796.4]
  wire [13:0] _T_66468; // @[Modules.scala 166:64:@12797.4]
  wire [13:0] buffer_3_624; // @[Modules.scala 166:64:@12798.4]
  wire [14:0] _T_66470; // @[Modules.scala 160:64:@12800.4]
  wire [13:0] _T_66471; // @[Modules.scala 160:64:@12801.4]
  wire [13:0] buffer_3_625; // @[Modules.scala 160:64:@12802.4]
  wire [14:0] _T_66473; // @[Modules.scala 172:66:@12804.4]
  wire [13:0] _T_66474; // @[Modules.scala 172:66:@12805.4]
  wire [13:0] buffer_3_626; // @[Modules.scala 172:66:@12806.4]
  wire [5:0] _T_66491; // @[Modules.scala 150:74:@12977.4]
  wire [5:0] _GEN_279; // @[Modules.scala 150:103:@12979.4]
  wire [6:0] _T_66494; // @[Modules.scala 150:103:@12979.4]
  wire [5:0] _T_66495; // @[Modules.scala 150:103:@12980.4]
  wire [5:0] _T_66496; // @[Modules.scala 150:103:@12981.4]
  wire [4:0] _T_66500; // @[Modules.scala 151:80:@12984.4]
  wire [5:0] _T_66501; // @[Modules.scala 150:103:@12985.4]
  wire [4:0] _T_66502; // @[Modules.scala 150:103:@12986.4]
  wire [4:0] _T_66503; // @[Modules.scala 150:103:@12987.4]
  wire [5:0] _T_66508; // @[Modules.scala 150:103:@12991.4]
  wire [4:0] _T_66509; // @[Modules.scala 150:103:@12992.4]
  wire [4:0] _T_66510; // @[Modules.scala 150:103:@12993.4]
  wire [6:0] _T_66522; // @[Modules.scala 150:103:@13003.4]
  wire [5:0] _T_66523; // @[Modules.scala 150:103:@13004.4]
  wire [5:0] _T_66524; // @[Modules.scala 150:103:@13005.4]
  wire [6:0] _T_66529; // @[Modules.scala 150:103:@13009.4]
  wire [5:0] _T_66530; // @[Modules.scala 150:103:@13010.4]
  wire [5:0] _T_66531; // @[Modules.scala 150:103:@13011.4]
  wire [5:0] _T_66543; // @[Modules.scala 150:103:@13021.4]
  wire [4:0] _T_66544; // @[Modules.scala 150:103:@13022.4]
  wire [4:0] _T_66545; // @[Modules.scala 150:103:@13023.4]
  wire [5:0] _GEN_281; // @[Modules.scala 150:103:@13027.4]
  wire [6:0] _T_66550; // @[Modules.scala 150:103:@13027.4]
  wire [5:0] _T_66551; // @[Modules.scala 150:103:@13028.4]
  wire [5:0] _T_66552; // @[Modules.scala 150:103:@13029.4]
  wire [5:0] _T_66564; // @[Modules.scala 150:103:@13039.4]
  wire [4:0] _T_66565; // @[Modules.scala 150:103:@13040.4]
  wire [4:0] _T_66566; // @[Modules.scala 150:103:@13041.4]
  wire [5:0] _T_66571; // @[Modules.scala 150:103:@13045.4]
  wire [4:0] _T_66572; // @[Modules.scala 150:103:@13046.4]
  wire [4:0] _T_66573; // @[Modules.scala 150:103:@13047.4]
  wire [4:0] _T_66603; // @[Modules.scala 150:74:@13073.4]
  wire [4:0] _T_66605; // @[Modules.scala 151:80:@13074.4]
  wire [5:0] _T_66606; // @[Modules.scala 150:103:@13075.4]
  wire [4:0] _T_66607; // @[Modules.scala 150:103:@13076.4]
  wire [4:0] _T_66608; // @[Modules.scala 150:103:@13077.4]
  wire [4:0] _T_66610; // @[Modules.scala 150:74:@13079.4]
  wire [5:0] _GEN_282; // @[Modules.scala 150:103:@13081.4]
  wire [6:0] _T_66613; // @[Modules.scala 150:103:@13081.4]
  wire [5:0] _T_66614; // @[Modules.scala 150:103:@13082.4]
  wire [5:0] _T_66615; // @[Modules.scala 150:103:@13083.4]
  wire [5:0] _T_66624; // @[Modules.scala 150:74:@13091.4]
  wire [5:0] _GEN_283; // @[Modules.scala 150:103:@13093.4]
  wire [6:0] _T_66627; // @[Modules.scala 150:103:@13093.4]
  wire [5:0] _T_66628; // @[Modules.scala 150:103:@13094.4]
  wire [5:0] _T_66629; // @[Modules.scala 150:103:@13095.4]
  wire [5:0] _GEN_284; // @[Modules.scala 150:103:@13147.4]
  wire [6:0] _T_66690; // @[Modules.scala 150:103:@13147.4]
  wire [5:0] _T_66691; // @[Modules.scala 150:103:@13148.4]
  wire [5:0] _T_66692; // @[Modules.scala 150:103:@13149.4]
  wire [6:0] _T_66697; // @[Modules.scala 150:103:@13153.4]
  wire [5:0] _T_66698; // @[Modules.scala 150:103:@13154.4]
  wire [5:0] _T_66699; // @[Modules.scala 150:103:@13155.4]
  wire [6:0] _T_66711; // @[Modules.scala 150:103:@13165.4]
  wire [5:0] _T_66712; // @[Modules.scala 150:103:@13166.4]
  wire [5:0] _T_66713; // @[Modules.scala 150:103:@13167.4]
  wire [6:0] _T_66718; // @[Modules.scala 150:103:@13171.4]
  wire [5:0] _T_66719; // @[Modules.scala 150:103:@13172.4]
  wire [5:0] _T_66720; // @[Modules.scala 150:103:@13173.4]
  wire [5:0] _T_66725; // @[Modules.scala 150:103:@13177.4]
  wire [4:0] _T_66726; // @[Modules.scala 150:103:@13178.4]
  wire [4:0] _T_66727; // @[Modules.scala 150:103:@13179.4]
  wire [5:0] _T_66732; // @[Modules.scala 150:103:@13183.4]
  wire [4:0] _T_66733; // @[Modules.scala 150:103:@13184.4]
  wire [4:0] _T_66734; // @[Modules.scala 150:103:@13185.4]
  wire [5:0] _T_66739; // @[Modules.scala 150:103:@13189.4]
  wire [4:0] _T_66740; // @[Modules.scala 150:103:@13190.4]
  wire [4:0] _T_66741; // @[Modules.scala 150:103:@13191.4]
  wire [4:0] _T_66750; // @[Modules.scala 150:74:@13199.4]
  wire [5:0] _GEN_287; // @[Modules.scala 150:103:@13201.4]
  wire [6:0] _T_66753; // @[Modules.scala 150:103:@13201.4]
  wire [5:0] _T_66754; // @[Modules.scala 150:103:@13202.4]
  wire [5:0] _T_66755; // @[Modules.scala 150:103:@13203.4]
  wire [5:0] _GEN_288; // @[Modules.scala 150:103:@13213.4]
  wire [6:0] _T_66767; // @[Modules.scala 150:103:@13213.4]
  wire [5:0] _T_66768; // @[Modules.scala 150:103:@13214.4]
  wire [5:0] _T_66769; // @[Modules.scala 150:103:@13215.4]
  wire [5:0] _T_66774; // @[Modules.scala 150:103:@13219.4]
  wire [4:0] _T_66775; // @[Modules.scala 150:103:@13220.4]
  wire [4:0] _T_66776; // @[Modules.scala 150:103:@13221.4]
  wire [6:0] _T_66781; // @[Modules.scala 150:103:@13225.4]
  wire [5:0] _T_66782; // @[Modules.scala 150:103:@13226.4]
  wire [5:0] _T_66783; // @[Modules.scala 150:103:@13227.4]
  wire [5:0] _GEN_290; // @[Modules.scala 150:103:@13231.4]
  wire [6:0] _T_66788; // @[Modules.scala 150:103:@13231.4]
  wire [5:0] _T_66789; // @[Modules.scala 150:103:@13232.4]
  wire [5:0] _T_66790; // @[Modules.scala 150:103:@13233.4]
  wire [5:0] _T_66823; // @[Modules.scala 150:103:@13261.4]
  wire [4:0] _T_66824; // @[Modules.scala 150:103:@13262.4]
  wire [4:0] _T_66825; // @[Modules.scala 150:103:@13263.4]
  wire [4:0] _T_66841; // @[Modules.scala 150:74:@13277.4]
  wire [5:0] _T_66844; // @[Modules.scala 150:103:@13279.4]
  wire [4:0] _T_66845; // @[Modules.scala 150:103:@13280.4]
  wire [4:0] _T_66846; // @[Modules.scala 150:103:@13281.4]
  wire [5:0] _T_66851; // @[Modules.scala 150:103:@13285.4]
  wire [4:0] _T_66852; // @[Modules.scala 150:103:@13286.4]
  wire [4:0] _T_66853; // @[Modules.scala 150:103:@13287.4]
  wire [5:0] _T_66865; // @[Modules.scala 150:103:@13297.4]
  wire [4:0] _T_66866; // @[Modules.scala 150:103:@13298.4]
  wire [4:0] _T_66867; // @[Modules.scala 150:103:@13299.4]
  wire [6:0] _T_66872; // @[Modules.scala 150:103:@13303.4]
  wire [5:0] _T_66873; // @[Modules.scala 150:103:@13304.4]
  wire [5:0] _T_66874; // @[Modules.scala 150:103:@13305.4]
  wire [6:0] _T_66879; // @[Modules.scala 150:103:@13309.4]
  wire [5:0] _T_66880; // @[Modules.scala 150:103:@13310.4]
  wire [5:0] _T_66881; // @[Modules.scala 150:103:@13311.4]
  wire [5:0] _T_66907; // @[Modules.scala 150:103:@13333.4]
  wire [4:0] _T_66908; // @[Modules.scala 150:103:@13334.4]
  wire [4:0] _T_66909; // @[Modules.scala 150:103:@13335.4]
  wire [6:0] _T_66914; // @[Modules.scala 150:103:@13339.4]
  wire [5:0] _T_66915; // @[Modules.scala 150:103:@13340.4]
  wire [5:0] _T_66916; // @[Modules.scala 150:103:@13341.4]
  wire [5:0] _T_66920; // @[Modules.scala 151:80:@13344.4]
  wire [6:0] _T_66921; // @[Modules.scala 150:103:@13345.4]
  wire [5:0] _T_66922; // @[Modules.scala 150:103:@13346.4]
  wire [5:0] _T_66923; // @[Modules.scala 150:103:@13347.4]
  wire [5:0] _T_66925; // @[Modules.scala 150:74:@13349.4]
  wire [5:0] _GEN_293; // @[Modules.scala 150:103:@13351.4]
  wire [6:0] _T_66928; // @[Modules.scala 150:103:@13351.4]
  wire [5:0] _T_66929; // @[Modules.scala 150:103:@13352.4]
  wire [5:0] _T_66930; // @[Modules.scala 150:103:@13353.4]
  wire [5:0] _T_66977; // @[Modules.scala 150:103:@13393.4]
  wire [4:0] _T_66978; // @[Modules.scala 150:103:@13394.4]
  wire [4:0] _T_66979; // @[Modules.scala 150:103:@13395.4]
  wire [6:0] _T_66984; // @[Modules.scala 150:103:@13399.4]
  wire [5:0] _T_66985; // @[Modules.scala 150:103:@13400.4]
  wire [5:0] _T_66986; // @[Modules.scala 150:103:@13401.4]
  wire [6:0] _T_66991; // @[Modules.scala 150:103:@13405.4]
  wire [5:0] _T_66992; // @[Modules.scala 150:103:@13406.4]
  wire [5:0] _T_66993; // @[Modules.scala 150:103:@13407.4]
  wire [5:0] _GEN_295; // @[Modules.scala 150:103:@13417.4]
  wire [6:0] _T_67005; // @[Modules.scala 150:103:@13417.4]
  wire [5:0] _T_67006; // @[Modules.scala 150:103:@13418.4]
  wire [5:0] _T_67007; // @[Modules.scala 150:103:@13419.4]
  wire [5:0] _GEN_296; // @[Modules.scala 150:103:@13435.4]
  wire [6:0] _T_67026; // @[Modules.scala 150:103:@13435.4]
  wire [5:0] _T_67027; // @[Modules.scala 150:103:@13436.4]
  wire [5:0] _T_67028; // @[Modules.scala 150:103:@13437.4]
  wire [6:0] _T_67033; // @[Modules.scala 150:103:@13441.4]
  wire [5:0] _T_67034; // @[Modules.scala 150:103:@13442.4]
  wire [5:0] _T_67035; // @[Modules.scala 150:103:@13443.4]
  wire [5:0] _GEN_297; // @[Modules.scala 150:103:@13447.4]
  wire [6:0] _T_67040; // @[Modules.scala 150:103:@13447.4]
  wire [5:0] _T_67041; // @[Modules.scala 150:103:@13448.4]
  wire [5:0] _T_67042; // @[Modules.scala 150:103:@13449.4]
  wire [5:0] _T_67053; // @[Modules.scala 151:80:@13458.4]
  wire [5:0] _GEN_298; // @[Modules.scala 150:103:@13459.4]
  wire [6:0] _T_67054; // @[Modules.scala 150:103:@13459.4]
  wire [5:0] _T_67055; // @[Modules.scala 150:103:@13460.4]
  wire [5:0] _T_67056; // @[Modules.scala 150:103:@13461.4]
  wire [5:0] _GEN_299; // @[Modules.scala 150:103:@13477.4]
  wire [6:0] _T_67075; // @[Modules.scala 150:103:@13477.4]
  wire [5:0] _T_67076; // @[Modules.scala 150:103:@13478.4]
  wire [5:0] _T_67077; // @[Modules.scala 150:103:@13479.4]
  wire [6:0] _T_67110; // @[Modules.scala 150:103:@13507.4]
  wire [5:0] _T_67111; // @[Modules.scala 150:103:@13508.4]
  wire [5:0] _T_67112; // @[Modules.scala 150:103:@13509.4]
  wire [5:0] _GEN_300; // @[Modules.scala 150:103:@13513.4]
  wire [6:0] _T_67117; // @[Modules.scala 150:103:@13513.4]
  wire [5:0] _T_67118; // @[Modules.scala 150:103:@13514.4]
  wire [5:0] _T_67119; // @[Modules.scala 150:103:@13515.4]
  wire [5:0] _T_67124; // @[Modules.scala 150:103:@13519.4]
  wire [4:0] _T_67125; // @[Modules.scala 150:103:@13520.4]
  wire [4:0] _T_67126; // @[Modules.scala 150:103:@13521.4]
  wire [5:0] _T_67130; // @[Modules.scala 151:80:@13524.4]
  wire [6:0] _T_67131; // @[Modules.scala 150:103:@13525.4]
  wire [5:0] _T_67132; // @[Modules.scala 150:103:@13526.4]
  wire [5:0] _T_67133; // @[Modules.scala 150:103:@13527.4]
  wire [5:0] _T_67135; // @[Modules.scala 150:74:@13529.4]
  wire [6:0] _T_67138; // @[Modules.scala 150:103:@13531.4]
  wire [5:0] _T_67139; // @[Modules.scala 150:103:@13532.4]
  wire [5:0] _T_67140; // @[Modules.scala 150:103:@13533.4]
  wire [6:0] _T_67145; // @[Modules.scala 150:103:@13537.4]
  wire [5:0] _T_67146; // @[Modules.scala 150:103:@13538.4]
  wire [5:0] _T_67147; // @[Modules.scala 150:103:@13539.4]
  wire [6:0] _T_67152; // @[Modules.scala 150:103:@13543.4]
  wire [5:0] _T_67153; // @[Modules.scala 150:103:@13544.4]
  wire [5:0] _T_67154; // @[Modules.scala 150:103:@13545.4]
  wire [6:0] _T_67187; // @[Modules.scala 150:103:@13573.4]
  wire [5:0] _T_67188; // @[Modules.scala 150:103:@13574.4]
  wire [5:0] _T_67189; // @[Modules.scala 150:103:@13575.4]
  wire [5:0] _T_67200; // @[Modules.scala 151:80:@13584.4]
  wire [6:0] _T_67201; // @[Modules.scala 150:103:@13585.4]
  wire [5:0] _T_67202; // @[Modules.scala 150:103:@13586.4]
  wire [5:0] _T_67203; // @[Modules.scala 150:103:@13587.4]
  wire [5:0] _GEN_302; // @[Modules.scala 150:103:@13591.4]
  wire [6:0] _T_67208; // @[Modules.scala 150:103:@13591.4]
  wire [5:0] _T_67209; // @[Modules.scala 150:103:@13592.4]
  wire [5:0] _T_67210; // @[Modules.scala 150:103:@13593.4]
  wire [6:0] _T_67215; // @[Modules.scala 150:103:@13597.4]
  wire [5:0] _T_67216; // @[Modules.scala 150:103:@13598.4]
  wire [5:0] _T_67217; // @[Modules.scala 150:103:@13599.4]
  wire [6:0] _T_67222; // @[Modules.scala 150:103:@13603.4]
  wire [5:0] _T_67223; // @[Modules.scala 150:103:@13604.4]
  wire [5:0] _T_67224; // @[Modules.scala 150:103:@13605.4]
  wire [5:0] _T_67247; // @[Modules.scala 150:74:@13625.4]
  wire [5:0] _GEN_304; // @[Modules.scala 150:103:@13627.4]
  wire [6:0] _T_67250; // @[Modules.scala 150:103:@13627.4]
  wire [5:0] _T_67251; // @[Modules.scala 150:103:@13628.4]
  wire [5:0] _T_67252; // @[Modules.scala 150:103:@13629.4]
  wire [5:0] _T_67264; // @[Modules.scala 150:103:@13639.4]
  wire [4:0] _T_67265; // @[Modules.scala 150:103:@13640.4]
  wire [4:0] _T_67266; // @[Modules.scala 150:103:@13641.4]
  wire [6:0] _T_67271; // @[Modules.scala 150:103:@13645.4]
  wire [5:0] _T_67272; // @[Modules.scala 150:103:@13646.4]
  wire [5:0] _T_67273; // @[Modules.scala 150:103:@13647.4]
  wire [6:0] _T_67278; // @[Modules.scala 150:103:@13651.4]
  wire [5:0] _T_67279; // @[Modules.scala 150:103:@13652.4]
  wire [5:0] _T_67280; // @[Modules.scala 150:103:@13653.4]
  wire [6:0] _T_67285; // @[Modules.scala 150:103:@13657.4]
  wire [5:0] _T_67286; // @[Modules.scala 150:103:@13658.4]
  wire [5:0] _T_67287; // @[Modules.scala 150:103:@13659.4]
  wire [6:0] _T_67299; // @[Modules.scala 150:103:@13669.4]
  wire [5:0] _T_67300; // @[Modules.scala 150:103:@13670.4]
  wire [5:0] _T_67301; // @[Modules.scala 150:103:@13671.4]
  wire [6:0] _T_67306; // @[Modules.scala 150:103:@13675.4]
  wire [5:0] _T_67307; // @[Modules.scala 150:103:@13676.4]
  wire [5:0] _T_67308; // @[Modules.scala 150:103:@13677.4]
  wire [5:0] _GEN_306; // @[Modules.scala 150:103:@13681.4]
  wire [6:0] _T_67313; // @[Modules.scala 150:103:@13681.4]
  wire [5:0] _T_67314; // @[Modules.scala 150:103:@13682.4]
  wire [5:0] _T_67315; // @[Modules.scala 150:103:@13683.4]
  wire [5:0] _T_67324; // @[Modules.scala 150:74:@13691.4]
  wire [5:0] _GEN_307; // @[Modules.scala 150:103:@13693.4]
  wire [6:0] _T_67327; // @[Modules.scala 150:103:@13693.4]
  wire [5:0] _T_67328; // @[Modules.scala 150:103:@13694.4]
  wire [5:0] _T_67329; // @[Modules.scala 150:103:@13695.4]
  wire [4:0] _T_67340; // @[Modules.scala 151:80:@13704.4]
  wire [5:0] _T_67341; // @[Modules.scala 150:103:@13705.4]
  wire [4:0] _T_67342; // @[Modules.scala 150:103:@13706.4]
  wire [4:0] _T_67343; // @[Modules.scala 150:103:@13707.4]
  wire [5:0] _GEN_308; // @[Modules.scala 150:103:@13711.4]
  wire [6:0] _T_67348; // @[Modules.scala 150:103:@13711.4]
  wire [5:0] _T_67349; // @[Modules.scala 150:103:@13712.4]
  wire [5:0] _T_67350; // @[Modules.scala 150:103:@13713.4]
  wire [5:0] _GEN_309; // @[Modules.scala 150:103:@13729.4]
  wire [6:0] _T_67369; // @[Modules.scala 150:103:@13729.4]
  wire [5:0] _T_67370; // @[Modules.scala 150:103:@13730.4]
  wire [5:0] _T_67371; // @[Modules.scala 150:103:@13731.4]
  wire [5:0] _GEN_310; // @[Modules.scala 150:103:@13741.4]
  wire [6:0] _T_67383; // @[Modules.scala 150:103:@13741.4]
  wire [5:0] _T_67384; // @[Modules.scala 150:103:@13742.4]
  wire [5:0] _T_67385; // @[Modules.scala 150:103:@13743.4]
  wire [5:0] _GEN_311; // @[Modules.scala 150:103:@13747.4]
  wire [6:0] _T_67390; // @[Modules.scala 150:103:@13747.4]
  wire [5:0] _T_67391; // @[Modules.scala 150:103:@13748.4]
  wire [5:0] _T_67392; // @[Modules.scala 150:103:@13749.4]
  wire [5:0] _GEN_312; // @[Modules.scala 150:103:@13753.4]
  wire [6:0] _T_67397; // @[Modules.scala 150:103:@13753.4]
  wire [5:0] _T_67398; // @[Modules.scala 150:103:@13754.4]
  wire [5:0] _T_67399; // @[Modules.scala 150:103:@13755.4]
  wire [6:0] _T_67411; // @[Modules.scala 150:103:@13765.4]
  wire [5:0] _T_67412; // @[Modules.scala 150:103:@13766.4]
  wire [5:0] _T_67413; // @[Modules.scala 150:103:@13767.4]
  wire [5:0] _T_67425; // @[Modules.scala 150:103:@13777.4]
  wire [4:0] _T_67426; // @[Modules.scala 150:103:@13778.4]
  wire [4:0] _T_67427; // @[Modules.scala 150:103:@13779.4]
  wire [5:0] _GEN_314; // @[Modules.scala 150:103:@13789.4]
  wire [6:0] _T_67439; // @[Modules.scala 150:103:@13789.4]
  wire [5:0] _T_67440; // @[Modules.scala 150:103:@13790.4]
  wire [5:0] _T_67441; // @[Modules.scala 150:103:@13791.4]
  wire [5:0] _GEN_316; // @[Modules.scala 150:103:@13813.4]
  wire [6:0] _T_67467; // @[Modules.scala 150:103:@13813.4]
  wire [5:0] _T_67468; // @[Modules.scala 150:103:@13814.4]
  wire [5:0] _T_67469; // @[Modules.scala 150:103:@13815.4]
  wire [6:0] _T_67474; // @[Modules.scala 150:103:@13819.4]
  wire [5:0] _T_67475; // @[Modules.scala 150:103:@13820.4]
  wire [5:0] _T_67476; // @[Modules.scala 150:103:@13821.4]
  wire [5:0] _GEN_317; // @[Modules.scala 150:103:@13831.4]
  wire [6:0] _T_67488; // @[Modules.scala 150:103:@13831.4]
  wire [5:0] _T_67489; // @[Modules.scala 150:103:@13832.4]
  wire [5:0] _T_67490; // @[Modules.scala 150:103:@13833.4]
  wire [5:0] _T_67502; // @[Modules.scala 150:103:@13843.4]
  wire [4:0] _T_67503; // @[Modules.scala 150:103:@13844.4]
  wire [4:0] _T_67504; // @[Modules.scala 150:103:@13845.4]
  wire [6:0] _T_67509; // @[Modules.scala 150:103:@13849.4]
  wire [5:0] _T_67510; // @[Modules.scala 150:103:@13850.4]
  wire [5:0] _T_67511; // @[Modules.scala 150:103:@13851.4]
  wire [6:0] _T_67516; // @[Modules.scala 150:103:@13855.4]
  wire [5:0] _T_67517; // @[Modules.scala 150:103:@13856.4]
  wire [5:0] _T_67518; // @[Modules.scala 150:103:@13857.4]
  wire [4:0] _T_67550; // @[Modules.scala 151:80:@13884.4]
  wire [5:0] _T_67551; // @[Modules.scala 150:103:@13885.4]
  wire [4:0] _T_67552; // @[Modules.scala 150:103:@13886.4]
  wire [4:0] _T_67553; // @[Modules.scala 150:103:@13887.4]
  wire [6:0] _T_67565; // @[Modules.scala 150:103:@13897.4]
  wire [5:0] _T_67566; // @[Modules.scala 150:103:@13898.4]
  wire [5:0] _T_67567; // @[Modules.scala 150:103:@13899.4]
  wire [5:0] _T_67585; // @[Modules.scala 151:80:@13914.4]
  wire [6:0] _T_67586; // @[Modules.scala 150:103:@13915.4]
  wire [5:0] _T_67587; // @[Modules.scala 150:103:@13916.4]
  wire [5:0] _T_67588; // @[Modules.scala 150:103:@13917.4]
  wire [4:0] _T_67597; // @[Modules.scala 150:74:@13925.4]
  wire [5:0] _GEN_321; // @[Modules.scala 150:103:@13927.4]
  wire [6:0] _T_67600; // @[Modules.scala 150:103:@13927.4]
  wire [5:0] _T_67601; // @[Modules.scala 150:103:@13928.4]
  wire [5:0] _T_67602; // @[Modules.scala 150:103:@13929.4]
  wire [5:0] _T_67614; // @[Modules.scala 150:103:@13939.4]
  wire [4:0] _T_67615; // @[Modules.scala 150:103:@13940.4]
  wire [4:0] _T_67616; // @[Modules.scala 150:103:@13941.4]
  wire [5:0] _T_67621; // @[Modules.scala 150:103:@13945.4]
  wire [4:0] _T_67622; // @[Modules.scala 150:103:@13946.4]
  wire [4:0] _T_67623; // @[Modules.scala 150:103:@13947.4]
  wire [6:0] _T_67628; // @[Modules.scala 150:103:@13951.4]
  wire [5:0] _T_67629; // @[Modules.scala 150:103:@13952.4]
  wire [5:0] _T_67630; // @[Modules.scala 150:103:@13953.4]
  wire [6:0] _T_67635; // @[Modules.scala 150:103:@13957.4]
  wire [5:0] _T_67636; // @[Modules.scala 150:103:@13958.4]
  wire [5:0] _T_67637; // @[Modules.scala 150:103:@13959.4]
  wire [5:0] _GEN_323; // @[Modules.scala 150:103:@13963.4]
  wire [6:0] _T_67642; // @[Modules.scala 150:103:@13963.4]
  wire [5:0] _T_67643; // @[Modules.scala 150:103:@13964.4]
  wire [5:0] _T_67644; // @[Modules.scala 150:103:@13965.4]
  wire [5:0] _GEN_324; // @[Modules.scala 150:103:@13981.4]
  wire [6:0] _T_67663; // @[Modules.scala 150:103:@13981.4]
  wire [5:0] _T_67664; // @[Modules.scala 150:103:@13982.4]
  wire [5:0] _T_67665; // @[Modules.scala 150:103:@13983.4]
  wire [5:0] _T_67670; // @[Modules.scala 150:103:@13987.4]
  wire [4:0] _T_67671; // @[Modules.scala 150:103:@13988.4]
  wire [4:0] _T_67672; // @[Modules.scala 150:103:@13989.4]
  wire [5:0] _GEN_325; // @[Modules.scala 150:103:@13993.4]
  wire [6:0] _T_67677; // @[Modules.scala 150:103:@13993.4]
  wire [5:0] _T_67678; // @[Modules.scala 150:103:@13994.4]
  wire [5:0] _T_67679; // @[Modules.scala 150:103:@13995.4]
  wire [5:0] _T_67684; // @[Modules.scala 150:103:@13999.4]
  wire [4:0] _T_67685; // @[Modules.scala 150:103:@14000.4]
  wire [4:0] _T_67686; // @[Modules.scala 150:103:@14001.4]
  wire [5:0] _T_67691; // @[Modules.scala 150:103:@14005.4]
  wire [4:0] _T_67692; // @[Modules.scala 150:103:@14006.4]
  wire [4:0] _T_67693; // @[Modules.scala 150:103:@14007.4]
  wire [4:0] _T_67695; // @[Modules.scala 150:74:@14009.4]
  wire [5:0] _T_67698; // @[Modules.scala 150:103:@14011.4]
  wire [4:0] _T_67699; // @[Modules.scala 150:103:@14012.4]
  wire [4:0] _T_67700; // @[Modules.scala 150:103:@14013.4]
  wire [6:0] _T_67705; // @[Modules.scala 150:103:@14017.4]
  wire [5:0] _T_67706; // @[Modules.scala 150:103:@14018.4]
  wire [5:0] _T_67707; // @[Modules.scala 150:103:@14019.4]
  wire [6:0] _T_67747; // @[Modules.scala 150:103:@14053.4]
  wire [5:0] _T_67748; // @[Modules.scala 150:103:@14054.4]
  wire [5:0] _T_67749; // @[Modules.scala 150:103:@14055.4]
  wire [5:0] _GEN_330; // @[Modules.scala 150:103:@14059.4]
  wire [6:0] _T_67754; // @[Modules.scala 150:103:@14059.4]
  wire [5:0] _T_67755; // @[Modules.scala 150:103:@14060.4]
  wire [5:0] _T_67756; // @[Modules.scala 150:103:@14061.4]
  wire [5:0] _GEN_331; // @[Modules.scala 150:103:@14065.4]
  wire [6:0] _T_67761; // @[Modules.scala 150:103:@14065.4]
  wire [5:0] _T_67762; // @[Modules.scala 150:103:@14066.4]
  wire [5:0] _T_67763; // @[Modules.scala 150:103:@14067.4]
  wire [5:0] _T_67765; // @[Modules.scala 150:74:@14069.4]
  wire [5:0] _T_67767; // @[Modules.scala 151:80:@14070.4]
  wire [6:0] _T_67768; // @[Modules.scala 150:103:@14071.4]
  wire [5:0] _T_67769; // @[Modules.scala 150:103:@14072.4]
  wire [5:0] _T_67770; // @[Modules.scala 150:103:@14073.4]
  wire [6:0] _T_67775; // @[Modules.scala 150:103:@14077.4]
  wire [5:0] _T_67776; // @[Modules.scala 150:103:@14078.4]
  wire [5:0] _T_67777; // @[Modules.scala 150:103:@14079.4]
  wire [6:0] _T_67796; // @[Modules.scala 150:103:@14095.4]
  wire [5:0] _T_67797; // @[Modules.scala 150:103:@14096.4]
  wire [5:0] _T_67798; // @[Modules.scala 150:103:@14097.4]
  wire [5:0] _T_67817; // @[Modules.scala 150:103:@14113.4]
  wire [4:0] _T_67818; // @[Modules.scala 150:103:@14114.4]
  wire [4:0] _T_67819; // @[Modules.scala 150:103:@14115.4]
  wire [5:0] _T_67824; // @[Modules.scala 150:103:@14119.4]
  wire [4:0] _T_67825; // @[Modules.scala 150:103:@14120.4]
  wire [4:0] _T_67826; // @[Modules.scala 150:103:@14121.4]
  wire [5:0] _T_67831; // @[Modules.scala 150:103:@14125.4]
  wire [4:0] _T_67832; // @[Modules.scala 150:103:@14126.4]
  wire [4:0] _T_67833; // @[Modules.scala 150:103:@14127.4]
  wire [6:0] _T_67845; // @[Modules.scala 150:103:@14137.4]
  wire [5:0] _T_67846; // @[Modules.scala 150:103:@14138.4]
  wire [5:0] _T_67847; // @[Modules.scala 150:103:@14139.4]
  wire [5:0] _GEN_335; // @[Modules.scala 150:103:@14161.4]
  wire [6:0] _T_67873; // @[Modules.scala 150:103:@14161.4]
  wire [5:0] _T_67874; // @[Modules.scala 150:103:@14162.4]
  wire [5:0] _T_67875; // @[Modules.scala 150:103:@14163.4]
  wire [5:0] _T_67901; // @[Modules.scala 150:103:@14185.4]
  wire [4:0] _T_67902; // @[Modules.scala 150:103:@14186.4]
  wire [4:0] _T_67903; // @[Modules.scala 150:103:@14187.4]
  wire [5:0] _GEN_336; // @[Modules.scala 150:103:@14191.4]
  wire [6:0] _T_67908; // @[Modules.scala 150:103:@14191.4]
  wire [5:0] _T_67909; // @[Modules.scala 150:103:@14192.4]
  wire [5:0] _T_67910; // @[Modules.scala 150:103:@14193.4]
  wire [4:0] _T_67928; // @[Modules.scala 151:80:@14208.4]
  wire [5:0] _T_67929; // @[Modules.scala 150:103:@14209.4]
  wire [4:0] _T_67930; // @[Modules.scala 150:103:@14210.4]
  wire [4:0] _T_67931; // @[Modules.scala 150:103:@14211.4]
  wire [5:0] _T_67943; // @[Modules.scala 150:103:@14221.4]
  wire [4:0] _T_67944; // @[Modules.scala 150:103:@14222.4]
  wire [4:0] _T_67945; // @[Modules.scala 150:103:@14223.4]
  wire [6:0] _T_67950; // @[Modules.scala 150:103:@14227.4]
  wire [5:0] _T_67951; // @[Modules.scala 150:103:@14228.4]
  wire [5:0] _T_67952; // @[Modules.scala 150:103:@14229.4]
  wire [5:0] _GEN_338; // @[Modules.scala 150:103:@14233.4]
  wire [6:0] _T_67957; // @[Modules.scala 150:103:@14233.4]
  wire [5:0] _T_67958; // @[Modules.scala 150:103:@14234.4]
  wire [5:0] _T_67959; // @[Modules.scala 150:103:@14235.4]
  wire [4:0] _T_67991; // @[Modules.scala 151:80:@14262.4]
  wire [5:0] _GEN_339; // @[Modules.scala 150:103:@14263.4]
  wire [6:0] _T_67992; // @[Modules.scala 150:103:@14263.4]
  wire [5:0] _T_67993; // @[Modules.scala 150:103:@14264.4]
  wire [5:0] _T_67994; // @[Modules.scala 150:103:@14265.4]
  wire [5:0] _T_67999; // @[Modules.scala 150:103:@14269.4]
  wire [4:0] _T_68000; // @[Modules.scala 150:103:@14270.4]
  wire [4:0] _T_68001; // @[Modules.scala 150:103:@14271.4]
  wire [5:0] _T_68006; // @[Modules.scala 150:103:@14275.4]
  wire [4:0] _T_68007; // @[Modules.scala 150:103:@14276.4]
  wire [4:0] _T_68008; // @[Modules.scala 150:103:@14277.4]
  wire [5:0] _GEN_340; // @[Modules.scala 150:103:@14287.4]
  wire [6:0] _T_68020; // @[Modules.scala 150:103:@14287.4]
  wire [5:0] _T_68021; // @[Modules.scala 150:103:@14288.4]
  wire [5:0] _T_68022; // @[Modules.scala 150:103:@14289.4]
  wire [5:0] _GEN_341; // @[Modules.scala 150:103:@14293.4]
  wire [6:0] _T_68027; // @[Modules.scala 150:103:@14293.4]
  wire [5:0] _T_68028; // @[Modules.scala 150:103:@14294.4]
  wire [5:0] _T_68029; // @[Modules.scala 150:103:@14295.4]
  wire [5:0] _GEN_342; // @[Modules.scala 150:103:@14299.4]
  wire [6:0] _T_68034; // @[Modules.scala 150:103:@14299.4]
  wire [5:0] _T_68035; // @[Modules.scala 150:103:@14300.4]
  wire [5:0] _T_68036; // @[Modules.scala 150:103:@14301.4]
  wire [4:0] _T_68038; // @[Modules.scala 150:74:@14303.4]
  wire [5:0] _T_68041; // @[Modules.scala 150:103:@14305.4]
  wire [4:0] _T_68042; // @[Modules.scala 150:103:@14306.4]
  wire [4:0] _T_68043; // @[Modules.scala 150:103:@14307.4]
  wire [6:0] _T_68069; // @[Modules.scala 150:103:@14329.4]
  wire [5:0] _T_68070; // @[Modules.scala 150:103:@14330.4]
  wire [5:0] _T_68071; // @[Modules.scala 150:103:@14331.4]
  wire [4:0] _T_68075; // @[Modules.scala 151:80:@14334.4]
  wire [5:0] _T_68076; // @[Modules.scala 150:103:@14335.4]
  wire [4:0] _T_68077; // @[Modules.scala 150:103:@14336.4]
  wire [4:0] _T_68078; // @[Modules.scala 150:103:@14337.4]
  wire [5:0] _T_68083; // @[Modules.scala 150:103:@14341.4]
  wire [4:0] _T_68084; // @[Modules.scala 150:103:@14342.4]
  wire [4:0] _T_68085; // @[Modules.scala 150:103:@14343.4]
  wire [5:0] _T_68090; // @[Modules.scala 150:103:@14347.4]
  wire [4:0] _T_68091; // @[Modules.scala 150:103:@14348.4]
  wire [4:0] _T_68092; // @[Modules.scala 150:103:@14349.4]
  wire [5:0] _T_68111; // @[Modules.scala 150:103:@14365.4]
  wire [4:0] _T_68112; // @[Modules.scala 150:103:@14366.4]
  wire [4:0] _T_68113; // @[Modules.scala 150:103:@14367.4]
  wire [5:0] _T_68118; // @[Modules.scala 150:103:@14371.4]
  wire [4:0] _T_68119; // @[Modules.scala 150:103:@14372.4]
  wire [4:0] _T_68120; // @[Modules.scala 150:103:@14373.4]
  wire [5:0] _T_68153; // @[Modules.scala 150:103:@14401.4]
  wire [4:0] _T_68154; // @[Modules.scala 150:103:@14402.4]
  wire [4:0] _T_68155; // @[Modules.scala 150:103:@14403.4]
  wire [4:0] _T_68171; // @[Modules.scala 150:74:@14417.4]
  wire [5:0] _T_68174; // @[Modules.scala 150:103:@14419.4]
  wire [4:0] _T_68175; // @[Modules.scala 150:103:@14420.4]
  wire [4:0] _T_68176; // @[Modules.scala 150:103:@14421.4]
  wire [5:0] _T_68181; // @[Modules.scala 150:103:@14425.4]
  wire [4:0] _T_68182; // @[Modules.scala 150:103:@14426.4]
  wire [4:0] _T_68183; // @[Modules.scala 150:103:@14427.4]
  wire [5:0] _GEN_344; // @[Modules.scala 150:103:@14431.4]
  wire [6:0] _T_68188; // @[Modules.scala 150:103:@14431.4]
  wire [5:0] _T_68189; // @[Modules.scala 150:103:@14432.4]
  wire [5:0] _T_68190; // @[Modules.scala 150:103:@14433.4]
  wire [4:0] _T_68194; // @[Modules.scala 151:80:@14436.4]
  wire [5:0] _GEN_345; // @[Modules.scala 150:103:@14437.4]
  wire [6:0] _T_68195; // @[Modules.scala 150:103:@14437.4]
  wire [5:0] _T_68196; // @[Modules.scala 150:103:@14438.4]
  wire [5:0] _T_68197; // @[Modules.scala 150:103:@14439.4]
  wire [5:0] _T_68202; // @[Modules.scala 150:103:@14443.4]
  wire [4:0] _T_68203; // @[Modules.scala 150:103:@14444.4]
  wire [4:0] _T_68204; // @[Modules.scala 150:103:@14445.4]
  wire [5:0] _T_68209; // @[Modules.scala 150:103:@14449.4]
  wire [4:0] _T_68210; // @[Modules.scala 150:103:@14450.4]
  wire [4:0] _T_68211; // @[Modules.scala 150:103:@14451.4]
  wire [5:0] _GEN_346; // @[Modules.scala 150:103:@14455.4]
  wire [6:0] _T_68216; // @[Modules.scala 150:103:@14455.4]
  wire [5:0] _T_68217; // @[Modules.scala 150:103:@14456.4]
  wire [5:0] _T_68218; // @[Modules.scala 150:103:@14457.4]
  wire [5:0] _T_68220; // @[Modules.scala 150:74:@14459.4]
  wire [5:0] _GEN_347; // @[Modules.scala 150:103:@14461.4]
  wire [6:0] _T_68223; // @[Modules.scala 150:103:@14461.4]
  wire [5:0] _T_68224; // @[Modules.scala 150:103:@14462.4]
  wire [5:0] _T_68225; // @[Modules.scala 150:103:@14463.4]
  wire [5:0] _GEN_348; // @[Modules.scala 150:103:@14479.4]
  wire [6:0] _T_68244; // @[Modules.scala 150:103:@14479.4]
  wire [5:0] _T_68245; // @[Modules.scala 150:103:@14480.4]
  wire [5:0] _T_68246; // @[Modules.scala 150:103:@14481.4]
  wire [5:0] _T_68251; // @[Modules.scala 150:103:@14485.4]
  wire [4:0] _T_68252; // @[Modules.scala 150:103:@14486.4]
  wire [4:0] _T_68253; // @[Modules.scala 150:103:@14487.4]
  wire [5:0] _T_68257; // @[Modules.scala 151:80:@14490.4]
  wire [5:0] _GEN_349; // @[Modules.scala 150:103:@14491.4]
  wire [6:0] _T_68258; // @[Modules.scala 150:103:@14491.4]
  wire [5:0] _T_68259; // @[Modules.scala 150:103:@14492.4]
  wire [5:0] _T_68260; // @[Modules.scala 150:103:@14493.4]
  wire [5:0] _GEN_351; // @[Modules.scala 150:103:@14509.4]
  wire [6:0] _T_68279; // @[Modules.scala 150:103:@14509.4]
  wire [5:0] _T_68280; // @[Modules.scala 150:103:@14510.4]
  wire [5:0] _T_68281; // @[Modules.scala 150:103:@14511.4]
  wire [5:0] _GEN_352; // @[Modules.scala 150:103:@14515.4]
  wire [6:0] _T_68286; // @[Modules.scala 150:103:@14515.4]
  wire [5:0] _T_68287; // @[Modules.scala 150:103:@14516.4]
  wire [5:0] _T_68288; // @[Modules.scala 150:103:@14517.4]
  wire [5:0] _T_68293; // @[Modules.scala 150:103:@14521.4]
  wire [4:0] _T_68294; // @[Modules.scala 150:103:@14522.4]
  wire [4:0] _T_68295; // @[Modules.scala 150:103:@14523.4]
  wire [5:0] _T_68300; // @[Modules.scala 150:103:@14527.4]
  wire [4:0] _T_68301; // @[Modules.scala 150:103:@14528.4]
  wire [4:0] _T_68302; // @[Modules.scala 150:103:@14529.4]
  wire [5:0] _GEN_353; // @[Modules.scala 150:103:@14545.4]
  wire [6:0] _T_68321; // @[Modules.scala 150:103:@14545.4]
  wire [5:0] _T_68322; // @[Modules.scala 150:103:@14546.4]
  wire [5:0] _T_68323; // @[Modules.scala 150:103:@14547.4]
  wire [6:0] _T_68335; // @[Modules.scala 150:103:@14557.4]
  wire [5:0] _T_68336; // @[Modules.scala 150:103:@14558.4]
  wire [5:0] _T_68337; // @[Modules.scala 150:103:@14559.4]
  wire [4:0] _T_68341; // @[Modules.scala 151:80:@14562.4]
  wire [5:0] _T_68342; // @[Modules.scala 150:103:@14563.4]
  wire [4:0] _T_68343; // @[Modules.scala 150:103:@14564.4]
  wire [4:0] _T_68344; // @[Modules.scala 150:103:@14565.4]
  wire [5:0] _T_68349; // @[Modules.scala 150:103:@14569.4]
  wire [4:0] _T_68350; // @[Modules.scala 150:103:@14570.4]
  wire [4:0] _T_68351; // @[Modules.scala 150:103:@14571.4]
  wire [5:0] _GEN_354; // @[Modules.scala 150:103:@14575.4]
  wire [6:0] _T_68356; // @[Modules.scala 150:103:@14575.4]
  wire [5:0] _T_68357; // @[Modules.scala 150:103:@14576.4]
  wire [5:0] _T_68358; // @[Modules.scala 150:103:@14577.4]
  wire [5:0] _T_68423; // @[Modules.scala 150:74:@14633.4]
  wire [6:0] _T_68426; // @[Modules.scala 150:103:@14635.4]
  wire [5:0] _T_68427; // @[Modules.scala 150:103:@14636.4]
  wire [5:0] _T_68428; // @[Modules.scala 150:103:@14637.4]
  wire [6:0] _T_68433; // @[Modules.scala 150:103:@14641.4]
  wire [5:0] _T_68434; // @[Modules.scala 150:103:@14642.4]
  wire [5:0] _T_68435; // @[Modules.scala 150:103:@14643.4]
  wire [6:0] _T_68447; // @[Modules.scala 150:103:@14653.4]
  wire [5:0] _T_68448; // @[Modules.scala 150:103:@14654.4]
  wire [5:0] _T_68449; // @[Modules.scala 150:103:@14655.4]
  wire [6:0] _T_68454; // @[Modules.scala 150:103:@14659.4]
  wire [5:0] _T_68455; // @[Modules.scala 150:103:@14660.4]
  wire [5:0] _T_68456; // @[Modules.scala 150:103:@14661.4]
  wire [6:0] _T_68461; // @[Modules.scala 150:103:@14665.4]
  wire [5:0] _T_68462; // @[Modules.scala 150:103:@14666.4]
  wire [5:0] _T_68463; // @[Modules.scala 150:103:@14667.4]
  wire [6:0] _T_68468; // @[Modules.scala 150:103:@14671.4]
  wire [5:0] _T_68469; // @[Modules.scala 150:103:@14672.4]
  wire [5:0] _T_68470; // @[Modules.scala 150:103:@14673.4]
  wire [6:0] _T_68475; // @[Modules.scala 150:103:@14677.4]
  wire [5:0] _T_68476; // @[Modules.scala 150:103:@14678.4]
  wire [5:0] _T_68477; // @[Modules.scala 150:103:@14679.4]
  wire [6:0] _T_68482; // @[Modules.scala 150:103:@14683.4]
  wire [5:0] _T_68483; // @[Modules.scala 150:103:@14684.4]
  wire [5:0] _T_68484; // @[Modules.scala 150:103:@14685.4]
  wire [6:0] _T_68489; // @[Modules.scala 150:103:@14689.4]
  wire [5:0] _T_68490; // @[Modules.scala 150:103:@14690.4]
  wire [5:0] _T_68491; // @[Modules.scala 150:103:@14691.4]
  wire [6:0] _T_68496; // @[Modules.scala 150:103:@14695.4]
  wire [5:0] _T_68497; // @[Modules.scala 150:103:@14696.4]
  wire [5:0] _T_68498; // @[Modules.scala 150:103:@14697.4]
  wire [5:0] _T_68500; // @[Modules.scala 150:74:@14699.4]
  wire [5:0] _T_68502; // @[Modules.scala 151:80:@14700.4]
  wire [6:0] _T_68503; // @[Modules.scala 150:103:@14701.4]
  wire [5:0] _T_68504; // @[Modules.scala 150:103:@14702.4]
  wire [5:0] _T_68505; // @[Modules.scala 150:103:@14703.4]
  wire [5:0] _T_68523; // @[Modules.scala 151:80:@14718.4]
  wire [6:0] _T_68524; // @[Modules.scala 150:103:@14719.4]
  wire [5:0] _T_68525; // @[Modules.scala 150:103:@14720.4]
  wire [5:0] _T_68526; // @[Modules.scala 150:103:@14721.4]
  wire [5:0] _GEN_356; // @[Modules.scala 150:103:@14743.4]
  wire [6:0] _T_68552; // @[Modules.scala 150:103:@14743.4]
  wire [5:0] _T_68553; // @[Modules.scala 150:103:@14744.4]
  wire [5:0] _T_68554; // @[Modules.scala 150:103:@14745.4]
  wire [13:0] buffer_4_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68574; // @[Modules.scala 160:64:@14765.4]
  wire [13:0] _T_68575; // @[Modules.scala 160:64:@14766.4]
  wire [13:0] buffer_4_301; // @[Modules.scala 160:64:@14767.4]
  wire [13:0] buffer_4_4; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68577; // @[Modules.scala 160:64:@14769.4]
  wire [13:0] _T_68578; // @[Modules.scala 160:64:@14770.4]
  wire [13:0] buffer_4_302; // @[Modules.scala 160:64:@14771.4]
  wire [13:0] buffer_4_6; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_7; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68580; // @[Modules.scala 160:64:@14773.4]
  wire [13:0] _T_68581; // @[Modules.scala 160:64:@14774.4]
  wire [13:0] buffer_4_303; // @[Modules.scala 160:64:@14775.4]
  wire [13:0] buffer_4_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68583; // @[Modules.scala 160:64:@14777.4]
  wire [13:0] _T_68584; // @[Modules.scala 160:64:@14778.4]
  wire [13:0] buffer_4_304; // @[Modules.scala 160:64:@14779.4]
  wire [13:0] buffer_4_10; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68586; // @[Modules.scala 160:64:@14781.4]
  wire [13:0] _T_68587; // @[Modules.scala 160:64:@14782.4]
  wire [13:0] buffer_4_305; // @[Modules.scala 160:64:@14783.4]
  wire [13:0] buffer_4_12; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68589; // @[Modules.scala 160:64:@14785.4]
  wire [13:0] _T_68590; // @[Modules.scala 160:64:@14786.4]
  wire [13:0] buffer_4_306; // @[Modules.scala 160:64:@14787.4]
  wire [14:0] _T_68595; // @[Modules.scala 160:64:@14793.4]
  wire [13:0] _T_68596; // @[Modules.scala 160:64:@14794.4]
  wire [13:0] buffer_4_308; // @[Modules.scala 160:64:@14795.4]
  wire [13:0] buffer_4_18; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_19; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68598; // @[Modules.scala 160:64:@14797.4]
  wire [13:0] _T_68599; // @[Modules.scala 160:64:@14798.4]
  wire [13:0] buffer_4_309; // @[Modules.scala 160:64:@14799.4]
  wire [13:0] buffer_4_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68601; // @[Modules.scala 160:64:@14801.4]
  wire [13:0] _T_68602; // @[Modules.scala 160:64:@14802.4]
  wire [13:0] buffer_4_310; // @[Modules.scala 160:64:@14803.4]
  wire [14:0] _T_68604; // @[Modules.scala 160:64:@14805.4]
  wire [13:0] _T_68605; // @[Modules.scala 160:64:@14806.4]
  wire [13:0] buffer_4_311; // @[Modules.scala 160:64:@14807.4]
  wire [14:0] _T_68607; // @[Modules.scala 160:64:@14809.4]
  wire [13:0] _T_68608; // @[Modules.scala 160:64:@14810.4]
  wire [13:0] buffer_4_312; // @[Modules.scala 160:64:@14811.4]
  wire [14:0] _T_68610; // @[Modules.scala 160:64:@14813.4]
  wire [13:0] _T_68611; // @[Modules.scala 160:64:@14814.4]
  wire [13:0] buffer_4_313; // @[Modules.scala 160:64:@14815.4]
  wire [14:0] _T_68613; // @[Modules.scala 160:64:@14817.4]
  wire [13:0] _T_68614; // @[Modules.scala 160:64:@14818.4]
  wire [13:0] buffer_4_314; // @[Modules.scala 160:64:@14819.4]
  wire [13:0] buffer_4_30; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_31; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68616; // @[Modules.scala 160:64:@14821.4]
  wire [13:0] _T_68617; // @[Modules.scala 160:64:@14822.4]
  wire [13:0] buffer_4_315; // @[Modules.scala 160:64:@14823.4]
  wire [13:0] buffer_4_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68619; // @[Modules.scala 160:64:@14825.4]
  wire [13:0] _T_68620; // @[Modules.scala 160:64:@14826.4]
  wire [13:0] buffer_4_316; // @[Modules.scala 160:64:@14827.4]
  wire [13:0] buffer_4_34; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68622; // @[Modules.scala 160:64:@14829.4]
  wire [13:0] _T_68623; // @[Modules.scala 160:64:@14830.4]
  wire [13:0] buffer_4_317; // @[Modules.scala 160:64:@14831.4]
  wire [13:0] buffer_4_36; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_37; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68625; // @[Modules.scala 160:64:@14833.4]
  wire [13:0] _T_68626; // @[Modules.scala 160:64:@14834.4]
  wire [13:0] buffer_4_318; // @[Modules.scala 160:64:@14835.4]
  wire [13:0] buffer_4_39; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68628; // @[Modules.scala 160:64:@14837.4]
  wire [13:0] _T_68629; // @[Modules.scala 160:64:@14838.4]
  wire [13:0] buffer_4_319; // @[Modules.scala 160:64:@14839.4]
  wire [13:0] buffer_4_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68631; // @[Modules.scala 160:64:@14841.4]
  wire [13:0] _T_68632; // @[Modules.scala 160:64:@14842.4]
  wire [13:0] buffer_4_320; // @[Modules.scala 160:64:@14843.4]
  wire [13:0] buffer_4_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68634; // @[Modules.scala 160:64:@14845.4]
  wire [13:0] _T_68635; // @[Modules.scala 160:64:@14846.4]
  wire [13:0] buffer_4_321; // @[Modules.scala 160:64:@14847.4]
  wire [13:0] buffer_4_44; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68637; // @[Modules.scala 160:64:@14849.4]
  wire [13:0] _T_68638; // @[Modules.scala 160:64:@14850.4]
  wire [13:0] buffer_4_322; // @[Modules.scala 160:64:@14851.4]
  wire [13:0] buffer_4_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68643; // @[Modules.scala 160:64:@14857.4]
  wire [13:0] _T_68644; // @[Modules.scala 160:64:@14858.4]
  wire [13:0] buffer_4_324; // @[Modules.scala 160:64:@14859.4]
  wire [13:0] buffer_4_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68649; // @[Modules.scala 160:64:@14865.4]
  wire [13:0] _T_68650; // @[Modules.scala 160:64:@14866.4]
  wire [13:0] buffer_4_326; // @[Modules.scala 160:64:@14867.4]
  wire [13:0] buffer_4_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68652; // @[Modules.scala 160:64:@14869.4]
  wire [13:0] _T_68653; // @[Modules.scala 160:64:@14870.4]
  wire [13:0] buffer_4_327; // @[Modules.scala 160:64:@14871.4]
  wire [13:0] buffer_4_56; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68655; // @[Modules.scala 160:64:@14873.4]
  wire [13:0] _T_68656; // @[Modules.scala 160:64:@14874.4]
  wire [13:0] buffer_4_328; // @[Modules.scala 160:64:@14875.4]
  wire [13:0] buffer_4_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68661; // @[Modules.scala 160:64:@14881.4]
  wire [13:0] _T_68662; // @[Modules.scala 160:64:@14882.4]
  wire [13:0] buffer_4_330; // @[Modules.scala 160:64:@14883.4]
  wire [13:0] buffer_4_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68664; // @[Modules.scala 160:64:@14885.4]
  wire [13:0] _T_68665; // @[Modules.scala 160:64:@14886.4]
  wire [13:0] buffer_4_331; // @[Modules.scala 160:64:@14887.4]
  wire [13:0] buffer_4_64; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68667; // @[Modules.scala 160:64:@14889.4]
  wire [13:0] _T_68668; // @[Modules.scala 160:64:@14890.4]
  wire [13:0] buffer_4_332; // @[Modules.scala 160:64:@14891.4]
  wire [14:0] _T_68670; // @[Modules.scala 160:64:@14893.4]
  wire [13:0] _T_68671; // @[Modules.scala 160:64:@14894.4]
  wire [13:0] buffer_4_333; // @[Modules.scala 160:64:@14895.4]
  wire [13:0] buffer_4_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68676; // @[Modules.scala 160:64:@14901.4]
  wire [13:0] _T_68677; // @[Modules.scala 160:64:@14902.4]
  wire [13:0] buffer_4_335; // @[Modules.scala 160:64:@14903.4]
  wire [13:0] buffer_4_72; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68679; // @[Modules.scala 160:64:@14905.4]
  wire [13:0] _T_68680; // @[Modules.scala 160:64:@14906.4]
  wire [13:0] buffer_4_336; // @[Modules.scala 160:64:@14907.4]
  wire [13:0] buffer_4_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68682; // @[Modules.scala 160:64:@14909.4]
  wire [13:0] _T_68683; // @[Modules.scala 160:64:@14910.4]
  wire [13:0] buffer_4_337; // @[Modules.scala 160:64:@14911.4]
  wire [13:0] buffer_4_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68688; // @[Modules.scala 160:64:@14917.4]
  wire [13:0] _T_68689; // @[Modules.scala 160:64:@14918.4]
  wire [13:0] buffer_4_339; // @[Modules.scala 160:64:@14919.4]
  wire [13:0] buffer_4_80; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68691; // @[Modules.scala 160:64:@14921.4]
  wire [13:0] _T_68692; // @[Modules.scala 160:64:@14922.4]
  wire [13:0] buffer_4_340; // @[Modules.scala 160:64:@14923.4]
  wire [13:0] buffer_4_82; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68694; // @[Modules.scala 160:64:@14925.4]
  wire [13:0] _T_68695; // @[Modules.scala 160:64:@14926.4]
  wire [13:0] buffer_4_341; // @[Modules.scala 160:64:@14927.4]
  wire [13:0] buffer_4_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68697; // @[Modules.scala 160:64:@14929.4]
  wire [13:0] _T_68698; // @[Modules.scala 160:64:@14930.4]
  wire [13:0] buffer_4_342; // @[Modules.scala 160:64:@14931.4]
  wire [13:0] buffer_4_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68706; // @[Modules.scala 160:64:@14941.4]
  wire [13:0] _T_68707; // @[Modules.scala 160:64:@14942.4]
  wire [13:0] buffer_4_345; // @[Modules.scala 160:64:@14943.4]
  wire [13:0] buffer_4_92; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68709; // @[Modules.scala 160:64:@14945.4]
  wire [13:0] _T_68710; // @[Modules.scala 160:64:@14946.4]
  wire [13:0] buffer_4_346; // @[Modules.scala 160:64:@14947.4]
  wire [13:0] buffer_4_94; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68712; // @[Modules.scala 160:64:@14949.4]
  wire [13:0] _T_68713; // @[Modules.scala 160:64:@14950.4]
  wire [13:0] buffer_4_347; // @[Modules.scala 160:64:@14951.4]
  wire [13:0] buffer_4_96; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68715; // @[Modules.scala 160:64:@14953.4]
  wire [13:0] _T_68716; // @[Modules.scala 160:64:@14954.4]
  wire [13:0] buffer_4_348; // @[Modules.scala 160:64:@14955.4]
  wire [13:0] buffer_4_101; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68721; // @[Modules.scala 160:64:@14961.4]
  wire [13:0] _T_68722; // @[Modules.scala 160:64:@14962.4]
  wire [13:0] buffer_4_350; // @[Modules.scala 160:64:@14963.4]
  wire [13:0] buffer_4_103; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68724; // @[Modules.scala 160:64:@14965.4]
  wire [13:0] _T_68725; // @[Modules.scala 160:64:@14966.4]
  wire [13:0] buffer_4_351; // @[Modules.scala 160:64:@14967.4]
  wire [13:0] buffer_4_104; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68727; // @[Modules.scala 160:64:@14969.4]
  wire [13:0] _T_68728; // @[Modules.scala 160:64:@14970.4]
  wire [13:0] buffer_4_352; // @[Modules.scala 160:64:@14971.4]
  wire [13:0] buffer_4_106; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68730; // @[Modules.scala 160:64:@14973.4]
  wire [13:0] _T_68731; // @[Modules.scala 160:64:@14974.4]
  wire [13:0] buffer_4_353; // @[Modules.scala 160:64:@14975.4]
  wire [14:0] _T_68733; // @[Modules.scala 160:64:@14977.4]
  wire [13:0] _T_68734; // @[Modules.scala 160:64:@14978.4]
  wire [13:0] buffer_4_354; // @[Modules.scala 160:64:@14979.4]
  wire [13:0] buffer_4_110; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68736; // @[Modules.scala 160:64:@14981.4]
  wire [13:0] _T_68737; // @[Modules.scala 160:64:@14982.4]
  wire [13:0] buffer_4_355; // @[Modules.scala 160:64:@14983.4]
  wire [13:0] buffer_4_112; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68739; // @[Modules.scala 160:64:@14985.4]
  wire [13:0] _T_68740; // @[Modules.scala 160:64:@14986.4]
  wire [13:0] buffer_4_356; // @[Modules.scala 160:64:@14987.4]
  wire [13:0] buffer_4_114; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68742; // @[Modules.scala 160:64:@14989.4]
  wire [13:0] _T_68743; // @[Modules.scala 160:64:@14990.4]
  wire [13:0] buffer_4_357; // @[Modules.scala 160:64:@14991.4]
  wire [13:0] buffer_4_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68745; // @[Modules.scala 160:64:@14993.4]
  wire [13:0] _T_68746; // @[Modules.scala 160:64:@14994.4]
  wire [13:0] buffer_4_358; // @[Modules.scala 160:64:@14995.4]
  wire [13:0] buffer_4_118; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_119; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68748; // @[Modules.scala 160:64:@14997.4]
  wire [13:0] _T_68749; // @[Modules.scala 160:64:@14998.4]
  wire [13:0] buffer_4_359; // @[Modules.scala 160:64:@14999.4]
  wire [13:0] buffer_4_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68751; // @[Modules.scala 160:64:@15001.4]
  wire [13:0] _T_68752; // @[Modules.scala 160:64:@15002.4]
  wire [13:0] buffer_4_360; // @[Modules.scala 160:64:@15003.4]
  wire [13:0] buffer_4_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68754; // @[Modules.scala 160:64:@15005.4]
  wire [13:0] _T_68755; // @[Modules.scala 160:64:@15006.4]
  wire [13:0] buffer_4_361; // @[Modules.scala 160:64:@15007.4]
  wire [13:0] buffer_4_124; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68757; // @[Modules.scala 160:64:@15009.4]
  wire [13:0] _T_68758; // @[Modules.scala 160:64:@15010.4]
  wire [13:0] buffer_4_362; // @[Modules.scala 160:64:@15011.4]
  wire [13:0] buffer_4_127; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68760; // @[Modules.scala 160:64:@15013.4]
  wire [13:0] _T_68761; // @[Modules.scala 160:64:@15014.4]
  wire [13:0] buffer_4_363; // @[Modules.scala 160:64:@15015.4]
  wire [13:0] buffer_4_129; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68763; // @[Modules.scala 160:64:@15017.4]
  wire [13:0] _T_68764; // @[Modules.scala 160:64:@15018.4]
  wire [13:0] buffer_4_364; // @[Modules.scala 160:64:@15019.4]
  wire [13:0] buffer_4_130; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68766; // @[Modules.scala 160:64:@15021.4]
  wire [13:0] _T_68767; // @[Modules.scala 160:64:@15022.4]
  wire [13:0] buffer_4_365; // @[Modules.scala 160:64:@15023.4]
  wire [13:0] buffer_4_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68769; // @[Modules.scala 160:64:@15025.4]
  wire [13:0] _T_68770; // @[Modules.scala 160:64:@15026.4]
  wire [13:0] buffer_4_366; // @[Modules.scala 160:64:@15027.4]
  wire [13:0] buffer_4_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68772; // @[Modules.scala 160:64:@15029.4]
  wire [13:0] _T_68773; // @[Modules.scala 160:64:@15030.4]
  wire [13:0] buffer_4_367; // @[Modules.scala 160:64:@15031.4]
  wire [13:0] buffer_4_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68775; // @[Modules.scala 160:64:@15033.4]
  wire [13:0] _T_68776; // @[Modules.scala 160:64:@15034.4]
  wire [13:0] buffer_4_368; // @[Modules.scala 160:64:@15035.4]
  wire [14:0] _T_68778; // @[Modules.scala 160:64:@15037.4]
  wire [13:0] _T_68779; // @[Modules.scala 160:64:@15038.4]
  wire [13:0] buffer_4_369; // @[Modules.scala 160:64:@15039.4]
  wire [13:0] buffer_4_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68781; // @[Modules.scala 160:64:@15041.4]
  wire [13:0] _T_68782; // @[Modules.scala 160:64:@15042.4]
  wire [13:0] buffer_4_370; // @[Modules.scala 160:64:@15043.4]
  wire [13:0] buffer_4_142; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68784; // @[Modules.scala 160:64:@15045.4]
  wire [13:0] _T_68785; // @[Modules.scala 160:64:@15046.4]
  wire [13:0] buffer_4_371; // @[Modules.scala 160:64:@15047.4]
  wire [13:0] buffer_4_144; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68787; // @[Modules.scala 160:64:@15049.4]
  wire [13:0] _T_68788; // @[Modules.scala 160:64:@15050.4]
  wire [13:0] buffer_4_372; // @[Modules.scala 160:64:@15051.4]
  wire [13:0] buffer_4_146; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68790; // @[Modules.scala 160:64:@15053.4]
  wire [13:0] _T_68791; // @[Modules.scala 160:64:@15054.4]
  wire [13:0] buffer_4_373; // @[Modules.scala 160:64:@15055.4]
  wire [13:0] buffer_4_148; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68793; // @[Modules.scala 160:64:@15057.4]
  wire [13:0] _T_68794; // @[Modules.scala 160:64:@15058.4]
  wire [13:0] buffer_4_374; // @[Modules.scala 160:64:@15059.4]
  wire [14:0] _T_68796; // @[Modules.scala 160:64:@15061.4]
  wire [13:0] _T_68797; // @[Modules.scala 160:64:@15062.4]
  wire [13:0] buffer_4_375; // @[Modules.scala 160:64:@15063.4]
  wire [13:0] buffer_4_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68799; // @[Modules.scala 160:64:@15065.4]
  wire [13:0] _T_68800; // @[Modules.scala 160:64:@15066.4]
  wire [13:0] buffer_4_376; // @[Modules.scala 160:64:@15067.4]
  wire [13:0] buffer_4_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68802; // @[Modules.scala 160:64:@15069.4]
  wire [13:0] _T_68803; // @[Modules.scala 160:64:@15070.4]
  wire [13:0] buffer_4_377; // @[Modules.scala 160:64:@15071.4]
  wire [14:0] _T_68805; // @[Modules.scala 160:64:@15073.4]
  wire [13:0] _T_68806; // @[Modules.scala 160:64:@15074.4]
  wire [13:0] buffer_4_378; // @[Modules.scala 160:64:@15075.4]
  wire [13:0] buffer_4_158; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68808; // @[Modules.scala 160:64:@15077.4]
  wire [13:0] _T_68809; // @[Modules.scala 160:64:@15078.4]
  wire [13:0] buffer_4_379; // @[Modules.scala 160:64:@15079.4]
  wire [13:0] buffer_4_160; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68811; // @[Modules.scala 160:64:@15081.4]
  wire [13:0] _T_68812; // @[Modules.scala 160:64:@15082.4]
  wire [13:0] buffer_4_380; // @[Modules.scala 160:64:@15083.4]
  wire [13:0] buffer_4_162; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_163; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68814; // @[Modules.scala 160:64:@15085.4]
  wire [13:0] _T_68815; // @[Modules.scala 160:64:@15086.4]
  wire [13:0] buffer_4_381; // @[Modules.scala 160:64:@15087.4]
  wire [13:0] buffer_4_164; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68817; // @[Modules.scala 160:64:@15089.4]
  wire [13:0] _T_68818; // @[Modules.scala 160:64:@15090.4]
  wire [13:0] buffer_4_382; // @[Modules.scala 160:64:@15091.4]
  wire [13:0] buffer_4_166; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68820; // @[Modules.scala 160:64:@15093.4]
  wire [13:0] _T_68821; // @[Modules.scala 160:64:@15094.4]
  wire [13:0] buffer_4_383; // @[Modules.scala 160:64:@15095.4]
  wire [13:0] buffer_4_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68823; // @[Modules.scala 160:64:@15097.4]
  wire [13:0] _T_68824; // @[Modules.scala 160:64:@15098.4]
  wire [13:0] buffer_4_384; // @[Modules.scala 160:64:@15099.4]
  wire [13:0] buffer_4_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68826; // @[Modules.scala 160:64:@15101.4]
  wire [13:0] _T_68827; // @[Modules.scala 160:64:@15102.4]
  wire [13:0] buffer_4_385; // @[Modules.scala 160:64:@15103.4]
  wire [13:0] buffer_4_172; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_173; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68829; // @[Modules.scala 160:64:@15105.4]
  wire [13:0] _T_68830; // @[Modules.scala 160:64:@15106.4]
  wire [13:0] buffer_4_386; // @[Modules.scala 160:64:@15107.4]
  wire [13:0] buffer_4_174; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68832; // @[Modules.scala 160:64:@15109.4]
  wire [13:0] _T_68833; // @[Modules.scala 160:64:@15110.4]
  wire [13:0] buffer_4_387; // @[Modules.scala 160:64:@15111.4]
  wire [14:0] _T_68838; // @[Modules.scala 160:64:@15117.4]
  wire [13:0] _T_68839; // @[Modules.scala 160:64:@15118.4]
  wire [13:0] buffer_4_389; // @[Modules.scala 160:64:@15119.4]
  wire [13:0] buffer_4_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68841; // @[Modules.scala 160:64:@15121.4]
  wire [13:0] _T_68842; // @[Modules.scala 160:64:@15122.4]
  wire [13:0] buffer_4_390; // @[Modules.scala 160:64:@15123.4]
  wire [13:0] buffer_4_182; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68844; // @[Modules.scala 160:64:@15125.4]
  wire [13:0] _T_68845; // @[Modules.scala 160:64:@15126.4]
  wire [13:0] buffer_4_391; // @[Modules.scala 160:64:@15127.4]
  wire [13:0] buffer_4_184; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68847; // @[Modules.scala 160:64:@15129.4]
  wire [13:0] _T_68848; // @[Modules.scala 160:64:@15130.4]
  wire [13:0] buffer_4_392; // @[Modules.scala 160:64:@15131.4]
  wire [13:0] buffer_4_188; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68853; // @[Modules.scala 160:64:@15137.4]
  wire [13:0] _T_68854; // @[Modules.scala 160:64:@15138.4]
  wire [13:0] buffer_4_394; // @[Modules.scala 160:64:@15139.4]
  wire [13:0] buffer_4_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68856; // @[Modules.scala 160:64:@15141.4]
  wire [13:0] _T_68857; // @[Modules.scala 160:64:@15142.4]
  wire [13:0] buffer_4_395; // @[Modules.scala 160:64:@15143.4]
  wire [13:0] buffer_4_192; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68859; // @[Modules.scala 160:64:@15145.4]
  wire [13:0] _T_68860; // @[Modules.scala 160:64:@15146.4]
  wire [13:0] buffer_4_396; // @[Modules.scala 160:64:@15147.4]
  wire [13:0] buffer_4_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68862; // @[Modules.scala 160:64:@15149.4]
  wire [13:0] _T_68863; // @[Modules.scala 160:64:@15150.4]
  wire [13:0] buffer_4_397; // @[Modules.scala 160:64:@15151.4]
  wire [13:0] buffer_4_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68868; // @[Modules.scala 160:64:@15157.4]
  wire [13:0] _T_68869; // @[Modules.scala 160:64:@15158.4]
  wire [13:0] buffer_4_399; // @[Modules.scala 160:64:@15159.4]
  wire [14:0] _T_68871; // @[Modules.scala 160:64:@15161.4]
  wire [13:0] _T_68872; // @[Modules.scala 160:64:@15162.4]
  wire [13:0] buffer_4_400; // @[Modules.scala 160:64:@15163.4]
  wire [13:0] buffer_4_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68874; // @[Modules.scala 160:64:@15165.4]
  wire [13:0] _T_68875; // @[Modules.scala 160:64:@15166.4]
  wire [13:0] buffer_4_401; // @[Modules.scala 160:64:@15167.4]
  wire [13:0] buffer_4_204; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68877; // @[Modules.scala 160:64:@15169.4]
  wire [13:0] _T_68878; // @[Modules.scala 160:64:@15170.4]
  wire [13:0] buffer_4_402; // @[Modules.scala 160:64:@15171.4]
  wire [13:0] buffer_4_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68880; // @[Modules.scala 160:64:@15173.4]
  wire [13:0] _T_68881; // @[Modules.scala 160:64:@15174.4]
  wire [13:0] buffer_4_403; // @[Modules.scala 160:64:@15175.4]
  wire [13:0] buffer_4_209; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68883; // @[Modules.scala 160:64:@15177.4]
  wire [13:0] _T_68884; // @[Modules.scala 160:64:@15178.4]
  wire [13:0] buffer_4_404; // @[Modules.scala 160:64:@15179.4]
  wire [13:0] buffer_4_210; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68886; // @[Modules.scala 160:64:@15181.4]
  wire [13:0] _T_68887; // @[Modules.scala 160:64:@15182.4]
  wire [13:0] buffer_4_405; // @[Modules.scala 160:64:@15183.4]
  wire [13:0] buffer_4_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68895; // @[Modules.scala 160:64:@15193.4]
  wire [13:0] _T_68896; // @[Modules.scala 160:64:@15194.4]
  wire [13:0] buffer_4_408; // @[Modules.scala 160:64:@15195.4]
  wire [13:0] buffer_4_218; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68898; // @[Modules.scala 160:64:@15197.4]
  wire [13:0] _T_68899; // @[Modules.scala 160:64:@15198.4]
  wire [13:0] buffer_4_409; // @[Modules.scala 160:64:@15199.4]
  wire [13:0] buffer_4_220; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_221; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68901; // @[Modules.scala 160:64:@15201.4]
  wire [13:0] _T_68902; // @[Modules.scala 160:64:@15202.4]
  wire [13:0] buffer_4_410; // @[Modules.scala 160:64:@15203.4]
  wire [13:0] buffer_4_222; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68904; // @[Modules.scala 160:64:@15205.4]
  wire [13:0] _T_68905; // @[Modules.scala 160:64:@15206.4]
  wire [13:0] buffer_4_411; // @[Modules.scala 160:64:@15207.4]
  wire [13:0] buffer_4_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68910; // @[Modules.scala 160:64:@15213.4]
  wire [13:0] _T_68911; // @[Modules.scala 160:64:@15214.4]
  wire [13:0] buffer_4_413; // @[Modules.scala 160:64:@15215.4]
  wire [13:0] buffer_4_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68913; // @[Modules.scala 160:64:@15217.4]
  wire [13:0] _T_68914; // @[Modules.scala 160:64:@15218.4]
  wire [13:0] buffer_4_414; // @[Modules.scala 160:64:@15219.4]
  wire [13:0] buffer_4_230; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68916; // @[Modules.scala 160:64:@15221.4]
  wire [13:0] _T_68917; // @[Modules.scala 160:64:@15222.4]
  wire [13:0] buffer_4_415; // @[Modules.scala 160:64:@15223.4]
  wire [13:0] buffer_4_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68919; // @[Modules.scala 160:64:@15225.4]
  wire [13:0] _T_68920; // @[Modules.scala 160:64:@15226.4]
  wire [13:0] buffer_4_416; // @[Modules.scala 160:64:@15227.4]
  wire [13:0] buffer_4_234; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68922; // @[Modules.scala 160:64:@15229.4]
  wire [13:0] _T_68923; // @[Modules.scala 160:64:@15230.4]
  wire [13:0] buffer_4_417; // @[Modules.scala 160:64:@15231.4]
  wire [13:0] buffer_4_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68928; // @[Modules.scala 160:64:@15237.4]
  wire [13:0] _T_68929; // @[Modules.scala 160:64:@15238.4]
  wire [13:0] buffer_4_419; // @[Modules.scala 160:64:@15239.4]
  wire [14:0] _T_68931; // @[Modules.scala 160:64:@15241.4]
  wire [13:0] _T_68932; // @[Modules.scala 160:64:@15242.4]
  wire [13:0] buffer_4_420; // @[Modules.scala 160:64:@15243.4]
  wire [13:0] buffer_4_242; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68934; // @[Modules.scala 160:64:@15245.4]
  wire [13:0] _T_68935; // @[Modules.scala 160:64:@15246.4]
  wire [13:0] buffer_4_421; // @[Modules.scala 160:64:@15247.4]
  wire [13:0] buffer_4_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68937; // @[Modules.scala 160:64:@15249.4]
  wire [13:0] _T_68938; // @[Modules.scala 160:64:@15250.4]
  wire [13:0] buffer_4_422; // @[Modules.scala 160:64:@15251.4]
  wire [13:0] buffer_4_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68940; // @[Modules.scala 160:64:@15253.4]
  wire [13:0] _T_68941; // @[Modules.scala 160:64:@15254.4]
  wire [13:0] buffer_4_423; // @[Modules.scala 160:64:@15255.4]
  wire [13:0] buffer_4_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68943; // @[Modules.scala 160:64:@15257.4]
  wire [13:0] _T_68944; // @[Modules.scala 160:64:@15258.4]
  wire [13:0] buffer_4_424; // @[Modules.scala 160:64:@15259.4]
  wire [13:0] buffer_4_252; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68949; // @[Modules.scala 160:64:@15265.4]
  wire [13:0] _T_68950; // @[Modules.scala 160:64:@15266.4]
  wire [13:0] buffer_4_426; // @[Modules.scala 160:64:@15267.4]
  wire [13:0] buffer_4_254; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68952; // @[Modules.scala 160:64:@15269.4]
  wire [13:0] _T_68953; // @[Modules.scala 160:64:@15270.4]
  wire [13:0] buffer_4_427; // @[Modules.scala 160:64:@15271.4]
  wire [13:0] buffer_4_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68955; // @[Modules.scala 160:64:@15273.4]
  wire [13:0] _T_68956; // @[Modules.scala 160:64:@15274.4]
  wire [13:0] buffer_4_428; // @[Modules.scala 160:64:@15275.4]
  wire [13:0] buffer_4_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68958; // @[Modules.scala 160:64:@15277.4]
  wire [13:0] _T_68959; // @[Modules.scala 160:64:@15278.4]
  wire [13:0] buffer_4_429; // @[Modules.scala 160:64:@15279.4]
  wire [13:0] buffer_4_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68961; // @[Modules.scala 160:64:@15281.4]
  wire [13:0] _T_68962; // @[Modules.scala 160:64:@15282.4]
  wire [13:0] buffer_4_430; // @[Modules.scala 160:64:@15283.4]
  wire [13:0] buffer_4_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68964; // @[Modules.scala 160:64:@15285.4]
  wire [13:0] _T_68965; // @[Modules.scala 160:64:@15286.4]
  wire [13:0] buffer_4_431; // @[Modules.scala 160:64:@15287.4]
  wire [13:0] buffer_4_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68967; // @[Modules.scala 160:64:@15289.4]
  wire [13:0] _T_68968; // @[Modules.scala 160:64:@15290.4]
  wire [13:0] buffer_4_432; // @[Modules.scala 160:64:@15291.4]
  wire [13:0] buffer_4_266; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_267; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68970; // @[Modules.scala 160:64:@15293.4]
  wire [13:0] _T_68971; // @[Modules.scala 160:64:@15294.4]
  wire [13:0] buffer_4_433; // @[Modules.scala 160:64:@15295.4]
  wire [13:0] buffer_4_268; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68973; // @[Modules.scala 160:64:@15297.4]
  wire [13:0] _T_68974; // @[Modules.scala 160:64:@15298.4]
  wire [13:0] buffer_4_434; // @[Modules.scala 160:64:@15299.4]
  wire [14:0] _T_68976; // @[Modules.scala 160:64:@15301.4]
  wire [13:0] _T_68977; // @[Modules.scala 160:64:@15302.4]
  wire [13:0] buffer_4_435; // @[Modules.scala 160:64:@15303.4]
  wire [14:0] _T_68979; // @[Modules.scala 160:64:@15305.4]
  wire [13:0] _T_68980; // @[Modules.scala 160:64:@15306.4]
  wire [13:0] buffer_4_436; // @[Modules.scala 160:64:@15307.4]
  wire [14:0] _T_68982; // @[Modules.scala 160:64:@15309.4]
  wire [13:0] _T_68983; // @[Modules.scala 160:64:@15310.4]
  wire [13:0] buffer_4_437; // @[Modules.scala 160:64:@15311.4]
  wire [13:0] buffer_4_278; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68988; // @[Modules.scala 160:64:@15317.4]
  wire [13:0] _T_68989; // @[Modules.scala 160:64:@15318.4]
  wire [13:0] buffer_4_439; // @[Modules.scala 160:64:@15319.4]
  wire [13:0] buffer_4_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68991; // @[Modules.scala 160:64:@15321.4]
  wire [13:0] _T_68992; // @[Modules.scala 160:64:@15322.4]
  wire [13:0] buffer_4_440; // @[Modules.scala 160:64:@15323.4]
  wire [13:0] buffer_4_282; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68994; // @[Modules.scala 160:64:@15325.4]
  wire [13:0] _T_68995; // @[Modules.scala 160:64:@15326.4]
  wire [13:0] buffer_4_441; // @[Modules.scala 160:64:@15327.4]
  wire [13:0] buffer_4_284; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_285; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_68997; // @[Modules.scala 160:64:@15329.4]
  wire [13:0] _T_68998; // @[Modules.scala 160:64:@15330.4]
  wire [13:0] buffer_4_442; // @[Modules.scala 160:64:@15331.4]
  wire [13:0] buffer_4_286; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_287; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_69000; // @[Modules.scala 160:64:@15333.4]
  wire [13:0] _T_69001; // @[Modules.scala 160:64:@15334.4]
  wire [13:0] buffer_4_443; // @[Modules.scala 160:64:@15335.4]
  wire [13:0] buffer_4_288; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_4_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_69003; // @[Modules.scala 160:64:@15337.4]
  wire [13:0] _T_69004; // @[Modules.scala 160:64:@15338.4]
  wire [13:0] buffer_4_444; // @[Modules.scala 160:64:@15339.4]
  wire [14:0] _T_69006; // @[Modules.scala 160:64:@15341.4]
  wire [13:0] _T_69007; // @[Modules.scala 160:64:@15342.4]
  wire [13:0] buffer_4_445; // @[Modules.scala 160:64:@15343.4]
  wire [13:0] buffer_4_292; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_69009; // @[Modules.scala 160:64:@15345.4]
  wire [13:0] _T_69010; // @[Modules.scala 160:64:@15346.4]
  wire [13:0] buffer_4_446; // @[Modules.scala 160:64:@15347.4]
  wire [13:0] buffer_4_296; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_69015; // @[Modules.scala 160:64:@15353.4]
  wire [13:0] _T_69016; // @[Modules.scala 160:64:@15354.4]
  wire [13:0] buffer_4_448; // @[Modules.scala 160:64:@15355.4]
  wire [14:0] _T_69021; // @[Modules.scala 160:64:@15361.4]
  wire [13:0] _T_69022; // @[Modules.scala 160:64:@15362.4]
  wire [13:0] buffer_4_450; // @[Modules.scala 160:64:@15363.4]
  wire [14:0] _T_69024; // @[Modules.scala 160:64:@15365.4]
  wire [13:0] _T_69025; // @[Modules.scala 160:64:@15366.4]
  wire [13:0] buffer_4_451; // @[Modules.scala 160:64:@15367.4]
  wire [14:0] _T_69027; // @[Modules.scala 160:64:@15369.4]
  wire [13:0] _T_69028; // @[Modules.scala 160:64:@15370.4]
  wire [13:0] buffer_4_452; // @[Modules.scala 160:64:@15371.4]
  wire [14:0] _T_69030; // @[Modules.scala 160:64:@15373.4]
  wire [13:0] _T_69031; // @[Modules.scala 160:64:@15374.4]
  wire [13:0] buffer_4_453; // @[Modules.scala 160:64:@15375.4]
  wire [14:0] _T_69033; // @[Modules.scala 160:64:@15377.4]
  wire [13:0] _T_69034; // @[Modules.scala 160:64:@15378.4]
  wire [13:0] buffer_4_454; // @[Modules.scala 160:64:@15379.4]
  wire [14:0] _T_69036; // @[Modules.scala 160:64:@15381.4]
  wire [13:0] _T_69037; // @[Modules.scala 160:64:@15382.4]
  wire [13:0] buffer_4_455; // @[Modules.scala 160:64:@15383.4]
  wire [14:0] _T_69039; // @[Modules.scala 160:64:@15385.4]
  wire [13:0] _T_69040; // @[Modules.scala 160:64:@15386.4]
  wire [13:0] buffer_4_456; // @[Modules.scala 160:64:@15387.4]
  wire [14:0] _T_69042; // @[Modules.scala 160:64:@15389.4]
  wire [13:0] _T_69043; // @[Modules.scala 160:64:@15390.4]
  wire [13:0] buffer_4_457; // @[Modules.scala 160:64:@15391.4]
  wire [14:0] _T_69045; // @[Modules.scala 160:64:@15393.4]
  wire [13:0] _T_69046; // @[Modules.scala 160:64:@15394.4]
  wire [13:0] buffer_4_458; // @[Modules.scala 160:64:@15395.4]
  wire [14:0] _T_69048; // @[Modules.scala 160:64:@15397.4]
  wire [13:0] _T_69049; // @[Modules.scala 160:64:@15398.4]
  wire [13:0] buffer_4_459; // @[Modules.scala 160:64:@15399.4]
  wire [14:0] _T_69051; // @[Modules.scala 160:64:@15401.4]
  wire [13:0] _T_69052; // @[Modules.scala 160:64:@15402.4]
  wire [13:0] buffer_4_460; // @[Modules.scala 160:64:@15403.4]
  wire [14:0] _T_69054; // @[Modules.scala 160:64:@15405.4]
  wire [13:0] _T_69055; // @[Modules.scala 160:64:@15406.4]
  wire [13:0] buffer_4_461; // @[Modules.scala 160:64:@15407.4]
  wire [14:0] _T_69057; // @[Modules.scala 160:64:@15409.4]
  wire [13:0] _T_69058; // @[Modules.scala 160:64:@15410.4]
  wire [13:0] buffer_4_462; // @[Modules.scala 160:64:@15411.4]
  wire [14:0] _T_69060; // @[Modules.scala 160:64:@15413.4]
  wire [13:0] _T_69061; // @[Modules.scala 160:64:@15414.4]
  wire [13:0] buffer_4_463; // @[Modules.scala 160:64:@15415.4]
  wire [14:0] _T_69063; // @[Modules.scala 160:64:@15417.4]
  wire [13:0] _T_69064; // @[Modules.scala 160:64:@15418.4]
  wire [13:0] buffer_4_464; // @[Modules.scala 160:64:@15419.4]
  wire [14:0] _T_69066; // @[Modules.scala 160:64:@15421.4]
  wire [13:0] _T_69067; // @[Modules.scala 160:64:@15422.4]
  wire [13:0] buffer_4_465; // @[Modules.scala 160:64:@15423.4]
  wire [14:0] _T_69069; // @[Modules.scala 160:64:@15425.4]
  wire [13:0] _T_69070; // @[Modules.scala 160:64:@15426.4]
  wire [13:0] buffer_4_466; // @[Modules.scala 160:64:@15427.4]
  wire [14:0] _T_69072; // @[Modules.scala 160:64:@15429.4]
  wire [13:0] _T_69073; // @[Modules.scala 160:64:@15430.4]
  wire [13:0] buffer_4_467; // @[Modules.scala 160:64:@15431.4]
  wire [14:0] _T_69075; // @[Modules.scala 160:64:@15433.4]
  wire [13:0] _T_69076; // @[Modules.scala 160:64:@15434.4]
  wire [13:0] buffer_4_468; // @[Modules.scala 160:64:@15435.4]
  wire [14:0] _T_69078; // @[Modules.scala 160:64:@15437.4]
  wire [13:0] _T_69079; // @[Modules.scala 160:64:@15438.4]
  wire [13:0] buffer_4_469; // @[Modules.scala 160:64:@15439.4]
  wire [14:0] _T_69081; // @[Modules.scala 160:64:@15441.4]
  wire [13:0] _T_69082; // @[Modules.scala 160:64:@15442.4]
  wire [13:0] buffer_4_470; // @[Modules.scala 160:64:@15443.4]
  wire [14:0] _T_69084; // @[Modules.scala 160:64:@15445.4]
  wire [13:0] _T_69085; // @[Modules.scala 160:64:@15446.4]
  wire [13:0] buffer_4_471; // @[Modules.scala 160:64:@15447.4]
  wire [14:0] _T_69087; // @[Modules.scala 160:64:@15449.4]
  wire [13:0] _T_69088; // @[Modules.scala 160:64:@15450.4]
  wire [13:0] buffer_4_472; // @[Modules.scala 160:64:@15451.4]
  wire [14:0] _T_69090; // @[Modules.scala 160:64:@15453.4]
  wire [13:0] _T_69091; // @[Modules.scala 160:64:@15454.4]
  wire [13:0] buffer_4_473; // @[Modules.scala 160:64:@15455.4]
  wire [14:0] _T_69093; // @[Modules.scala 160:64:@15457.4]
  wire [13:0] _T_69094; // @[Modules.scala 160:64:@15458.4]
  wire [13:0] buffer_4_474; // @[Modules.scala 160:64:@15459.4]
  wire [14:0] _T_69096; // @[Modules.scala 160:64:@15461.4]
  wire [13:0] _T_69097; // @[Modules.scala 160:64:@15462.4]
  wire [13:0] buffer_4_475; // @[Modules.scala 160:64:@15463.4]
  wire [14:0] _T_69099; // @[Modules.scala 160:64:@15465.4]
  wire [13:0] _T_69100; // @[Modules.scala 160:64:@15466.4]
  wire [13:0] buffer_4_476; // @[Modules.scala 160:64:@15467.4]
  wire [14:0] _T_69102; // @[Modules.scala 160:64:@15469.4]
  wire [13:0] _T_69103; // @[Modules.scala 160:64:@15470.4]
  wire [13:0] buffer_4_477; // @[Modules.scala 160:64:@15471.4]
  wire [14:0] _T_69105; // @[Modules.scala 160:64:@15473.4]
  wire [13:0] _T_69106; // @[Modules.scala 160:64:@15474.4]
  wire [13:0] buffer_4_478; // @[Modules.scala 160:64:@15475.4]
  wire [14:0] _T_69108; // @[Modules.scala 160:64:@15477.4]
  wire [13:0] _T_69109; // @[Modules.scala 160:64:@15478.4]
  wire [13:0] buffer_4_479; // @[Modules.scala 160:64:@15479.4]
  wire [14:0] _T_69111; // @[Modules.scala 160:64:@15481.4]
  wire [13:0] _T_69112; // @[Modules.scala 160:64:@15482.4]
  wire [13:0] buffer_4_480; // @[Modules.scala 160:64:@15483.4]
  wire [14:0] _T_69114; // @[Modules.scala 160:64:@15485.4]
  wire [13:0] _T_69115; // @[Modules.scala 160:64:@15486.4]
  wire [13:0] buffer_4_481; // @[Modules.scala 160:64:@15487.4]
  wire [14:0] _T_69117; // @[Modules.scala 160:64:@15489.4]
  wire [13:0] _T_69118; // @[Modules.scala 160:64:@15490.4]
  wire [13:0] buffer_4_482; // @[Modules.scala 160:64:@15491.4]
  wire [14:0] _T_69120; // @[Modules.scala 160:64:@15493.4]
  wire [13:0] _T_69121; // @[Modules.scala 160:64:@15494.4]
  wire [13:0] buffer_4_483; // @[Modules.scala 160:64:@15495.4]
  wire [14:0] _T_69123; // @[Modules.scala 160:64:@15497.4]
  wire [13:0] _T_69124; // @[Modules.scala 160:64:@15498.4]
  wire [13:0] buffer_4_484; // @[Modules.scala 160:64:@15499.4]
  wire [14:0] _T_69126; // @[Modules.scala 160:64:@15501.4]
  wire [13:0] _T_69127; // @[Modules.scala 160:64:@15502.4]
  wire [13:0] buffer_4_485; // @[Modules.scala 160:64:@15503.4]
  wire [14:0] _T_69129; // @[Modules.scala 160:64:@15505.4]
  wire [13:0] _T_69130; // @[Modules.scala 160:64:@15506.4]
  wire [13:0] buffer_4_486; // @[Modules.scala 160:64:@15507.4]
  wire [14:0] _T_69132; // @[Modules.scala 160:64:@15509.4]
  wire [13:0] _T_69133; // @[Modules.scala 160:64:@15510.4]
  wire [13:0] buffer_4_487; // @[Modules.scala 160:64:@15511.4]
  wire [14:0] _T_69135; // @[Modules.scala 160:64:@15513.4]
  wire [13:0] _T_69136; // @[Modules.scala 160:64:@15514.4]
  wire [13:0] buffer_4_488; // @[Modules.scala 160:64:@15515.4]
  wire [14:0] _T_69138; // @[Modules.scala 160:64:@15517.4]
  wire [13:0] _T_69139; // @[Modules.scala 160:64:@15518.4]
  wire [13:0] buffer_4_489; // @[Modules.scala 160:64:@15519.4]
  wire [14:0] _T_69141; // @[Modules.scala 160:64:@15521.4]
  wire [13:0] _T_69142; // @[Modules.scala 160:64:@15522.4]
  wire [13:0] buffer_4_490; // @[Modules.scala 160:64:@15523.4]
  wire [14:0] _T_69144; // @[Modules.scala 160:64:@15525.4]
  wire [13:0] _T_69145; // @[Modules.scala 160:64:@15526.4]
  wire [13:0] buffer_4_491; // @[Modules.scala 160:64:@15527.4]
  wire [14:0] _T_69147; // @[Modules.scala 160:64:@15529.4]
  wire [13:0] _T_69148; // @[Modules.scala 160:64:@15530.4]
  wire [13:0] buffer_4_492; // @[Modules.scala 160:64:@15531.4]
  wire [14:0] _T_69150; // @[Modules.scala 160:64:@15533.4]
  wire [13:0] _T_69151; // @[Modules.scala 160:64:@15534.4]
  wire [13:0] buffer_4_493; // @[Modules.scala 160:64:@15535.4]
  wire [14:0] _T_69153; // @[Modules.scala 160:64:@15537.4]
  wire [13:0] _T_69154; // @[Modules.scala 160:64:@15538.4]
  wire [13:0] buffer_4_494; // @[Modules.scala 160:64:@15539.4]
  wire [14:0] _T_69156; // @[Modules.scala 160:64:@15541.4]
  wire [13:0] _T_69157; // @[Modules.scala 160:64:@15542.4]
  wire [13:0] buffer_4_495; // @[Modules.scala 160:64:@15543.4]
  wire [14:0] _T_69159; // @[Modules.scala 160:64:@15545.4]
  wire [13:0] _T_69160; // @[Modules.scala 160:64:@15546.4]
  wire [13:0] buffer_4_496; // @[Modules.scala 160:64:@15547.4]
  wire [14:0] _T_69162; // @[Modules.scala 160:64:@15549.4]
  wire [13:0] _T_69163; // @[Modules.scala 160:64:@15550.4]
  wire [13:0] buffer_4_497; // @[Modules.scala 160:64:@15551.4]
  wire [14:0] _T_69165; // @[Modules.scala 160:64:@15553.4]
  wire [13:0] _T_69166; // @[Modules.scala 160:64:@15554.4]
  wire [13:0] buffer_4_498; // @[Modules.scala 160:64:@15555.4]
  wire [14:0] _T_69168; // @[Modules.scala 160:64:@15557.4]
  wire [13:0] _T_69169; // @[Modules.scala 160:64:@15558.4]
  wire [13:0] buffer_4_499; // @[Modules.scala 160:64:@15559.4]
  wire [14:0] _T_69171; // @[Modules.scala 160:64:@15561.4]
  wire [13:0] _T_69172; // @[Modules.scala 160:64:@15562.4]
  wire [13:0] buffer_4_500; // @[Modules.scala 160:64:@15563.4]
  wire [14:0] _T_69174; // @[Modules.scala 160:64:@15565.4]
  wire [13:0] _T_69175; // @[Modules.scala 160:64:@15566.4]
  wire [13:0] buffer_4_501; // @[Modules.scala 160:64:@15567.4]
  wire [14:0] _T_69177; // @[Modules.scala 160:64:@15569.4]
  wire [13:0] _T_69178; // @[Modules.scala 160:64:@15570.4]
  wire [13:0] buffer_4_502; // @[Modules.scala 160:64:@15571.4]
  wire [14:0] _T_69183; // @[Modules.scala 160:64:@15577.4]
  wire [13:0] _T_69184; // @[Modules.scala 160:64:@15578.4]
  wire [13:0] buffer_4_504; // @[Modules.scala 160:64:@15579.4]
  wire [14:0] _T_69186; // @[Modules.scala 160:64:@15581.4]
  wire [13:0] _T_69187; // @[Modules.scala 160:64:@15582.4]
  wire [13:0] buffer_4_505; // @[Modules.scala 160:64:@15583.4]
  wire [14:0] _T_69189; // @[Modules.scala 160:64:@15585.4]
  wire [13:0] _T_69190; // @[Modules.scala 160:64:@15586.4]
  wire [13:0] buffer_4_506; // @[Modules.scala 160:64:@15587.4]
  wire [14:0] _T_69192; // @[Modules.scala 160:64:@15589.4]
  wire [13:0] _T_69193; // @[Modules.scala 160:64:@15590.4]
  wire [13:0] buffer_4_507; // @[Modules.scala 160:64:@15591.4]
  wire [14:0] _T_69195; // @[Modules.scala 160:64:@15593.4]
  wire [13:0] _T_69196; // @[Modules.scala 160:64:@15594.4]
  wire [13:0] buffer_4_508; // @[Modules.scala 160:64:@15595.4]
  wire [14:0] _T_69198; // @[Modules.scala 160:64:@15597.4]
  wire [13:0] _T_69199; // @[Modules.scala 160:64:@15598.4]
  wire [13:0] buffer_4_509; // @[Modules.scala 160:64:@15599.4]
  wire [14:0] _T_69201; // @[Modules.scala 160:64:@15601.4]
  wire [13:0] _T_69202; // @[Modules.scala 160:64:@15602.4]
  wire [13:0] buffer_4_510; // @[Modules.scala 160:64:@15603.4]
  wire [14:0] _T_69204; // @[Modules.scala 160:64:@15605.4]
  wire [13:0] _T_69205; // @[Modules.scala 160:64:@15606.4]
  wire [13:0] buffer_4_511; // @[Modules.scala 160:64:@15607.4]
  wire [14:0] _T_69207; // @[Modules.scala 160:64:@15609.4]
  wire [13:0] _T_69208; // @[Modules.scala 160:64:@15610.4]
  wire [13:0] buffer_4_512; // @[Modules.scala 160:64:@15611.4]
  wire [14:0] _T_69210; // @[Modules.scala 160:64:@15613.4]
  wire [13:0] _T_69211; // @[Modules.scala 160:64:@15614.4]
  wire [13:0] buffer_4_513; // @[Modules.scala 160:64:@15615.4]
  wire [14:0] _T_69213; // @[Modules.scala 160:64:@15617.4]
  wire [13:0] _T_69214; // @[Modules.scala 160:64:@15618.4]
  wire [13:0] buffer_4_514; // @[Modules.scala 160:64:@15619.4]
  wire [14:0] _T_69216; // @[Modules.scala 160:64:@15621.4]
  wire [13:0] _T_69217; // @[Modules.scala 160:64:@15622.4]
  wire [13:0] buffer_4_515; // @[Modules.scala 160:64:@15623.4]
  wire [14:0] _T_69219; // @[Modules.scala 160:64:@15625.4]
  wire [13:0] _T_69220; // @[Modules.scala 160:64:@15626.4]
  wire [13:0] buffer_4_516; // @[Modules.scala 160:64:@15627.4]
  wire [14:0] _T_69222; // @[Modules.scala 160:64:@15629.4]
  wire [13:0] _T_69223; // @[Modules.scala 160:64:@15630.4]
  wire [13:0] buffer_4_517; // @[Modules.scala 160:64:@15631.4]
  wire [14:0] _T_69225; // @[Modules.scala 160:64:@15633.4]
  wire [13:0] _T_69226; // @[Modules.scala 160:64:@15634.4]
  wire [13:0] buffer_4_518; // @[Modules.scala 160:64:@15635.4]
  wire [14:0] _T_69228; // @[Modules.scala 160:64:@15637.4]
  wire [13:0] _T_69229; // @[Modules.scala 160:64:@15638.4]
  wire [13:0] buffer_4_519; // @[Modules.scala 160:64:@15639.4]
  wire [14:0] _T_69231; // @[Modules.scala 160:64:@15641.4]
  wire [13:0] _T_69232; // @[Modules.scala 160:64:@15642.4]
  wire [13:0] buffer_4_520; // @[Modules.scala 160:64:@15643.4]
  wire [14:0] _T_69234; // @[Modules.scala 160:64:@15645.4]
  wire [13:0] _T_69235; // @[Modules.scala 160:64:@15646.4]
  wire [13:0] buffer_4_521; // @[Modules.scala 160:64:@15647.4]
  wire [14:0] _T_69237; // @[Modules.scala 160:64:@15649.4]
  wire [13:0] _T_69238; // @[Modules.scala 160:64:@15650.4]
  wire [13:0] buffer_4_522; // @[Modules.scala 160:64:@15651.4]
  wire [14:0] _T_69240; // @[Modules.scala 160:64:@15653.4]
  wire [13:0] _T_69241; // @[Modules.scala 160:64:@15654.4]
  wire [13:0] buffer_4_523; // @[Modules.scala 160:64:@15655.4]
  wire [14:0] _T_69243; // @[Modules.scala 160:64:@15657.4]
  wire [13:0] _T_69244; // @[Modules.scala 160:64:@15658.4]
  wire [13:0] buffer_4_524; // @[Modules.scala 160:64:@15659.4]
  wire [14:0] _T_69246; // @[Modules.scala 166:64:@15661.4]
  wire [13:0] _T_69247; // @[Modules.scala 166:64:@15662.4]
  wire [13:0] buffer_4_525; // @[Modules.scala 166:64:@15663.4]
  wire [14:0] _T_69249; // @[Modules.scala 166:64:@15665.4]
  wire [13:0] _T_69250; // @[Modules.scala 166:64:@15666.4]
  wire [13:0] buffer_4_526; // @[Modules.scala 166:64:@15667.4]
  wire [14:0] _T_69252; // @[Modules.scala 166:64:@15669.4]
  wire [13:0] _T_69253; // @[Modules.scala 166:64:@15670.4]
  wire [13:0] buffer_4_527; // @[Modules.scala 166:64:@15671.4]
  wire [14:0] _T_69255; // @[Modules.scala 166:64:@15673.4]
  wire [13:0] _T_69256; // @[Modules.scala 166:64:@15674.4]
  wire [13:0] buffer_4_528; // @[Modules.scala 166:64:@15675.4]
  wire [14:0] _T_69258; // @[Modules.scala 166:64:@15677.4]
  wire [13:0] _T_69259; // @[Modules.scala 166:64:@15678.4]
  wire [13:0] buffer_4_529; // @[Modules.scala 166:64:@15679.4]
  wire [14:0] _T_69261; // @[Modules.scala 166:64:@15681.4]
  wire [13:0] _T_69262; // @[Modules.scala 166:64:@15682.4]
  wire [13:0] buffer_4_530; // @[Modules.scala 166:64:@15683.4]
  wire [14:0] _T_69264; // @[Modules.scala 166:64:@15685.4]
  wire [13:0] _T_69265; // @[Modules.scala 166:64:@15686.4]
  wire [13:0] buffer_4_531; // @[Modules.scala 166:64:@15687.4]
  wire [14:0] _T_69267; // @[Modules.scala 166:64:@15689.4]
  wire [13:0] _T_69268; // @[Modules.scala 166:64:@15690.4]
  wire [13:0] buffer_4_532; // @[Modules.scala 166:64:@15691.4]
  wire [14:0] _T_69270; // @[Modules.scala 166:64:@15693.4]
  wire [13:0] _T_69271; // @[Modules.scala 166:64:@15694.4]
  wire [13:0] buffer_4_533; // @[Modules.scala 166:64:@15695.4]
  wire [14:0] _T_69273; // @[Modules.scala 166:64:@15697.4]
  wire [13:0] _T_69274; // @[Modules.scala 166:64:@15698.4]
  wire [13:0] buffer_4_534; // @[Modules.scala 166:64:@15699.4]
  wire [14:0] _T_69276; // @[Modules.scala 166:64:@15701.4]
  wire [13:0] _T_69277; // @[Modules.scala 166:64:@15702.4]
  wire [13:0] buffer_4_535; // @[Modules.scala 166:64:@15703.4]
  wire [14:0] _T_69279; // @[Modules.scala 166:64:@15705.4]
  wire [13:0] _T_69280; // @[Modules.scala 166:64:@15706.4]
  wire [13:0] buffer_4_536; // @[Modules.scala 166:64:@15707.4]
  wire [14:0] _T_69282; // @[Modules.scala 166:64:@15709.4]
  wire [13:0] _T_69283; // @[Modules.scala 166:64:@15710.4]
  wire [13:0] buffer_4_537; // @[Modules.scala 166:64:@15711.4]
  wire [14:0] _T_69285; // @[Modules.scala 166:64:@15713.4]
  wire [13:0] _T_69286; // @[Modules.scala 166:64:@15714.4]
  wire [13:0] buffer_4_538; // @[Modules.scala 166:64:@15715.4]
  wire [14:0] _T_69288; // @[Modules.scala 166:64:@15717.4]
  wire [13:0] _T_69289; // @[Modules.scala 166:64:@15718.4]
  wire [13:0] buffer_4_539; // @[Modules.scala 166:64:@15719.4]
  wire [14:0] _T_69291; // @[Modules.scala 166:64:@15721.4]
  wire [13:0] _T_69292; // @[Modules.scala 166:64:@15722.4]
  wire [13:0] buffer_4_540; // @[Modules.scala 166:64:@15723.4]
  wire [14:0] _T_69294; // @[Modules.scala 166:64:@15725.4]
  wire [13:0] _T_69295; // @[Modules.scala 166:64:@15726.4]
  wire [13:0] buffer_4_541; // @[Modules.scala 166:64:@15727.4]
  wire [14:0] _T_69297; // @[Modules.scala 166:64:@15729.4]
  wire [13:0] _T_69298; // @[Modules.scala 166:64:@15730.4]
  wire [13:0] buffer_4_542; // @[Modules.scala 166:64:@15731.4]
  wire [14:0] _T_69300; // @[Modules.scala 166:64:@15733.4]
  wire [13:0] _T_69301; // @[Modules.scala 166:64:@15734.4]
  wire [13:0] buffer_4_543; // @[Modules.scala 166:64:@15735.4]
  wire [14:0] _T_69303; // @[Modules.scala 166:64:@15737.4]
  wire [13:0] _T_69304; // @[Modules.scala 166:64:@15738.4]
  wire [13:0] buffer_4_544; // @[Modules.scala 166:64:@15739.4]
  wire [14:0] _T_69306; // @[Modules.scala 166:64:@15741.4]
  wire [13:0] _T_69307; // @[Modules.scala 166:64:@15742.4]
  wire [13:0] buffer_4_545; // @[Modules.scala 166:64:@15743.4]
  wire [14:0] _T_69309; // @[Modules.scala 166:64:@15745.4]
  wire [13:0] _T_69310; // @[Modules.scala 166:64:@15746.4]
  wire [13:0] buffer_4_546; // @[Modules.scala 166:64:@15747.4]
  wire [14:0] _T_69312; // @[Modules.scala 166:64:@15749.4]
  wire [13:0] _T_69313; // @[Modules.scala 166:64:@15750.4]
  wire [13:0] buffer_4_547; // @[Modules.scala 166:64:@15751.4]
  wire [14:0] _T_69315; // @[Modules.scala 166:64:@15753.4]
  wire [13:0] _T_69316; // @[Modules.scala 166:64:@15754.4]
  wire [13:0] buffer_4_548; // @[Modules.scala 166:64:@15755.4]
  wire [14:0] _T_69318; // @[Modules.scala 166:64:@15757.4]
  wire [13:0] _T_69319; // @[Modules.scala 166:64:@15758.4]
  wire [13:0] buffer_4_549; // @[Modules.scala 166:64:@15759.4]
  wire [14:0] _T_69321; // @[Modules.scala 166:64:@15761.4]
  wire [13:0] _T_69322; // @[Modules.scala 166:64:@15762.4]
  wire [13:0] buffer_4_550; // @[Modules.scala 166:64:@15763.4]
  wire [14:0] _T_69324; // @[Modules.scala 166:64:@15765.4]
  wire [13:0] _T_69325; // @[Modules.scala 166:64:@15766.4]
  wire [13:0] buffer_4_551; // @[Modules.scala 166:64:@15767.4]
  wire [14:0] _T_69327; // @[Modules.scala 166:64:@15769.4]
  wire [13:0] _T_69328; // @[Modules.scala 166:64:@15770.4]
  wire [13:0] buffer_4_552; // @[Modules.scala 166:64:@15771.4]
  wire [14:0] _T_69330; // @[Modules.scala 166:64:@15773.4]
  wire [13:0] _T_69331; // @[Modules.scala 166:64:@15774.4]
  wire [13:0] buffer_4_553; // @[Modules.scala 166:64:@15775.4]
  wire [14:0] _T_69333; // @[Modules.scala 166:64:@15777.4]
  wire [13:0] _T_69334; // @[Modules.scala 166:64:@15778.4]
  wire [13:0] buffer_4_554; // @[Modules.scala 166:64:@15779.4]
  wire [14:0] _T_69336; // @[Modules.scala 166:64:@15781.4]
  wire [13:0] _T_69337; // @[Modules.scala 166:64:@15782.4]
  wire [13:0] buffer_4_555; // @[Modules.scala 166:64:@15783.4]
  wire [14:0] _T_69339; // @[Modules.scala 166:64:@15785.4]
  wire [13:0] _T_69340; // @[Modules.scala 166:64:@15786.4]
  wire [13:0] buffer_4_556; // @[Modules.scala 166:64:@15787.4]
  wire [14:0] _T_69342; // @[Modules.scala 166:64:@15789.4]
  wire [13:0] _T_69343; // @[Modules.scala 166:64:@15790.4]
  wire [13:0] buffer_4_557; // @[Modules.scala 166:64:@15791.4]
  wire [14:0] _T_69345; // @[Modules.scala 166:64:@15793.4]
  wire [13:0] _T_69346; // @[Modules.scala 166:64:@15794.4]
  wire [13:0] buffer_4_558; // @[Modules.scala 166:64:@15795.4]
  wire [14:0] _T_69348; // @[Modules.scala 166:64:@15797.4]
  wire [13:0] _T_69349; // @[Modules.scala 166:64:@15798.4]
  wire [13:0] buffer_4_559; // @[Modules.scala 166:64:@15799.4]
  wire [14:0] _T_69351; // @[Modules.scala 166:64:@15801.4]
  wire [13:0] _T_69352; // @[Modules.scala 166:64:@15802.4]
  wire [13:0] buffer_4_560; // @[Modules.scala 166:64:@15803.4]
  wire [14:0] _T_69354; // @[Modules.scala 166:64:@15805.4]
  wire [13:0] _T_69355; // @[Modules.scala 166:64:@15806.4]
  wire [13:0] buffer_4_561; // @[Modules.scala 166:64:@15807.4]
  wire [14:0] _T_69357; // @[Modules.scala 166:64:@15809.4]
  wire [13:0] _T_69358; // @[Modules.scala 166:64:@15810.4]
  wire [13:0] buffer_4_562; // @[Modules.scala 166:64:@15811.4]
  wire [14:0] _T_69360; // @[Modules.scala 166:64:@15813.4]
  wire [13:0] _T_69361; // @[Modules.scala 166:64:@15814.4]
  wire [13:0] buffer_4_563; // @[Modules.scala 166:64:@15815.4]
  wire [14:0] _T_69363; // @[Modules.scala 166:64:@15817.4]
  wire [13:0] _T_69364; // @[Modules.scala 166:64:@15818.4]
  wire [13:0] buffer_4_564; // @[Modules.scala 166:64:@15819.4]
  wire [14:0] _T_69366; // @[Modules.scala 166:64:@15821.4]
  wire [13:0] _T_69367; // @[Modules.scala 166:64:@15822.4]
  wire [13:0] buffer_4_565; // @[Modules.scala 166:64:@15823.4]
  wire [14:0] _T_69369; // @[Modules.scala 166:64:@15825.4]
  wire [13:0] _T_69370; // @[Modules.scala 166:64:@15826.4]
  wire [13:0] buffer_4_566; // @[Modules.scala 166:64:@15827.4]
  wire [14:0] _T_69372; // @[Modules.scala 166:64:@15829.4]
  wire [13:0] _T_69373; // @[Modules.scala 166:64:@15830.4]
  wire [13:0] buffer_4_567; // @[Modules.scala 166:64:@15831.4]
  wire [14:0] _T_69375; // @[Modules.scala 166:64:@15833.4]
  wire [13:0] _T_69376; // @[Modules.scala 166:64:@15834.4]
  wire [13:0] buffer_4_568; // @[Modules.scala 166:64:@15835.4]
  wire [14:0] _T_69378; // @[Modules.scala 166:64:@15837.4]
  wire [13:0] _T_69379; // @[Modules.scala 166:64:@15838.4]
  wire [13:0] buffer_4_569; // @[Modules.scala 166:64:@15839.4]
  wire [14:0] _T_69381; // @[Modules.scala 166:64:@15841.4]
  wire [13:0] _T_69382; // @[Modules.scala 166:64:@15842.4]
  wire [13:0] buffer_4_570; // @[Modules.scala 166:64:@15843.4]
  wire [14:0] _T_69384; // @[Modules.scala 166:64:@15845.4]
  wire [13:0] _T_69385; // @[Modules.scala 166:64:@15846.4]
  wire [13:0] buffer_4_571; // @[Modules.scala 166:64:@15847.4]
  wire [14:0] _T_69387; // @[Modules.scala 166:64:@15849.4]
  wire [13:0] _T_69388; // @[Modules.scala 166:64:@15850.4]
  wire [13:0] buffer_4_572; // @[Modules.scala 166:64:@15851.4]
  wire [14:0] _T_69390; // @[Modules.scala 166:64:@15853.4]
  wire [13:0] _T_69391; // @[Modules.scala 166:64:@15854.4]
  wire [13:0] buffer_4_573; // @[Modules.scala 166:64:@15855.4]
  wire [14:0] _T_69393; // @[Modules.scala 166:64:@15857.4]
  wire [13:0] _T_69394; // @[Modules.scala 166:64:@15858.4]
  wire [13:0] buffer_4_574; // @[Modules.scala 166:64:@15859.4]
  wire [14:0] _T_69396; // @[Modules.scala 166:64:@15861.4]
  wire [13:0] _T_69397; // @[Modules.scala 166:64:@15862.4]
  wire [13:0] buffer_4_575; // @[Modules.scala 166:64:@15863.4]
  wire [14:0] _T_69399; // @[Modules.scala 166:64:@15865.4]
  wire [13:0] _T_69400; // @[Modules.scala 166:64:@15866.4]
  wire [13:0] buffer_4_576; // @[Modules.scala 166:64:@15867.4]
  wire [14:0] _T_69402; // @[Modules.scala 166:64:@15869.4]
  wire [13:0] _T_69403; // @[Modules.scala 166:64:@15870.4]
  wire [13:0] buffer_4_577; // @[Modules.scala 166:64:@15871.4]
  wire [14:0] _T_69405; // @[Modules.scala 166:64:@15873.4]
  wire [13:0] _T_69406; // @[Modules.scala 166:64:@15874.4]
  wire [13:0] buffer_4_578; // @[Modules.scala 166:64:@15875.4]
  wire [14:0] _T_69408; // @[Modules.scala 166:64:@15877.4]
  wire [13:0] _T_69409; // @[Modules.scala 166:64:@15878.4]
  wire [13:0] buffer_4_579; // @[Modules.scala 166:64:@15879.4]
  wire [14:0] _T_69411; // @[Modules.scala 172:66:@15881.4]
  wire [13:0] _T_69412; // @[Modules.scala 172:66:@15882.4]
  wire [13:0] buffer_4_580; // @[Modules.scala 172:66:@15883.4]
  wire [14:0] _T_69414; // @[Modules.scala 166:64:@15885.4]
  wire [13:0] _T_69415; // @[Modules.scala 166:64:@15886.4]
  wire [13:0] buffer_4_581; // @[Modules.scala 166:64:@15887.4]
  wire [14:0] _T_69417; // @[Modules.scala 166:64:@15889.4]
  wire [13:0] _T_69418; // @[Modules.scala 166:64:@15890.4]
  wire [13:0] buffer_4_582; // @[Modules.scala 166:64:@15891.4]
  wire [14:0] _T_69420; // @[Modules.scala 166:64:@15893.4]
  wire [13:0] _T_69421; // @[Modules.scala 166:64:@15894.4]
  wire [13:0] buffer_4_583; // @[Modules.scala 166:64:@15895.4]
  wire [14:0] _T_69423; // @[Modules.scala 166:64:@15897.4]
  wire [13:0] _T_69424; // @[Modules.scala 166:64:@15898.4]
  wire [13:0] buffer_4_584; // @[Modules.scala 166:64:@15899.4]
  wire [14:0] _T_69426; // @[Modules.scala 166:64:@15901.4]
  wire [13:0] _T_69427; // @[Modules.scala 166:64:@15902.4]
  wire [13:0] buffer_4_585; // @[Modules.scala 166:64:@15903.4]
  wire [14:0] _T_69429; // @[Modules.scala 166:64:@15905.4]
  wire [13:0] _T_69430; // @[Modules.scala 166:64:@15906.4]
  wire [13:0] buffer_4_586; // @[Modules.scala 166:64:@15907.4]
  wire [14:0] _T_69432; // @[Modules.scala 166:64:@15909.4]
  wire [13:0] _T_69433; // @[Modules.scala 166:64:@15910.4]
  wire [13:0] buffer_4_587; // @[Modules.scala 166:64:@15911.4]
  wire [14:0] _T_69435; // @[Modules.scala 166:64:@15913.4]
  wire [13:0] _T_69436; // @[Modules.scala 166:64:@15914.4]
  wire [13:0] buffer_4_588; // @[Modules.scala 166:64:@15915.4]
  wire [14:0] _T_69438; // @[Modules.scala 166:64:@15917.4]
  wire [13:0] _T_69439; // @[Modules.scala 166:64:@15918.4]
  wire [13:0] buffer_4_589; // @[Modules.scala 166:64:@15919.4]
  wire [14:0] _T_69441; // @[Modules.scala 166:64:@15921.4]
  wire [13:0] _T_69442; // @[Modules.scala 166:64:@15922.4]
  wire [13:0] buffer_4_590; // @[Modules.scala 166:64:@15923.4]
  wire [14:0] _T_69444; // @[Modules.scala 166:64:@15925.4]
  wire [13:0] _T_69445; // @[Modules.scala 166:64:@15926.4]
  wire [13:0] buffer_4_591; // @[Modules.scala 166:64:@15927.4]
  wire [14:0] _T_69447; // @[Modules.scala 166:64:@15929.4]
  wire [13:0] _T_69448; // @[Modules.scala 166:64:@15930.4]
  wire [13:0] buffer_4_592; // @[Modules.scala 166:64:@15931.4]
  wire [14:0] _T_69450; // @[Modules.scala 166:64:@15933.4]
  wire [13:0] _T_69451; // @[Modules.scala 166:64:@15934.4]
  wire [13:0] buffer_4_593; // @[Modules.scala 166:64:@15935.4]
  wire [14:0] _T_69453; // @[Modules.scala 172:66:@15937.4]
  wire [13:0] _T_69454; // @[Modules.scala 172:66:@15938.4]
  wire [13:0] buffer_4_594; // @[Modules.scala 172:66:@15939.4]
  wire [14:0] _T_69456; // @[Modules.scala 166:64:@15941.4]
  wire [13:0] _T_69457; // @[Modules.scala 166:64:@15942.4]
  wire [13:0] buffer_4_595; // @[Modules.scala 166:64:@15943.4]
  wire [14:0] _T_69459; // @[Modules.scala 166:64:@15945.4]
  wire [13:0] _T_69460; // @[Modules.scala 166:64:@15946.4]
  wire [13:0] buffer_4_596; // @[Modules.scala 166:64:@15947.4]
  wire [14:0] _T_69462; // @[Modules.scala 160:64:@15949.4]
  wire [13:0] _T_69463; // @[Modules.scala 160:64:@15950.4]
  wire [13:0] buffer_4_597; // @[Modules.scala 160:64:@15951.4]
  wire [14:0] _T_69465; // @[Modules.scala 172:66:@15953.4]
  wire [13:0] _T_69466; // @[Modules.scala 172:66:@15954.4]
  wire [13:0] buffer_4_598; // @[Modules.scala 172:66:@15955.4]
  wire [5:0] _T_69469; // @[Modules.scala 143:74:@16142.4]
  wire [4:0] _T_69471; // @[Modules.scala 144:80:@16143.4]
  wire [5:0] _GEN_357; // @[Modules.scala 143:103:@16144.4]
  wire [6:0] _T_69472; // @[Modules.scala 143:103:@16144.4]
  wire [5:0] _T_69473; // @[Modules.scala 143:103:@16145.4]
  wire [5:0] _T_69474; // @[Modules.scala 143:103:@16146.4]
  wire [6:0] _T_69500; // @[Modules.scala 143:103:@16168.4]
  wire [5:0] _T_69501; // @[Modules.scala 143:103:@16169.4]
  wire [5:0] _T_69502; // @[Modules.scala 143:103:@16170.4]
  wire [5:0] _T_69514; // @[Modules.scala 143:103:@16180.4]
  wire [4:0] _T_69515; // @[Modules.scala 143:103:@16181.4]
  wire [4:0] _T_69516; // @[Modules.scala 143:103:@16182.4]
  wire [5:0] _GEN_359; // @[Modules.scala 143:103:@16198.4]
  wire [6:0] _T_69535; // @[Modules.scala 143:103:@16198.4]
  wire [5:0] _T_69536; // @[Modules.scala 143:103:@16199.4]
  wire [5:0] _T_69537; // @[Modules.scala 143:103:@16200.4]
  wire [4:0] _T_69548; // @[Modules.scala 144:80:@16209.4]
  wire [5:0] _GEN_360; // @[Modules.scala 143:103:@16210.4]
  wire [6:0] _T_69549; // @[Modules.scala 143:103:@16210.4]
  wire [5:0] _T_69550; // @[Modules.scala 143:103:@16211.4]
  wire [5:0] _T_69551; // @[Modules.scala 143:103:@16212.4]
  wire [6:0] _T_69556; // @[Modules.scala 143:103:@16216.4]
  wire [5:0] _T_69557; // @[Modules.scala 143:103:@16217.4]
  wire [5:0] _T_69558; // @[Modules.scala 143:103:@16218.4]
  wire [6:0] _T_69619; // @[Modules.scala 143:103:@16270.4]
  wire [5:0] _T_69620; // @[Modules.scala 143:103:@16271.4]
  wire [5:0] _T_69621; // @[Modules.scala 143:103:@16272.4]
  wire [5:0] _GEN_364; // @[Modules.scala 143:103:@16288.4]
  wire [6:0] _T_69640; // @[Modules.scala 143:103:@16288.4]
  wire [5:0] _T_69641; // @[Modules.scala 143:103:@16289.4]
  wire [5:0] _T_69642; // @[Modules.scala 143:103:@16290.4]
  wire [5:0] _T_69661; // @[Modules.scala 143:103:@16306.4]
  wire [4:0] _T_69662; // @[Modules.scala 143:103:@16307.4]
  wire [4:0] _T_69663; // @[Modules.scala 143:103:@16308.4]
  wire [5:0] _T_69668; // @[Modules.scala 143:103:@16312.4]
  wire [4:0] _T_69669; // @[Modules.scala 143:103:@16313.4]
  wire [4:0] _T_69670; // @[Modules.scala 143:103:@16314.4]
  wire [5:0] _T_69696; // @[Modules.scala 143:103:@16336.4]
  wire [4:0] _T_69697; // @[Modules.scala 143:103:@16337.4]
  wire [4:0] _T_69698; // @[Modules.scala 143:103:@16338.4]
  wire [5:0] _T_69703; // @[Modules.scala 143:103:@16342.4]
  wire [4:0] _T_69704; // @[Modules.scala 143:103:@16343.4]
  wire [4:0] _T_69705; // @[Modules.scala 143:103:@16344.4]
  wire [5:0] _GEN_365; // @[Modules.scala 143:103:@16348.4]
  wire [6:0] _T_69710; // @[Modules.scala 143:103:@16348.4]
  wire [5:0] _T_69711; // @[Modules.scala 143:103:@16349.4]
  wire [5:0] _T_69712; // @[Modules.scala 143:103:@16350.4]
  wire [6:0] _T_69724; // @[Modules.scala 143:103:@16360.4]
  wire [5:0] _T_69725; // @[Modules.scala 143:103:@16361.4]
  wire [5:0] _T_69726; // @[Modules.scala 143:103:@16362.4]
  wire [5:0] _T_69749; // @[Modules.scala 143:74:@16382.4]
  wire [6:0] _T_69752; // @[Modules.scala 143:103:@16384.4]
  wire [5:0] _T_69753; // @[Modules.scala 143:103:@16385.4]
  wire [5:0] _T_69754; // @[Modules.scala 143:103:@16386.4]
  wire [4:0] _T_69763; // @[Modules.scala 143:74:@16394.4]
  wire [4:0] _T_69765; // @[Modules.scala 144:80:@16395.4]
  wire [5:0] _T_69766; // @[Modules.scala 143:103:@16396.4]
  wire [4:0] _T_69767; // @[Modules.scala 143:103:@16397.4]
  wire [4:0] _T_69768; // @[Modules.scala 143:103:@16398.4]
  wire [4:0] _T_69770; // @[Modules.scala 143:74:@16400.4]
  wire [5:0] _T_69773; // @[Modules.scala 143:103:@16402.4]
  wire [4:0] _T_69774; // @[Modules.scala 143:103:@16403.4]
  wire [4:0] _T_69775; // @[Modules.scala 143:103:@16404.4]
  wire [5:0] _GEN_366; // @[Modules.scala 143:103:@16408.4]
  wire [6:0] _T_69780; // @[Modules.scala 143:103:@16408.4]
  wire [5:0] _T_69781; // @[Modules.scala 143:103:@16409.4]
  wire [5:0] _T_69782; // @[Modules.scala 143:103:@16410.4]
  wire [6:0] _T_69794; // @[Modules.scala 143:103:@16420.4]
  wire [5:0] _T_69795; // @[Modules.scala 143:103:@16421.4]
  wire [5:0] _T_69796; // @[Modules.scala 143:103:@16422.4]
  wire [5:0] _T_69819; // @[Modules.scala 143:74:@16442.4]
  wire [6:0] _T_69822; // @[Modules.scala 143:103:@16444.4]
  wire [5:0] _T_69823; // @[Modules.scala 143:103:@16445.4]
  wire [5:0] _T_69824; // @[Modules.scala 143:103:@16446.4]
  wire [5:0] _T_69826; // @[Modules.scala 143:74:@16448.4]
  wire [5:0] _T_69828; // @[Modules.scala 144:80:@16449.4]
  wire [6:0] _T_69829; // @[Modules.scala 143:103:@16450.4]
  wire [5:0] _T_69830; // @[Modules.scala 143:103:@16451.4]
  wire [5:0] _T_69831; // @[Modules.scala 143:103:@16452.4]
  wire [5:0] _T_69833; // @[Modules.scala 143:74:@16454.4]
  wire [5:0] _GEN_369; // @[Modules.scala 143:103:@16456.4]
  wire [6:0] _T_69836; // @[Modules.scala 143:103:@16456.4]
  wire [5:0] _T_69837; // @[Modules.scala 143:103:@16457.4]
  wire [5:0] _T_69838; // @[Modules.scala 143:103:@16458.4]
  wire [5:0] _T_69843; // @[Modules.scala 143:103:@16462.4]
  wire [4:0] _T_69844; // @[Modules.scala 143:103:@16463.4]
  wire [4:0] _T_69845; // @[Modules.scala 143:103:@16464.4]
  wire [5:0] _GEN_370; // @[Modules.scala 143:103:@16474.4]
  wire [6:0] _T_69857; // @[Modules.scala 143:103:@16474.4]
  wire [5:0] _T_69858; // @[Modules.scala 143:103:@16475.4]
  wire [5:0] _T_69859; // @[Modules.scala 143:103:@16476.4]
  wire [5:0] _T_69878; // @[Modules.scala 143:103:@16492.4]
  wire [4:0] _T_69879; // @[Modules.scala 143:103:@16493.4]
  wire [4:0] _T_69880; // @[Modules.scala 143:103:@16494.4]
  wire [5:0] _GEN_373; // @[Modules.scala 143:103:@16498.4]
  wire [6:0] _T_69885; // @[Modules.scala 143:103:@16498.4]
  wire [5:0] _T_69886; // @[Modules.scala 143:103:@16499.4]
  wire [5:0] _T_69887; // @[Modules.scala 143:103:@16500.4]
  wire [5:0] _T_69891; // @[Modules.scala 144:80:@16503.4]
  wire [6:0] _T_69892; // @[Modules.scala 143:103:@16504.4]
  wire [5:0] _T_69893; // @[Modules.scala 143:103:@16505.4]
  wire [5:0] _T_69894; // @[Modules.scala 143:103:@16506.4]
  wire [6:0] _T_69899; // @[Modules.scala 143:103:@16510.4]
  wire [5:0] _T_69900; // @[Modules.scala 143:103:@16511.4]
  wire [5:0] _T_69901; // @[Modules.scala 143:103:@16512.4]
  wire [6:0] _T_69913; // @[Modules.scala 143:103:@16522.4]
  wire [5:0] _T_69914; // @[Modules.scala 143:103:@16523.4]
  wire [5:0] _T_69915; // @[Modules.scala 143:103:@16524.4]
  wire [6:0] _T_69920; // @[Modules.scala 143:103:@16528.4]
  wire [5:0] _T_69921; // @[Modules.scala 143:103:@16529.4]
  wire [5:0] _T_69922; // @[Modules.scala 143:103:@16530.4]
  wire [5:0] _T_69924; // @[Modules.scala 143:74:@16532.4]
  wire [6:0] _T_69927; // @[Modules.scala 143:103:@16534.4]
  wire [5:0] _T_69928; // @[Modules.scala 143:103:@16535.4]
  wire [5:0] _T_69929; // @[Modules.scala 143:103:@16536.4]
  wire [5:0] _GEN_375; // @[Modules.scala 143:103:@16540.4]
  wire [6:0] _T_69934; // @[Modules.scala 143:103:@16540.4]
  wire [5:0] _T_69935; // @[Modules.scala 143:103:@16541.4]
  wire [5:0] _T_69936; // @[Modules.scala 143:103:@16542.4]
  wire [5:0] _T_69938; // @[Modules.scala 143:74:@16544.4]
  wire [6:0] _T_69941; // @[Modules.scala 143:103:@16546.4]
  wire [5:0] _T_69942; // @[Modules.scala 143:103:@16547.4]
  wire [5:0] _T_69943; // @[Modules.scala 143:103:@16548.4]
  wire [4:0] _T_69947; // @[Modules.scala 144:80:@16551.4]
  wire [5:0] _T_69948; // @[Modules.scala 143:103:@16552.4]
  wire [4:0] _T_69949; // @[Modules.scala 143:103:@16553.4]
  wire [4:0] _T_69950; // @[Modules.scala 143:103:@16554.4]
  wire [6:0] _T_69955; // @[Modules.scala 143:103:@16558.4]
  wire [5:0] _T_69956; // @[Modules.scala 143:103:@16559.4]
  wire [5:0] _T_69957; // @[Modules.scala 143:103:@16560.4]
  wire [5:0] _GEN_377; // @[Modules.scala 143:103:@16564.4]
  wire [6:0] _T_69962; // @[Modules.scala 143:103:@16564.4]
  wire [5:0] _T_69963; // @[Modules.scala 143:103:@16565.4]
  wire [5:0] _T_69964; // @[Modules.scala 143:103:@16566.4]
  wire [5:0] _T_69968; // @[Modules.scala 144:80:@16569.4]
  wire [6:0] _T_69969; // @[Modules.scala 143:103:@16570.4]
  wire [5:0] _T_69970; // @[Modules.scala 143:103:@16571.4]
  wire [5:0] _T_69971; // @[Modules.scala 143:103:@16572.4]
  wire [5:0] _T_69973; // @[Modules.scala 143:74:@16574.4]
  wire [6:0] _T_69976; // @[Modules.scala 143:103:@16576.4]
  wire [5:0] _T_69977; // @[Modules.scala 143:103:@16577.4]
  wire [5:0] _T_69978; // @[Modules.scala 143:103:@16578.4]
  wire [6:0] _T_70004; // @[Modules.scala 143:103:@16600.4]
  wire [5:0] _T_70005; // @[Modules.scala 143:103:@16601.4]
  wire [5:0] _T_70006; // @[Modules.scala 143:103:@16602.4]
  wire [5:0] _T_70010; // @[Modules.scala 144:80:@16605.4]
  wire [6:0] _T_70011; // @[Modules.scala 143:103:@16606.4]
  wire [5:0] _T_70012; // @[Modules.scala 143:103:@16607.4]
  wire [5:0] _T_70013; // @[Modules.scala 143:103:@16608.4]
  wire [5:0] _GEN_378; // @[Modules.scala 143:103:@16624.4]
  wire [6:0] _T_70032; // @[Modules.scala 143:103:@16624.4]
  wire [5:0] _T_70033; // @[Modules.scala 143:103:@16625.4]
  wire [5:0] _T_70034; // @[Modules.scala 143:103:@16626.4]
  wire [4:0] _T_70036; // @[Modules.scala 143:74:@16628.4]
  wire [5:0] _GEN_379; // @[Modules.scala 143:103:@16630.4]
  wire [6:0] _T_70039; // @[Modules.scala 143:103:@16630.4]
  wire [5:0] _T_70040; // @[Modules.scala 143:103:@16631.4]
  wire [5:0] _T_70041; // @[Modules.scala 143:103:@16632.4]
  wire [5:0] _T_70057; // @[Modules.scala 143:74:@16646.4]
  wire [5:0] _T_70059; // @[Modules.scala 144:80:@16647.4]
  wire [6:0] _T_70060; // @[Modules.scala 143:103:@16648.4]
  wire [5:0] _T_70061; // @[Modules.scala 143:103:@16649.4]
  wire [5:0] _T_70062; // @[Modules.scala 143:103:@16650.4]
  wire [6:0] _T_70067; // @[Modules.scala 143:103:@16654.4]
  wire [5:0] _T_70068; // @[Modules.scala 143:103:@16655.4]
  wire [5:0] _T_70069; // @[Modules.scala 143:103:@16656.4]
  wire [5:0] _T_70099; // @[Modules.scala 143:74:@16682.4]
  wire [6:0] _T_70102; // @[Modules.scala 143:103:@16684.4]
  wire [5:0] _T_70103; // @[Modules.scala 143:103:@16685.4]
  wire [5:0] _T_70104; // @[Modules.scala 143:103:@16686.4]
  wire [6:0] _T_70109; // @[Modules.scala 143:103:@16690.4]
  wire [5:0] _T_70110; // @[Modules.scala 143:103:@16691.4]
  wire [5:0] _T_70111; // @[Modules.scala 143:103:@16692.4]
  wire [6:0] _T_70116; // @[Modules.scala 143:103:@16696.4]
  wire [5:0] _T_70117; // @[Modules.scala 143:103:@16697.4]
  wire [5:0] _T_70118; // @[Modules.scala 143:103:@16698.4]
  wire [6:0] _T_70123; // @[Modules.scala 143:103:@16702.4]
  wire [5:0] _T_70124; // @[Modules.scala 143:103:@16703.4]
  wire [5:0] _T_70125; // @[Modules.scala 143:103:@16704.4]
  wire [6:0] _T_70137; // @[Modules.scala 143:103:@16714.4]
  wire [5:0] _T_70138; // @[Modules.scala 143:103:@16715.4]
  wire [5:0] _T_70139; // @[Modules.scala 143:103:@16716.4]
  wire [5:0] _T_70143; // @[Modules.scala 144:80:@16719.4]
  wire [6:0] _T_70144; // @[Modules.scala 143:103:@16720.4]
  wire [5:0] _T_70145; // @[Modules.scala 143:103:@16721.4]
  wire [5:0] _T_70146; // @[Modules.scala 143:103:@16722.4]
  wire [5:0] _T_70148; // @[Modules.scala 143:74:@16724.4]
  wire [6:0] _T_70151; // @[Modules.scala 143:103:@16726.4]
  wire [5:0] _T_70152; // @[Modules.scala 143:103:@16727.4]
  wire [5:0] _T_70153; // @[Modules.scala 143:103:@16728.4]
  wire [6:0] _T_70158; // @[Modules.scala 143:103:@16732.4]
  wire [5:0] _T_70159; // @[Modules.scala 143:103:@16733.4]
  wire [5:0] _T_70160; // @[Modules.scala 143:103:@16734.4]
  wire [6:0] _T_70186; // @[Modules.scala 143:103:@16756.4]
  wire [5:0] _T_70187; // @[Modules.scala 143:103:@16757.4]
  wire [5:0] _T_70188; // @[Modules.scala 143:103:@16758.4]
  wire [5:0] _T_70192; // @[Modules.scala 144:80:@16761.4]
  wire [6:0] _T_70193; // @[Modules.scala 143:103:@16762.4]
  wire [5:0] _T_70194; // @[Modules.scala 143:103:@16763.4]
  wire [5:0] _T_70195; // @[Modules.scala 143:103:@16764.4]
  wire [6:0] _T_70200; // @[Modules.scala 143:103:@16768.4]
  wire [5:0] _T_70201; // @[Modules.scala 143:103:@16769.4]
  wire [5:0] _T_70202; // @[Modules.scala 143:103:@16770.4]
  wire [6:0] _T_70207; // @[Modules.scala 143:103:@16774.4]
  wire [5:0] _T_70208; // @[Modules.scala 143:103:@16775.4]
  wire [5:0] _T_70209; // @[Modules.scala 143:103:@16776.4]
  wire [5:0] _T_70213; // @[Modules.scala 144:80:@16779.4]
  wire [6:0] _T_70214; // @[Modules.scala 143:103:@16780.4]
  wire [5:0] _T_70215; // @[Modules.scala 143:103:@16781.4]
  wire [5:0] _T_70216; // @[Modules.scala 143:103:@16782.4]
  wire [4:0] _T_70220; // @[Modules.scala 144:80:@16785.4]
  wire [5:0] _GEN_380; // @[Modules.scala 143:103:@16786.4]
  wire [6:0] _T_70221; // @[Modules.scala 143:103:@16786.4]
  wire [5:0] _T_70222; // @[Modules.scala 143:103:@16787.4]
  wire [5:0] _T_70223; // @[Modules.scala 143:103:@16788.4]
  wire [6:0] _T_70235; // @[Modules.scala 143:103:@16798.4]
  wire [5:0] _T_70236; // @[Modules.scala 143:103:@16799.4]
  wire [5:0] _T_70237; // @[Modules.scala 143:103:@16800.4]
  wire [6:0] _T_70242; // @[Modules.scala 143:103:@16804.4]
  wire [5:0] _T_70243; // @[Modules.scala 143:103:@16805.4]
  wire [5:0] _T_70244; // @[Modules.scala 143:103:@16806.4]
  wire [6:0] _T_70249; // @[Modules.scala 143:103:@16810.4]
  wire [5:0] _T_70250; // @[Modules.scala 143:103:@16811.4]
  wire [5:0] _T_70251; // @[Modules.scala 143:103:@16812.4]
  wire [6:0] _T_70256; // @[Modules.scala 143:103:@16816.4]
  wire [5:0] _T_70257; // @[Modules.scala 143:103:@16817.4]
  wire [5:0] _T_70258; // @[Modules.scala 143:103:@16818.4]
  wire [6:0] _T_70270; // @[Modules.scala 143:103:@16828.4]
  wire [5:0] _T_70271; // @[Modules.scala 143:103:@16829.4]
  wire [5:0] _T_70272; // @[Modules.scala 143:103:@16830.4]
  wire [6:0] _T_70277; // @[Modules.scala 143:103:@16834.4]
  wire [5:0] _T_70278; // @[Modules.scala 143:103:@16835.4]
  wire [5:0] _T_70279; // @[Modules.scala 143:103:@16836.4]
  wire [5:0] _T_70281; // @[Modules.scala 143:74:@16838.4]
  wire [6:0] _T_70284; // @[Modules.scala 143:103:@16840.4]
  wire [5:0] _T_70285; // @[Modules.scala 143:103:@16841.4]
  wire [5:0] _T_70286; // @[Modules.scala 143:103:@16842.4]
  wire [6:0] _T_70291; // @[Modules.scala 143:103:@16846.4]
  wire [5:0] _T_70292; // @[Modules.scala 143:103:@16847.4]
  wire [5:0] _T_70293; // @[Modules.scala 143:103:@16848.4]
  wire [5:0] _T_70319; // @[Modules.scala 143:103:@16870.4]
  wire [4:0] _T_70320; // @[Modules.scala 143:103:@16871.4]
  wire [4:0] _T_70321; // @[Modules.scala 143:103:@16872.4]
  wire [5:0] _GEN_382; // @[Modules.scala 143:103:@16876.4]
  wire [6:0] _T_70326; // @[Modules.scala 143:103:@16876.4]
  wire [5:0] _T_70327; // @[Modules.scala 143:103:@16877.4]
  wire [5:0] _T_70328; // @[Modules.scala 143:103:@16878.4]
  wire [6:0] _T_70333; // @[Modules.scala 143:103:@16882.4]
  wire [5:0] _T_70334; // @[Modules.scala 143:103:@16883.4]
  wire [5:0] _T_70335; // @[Modules.scala 143:103:@16884.4]
  wire [6:0] _T_70340; // @[Modules.scala 143:103:@16888.4]
  wire [5:0] _T_70341; // @[Modules.scala 143:103:@16889.4]
  wire [5:0] _T_70342; // @[Modules.scala 143:103:@16890.4]
  wire [5:0] _T_70347; // @[Modules.scala 143:103:@16894.4]
  wire [4:0] _T_70348; // @[Modules.scala 143:103:@16895.4]
  wire [4:0] _T_70349; // @[Modules.scala 143:103:@16896.4]
  wire [5:0] _T_70351; // @[Modules.scala 143:74:@16898.4]
  wire [5:0] _T_70353; // @[Modules.scala 144:80:@16899.4]
  wire [6:0] _T_70354; // @[Modules.scala 143:103:@16900.4]
  wire [5:0] _T_70355; // @[Modules.scala 143:103:@16901.4]
  wire [5:0] _T_70356; // @[Modules.scala 143:103:@16902.4]
  wire [5:0] _T_70368; // @[Modules.scala 143:103:@16912.4]
  wire [4:0] _T_70369; // @[Modules.scala 143:103:@16913.4]
  wire [4:0] _T_70370; // @[Modules.scala 143:103:@16914.4]
  wire [6:0] _T_70382; // @[Modules.scala 143:103:@16924.4]
  wire [5:0] _T_70383; // @[Modules.scala 143:103:@16925.4]
  wire [5:0] _T_70384; // @[Modules.scala 143:103:@16926.4]
  wire [5:0] _GEN_384; // @[Modules.scala 143:103:@16942.4]
  wire [6:0] _T_70403; // @[Modules.scala 143:103:@16942.4]
  wire [5:0] _T_70404; // @[Modules.scala 143:103:@16943.4]
  wire [5:0] _T_70405; // @[Modules.scala 143:103:@16944.4]
  wire [5:0] _T_70410; // @[Modules.scala 143:103:@16948.4]
  wire [4:0] _T_70411; // @[Modules.scala 143:103:@16949.4]
  wire [4:0] _T_70412; // @[Modules.scala 143:103:@16950.4]
  wire [4:0] _T_70414; // @[Modules.scala 143:74:@16952.4]
  wire [5:0] _T_70417; // @[Modules.scala 143:103:@16954.4]
  wire [4:0] _T_70418; // @[Modules.scala 143:103:@16955.4]
  wire [4:0] _T_70419; // @[Modules.scala 143:103:@16956.4]
  wire [6:0] _T_70466; // @[Modules.scala 143:103:@16996.4]
  wire [5:0] _T_70467; // @[Modules.scala 143:103:@16997.4]
  wire [5:0] _T_70468; // @[Modules.scala 143:103:@16998.4]
  wire [5:0] _T_70473; // @[Modules.scala 143:103:@17002.4]
  wire [4:0] _T_70474; // @[Modules.scala 143:103:@17003.4]
  wire [4:0] _T_70475; // @[Modules.scala 143:103:@17004.4]
  wire [5:0] _T_70480; // @[Modules.scala 143:103:@17008.4]
  wire [4:0] _T_70481; // @[Modules.scala 143:103:@17009.4]
  wire [4:0] _T_70482; // @[Modules.scala 143:103:@17010.4]
  wire [6:0] _T_70487; // @[Modules.scala 143:103:@17014.4]
  wire [5:0] _T_70488; // @[Modules.scala 143:103:@17015.4]
  wire [5:0] _T_70489; // @[Modules.scala 143:103:@17016.4]
  wire [4:0] _T_70491; // @[Modules.scala 143:74:@17018.4]
  wire [5:0] _GEN_387; // @[Modules.scala 143:103:@17020.4]
  wire [6:0] _T_70494; // @[Modules.scala 143:103:@17020.4]
  wire [5:0] _T_70495; // @[Modules.scala 143:103:@17021.4]
  wire [5:0] _T_70496; // @[Modules.scala 143:103:@17022.4]
  wire [5:0] _GEN_388; // @[Modules.scala 143:103:@17026.4]
  wire [6:0] _T_70501; // @[Modules.scala 143:103:@17026.4]
  wire [5:0] _T_70502; // @[Modules.scala 143:103:@17027.4]
  wire [5:0] _T_70503; // @[Modules.scala 143:103:@17028.4]
  wire [5:0] _GEN_389; // @[Modules.scala 143:103:@17038.4]
  wire [6:0] _T_70515; // @[Modules.scala 143:103:@17038.4]
  wire [5:0] _T_70516; // @[Modules.scala 143:103:@17039.4]
  wire [5:0] _T_70517; // @[Modules.scala 143:103:@17040.4]
  wire [6:0] _T_70522; // @[Modules.scala 143:103:@17044.4]
  wire [5:0] _T_70523; // @[Modules.scala 143:103:@17045.4]
  wire [5:0] _T_70524; // @[Modules.scala 143:103:@17046.4]
  wire [5:0] _T_70529; // @[Modules.scala 143:103:@17050.4]
  wire [4:0] _T_70530; // @[Modules.scala 143:103:@17051.4]
  wire [4:0] _T_70531; // @[Modules.scala 143:103:@17052.4]
  wire [4:0] _T_70533; // @[Modules.scala 143:74:@17054.4]
  wire [5:0] _T_70536; // @[Modules.scala 143:103:@17056.4]
  wire [4:0] _T_70537; // @[Modules.scala 143:103:@17057.4]
  wire [4:0] _T_70538; // @[Modules.scala 143:103:@17058.4]
  wire [5:0] _T_70543; // @[Modules.scala 143:103:@17062.4]
  wire [4:0] _T_70544; // @[Modules.scala 143:103:@17063.4]
  wire [4:0] _T_70545; // @[Modules.scala 143:103:@17064.4]
  wire [5:0] _T_70550; // @[Modules.scala 143:103:@17068.4]
  wire [4:0] _T_70551; // @[Modules.scala 143:103:@17069.4]
  wire [4:0] _T_70552; // @[Modules.scala 143:103:@17070.4]
  wire [5:0] _T_70557; // @[Modules.scala 143:103:@17074.4]
  wire [4:0] _T_70558; // @[Modules.scala 143:103:@17075.4]
  wire [4:0] _T_70559; // @[Modules.scala 143:103:@17076.4]
  wire [4:0] _T_70570; // @[Modules.scala 144:80:@17085.4]
  wire [5:0] _T_70571; // @[Modules.scala 143:103:@17086.4]
  wire [4:0] _T_70572; // @[Modules.scala 143:103:@17087.4]
  wire [4:0] _T_70573; // @[Modules.scala 143:103:@17088.4]
  wire [4:0] _T_70575; // @[Modules.scala 143:74:@17090.4]
  wire [5:0] _GEN_390; // @[Modules.scala 143:103:@17092.4]
  wire [6:0] _T_70578; // @[Modules.scala 143:103:@17092.4]
  wire [5:0] _T_70579; // @[Modules.scala 143:103:@17093.4]
  wire [5:0] _T_70580; // @[Modules.scala 143:103:@17094.4]
  wire [4:0] _T_70584; // @[Modules.scala 144:80:@17097.4]
  wire [5:0] _GEN_391; // @[Modules.scala 143:103:@17098.4]
  wire [6:0] _T_70585; // @[Modules.scala 143:103:@17098.4]
  wire [5:0] _T_70586; // @[Modules.scala 143:103:@17099.4]
  wire [5:0] _T_70587; // @[Modules.scala 143:103:@17100.4]
  wire [4:0] _T_70589; // @[Modules.scala 143:74:@17102.4]
  wire [5:0] _T_70592; // @[Modules.scala 143:103:@17104.4]
  wire [4:0] _T_70593; // @[Modules.scala 143:103:@17105.4]
  wire [4:0] _T_70594; // @[Modules.scala 143:103:@17106.4]
  wire [5:0] _T_70599; // @[Modules.scala 143:103:@17110.4]
  wire [4:0] _T_70600; // @[Modules.scala 143:103:@17111.4]
  wire [4:0] _T_70601; // @[Modules.scala 143:103:@17112.4]
  wire [5:0] _T_70605; // @[Modules.scala 144:80:@17115.4]
  wire [5:0] _GEN_392; // @[Modules.scala 143:103:@17116.4]
  wire [6:0] _T_70606; // @[Modules.scala 143:103:@17116.4]
  wire [5:0] _T_70607; // @[Modules.scala 143:103:@17117.4]
  wire [5:0] _T_70608; // @[Modules.scala 143:103:@17118.4]
  wire [6:0] _T_70613; // @[Modules.scala 143:103:@17122.4]
  wire [5:0] _T_70614; // @[Modules.scala 143:103:@17123.4]
  wire [5:0] _T_70615; // @[Modules.scala 143:103:@17124.4]
  wire [6:0] _T_70620; // @[Modules.scala 143:103:@17128.4]
  wire [5:0] _T_70621; // @[Modules.scala 143:103:@17129.4]
  wire [5:0] _T_70622; // @[Modules.scala 143:103:@17130.4]
  wire [4:0] _T_70626; // @[Modules.scala 144:80:@17133.4]
  wire [5:0] _T_70627; // @[Modules.scala 143:103:@17134.4]
  wire [4:0] _T_70628; // @[Modules.scala 143:103:@17135.4]
  wire [4:0] _T_70629; // @[Modules.scala 143:103:@17136.4]
  wire [5:0] _T_70634; // @[Modules.scala 143:103:@17140.4]
  wire [4:0] _T_70635; // @[Modules.scala 143:103:@17141.4]
  wire [4:0] _T_70636; // @[Modules.scala 143:103:@17142.4]
  wire [5:0] _T_70641; // @[Modules.scala 143:103:@17146.4]
  wire [4:0] _T_70642; // @[Modules.scala 143:103:@17147.4]
  wire [4:0] _T_70643; // @[Modules.scala 143:103:@17148.4]
  wire [5:0] _GEN_394; // @[Modules.scala 143:103:@17152.4]
  wire [6:0] _T_70648; // @[Modules.scala 143:103:@17152.4]
  wire [5:0] _T_70649; // @[Modules.scala 143:103:@17153.4]
  wire [5:0] _T_70650; // @[Modules.scala 143:103:@17154.4]
  wire [4:0] _T_70661; // @[Modules.scala 144:80:@17163.4]
  wire [5:0] _T_70662; // @[Modules.scala 143:103:@17164.4]
  wire [4:0] _T_70663; // @[Modules.scala 143:103:@17165.4]
  wire [4:0] _T_70664; // @[Modules.scala 143:103:@17166.4]
  wire [4:0] _T_70666; // @[Modules.scala 143:74:@17168.4]
  wire [5:0] _GEN_395; // @[Modules.scala 143:103:@17170.4]
  wire [6:0] _T_70669; // @[Modules.scala 143:103:@17170.4]
  wire [5:0] _T_70670; // @[Modules.scala 143:103:@17171.4]
  wire [5:0] _T_70671; // @[Modules.scala 143:103:@17172.4]
  wire [6:0] _T_70704; // @[Modules.scala 143:103:@17200.4]
  wire [5:0] _T_70705; // @[Modules.scala 143:103:@17201.4]
  wire [5:0] _T_70706; // @[Modules.scala 143:103:@17202.4]
  wire [6:0] _T_70718; // @[Modules.scala 143:103:@17212.4]
  wire [5:0] _T_70719; // @[Modules.scala 143:103:@17213.4]
  wire [5:0] _T_70720; // @[Modules.scala 143:103:@17214.4]
  wire [6:0] _T_70725; // @[Modules.scala 143:103:@17218.4]
  wire [5:0] _T_70726; // @[Modules.scala 143:103:@17219.4]
  wire [5:0] _T_70727; // @[Modules.scala 143:103:@17220.4]
  wire [5:0] _GEN_400; // @[Modules.scala 143:103:@17224.4]
  wire [6:0] _T_70732; // @[Modules.scala 143:103:@17224.4]
  wire [5:0] _T_70733; // @[Modules.scala 143:103:@17225.4]
  wire [5:0] _T_70734; // @[Modules.scala 143:103:@17226.4]
  wire [5:0] _T_70739; // @[Modules.scala 143:103:@17230.4]
  wire [4:0] _T_70740; // @[Modules.scala 143:103:@17231.4]
  wire [4:0] _T_70741; // @[Modules.scala 143:103:@17232.4]
  wire [5:0] _GEN_402; // @[Modules.scala 143:103:@17248.4]
  wire [6:0] _T_70760; // @[Modules.scala 143:103:@17248.4]
  wire [5:0] _T_70761; // @[Modules.scala 143:103:@17249.4]
  wire [5:0] _T_70762; // @[Modules.scala 143:103:@17250.4]
  wire [5:0] _T_70766; // @[Modules.scala 144:80:@17253.4]
  wire [6:0] _T_70767; // @[Modules.scala 143:103:@17254.4]
  wire [5:0] _T_70768; // @[Modules.scala 143:103:@17255.4]
  wire [5:0] _T_70769; // @[Modules.scala 143:103:@17256.4]
  wire [4:0] _T_70780; // @[Modules.scala 144:80:@17265.4]
  wire [5:0] _GEN_404; // @[Modules.scala 143:103:@17266.4]
  wire [6:0] _T_70781; // @[Modules.scala 143:103:@17266.4]
  wire [5:0] _T_70782; // @[Modules.scala 143:103:@17267.4]
  wire [5:0] _T_70783; // @[Modules.scala 143:103:@17268.4]
  wire [5:0] _T_70799; // @[Modules.scala 143:74:@17282.4]
  wire [6:0] _T_70802; // @[Modules.scala 143:103:@17284.4]
  wire [5:0] _T_70803; // @[Modules.scala 143:103:@17285.4]
  wire [5:0] _T_70804; // @[Modules.scala 143:103:@17286.4]
  wire [5:0] _T_70809; // @[Modules.scala 143:103:@17290.4]
  wire [4:0] _T_70810; // @[Modules.scala 143:103:@17291.4]
  wire [4:0] _T_70811; // @[Modules.scala 143:103:@17292.4]
  wire [4:0] _T_70815; // @[Modules.scala 144:80:@17295.4]
  wire [5:0] _T_70816; // @[Modules.scala 143:103:@17296.4]
  wire [4:0] _T_70817; // @[Modules.scala 143:103:@17297.4]
  wire [4:0] _T_70818; // @[Modules.scala 143:103:@17298.4]
  wire [5:0] _T_70829; // @[Modules.scala 144:80:@17307.4]
  wire [6:0] _T_70830; // @[Modules.scala 143:103:@17308.4]
  wire [5:0] _T_70831; // @[Modules.scala 143:103:@17309.4]
  wire [5:0] _T_70832; // @[Modules.scala 143:103:@17310.4]
  wire [6:0] _T_70837; // @[Modules.scala 143:103:@17314.4]
  wire [5:0] _T_70838; // @[Modules.scala 143:103:@17315.4]
  wire [5:0] _T_70839; // @[Modules.scala 143:103:@17316.4]
  wire [6:0] _T_70844; // @[Modules.scala 143:103:@17320.4]
  wire [5:0] _T_70845; // @[Modules.scala 143:103:@17321.4]
  wire [5:0] _T_70846; // @[Modules.scala 143:103:@17322.4]
  wire [4:0] _T_70855; // @[Modules.scala 143:74:@17330.4]
  wire [5:0] _GEN_406; // @[Modules.scala 143:103:@17332.4]
  wire [6:0] _T_70858; // @[Modules.scala 143:103:@17332.4]
  wire [5:0] _T_70859; // @[Modules.scala 143:103:@17333.4]
  wire [5:0] _T_70860; // @[Modules.scala 143:103:@17334.4]
  wire [6:0] _T_70872; // @[Modules.scala 143:103:@17344.4]
  wire [5:0] _T_70873; // @[Modules.scala 143:103:@17345.4]
  wire [5:0] _T_70874; // @[Modules.scala 143:103:@17346.4]
  wire [5:0] _T_70876; // @[Modules.scala 143:74:@17348.4]
  wire [6:0] _T_70879; // @[Modules.scala 143:103:@17350.4]
  wire [5:0] _T_70880; // @[Modules.scala 143:103:@17351.4]
  wire [5:0] _T_70881; // @[Modules.scala 143:103:@17352.4]
  wire [4:0] _T_70897; // @[Modules.scala 143:74:@17366.4]
  wire [5:0] _GEN_408; // @[Modules.scala 143:103:@17368.4]
  wire [6:0] _T_70900; // @[Modules.scala 143:103:@17368.4]
  wire [5:0] _T_70901; // @[Modules.scala 143:103:@17369.4]
  wire [5:0] _T_70902; // @[Modules.scala 143:103:@17370.4]
  wire [5:0] _T_70904; // @[Modules.scala 143:74:@17372.4]
  wire [6:0] _T_70907; // @[Modules.scala 143:103:@17374.4]
  wire [5:0] _T_70908; // @[Modules.scala 143:103:@17375.4]
  wire [5:0] _T_70909; // @[Modules.scala 143:103:@17376.4]
  wire [5:0] _T_70911; // @[Modules.scala 143:74:@17378.4]
  wire [5:0] _GEN_409; // @[Modules.scala 143:103:@17380.4]
  wire [6:0] _T_70914; // @[Modules.scala 143:103:@17380.4]
  wire [5:0] _T_70915; // @[Modules.scala 143:103:@17381.4]
  wire [5:0] _T_70916; // @[Modules.scala 143:103:@17382.4]
  wire [5:0] _T_70918; // @[Modules.scala 143:74:@17384.4]
  wire [6:0] _T_70921; // @[Modules.scala 143:103:@17386.4]
  wire [5:0] _T_70922; // @[Modules.scala 143:103:@17387.4]
  wire [5:0] _T_70923; // @[Modules.scala 143:103:@17388.4]
  wire [6:0] _T_70928; // @[Modules.scala 143:103:@17392.4]
  wire [5:0] _T_70929; // @[Modules.scala 143:103:@17393.4]
  wire [5:0] _T_70930; // @[Modules.scala 143:103:@17394.4]
  wire [6:0] _T_70935; // @[Modules.scala 143:103:@17398.4]
  wire [5:0] _T_70936; // @[Modules.scala 143:103:@17399.4]
  wire [5:0] _T_70937; // @[Modules.scala 143:103:@17400.4]
  wire [5:0] _T_70960; // @[Modules.scala 143:74:@17420.4]
  wire [6:0] _T_70963; // @[Modules.scala 143:103:@17422.4]
  wire [5:0] _T_70964; // @[Modules.scala 143:103:@17423.4]
  wire [5:0] _T_70965; // @[Modules.scala 143:103:@17424.4]
  wire [5:0] _GEN_411; // @[Modules.scala 143:103:@17428.4]
  wire [6:0] _T_70970; // @[Modules.scala 143:103:@17428.4]
  wire [5:0] _T_70971; // @[Modules.scala 143:103:@17429.4]
  wire [5:0] _T_70972; // @[Modules.scala 143:103:@17430.4]
  wire [5:0] _T_70977; // @[Modules.scala 143:103:@17434.4]
  wire [4:0] _T_70978; // @[Modules.scala 143:103:@17435.4]
  wire [4:0] _T_70979; // @[Modules.scala 143:103:@17436.4]
  wire [5:0] _T_70984; // @[Modules.scala 143:103:@17440.4]
  wire [4:0] _T_70985; // @[Modules.scala 143:103:@17441.4]
  wire [4:0] _T_70986; // @[Modules.scala 143:103:@17442.4]
  wire [5:0] _T_70990; // @[Modules.scala 144:80:@17445.4]
  wire [6:0] _T_70991; // @[Modules.scala 143:103:@17446.4]
  wire [5:0] _T_70992; // @[Modules.scala 143:103:@17447.4]
  wire [5:0] _T_70993; // @[Modules.scala 143:103:@17448.4]
  wire [5:0] _T_71002; // @[Modules.scala 143:74:@17456.4]
  wire [5:0] _T_71004; // @[Modules.scala 144:80:@17457.4]
  wire [6:0] _T_71005; // @[Modules.scala 143:103:@17458.4]
  wire [5:0] _T_71006; // @[Modules.scala 143:103:@17459.4]
  wire [5:0] _T_71007; // @[Modules.scala 143:103:@17460.4]
  wire [5:0] _T_71009; // @[Modules.scala 143:74:@17462.4]
  wire [6:0] _T_71012; // @[Modules.scala 143:103:@17464.4]
  wire [5:0] _T_71013; // @[Modules.scala 143:103:@17465.4]
  wire [5:0] _T_71014; // @[Modules.scala 143:103:@17466.4]
  wire [5:0] _T_71026; // @[Modules.scala 143:103:@17476.4]
  wire [4:0] _T_71027; // @[Modules.scala 143:103:@17477.4]
  wire [4:0] _T_71028; // @[Modules.scala 143:103:@17478.4]
  wire [6:0] _T_71040; // @[Modules.scala 143:103:@17488.4]
  wire [5:0] _T_71041; // @[Modules.scala 143:103:@17489.4]
  wire [5:0] _T_71042; // @[Modules.scala 143:103:@17490.4]
  wire [6:0] _T_71047; // @[Modules.scala 143:103:@17494.4]
  wire [5:0] _T_71048; // @[Modules.scala 143:103:@17495.4]
  wire [5:0] _T_71049; // @[Modules.scala 143:103:@17496.4]
  wire [5:0] _GEN_414; // @[Modules.scala 143:103:@17506.4]
  wire [6:0] _T_71061; // @[Modules.scala 143:103:@17506.4]
  wire [5:0] _T_71062; // @[Modules.scala 143:103:@17507.4]
  wire [5:0] _T_71063; // @[Modules.scala 143:103:@17508.4]
  wire [5:0] _T_71068; // @[Modules.scala 143:103:@17512.4]
  wire [4:0] _T_71069; // @[Modules.scala 143:103:@17513.4]
  wire [4:0] _T_71070; // @[Modules.scala 143:103:@17514.4]
  wire [5:0] _T_71075; // @[Modules.scala 143:103:@17518.4]
  wire [4:0] _T_71076; // @[Modules.scala 143:103:@17519.4]
  wire [4:0] _T_71077; // @[Modules.scala 143:103:@17520.4]
  wire [6:0] _T_71082; // @[Modules.scala 143:103:@17524.4]
  wire [5:0] _T_71083; // @[Modules.scala 143:103:@17525.4]
  wire [5:0] _T_71084; // @[Modules.scala 143:103:@17526.4]
  wire [5:0] _T_71088; // @[Modules.scala 144:80:@17529.4]
  wire [6:0] _T_71089; // @[Modules.scala 143:103:@17530.4]
  wire [5:0] _T_71090; // @[Modules.scala 143:103:@17531.4]
  wire [5:0] _T_71091; // @[Modules.scala 143:103:@17532.4]
  wire [6:0] _T_71096; // @[Modules.scala 143:103:@17536.4]
  wire [5:0] _T_71097; // @[Modules.scala 143:103:@17537.4]
  wire [5:0] _T_71098; // @[Modules.scala 143:103:@17538.4]
  wire [4:0] _T_71116; // @[Modules.scala 144:80:@17553.4]
  wire [5:0] _GEN_416; // @[Modules.scala 143:103:@17554.4]
  wire [6:0] _T_71117; // @[Modules.scala 143:103:@17554.4]
  wire [5:0] _T_71118; // @[Modules.scala 143:103:@17555.4]
  wire [5:0] _T_71119; // @[Modules.scala 143:103:@17556.4]
  wire [6:0] _T_71124; // @[Modules.scala 143:103:@17560.4]
  wire [5:0] _T_71125; // @[Modules.scala 143:103:@17561.4]
  wire [5:0] _T_71126; // @[Modules.scala 143:103:@17562.4]
  wire [6:0] _T_71131; // @[Modules.scala 143:103:@17566.4]
  wire [5:0] _T_71132; // @[Modules.scala 143:103:@17567.4]
  wire [5:0] _T_71133; // @[Modules.scala 143:103:@17568.4]
  wire [5:0] _T_71137; // @[Modules.scala 144:80:@17571.4]
  wire [6:0] _T_71138; // @[Modules.scala 143:103:@17572.4]
  wire [5:0] _T_71139; // @[Modules.scala 143:103:@17573.4]
  wire [5:0] _T_71140; // @[Modules.scala 143:103:@17574.4]
  wire [5:0] _GEN_417; // @[Modules.scala 143:103:@17578.4]
  wire [6:0] _T_71145; // @[Modules.scala 143:103:@17578.4]
  wire [5:0] _T_71146; // @[Modules.scala 143:103:@17579.4]
  wire [5:0] _T_71147; // @[Modules.scala 143:103:@17580.4]
  wire [4:0] _T_71151; // @[Modules.scala 144:80:@17583.4]
  wire [5:0] _T_71152; // @[Modules.scala 143:103:@17584.4]
  wire [4:0] _T_71153; // @[Modules.scala 143:103:@17585.4]
  wire [4:0] _T_71154; // @[Modules.scala 143:103:@17586.4]
  wire [5:0] _T_71159; // @[Modules.scala 143:103:@17590.4]
  wire [4:0] _T_71160; // @[Modules.scala 143:103:@17591.4]
  wire [4:0] _T_71161; // @[Modules.scala 143:103:@17592.4]
  wire [4:0] _T_71163; // @[Modules.scala 143:74:@17594.4]
  wire [5:0] _T_71166; // @[Modules.scala 143:103:@17596.4]
  wire [4:0] _T_71167; // @[Modules.scala 143:103:@17597.4]
  wire [4:0] _T_71168; // @[Modules.scala 143:103:@17598.4]
  wire [5:0] _T_71173; // @[Modules.scala 143:103:@17602.4]
  wire [4:0] _T_71174; // @[Modules.scala 143:103:@17603.4]
  wire [4:0] _T_71175; // @[Modules.scala 143:103:@17604.4]
  wire [5:0] _T_71179; // @[Modules.scala 144:80:@17607.4]
  wire [6:0] _T_71180; // @[Modules.scala 143:103:@17608.4]
  wire [5:0] _T_71181; // @[Modules.scala 143:103:@17609.4]
  wire [5:0] _T_71182; // @[Modules.scala 143:103:@17610.4]
  wire [6:0] _T_71187; // @[Modules.scala 143:103:@17614.4]
  wire [5:0] _T_71188; // @[Modules.scala 143:103:@17615.4]
  wire [5:0] _T_71189; // @[Modules.scala 143:103:@17616.4]
  wire [6:0] _T_71194; // @[Modules.scala 143:103:@17620.4]
  wire [5:0] _T_71195; // @[Modules.scala 143:103:@17621.4]
  wire [5:0] _T_71196; // @[Modules.scala 143:103:@17622.4]
  wire [5:0] _T_71201; // @[Modules.scala 143:103:@17626.4]
  wire [4:0] _T_71202; // @[Modules.scala 143:103:@17627.4]
  wire [4:0] _T_71203; // @[Modules.scala 143:103:@17628.4]
  wire [6:0] _T_71208; // @[Modules.scala 143:103:@17632.4]
  wire [5:0] _T_71209; // @[Modules.scala 143:103:@17633.4]
  wire [5:0] _T_71210; // @[Modules.scala 143:103:@17634.4]
  wire [5:0] _T_71221; // @[Modules.scala 144:80:@17643.4]
  wire [5:0] _GEN_418; // @[Modules.scala 143:103:@17644.4]
  wire [6:0] _T_71222; // @[Modules.scala 143:103:@17644.4]
  wire [5:0] _T_71223; // @[Modules.scala 143:103:@17645.4]
  wire [5:0] _T_71224; // @[Modules.scala 143:103:@17646.4]
  wire [5:0] _T_71235; // @[Modules.scala 144:80:@17655.4]
  wire [6:0] _T_71236; // @[Modules.scala 143:103:@17656.4]
  wire [5:0] _T_71237; // @[Modules.scala 143:103:@17657.4]
  wire [5:0] _T_71238; // @[Modules.scala 143:103:@17658.4]
  wire [5:0] _T_71240; // @[Modules.scala 143:74:@17660.4]
  wire [5:0] _T_71242; // @[Modules.scala 144:80:@17661.4]
  wire [6:0] _T_71243; // @[Modules.scala 143:103:@17662.4]
  wire [5:0] _T_71244; // @[Modules.scala 143:103:@17663.4]
  wire [5:0] _T_71245; // @[Modules.scala 143:103:@17664.4]
  wire [5:0] _T_71247; // @[Modules.scala 143:74:@17666.4]
  wire [6:0] _T_71250; // @[Modules.scala 143:103:@17668.4]
  wire [5:0] _T_71251; // @[Modules.scala 143:103:@17669.4]
  wire [5:0] _T_71252; // @[Modules.scala 143:103:@17670.4]
  wire [5:0] _GEN_419; // @[Modules.scala 143:103:@17674.4]
  wire [6:0] _T_71257; // @[Modules.scala 143:103:@17674.4]
  wire [5:0] _T_71258; // @[Modules.scala 143:103:@17675.4]
  wire [5:0] _T_71259; // @[Modules.scala 143:103:@17676.4]
  wire [6:0] _T_71264; // @[Modules.scala 143:103:@17680.4]
  wire [5:0] _T_71265; // @[Modules.scala 143:103:@17681.4]
  wire [5:0] _T_71266; // @[Modules.scala 143:103:@17682.4]
  wire [6:0] _T_71271; // @[Modules.scala 143:103:@17686.4]
  wire [5:0] _T_71272; // @[Modules.scala 143:103:@17687.4]
  wire [5:0] _T_71273; // @[Modules.scala 143:103:@17688.4]
  wire [5:0] _T_71278; // @[Modules.scala 143:103:@17692.4]
  wire [4:0] _T_71279; // @[Modules.scala 143:103:@17693.4]
  wire [4:0] _T_71280; // @[Modules.scala 143:103:@17694.4]
  wire [6:0] _T_71285; // @[Modules.scala 143:103:@17698.4]
  wire [5:0] _T_71286; // @[Modules.scala 143:103:@17699.4]
  wire [5:0] _T_71287; // @[Modules.scala 143:103:@17700.4]
  wire [5:0] _T_71299; // @[Modules.scala 143:103:@17710.4]
  wire [4:0] _T_71300; // @[Modules.scala 143:103:@17711.4]
  wire [4:0] _T_71301; // @[Modules.scala 143:103:@17712.4]
  wire [5:0] _T_71303; // @[Modules.scala 143:74:@17714.4]
  wire [6:0] _T_71306; // @[Modules.scala 143:103:@17716.4]
  wire [5:0] _T_71307; // @[Modules.scala 143:103:@17717.4]
  wire [5:0] _T_71308; // @[Modules.scala 143:103:@17718.4]
  wire [5:0] _T_71317; // @[Modules.scala 143:74:@17726.4]
  wire [6:0] _T_71320; // @[Modules.scala 143:103:@17728.4]
  wire [5:0] _T_71321; // @[Modules.scala 143:103:@17729.4]
  wire [5:0] _T_71322; // @[Modules.scala 143:103:@17730.4]
  wire [6:0] _T_71327; // @[Modules.scala 143:103:@17734.4]
  wire [5:0] _T_71328; // @[Modules.scala 143:103:@17735.4]
  wire [5:0] _T_71329; // @[Modules.scala 143:103:@17736.4]
  wire [6:0] _T_71334; // @[Modules.scala 143:103:@17740.4]
  wire [5:0] _T_71335; // @[Modules.scala 143:103:@17741.4]
  wire [5:0] _T_71336; // @[Modules.scala 143:103:@17742.4]
  wire [5:0] _T_71348; // @[Modules.scala 143:103:@17752.4]
  wire [4:0] _T_71349; // @[Modules.scala 143:103:@17753.4]
  wire [4:0] _T_71350; // @[Modules.scala 143:103:@17754.4]
  wire [4:0] _T_71354; // @[Modules.scala 144:80:@17757.4]
  wire [5:0] _T_71355; // @[Modules.scala 143:103:@17758.4]
  wire [4:0] _T_71356; // @[Modules.scala 143:103:@17759.4]
  wire [4:0] _T_71357; // @[Modules.scala 143:103:@17760.4]
  wire [6:0] _T_71362; // @[Modules.scala 143:103:@17764.4]
  wire [5:0] _T_71363; // @[Modules.scala 143:103:@17765.4]
  wire [5:0] _T_71364; // @[Modules.scala 143:103:@17766.4]
  wire [6:0] _T_71369; // @[Modules.scala 143:103:@17770.4]
  wire [5:0] _T_71370; // @[Modules.scala 143:103:@17771.4]
  wire [5:0] _T_71371; // @[Modules.scala 143:103:@17772.4]
  wire [6:0] _T_71383; // @[Modules.scala 143:103:@17782.4]
  wire [5:0] _T_71384; // @[Modules.scala 143:103:@17783.4]
  wire [5:0] _T_71385; // @[Modules.scala 143:103:@17784.4]
  wire [5:0] _T_71389; // @[Modules.scala 144:80:@17787.4]
  wire [6:0] _T_71390; // @[Modules.scala 143:103:@17788.4]
  wire [5:0] _T_71391; // @[Modules.scala 143:103:@17789.4]
  wire [5:0] _T_71392; // @[Modules.scala 143:103:@17790.4]
  wire [5:0] _T_71394; // @[Modules.scala 143:74:@17792.4]
  wire [5:0] _T_71396; // @[Modules.scala 144:80:@17793.4]
  wire [6:0] _T_71397; // @[Modules.scala 143:103:@17794.4]
  wire [5:0] _T_71398; // @[Modules.scala 143:103:@17795.4]
  wire [5:0] _T_71399; // @[Modules.scala 143:103:@17796.4]
  wire [6:0] _T_71404; // @[Modules.scala 143:103:@17800.4]
  wire [5:0] _T_71405; // @[Modules.scala 143:103:@17801.4]
  wire [5:0] _T_71406; // @[Modules.scala 143:103:@17802.4]
  wire [6:0] _T_71411; // @[Modules.scala 143:103:@17806.4]
  wire [5:0] _T_71412; // @[Modules.scala 143:103:@17807.4]
  wire [5:0] _T_71413; // @[Modules.scala 143:103:@17808.4]
  wire [5:0] _GEN_423; // @[Modules.scala 143:103:@17824.4]
  wire [6:0] _T_71432; // @[Modules.scala 143:103:@17824.4]
  wire [5:0] _T_71433; // @[Modules.scala 143:103:@17825.4]
  wire [5:0] _T_71434; // @[Modules.scala 143:103:@17826.4]
  wire [6:0] _T_71446; // @[Modules.scala 143:103:@17836.4]
  wire [5:0] _T_71447; // @[Modules.scala 143:103:@17837.4]
  wire [5:0] _T_71448; // @[Modules.scala 143:103:@17838.4]
  wire [6:0] _T_71509; // @[Modules.scala 143:103:@17890.4]
  wire [5:0] _T_71510; // @[Modules.scala 143:103:@17891.4]
  wire [5:0] _T_71511; // @[Modules.scala 143:103:@17892.4]
  wire [4:0] _T_71515; // @[Modules.scala 144:80:@17895.4]
  wire [5:0] _T_71516; // @[Modules.scala 143:103:@17896.4]
  wire [4:0] _T_71517; // @[Modules.scala 143:103:@17897.4]
  wire [4:0] _T_71518; // @[Modules.scala 143:103:@17898.4]
  wire [4:0] _T_71520; // @[Modules.scala 143:74:@17900.4]
  wire [5:0] _GEN_424; // @[Modules.scala 143:103:@17902.4]
  wire [6:0] _T_71523; // @[Modules.scala 143:103:@17902.4]
  wire [5:0] _T_71524; // @[Modules.scala 143:103:@17903.4]
  wire [5:0] _T_71525; // @[Modules.scala 143:103:@17904.4]
  wire [6:0] _T_71586; // @[Modules.scala 143:103:@17956.4]
  wire [5:0] _T_71587; // @[Modules.scala 143:103:@17957.4]
  wire [5:0] _T_71588; // @[Modules.scala 143:103:@17958.4]
  wire [6:0] _T_71593; // @[Modules.scala 143:103:@17962.4]
  wire [5:0] _T_71594; // @[Modules.scala 143:103:@17963.4]
  wire [5:0] _T_71595; // @[Modules.scala 143:103:@17964.4]
  wire [5:0] _T_71600; // @[Modules.scala 143:103:@17968.4]
  wire [4:0] _T_71601; // @[Modules.scala 143:103:@17969.4]
  wire [4:0] _T_71602; // @[Modules.scala 143:103:@17970.4]
  wire [6:0] _T_71607; // @[Modules.scala 143:103:@17974.4]
  wire [5:0] _T_71608; // @[Modules.scala 143:103:@17975.4]
  wire [5:0] _T_71609; // @[Modules.scala 143:103:@17976.4]
  wire [6:0] _T_71614; // @[Modules.scala 143:103:@17980.4]
  wire [5:0] _T_71615; // @[Modules.scala 143:103:@17981.4]
  wire [5:0] _T_71616; // @[Modules.scala 143:103:@17982.4]
  wire [6:0] _T_71621; // @[Modules.scala 143:103:@17986.4]
  wire [5:0] _T_71622; // @[Modules.scala 143:103:@17987.4]
  wire [5:0] _T_71623; // @[Modules.scala 143:103:@17988.4]
  wire [5:0] _T_71625; // @[Modules.scala 143:74:@17990.4]
  wire [6:0] _T_71628; // @[Modules.scala 143:103:@17992.4]
  wire [5:0] _T_71629; // @[Modules.scala 143:103:@17993.4]
  wire [5:0] _T_71630; // @[Modules.scala 143:103:@17994.4]
  wire [6:0] _T_71649; // @[Modules.scala 143:103:@18010.4]
  wire [5:0] _T_71650; // @[Modules.scala 143:103:@18011.4]
  wire [5:0] _T_71651; // @[Modules.scala 143:103:@18012.4]
  wire [5:0] _GEN_425; // @[Modules.scala 143:103:@18022.4]
  wire [6:0] _T_71663; // @[Modules.scala 143:103:@18022.4]
  wire [5:0] _T_71664; // @[Modules.scala 143:103:@18023.4]
  wire [5:0] _T_71665; // @[Modules.scala 143:103:@18024.4]
  wire [13:0] buffer_5_0; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71666; // @[Modules.scala 160:64:@18026.4]
  wire [13:0] _T_71667; // @[Modules.scala 160:64:@18027.4]
  wire [13:0] buffer_5_314; // @[Modules.scala 160:64:@18028.4]
  wire [14:0] _T_71669; // @[Modules.scala 160:64:@18030.4]
  wire [13:0] _T_71670; // @[Modules.scala 160:64:@18031.4]
  wire [13:0] buffer_5_315; // @[Modules.scala 160:64:@18032.4]
  wire [13:0] buffer_5_4; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71672; // @[Modules.scala 160:64:@18034.4]
  wire [13:0] _T_71673; // @[Modules.scala 160:64:@18035.4]
  wire [13:0] buffer_5_316; // @[Modules.scala 160:64:@18036.4]
  wire [13:0] buffer_5_6; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71675; // @[Modules.scala 160:64:@18038.4]
  wire [13:0] _T_71676; // @[Modules.scala 160:64:@18039.4]
  wire [13:0] buffer_5_317; // @[Modules.scala 160:64:@18040.4]
  wire [13:0] buffer_5_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71678; // @[Modules.scala 160:64:@18042.4]
  wire [13:0] _T_71679; // @[Modules.scala 160:64:@18043.4]
  wire [13:0] buffer_5_318; // @[Modules.scala 160:64:@18044.4]
  wire [13:0] buffer_5_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71681; // @[Modules.scala 160:64:@18046.4]
  wire [13:0] _T_71682; // @[Modules.scala 160:64:@18047.4]
  wire [13:0] buffer_5_319; // @[Modules.scala 160:64:@18048.4]
  wire [13:0] buffer_5_12; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71684; // @[Modules.scala 160:64:@18050.4]
  wire [13:0] _T_71685; // @[Modules.scala 160:64:@18051.4]
  wire [13:0] buffer_5_320; // @[Modules.scala 160:64:@18052.4]
  wire [13:0] buffer_5_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71696; // @[Modules.scala 160:64:@18066.4]
  wire [13:0] _T_71697; // @[Modules.scala 160:64:@18067.4]
  wire [13:0] buffer_5_324; // @[Modules.scala 160:64:@18068.4]
  wire [13:0] buffer_5_24; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71702; // @[Modules.scala 160:64:@18074.4]
  wire [13:0] _T_71703; // @[Modules.scala 160:64:@18075.4]
  wire [13:0] buffer_5_326; // @[Modules.scala 160:64:@18076.4]
  wire [13:0] buffer_5_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71705; // @[Modules.scala 160:64:@18078.4]
  wire [13:0] _T_71706; // @[Modules.scala 160:64:@18079.4]
  wire [13:0] buffer_5_327; // @[Modules.scala 160:64:@18080.4]
  wire [13:0] buffer_5_28; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71708; // @[Modules.scala 160:64:@18082.4]
  wire [13:0] _T_71709; // @[Modules.scala 160:64:@18083.4]
  wire [13:0] buffer_5_328; // @[Modules.scala 160:64:@18084.4]
  wire [13:0] buffer_5_32; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71714; // @[Modules.scala 160:64:@18090.4]
  wire [13:0] _T_71715; // @[Modules.scala 160:64:@18091.4]
  wire [13:0] buffer_5_330; // @[Modules.scala 160:64:@18092.4]
  wire [13:0] buffer_5_34; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71717; // @[Modules.scala 160:64:@18094.4]
  wire [13:0] _T_71718; // @[Modules.scala 160:64:@18095.4]
  wire [13:0] buffer_5_331; // @[Modules.scala 160:64:@18096.4]
  wire [13:0] buffer_5_36; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71720; // @[Modules.scala 160:64:@18098.4]
  wire [13:0] _T_71721; // @[Modules.scala 160:64:@18099.4]
  wire [13:0] buffer_5_332; // @[Modules.scala 160:64:@18100.4]
  wire [14:0] _T_71723; // @[Modules.scala 160:64:@18102.4]
  wire [13:0] _T_71724; // @[Modules.scala 160:64:@18103.4]
  wire [13:0] buffer_5_333; // @[Modules.scala 160:64:@18104.4]
  wire [13:0] buffer_5_40; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71726; // @[Modules.scala 160:64:@18106.4]
  wire [13:0] _T_71727; // @[Modules.scala 160:64:@18107.4]
  wire [13:0] buffer_5_334; // @[Modules.scala 160:64:@18108.4]
  wire [13:0] buffer_5_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71729; // @[Modules.scala 160:64:@18110.4]
  wire [13:0] _T_71730; // @[Modules.scala 160:64:@18111.4]
  wire [13:0] buffer_5_335; // @[Modules.scala 160:64:@18112.4]
  wire [13:0] buffer_5_44; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71732; // @[Modules.scala 160:64:@18114.4]
  wire [13:0] _T_71733; // @[Modules.scala 160:64:@18115.4]
  wire [13:0] buffer_5_336; // @[Modules.scala 160:64:@18116.4]
  wire [13:0] buffer_5_46; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71735; // @[Modules.scala 160:64:@18118.4]
  wire [13:0] _T_71736; // @[Modules.scala 160:64:@18119.4]
  wire [13:0] buffer_5_337; // @[Modules.scala 160:64:@18120.4]
  wire [13:0] buffer_5_50; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71741; // @[Modules.scala 160:64:@18126.4]
  wire [13:0] _T_71742; // @[Modules.scala 160:64:@18127.4]
  wire [13:0] buffer_5_339; // @[Modules.scala 160:64:@18128.4]
  wire [13:0] buffer_5_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71744; // @[Modules.scala 160:64:@18130.4]
  wire [13:0] _T_71745; // @[Modules.scala 160:64:@18131.4]
  wire [13:0] buffer_5_340; // @[Modules.scala 160:64:@18132.4]
  wire [13:0] buffer_5_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71747; // @[Modules.scala 160:64:@18134.4]
  wire [13:0] _T_71748; // @[Modules.scala 160:64:@18135.4]
  wire [13:0] buffer_5_341; // @[Modules.scala 160:64:@18136.4]
  wire [14:0] _T_71750; // @[Modules.scala 160:64:@18138.4]
  wire [13:0] _T_71751; // @[Modules.scala 160:64:@18139.4]
  wire [13:0] buffer_5_342; // @[Modules.scala 160:64:@18140.4]
  wire [13:0] buffer_5_58; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71753; // @[Modules.scala 160:64:@18142.4]
  wire [13:0] _T_71754; // @[Modules.scala 160:64:@18143.4]
  wire [13:0] buffer_5_343; // @[Modules.scala 160:64:@18144.4]
  wire [13:0] buffer_5_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71756; // @[Modules.scala 160:64:@18146.4]
  wire [13:0] _T_71757; // @[Modules.scala 160:64:@18147.4]
  wire [13:0] buffer_5_344; // @[Modules.scala 160:64:@18148.4]
  wire [13:0] buffer_5_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71759; // @[Modules.scala 160:64:@18150.4]
  wire [13:0] _T_71760; // @[Modules.scala 160:64:@18151.4]
  wire [13:0] buffer_5_345; // @[Modules.scala 160:64:@18152.4]
  wire [13:0] buffer_5_64; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_65; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71762; // @[Modules.scala 160:64:@18154.4]
  wire [13:0] _T_71763; // @[Modules.scala 160:64:@18155.4]
  wire [13:0] buffer_5_346; // @[Modules.scala 160:64:@18156.4]
  wire [13:0] buffer_5_66; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71765; // @[Modules.scala 160:64:@18158.4]
  wire [13:0] _T_71766; // @[Modules.scala 160:64:@18159.4]
  wire [13:0] buffer_5_347; // @[Modules.scala 160:64:@18160.4]
  wire [13:0] buffer_5_68; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71768; // @[Modules.scala 160:64:@18162.4]
  wire [13:0] _T_71769; // @[Modules.scala 160:64:@18163.4]
  wire [13:0] buffer_5_348; // @[Modules.scala 160:64:@18164.4]
  wire [13:0] buffer_5_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71771; // @[Modules.scala 160:64:@18166.4]
  wire [13:0] _T_71772; // @[Modules.scala 160:64:@18167.4]
  wire [13:0] buffer_5_349; // @[Modules.scala 160:64:@18168.4]
  wire [13:0] buffer_5_72; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71774; // @[Modules.scala 160:64:@18170.4]
  wire [13:0] _T_71775; // @[Modules.scala 160:64:@18171.4]
  wire [13:0] buffer_5_350; // @[Modules.scala 160:64:@18172.4]
  wire [13:0] buffer_5_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71780; // @[Modules.scala 160:64:@18178.4]
  wire [13:0] _T_71781; // @[Modules.scala 160:64:@18179.4]
  wire [13:0] buffer_5_352; // @[Modules.scala 160:64:@18180.4]
  wire [14:0] _T_71783; // @[Modules.scala 160:64:@18182.4]
  wire [13:0] _T_71784; // @[Modules.scala 160:64:@18183.4]
  wire [13:0] buffer_5_353; // @[Modules.scala 160:64:@18184.4]
  wire [13:0] buffer_5_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71786; // @[Modules.scala 160:64:@18186.4]
  wire [13:0] _T_71787; // @[Modules.scala 160:64:@18187.4]
  wire [13:0] buffer_5_354; // @[Modules.scala 160:64:@18188.4]
  wire [13:0] buffer_5_84; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71792; // @[Modules.scala 160:64:@18194.4]
  wire [13:0] _T_71793; // @[Modules.scala 160:64:@18195.4]
  wire [13:0] buffer_5_356; // @[Modules.scala 160:64:@18196.4]
  wire [13:0] buffer_5_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71801; // @[Modules.scala 160:64:@18206.4]
  wire [13:0] _T_71802; // @[Modules.scala 160:64:@18207.4]
  wire [13:0] buffer_5_359; // @[Modules.scala 160:64:@18208.4]
  wire [13:0] buffer_5_92; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71804; // @[Modules.scala 160:64:@18210.4]
  wire [13:0] _T_71805; // @[Modules.scala 160:64:@18211.4]
  wire [13:0] buffer_5_360; // @[Modules.scala 160:64:@18212.4]
  wire [13:0] buffer_5_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71807; // @[Modules.scala 160:64:@18214.4]
  wire [13:0] _T_71808; // @[Modules.scala 160:64:@18215.4]
  wire [13:0] buffer_5_361; // @[Modules.scala 160:64:@18216.4]
  wire [13:0] buffer_5_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71810; // @[Modules.scala 160:64:@18218.4]
  wire [13:0] _T_71811; // @[Modules.scala 160:64:@18219.4]
  wire [13:0] buffer_5_362; // @[Modules.scala 160:64:@18220.4]
  wire [13:0] buffer_5_98; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71813; // @[Modules.scala 160:64:@18222.4]
  wire [13:0] _T_71814; // @[Modules.scala 160:64:@18223.4]
  wire [13:0] buffer_5_363; // @[Modules.scala 160:64:@18224.4]
  wire [13:0] buffer_5_102; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_103; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71819; // @[Modules.scala 160:64:@18230.4]
  wire [13:0] _T_71820; // @[Modules.scala 160:64:@18231.4]
  wire [13:0] buffer_5_365; // @[Modules.scala 160:64:@18232.4]
  wire [13:0] buffer_5_104; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71822; // @[Modules.scala 160:64:@18234.4]
  wire [13:0] _T_71823; // @[Modules.scala 160:64:@18235.4]
  wire [13:0] buffer_5_366; // @[Modules.scala 160:64:@18236.4]
  wire [13:0] buffer_5_106; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71825; // @[Modules.scala 160:64:@18238.4]
  wire [13:0] _T_71826; // @[Modules.scala 160:64:@18239.4]
  wire [13:0] buffer_5_367; // @[Modules.scala 160:64:@18240.4]
  wire [13:0] buffer_5_109; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71828; // @[Modules.scala 160:64:@18242.4]
  wire [13:0] _T_71829; // @[Modules.scala 160:64:@18243.4]
  wire [13:0] buffer_5_368; // @[Modules.scala 160:64:@18244.4]
  wire [13:0] buffer_5_110; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71831; // @[Modules.scala 160:64:@18246.4]
  wire [13:0] _T_71832; // @[Modules.scala 160:64:@18247.4]
  wire [13:0] buffer_5_369; // @[Modules.scala 160:64:@18248.4]
  wire [13:0] buffer_5_112; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71834; // @[Modules.scala 160:64:@18250.4]
  wire [13:0] _T_71835; // @[Modules.scala 160:64:@18251.4]
  wire [13:0] buffer_5_370; // @[Modules.scala 160:64:@18252.4]
  wire [13:0] buffer_5_114; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71837; // @[Modules.scala 160:64:@18254.4]
  wire [13:0] _T_71838; // @[Modules.scala 160:64:@18255.4]
  wire [13:0] buffer_5_371; // @[Modules.scala 160:64:@18256.4]
  wire [13:0] buffer_5_116; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71840; // @[Modules.scala 160:64:@18258.4]
  wire [13:0] _T_71841; // @[Modules.scala 160:64:@18259.4]
  wire [13:0] buffer_5_372; // @[Modules.scala 160:64:@18260.4]
  wire [13:0] buffer_5_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71846; // @[Modules.scala 160:64:@18266.4]
  wire [13:0] _T_71847; // @[Modules.scala 160:64:@18267.4]
  wire [13:0] buffer_5_374; // @[Modules.scala 160:64:@18268.4]
  wire [13:0] buffer_5_122; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71849; // @[Modules.scala 160:64:@18270.4]
  wire [13:0] _T_71850; // @[Modules.scala 160:64:@18271.4]
  wire [13:0] buffer_5_375; // @[Modules.scala 160:64:@18272.4]
  wire [13:0] buffer_5_124; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71852; // @[Modules.scala 160:64:@18274.4]
  wire [13:0] _T_71853; // @[Modules.scala 160:64:@18275.4]
  wire [13:0] buffer_5_376; // @[Modules.scala 160:64:@18276.4]
  wire [13:0] buffer_5_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71855; // @[Modules.scala 160:64:@18278.4]
  wire [13:0] _T_71856; // @[Modules.scala 160:64:@18279.4]
  wire [13:0] buffer_5_377; // @[Modules.scala 160:64:@18280.4]
  wire [13:0] buffer_5_128; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71858; // @[Modules.scala 160:64:@18282.4]
  wire [13:0] _T_71859; // @[Modules.scala 160:64:@18283.4]
  wire [13:0] buffer_5_378; // @[Modules.scala 160:64:@18284.4]
  wire [13:0] buffer_5_130; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71861; // @[Modules.scala 160:64:@18286.4]
  wire [13:0] _T_71862; // @[Modules.scala 160:64:@18287.4]
  wire [13:0] buffer_5_379; // @[Modules.scala 160:64:@18288.4]
  wire [13:0] buffer_5_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71864; // @[Modules.scala 160:64:@18290.4]
  wire [13:0] _T_71865; // @[Modules.scala 160:64:@18291.4]
  wire [13:0] buffer_5_380; // @[Modules.scala 160:64:@18292.4]
  wire [13:0] buffer_5_134; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71867; // @[Modules.scala 160:64:@18294.4]
  wire [13:0] _T_71868; // @[Modules.scala 160:64:@18295.4]
  wire [13:0] buffer_5_381; // @[Modules.scala 160:64:@18296.4]
  wire [14:0] _T_71870; // @[Modules.scala 160:64:@18298.4]
  wire [13:0] _T_71871; // @[Modules.scala 160:64:@18299.4]
  wire [13:0] buffer_5_382; // @[Modules.scala 160:64:@18300.4]
  wire [14:0] _T_71876; // @[Modules.scala 160:64:@18306.4]
  wire [13:0] _T_71877; // @[Modules.scala 160:64:@18307.4]
  wire [13:0] buffer_5_384; // @[Modules.scala 160:64:@18308.4]
  wire [13:0] buffer_5_142; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_143; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71879; // @[Modules.scala 160:64:@18310.4]
  wire [13:0] _T_71880; // @[Modules.scala 160:64:@18311.4]
  wire [13:0] buffer_5_385; // @[Modules.scala 160:64:@18312.4]
  wire [13:0] buffer_5_144; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71882; // @[Modules.scala 160:64:@18314.4]
  wire [13:0] _T_71883; // @[Modules.scala 160:64:@18315.4]
  wire [13:0] buffer_5_386; // @[Modules.scala 160:64:@18316.4]
  wire [13:0] buffer_5_146; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71885; // @[Modules.scala 160:64:@18318.4]
  wire [13:0] _T_71886; // @[Modules.scala 160:64:@18319.4]
  wire [13:0] buffer_5_387; // @[Modules.scala 160:64:@18320.4]
  wire [13:0] buffer_5_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71888; // @[Modules.scala 160:64:@18322.4]
  wire [13:0] _T_71889; // @[Modules.scala 160:64:@18323.4]
  wire [13:0] buffer_5_388; // @[Modules.scala 160:64:@18324.4]
  wire [13:0] buffer_5_150; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71891; // @[Modules.scala 160:64:@18326.4]
  wire [13:0] _T_71892; // @[Modules.scala 160:64:@18327.4]
  wire [13:0] buffer_5_389; // @[Modules.scala 160:64:@18328.4]
  wire [13:0] buffer_5_152; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71894; // @[Modules.scala 160:64:@18330.4]
  wire [13:0] _T_71895; // @[Modules.scala 160:64:@18331.4]
  wire [13:0] buffer_5_390; // @[Modules.scala 160:64:@18332.4]
  wire [13:0] buffer_5_154; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71897; // @[Modules.scala 160:64:@18334.4]
  wire [13:0] _T_71898; // @[Modules.scala 160:64:@18335.4]
  wire [13:0] buffer_5_391; // @[Modules.scala 160:64:@18336.4]
  wire [13:0] buffer_5_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71900; // @[Modules.scala 160:64:@18338.4]
  wire [13:0] _T_71901; // @[Modules.scala 160:64:@18339.4]
  wire [13:0] buffer_5_392; // @[Modules.scala 160:64:@18340.4]
  wire [13:0] buffer_5_158; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71903; // @[Modules.scala 160:64:@18342.4]
  wire [13:0] _T_71904; // @[Modules.scala 160:64:@18343.4]
  wire [13:0] buffer_5_393; // @[Modules.scala 160:64:@18344.4]
  wire [13:0] buffer_5_160; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71906; // @[Modules.scala 160:64:@18346.4]
  wire [13:0] _T_71907; // @[Modules.scala 160:64:@18347.4]
  wire [13:0] buffer_5_394; // @[Modules.scala 160:64:@18348.4]
  wire [13:0] buffer_5_162; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_163; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71909; // @[Modules.scala 160:64:@18350.4]
  wire [13:0] _T_71910; // @[Modules.scala 160:64:@18351.4]
  wire [13:0] buffer_5_395; // @[Modules.scala 160:64:@18352.4]
  wire [13:0] buffer_5_164; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71912; // @[Modules.scala 160:64:@18354.4]
  wire [13:0] _T_71913; // @[Modules.scala 160:64:@18355.4]
  wire [13:0] buffer_5_396; // @[Modules.scala 160:64:@18356.4]
  wire [13:0] buffer_5_166; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71915; // @[Modules.scala 160:64:@18358.4]
  wire [13:0] _T_71916; // @[Modules.scala 160:64:@18359.4]
  wire [13:0] buffer_5_397; // @[Modules.scala 160:64:@18360.4]
  wire [13:0] buffer_5_168; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71918; // @[Modules.scala 160:64:@18362.4]
  wire [13:0] _T_71919; // @[Modules.scala 160:64:@18363.4]
  wire [13:0] buffer_5_398; // @[Modules.scala 160:64:@18364.4]
  wire [13:0] buffer_5_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71921; // @[Modules.scala 160:64:@18366.4]
  wire [13:0] _T_71922; // @[Modules.scala 160:64:@18367.4]
  wire [13:0] buffer_5_399; // @[Modules.scala 160:64:@18368.4]
  wire [13:0] buffer_5_176; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71930; // @[Modules.scala 160:64:@18378.4]
  wire [13:0] _T_71931; // @[Modules.scala 160:64:@18379.4]
  wire [13:0] buffer_5_402; // @[Modules.scala 160:64:@18380.4]
  wire [13:0] buffer_5_178; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_179; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71933; // @[Modules.scala 160:64:@18382.4]
  wire [13:0] _T_71934; // @[Modules.scala 160:64:@18383.4]
  wire [13:0] buffer_5_403; // @[Modules.scala 160:64:@18384.4]
  wire [13:0] buffer_5_180; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71936; // @[Modules.scala 160:64:@18386.4]
  wire [13:0] _T_71937; // @[Modules.scala 160:64:@18387.4]
  wire [13:0] buffer_5_404; // @[Modules.scala 160:64:@18388.4]
  wire [14:0] _T_71939; // @[Modules.scala 160:64:@18390.4]
  wire [13:0] _T_71940; // @[Modules.scala 160:64:@18391.4]
  wire [13:0] buffer_5_405; // @[Modules.scala 160:64:@18392.4]
  wire [13:0] buffer_5_184; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71942; // @[Modules.scala 160:64:@18394.4]
  wire [13:0] _T_71943; // @[Modules.scala 160:64:@18395.4]
  wire [13:0] buffer_5_406; // @[Modules.scala 160:64:@18396.4]
  wire [13:0] buffer_5_187; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71945; // @[Modules.scala 160:64:@18398.4]
  wire [13:0] _T_71946; // @[Modules.scala 160:64:@18399.4]
  wire [13:0] buffer_5_407; // @[Modules.scala 160:64:@18400.4]
  wire [13:0] buffer_5_190; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71951; // @[Modules.scala 160:64:@18406.4]
  wire [13:0] _T_71952; // @[Modules.scala 160:64:@18407.4]
  wire [13:0] buffer_5_409; // @[Modules.scala 160:64:@18408.4]
  wire [13:0] buffer_5_192; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71954; // @[Modules.scala 160:64:@18410.4]
  wire [13:0] _T_71955; // @[Modules.scala 160:64:@18411.4]
  wire [13:0] buffer_5_410; // @[Modules.scala 160:64:@18412.4]
  wire [13:0] buffer_5_194; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71957; // @[Modules.scala 160:64:@18414.4]
  wire [13:0] _T_71958; // @[Modules.scala 160:64:@18415.4]
  wire [13:0] buffer_5_411; // @[Modules.scala 160:64:@18416.4]
  wire [13:0] buffer_5_196; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71960; // @[Modules.scala 160:64:@18418.4]
  wire [13:0] _T_71961; // @[Modules.scala 160:64:@18419.4]
  wire [13:0] buffer_5_412; // @[Modules.scala 160:64:@18420.4]
  wire [13:0] buffer_5_198; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71963; // @[Modules.scala 160:64:@18422.4]
  wire [13:0] _T_71964; // @[Modules.scala 160:64:@18423.4]
  wire [13:0] buffer_5_413; // @[Modules.scala 160:64:@18424.4]
  wire [13:0] buffer_5_200; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71966; // @[Modules.scala 160:64:@18426.4]
  wire [13:0] _T_71967; // @[Modules.scala 160:64:@18427.4]
  wire [13:0] buffer_5_414; // @[Modules.scala 160:64:@18428.4]
  wire [14:0] _T_71969; // @[Modules.scala 160:64:@18430.4]
  wire [13:0] _T_71970; // @[Modules.scala 160:64:@18431.4]
  wire [13:0] buffer_5_415; // @[Modules.scala 160:64:@18432.4]
  wire [13:0] buffer_5_204; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71972; // @[Modules.scala 160:64:@18434.4]
  wire [13:0] _T_71973; // @[Modules.scala 160:64:@18435.4]
  wire [13:0] buffer_5_416; // @[Modules.scala 160:64:@18436.4]
  wire [13:0] buffer_5_206; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71975; // @[Modules.scala 160:64:@18438.4]
  wire [13:0] _T_71976; // @[Modules.scala 160:64:@18439.4]
  wire [13:0] buffer_5_417; // @[Modules.scala 160:64:@18440.4]
  wire [13:0] buffer_5_208; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_209; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71978; // @[Modules.scala 160:64:@18442.4]
  wire [13:0] _T_71979; // @[Modules.scala 160:64:@18443.4]
  wire [13:0] buffer_5_418; // @[Modules.scala 160:64:@18444.4]
  wire [14:0] _T_71981; // @[Modules.scala 160:64:@18446.4]
  wire [13:0] _T_71982; // @[Modules.scala 160:64:@18447.4]
  wire [13:0] buffer_5_419; // @[Modules.scala 160:64:@18448.4]
  wire [13:0] buffer_5_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71984; // @[Modules.scala 160:64:@18450.4]
  wire [13:0] _T_71985; // @[Modules.scala 160:64:@18451.4]
  wire [13:0] buffer_5_420; // @[Modules.scala 160:64:@18452.4]
  wire [13:0] buffer_5_214; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71987; // @[Modules.scala 160:64:@18454.4]
  wire [13:0] _T_71988; // @[Modules.scala 160:64:@18455.4]
  wire [13:0] buffer_5_421; // @[Modules.scala 160:64:@18456.4]
  wire [13:0] buffer_5_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71990; // @[Modules.scala 160:64:@18458.4]
  wire [13:0] _T_71991; // @[Modules.scala 160:64:@18459.4]
  wire [13:0] buffer_5_422; // @[Modules.scala 160:64:@18460.4]
  wire [13:0] buffer_5_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71993; // @[Modules.scala 160:64:@18462.4]
  wire [13:0] _T_71994; // @[Modules.scala 160:64:@18463.4]
  wire [13:0] buffer_5_423; // @[Modules.scala 160:64:@18464.4]
  wire [13:0] buffer_5_220; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71996; // @[Modules.scala 160:64:@18466.4]
  wire [13:0] _T_71997; // @[Modules.scala 160:64:@18467.4]
  wire [13:0] buffer_5_424; // @[Modules.scala 160:64:@18468.4]
  wire [13:0] buffer_5_222; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_71999; // @[Modules.scala 160:64:@18470.4]
  wire [13:0] _T_72000; // @[Modules.scala 160:64:@18471.4]
  wire [13:0] buffer_5_425; // @[Modules.scala 160:64:@18472.4]
  wire [13:0] buffer_5_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72002; // @[Modules.scala 160:64:@18474.4]
  wire [13:0] _T_72003; // @[Modules.scala 160:64:@18475.4]
  wire [13:0] buffer_5_426; // @[Modules.scala 160:64:@18476.4]
  wire [13:0] buffer_5_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72005; // @[Modules.scala 160:64:@18478.4]
  wire [13:0] _T_72006; // @[Modules.scala 160:64:@18479.4]
  wire [13:0] buffer_5_427; // @[Modules.scala 160:64:@18480.4]
  wire [13:0] buffer_5_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72008; // @[Modules.scala 160:64:@18482.4]
  wire [13:0] _T_72009; // @[Modules.scala 160:64:@18483.4]
  wire [13:0] buffer_5_428; // @[Modules.scala 160:64:@18484.4]
  wire [13:0] buffer_5_230; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72011; // @[Modules.scala 160:64:@18486.4]
  wire [13:0] _T_72012; // @[Modules.scala 160:64:@18487.4]
  wire [13:0] buffer_5_429; // @[Modules.scala 160:64:@18488.4]
  wire [13:0] buffer_5_232; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72014; // @[Modules.scala 160:64:@18490.4]
  wire [13:0] _T_72015; // @[Modules.scala 160:64:@18491.4]
  wire [13:0] buffer_5_430; // @[Modules.scala 160:64:@18492.4]
  wire [13:0] buffer_5_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72017; // @[Modules.scala 160:64:@18494.4]
  wire [13:0] _T_72018; // @[Modules.scala 160:64:@18495.4]
  wire [13:0] buffer_5_431; // @[Modules.scala 160:64:@18496.4]
  wire [13:0] buffer_5_236; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72020; // @[Modules.scala 160:64:@18498.4]
  wire [13:0] _T_72021; // @[Modules.scala 160:64:@18499.4]
  wire [13:0] buffer_5_432; // @[Modules.scala 160:64:@18500.4]
  wire [13:0] buffer_5_238; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72023; // @[Modules.scala 160:64:@18502.4]
  wire [13:0] _T_72024; // @[Modules.scala 160:64:@18503.4]
  wire [13:0] buffer_5_433; // @[Modules.scala 160:64:@18504.4]
  wire [13:0] buffer_5_240; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72026; // @[Modules.scala 160:64:@18506.4]
  wire [13:0] _T_72027; // @[Modules.scala 160:64:@18507.4]
  wire [13:0] buffer_5_434; // @[Modules.scala 160:64:@18508.4]
  wire [13:0] buffer_5_242; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72029; // @[Modules.scala 160:64:@18510.4]
  wire [13:0] _T_72030; // @[Modules.scala 160:64:@18511.4]
  wire [13:0] buffer_5_435; // @[Modules.scala 160:64:@18512.4]
  wire [13:0] buffer_5_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72032; // @[Modules.scala 160:64:@18514.4]
  wire [13:0] _T_72033; // @[Modules.scala 160:64:@18515.4]
  wire [13:0] buffer_5_436; // @[Modules.scala 160:64:@18516.4]
  wire [13:0] buffer_5_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72035; // @[Modules.scala 160:64:@18518.4]
  wire [13:0] _T_72036; // @[Modules.scala 160:64:@18519.4]
  wire [13:0] buffer_5_437; // @[Modules.scala 160:64:@18520.4]
  wire [13:0] buffer_5_248; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72038; // @[Modules.scala 160:64:@18522.4]
  wire [13:0] _T_72039; // @[Modules.scala 160:64:@18523.4]
  wire [13:0] buffer_5_438; // @[Modules.scala 160:64:@18524.4]
  wire [13:0] buffer_5_250; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72041; // @[Modules.scala 160:64:@18526.4]
  wire [13:0] _T_72042; // @[Modules.scala 160:64:@18527.4]
  wire [13:0] buffer_5_439; // @[Modules.scala 160:64:@18528.4]
  wire [13:0] buffer_5_252; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72044; // @[Modules.scala 160:64:@18530.4]
  wire [13:0] _T_72045; // @[Modules.scala 160:64:@18531.4]
  wire [13:0] buffer_5_440; // @[Modules.scala 160:64:@18532.4]
  wire [13:0] buffer_5_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72047; // @[Modules.scala 160:64:@18534.4]
  wire [13:0] _T_72048; // @[Modules.scala 160:64:@18535.4]
  wire [13:0] buffer_5_441; // @[Modules.scala 160:64:@18536.4]
  wire [13:0] buffer_5_256; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72050; // @[Modules.scala 160:64:@18538.4]
  wire [13:0] _T_72051; // @[Modules.scala 160:64:@18539.4]
  wire [13:0] buffer_5_442; // @[Modules.scala 160:64:@18540.4]
  wire [13:0] buffer_5_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72053; // @[Modules.scala 160:64:@18542.4]
  wire [13:0] _T_72054; // @[Modules.scala 160:64:@18543.4]
  wire [13:0] buffer_5_443; // @[Modules.scala 160:64:@18544.4]
  wire [13:0] buffer_5_261; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72056; // @[Modules.scala 160:64:@18546.4]
  wire [13:0] _T_72057; // @[Modules.scala 160:64:@18547.4]
  wire [13:0] buffer_5_444; // @[Modules.scala 160:64:@18548.4]
  wire [13:0] buffer_5_262; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72059; // @[Modules.scala 160:64:@18550.4]
  wire [13:0] _T_72060; // @[Modules.scala 160:64:@18551.4]
  wire [13:0] buffer_5_445; // @[Modules.scala 160:64:@18552.4]
  wire [13:0] buffer_5_264; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72062; // @[Modules.scala 160:64:@18554.4]
  wire [13:0] _T_72063; // @[Modules.scala 160:64:@18555.4]
  wire [13:0] buffer_5_446; // @[Modules.scala 160:64:@18556.4]
  wire [13:0] buffer_5_266; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72065; // @[Modules.scala 160:64:@18558.4]
  wire [13:0] _T_72066; // @[Modules.scala 160:64:@18559.4]
  wire [13:0] buffer_5_447; // @[Modules.scala 160:64:@18560.4]
  wire [13:0] buffer_5_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72068; // @[Modules.scala 160:64:@18562.4]
  wire [13:0] _T_72069; // @[Modules.scala 160:64:@18563.4]
  wire [13:0] buffer_5_448; // @[Modules.scala 160:64:@18564.4]
  wire [13:0] buffer_5_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72071; // @[Modules.scala 160:64:@18566.4]
  wire [13:0] _T_72072; // @[Modules.scala 160:64:@18567.4]
  wire [13:0] buffer_5_449; // @[Modules.scala 160:64:@18568.4]
  wire [13:0] buffer_5_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72074; // @[Modules.scala 160:64:@18570.4]
  wire [13:0] _T_72075; // @[Modules.scala 160:64:@18571.4]
  wire [13:0] buffer_5_450; // @[Modules.scala 160:64:@18572.4]
  wire [13:0] buffer_5_274; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_275; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72077; // @[Modules.scala 160:64:@18574.4]
  wire [13:0] _T_72078; // @[Modules.scala 160:64:@18575.4]
  wire [13:0] buffer_5_451; // @[Modules.scala 160:64:@18576.4]
  wire [13:0] buffer_5_276; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_277; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72080; // @[Modules.scala 160:64:@18578.4]
  wire [13:0] _T_72081; // @[Modules.scala 160:64:@18579.4]
  wire [13:0] buffer_5_452; // @[Modules.scala 160:64:@18580.4]
  wire [13:0] buffer_5_280; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72086; // @[Modules.scala 160:64:@18586.4]
  wire [13:0] _T_72087; // @[Modules.scala 160:64:@18587.4]
  wire [13:0] buffer_5_454; // @[Modules.scala 160:64:@18588.4]
  wire [13:0] buffer_5_282; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72089; // @[Modules.scala 160:64:@18590.4]
  wire [13:0] _T_72090; // @[Modules.scala 160:64:@18591.4]
  wire [13:0] buffer_5_455; // @[Modules.scala 160:64:@18592.4]
  wire [13:0] buffer_5_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72101; // @[Modules.scala 160:64:@18606.4]
  wire [13:0] _T_72102; // @[Modules.scala 160:64:@18607.4]
  wire [13:0] buffer_5_459; // @[Modules.scala 160:64:@18608.4]
  wire [13:0] buffer_5_292; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72104; // @[Modules.scala 160:64:@18610.4]
  wire [13:0] _T_72105; // @[Modules.scala 160:64:@18611.4]
  wire [13:0] buffer_5_460; // @[Modules.scala 160:64:@18612.4]
  wire [14:0] _T_72110; // @[Modules.scala 160:64:@18618.4]
  wire [13:0] _T_72111; // @[Modules.scala 160:64:@18619.4]
  wire [13:0] buffer_5_462; // @[Modules.scala 160:64:@18620.4]
  wire [13:0] buffer_5_302; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72119; // @[Modules.scala 160:64:@18630.4]
  wire [13:0] _T_72120; // @[Modules.scala 160:64:@18631.4]
  wire [13:0] buffer_5_465; // @[Modules.scala 160:64:@18632.4]
  wire [13:0] buffer_5_304; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_305; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72122; // @[Modules.scala 160:64:@18634.4]
  wire [13:0] _T_72123; // @[Modules.scala 160:64:@18635.4]
  wire [13:0] buffer_5_466; // @[Modules.scala 160:64:@18636.4]
  wire [13:0] buffer_5_306; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_5_307; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72125; // @[Modules.scala 160:64:@18638.4]
  wire [13:0] _T_72126; // @[Modules.scala 160:64:@18639.4]
  wire [13:0] buffer_5_467; // @[Modules.scala 160:64:@18640.4]
  wire [13:0] buffer_5_308; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72128; // @[Modules.scala 160:64:@18642.4]
  wire [13:0] _T_72129; // @[Modules.scala 160:64:@18643.4]
  wire [13:0] buffer_5_468; // @[Modules.scala 160:64:@18644.4]
  wire [13:0] buffer_5_311; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72131; // @[Modules.scala 160:64:@18646.4]
  wire [13:0] _T_72132; // @[Modules.scala 160:64:@18647.4]
  wire [13:0] buffer_5_469; // @[Modules.scala 160:64:@18648.4]
  wire [13:0] buffer_5_313; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_72134; // @[Modules.scala 160:64:@18650.4]
  wire [13:0] _T_72135; // @[Modules.scala 160:64:@18651.4]
  wire [13:0] buffer_5_470; // @[Modules.scala 160:64:@18652.4]
  wire [14:0] _T_72137; // @[Modules.scala 166:64:@18654.4]
  wire [13:0] _T_72138; // @[Modules.scala 166:64:@18655.4]
  wire [13:0] buffer_5_471; // @[Modules.scala 166:64:@18656.4]
  wire [14:0] _T_72140; // @[Modules.scala 166:64:@18658.4]
  wire [13:0] _T_72141; // @[Modules.scala 166:64:@18659.4]
  wire [13:0] buffer_5_472; // @[Modules.scala 166:64:@18660.4]
  wire [14:0] _T_72143; // @[Modules.scala 166:64:@18662.4]
  wire [13:0] _T_72144; // @[Modules.scala 166:64:@18663.4]
  wire [13:0] buffer_5_473; // @[Modules.scala 166:64:@18664.4]
  wire [14:0] _T_72146; // @[Modules.scala 166:64:@18666.4]
  wire [13:0] _T_72147; // @[Modules.scala 166:64:@18667.4]
  wire [13:0] buffer_5_474; // @[Modules.scala 166:64:@18668.4]
  wire [14:0] _T_72149; // @[Modules.scala 166:64:@18670.4]
  wire [13:0] _T_72150; // @[Modules.scala 166:64:@18671.4]
  wire [13:0] buffer_5_475; // @[Modules.scala 166:64:@18672.4]
  wire [14:0] _T_72152; // @[Modules.scala 166:64:@18674.4]
  wire [13:0] _T_72153; // @[Modules.scala 166:64:@18675.4]
  wire [13:0] buffer_5_476; // @[Modules.scala 166:64:@18676.4]
  wire [14:0] _T_72155; // @[Modules.scala 166:64:@18678.4]
  wire [13:0] _T_72156; // @[Modules.scala 166:64:@18679.4]
  wire [13:0] buffer_5_477; // @[Modules.scala 166:64:@18680.4]
  wire [14:0] _T_72158; // @[Modules.scala 166:64:@18682.4]
  wire [13:0] _T_72159; // @[Modules.scala 166:64:@18683.4]
  wire [13:0] buffer_5_478; // @[Modules.scala 166:64:@18684.4]
  wire [14:0] _T_72161; // @[Modules.scala 166:64:@18686.4]
  wire [13:0] _T_72162; // @[Modules.scala 166:64:@18687.4]
  wire [13:0] buffer_5_479; // @[Modules.scala 166:64:@18688.4]
  wire [14:0] _T_72164; // @[Modules.scala 166:64:@18690.4]
  wire [13:0] _T_72165; // @[Modules.scala 166:64:@18691.4]
  wire [13:0] buffer_5_480; // @[Modules.scala 166:64:@18692.4]
  wire [14:0] _T_72167; // @[Modules.scala 166:64:@18694.4]
  wire [13:0] _T_72168; // @[Modules.scala 166:64:@18695.4]
  wire [13:0] buffer_5_481; // @[Modules.scala 166:64:@18696.4]
  wire [14:0] _T_72170; // @[Modules.scala 166:64:@18698.4]
  wire [13:0] _T_72171; // @[Modules.scala 166:64:@18699.4]
  wire [13:0] buffer_5_482; // @[Modules.scala 166:64:@18700.4]
  wire [14:0] _T_72173; // @[Modules.scala 166:64:@18702.4]
  wire [13:0] _T_72174; // @[Modules.scala 166:64:@18703.4]
  wire [13:0] buffer_5_483; // @[Modules.scala 166:64:@18704.4]
  wire [14:0] _T_72176; // @[Modules.scala 166:64:@18706.4]
  wire [13:0] _T_72177; // @[Modules.scala 166:64:@18707.4]
  wire [13:0] buffer_5_484; // @[Modules.scala 166:64:@18708.4]
  wire [14:0] _T_72179; // @[Modules.scala 166:64:@18710.4]
  wire [13:0] _T_72180; // @[Modules.scala 166:64:@18711.4]
  wire [13:0] buffer_5_485; // @[Modules.scala 166:64:@18712.4]
  wire [14:0] _T_72182; // @[Modules.scala 166:64:@18714.4]
  wire [13:0] _T_72183; // @[Modules.scala 166:64:@18715.4]
  wire [13:0] buffer_5_486; // @[Modules.scala 166:64:@18716.4]
  wire [14:0] _T_72185; // @[Modules.scala 166:64:@18718.4]
  wire [13:0] _T_72186; // @[Modules.scala 166:64:@18719.4]
  wire [13:0] buffer_5_487; // @[Modules.scala 166:64:@18720.4]
  wire [14:0] _T_72188; // @[Modules.scala 166:64:@18722.4]
  wire [13:0] _T_72189; // @[Modules.scala 166:64:@18723.4]
  wire [13:0] buffer_5_488; // @[Modules.scala 166:64:@18724.4]
  wire [14:0] _T_72191; // @[Modules.scala 166:64:@18726.4]
  wire [13:0] _T_72192; // @[Modules.scala 166:64:@18727.4]
  wire [13:0] buffer_5_489; // @[Modules.scala 166:64:@18728.4]
  wire [14:0] _T_72194; // @[Modules.scala 166:64:@18730.4]
  wire [13:0] _T_72195; // @[Modules.scala 166:64:@18731.4]
  wire [13:0] buffer_5_490; // @[Modules.scala 166:64:@18732.4]
  wire [14:0] _T_72197; // @[Modules.scala 166:64:@18734.4]
  wire [13:0] _T_72198; // @[Modules.scala 166:64:@18735.4]
  wire [13:0] buffer_5_491; // @[Modules.scala 166:64:@18736.4]
  wire [14:0] _T_72200; // @[Modules.scala 166:64:@18738.4]
  wire [13:0] _T_72201; // @[Modules.scala 166:64:@18739.4]
  wire [13:0] buffer_5_492; // @[Modules.scala 166:64:@18740.4]
  wire [14:0] _T_72203; // @[Modules.scala 166:64:@18742.4]
  wire [13:0] _T_72204; // @[Modules.scala 166:64:@18743.4]
  wire [13:0] buffer_5_493; // @[Modules.scala 166:64:@18744.4]
  wire [14:0] _T_72206; // @[Modules.scala 166:64:@18746.4]
  wire [13:0] _T_72207; // @[Modules.scala 166:64:@18747.4]
  wire [13:0] buffer_5_494; // @[Modules.scala 166:64:@18748.4]
  wire [14:0] _T_72209; // @[Modules.scala 166:64:@18750.4]
  wire [13:0] _T_72210; // @[Modules.scala 166:64:@18751.4]
  wire [13:0] buffer_5_495; // @[Modules.scala 166:64:@18752.4]
  wire [14:0] _T_72212; // @[Modules.scala 166:64:@18754.4]
  wire [13:0] _T_72213; // @[Modules.scala 166:64:@18755.4]
  wire [13:0] buffer_5_496; // @[Modules.scala 166:64:@18756.4]
  wire [14:0] _T_72215; // @[Modules.scala 166:64:@18758.4]
  wire [13:0] _T_72216; // @[Modules.scala 166:64:@18759.4]
  wire [13:0] buffer_5_497; // @[Modules.scala 166:64:@18760.4]
  wire [14:0] _T_72218; // @[Modules.scala 166:64:@18762.4]
  wire [13:0] _T_72219; // @[Modules.scala 166:64:@18763.4]
  wire [13:0] buffer_5_498; // @[Modules.scala 166:64:@18764.4]
  wire [14:0] _T_72221; // @[Modules.scala 166:64:@18766.4]
  wire [13:0] _T_72222; // @[Modules.scala 166:64:@18767.4]
  wire [13:0] buffer_5_499; // @[Modules.scala 166:64:@18768.4]
  wire [14:0] _T_72224; // @[Modules.scala 166:64:@18770.4]
  wire [13:0] _T_72225; // @[Modules.scala 166:64:@18771.4]
  wire [13:0] buffer_5_500; // @[Modules.scala 166:64:@18772.4]
  wire [14:0] _T_72227; // @[Modules.scala 166:64:@18774.4]
  wire [13:0] _T_72228; // @[Modules.scala 166:64:@18775.4]
  wire [13:0] buffer_5_501; // @[Modules.scala 166:64:@18776.4]
  wire [14:0] _T_72230; // @[Modules.scala 166:64:@18778.4]
  wire [13:0] _T_72231; // @[Modules.scala 166:64:@18779.4]
  wire [13:0] buffer_5_502; // @[Modules.scala 166:64:@18780.4]
  wire [14:0] _T_72233; // @[Modules.scala 166:64:@18782.4]
  wire [13:0] _T_72234; // @[Modules.scala 166:64:@18783.4]
  wire [13:0] buffer_5_503; // @[Modules.scala 166:64:@18784.4]
  wire [14:0] _T_72236; // @[Modules.scala 166:64:@18786.4]
  wire [13:0] _T_72237; // @[Modules.scala 166:64:@18787.4]
  wire [13:0] buffer_5_504; // @[Modules.scala 166:64:@18788.4]
  wire [14:0] _T_72239; // @[Modules.scala 166:64:@18790.4]
  wire [13:0] _T_72240; // @[Modules.scala 166:64:@18791.4]
  wire [13:0] buffer_5_505; // @[Modules.scala 166:64:@18792.4]
  wire [14:0] _T_72242; // @[Modules.scala 166:64:@18794.4]
  wire [13:0] _T_72243; // @[Modules.scala 166:64:@18795.4]
  wire [13:0] buffer_5_506; // @[Modules.scala 166:64:@18796.4]
  wire [14:0] _T_72245; // @[Modules.scala 166:64:@18798.4]
  wire [13:0] _T_72246; // @[Modules.scala 166:64:@18799.4]
  wire [13:0] buffer_5_507; // @[Modules.scala 166:64:@18800.4]
  wire [14:0] _T_72248; // @[Modules.scala 166:64:@18802.4]
  wire [13:0] _T_72249; // @[Modules.scala 166:64:@18803.4]
  wire [13:0] buffer_5_508; // @[Modules.scala 166:64:@18804.4]
  wire [14:0] _T_72251; // @[Modules.scala 166:64:@18806.4]
  wire [13:0] _T_72252; // @[Modules.scala 166:64:@18807.4]
  wire [13:0] buffer_5_509; // @[Modules.scala 166:64:@18808.4]
  wire [14:0] _T_72254; // @[Modules.scala 166:64:@18810.4]
  wire [13:0] _T_72255; // @[Modules.scala 166:64:@18811.4]
  wire [13:0] buffer_5_510; // @[Modules.scala 166:64:@18812.4]
  wire [14:0] _T_72257; // @[Modules.scala 166:64:@18814.4]
  wire [13:0] _T_72258; // @[Modules.scala 166:64:@18815.4]
  wire [13:0] buffer_5_511; // @[Modules.scala 166:64:@18816.4]
  wire [14:0] _T_72260; // @[Modules.scala 166:64:@18818.4]
  wire [13:0] _T_72261; // @[Modules.scala 166:64:@18819.4]
  wire [13:0] buffer_5_512; // @[Modules.scala 166:64:@18820.4]
  wire [14:0] _T_72263; // @[Modules.scala 166:64:@18822.4]
  wire [13:0] _T_72264; // @[Modules.scala 166:64:@18823.4]
  wire [13:0] buffer_5_513; // @[Modules.scala 166:64:@18824.4]
  wire [14:0] _T_72266; // @[Modules.scala 166:64:@18826.4]
  wire [13:0] _T_72267; // @[Modules.scala 166:64:@18827.4]
  wire [13:0] buffer_5_514; // @[Modules.scala 166:64:@18828.4]
  wire [14:0] _T_72269; // @[Modules.scala 166:64:@18830.4]
  wire [13:0] _T_72270; // @[Modules.scala 166:64:@18831.4]
  wire [13:0] buffer_5_515; // @[Modules.scala 166:64:@18832.4]
  wire [14:0] _T_72272; // @[Modules.scala 166:64:@18834.4]
  wire [13:0] _T_72273; // @[Modules.scala 166:64:@18835.4]
  wire [13:0] buffer_5_516; // @[Modules.scala 166:64:@18836.4]
  wire [14:0] _T_72275; // @[Modules.scala 166:64:@18838.4]
  wire [13:0] _T_72276; // @[Modules.scala 166:64:@18839.4]
  wire [13:0] buffer_5_517; // @[Modules.scala 166:64:@18840.4]
  wire [14:0] _T_72278; // @[Modules.scala 166:64:@18842.4]
  wire [13:0] _T_72279; // @[Modules.scala 166:64:@18843.4]
  wire [13:0] buffer_5_518; // @[Modules.scala 166:64:@18844.4]
  wire [14:0] _T_72281; // @[Modules.scala 166:64:@18846.4]
  wire [13:0] _T_72282; // @[Modules.scala 166:64:@18847.4]
  wire [13:0] buffer_5_519; // @[Modules.scala 166:64:@18848.4]
  wire [14:0] _T_72284; // @[Modules.scala 166:64:@18850.4]
  wire [13:0] _T_72285; // @[Modules.scala 166:64:@18851.4]
  wire [13:0] buffer_5_520; // @[Modules.scala 166:64:@18852.4]
  wire [14:0] _T_72287; // @[Modules.scala 166:64:@18854.4]
  wire [13:0] _T_72288; // @[Modules.scala 166:64:@18855.4]
  wire [13:0] buffer_5_521; // @[Modules.scala 166:64:@18856.4]
  wire [14:0] _T_72290; // @[Modules.scala 166:64:@18858.4]
  wire [13:0] _T_72291; // @[Modules.scala 166:64:@18859.4]
  wire [13:0] buffer_5_522; // @[Modules.scala 166:64:@18860.4]
  wire [14:0] _T_72293; // @[Modules.scala 166:64:@18862.4]
  wire [13:0] _T_72294; // @[Modules.scala 166:64:@18863.4]
  wire [13:0] buffer_5_523; // @[Modules.scala 166:64:@18864.4]
  wire [14:0] _T_72296; // @[Modules.scala 166:64:@18866.4]
  wire [13:0] _T_72297; // @[Modules.scala 166:64:@18867.4]
  wire [13:0] buffer_5_524; // @[Modules.scala 166:64:@18868.4]
  wire [14:0] _T_72299; // @[Modules.scala 166:64:@18870.4]
  wire [13:0] _T_72300; // @[Modules.scala 166:64:@18871.4]
  wire [13:0] buffer_5_525; // @[Modules.scala 166:64:@18872.4]
  wire [14:0] _T_72302; // @[Modules.scala 166:64:@18874.4]
  wire [13:0] _T_72303; // @[Modules.scala 166:64:@18875.4]
  wire [13:0] buffer_5_526; // @[Modules.scala 166:64:@18876.4]
  wire [14:0] _T_72305; // @[Modules.scala 166:64:@18878.4]
  wire [13:0] _T_72306; // @[Modules.scala 166:64:@18879.4]
  wire [13:0] buffer_5_527; // @[Modules.scala 166:64:@18880.4]
  wire [14:0] _T_72308; // @[Modules.scala 166:64:@18882.4]
  wire [13:0] _T_72309; // @[Modules.scala 166:64:@18883.4]
  wire [13:0] buffer_5_528; // @[Modules.scala 166:64:@18884.4]
  wire [14:0] _T_72311; // @[Modules.scala 166:64:@18886.4]
  wire [13:0] _T_72312; // @[Modules.scala 166:64:@18887.4]
  wire [13:0] buffer_5_529; // @[Modules.scala 166:64:@18888.4]
  wire [14:0] _T_72314; // @[Modules.scala 166:64:@18890.4]
  wire [13:0] _T_72315; // @[Modules.scala 166:64:@18891.4]
  wire [13:0] buffer_5_530; // @[Modules.scala 166:64:@18892.4]
  wire [14:0] _T_72317; // @[Modules.scala 166:64:@18894.4]
  wire [13:0] _T_72318; // @[Modules.scala 166:64:@18895.4]
  wire [13:0] buffer_5_531; // @[Modules.scala 166:64:@18896.4]
  wire [14:0] _T_72320; // @[Modules.scala 166:64:@18898.4]
  wire [13:0] _T_72321; // @[Modules.scala 166:64:@18899.4]
  wire [13:0] buffer_5_532; // @[Modules.scala 166:64:@18900.4]
  wire [14:0] _T_72323; // @[Modules.scala 166:64:@18902.4]
  wire [13:0] _T_72324; // @[Modules.scala 166:64:@18903.4]
  wire [13:0] buffer_5_533; // @[Modules.scala 166:64:@18904.4]
  wire [14:0] _T_72326; // @[Modules.scala 166:64:@18906.4]
  wire [13:0] _T_72327; // @[Modules.scala 166:64:@18907.4]
  wire [13:0] buffer_5_534; // @[Modules.scala 166:64:@18908.4]
  wire [14:0] _T_72329; // @[Modules.scala 166:64:@18910.4]
  wire [13:0] _T_72330; // @[Modules.scala 166:64:@18911.4]
  wire [13:0] buffer_5_535; // @[Modules.scala 166:64:@18912.4]
  wire [14:0] _T_72332; // @[Modules.scala 166:64:@18914.4]
  wire [13:0] _T_72333; // @[Modules.scala 166:64:@18915.4]
  wire [13:0] buffer_5_536; // @[Modules.scala 166:64:@18916.4]
  wire [14:0] _T_72335; // @[Modules.scala 166:64:@18918.4]
  wire [13:0] _T_72336; // @[Modules.scala 166:64:@18919.4]
  wire [13:0] buffer_5_537; // @[Modules.scala 166:64:@18920.4]
  wire [14:0] _T_72338; // @[Modules.scala 166:64:@18922.4]
  wire [13:0] _T_72339; // @[Modules.scala 166:64:@18923.4]
  wire [13:0] buffer_5_538; // @[Modules.scala 166:64:@18924.4]
  wire [14:0] _T_72341; // @[Modules.scala 166:64:@18926.4]
  wire [13:0] _T_72342; // @[Modules.scala 166:64:@18927.4]
  wire [13:0] buffer_5_539; // @[Modules.scala 166:64:@18928.4]
  wire [14:0] _T_72344; // @[Modules.scala 166:64:@18930.4]
  wire [13:0] _T_72345; // @[Modules.scala 166:64:@18931.4]
  wire [13:0] buffer_5_540; // @[Modules.scala 166:64:@18932.4]
  wire [14:0] _T_72347; // @[Modules.scala 166:64:@18934.4]
  wire [13:0] _T_72348; // @[Modules.scala 166:64:@18935.4]
  wire [13:0] buffer_5_541; // @[Modules.scala 166:64:@18936.4]
  wire [14:0] _T_72350; // @[Modules.scala 166:64:@18938.4]
  wire [13:0] _T_72351; // @[Modules.scala 166:64:@18939.4]
  wire [13:0] buffer_5_542; // @[Modules.scala 166:64:@18940.4]
  wire [14:0] _T_72353; // @[Modules.scala 166:64:@18942.4]
  wire [13:0] _T_72354; // @[Modules.scala 166:64:@18943.4]
  wire [13:0] buffer_5_543; // @[Modules.scala 166:64:@18944.4]
  wire [14:0] _T_72356; // @[Modules.scala 166:64:@18946.4]
  wire [13:0] _T_72357; // @[Modules.scala 166:64:@18947.4]
  wire [13:0] buffer_5_544; // @[Modules.scala 166:64:@18948.4]
  wire [14:0] _T_72359; // @[Modules.scala 166:64:@18950.4]
  wire [13:0] _T_72360; // @[Modules.scala 166:64:@18951.4]
  wire [13:0] buffer_5_545; // @[Modules.scala 166:64:@18952.4]
  wire [14:0] _T_72362; // @[Modules.scala 166:64:@18954.4]
  wire [13:0] _T_72363; // @[Modules.scala 166:64:@18955.4]
  wire [13:0] buffer_5_546; // @[Modules.scala 166:64:@18956.4]
  wire [14:0] _T_72365; // @[Modules.scala 166:64:@18958.4]
  wire [13:0] _T_72366; // @[Modules.scala 166:64:@18959.4]
  wire [13:0] buffer_5_547; // @[Modules.scala 166:64:@18960.4]
  wire [14:0] _T_72368; // @[Modules.scala 166:64:@18962.4]
  wire [13:0] _T_72369; // @[Modules.scala 166:64:@18963.4]
  wire [13:0] buffer_5_548; // @[Modules.scala 166:64:@18964.4]
  wire [14:0] _T_72371; // @[Modules.scala 160:64:@18966.4]
  wire [13:0] _T_72372; // @[Modules.scala 160:64:@18967.4]
  wire [13:0] buffer_5_549; // @[Modules.scala 160:64:@18968.4]
  wire [14:0] _T_72374; // @[Modules.scala 160:64:@18970.4]
  wire [13:0] _T_72375; // @[Modules.scala 160:64:@18971.4]
  wire [13:0] buffer_5_550; // @[Modules.scala 160:64:@18972.4]
  wire [14:0] _T_72377; // @[Modules.scala 160:64:@18974.4]
  wire [13:0] _T_72378; // @[Modules.scala 160:64:@18975.4]
  wire [13:0] buffer_5_551; // @[Modules.scala 160:64:@18976.4]
  wire [14:0] _T_72380; // @[Modules.scala 160:64:@18978.4]
  wire [13:0] _T_72381; // @[Modules.scala 160:64:@18979.4]
  wire [13:0] buffer_5_552; // @[Modules.scala 160:64:@18980.4]
  wire [14:0] _T_72383; // @[Modules.scala 160:64:@18982.4]
  wire [13:0] _T_72384; // @[Modules.scala 160:64:@18983.4]
  wire [13:0] buffer_5_553; // @[Modules.scala 160:64:@18984.4]
  wire [14:0] _T_72386; // @[Modules.scala 160:64:@18986.4]
  wire [13:0] _T_72387; // @[Modules.scala 160:64:@18987.4]
  wire [13:0] buffer_5_554; // @[Modules.scala 160:64:@18988.4]
  wire [14:0] _T_72389; // @[Modules.scala 160:64:@18990.4]
  wire [13:0] _T_72390; // @[Modules.scala 160:64:@18991.4]
  wire [13:0] buffer_5_555; // @[Modules.scala 160:64:@18992.4]
  wire [14:0] _T_72392; // @[Modules.scala 160:64:@18994.4]
  wire [13:0] _T_72393; // @[Modules.scala 160:64:@18995.4]
  wire [13:0] buffer_5_556; // @[Modules.scala 160:64:@18996.4]
  wire [14:0] _T_72395; // @[Modules.scala 160:64:@18998.4]
  wire [13:0] _T_72396; // @[Modules.scala 160:64:@18999.4]
  wire [13:0] buffer_5_557; // @[Modules.scala 160:64:@19000.4]
  wire [14:0] _T_72398; // @[Modules.scala 160:64:@19002.4]
  wire [13:0] _T_72399; // @[Modules.scala 160:64:@19003.4]
  wire [13:0] buffer_5_558; // @[Modules.scala 160:64:@19004.4]
  wire [14:0] _T_72401; // @[Modules.scala 160:64:@19006.4]
  wire [13:0] _T_72402; // @[Modules.scala 160:64:@19007.4]
  wire [13:0] buffer_5_559; // @[Modules.scala 160:64:@19008.4]
  wire [14:0] _T_72404; // @[Modules.scala 160:64:@19010.4]
  wire [13:0] _T_72405; // @[Modules.scala 160:64:@19011.4]
  wire [13:0] buffer_5_560; // @[Modules.scala 160:64:@19012.4]
  wire [14:0] _T_72407; // @[Modules.scala 160:64:@19014.4]
  wire [13:0] _T_72408; // @[Modules.scala 160:64:@19015.4]
  wire [13:0] buffer_5_561; // @[Modules.scala 160:64:@19016.4]
  wire [14:0] _T_72410; // @[Modules.scala 160:64:@19018.4]
  wire [13:0] _T_72411; // @[Modules.scala 160:64:@19019.4]
  wire [13:0] buffer_5_562; // @[Modules.scala 160:64:@19020.4]
  wire [14:0] _T_72413; // @[Modules.scala 160:64:@19022.4]
  wire [13:0] _T_72414; // @[Modules.scala 160:64:@19023.4]
  wire [13:0] buffer_5_563; // @[Modules.scala 160:64:@19024.4]
  wire [14:0] _T_72416; // @[Modules.scala 160:64:@19026.4]
  wire [13:0] _T_72417; // @[Modules.scala 160:64:@19027.4]
  wire [13:0] buffer_5_564; // @[Modules.scala 160:64:@19028.4]
  wire [14:0] _T_72419; // @[Modules.scala 160:64:@19030.4]
  wire [13:0] _T_72420; // @[Modules.scala 160:64:@19031.4]
  wire [13:0] buffer_5_565; // @[Modules.scala 160:64:@19032.4]
  wire [14:0] _T_72422; // @[Modules.scala 160:64:@19034.4]
  wire [13:0] _T_72423; // @[Modules.scala 160:64:@19035.4]
  wire [13:0] buffer_5_566; // @[Modules.scala 160:64:@19036.4]
  wire [14:0] _T_72425; // @[Modules.scala 160:64:@19038.4]
  wire [13:0] _T_72426; // @[Modules.scala 160:64:@19039.4]
  wire [13:0] buffer_5_567; // @[Modules.scala 160:64:@19040.4]
  wire [14:0] _T_72428; // @[Modules.scala 160:64:@19042.4]
  wire [13:0] _T_72429; // @[Modules.scala 160:64:@19043.4]
  wire [13:0] buffer_5_568; // @[Modules.scala 160:64:@19044.4]
  wire [14:0] _T_72431; // @[Modules.scala 160:64:@19046.4]
  wire [13:0] _T_72432; // @[Modules.scala 160:64:@19047.4]
  wire [13:0] buffer_5_569; // @[Modules.scala 160:64:@19048.4]
  wire [14:0] _T_72434; // @[Modules.scala 160:64:@19050.4]
  wire [13:0] _T_72435; // @[Modules.scala 160:64:@19051.4]
  wire [13:0] buffer_5_570; // @[Modules.scala 160:64:@19052.4]
  wire [14:0] _T_72437; // @[Modules.scala 160:64:@19054.4]
  wire [13:0] _T_72438; // @[Modules.scala 160:64:@19055.4]
  wire [13:0] buffer_5_571; // @[Modules.scala 160:64:@19056.4]
  wire [14:0] _T_72440; // @[Modules.scala 160:64:@19058.4]
  wire [13:0] _T_72441; // @[Modules.scala 160:64:@19059.4]
  wire [13:0] buffer_5_572; // @[Modules.scala 160:64:@19060.4]
  wire [14:0] _T_72443; // @[Modules.scala 160:64:@19062.4]
  wire [13:0] _T_72444; // @[Modules.scala 160:64:@19063.4]
  wire [13:0] buffer_5_573; // @[Modules.scala 160:64:@19064.4]
  wire [14:0] _T_72446; // @[Modules.scala 160:64:@19066.4]
  wire [13:0] _T_72447; // @[Modules.scala 160:64:@19067.4]
  wire [13:0] buffer_5_574; // @[Modules.scala 160:64:@19068.4]
  wire [14:0] _T_72449; // @[Modules.scala 160:64:@19070.4]
  wire [13:0] _T_72450; // @[Modules.scala 160:64:@19071.4]
  wire [13:0] buffer_5_575; // @[Modules.scala 160:64:@19072.4]
  wire [14:0] _T_72452; // @[Modules.scala 160:64:@19074.4]
  wire [13:0] _T_72453; // @[Modules.scala 160:64:@19075.4]
  wire [13:0] buffer_5_576; // @[Modules.scala 160:64:@19076.4]
  wire [14:0] _T_72455; // @[Modules.scala 160:64:@19078.4]
  wire [13:0] _T_72456; // @[Modules.scala 160:64:@19079.4]
  wire [13:0] buffer_5_577; // @[Modules.scala 160:64:@19080.4]
  wire [14:0] _T_72458; // @[Modules.scala 160:64:@19082.4]
  wire [13:0] _T_72459; // @[Modules.scala 160:64:@19083.4]
  wire [13:0] buffer_5_578; // @[Modules.scala 160:64:@19084.4]
  wire [14:0] _T_72461; // @[Modules.scala 160:64:@19086.4]
  wire [13:0] _T_72462; // @[Modules.scala 160:64:@19087.4]
  wire [13:0] buffer_5_579; // @[Modules.scala 160:64:@19088.4]
  wire [14:0] _T_72464; // @[Modules.scala 160:64:@19090.4]
  wire [13:0] _T_72465; // @[Modules.scala 160:64:@19091.4]
  wire [13:0] buffer_5_580; // @[Modules.scala 160:64:@19092.4]
  wire [14:0] _T_72467; // @[Modules.scala 160:64:@19094.4]
  wire [13:0] _T_72468; // @[Modules.scala 160:64:@19095.4]
  wire [13:0] buffer_5_581; // @[Modules.scala 160:64:@19096.4]
  wire [14:0] _T_72470; // @[Modules.scala 160:64:@19098.4]
  wire [13:0] _T_72471; // @[Modules.scala 160:64:@19099.4]
  wire [13:0] buffer_5_582; // @[Modules.scala 160:64:@19100.4]
  wire [14:0] _T_72473; // @[Modules.scala 160:64:@19102.4]
  wire [13:0] _T_72474; // @[Modules.scala 160:64:@19103.4]
  wire [13:0] buffer_5_583; // @[Modules.scala 160:64:@19104.4]
  wire [14:0] _T_72476; // @[Modules.scala 160:64:@19106.4]
  wire [13:0] _T_72477; // @[Modules.scala 160:64:@19107.4]
  wire [13:0] buffer_5_584; // @[Modules.scala 160:64:@19108.4]
  wire [14:0] _T_72479; // @[Modules.scala 160:64:@19110.4]
  wire [13:0] _T_72480; // @[Modules.scala 160:64:@19111.4]
  wire [13:0] buffer_5_585; // @[Modules.scala 160:64:@19112.4]
  wire [14:0] _T_72482; // @[Modules.scala 160:64:@19114.4]
  wire [13:0] _T_72483; // @[Modules.scala 160:64:@19115.4]
  wire [13:0] buffer_5_586; // @[Modules.scala 160:64:@19116.4]
  wire [14:0] _T_72485; // @[Modules.scala 160:64:@19118.4]
  wire [13:0] _T_72486; // @[Modules.scala 160:64:@19119.4]
  wire [13:0] buffer_5_587; // @[Modules.scala 160:64:@19120.4]
  wire [14:0] _T_72488; // @[Modules.scala 166:64:@19122.4]
  wire [13:0] _T_72489; // @[Modules.scala 166:64:@19123.4]
  wire [13:0] buffer_5_588; // @[Modules.scala 166:64:@19124.4]
  wire [14:0] _T_72491; // @[Modules.scala 166:64:@19126.4]
  wire [13:0] _T_72492; // @[Modules.scala 166:64:@19127.4]
  wire [13:0] buffer_5_589; // @[Modules.scala 166:64:@19128.4]
  wire [14:0] _T_72494; // @[Modules.scala 166:64:@19130.4]
  wire [13:0] _T_72495; // @[Modules.scala 166:64:@19131.4]
  wire [13:0] buffer_5_590; // @[Modules.scala 166:64:@19132.4]
  wire [14:0] _T_72497; // @[Modules.scala 166:64:@19134.4]
  wire [13:0] _T_72498; // @[Modules.scala 166:64:@19135.4]
  wire [13:0] buffer_5_591; // @[Modules.scala 166:64:@19136.4]
  wire [14:0] _T_72500; // @[Modules.scala 166:64:@19138.4]
  wire [13:0] _T_72501; // @[Modules.scala 166:64:@19139.4]
  wire [13:0] buffer_5_592; // @[Modules.scala 166:64:@19140.4]
  wire [14:0] _T_72503; // @[Modules.scala 166:64:@19142.4]
  wire [13:0] _T_72504; // @[Modules.scala 166:64:@19143.4]
  wire [13:0] buffer_5_593; // @[Modules.scala 166:64:@19144.4]
  wire [14:0] _T_72506; // @[Modules.scala 166:64:@19146.4]
  wire [13:0] _T_72507; // @[Modules.scala 166:64:@19147.4]
  wire [13:0] buffer_5_594; // @[Modules.scala 166:64:@19148.4]
  wire [14:0] _T_72509; // @[Modules.scala 166:64:@19150.4]
  wire [13:0] _T_72510; // @[Modules.scala 166:64:@19151.4]
  wire [13:0] buffer_5_595; // @[Modules.scala 166:64:@19152.4]
  wire [14:0] _T_72512; // @[Modules.scala 166:64:@19154.4]
  wire [13:0] _T_72513; // @[Modules.scala 166:64:@19155.4]
  wire [13:0] buffer_5_596; // @[Modules.scala 166:64:@19156.4]
  wire [14:0] _T_72515; // @[Modules.scala 166:64:@19158.4]
  wire [13:0] _T_72516; // @[Modules.scala 166:64:@19159.4]
  wire [13:0] buffer_5_597; // @[Modules.scala 166:64:@19160.4]
  wire [14:0] _T_72518; // @[Modules.scala 166:64:@19162.4]
  wire [13:0] _T_72519; // @[Modules.scala 166:64:@19163.4]
  wire [13:0] buffer_5_598; // @[Modules.scala 166:64:@19164.4]
  wire [14:0] _T_72521; // @[Modules.scala 166:64:@19166.4]
  wire [13:0] _T_72522; // @[Modules.scala 166:64:@19167.4]
  wire [13:0] buffer_5_599; // @[Modules.scala 166:64:@19168.4]
  wire [14:0] _T_72524; // @[Modules.scala 166:64:@19170.4]
  wire [13:0] _T_72525; // @[Modules.scala 166:64:@19171.4]
  wire [13:0] buffer_5_600; // @[Modules.scala 166:64:@19172.4]
  wire [14:0] _T_72527; // @[Modules.scala 166:64:@19174.4]
  wire [13:0] _T_72528; // @[Modules.scala 166:64:@19175.4]
  wire [13:0] buffer_5_601; // @[Modules.scala 166:64:@19176.4]
  wire [14:0] _T_72530; // @[Modules.scala 166:64:@19178.4]
  wire [13:0] _T_72531; // @[Modules.scala 166:64:@19179.4]
  wire [13:0] buffer_5_602; // @[Modules.scala 166:64:@19180.4]
  wire [14:0] _T_72533; // @[Modules.scala 166:64:@19182.4]
  wire [13:0] _T_72534; // @[Modules.scala 166:64:@19183.4]
  wire [13:0] buffer_5_603; // @[Modules.scala 166:64:@19184.4]
  wire [14:0] _T_72536; // @[Modules.scala 166:64:@19186.4]
  wire [13:0] _T_72537; // @[Modules.scala 166:64:@19187.4]
  wire [13:0] buffer_5_604; // @[Modules.scala 166:64:@19188.4]
  wire [14:0] _T_72539; // @[Modules.scala 166:64:@19190.4]
  wire [13:0] _T_72540; // @[Modules.scala 166:64:@19191.4]
  wire [13:0] buffer_5_605; // @[Modules.scala 166:64:@19192.4]
  wire [14:0] _T_72542; // @[Modules.scala 166:64:@19194.4]
  wire [13:0] _T_72543; // @[Modules.scala 166:64:@19195.4]
  wire [13:0] buffer_5_606; // @[Modules.scala 166:64:@19196.4]
  wire [14:0] _T_72545; // @[Modules.scala 172:66:@19198.4]
  wire [13:0] _T_72546; // @[Modules.scala 172:66:@19199.4]
  wire [13:0] buffer_5_607; // @[Modules.scala 172:66:@19200.4]
  wire [14:0] _T_72548; // @[Modules.scala 160:64:@19202.4]
  wire [13:0] _T_72549; // @[Modules.scala 160:64:@19203.4]
  wire [13:0] buffer_5_608; // @[Modules.scala 160:64:@19204.4]
  wire [14:0] _T_72551; // @[Modules.scala 160:64:@19206.4]
  wire [13:0] _T_72552; // @[Modules.scala 160:64:@19207.4]
  wire [13:0] buffer_5_609; // @[Modules.scala 160:64:@19208.4]
  wire [14:0] _T_72554; // @[Modules.scala 160:64:@19210.4]
  wire [13:0] _T_72555; // @[Modules.scala 160:64:@19211.4]
  wire [13:0] buffer_5_610; // @[Modules.scala 160:64:@19212.4]
  wire [14:0] _T_72557; // @[Modules.scala 160:64:@19214.4]
  wire [13:0] _T_72558; // @[Modules.scala 160:64:@19215.4]
  wire [13:0] buffer_5_611; // @[Modules.scala 160:64:@19216.4]
  wire [14:0] _T_72560; // @[Modules.scala 160:64:@19218.4]
  wire [13:0] _T_72561; // @[Modules.scala 160:64:@19219.4]
  wire [13:0] buffer_5_612; // @[Modules.scala 160:64:@19220.4]
  wire [14:0] _T_72563; // @[Modules.scala 160:64:@19222.4]
  wire [13:0] _T_72564; // @[Modules.scala 160:64:@19223.4]
  wire [13:0] buffer_5_613; // @[Modules.scala 160:64:@19224.4]
  wire [14:0] _T_72566; // @[Modules.scala 160:64:@19226.4]
  wire [13:0] _T_72567; // @[Modules.scala 160:64:@19227.4]
  wire [13:0] buffer_5_614; // @[Modules.scala 160:64:@19228.4]
  wire [14:0] _T_72569; // @[Modules.scala 160:64:@19230.4]
  wire [13:0] _T_72570; // @[Modules.scala 160:64:@19231.4]
  wire [13:0] buffer_5_615; // @[Modules.scala 160:64:@19232.4]
  wire [14:0] _T_72572; // @[Modules.scala 160:64:@19234.4]
  wire [13:0] _T_72573; // @[Modules.scala 160:64:@19235.4]
  wire [13:0] buffer_5_616; // @[Modules.scala 160:64:@19236.4]
  wire [14:0] _T_72575; // @[Modules.scala 160:64:@19238.4]
  wire [13:0] _T_72576; // @[Modules.scala 160:64:@19239.4]
  wire [13:0] buffer_5_617; // @[Modules.scala 160:64:@19240.4]
  wire [14:0] _T_72578; // @[Modules.scala 160:64:@19242.4]
  wire [13:0] _T_72579; // @[Modules.scala 160:64:@19243.4]
  wire [13:0] buffer_5_618; // @[Modules.scala 160:64:@19244.4]
  wire [14:0] _T_72581; // @[Modules.scala 160:64:@19246.4]
  wire [13:0] _T_72582; // @[Modules.scala 160:64:@19247.4]
  wire [13:0] buffer_5_619; // @[Modules.scala 160:64:@19248.4]
  wire [14:0] _T_72584; // @[Modules.scala 160:64:@19250.4]
  wire [13:0] _T_72585; // @[Modules.scala 160:64:@19251.4]
  wire [13:0] buffer_5_620; // @[Modules.scala 160:64:@19252.4]
  wire [14:0] _T_72587; // @[Modules.scala 160:64:@19254.4]
  wire [13:0] _T_72588; // @[Modules.scala 160:64:@19255.4]
  wire [13:0] buffer_5_621; // @[Modules.scala 160:64:@19256.4]
  wire [14:0] _T_72590; // @[Modules.scala 160:64:@19258.4]
  wire [13:0] _T_72591; // @[Modules.scala 160:64:@19259.4]
  wire [13:0] buffer_5_622; // @[Modules.scala 160:64:@19260.4]
  wire [14:0] _T_72593; // @[Modules.scala 166:64:@19262.4]
  wire [13:0] _T_72594; // @[Modules.scala 166:64:@19263.4]
  wire [13:0] buffer_5_623; // @[Modules.scala 166:64:@19264.4]
  wire [14:0] _T_72596; // @[Modules.scala 166:64:@19266.4]
  wire [13:0] _T_72597; // @[Modules.scala 166:64:@19267.4]
  wire [13:0] buffer_5_624; // @[Modules.scala 166:64:@19268.4]
  wire [14:0] _T_72599; // @[Modules.scala 160:64:@19270.4]
  wire [13:0] _T_72600; // @[Modules.scala 160:64:@19271.4]
  wire [13:0] buffer_5_625; // @[Modules.scala 160:64:@19272.4]
  wire [14:0] _T_72602; // @[Modules.scala 172:66:@19274.4]
  wire [13:0] _T_72603; // @[Modules.scala 172:66:@19275.4]
  wire [13:0] buffer_5_626; // @[Modules.scala 172:66:@19276.4]
  wire [4:0] _T_72620; // @[Modules.scala 143:74:@19447.4]
  wire [5:0] _GEN_426; // @[Modules.scala 143:103:@19449.4]
  wire [6:0] _T_72623; // @[Modules.scala 143:103:@19449.4]
  wire [5:0] _T_72624; // @[Modules.scala 143:103:@19450.4]
  wire [5:0] _T_72625; // @[Modules.scala 143:103:@19451.4]
  wire [5:0] _T_72630; // @[Modules.scala 143:103:@19455.4]
  wire [4:0] _T_72631; // @[Modules.scala 143:103:@19456.4]
  wire [4:0] _T_72632; // @[Modules.scala 143:103:@19457.4]
  wire [5:0] _T_72637; // @[Modules.scala 143:103:@19461.4]
  wire [4:0] _T_72638; // @[Modules.scala 143:103:@19462.4]
  wire [4:0] _T_72639; // @[Modules.scala 143:103:@19463.4]
  wire [6:0] _T_72665; // @[Modules.scala 143:103:@19485.4]
  wire [5:0] _T_72666; // @[Modules.scala 143:103:@19486.4]
  wire [5:0] _T_72667; // @[Modules.scala 143:103:@19487.4]
  wire [6:0] _T_72672; // @[Modules.scala 143:103:@19491.4]
  wire [5:0] _T_72673; // @[Modules.scala 143:103:@19492.4]
  wire [5:0] _T_72674; // @[Modules.scala 143:103:@19493.4]
  wire [6:0] _T_72679; // @[Modules.scala 143:103:@19497.4]
  wire [5:0] _T_72680; // @[Modules.scala 143:103:@19498.4]
  wire [5:0] _T_72681; // @[Modules.scala 143:103:@19499.4]
  wire [6:0] _T_72686; // @[Modules.scala 143:103:@19503.4]
  wire [5:0] _T_72687; // @[Modules.scala 143:103:@19504.4]
  wire [5:0] _T_72688; // @[Modules.scala 143:103:@19505.4]
  wire [5:0] _T_72749; // @[Modules.scala 143:103:@19557.4]
  wire [4:0] _T_72750; // @[Modules.scala 143:103:@19558.4]
  wire [4:0] _T_72751; // @[Modules.scala 143:103:@19559.4]
  wire [5:0] _T_72756; // @[Modules.scala 143:103:@19563.4]
  wire [4:0] _T_72757; // @[Modules.scala 143:103:@19564.4]
  wire [4:0] _T_72758; // @[Modules.scala 143:103:@19565.4]
  wire [5:0] _GEN_431; // @[Modules.scala 143:103:@19569.4]
  wire [6:0] _T_72763; // @[Modules.scala 143:103:@19569.4]
  wire [5:0] _T_72764; // @[Modules.scala 143:103:@19570.4]
  wire [5:0] _T_72765; // @[Modules.scala 143:103:@19571.4]
  wire [6:0] _T_72784; // @[Modules.scala 143:103:@19587.4]
  wire [5:0] _T_72785; // @[Modules.scala 143:103:@19588.4]
  wire [5:0] _T_72786; // @[Modules.scala 143:103:@19589.4]
  wire [6:0] _T_72791; // @[Modules.scala 143:103:@19593.4]
  wire [5:0] _T_72792; // @[Modules.scala 143:103:@19594.4]
  wire [5:0] _T_72793; // @[Modules.scala 143:103:@19595.4]
  wire [5:0] _GEN_433; // @[Modules.scala 143:103:@19611.4]
  wire [6:0] _T_72812; // @[Modules.scala 143:103:@19611.4]
  wire [5:0] _T_72813; // @[Modules.scala 143:103:@19612.4]
  wire [5:0] _T_72814; // @[Modules.scala 143:103:@19613.4]
  wire [5:0] _GEN_434; // @[Modules.scala 143:103:@19617.4]
  wire [6:0] _T_72819; // @[Modules.scala 143:103:@19617.4]
  wire [5:0] _T_72820; // @[Modules.scala 143:103:@19618.4]
  wire [5:0] _T_72821; // @[Modules.scala 143:103:@19619.4]
  wire [5:0] _GEN_436; // @[Modules.scala 143:103:@19635.4]
  wire [6:0] _T_72840; // @[Modules.scala 143:103:@19635.4]
  wire [5:0] _T_72841; // @[Modules.scala 143:103:@19636.4]
  wire [5:0] _T_72842; // @[Modules.scala 143:103:@19637.4]
  wire [6:0] _T_72854; // @[Modules.scala 143:103:@19647.4]
  wire [5:0] _T_72855; // @[Modules.scala 143:103:@19648.4]
  wire [5:0] _T_72856; // @[Modules.scala 143:103:@19649.4]
  wire [6:0] _T_72882; // @[Modules.scala 143:103:@19671.4]
  wire [5:0] _T_72883; // @[Modules.scala 143:103:@19672.4]
  wire [5:0] _T_72884; // @[Modules.scala 143:103:@19673.4]
  wire [6:0] _T_72917; // @[Modules.scala 143:103:@19701.4]
  wire [5:0] _T_72918; // @[Modules.scala 143:103:@19702.4]
  wire [5:0] _T_72919; // @[Modules.scala 143:103:@19703.4]
  wire [6:0] _T_72924; // @[Modules.scala 143:103:@19707.4]
  wire [5:0] _T_72925; // @[Modules.scala 143:103:@19708.4]
  wire [5:0] _T_72926; // @[Modules.scala 143:103:@19709.4]
  wire [6:0] _T_72931; // @[Modules.scala 143:103:@19713.4]
  wire [5:0] _T_72932; // @[Modules.scala 143:103:@19714.4]
  wire [5:0] _T_72933; // @[Modules.scala 143:103:@19715.4]
  wire [6:0] _T_72959; // @[Modules.scala 143:103:@19737.4]
  wire [5:0] _T_72960; // @[Modules.scala 143:103:@19738.4]
  wire [5:0] _T_72961; // @[Modules.scala 143:103:@19739.4]
  wire [6:0] _T_72966; // @[Modules.scala 143:103:@19743.4]
  wire [5:0] _T_72967; // @[Modules.scala 143:103:@19744.4]
  wire [5:0] _T_72968; // @[Modules.scala 143:103:@19745.4]
  wire [6:0] _T_73001; // @[Modules.scala 143:103:@19773.4]
  wire [5:0] _T_73002; // @[Modules.scala 143:103:@19774.4]
  wire [5:0] _T_73003; // @[Modules.scala 143:103:@19775.4]
  wire [6:0] _T_73008; // @[Modules.scala 143:103:@19779.4]
  wire [5:0] _T_73009; // @[Modules.scala 143:103:@19780.4]
  wire [5:0] _T_73010; // @[Modules.scala 143:103:@19781.4]
  wire [6:0] _T_73015; // @[Modules.scala 143:103:@19785.4]
  wire [5:0] _T_73016; // @[Modules.scala 143:103:@19786.4]
  wire [5:0] _T_73017; // @[Modules.scala 143:103:@19787.4]
  wire [5:0] _T_73021; // @[Modules.scala 144:80:@19790.4]
  wire [6:0] _T_73022; // @[Modules.scala 143:103:@19791.4]
  wire [5:0] _T_73023; // @[Modules.scala 143:103:@19792.4]
  wire [5:0] _T_73024; // @[Modules.scala 143:103:@19793.4]
  wire [6:0] _T_73029; // @[Modules.scala 143:103:@19797.4]
  wire [5:0] _T_73030; // @[Modules.scala 143:103:@19798.4]
  wire [5:0] _T_73031; // @[Modules.scala 143:103:@19799.4]
  wire [6:0] _T_73036; // @[Modules.scala 143:103:@19803.4]
  wire [5:0] _T_73037; // @[Modules.scala 143:103:@19804.4]
  wire [5:0] _T_73038; // @[Modules.scala 143:103:@19805.4]
  wire [5:0] _GEN_443; // @[Modules.scala 143:103:@19809.4]
  wire [6:0] _T_73043; // @[Modules.scala 143:103:@19809.4]
  wire [5:0] _T_73044; // @[Modules.scala 143:103:@19810.4]
  wire [5:0] _T_73045; // @[Modules.scala 143:103:@19811.4]
  wire [5:0] _T_73049; // @[Modules.scala 144:80:@19814.4]
  wire [6:0] _T_73050; // @[Modules.scala 143:103:@19815.4]
  wire [5:0] _T_73051; // @[Modules.scala 143:103:@19816.4]
  wire [5:0] _T_73052; // @[Modules.scala 143:103:@19817.4]
  wire [6:0] _T_73071; // @[Modules.scala 143:103:@19833.4]
  wire [5:0] _T_73072; // @[Modules.scala 143:103:@19834.4]
  wire [5:0] _T_73073; // @[Modules.scala 143:103:@19835.4]
  wire [6:0] _T_73078; // @[Modules.scala 143:103:@19839.4]
  wire [5:0] _T_73079; // @[Modules.scala 143:103:@19840.4]
  wire [5:0] _T_73080; // @[Modules.scala 143:103:@19841.4]
  wire [6:0] _T_73092; // @[Modules.scala 143:103:@19851.4]
  wire [5:0] _T_73093; // @[Modules.scala 143:103:@19852.4]
  wire [5:0] _T_73094; // @[Modules.scala 143:103:@19853.4]
  wire [6:0] _T_73099; // @[Modules.scala 143:103:@19857.4]
  wire [5:0] _T_73100; // @[Modules.scala 143:103:@19858.4]
  wire [5:0] _T_73101; // @[Modules.scala 143:103:@19859.4]
  wire [6:0] _T_73106; // @[Modules.scala 143:103:@19863.4]
  wire [5:0] _T_73107; // @[Modules.scala 143:103:@19864.4]
  wire [5:0] _T_73108; // @[Modules.scala 143:103:@19865.4]
  wire [5:0] _T_73120; // @[Modules.scala 143:103:@19875.4]
  wire [4:0] _T_73121; // @[Modules.scala 143:103:@19876.4]
  wire [4:0] _T_73122; // @[Modules.scala 143:103:@19877.4]
  wire [6:0] _T_73127; // @[Modules.scala 143:103:@19881.4]
  wire [5:0] _T_73128; // @[Modules.scala 143:103:@19882.4]
  wire [5:0] _T_73129; // @[Modules.scala 143:103:@19883.4]
  wire [5:0] _GEN_446; // @[Modules.scala 143:103:@19887.4]
  wire [6:0] _T_73134; // @[Modules.scala 143:103:@19887.4]
  wire [5:0] _T_73135; // @[Modules.scala 143:103:@19888.4]
  wire [5:0] _T_73136; // @[Modules.scala 143:103:@19889.4]
  wire [5:0] _T_73141; // @[Modules.scala 143:103:@19893.4]
  wire [4:0] _T_73142; // @[Modules.scala 143:103:@19894.4]
  wire [4:0] _T_73143; // @[Modules.scala 143:103:@19895.4]
  wire [5:0] _T_73148; // @[Modules.scala 143:103:@19899.4]
  wire [4:0] _T_73149; // @[Modules.scala 143:103:@19900.4]
  wire [4:0] _T_73150; // @[Modules.scala 143:103:@19901.4]
  wire [6:0] _T_73155; // @[Modules.scala 143:103:@19905.4]
  wire [5:0] _T_73156; // @[Modules.scala 143:103:@19906.4]
  wire [5:0] _T_73157; // @[Modules.scala 143:103:@19907.4]
  wire [6:0] _T_73176; // @[Modules.scala 143:103:@19923.4]
  wire [5:0] _T_73177; // @[Modules.scala 143:103:@19924.4]
  wire [5:0] _T_73178; // @[Modules.scala 143:103:@19925.4]
  wire [6:0] _T_73183; // @[Modules.scala 143:103:@19929.4]
  wire [5:0] _T_73184; // @[Modules.scala 143:103:@19930.4]
  wire [5:0] _T_73185; // @[Modules.scala 143:103:@19931.4]
  wire [5:0] _GEN_450; // @[Modules.scala 143:103:@19965.4]
  wire [6:0] _T_73225; // @[Modules.scala 143:103:@19965.4]
  wire [5:0] _T_73226; // @[Modules.scala 143:103:@19966.4]
  wire [5:0] _T_73227; // @[Modules.scala 143:103:@19967.4]
  wire [5:0] _GEN_451; // @[Modules.scala 143:103:@19977.4]
  wire [6:0] _T_73239; // @[Modules.scala 143:103:@19977.4]
  wire [5:0] _T_73240; // @[Modules.scala 143:103:@19978.4]
  wire [5:0] _T_73241; // @[Modules.scala 143:103:@19979.4]
  wire [5:0] _GEN_452; // @[Modules.scala 143:103:@20001.4]
  wire [6:0] _T_73267; // @[Modules.scala 143:103:@20001.4]
  wire [5:0] _T_73268; // @[Modules.scala 143:103:@20002.4]
  wire [5:0] _T_73269; // @[Modules.scala 143:103:@20003.4]
  wire [5:0] _T_73274; // @[Modules.scala 143:103:@20007.4]
  wire [4:0] _T_73275; // @[Modules.scala 143:103:@20008.4]
  wire [4:0] _T_73276; // @[Modules.scala 143:103:@20009.4]
  wire [5:0] _T_73281; // @[Modules.scala 143:103:@20013.4]
  wire [4:0] _T_73282; // @[Modules.scala 143:103:@20014.4]
  wire [4:0] _T_73283; // @[Modules.scala 143:103:@20015.4]
  wire [5:0] _GEN_453; // @[Modules.scala 143:103:@20019.4]
  wire [6:0] _T_73288; // @[Modules.scala 143:103:@20019.4]
  wire [5:0] _T_73289; // @[Modules.scala 143:103:@20020.4]
  wire [5:0] _T_73290; // @[Modules.scala 143:103:@20021.4]
  wire [5:0] _GEN_454; // @[Modules.scala 143:103:@20037.4]
  wire [6:0] _T_73309; // @[Modules.scala 143:103:@20037.4]
  wire [5:0] _T_73310; // @[Modules.scala 143:103:@20038.4]
  wire [5:0] _T_73311; // @[Modules.scala 143:103:@20039.4]
  wire [5:0] _T_73316; // @[Modules.scala 143:103:@20043.4]
  wire [4:0] _T_73317; // @[Modules.scala 143:103:@20044.4]
  wire [4:0] _T_73318; // @[Modules.scala 143:103:@20045.4]
  wire [5:0] _GEN_455; // @[Modules.scala 143:103:@20049.4]
  wire [6:0] _T_73323; // @[Modules.scala 143:103:@20049.4]
  wire [5:0] _T_73324; // @[Modules.scala 143:103:@20050.4]
  wire [5:0] _T_73325; // @[Modules.scala 143:103:@20051.4]
  wire [6:0] _T_73344; // @[Modules.scala 143:103:@20067.4]
  wire [5:0] _T_73345; // @[Modules.scala 143:103:@20068.4]
  wire [5:0] _T_73346; // @[Modules.scala 143:103:@20069.4]
  wire [6:0] _T_73386; // @[Modules.scala 143:103:@20103.4]
  wire [5:0] _T_73387; // @[Modules.scala 143:103:@20104.4]
  wire [5:0] _T_73388; // @[Modules.scala 143:103:@20105.4]
  wire [5:0] _GEN_457; // @[Modules.scala 143:103:@20109.4]
  wire [6:0] _T_73393; // @[Modules.scala 143:103:@20109.4]
  wire [5:0] _T_73394; // @[Modules.scala 143:103:@20110.4]
  wire [5:0] _T_73395; // @[Modules.scala 143:103:@20111.4]
  wire [5:0] _GEN_458; // @[Modules.scala 143:103:@20121.4]
  wire [6:0] _T_73407; // @[Modules.scala 143:103:@20121.4]
  wire [5:0] _T_73408; // @[Modules.scala 143:103:@20122.4]
  wire [5:0] _T_73409; // @[Modules.scala 143:103:@20123.4]
  wire [5:0] _GEN_459; // @[Modules.scala 143:103:@20145.4]
  wire [6:0] _T_73435; // @[Modules.scala 143:103:@20145.4]
  wire [5:0] _T_73436; // @[Modules.scala 143:103:@20146.4]
  wire [5:0] _T_73437; // @[Modules.scala 143:103:@20147.4]
  wire [6:0] _T_73463; // @[Modules.scala 143:103:@20169.4]
  wire [5:0] _T_73464; // @[Modules.scala 143:103:@20170.4]
  wire [5:0] _T_73465; // @[Modules.scala 143:103:@20171.4]
  wire [6:0] _T_73505; // @[Modules.scala 143:103:@20205.4]
  wire [5:0] _T_73506; // @[Modules.scala 143:103:@20206.4]
  wire [5:0] _T_73507; // @[Modules.scala 143:103:@20207.4]
  wire [5:0] _GEN_461; // @[Modules.scala 143:103:@20217.4]
  wire [6:0] _T_73519; // @[Modules.scala 143:103:@20217.4]
  wire [5:0] _T_73520; // @[Modules.scala 143:103:@20218.4]
  wire [5:0] _T_73521; // @[Modules.scala 143:103:@20219.4]
  wire [6:0] _T_73554; // @[Modules.scala 143:103:@20247.4]
  wire [5:0] _T_73555; // @[Modules.scala 143:103:@20248.4]
  wire [5:0] _T_73556; // @[Modules.scala 143:103:@20249.4]
  wire [6:0] _T_73561; // @[Modules.scala 143:103:@20253.4]
  wire [5:0] _T_73562; // @[Modules.scala 143:103:@20254.4]
  wire [5:0] _T_73563; // @[Modules.scala 143:103:@20255.4]
  wire [4:0] _T_73565; // @[Modules.scala 143:74:@20257.4]
  wire [5:0] _GEN_463; // @[Modules.scala 143:103:@20259.4]
  wire [6:0] _T_73568; // @[Modules.scala 143:103:@20259.4]
  wire [5:0] _T_73569; // @[Modules.scala 143:103:@20260.4]
  wire [5:0] _T_73570; // @[Modules.scala 143:103:@20261.4]
  wire [6:0] _T_73589; // @[Modules.scala 143:103:@20277.4]
  wire [5:0] _T_73590; // @[Modules.scala 143:103:@20278.4]
  wire [5:0] _T_73591; // @[Modules.scala 143:103:@20279.4]
  wire [6:0] _T_73596; // @[Modules.scala 143:103:@20283.4]
  wire [5:0] _T_73597; // @[Modules.scala 143:103:@20284.4]
  wire [5:0] _T_73598; // @[Modules.scala 143:103:@20285.4]
  wire [5:0] _GEN_466; // @[Modules.scala 143:103:@20301.4]
  wire [6:0] _T_73617; // @[Modules.scala 143:103:@20301.4]
  wire [5:0] _T_73618; // @[Modules.scala 143:103:@20302.4]
  wire [5:0] _T_73619; // @[Modules.scala 143:103:@20303.4]
  wire [5:0] _T_73652; // @[Modules.scala 143:103:@20331.4]
  wire [4:0] _T_73653; // @[Modules.scala 143:103:@20332.4]
  wire [4:0] _T_73654; // @[Modules.scala 143:103:@20333.4]
  wire [4:0] _T_73663; // @[Modules.scala 143:74:@20341.4]
  wire [5:0] _T_73666; // @[Modules.scala 143:103:@20343.4]
  wire [4:0] _T_73667; // @[Modules.scala 143:103:@20344.4]
  wire [4:0] _T_73668; // @[Modules.scala 143:103:@20345.4]
  wire [5:0] _T_73764; // @[Modules.scala 143:103:@20427.4]
  wire [4:0] _T_73765; // @[Modules.scala 143:103:@20428.4]
  wire [4:0] _T_73766; // @[Modules.scala 143:103:@20429.4]
  wire [5:0] _GEN_469; // @[Modules.scala 143:103:@20451.4]
  wire [6:0] _T_73792; // @[Modules.scala 143:103:@20451.4]
  wire [5:0] _T_73793; // @[Modules.scala 143:103:@20452.4]
  wire [5:0] _T_73794; // @[Modules.scala 143:103:@20453.4]
  wire [6:0] _T_73806; // @[Modules.scala 143:103:@20463.4]
  wire [5:0] _T_73807; // @[Modules.scala 143:103:@20464.4]
  wire [5:0] _T_73808; // @[Modules.scala 143:103:@20465.4]
  wire [6:0] _T_73834; // @[Modules.scala 143:103:@20487.4]
  wire [5:0] _T_73835; // @[Modules.scala 143:103:@20488.4]
  wire [5:0] _T_73836; // @[Modules.scala 143:103:@20489.4]
  wire [5:0] _T_73848; // @[Modules.scala 143:103:@20499.4]
  wire [4:0] _T_73849; // @[Modules.scala 143:103:@20500.4]
  wire [4:0] _T_73850; // @[Modules.scala 143:103:@20501.4]
  wire [5:0] _GEN_471; // @[Modules.scala 143:103:@20505.4]
  wire [6:0] _T_73855; // @[Modules.scala 143:103:@20505.4]
  wire [5:0] _T_73856; // @[Modules.scala 143:103:@20506.4]
  wire [5:0] _T_73857; // @[Modules.scala 143:103:@20507.4]
  wire [6:0] _T_73869; // @[Modules.scala 143:103:@20517.4]
  wire [5:0] _T_73870; // @[Modules.scala 143:103:@20518.4]
  wire [5:0] _T_73871; // @[Modules.scala 143:103:@20519.4]
  wire [6:0] _T_73890; // @[Modules.scala 143:103:@20535.4]
  wire [5:0] _T_73891; // @[Modules.scala 143:103:@20536.4]
  wire [5:0] _T_73892; // @[Modules.scala 143:103:@20537.4]
  wire [6:0] _T_73904; // @[Modules.scala 143:103:@20547.4]
  wire [5:0] _T_73905; // @[Modules.scala 143:103:@20548.4]
  wire [5:0] _T_73906; // @[Modules.scala 143:103:@20549.4]
  wire [6:0] _T_73925; // @[Modules.scala 143:103:@20565.4]
  wire [5:0] _T_73926; // @[Modules.scala 143:103:@20566.4]
  wire [5:0] _T_73927; // @[Modules.scala 143:103:@20567.4]
  wire [6:0] _T_73932; // @[Modules.scala 143:103:@20571.4]
  wire [5:0] _T_73933; // @[Modules.scala 143:103:@20572.4]
  wire [5:0] _T_73934; // @[Modules.scala 143:103:@20573.4]
  wire [5:0] _T_73936; // @[Modules.scala 143:74:@20575.4]
  wire [6:0] _T_73939; // @[Modules.scala 143:103:@20577.4]
  wire [5:0] _T_73940; // @[Modules.scala 143:103:@20578.4]
  wire [5:0] _T_73941; // @[Modules.scala 143:103:@20579.4]
  wire [6:0] _T_73953; // @[Modules.scala 143:103:@20589.4]
  wire [5:0] _T_73954; // @[Modules.scala 143:103:@20590.4]
  wire [5:0] _T_73955; // @[Modules.scala 143:103:@20591.4]
  wire [6:0] _T_73960; // @[Modules.scala 143:103:@20595.4]
  wire [5:0] _T_73961; // @[Modules.scala 143:103:@20596.4]
  wire [5:0] _T_73962; // @[Modules.scala 143:103:@20597.4]
  wire [6:0] _T_73967; // @[Modules.scala 143:103:@20601.4]
  wire [5:0] _T_73968; // @[Modules.scala 143:103:@20602.4]
  wire [5:0] _T_73969; // @[Modules.scala 143:103:@20603.4]
  wire [6:0] _T_73974; // @[Modules.scala 143:103:@20607.4]
  wire [5:0] _T_73975; // @[Modules.scala 143:103:@20608.4]
  wire [5:0] _T_73976; // @[Modules.scala 143:103:@20609.4]
  wire [5:0] _GEN_473; // @[Modules.scala 143:103:@20625.4]
  wire [6:0] _T_73995; // @[Modules.scala 143:103:@20625.4]
  wire [5:0] _T_73996; // @[Modules.scala 143:103:@20626.4]
  wire [5:0] _T_73997; // @[Modules.scala 143:103:@20627.4]
  wire [6:0] _T_74009; // @[Modules.scala 143:103:@20637.4]
  wire [5:0] _T_74010; // @[Modules.scala 143:103:@20638.4]
  wire [5:0] _T_74011; // @[Modules.scala 143:103:@20639.4]
  wire [6:0] _T_74023; // @[Modules.scala 143:103:@20649.4]
  wire [5:0] _T_74024; // @[Modules.scala 143:103:@20650.4]
  wire [5:0] _T_74025; // @[Modules.scala 143:103:@20651.4]
  wire [5:0] _GEN_475; // @[Modules.scala 143:103:@20703.4]
  wire [6:0] _T_74086; // @[Modules.scala 143:103:@20703.4]
  wire [5:0] _T_74087; // @[Modules.scala 143:103:@20704.4]
  wire [5:0] _T_74088; // @[Modules.scala 143:103:@20705.4]
  wire [6:0] _T_74093; // @[Modules.scala 143:103:@20709.4]
  wire [5:0] _T_74094; // @[Modules.scala 143:103:@20710.4]
  wire [5:0] _T_74095; // @[Modules.scala 143:103:@20711.4]
  wire [6:0] _T_74100; // @[Modules.scala 143:103:@20715.4]
  wire [5:0] _T_74101; // @[Modules.scala 143:103:@20716.4]
  wire [5:0] _T_74102; // @[Modules.scala 143:103:@20717.4]
  wire [5:0] _GEN_478; // @[Modules.scala 143:103:@20757.4]
  wire [6:0] _T_74149; // @[Modules.scala 143:103:@20757.4]
  wire [5:0] _T_74150; // @[Modules.scala 143:103:@20758.4]
  wire [5:0] _T_74151; // @[Modules.scala 143:103:@20759.4]
  wire [6:0] _T_74170; // @[Modules.scala 143:103:@20775.4]
  wire [5:0] _T_74171; // @[Modules.scala 143:103:@20776.4]
  wire [5:0] _T_74172; // @[Modules.scala 143:103:@20777.4]
  wire [6:0] _T_74177; // @[Modules.scala 143:103:@20781.4]
  wire [5:0] _T_74178; // @[Modules.scala 143:103:@20782.4]
  wire [5:0] _T_74179; // @[Modules.scala 143:103:@20783.4]
  wire [6:0] _T_74184; // @[Modules.scala 143:103:@20787.4]
  wire [5:0] _T_74185; // @[Modules.scala 143:103:@20788.4]
  wire [5:0] _T_74186; // @[Modules.scala 143:103:@20789.4]
  wire [5:0] _T_74191; // @[Modules.scala 143:103:@20793.4]
  wire [4:0] _T_74192; // @[Modules.scala 143:103:@20794.4]
  wire [4:0] _T_74193; // @[Modules.scala 143:103:@20795.4]
  wire [5:0] _GEN_479; // @[Modules.scala 143:103:@20799.4]
  wire [6:0] _T_74198; // @[Modules.scala 143:103:@20799.4]
  wire [5:0] _T_74199; // @[Modules.scala 143:103:@20800.4]
  wire [5:0] _T_74200; // @[Modules.scala 143:103:@20801.4]
  wire [6:0] _T_74205; // @[Modules.scala 143:103:@20805.4]
  wire [5:0] _T_74206; // @[Modules.scala 143:103:@20806.4]
  wire [5:0] _T_74207; // @[Modules.scala 143:103:@20807.4]
  wire [6:0] _T_74212; // @[Modules.scala 143:103:@20811.4]
  wire [5:0] _T_74213; // @[Modules.scala 143:103:@20812.4]
  wire [5:0] _T_74214; // @[Modules.scala 143:103:@20813.4]
  wire [5:0] _GEN_481; // @[Modules.scala 143:103:@20817.4]
  wire [6:0] _T_74219; // @[Modules.scala 143:103:@20817.4]
  wire [5:0] _T_74220; // @[Modules.scala 143:103:@20818.4]
  wire [5:0] _T_74221; // @[Modules.scala 143:103:@20819.4]
  wire [5:0] _GEN_482; // @[Modules.scala 143:103:@20835.4]
  wire [6:0] _T_74240; // @[Modules.scala 143:103:@20835.4]
  wire [5:0] _T_74241; // @[Modules.scala 143:103:@20836.4]
  wire [5:0] _T_74242; // @[Modules.scala 143:103:@20837.4]
  wire [5:0] _T_74260; // @[Modules.scala 144:80:@20852.4]
  wire [6:0] _T_74261; // @[Modules.scala 143:103:@20853.4]
  wire [5:0] _T_74262; // @[Modules.scala 143:103:@20854.4]
  wire [5:0] _T_74263; // @[Modules.scala 143:103:@20855.4]
  wire [6:0] _T_74289; // @[Modules.scala 143:103:@20877.4]
  wire [5:0] _T_74290; // @[Modules.scala 143:103:@20878.4]
  wire [5:0] _T_74291; // @[Modules.scala 143:103:@20879.4]
  wire [6:0] _T_74296; // @[Modules.scala 143:103:@20883.4]
  wire [5:0] _T_74297; // @[Modules.scala 143:103:@20884.4]
  wire [5:0] _T_74298; // @[Modules.scala 143:103:@20885.4]
  wire [6:0] _T_74310; // @[Modules.scala 143:103:@20895.4]
  wire [5:0] _T_74311; // @[Modules.scala 143:103:@20896.4]
  wire [5:0] _T_74312; // @[Modules.scala 143:103:@20897.4]
  wire [5:0] _T_74317; // @[Modules.scala 143:103:@20901.4]
  wire [4:0] _T_74318; // @[Modules.scala 143:103:@20902.4]
  wire [4:0] _T_74319; // @[Modules.scala 143:103:@20903.4]
  wire [5:0] _T_74323; // @[Modules.scala 144:80:@20906.4]
  wire [5:0] _GEN_485; // @[Modules.scala 143:103:@20907.4]
  wire [6:0] _T_74324; // @[Modules.scala 143:103:@20907.4]
  wire [5:0] _T_74325; // @[Modules.scala 143:103:@20908.4]
  wire [5:0] _T_74326; // @[Modules.scala 143:103:@20909.4]
  wire [5:0] _T_74330; // @[Modules.scala 144:80:@20912.4]
  wire [6:0] _T_74331; // @[Modules.scala 143:103:@20913.4]
  wire [5:0] _T_74332; // @[Modules.scala 143:103:@20914.4]
  wire [5:0] _T_74333; // @[Modules.scala 143:103:@20915.4]
  wire [6:0] _T_74338; // @[Modules.scala 143:103:@20919.4]
  wire [5:0] _T_74339; // @[Modules.scala 143:103:@20920.4]
  wire [5:0] _T_74340; // @[Modules.scala 143:103:@20921.4]
  wire [5:0] _GEN_486; // @[Modules.scala 143:103:@20925.4]
  wire [6:0] _T_74345; // @[Modules.scala 143:103:@20925.4]
  wire [5:0] _T_74346; // @[Modules.scala 143:103:@20926.4]
  wire [5:0] _T_74347; // @[Modules.scala 143:103:@20927.4]
  wire [6:0] _T_74352; // @[Modules.scala 143:103:@20931.4]
  wire [5:0] _T_74353; // @[Modules.scala 143:103:@20932.4]
  wire [5:0] _T_74354; // @[Modules.scala 143:103:@20933.4]
  wire [5:0] _T_74359; // @[Modules.scala 143:103:@20937.4]
  wire [4:0] _T_74360; // @[Modules.scala 143:103:@20938.4]
  wire [4:0] _T_74361; // @[Modules.scala 143:103:@20939.4]
  wire [6:0] _T_74366; // @[Modules.scala 143:103:@20943.4]
  wire [5:0] _T_74367; // @[Modules.scala 143:103:@20944.4]
  wire [5:0] _T_74368; // @[Modules.scala 143:103:@20945.4]
  wire [6:0] _T_74373; // @[Modules.scala 143:103:@20949.4]
  wire [5:0] _T_74374; // @[Modules.scala 143:103:@20950.4]
  wire [5:0] _T_74375; // @[Modules.scala 143:103:@20951.4]
  wire [6:0] _T_74380; // @[Modules.scala 143:103:@20955.4]
  wire [5:0] _T_74381; // @[Modules.scala 143:103:@20956.4]
  wire [5:0] _T_74382; // @[Modules.scala 143:103:@20957.4]
  wire [6:0] _T_74408; // @[Modules.scala 143:103:@20979.4]
  wire [5:0] _T_74409; // @[Modules.scala 143:103:@20980.4]
  wire [5:0] _T_74410; // @[Modules.scala 143:103:@20981.4]
  wire [6:0] _T_74415; // @[Modules.scala 143:103:@20985.4]
  wire [5:0] _T_74416; // @[Modules.scala 143:103:@20986.4]
  wire [5:0] _T_74417; // @[Modules.scala 143:103:@20987.4]
  wire [6:0] _T_74422; // @[Modules.scala 143:103:@20991.4]
  wire [5:0] _T_74423; // @[Modules.scala 143:103:@20992.4]
  wire [5:0] _T_74424; // @[Modules.scala 143:103:@20993.4]
  wire [6:0] _T_74429; // @[Modules.scala 143:103:@20997.4]
  wire [5:0] _T_74430; // @[Modules.scala 143:103:@20998.4]
  wire [5:0] _T_74431; // @[Modules.scala 143:103:@20999.4]
  wire [6:0] _T_74450; // @[Modules.scala 143:103:@21015.4]
  wire [5:0] _T_74451; // @[Modules.scala 143:103:@21016.4]
  wire [5:0] _T_74452; // @[Modules.scala 143:103:@21017.4]
  wire [5:0] _GEN_490; // @[Modules.scala 143:103:@21021.4]
  wire [6:0] _T_74457; // @[Modules.scala 143:103:@21021.4]
  wire [5:0] _T_74458; // @[Modules.scala 143:103:@21022.4]
  wire [5:0] _T_74459; // @[Modules.scala 143:103:@21023.4]
  wire [5:0] _T_74464; // @[Modules.scala 143:103:@21027.4]
  wire [4:0] _T_74465; // @[Modules.scala 143:103:@21028.4]
  wire [4:0] _T_74466; // @[Modules.scala 143:103:@21029.4]
  wire [5:0] _T_74485; // @[Modules.scala 143:103:@21045.4]
  wire [4:0] _T_74486; // @[Modules.scala 143:103:@21046.4]
  wire [4:0] _T_74487; // @[Modules.scala 143:103:@21047.4]
  wire [5:0] _T_74492; // @[Modules.scala 143:103:@21051.4]
  wire [4:0] _T_74493; // @[Modules.scala 143:103:@21052.4]
  wire [4:0] _T_74494; // @[Modules.scala 143:103:@21053.4]
  wire [6:0] _T_74499; // @[Modules.scala 143:103:@21057.4]
  wire [5:0] _T_74500; // @[Modules.scala 143:103:@21058.4]
  wire [5:0] _T_74501; // @[Modules.scala 143:103:@21059.4]
  wire [6:0] _T_74506; // @[Modules.scala 143:103:@21063.4]
  wire [5:0] _T_74507; // @[Modules.scala 143:103:@21064.4]
  wire [5:0] _T_74508; // @[Modules.scala 143:103:@21065.4]
  wire [6:0] _T_74513; // @[Modules.scala 143:103:@21069.4]
  wire [5:0] _T_74514; // @[Modules.scala 143:103:@21070.4]
  wire [5:0] _T_74515; // @[Modules.scala 143:103:@21071.4]
  wire [6:0] _T_74520; // @[Modules.scala 143:103:@21075.4]
  wire [5:0] _T_74521; // @[Modules.scala 143:103:@21076.4]
  wire [5:0] _T_74522; // @[Modules.scala 143:103:@21077.4]
  wire [6:0] _T_74527; // @[Modules.scala 143:103:@21081.4]
  wire [5:0] _T_74528; // @[Modules.scala 143:103:@21082.4]
  wire [5:0] _T_74529; // @[Modules.scala 143:103:@21083.4]
  wire [5:0] _T_74555; // @[Modules.scala 143:103:@21105.4]
  wire [4:0] _T_74556; // @[Modules.scala 143:103:@21106.4]
  wire [4:0] _T_74557; // @[Modules.scala 143:103:@21107.4]
  wire [5:0] _T_74562; // @[Modules.scala 143:103:@21111.4]
  wire [4:0] _T_74563; // @[Modules.scala 143:103:@21112.4]
  wire [4:0] _T_74564; // @[Modules.scala 143:103:@21113.4]
  wire [5:0] _T_74569; // @[Modules.scala 143:103:@21117.4]
  wire [4:0] _T_74570; // @[Modules.scala 143:103:@21118.4]
  wire [4:0] _T_74571; // @[Modules.scala 143:103:@21119.4]
  wire [6:0] _T_74583; // @[Modules.scala 143:103:@21129.4]
  wire [5:0] _T_74584; // @[Modules.scala 143:103:@21130.4]
  wire [5:0] _T_74585; // @[Modules.scala 143:103:@21131.4]
  wire [6:0] _T_74590; // @[Modules.scala 143:103:@21135.4]
  wire [5:0] _T_74591; // @[Modules.scala 143:103:@21136.4]
  wire [5:0] _T_74592; // @[Modules.scala 143:103:@21137.4]
  wire [6:0] _T_74597; // @[Modules.scala 143:103:@21141.4]
  wire [5:0] _T_74598; // @[Modules.scala 143:103:@21142.4]
  wire [5:0] _T_74599; // @[Modules.scala 143:103:@21143.4]
  wire [6:0] _T_74604; // @[Modules.scala 143:103:@21147.4]
  wire [5:0] _T_74605; // @[Modules.scala 143:103:@21148.4]
  wire [5:0] _T_74606; // @[Modules.scala 143:103:@21149.4]
  wire [6:0] _T_74611; // @[Modules.scala 143:103:@21153.4]
  wire [5:0] _T_74612; // @[Modules.scala 143:103:@21154.4]
  wire [5:0] _T_74613; // @[Modules.scala 143:103:@21155.4]
  wire [6:0] _T_74632; // @[Modules.scala 143:103:@21171.4]
  wire [5:0] _T_74633; // @[Modules.scala 143:103:@21172.4]
  wire [5:0] _T_74634; // @[Modules.scala 143:103:@21173.4]
  wire [5:0] _T_74646; // @[Modules.scala 143:103:@21183.4]
  wire [4:0] _T_74647; // @[Modules.scala 143:103:@21184.4]
  wire [4:0] _T_74648; // @[Modules.scala 143:103:@21185.4]
  wire [5:0] _T_74653; // @[Modules.scala 143:103:@21189.4]
  wire [4:0] _T_74654; // @[Modules.scala 143:103:@21190.4]
  wire [4:0] _T_74655; // @[Modules.scala 143:103:@21191.4]
  wire [5:0] _T_74660; // @[Modules.scala 143:103:@21195.4]
  wire [4:0] _T_74661; // @[Modules.scala 143:103:@21196.4]
  wire [4:0] _T_74662; // @[Modules.scala 143:103:@21197.4]
  wire [5:0] _GEN_492; // @[Modules.scala 143:103:@21201.4]
  wire [6:0] _T_74667; // @[Modules.scala 143:103:@21201.4]
  wire [5:0] _T_74668; // @[Modules.scala 143:103:@21202.4]
  wire [5:0] _T_74669; // @[Modules.scala 143:103:@21203.4]
  wire [6:0] _T_74674; // @[Modules.scala 143:103:@21207.4]
  wire [5:0] _T_74675; // @[Modules.scala 143:103:@21208.4]
  wire [5:0] _T_74676; // @[Modules.scala 143:103:@21209.4]
  wire [5:0] _GEN_494; // @[Modules.scala 143:103:@21213.4]
  wire [6:0] _T_74681; // @[Modules.scala 143:103:@21213.4]
  wire [5:0] _T_74682; // @[Modules.scala 143:103:@21214.4]
  wire [5:0] _T_74683; // @[Modules.scala 143:103:@21215.4]
  wire [6:0] _T_74730; // @[Modules.scala 143:103:@21255.4]
  wire [5:0] _T_74731; // @[Modules.scala 143:103:@21256.4]
  wire [5:0] _T_74732; // @[Modules.scala 143:103:@21257.4]
  wire [5:0] _T_74737; // @[Modules.scala 143:103:@21261.4]
  wire [4:0] _T_74738; // @[Modules.scala 143:103:@21262.4]
  wire [4:0] _T_74739; // @[Modules.scala 143:103:@21263.4]
  wire [5:0] _GEN_497; // @[Modules.scala 143:103:@21327.4]
  wire [6:0] _T_74814; // @[Modules.scala 143:103:@21327.4]
  wire [5:0] _T_74815; // @[Modules.scala 143:103:@21328.4]
  wire [5:0] _T_74816; // @[Modules.scala 143:103:@21329.4]
  wire [13:0] buffer_6_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74820; // @[Modules.scala 160:64:@21335.4]
  wire [13:0] _T_74821; // @[Modules.scala 160:64:@21336.4]
  wire [13:0] buffer_6_317; // @[Modules.scala 160:64:@21337.4]
  wire [13:0] buffer_6_4; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74823; // @[Modules.scala 160:64:@21339.4]
  wire [13:0] _T_74824; // @[Modules.scala 160:64:@21340.4]
  wire [13:0] buffer_6_318; // @[Modules.scala 160:64:@21341.4]
  wire [13:0] buffer_6_8; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74829; // @[Modules.scala 160:64:@21347.4]
  wire [13:0] _T_74830; // @[Modules.scala 160:64:@21348.4]
  wire [13:0] buffer_6_320; // @[Modules.scala 160:64:@21349.4]
  wire [13:0] buffer_6_10; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74832; // @[Modules.scala 160:64:@21351.4]
  wire [13:0] _T_74833; // @[Modules.scala 160:64:@21352.4]
  wire [13:0] buffer_6_321; // @[Modules.scala 160:64:@21353.4]
  wire [14:0] _T_74835; // @[Modules.scala 160:64:@21355.4]
  wire [13:0] _T_74836; // @[Modules.scala 160:64:@21356.4]
  wire [13:0] buffer_6_322; // @[Modules.scala 160:64:@21357.4]
  wire [13:0] buffer_6_20; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74847; // @[Modules.scala 160:64:@21371.4]
  wire [13:0] _T_74848; // @[Modules.scala 160:64:@21372.4]
  wire [13:0] buffer_6_326; // @[Modules.scala 160:64:@21373.4]
  wire [13:0] buffer_6_22; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74850; // @[Modules.scala 160:64:@21375.4]
  wire [13:0] _T_74851; // @[Modules.scala 160:64:@21376.4]
  wire [13:0] buffer_6_327; // @[Modules.scala 160:64:@21377.4]
  wire [13:0] buffer_6_25; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74853; // @[Modules.scala 160:64:@21379.4]
  wire [13:0] _T_74854; // @[Modules.scala 160:64:@21380.4]
  wire [13:0] buffer_6_328; // @[Modules.scala 160:64:@21381.4]
  wire [13:0] buffer_6_26; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74856; // @[Modules.scala 160:64:@21383.4]
  wire [13:0] _T_74857; // @[Modules.scala 160:64:@21384.4]
  wire [13:0] buffer_6_329; // @[Modules.scala 160:64:@21385.4]
  wire [13:0] buffer_6_29; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74859; // @[Modules.scala 160:64:@21387.4]
  wire [13:0] _T_74860; // @[Modules.scala 160:64:@21388.4]
  wire [13:0] buffer_6_330; // @[Modules.scala 160:64:@21389.4]
  wire [13:0] buffer_6_30; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74862; // @[Modules.scala 160:64:@21391.4]
  wire [13:0] _T_74863; // @[Modules.scala 160:64:@21392.4]
  wire [13:0] buffer_6_331; // @[Modules.scala 160:64:@21393.4]
  wire [13:0] buffer_6_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74865; // @[Modules.scala 160:64:@21395.4]
  wire [13:0] _T_74866; // @[Modules.scala 160:64:@21396.4]
  wire [13:0] buffer_6_332; // @[Modules.scala 160:64:@21397.4]
  wire [13:0] buffer_6_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74868; // @[Modules.scala 160:64:@21399.4]
  wire [13:0] _T_74869; // @[Modules.scala 160:64:@21400.4]
  wire [13:0] buffer_6_333; // @[Modules.scala 160:64:@21401.4]
  wire [13:0] buffer_6_39; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74874; // @[Modules.scala 160:64:@21407.4]
  wire [13:0] _T_74875; // @[Modules.scala 160:64:@21408.4]
  wire [13:0] buffer_6_335; // @[Modules.scala 160:64:@21409.4]
  wire [13:0] buffer_6_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74883; // @[Modules.scala 160:64:@21419.4]
  wire [13:0] _T_74884; // @[Modules.scala 160:64:@21420.4]
  wire [13:0] buffer_6_338; // @[Modules.scala 160:64:@21421.4]
  wire [13:0] buffer_6_46; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74886; // @[Modules.scala 160:64:@21423.4]
  wire [13:0] _T_74887; // @[Modules.scala 160:64:@21424.4]
  wire [13:0] buffer_6_339; // @[Modules.scala 160:64:@21425.4]
  wire [13:0] buffer_6_50; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74892; // @[Modules.scala 160:64:@21431.4]
  wire [13:0] _T_74893; // @[Modules.scala 160:64:@21432.4]
  wire [13:0] buffer_6_341; // @[Modules.scala 160:64:@21433.4]
  wire [14:0] _T_74895; // @[Modules.scala 160:64:@21435.4]
  wire [13:0] _T_74896; // @[Modules.scala 160:64:@21436.4]
  wire [13:0] buffer_6_342; // @[Modules.scala 160:64:@21437.4]
  wire [14:0] _T_74898; // @[Modules.scala 160:64:@21439.4]
  wire [13:0] _T_74899; // @[Modules.scala 160:64:@21440.4]
  wire [13:0] buffer_6_343; // @[Modules.scala 160:64:@21441.4]
  wire [13:0] buffer_6_56; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74901; // @[Modules.scala 160:64:@21443.4]
  wire [13:0] _T_74902; // @[Modules.scala 160:64:@21444.4]
  wire [13:0] buffer_6_344; // @[Modules.scala 160:64:@21445.4]
  wire [13:0] buffer_6_58; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74904; // @[Modules.scala 160:64:@21447.4]
  wire [13:0] _T_74905; // @[Modules.scala 160:64:@21448.4]
  wire [13:0] buffer_6_345; // @[Modules.scala 160:64:@21449.4]
  wire [13:0] buffer_6_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74907; // @[Modules.scala 160:64:@21451.4]
  wire [13:0] _T_74908; // @[Modules.scala 160:64:@21452.4]
  wire [13:0] buffer_6_346; // @[Modules.scala 160:64:@21453.4]
  wire [13:0] buffer_6_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74910; // @[Modules.scala 160:64:@21455.4]
  wire [13:0] _T_74911; // @[Modules.scala 160:64:@21456.4]
  wire [13:0] buffer_6_347; // @[Modules.scala 160:64:@21457.4]
  wire [13:0] buffer_6_66; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74916; // @[Modules.scala 160:64:@21463.4]
  wire [13:0] _T_74917; // @[Modules.scala 160:64:@21464.4]
  wire [13:0] buffer_6_349; // @[Modules.scala 160:64:@21465.4]
  wire [13:0] buffer_6_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74919; // @[Modules.scala 160:64:@21467.4]
  wire [13:0] _T_74920; // @[Modules.scala 160:64:@21468.4]
  wire [13:0] buffer_6_350; // @[Modules.scala 160:64:@21469.4]
  wire [13:0] buffer_6_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74922; // @[Modules.scala 160:64:@21471.4]
  wire [13:0] _T_74923; // @[Modules.scala 160:64:@21472.4]
  wire [13:0] buffer_6_351; // @[Modules.scala 160:64:@21473.4]
  wire [13:0] buffer_6_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74925; // @[Modules.scala 160:64:@21475.4]
  wire [13:0] _T_74926; // @[Modules.scala 160:64:@21476.4]
  wire [13:0] buffer_6_352; // @[Modules.scala 160:64:@21477.4]
  wire [13:0] buffer_6_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74928; // @[Modules.scala 160:64:@21479.4]
  wire [13:0] _T_74929; // @[Modules.scala 160:64:@21480.4]
  wire [13:0] buffer_6_353; // @[Modules.scala 160:64:@21481.4]
  wire [13:0] buffer_6_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74931; // @[Modules.scala 160:64:@21483.4]
  wire [13:0] _T_74932; // @[Modules.scala 160:64:@21484.4]
  wire [13:0] buffer_6_354; // @[Modules.scala 160:64:@21485.4]
  wire [13:0] buffer_6_78; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74934; // @[Modules.scala 160:64:@21487.4]
  wire [13:0] _T_74935; // @[Modules.scala 160:64:@21488.4]
  wire [13:0] buffer_6_355; // @[Modules.scala 160:64:@21489.4]
  wire [13:0] buffer_6_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74937; // @[Modules.scala 160:64:@21491.4]
  wire [13:0] _T_74938; // @[Modules.scala 160:64:@21492.4]
  wire [13:0] buffer_6_356; // @[Modules.scala 160:64:@21493.4]
  wire [13:0] buffer_6_82; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74940; // @[Modules.scala 160:64:@21495.4]
  wire [13:0] _T_74941; // @[Modules.scala 160:64:@21496.4]
  wire [13:0] buffer_6_357; // @[Modules.scala 160:64:@21497.4]
  wire [13:0] buffer_6_88; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74949; // @[Modules.scala 160:64:@21507.4]
  wire [13:0] _T_74950; // @[Modules.scala 160:64:@21508.4]
  wire [13:0] buffer_6_360; // @[Modules.scala 160:64:@21509.4]
  wire [13:0] buffer_6_90; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74952; // @[Modules.scala 160:64:@21511.4]
  wire [13:0] _T_74953; // @[Modules.scala 160:64:@21512.4]
  wire [13:0] buffer_6_361; // @[Modules.scala 160:64:@21513.4]
  wire [13:0] buffer_6_94; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74958; // @[Modules.scala 160:64:@21519.4]
  wire [13:0] _T_74959; // @[Modules.scala 160:64:@21520.4]
  wire [13:0] buffer_6_363; // @[Modules.scala 160:64:@21521.4]
  wire [13:0] buffer_6_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74961; // @[Modules.scala 160:64:@21523.4]
  wire [13:0] _T_74962; // @[Modules.scala 160:64:@21524.4]
  wire [13:0] buffer_6_364; // @[Modules.scala 160:64:@21525.4]
  wire [14:0] _T_74964; // @[Modules.scala 160:64:@21527.4]
  wire [13:0] _T_74965; // @[Modules.scala 160:64:@21528.4]
  wire [13:0] buffer_6_365; // @[Modules.scala 160:64:@21529.4]
  wire [13:0] buffer_6_100; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_101; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74967; // @[Modules.scala 160:64:@21531.4]
  wire [13:0] _T_74968; // @[Modules.scala 160:64:@21532.4]
  wire [13:0] buffer_6_366; // @[Modules.scala 160:64:@21533.4]
  wire [13:0] buffer_6_102; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74970; // @[Modules.scala 160:64:@21535.4]
  wire [13:0] _T_74971; // @[Modules.scala 160:64:@21536.4]
  wire [13:0] buffer_6_367; // @[Modules.scala 160:64:@21537.4]
  wire [13:0] buffer_6_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74973; // @[Modules.scala 160:64:@21539.4]
  wire [13:0] _T_74974; // @[Modules.scala 160:64:@21540.4]
  wire [13:0] buffer_6_368; // @[Modules.scala 160:64:@21541.4]
  wire [14:0] _T_74976; // @[Modules.scala 160:64:@21543.4]
  wire [13:0] _T_74977; // @[Modules.scala 160:64:@21544.4]
  wire [13:0] buffer_6_369; // @[Modules.scala 160:64:@21545.4]
  wire [14:0] _T_74979; // @[Modules.scala 160:64:@21547.4]
  wire [13:0] _T_74980; // @[Modules.scala 160:64:@21548.4]
  wire [13:0] buffer_6_370; // @[Modules.scala 160:64:@21549.4]
  wire [13:0] buffer_6_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74982; // @[Modules.scala 160:64:@21551.4]
  wire [13:0] _T_74983; // @[Modules.scala 160:64:@21552.4]
  wire [13:0] buffer_6_371; // @[Modules.scala 160:64:@21553.4]
  wire [13:0] buffer_6_112; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74985; // @[Modules.scala 160:64:@21555.4]
  wire [13:0] _T_74986; // @[Modules.scala 160:64:@21556.4]
  wire [13:0] buffer_6_372; // @[Modules.scala 160:64:@21557.4]
  wire [13:0] buffer_6_114; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74988; // @[Modules.scala 160:64:@21559.4]
  wire [13:0] _T_74989; // @[Modules.scala 160:64:@21560.4]
  wire [13:0] buffer_6_373; // @[Modules.scala 160:64:@21561.4]
  wire [14:0] _T_74991; // @[Modules.scala 160:64:@21563.4]
  wire [13:0] _T_74992; // @[Modules.scala 160:64:@21564.4]
  wire [13:0] buffer_6_374; // @[Modules.scala 160:64:@21565.4]
  wire [13:0] buffer_6_118; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_74994; // @[Modules.scala 160:64:@21567.4]
  wire [13:0] _T_74995; // @[Modules.scala 160:64:@21568.4]
  wire [13:0] buffer_6_375; // @[Modules.scala 160:64:@21569.4]
  wire [14:0] _T_74997; // @[Modules.scala 160:64:@21571.4]
  wire [13:0] _T_74998; // @[Modules.scala 160:64:@21572.4]
  wire [13:0] buffer_6_376; // @[Modules.scala 160:64:@21573.4]
  wire [13:0] buffer_6_122; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75000; // @[Modules.scala 160:64:@21575.4]
  wire [13:0] _T_75001; // @[Modules.scala 160:64:@21576.4]
  wire [13:0] buffer_6_377; // @[Modules.scala 160:64:@21577.4]
  wire [14:0] _T_75003; // @[Modules.scala 160:64:@21579.4]
  wire [13:0] _T_75004; // @[Modules.scala 160:64:@21580.4]
  wire [13:0] buffer_6_378; // @[Modules.scala 160:64:@21581.4]
  wire [14:0] _T_75006; // @[Modules.scala 160:64:@21583.4]
  wire [13:0] _T_75007; // @[Modules.scala 160:64:@21584.4]
  wire [13:0] buffer_6_379; // @[Modules.scala 160:64:@21585.4]
  wire [13:0] buffer_6_128; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75009; // @[Modules.scala 160:64:@21587.4]
  wire [13:0] _T_75010; // @[Modules.scala 160:64:@21588.4]
  wire [13:0] buffer_6_380; // @[Modules.scala 160:64:@21589.4]
  wire [13:0] buffer_6_130; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75012; // @[Modules.scala 160:64:@21591.4]
  wire [13:0] _T_75013; // @[Modules.scala 160:64:@21592.4]
  wire [13:0] buffer_6_381; // @[Modules.scala 160:64:@21593.4]
  wire [14:0] _T_75015; // @[Modules.scala 160:64:@21595.4]
  wire [13:0] _T_75016; // @[Modules.scala 160:64:@21596.4]
  wire [13:0] buffer_6_382; // @[Modules.scala 160:64:@21597.4]
  wire [13:0] buffer_6_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75018; // @[Modules.scala 160:64:@21599.4]
  wire [13:0] _T_75019; // @[Modules.scala 160:64:@21600.4]
  wire [13:0] buffer_6_383; // @[Modules.scala 160:64:@21601.4]
  wire [13:0] buffer_6_136; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75021; // @[Modules.scala 160:64:@21603.4]
  wire [13:0] _T_75022; // @[Modules.scala 160:64:@21604.4]
  wire [13:0] buffer_6_384; // @[Modules.scala 160:64:@21605.4]
  wire [13:0] buffer_6_140; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75027; // @[Modules.scala 160:64:@21611.4]
  wire [13:0] _T_75028; // @[Modules.scala 160:64:@21612.4]
  wire [13:0] buffer_6_386; // @[Modules.scala 160:64:@21613.4]
  wire [13:0] buffer_6_144; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75033; // @[Modules.scala 160:64:@21619.4]
  wire [13:0] _T_75034; // @[Modules.scala 160:64:@21620.4]
  wire [13:0] buffer_6_388; // @[Modules.scala 160:64:@21621.4]
  wire [13:0] buffer_6_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75039; // @[Modules.scala 160:64:@21627.4]
  wire [13:0] _T_75040; // @[Modules.scala 160:64:@21628.4]
  wire [13:0] buffer_6_390; // @[Modules.scala 160:64:@21629.4]
  wire [13:0] buffer_6_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75042; // @[Modules.scala 160:64:@21631.4]
  wire [13:0] _T_75043; // @[Modules.scala 160:64:@21632.4]
  wire [13:0] buffer_6_391; // @[Modules.scala 160:64:@21633.4]
  wire [14:0] _T_75045; // @[Modules.scala 160:64:@21635.4]
  wire [13:0] _T_75046; // @[Modules.scala 160:64:@21636.4]
  wire [13:0] buffer_6_392; // @[Modules.scala 160:64:@21637.4]
  wire [14:0] _T_75048; // @[Modules.scala 160:64:@21639.4]
  wire [13:0] _T_75049; // @[Modules.scala 160:64:@21640.4]
  wire [13:0] buffer_6_393; // @[Modules.scala 160:64:@21641.4]
  wire [14:0] _T_75051; // @[Modules.scala 160:64:@21643.4]
  wire [13:0] _T_75052; // @[Modules.scala 160:64:@21644.4]
  wire [13:0] buffer_6_394; // @[Modules.scala 160:64:@21645.4]
  wire [14:0] _T_75054; // @[Modules.scala 160:64:@21647.4]
  wire [13:0] _T_75055; // @[Modules.scala 160:64:@21648.4]
  wire [13:0] buffer_6_395; // @[Modules.scala 160:64:@21649.4]
  wire [14:0] _T_75057; // @[Modules.scala 160:64:@21651.4]
  wire [13:0] _T_75058; // @[Modules.scala 160:64:@21652.4]
  wire [13:0] buffer_6_396; // @[Modules.scala 160:64:@21653.4]
  wire [14:0] _T_75060; // @[Modules.scala 160:64:@21655.4]
  wire [13:0] _T_75061; // @[Modules.scala 160:64:@21656.4]
  wire [13:0] buffer_6_397; // @[Modules.scala 160:64:@21657.4]
  wire [13:0] buffer_6_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75063; // @[Modules.scala 160:64:@21659.4]
  wire [13:0] _T_75064; // @[Modules.scala 160:64:@21660.4]
  wire [13:0] buffer_6_398; // @[Modules.scala 160:64:@21661.4]
  wire [14:0] _T_75066; // @[Modules.scala 160:64:@21663.4]
  wire [13:0] _T_75067; // @[Modules.scala 160:64:@21664.4]
  wire [13:0] buffer_6_399; // @[Modules.scala 160:64:@21665.4]
  wire [13:0] buffer_6_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75069; // @[Modules.scala 160:64:@21667.4]
  wire [13:0] _T_75070; // @[Modules.scala 160:64:@21668.4]
  wire [13:0] buffer_6_400; // @[Modules.scala 160:64:@21669.4]
  wire [13:0] buffer_6_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75072; // @[Modules.scala 160:64:@21671.4]
  wire [13:0] _T_75073; // @[Modules.scala 160:64:@21672.4]
  wire [13:0] buffer_6_401; // @[Modules.scala 160:64:@21673.4]
  wire [14:0] _T_75075; // @[Modules.scala 160:64:@21675.4]
  wire [13:0] _T_75076; // @[Modules.scala 160:64:@21676.4]
  wire [13:0] buffer_6_402; // @[Modules.scala 160:64:@21677.4]
  wire [13:0] buffer_6_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75078; // @[Modules.scala 160:64:@21679.4]
  wire [13:0] _T_75079; // @[Modules.scala 160:64:@21680.4]
  wire [13:0] buffer_6_403; // @[Modules.scala 160:64:@21681.4]
  wire [13:0] buffer_6_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75081; // @[Modules.scala 160:64:@21683.4]
  wire [13:0] _T_75082; // @[Modules.scala 160:64:@21684.4]
  wire [13:0] buffer_6_404; // @[Modules.scala 160:64:@21685.4]
  wire [13:0] buffer_6_178; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75084; // @[Modules.scala 160:64:@21687.4]
  wire [13:0] _T_75085; // @[Modules.scala 160:64:@21688.4]
  wire [13:0] buffer_6_405; // @[Modules.scala 160:64:@21689.4]
  wire [13:0] buffer_6_180; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75087; // @[Modules.scala 160:64:@21691.4]
  wire [13:0] _T_75088; // @[Modules.scala 160:64:@21692.4]
  wire [13:0] buffer_6_406; // @[Modules.scala 160:64:@21693.4]
  wire [13:0] buffer_6_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75090; // @[Modules.scala 160:64:@21695.4]
  wire [13:0] _T_75091; // @[Modules.scala 160:64:@21696.4]
  wire [13:0] buffer_6_407; // @[Modules.scala 160:64:@21697.4]
  wire [13:0] buffer_6_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75093; // @[Modules.scala 160:64:@21699.4]
  wire [13:0] _T_75094; // @[Modules.scala 160:64:@21700.4]
  wire [13:0] buffer_6_408; // @[Modules.scala 160:64:@21701.4]
  wire [14:0] _T_75096; // @[Modules.scala 160:64:@21703.4]
  wire [13:0] _T_75097; // @[Modules.scala 160:64:@21704.4]
  wire [13:0] buffer_6_409; // @[Modules.scala 160:64:@21705.4]
  wire [13:0] buffer_6_188; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75099; // @[Modules.scala 160:64:@21707.4]
  wire [13:0] _T_75100; // @[Modules.scala 160:64:@21708.4]
  wire [13:0] buffer_6_410; // @[Modules.scala 160:64:@21709.4]
  wire [13:0] buffer_6_190; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75102; // @[Modules.scala 160:64:@21711.4]
  wire [13:0] _T_75103; // @[Modules.scala 160:64:@21712.4]
  wire [13:0] buffer_6_411; // @[Modules.scala 160:64:@21713.4]
  wire [13:0] buffer_6_192; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75105; // @[Modules.scala 160:64:@21715.4]
  wire [13:0] _T_75106; // @[Modules.scala 160:64:@21716.4]
  wire [13:0] buffer_6_412; // @[Modules.scala 160:64:@21717.4]
  wire [13:0] buffer_6_194; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75108; // @[Modules.scala 160:64:@21719.4]
  wire [13:0] _T_75109; // @[Modules.scala 160:64:@21720.4]
  wire [13:0] buffer_6_413; // @[Modules.scala 160:64:@21721.4]
  wire [14:0] _T_75111; // @[Modules.scala 160:64:@21723.4]
  wire [13:0] _T_75112; // @[Modules.scala 160:64:@21724.4]
  wire [13:0] buffer_6_414; // @[Modules.scala 160:64:@21725.4]
  wire [13:0] buffer_6_198; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75114; // @[Modules.scala 160:64:@21727.4]
  wire [13:0] _T_75115; // @[Modules.scala 160:64:@21728.4]
  wire [13:0] buffer_6_415; // @[Modules.scala 160:64:@21729.4]
  wire [13:0] buffer_6_200; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75117; // @[Modules.scala 160:64:@21731.4]
  wire [13:0] _T_75118; // @[Modules.scala 160:64:@21732.4]
  wire [13:0] buffer_6_416; // @[Modules.scala 160:64:@21733.4]
  wire [13:0] buffer_6_202; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75120; // @[Modules.scala 160:64:@21735.4]
  wire [13:0] _T_75121; // @[Modules.scala 160:64:@21736.4]
  wire [13:0] buffer_6_417; // @[Modules.scala 160:64:@21737.4]
  wire [14:0] _T_75123; // @[Modules.scala 160:64:@21739.4]
  wire [13:0] _T_75124; // @[Modules.scala 160:64:@21740.4]
  wire [13:0] buffer_6_418; // @[Modules.scala 160:64:@21741.4]
  wire [14:0] _T_75126; // @[Modules.scala 160:64:@21743.4]
  wire [13:0] _T_75127; // @[Modules.scala 160:64:@21744.4]
  wire [13:0] buffer_6_419; // @[Modules.scala 160:64:@21745.4]
  wire [14:0] _T_75129; // @[Modules.scala 160:64:@21747.4]
  wire [13:0] _T_75130; // @[Modules.scala 160:64:@21748.4]
  wire [13:0] buffer_6_420; // @[Modules.scala 160:64:@21749.4]
  wire [13:0] buffer_6_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75132; // @[Modules.scala 160:64:@21751.4]
  wire [13:0] _T_75133; // @[Modules.scala 160:64:@21752.4]
  wire [13:0] buffer_6_421; // @[Modules.scala 160:64:@21753.4]
  wire [13:0] buffer_6_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75135; // @[Modules.scala 160:64:@21755.4]
  wire [13:0] _T_75136; // @[Modules.scala 160:64:@21756.4]
  wire [13:0] buffer_6_422; // @[Modules.scala 160:64:@21757.4]
  wire [13:0] buffer_6_220; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75147; // @[Modules.scala 160:64:@21771.4]
  wire [13:0] _T_75148; // @[Modules.scala 160:64:@21772.4]
  wire [13:0] buffer_6_426; // @[Modules.scala 160:64:@21773.4]
  wire [13:0] buffer_6_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75150; // @[Modules.scala 160:64:@21775.4]
  wire [13:0] _T_75151; // @[Modules.scala 160:64:@21776.4]
  wire [13:0] buffer_6_427; // @[Modules.scala 160:64:@21777.4]
  wire [13:0] buffer_6_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75153; // @[Modules.scala 160:64:@21779.4]
  wire [13:0] _T_75154; // @[Modules.scala 160:64:@21780.4]
  wire [13:0] buffer_6_428; // @[Modules.scala 160:64:@21781.4]
  wire [13:0] buffer_6_226; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75156; // @[Modules.scala 160:64:@21783.4]
  wire [13:0] _T_75157; // @[Modules.scala 160:64:@21784.4]
  wire [13:0] buffer_6_429; // @[Modules.scala 160:64:@21785.4]
  wire [13:0] buffer_6_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75159; // @[Modules.scala 160:64:@21787.4]
  wire [13:0] _T_75160; // @[Modules.scala 160:64:@21788.4]
  wire [13:0] buffer_6_430; // @[Modules.scala 160:64:@21789.4]
  wire [13:0] buffer_6_230; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75162; // @[Modules.scala 160:64:@21791.4]
  wire [13:0] _T_75163; // @[Modules.scala 160:64:@21792.4]
  wire [13:0] buffer_6_431; // @[Modules.scala 160:64:@21793.4]
  wire [13:0] buffer_6_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75165; // @[Modules.scala 160:64:@21795.4]
  wire [13:0] _T_75166; // @[Modules.scala 160:64:@21796.4]
  wire [13:0] buffer_6_432; // @[Modules.scala 160:64:@21797.4]
  wire [14:0] _T_75168; // @[Modules.scala 160:64:@21799.4]
  wire [13:0] _T_75169; // @[Modules.scala 160:64:@21800.4]
  wire [13:0] buffer_6_433; // @[Modules.scala 160:64:@21801.4]
  wire [13:0] buffer_6_236; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75171; // @[Modules.scala 160:64:@21803.4]
  wire [13:0] _T_75172; // @[Modules.scala 160:64:@21804.4]
  wire [13:0] buffer_6_434; // @[Modules.scala 160:64:@21805.4]
  wire [14:0] _T_75174; // @[Modules.scala 160:64:@21807.4]
  wire [13:0] _T_75175; // @[Modules.scala 160:64:@21808.4]
  wire [13:0] buffer_6_435; // @[Modules.scala 160:64:@21809.4]
  wire [13:0] buffer_6_240; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75177; // @[Modules.scala 160:64:@21811.4]
  wire [13:0] _T_75178; // @[Modules.scala 160:64:@21812.4]
  wire [13:0] buffer_6_436; // @[Modules.scala 160:64:@21813.4]
  wire [13:0] buffer_6_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75180; // @[Modules.scala 160:64:@21815.4]
  wire [13:0] _T_75181; // @[Modules.scala 160:64:@21816.4]
  wire [13:0] buffer_6_437; // @[Modules.scala 160:64:@21817.4]
  wire [13:0] buffer_6_244; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75183; // @[Modules.scala 160:64:@21819.4]
  wire [13:0] _T_75184; // @[Modules.scala 160:64:@21820.4]
  wire [13:0] buffer_6_438; // @[Modules.scala 160:64:@21821.4]
  wire [13:0] buffer_6_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75186; // @[Modules.scala 160:64:@21823.4]
  wire [13:0] _T_75187; // @[Modules.scala 160:64:@21824.4]
  wire [13:0] buffer_6_439; // @[Modules.scala 160:64:@21825.4]
  wire [13:0] buffer_6_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75189; // @[Modules.scala 160:64:@21827.4]
  wire [13:0] _T_75190; // @[Modules.scala 160:64:@21828.4]
  wire [13:0] buffer_6_440; // @[Modules.scala 160:64:@21829.4]
  wire [13:0] buffer_6_250; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75192; // @[Modules.scala 160:64:@21831.4]
  wire [13:0] _T_75193; // @[Modules.scala 160:64:@21832.4]
  wire [13:0] buffer_6_441; // @[Modules.scala 160:64:@21833.4]
  wire [13:0] buffer_6_252; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75195; // @[Modules.scala 160:64:@21835.4]
  wire [13:0] _T_75196; // @[Modules.scala 160:64:@21836.4]
  wire [13:0] buffer_6_442; // @[Modules.scala 160:64:@21837.4]
  wire [14:0] _T_75198; // @[Modules.scala 160:64:@21839.4]
  wire [13:0] _T_75199; // @[Modules.scala 160:64:@21840.4]
  wire [13:0] buffer_6_443; // @[Modules.scala 160:64:@21841.4]
  wire [13:0] buffer_6_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75201; // @[Modules.scala 160:64:@21843.4]
  wire [13:0] _T_75202; // @[Modules.scala 160:64:@21844.4]
  wire [13:0] buffer_6_444; // @[Modules.scala 160:64:@21845.4]
  wire [13:0] buffer_6_258; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75204; // @[Modules.scala 160:64:@21847.4]
  wire [13:0] _T_75205; // @[Modules.scala 160:64:@21848.4]
  wire [13:0] buffer_6_445; // @[Modules.scala 160:64:@21849.4]
  wire [13:0] buffer_6_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75207; // @[Modules.scala 160:64:@21851.4]
  wire [13:0] _T_75208; // @[Modules.scala 160:64:@21852.4]
  wire [13:0] buffer_6_446; // @[Modules.scala 160:64:@21853.4]
  wire [13:0] buffer_6_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75210; // @[Modules.scala 160:64:@21855.4]
  wire [13:0] _T_75211; // @[Modules.scala 160:64:@21856.4]
  wire [13:0] buffer_6_447; // @[Modules.scala 160:64:@21857.4]
  wire [13:0] buffer_6_264; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75213; // @[Modules.scala 160:64:@21859.4]
  wire [13:0] _T_75214; // @[Modules.scala 160:64:@21860.4]
  wire [13:0] buffer_6_448; // @[Modules.scala 160:64:@21861.4]
  wire [13:0] buffer_6_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75219; // @[Modules.scala 160:64:@21867.4]
  wire [13:0] _T_75220; // @[Modules.scala 160:64:@21868.4]
  wire [13:0] buffer_6_450; // @[Modules.scala 160:64:@21869.4]
  wire [13:0] buffer_6_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75222; // @[Modules.scala 160:64:@21871.4]
  wire [13:0] _T_75223; // @[Modules.scala 160:64:@21872.4]
  wire [13:0] buffer_6_451; // @[Modules.scala 160:64:@21873.4]
  wire [13:0] buffer_6_272; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75225; // @[Modules.scala 160:64:@21875.4]
  wire [13:0] _T_75226; // @[Modules.scala 160:64:@21876.4]
  wire [13:0] buffer_6_452; // @[Modules.scala 160:64:@21877.4]
  wire [13:0] buffer_6_274; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75228; // @[Modules.scala 160:64:@21879.4]
  wire [13:0] _T_75229; // @[Modules.scala 160:64:@21880.4]
  wire [13:0] buffer_6_453; // @[Modules.scala 160:64:@21881.4]
  wire [14:0] _T_75231; // @[Modules.scala 160:64:@21883.4]
  wire [13:0] _T_75232; // @[Modules.scala 160:64:@21884.4]
  wire [13:0] buffer_6_454; // @[Modules.scala 160:64:@21885.4]
  wire [13:0] buffer_6_278; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75234; // @[Modules.scala 160:64:@21887.4]
  wire [13:0] _T_75235; // @[Modules.scala 160:64:@21888.4]
  wire [13:0] buffer_6_455; // @[Modules.scala 160:64:@21889.4]
  wire [13:0] buffer_6_280; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75237; // @[Modules.scala 160:64:@21891.4]
  wire [13:0] _T_75238; // @[Modules.scala 160:64:@21892.4]
  wire [13:0] buffer_6_456; // @[Modules.scala 160:64:@21893.4]
  wire [13:0] buffer_6_282; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75240; // @[Modules.scala 160:64:@21895.4]
  wire [13:0] _T_75241; // @[Modules.scala 160:64:@21896.4]
  wire [13:0] buffer_6_457; // @[Modules.scala 160:64:@21897.4]
  wire [13:0] buffer_6_284; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_285; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75243; // @[Modules.scala 160:64:@21899.4]
  wire [13:0] _T_75244; // @[Modules.scala 160:64:@21900.4]
  wire [13:0] buffer_6_458; // @[Modules.scala 160:64:@21901.4]
  wire [13:0] buffer_6_286; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75246; // @[Modules.scala 160:64:@21903.4]
  wire [13:0] _T_75247; // @[Modules.scala 160:64:@21904.4]
  wire [13:0] buffer_6_459; // @[Modules.scala 160:64:@21905.4]
  wire [13:0] buffer_6_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75249; // @[Modules.scala 160:64:@21907.4]
  wire [13:0] _T_75250; // @[Modules.scala 160:64:@21908.4]
  wire [13:0] buffer_6_460; // @[Modules.scala 160:64:@21909.4]
  wire [13:0] buffer_6_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75252; // @[Modules.scala 160:64:@21911.4]
  wire [13:0] _T_75253; // @[Modules.scala 160:64:@21912.4]
  wire [13:0] buffer_6_461; // @[Modules.scala 160:64:@21913.4]
  wire [13:0] buffer_6_292; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75255; // @[Modules.scala 160:64:@21915.4]
  wire [13:0] _T_75256; // @[Modules.scala 160:64:@21916.4]
  wire [13:0] buffer_6_462; // @[Modules.scala 160:64:@21917.4]
  wire [13:0] buffer_6_294; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_6_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75258; // @[Modules.scala 160:64:@21919.4]
  wire [13:0] _T_75259; // @[Modules.scala 160:64:@21920.4]
  wire [13:0] buffer_6_463; // @[Modules.scala 160:64:@21921.4]
  wire [13:0] buffer_6_296; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75261; // @[Modules.scala 160:64:@21923.4]
  wire [13:0] _T_75262; // @[Modules.scala 160:64:@21924.4]
  wire [13:0] buffer_6_464; // @[Modules.scala 160:64:@21925.4]
  wire [13:0] buffer_6_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75270; // @[Modules.scala 160:64:@21935.4]
  wire [13:0] _T_75271; // @[Modules.scala 160:64:@21936.4]
  wire [13:0] buffer_6_467; // @[Modules.scala 160:64:@21937.4]
  wire [13:0] buffer_6_304; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75273; // @[Modules.scala 160:64:@21939.4]
  wire [13:0] _T_75274; // @[Modules.scala 160:64:@21940.4]
  wire [13:0] buffer_6_468; // @[Modules.scala 160:64:@21941.4]
  wire [14:0] _T_75276; // @[Modules.scala 160:64:@21943.4]
  wire [13:0] _T_75277; // @[Modules.scala 160:64:@21944.4]
  wire [13:0] buffer_6_469; // @[Modules.scala 160:64:@21945.4]
  wire [14:0] _T_75279; // @[Modules.scala 160:64:@21947.4]
  wire [13:0] _T_75280; // @[Modules.scala 160:64:@21948.4]
  wire [13:0] buffer_6_470; // @[Modules.scala 160:64:@21949.4]
  wire [14:0] _T_75282; // @[Modules.scala 160:64:@21951.4]
  wire [13:0] _T_75283; // @[Modules.scala 160:64:@21952.4]
  wire [13:0] buffer_6_471; // @[Modules.scala 160:64:@21953.4]
  wire [14:0] _T_75285; // @[Modules.scala 160:64:@21955.4]
  wire [13:0] _T_75286; // @[Modules.scala 160:64:@21956.4]
  wire [13:0] buffer_6_472; // @[Modules.scala 160:64:@21957.4]
  wire [13:0] buffer_6_315; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_75288; // @[Modules.scala 160:64:@21959.4]
  wire [13:0] _T_75289; // @[Modules.scala 160:64:@21960.4]
  wire [13:0] buffer_6_473; // @[Modules.scala 160:64:@21961.4]
  wire [14:0] _T_75291; // @[Modules.scala 160:64:@21963.4]
  wire [13:0] _T_75292; // @[Modules.scala 160:64:@21964.4]
  wire [13:0] buffer_6_474; // @[Modules.scala 160:64:@21965.4]
  wire [14:0] _T_75294; // @[Modules.scala 160:64:@21967.4]
  wire [13:0] _T_75295; // @[Modules.scala 160:64:@21968.4]
  wire [13:0] buffer_6_475; // @[Modules.scala 160:64:@21969.4]
  wire [14:0] _T_75297; // @[Modules.scala 160:64:@21971.4]
  wire [13:0] _T_75298; // @[Modules.scala 160:64:@21972.4]
  wire [13:0] buffer_6_476; // @[Modules.scala 160:64:@21973.4]
  wire [14:0] _T_75300; // @[Modules.scala 160:64:@21975.4]
  wire [13:0] _T_75301; // @[Modules.scala 160:64:@21976.4]
  wire [13:0] buffer_6_477; // @[Modules.scala 160:64:@21977.4]
  wire [14:0] _T_75306; // @[Modules.scala 160:64:@21983.4]
  wire [13:0] _T_75307; // @[Modules.scala 160:64:@21984.4]
  wire [13:0] buffer_6_479; // @[Modules.scala 160:64:@21985.4]
  wire [14:0] _T_75309; // @[Modules.scala 160:64:@21987.4]
  wire [13:0] _T_75310; // @[Modules.scala 160:64:@21988.4]
  wire [13:0] buffer_6_480; // @[Modules.scala 160:64:@21989.4]
  wire [14:0] _T_75312; // @[Modules.scala 160:64:@21991.4]
  wire [13:0] _T_75313; // @[Modules.scala 160:64:@21992.4]
  wire [13:0] buffer_6_481; // @[Modules.scala 160:64:@21993.4]
  wire [14:0] _T_75315; // @[Modules.scala 160:64:@21995.4]
  wire [13:0] _T_75316; // @[Modules.scala 160:64:@21996.4]
  wire [13:0] buffer_6_482; // @[Modules.scala 160:64:@21997.4]
  wire [14:0] _T_75318; // @[Modules.scala 160:64:@21999.4]
  wire [13:0] _T_75319; // @[Modules.scala 160:64:@22000.4]
  wire [13:0] buffer_6_483; // @[Modules.scala 160:64:@22001.4]
  wire [14:0] _T_75321; // @[Modules.scala 160:64:@22003.4]
  wire [13:0] _T_75322; // @[Modules.scala 160:64:@22004.4]
  wire [13:0] buffer_6_484; // @[Modules.scala 160:64:@22005.4]
  wire [14:0] _T_75324; // @[Modules.scala 160:64:@22007.4]
  wire [13:0] _T_75325; // @[Modules.scala 160:64:@22008.4]
  wire [13:0] buffer_6_485; // @[Modules.scala 160:64:@22009.4]
  wire [14:0] _T_75327; // @[Modules.scala 160:64:@22011.4]
  wire [13:0] _T_75328; // @[Modules.scala 160:64:@22012.4]
  wire [13:0] buffer_6_486; // @[Modules.scala 160:64:@22013.4]
  wire [14:0] _T_75330; // @[Modules.scala 160:64:@22015.4]
  wire [13:0] _T_75331; // @[Modules.scala 160:64:@22016.4]
  wire [13:0] buffer_6_487; // @[Modules.scala 160:64:@22017.4]
  wire [14:0] _T_75333; // @[Modules.scala 160:64:@22019.4]
  wire [13:0] _T_75334; // @[Modules.scala 160:64:@22020.4]
  wire [13:0] buffer_6_488; // @[Modules.scala 160:64:@22021.4]
  wire [14:0] _T_75336; // @[Modules.scala 160:64:@22023.4]
  wire [13:0] _T_75337; // @[Modules.scala 160:64:@22024.4]
  wire [13:0] buffer_6_489; // @[Modules.scala 160:64:@22025.4]
  wire [14:0] _T_75339; // @[Modules.scala 160:64:@22027.4]
  wire [13:0] _T_75340; // @[Modules.scala 160:64:@22028.4]
  wire [13:0] buffer_6_490; // @[Modules.scala 160:64:@22029.4]
  wire [14:0] _T_75342; // @[Modules.scala 160:64:@22031.4]
  wire [13:0] _T_75343; // @[Modules.scala 160:64:@22032.4]
  wire [13:0] buffer_6_491; // @[Modules.scala 160:64:@22033.4]
  wire [14:0] _T_75345; // @[Modules.scala 160:64:@22035.4]
  wire [13:0] _T_75346; // @[Modules.scala 160:64:@22036.4]
  wire [13:0] buffer_6_492; // @[Modules.scala 160:64:@22037.4]
  wire [14:0] _T_75348; // @[Modules.scala 160:64:@22039.4]
  wire [13:0] _T_75349; // @[Modules.scala 160:64:@22040.4]
  wire [13:0] buffer_6_493; // @[Modules.scala 160:64:@22041.4]
  wire [14:0] _T_75351; // @[Modules.scala 160:64:@22043.4]
  wire [13:0] _T_75352; // @[Modules.scala 160:64:@22044.4]
  wire [13:0] buffer_6_494; // @[Modules.scala 160:64:@22045.4]
  wire [14:0] _T_75354; // @[Modules.scala 160:64:@22047.4]
  wire [13:0] _T_75355; // @[Modules.scala 160:64:@22048.4]
  wire [13:0] buffer_6_495; // @[Modules.scala 160:64:@22049.4]
  wire [14:0] _T_75357; // @[Modules.scala 160:64:@22051.4]
  wire [13:0] _T_75358; // @[Modules.scala 160:64:@22052.4]
  wire [13:0] buffer_6_496; // @[Modules.scala 160:64:@22053.4]
  wire [14:0] _T_75360; // @[Modules.scala 160:64:@22055.4]
  wire [13:0] _T_75361; // @[Modules.scala 160:64:@22056.4]
  wire [13:0] buffer_6_497; // @[Modules.scala 160:64:@22057.4]
  wire [14:0] _T_75363; // @[Modules.scala 160:64:@22059.4]
  wire [13:0] _T_75364; // @[Modules.scala 160:64:@22060.4]
  wire [13:0] buffer_6_498; // @[Modules.scala 160:64:@22061.4]
  wire [14:0] _T_75366; // @[Modules.scala 160:64:@22063.4]
  wire [13:0] _T_75367; // @[Modules.scala 160:64:@22064.4]
  wire [13:0] buffer_6_499; // @[Modules.scala 160:64:@22065.4]
  wire [14:0] _T_75369; // @[Modules.scala 160:64:@22067.4]
  wire [13:0] _T_75370; // @[Modules.scala 160:64:@22068.4]
  wire [13:0] buffer_6_500; // @[Modules.scala 160:64:@22069.4]
  wire [14:0] _T_75372; // @[Modules.scala 160:64:@22071.4]
  wire [13:0] _T_75373; // @[Modules.scala 160:64:@22072.4]
  wire [13:0] buffer_6_501; // @[Modules.scala 160:64:@22073.4]
  wire [14:0] _T_75375; // @[Modules.scala 160:64:@22075.4]
  wire [13:0] _T_75376; // @[Modules.scala 160:64:@22076.4]
  wire [13:0] buffer_6_502; // @[Modules.scala 160:64:@22077.4]
  wire [14:0] _T_75378; // @[Modules.scala 160:64:@22079.4]
  wire [13:0] _T_75379; // @[Modules.scala 160:64:@22080.4]
  wire [13:0] buffer_6_503; // @[Modules.scala 160:64:@22081.4]
  wire [14:0] _T_75381; // @[Modules.scala 160:64:@22083.4]
  wire [13:0] _T_75382; // @[Modules.scala 160:64:@22084.4]
  wire [13:0] buffer_6_504; // @[Modules.scala 160:64:@22085.4]
  wire [14:0] _T_75384; // @[Modules.scala 160:64:@22087.4]
  wire [13:0] _T_75385; // @[Modules.scala 160:64:@22088.4]
  wire [13:0] buffer_6_505; // @[Modules.scala 160:64:@22089.4]
  wire [14:0] _T_75387; // @[Modules.scala 160:64:@22091.4]
  wire [13:0] _T_75388; // @[Modules.scala 160:64:@22092.4]
  wire [13:0] buffer_6_506; // @[Modules.scala 160:64:@22093.4]
  wire [14:0] _T_75390; // @[Modules.scala 160:64:@22095.4]
  wire [13:0] _T_75391; // @[Modules.scala 160:64:@22096.4]
  wire [13:0] buffer_6_507; // @[Modules.scala 160:64:@22097.4]
  wire [14:0] _T_75393; // @[Modules.scala 160:64:@22099.4]
  wire [13:0] _T_75394; // @[Modules.scala 160:64:@22100.4]
  wire [13:0] buffer_6_508; // @[Modules.scala 160:64:@22101.4]
  wire [14:0] _T_75396; // @[Modules.scala 160:64:@22103.4]
  wire [13:0] _T_75397; // @[Modules.scala 160:64:@22104.4]
  wire [13:0] buffer_6_509; // @[Modules.scala 160:64:@22105.4]
  wire [14:0] _T_75399; // @[Modules.scala 160:64:@22107.4]
  wire [13:0] _T_75400; // @[Modules.scala 160:64:@22108.4]
  wire [13:0] buffer_6_510; // @[Modules.scala 160:64:@22109.4]
  wire [14:0] _T_75402; // @[Modules.scala 160:64:@22111.4]
  wire [13:0] _T_75403; // @[Modules.scala 160:64:@22112.4]
  wire [13:0] buffer_6_511; // @[Modules.scala 160:64:@22113.4]
  wire [14:0] _T_75405; // @[Modules.scala 160:64:@22115.4]
  wire [13:0] _T_75406; // @[Modules.scala 160:64:@22116.4]
  wire [13:0] buffer_6_512; // @[Modules.scala 160:64:@22117.4]
  wire [14:0] _T_75408; // @[Modules.scala 160:64:@22119.4]
  wire [13:0] _T_75409; // @[Modules.scala 160:64:@22120.4]
  wire [13:0] buffer_6_513; // @[Modules.scala 160:64:@22121.4]
  wire [14:0] _T_75411; // @[Modules.scala 160:64:@22123.4]
  wire [13:0] _T_75412; // @[Modules.scala 160:64:@22124.4]
  wire [13:0] buffer_6_514; // @[Modules.scala 160:64:@22125.4]
  wire [14:0] _T_75414; // @[Modules.scala 160:64:@22127.4]
  wire [13:0] _T_75415; // @[Modules.scala 160:64:@22128.4]
  wire [13:0] buffer_6_515; // @[Modules.scala 160:64:@22129.4]
  wire [14:0] _T_75417; // @[Modules.scala 160:64:@22131.4]
  wire [13:0] _T_75418; // @[Modules.scala 160:64:@22132.4]
  wire [13:0] buffer_6_516; // @[Modules.scala 160:64:@22133.4]
  wire [14:0] _T_75420; // @[Modules.scala 160:64:@22135.4]
  wire [13:0] _T_75421; // @[Modules.scala 160:64:@22136.4]
  wire [13:0] buffer_6_517; // @[Modules.scala 160:64:@22137.4]
  wire [14:0] _T_75423; // @[Modules.scala 160:64:@22139.4]
  wire [13:0] _T_75424; // @[Modules.scala 160:64:@22140.4]
  wire [13:0] buffer_6_518; // @[Modules.scala 160:64:@22141.4]
  wire [14:0] _T_75426; // @[Modules.scala 160:64:@22143.4]
  wire [13:0] _T_75427; // @[Modules.scala 160:64:@22144.4]
  wire [13:0] buffer_6_519; // @[Modules.scala 160:64:@22145.4]
  wire [14:0] _T_75429; // @[Modules.scala 160:64:@22147.4]
  wire [13:0] _T_75430; // @[Modules.scala 160:64:@22148.4]
  wire [13:0] buffer_6_520; // @[Modules.scala 160:64:@22149.4]
  wire [14:0] _T_75432; // @[Modules.scala 160:64:@22151.4]
  wire [13:0] _T_75433; // @[Modules.scala 160:64:@22152.4]
  wire [13:0] buffer_6_521; // @[Modules.scala 160:64:@22153.4]
  wire [14:0] _T_75435; // @[Modules.scala 160:64:@22155.4]
  wire [13:0] _T_75436; // @[Modules.scala 160:64:@22156.4]
  wire [13:0] buffer_6_522; // @[Modules.scala 160:64:@22157.4]
  wire [14:0] _T_75438; // @[Modules.scala 160:64:@22159.4]
  wire [13:0] _T_75439; // @[Modules.scala 160:64:@22160.4]
  wire [13:0] buffer_6_523; // @[Modules.scala 160:64:@22161.4]
  wire [14:0] _T_75441; // @[Modules.scala 160:64:@22163.4]
  wire [13:0] _T_75442; // @[Modules.scala 160:64:@22164.4]
  wire [13:0] buffer_6_524; // @[Modules.scala 160:64:@22165.4]
  wire [14:0] _T_75444; // @[Modules.scala 160:64:@22167.4]
  wire [13:0] _T_75445; // @[Modules.scala 160:64:@22168.4]
  wire [13:0] buffer_6_525; // @[Modules.scala 160:64:@22169.4]
  wire [14:0] _T_75447; // @[Modules.scala 160:64:@22171.4]
  wire [13:0] _T_75448; // @[Modules.scala 160:64:@22172.4]
  wire [13:0] buffer_6_526; // @[Modules.scala 160:64:@22173.4]
  wire [14:0] _T_75450; // @[Modules.scala 160:64:@22175.4]
  wire [13:0] _T_75451; // @[Modules.scala 160:64:@22176.4]
  wire [13:0] buffer_6_527; // @[Modules.scala 160:64:@22177.4]
  wire [14:0] _T_75453; // @[Modules.scala 160:64:@22179.4]
  wire [13:0] _T_75454; // @[Modules.scala 160:64:@22180.4]
  wire [13:0] buffer_6_528; // @[Modules.scala 160:64:@22181.4]
  wire [14:0] _T_75456; // @[Modules.scala 160:64:@22183.4]
  wire [13:0] _T_75457; // @[Modules.scala 160:64:@22184.4]
  wire [13:0] buffer_6_529; // @[Modules.scala 160:64:@22185.4]
  wire [14:0] _T_75459; // @[Modules.scala 160:64:@22187.4]
  wire [13:0] _T_75460; // @[Modules.scala 160:64:@22188.4]
  wire [13:0] buffer_6_530; // @[Modules.scala 160:64:@22189.4]
  wire [14:0] _T_75462; // @[Modules.scala 160:64:@22191.4]
  wire [13:0] _T_75463; // @[Modules.scala 160:64:@22192.4]
  wire [13:0] buffer_6_531; // @[Modules.scala 160:64:@22193.4]
  wire [14:0] _T_75465; // @[Modules.scala 160:64:@22195.4]
  wire [13:0] _T_75466; // @[Modules.scala 160:64:@22196.4]
  wire [13:0] buffer_6_532; // @[Modules.scala 160:64:@22197.4]
  wire [14:0] _T_75468; // @[Modules.scala 160:64:@22199.4]
  wire [13:0] _T_75469; // @[Modules.scala 160:64:@22200.4]
  wire [13:0] buffer_6_533; // @[Modules.scala 160:64:@22201.4]
  wire [14:0] _T_75471; // @[Modules.scala 160:64:@22203.4]
  wire [13:0] _T_75472; // @[Modules.scala 160:64:@22204.4]
  wire [13:0] buffer_6_534; // @[Modules.scala 160:64:@22205.4]
  wire [14:0] _T_75474; // @[Modules.scala 160:64:@22207.4]
  wire [13:0] _T_75475; // @[Modules.scala 160:64:@22208.4]
  wire [13:0] buffer_6_535; // @[Modules.scala 160:64:@22209.4]
  wire [14:0] _T_75477; // @[Modules.scala 160:64:@22211.4]
  wire [13:0] _T_75478; // @[Modules.scala 160:64:@22212.4]
  wire [13:0] buffer_6_536; // @[Modules.scala 160:64:@22213.4]
  wire [14:0] _T_75480; // @[Modules.scala 160:64:@22215.4]
  wire [13:0] _T_75481; // @[Modules.scala 160:64:@22216.4]
  wire [13:0] buffer_6_537; // @[Modules.scala 160:64:@22217.4]
  wire [14:0] _T_75483; // @[Modules.scala 160:64:@22219.4]
  wire [13:0] _T_75484; // @[Modules.scala 160:64:@22220.4]
  wire [13:0] buffer_6_538; // @[Modules.scala 160:64:@22221.4]
  wire [14:0] _T_75486; // @[Modules.scala 160:64:@22223.4]
  wire [13:0] _T_75487; // @[Modules.scala 160:64:@22224.4]
  wire [13:0] buffer_6_539; // @[Modules.scala 160:64:@22225.4]
  wire [14:0] _T_75489; // @[Modules.scala 160:64:@22227.4]
  wire [13:0] _T_75490; // @[Modules.scala 160:64:@22228.4]
  wire [13:0] buffer_6_540; // @[Modules.scala 160:64:@22229.4]
  wire [14:0] _T_75492; // @[Modules.scala 160:64:@22231.4]
  wire [13:0] _T_75493; // @[Modules.scala 160:64:@22232.4]
  wire [13:0] buffer_6_541; // @[Modules.scala 160:64:@22233.4]
  wire [14:0] _T_75495; // @[Modules.scala 160:64:@22235.4]
  wire [13:0] _T_75496; // @[Modules.scala 160:64:@22236.4]
  wire [13:0] buffer_6_542; // @[Modules.scala 160:64:@22237.4]
  wire [14:0] _T_75498; // @[Modules.scala 160:64:@22239.4]
  wire [13:0] _T_75499; // @[Modules.scala 160:64:@22240.4]
  wire [13:0] buffer_6_543; // @[Modules.scala 160:64:@22241.4]
  wire [14:0] _T_75501; // @[Modules.scala 160:64:@22243.4]
  wire [13:0] _T_75502; // @[Modules.scala 160:64:@22244.4]
  wire [13:0] buffer_6_544; // @[Modules.scala 160:64:@22245.4]
  wire [14:0] _T_75504; // @[Modules.scala 160:64:@22247.4]
  wire [13:0] _T_75505; // @[Modules.scala 160:64:@22248.4]
  wire [13:0] buffer_6_545; // @[Modules.scala 160:64:@22249.4]
  wire [14:0] _T_75507; // @[Modules.scala 160:64:@22251.4]
  wire [13:0] _T_75508; // @[Modules.scala 160:64:@22252.4]
  wire [13:0] buffer_6_546; // @[Modules.scala 160:64:@22253.4]
  wire [14:0] _T_75510; // @[Modules.scala 160:64:@22255.4]
  wire [13:0] _T_75511; // @[Modules.scala 160:64:@22256.4]
  wire [13:0] buffer_6_547; // @[Modules.scala 160:64:@22257.4]
  wire [14:0] _T_75513; // @[Modules.scala 160:64:@22259.4]
  wire [13:0] _T_75514; // @[Modules.scala 160:64:@22260.4]
  wire [13:0] buffer_6_548; // @[Modules.scala 160:64:@22261.4]
  wire [14:0] _T_75516; // @[Modules.scala 160:64:@22263.4]
  wire [13:0] _T_75517; // @[Modules.scala 160:64:@22264.4]
  wire [13:0] buffer_6_549; // @[Modules.scala 160:64:@22265.4]
  wire [14:0] _T_75519; // @[Modules.scala 160:64:@22267.4]
  wire [13:0] _T_75520; // @[Modules.scala 160:64:@22268.4]
  wire [13:0] buffer_6_550; // @[Modules.scala 160:64:@22269.4]
  wire [14:0] _T_75522; // @[Modules.scala 160:64:@22271.4]
  wire [13:0] _T_75523; // @[Modules.scala 160:64:@22272.4]
  wire [13:0] buffer_6_551; // @[Modules.scala 160:64:@22273.4]
  wire [14:0] _T_75525; // @[Modules.scala 160:64:@22275.4]
  wire [13:0] _T_75526; // @[Modules.scala 160:64:@22276.4]
  wire [13:0] buffer_6_552; // @[Modules.scala 160:64:@22277.4]
  wire [14:0] _T_75528; // @[Modules.scala 166:64:@22279.4]
  wire [13:0] _T_75529; // @[Modules.scala 166:64:@22280.4]
  wire [13:0] buffer_6_553; // @[Modules.scala 166:64:@22281.4]
  wire [14:0] _T_75531; // @[Modules.scala 166:64:@22283.4]
  wire [13:0] _T_75532; // @[Modules.scala 166:64:@22284.4]
  wire [13:0] buffer_6_554; // @[Modules.scala 166:64:@22285.4]
  wire [14:0] _T_75534; // @[Modules.scala 166:64:@22287.4]
  wire [13:0] _T_75535; // @[Modules.scala 166:64:@22288.4]
  wire [13:0] buffer_6_555; // @[Modules.scala 166:64:@22289.4]
  wire [14:0] _T_75537; // @[Modules.scala 166:64:@22291.4]
  wire [13:0] _T_75538; // @[Modules.scala 166:64:@22292.4]
  wire [13:0] buffer_6_556; // @[Modules.scala 166:64:@22293.4]
  wire [14:0] _T_75540; // @[Modules.scala 166:64:@22295.4]
  wire [13:0] _T_75541; // @[Modules.scala 166:64:@22296.4]
  wire [13:0] buffer_6_557; // @[Modules.scala 166:64:@22297.4]
  wire [14:0] _T_75543; // @[Modules.scala 166:64:@22299.4]
  wire [13:0] _T_75544; // @[Modules.scala 166:64:@22300.4]
  wire [13:0] buffer_6_558; // @[Modules.scala 166:64:@22301.4]
  wire [14:0] _T_75546; // @[Modules.scala 166:64:@22303.4]
  wire [13:0] _T_75547; // @[Modules.scala 166:64:@22304.4]
  wire [13:0] buffer_6_559; // @[Modules.scala 166:64:@22305.4]
  wire [14:0] _T_75549; // @[Modules.scala 166:64:@22307.4]
  wire [13:0] _T_75550; // @[Modules.scala 166:64:@22308.4]
  wire [13:0] buffer_6_560; // @[Modules.scala 166:64:@22309.4]
  wire [14:0] _T_75552; // @[Modules.scala 166:64:@22311.4]
  wire [13:0] _T_75553; // @[Modules.scala 166:64:@22312.4]
  wire [13:0] buffer_6_561; // @[Modules.scala 166:64:@22313.4]
  wire [14:0] _T_75555; // @[Modules.scala 166:64:@22315.4]
  wire [13:0] _T_75556; // @[Modules.scala 166:64:@22316.4]
  wire [13:0] buffer_6_562; // @[Modules.scala 166:64:@22317.4]
  wire [14:0] _T_75558; // @[Modules.scala 166:64:@22319.4]
  wire [13:0] _T_75559; // @[Modules.scala 166:64:@22320.4]
  wire [13:0] buffer_6_563; // @[Modules.scala 166:64:@22321.4]
  wire [14:0] _T_75561; // @[Modules.scala 166:64:@22323.4]
  wire [13:0] _T_75562; // @[Modules.scala 166:64:@22324.4]
  wire [13:0] buffer_6_564; // @[Modules.scala 166:64:@22325.4]
  wire [14:0] _T_75564; // @[Modules.scala 166:64:@22327.4]
  wire [13:0] _T_75565; // @[Modules.scala 166:64:@22328.4]
  wire [13:0] buffer_6_565; // @[Modules.scala 166:64:@22329.4]
  wire [14:0] _T_75567; // @[Modules.scala 166:64:@22331.4]
  wire [13:0] _T_75568; // @[Modules.scala 166:64:@22332.4]
  wire [13:0] buffer_6_566; // @[Modules.scala 166:64:@22333.4]
  wire [14:0] _T_75570; // @[Modules.scala 166:64:@22335.4]
  wire [13:0] _T_75571; // @[Modules.scala 166:64:@22336.4]
  wire [13:0] buffer_6_567; // @[Modules.scala 166:64:@22337.4]
  wire [14:0] _T_75573; // @[Modules.scala 166:64:@22339.4]
  wire [13:0] _T_75574; // @[Modules.scala 166:64:@22340.4]
  wire [13:0] buffer_6_568; // @[Modules.scala 166:64:@22341.4]
  wire [14:0] _T_75576; // @[Modules.scala 166:64:@22343.4]
  wire [13:0] _T_75577; // @[Modules.scala 166:64:@22344.4]
  wire [13:0] buffer_6_569; // @[Modules.scala 166:64:@22345.4]
  wire [14:0] _T_75579; // @[Modules.scala 166:64:@22347.4]
  wire [13:0] _T_75580; // @[Modules.scala 166:64:@22348.4]
  wire [13:0] buffer_6_570; // @[Modules.scala 166:64:@22349.4]
  wire [14:0] _T_75582; // @[Modules.scala 166:64:@22351.4]
  wire [13:0] _T_75583; // @[Modules.scala 166:64:@22352.4]
  wire [13:0] buffer_6_571; // @[Modules.scala 166:64:@22353.4]
  wire [14:0] _T_75585; // @[Modules.scala 166:64:@22355.4]
  wire [13:0] _T_75586; // @[Modules.scala 166:64:@22356.4]
  wire [13:0] buffer_6_572; // @[Modules.scala 166:64:@22357.4]
  wire [14:0] _T_75588; // @[Modules.scala 166:64:@22359.4]
  wire [13:0] _T_75589; // @[Modules.scala 166:64:@22360.4]
  wire [13:0] buffer_6_573; // @[Modules.scala 166:64:@22361.4]
  wire [14:0] _T_75591; // @[Modules.scala 166:64:@22363.4]
  wire [13:0] _T_75592; // @[Modules.scala 166:64:@22364.4]
  wire [13:0] buffer_6_574; // @[Modules.scala 166:64:@22365.4]
  wire [14:0] _T_75594; // @[Modules.scala 166:64:@22367.4]
  wire [13:0] _T_75595; // @[Modules.scala 166:64:@22368.4]
  wire [13:0] buffer_6_575; // @[Modules.scala 166:64:@22369.4]
  wire [14:0] _T_75597; // @[Modules.scala 166:64:@22371.4]
  wire [13:0] _T_75598; // @[Modules.scala 166:64:@22372.4]
  wire [13:0] buffer_6_576; // @[Modules.scala 166:64:@22373.4]
  wire [14:0] _T_75600; // @[Modules.scala 166:64:@22375.4]
  wire [13:0] _T_75601; // @[Modules.scala 166:64:@22376.4]
  wire [13:0] buffer_6_577; // @[Modules.scala 166:64:@22377.4]
  wire [14:0] _T_75603; // @[Modules.scala 166:64:@22379.4]
  wire [13:0] _T_75604; // @[Modules.scala 166:64:@22380.4]
  wire [13:0] buffer_6_578; // @[Modules.scala 166:64:@22381.4]
  wire [14:0] _T_75606; // @[Modules.scala 166:64:@22383.4]
  wire [13:0] _T_75607; // @[Modules.scala 166:64:@22384.4]
  wire [13:0] buffer_6_579; // @[Modules.scala 166:64:@22385.4]
  wire [14:0] _T_75609; // @[Modules.scala 166:64:@22387.4]
  wire [13:0] _T_75610; // @[Modules.scala 166:64:@22388.4]
  wire [13:0] buffer_6_580; // @[Modules.scala 166:64:@22389.4]
  wire [14:0] _T_75612; // @[Modules.scala 166:64:@22391.4]
  wire [13:0] _T_75613; // @[Modules.scala 166:64:@22392.4]
  wire [13:0] buffer_6_581; // @[Modules.scala 166:64:@22393.4]
  wire [14:0] _T_75615; // @[Modules.scala 166:64:@22395.4]
  wire [13:0] _T_75616; // @[Modules.scala 166:64:@22396.4]
  wire [13:0] buffer_6_582; // @[Modules.scala 166:64:@22397.4]
  wire [14:0] _T_75618; // @[Modules.scala 166:64:@22399.4]
  wire [13:0] _T_75619; // @[Modules.scala 166:64:@22400.4]
  wire [13:0] buffer_6_583; // @[Modules.scala 166:64:@22401.4]
  wire [14:0] _T_75621; // @[Modules.scala 166:64:@22403.4]
  wire [13:0] _T_75622; // @[Modules.scala 166:64:@22404.4]
  wire [13:0] buffer_6_584; // @[Modules.scala 166:64:@22405.4]
  wire [14:0] _T_75624; // @[Modules.scala 166:64:@22407.4]
  wire [13:0] _T_75625; // @[Modules.scala 166:64:@22408.4]
  wire [13:0] buffer_6_585; // @[Modules.scala 166:64:@22409.4]
  wire [14:0] _T_75627; // @[Modules.scala 166:64:@22411.4]
  wire [13:0] _T_75628; // @[Modules.scala 166:64:@22412.4]
  wire [13:0] buffer_6_586; // @[Modules.scala 166:64:@22413.4]
  wire [14:0] _T_75630; // @[Modules.scala 166:64:@22415.4]
  wire [13:0] _T_75631; // @[Modules.scala 166:64:@22416.4]
  wire [13:0] buffer_6_587; // @[Modules.scala 166:64:@22417.4]
  wire [14:0] _T_75633; // @[Modules.scala 166:64:@22419.4]
  wire [13:0] _T_75634; // @[Modules.scala 166:64:@22420.4]
  wire [13:0] buffer_6_588; // @[Modules.scala 166:64:@22421.4]
  wire [14:0] _T_75636; // @[Modules.scala 166:64:@22423.4]
  wire [13:0] _T_75637; // @[Modules.scala 166:64:@22424.4]
  wire [13:0] buffer_6_589; // @[Modules.scala 166:64:@22425.4]
  wire [14:0] _T_75639; // @[Modules.scala 166:64:@22427.4]
  wire [13:0] _T_75640; // @[Modules.scala 166:64:@22428.4]
  wire [13:0] buffer_6_590; // @[Modules.scala 166:64:@22429.4]
  wire [14:0] _T_75642; // @[Modules.scala 166:64:@22431.4]
  wire [13:0] _T_75643; // @[Modules.scala 166:64:@22432.4]
  wire [13:0] buffer_6_591; // @[Modules.scala 166:64:@22433.4]
  wire [14:0] _T_75645; // @[Modules.scala 166:64:@22435.4]
  wire [13:0] _T_75646; // @[Modules.scala 166:64:@22436.4]
  wire [13:0] buffer_6_592; // @[Modules.scala 166:64:@22437.4]
  wire [14:0] _T_75648; // @[Modules.scala 166:64:@22439.4]
  wire [13:0] _T_75649; // @[Modules.scala 166:64:@22440.4]
  wire [13:0] buffer_6_593; // @[Modules.scala 166:64:@22441.4]
  wire [14:0] _T_75651; // @[Modules.scala 166:64:@22443.4]
  wire [13:0] _T_75652; // @[Modules.scala 166:64:@22444.4]
  wire [13:0] buffer_6_594; // @[Modules.scala 166:64:@22445.4]
  wire [14:0] _T_75654; // @[Modules.scala 166:64:@22447.4]
  wire [13:0] _T_75655; // @[Modules.scala 166:64:@22448.4]
  wire [13:0] buffer_6_595; // @[Modules.scala 166:64:@22449.4]
  wire [14:0] _T_75657; // @[Modules.scala 166:64:@22451.4]
  wire [13:0] _T_75658; // @[Modules.scala 166:64:@22452.4]
  wire [13:0] buffer_6_596; // @[Modules.scala 166:64:@22453.4]
  wire [14:0] _T_75660; // @[Modules.scala 166:64:@22455.4]
  wire [13:0] _T_75661; // @[Modules.scala 166:64:@22456.4]
  wire [13:0] buffer_6_597; // @[Modules.scala 166:64:@22457.4]
  wire [14:0] _T_75663; // @[Modules.scala 166:64:@22459.4]
  wire [13:0] _T_75664; // @[Modules.scala 166:64:@22460.4]
  wire [13:0] buffer_6_598; // @[Modules.scala 166:64:@22461.4]
  wire [14:0] _T_75666; // @[Modules.scala 166:64:@22463.4]
  wire [13:0] _T_75667; // @[Modules.scala 166:64:@22464.4]
  wire [13:0] buffer_6_599; // @[Modules.scala 166:64:@22465.4]
  wire [14:0] _T_75669; // @[Modules.scala 166:64:@22467.4]
  wire [13:0] _T_75670; // @[Modules.scala 166:64:@22468.4]
  wire [13:0] buffer_6_600; // @[Modules.scala 166:64:@22469.4]
  wire [14:0] _T_75672; // @[Modules.scala 166:64:@22471.4]
  wire [13:0] _T_75673; // @[Modules.scala 166:64:@22472.4]
  wire [13:0] buffer_6_601; // @[Modules.scala 166:64:@22473.4]
  wire [14:0] _T_75675; // @[Modules.scala 166:64:@22475.4]
  wire [13:0] _T_75676; // @[Modules.scala 166:64:@22476.4]
  wire [13:0] buffer_6_602; // @[Modules.scala 166:64:@22477.4]
  wire [14:0] _T_75678; // @[Modules.scala 166:64:@22479.4]
  wire [13:0] _T_75679; // @[Modules.scala 166:64:@22480.4]
  wire [13:0] buffer_6_603; // @[Modules.scala 166:64:@22481.4]
  wire [14:0] _T_75681; // @[Modules.scala 166:64:@22483.4]
  wire [13:0] _T_75682; // @[Modules.scala 166:64:@22484.4]
  wire [13:0] buffer_6_604; // @[Modules.scala 166:64:@22485.4]
  wire [14:0] _T_75684; // @[Modules.scala 166:64:@22487.4]
  wire [13:0] _T_75685; // @[Modules.scala 166:64:@22488.4]
  wire [13:0] buffer_6_605; // @[Modules.scala 166:64:@22489.4]
  wire [14:0] _T_75687; // @[Modules.scala 166:64:@22491.4]
  wire [13:0] _T_75688; // @[Modules.scala 166:64:@22492.4]
  wire [13:0] buffer_6_606; // @[Modules.scala 166:64:@22493.4]
  wire [14:0] _T_75690; // @[Modules.scala 166:64:@22495.4]
  wire [13:0] _T_75691; // @[Modules.scala 166:64:@22496.4]
  wire [13:0] buffer_6_607; // @[Modules.scala 166:64:@22497.4]
  wire [14:0] _T_75693; // @[Modules.scala 166:64:@22499.4]
  wire [13:0] _T_75694; // @[Modules.scala 166:64:@22500.4]
  wire [13:0] buffer_6_608; // @[Modules.scala 166:64:@22501.4]
  wire [14:0] _T_75696; // @[Modules.scala 166:64:@22503.4]
  wire [13:0] _T_75697; // @[Modules.scala 166:64:@22504.4]
  wire [13:0] buffer_6_609; // @[Modules.scala 166:64:@22505.4]
  wire [14:0] _T_75699; // @[Modules.scala 166:64:@22507.4]
  wire [13:0] _T_75700; // @[Modules.scala 166:64:@22508.4]
  wire [13:0] buffer_6_610; // @[Modules.scala 166:64:@22509.4]
  wire [14:0] _T_75702; // @[Modules.scala 172:66:@22511.4]
  wire [13:0] _T_75703; // @[Modules.scala 172:66:@22512.4]
  wire [13:0] buffer_6_611; // @[Modules.scala 172:66:@22513.4]
  wire [14:0] _T_75705; // @[Modules.scala 160:64:@22515.4]
  wire [13:0] _T_75706; // @[Modules.scala 160:64:@22516.4]
  wire [13:0] buffer_6_612; // @[Modules.scala 160:64:@22517.4]
  wire [14:0] _T_75708; // @[Modules.scala 160:64:@22519.4]
  wire [13:0] _T_75709; // @[Modules.scala 160:64:@22520.4]
  wire [13:0] buffer_6_613; // @[Modules.scala 160:64:@22521.4]
  wire [14:0] _T_75711; // @[Modules.scala 160:64:@22523.4]
  wire [13:0] _T_75712; // @[Modules.scala 160:64:@22524.4]
  wire [13:0] buffer_6_614; // @[Modules.scala 160:64:@22525.4]
  wire [14:0] _T_75714; // @[Modules.scala 160:64:@22527.4]
  wire [13:0] _T_75715; // @[Modules.scala 160:64:@22528.4]
  wire [13:0] buffer_6_615; // @[Modules.scala 160:64:@22529.4]
  wire [14:0] _T_75717; // @[Modules.scala 160:64:@22531.4]
  wire [13:0] _T_75718; // @[Modules.scala 160:64:@22532.4]
  wire [13:0] buffer_6_616; // @[Modules.scala 160:64:@22533.4]
  wire [14:0] _T_75720; // @[Modules.scala 160:64:@22535.4]
  wire [13:0] _T_75721; // @[Modules.scala 160:64:@22536.4]
  wire [13:0] buffer_6_617; // @[Modules.scala 160:64:@22537.4]
  wire [14:0] _T_75723; // @[Modules.scala 160:64:@22539.4]
  wire [13:0] _T_75724; // @[Modules.scala 160:64:@22540.4]
  wire [13:0] buffer_6_618; // @[Modules.scala 160:64:@22541.4]
  wire [14:0] _T_75726; // @[Modules.scala 160:64:@22543.4]
  wire [13:0] _T_75727; // @[Modules.scala 160:64:@22544.4]
  wire [13:0] buffer_6_619; // @[Modules.scala 160:64:@22545.4]
  wire [14:0] _T_75729; // @[Modules.scala 160:64:@22547.4]
  wire [13:0] _T_75730; // @[Modules.scala 160:64:@22548.4]
  wire [13:0] buffer_6_620; // @[Modules.scala 160:64:@22549.4]
  wire [14:0] _T_75732; // @[Modules.scala 160:64:@22551.4]
  wire [13:0] _T_75733; // @[Modules.scala 160:64:@22552.4]
  wire [13:0] buffer_6_621; // @[Modules.scala 160:64:@22553.4]
  wire [14:0] _T_75735; // @[Modules.scala 160:64:@22555.4]
  wire [13:0] _T_75736; // @[Modules.scala 160:64:@22556.4]
  wire [13:0] buffer_6_622; // @[Modules.scala 160:64:@22557.4]
  wire [14:0] _T_75738; // @[Modules.scala 160:64:@22559.4]
  wire [13:0] _T_75739; // @[Modules.scala 160:64:@22560.4]
  wire [13:0] buffer_6_623; // @[Modules.scala 160:64:@22561.4]
  wire [14:0] _T_75741; // @[Modules.scala 160:64:@22563.4]
  wire [13:0] _T_75742; // @[Modules.scala 160:64:@22564.4]
  wire [13:0] buffer_6_624; // @[Modules.scala 160:64:@22565.4]
  wire [14:0] _T_75744; // @[Modules.scala 160:64:@22567.4]
  wire [13:0] _T_75745; // @[Modules.scala 160:64:@22568.4]
  wire [13:0] buffer_6_625; // @[Modules.scala 160:64:@22569.4]
  wire [14:0] _T_75747; // @[Modules.scala 160:64:@22571.4]
  wire [13:0] _T_75748; // @[Modules.scala 160:64:@22572.4]
  wire [13:0] buffer_6_626; // @[Modules.scala 160:64:@22573.4]
  wire [14:0] _T_75750; // @[Modules.scala 166:64:@22575.4]
  wire [13:0] _T_75751; // @[Modules.scala 166:64:@22576.4]
  wire [13:0] buffer_6_627; // @[Modules.scala 166:64:@22577.4]
  wire [14:0] _T_75753; // @[Modules.scala 166:64:@22579.4]
  wire [13:0] _T_75754; // @[Modules.scala 166:64:@22580.4]
  wire [13:0] buffer_6_628; // @[Modules.scala 166:64:@22581.4]
  wire [14:0] _T_75756; // @[Modules.scala 160:64:@22583.4]
  wire [13:0] _T_75757; // @[Modules.scala 160:64:@22584.4]
  wire [13:0] buffer_6_629; // @[Modules.scala 160:64:@22585.4]
  wire [14:0] _T_75759; // @[Modules.scala 172:66:@22587.4]
  wire [13:0] _T_75760; // @[Modules.scala 172:66:@22588.4]
  wire [13:0] buffer_6_630; // @[Modules.scala 172:66:@22589.4]
  wire [4:0] _T_75763; // @[Modules.scala 143:74:@22744.4]
  wire [5:0] _T_75766; // @[Modules.scala 143:103:@22746.4]
  wire [4:0] _T_75767; // @[Modules.scala 143:103:@22747.4]
  wire [4:0] _T_75768; // @[Modules.scala 143:103:@22748.4]
  wire [5:0] _GEN_498; // @[Modules.scala 143:103:@22770.4]
  wire [6:0] _T_75794; // @[Modules.scala 143:103:@22770.4]
  wire [5:0] _T_75795; // @[Modules.scala 143:103:@22771.4]
  wire [5:0] _T_75796; // @[Modules.scala 143:103:@22772.4]
  wire [5:0] _T_75829; // @[Modules.scala 143:103:@22800.4]
  wire [4:0] _T_75830; // @[Modules.scala 143:103:@22801.4]
  wire [4:0] _T_75831; // @[Modules.scala 143:103:@22802.4]
  wire [6:0] _T_75857; // @[Modules.scala 143:103:@22824.4]
  wire [5:0] _T_75858; // @[Modules.scala 143:103:@22825.4]
  wire [5:0] _T_75859; // @[Modules.scala 143:103:@22826.4]
  wire [6:0] _T_75906; // @[Modules.scala 143:103:@22866.4]
  wire [5:0] _T_75907; // @[Modules.scala 143:103:@22867.4]
  wire [5:0] _T_75908; // @[Modules.scala 143:103:@22868.4]
  wire [6:0] _T_75920; // @[Modules.scala 143:103:@22878.4]
  wire [5:0] _T_75921; // @[Modules.scala 143:103:@22879.4]
  wire [5:0] _T_75922; // @[Modules.scala 143:103:@22880.4]
  wire [5:0] _GEN_502; // @[Modules.scala 143:103:@22890.4]
  wire [6:0] _T_75934; // @[Modules.scala 143:103:@22890.4]
  wire [5:0] _T_75935; // @[Modules.scala 143:103:@22891.4]
  wire [5:0] _T_75936; // @[Modules.scala 143:103:@22892.4]
  wire [5:0] _GEN_503; // @[Modules.scala 143:103:@22944.4]
  wire [6:0] _T_75997; // @[Modules.scala 143:103:@22944.4]
  wire [5:0] _T_75998; // @[Modules.scala 143:103:@22945.4]
  wire [5:0] _T_75999; // @[Modules.scala 143:103:@22946.4]
  wire [5:0] _GEN_505; // @[Modules.scala 143:103:@22956.4]
  wire [6:0] _T_76011; // @[Modules.scala 143:103:@22956.4]
  wire [5:0] _T_76012; // @[Modules.scala 143:103:@22957.4]
  wire [5:0] _T_76013; // @[Modules.scala 143:103:@22958.4]
  wire [5:0] _GEN_506; // @[Modules.scala 143:103:@22974.4]
  wire [6:0] _T_76032; // @[Modules.scala 143:103:@22974.4]
  wire [5:0] _T_76033; // @[Modules.scala 143:103:@22975.4]
  wire [5:0] _T_76034; // @[Modules.scala 143:103:@22976.4]
  wire [5:0] _T_76046; // @[Modules.scala 143:103:@22986.4]
  wire [4:0] _T_76047; // @[Modules.scala 143:103:@22987.4]
  wire [4:0] _T_76048; // @[Modules.scala 143:103:@22988.4]
  wire [4:0] _T_76052; // @[Modules.scala 144:80:@22991.4]
  wire [5:0] _T_76053; // @[Modules.scala 143:103:@22992.4]
  wire [4:0] _T_76054; // @[Modules.scala 143:103:@22993.4]
  wire [4:0] _T_76055; // @[Modules.scala 143:103:@22994.4]
  wire [4:0] _T_76057; // @[Modules.scala 143:74:@22996.4]
  wire [5:0] _T_76060; // @[Modules.scala 143:103:@22998.4]
  wire [4:0] _T_76061; // @[Modules.scala 143:103:@22999.4]
  wire [4:0] _T_76062; // @[Modules.scala 143:103:@23000.4]
  wire [5:0] _GEN_507; // @[Modules.scala 143:103:@23004.4]
  wire [6:0] _T_76067; // @[Modules.scala 143:103:@23004.4]
  wire [5:0] _T_76068; // @[Modules.scala 143:103:@23005.4]
  wire [5:0] _T_76069; // @[Modules.scala 143:103:@23006.4]
  wire [6:0] _T_76081; // @[Modules.scala 143:103:@23016.4]
  wire [5:0] _T_76082; // @[Modules.scala 143:103:@23017.4]
  wire [5:0] _T_76083; // @[Modules.scala 143:103:@23018.4]
  wire [5:0] _GEN_509; // @[Modules.scala 143:103:@23040.4]
  wire [6:0] _T_76109; // @[Modules.scala 143:103:@23040.4]
  wire [5:0] _T_76110; // @[Modules.scala 143:103:@23041.4]
  wire [5:0] _T_76111; // @[Modules.scala 143:103:@23042.4]
  wire [5:0] _T_76122; // @[Modules.scala 144:80:@23051.4]
  wire [6:0] _T_76123; // @[Modules.scala 143:103:@23052.4]
  wire [5:0] _T_76124; // @[Modules.scala 143:103:@23053.4]
  wire [5:0] _T_76125; // @[Modules.scala 143:103:@23054.4]
  wire [6:0] _T_76130; // @[Modules.scala 143:103:@23058.4]
  wire [5:0] _T_76131; // @[Modules.scala 143:103:@23059.4]
  wire [5:0] _T_76132; // @[Modules.scala 143:103:@23060.4]
  wire [6:0] _T_76137; // @[Modules.scala 143:103:@23064.4]
  wire [5:0] _T_76138; // @[Modules.scala 143:103:@23065.4]
  wire [5:0] _T_76139; // @[Modules.scala 143:103:@23066.4]
  wire [6:0] _T_76144; // @[Modules.scala 143:103:@23070.4]
  wire [5:0] _T_76145; // @[Modules.scala 143:103:@23071.4]
  wire [5:0] _T_76146; // @[Modules.scala 143:103:@23072.4]
  wire [5:0] _T_76150; // @[Modules.scala 144:80:@23075.4]
  wire [6:0] _T_76151; // @[Modules.scala 143:103:@23076.4]
  wire [5:0] _T_76152; // @[Modules.scala 143:103:@23077.4]
  wire [5:0] _T_76153; // @[Modules.scala 143:103:@23078.4]
  wire [6:0] _T_76165; // @[Modules.scala 143:103:@23088.4]
  wire [5:0] _T_76166; // @[Modules.scala 143:103:@23089.4]
  wire [5:0] _T_76167; // @[Modules.scala 143:103:@23090.4]
  wire [5:0] _T_76186; // @[Modules.scala 143:103:@23106.4]
  wire [4:0] _T_76187; // @[Modules.scala 143:103:@23107.4]
  wire [4:0] _T_76188; // @[Modules.scala 143:103:@23108.4]
  wire [5:0] _GEN_513; // @[Modules.scala 143:103:@23124.4]
  wire [6:0] _T_76207; // @[Modules.scala 143:103:@23124.4]
  wire [5:0] _T_76208; // @[Modules.scala 143:103:@23125.4]
  wire [5:0] _T_76209; // @[Modules.scala 143:103:@23126.4]
  wire [6:0] _T_76228; // @[Modules.scala 143:103:@23142.4]
  wire [5:0] _T_76229; // @[Modules.scala 143:103:@23143.4]
  wire [5:0] _T_76230; // @[Modules.scala 143:103:@23144.4]
  wire [6:0] _T_76242; // @[Modules.scala 143:103:@23154.4]
  wire [5:0] _T_76243; // @[Modules.scala 143:103:@23155.4]
  wire [5:0] _T_76244; // @[Modules.scala 143:103:@23156.4]
  wire [6:0] _T_76284; // @[Modules.scala 143:103:@23190.4]
  wire [5:0] _T_76285; // @[Modules.scala 143:103:@23191.4]
  wire [5:0] _T_76286; // @[Modules.scala 143:103:@23192.4]
  wire [6:0] _T_76291; // @[Modules.scala 143:103:@23196.4]
  wire [5:0] _T_76292; // @[Modules.scala 143:103:@23197.4]
  wire [5:0] _T_76293; // @[Modules.scala 143:103:@23198.4]
  wire [6:0] _T_76298; // @[Modules.scala 143:103:@23202.4]
  wire [5:0] _T_76299; // @[Modules.scala 143:103:@23203.4]
  wire [5:0] _T_76300; // @[Modules.scala 143:103:@23204.4]
  wire [6:0] _T_76305; // @[Modules.scala 143:103:@23208.4]
  wire [5:0] _T_76306; // @[Modules.scala 143:103:@23209.4]
  wire [5:0] _T_76307; // @[Modules.scala 143:103:@23210.4]
  wire [6:0] _T_76340; // @[Modules.scala 143:103:@23238.4]
  wire [5:0] _T_76341; // @[Modules.scala 143:103:@23239.4]
  wire [5:0] _T_76342; // @[Modules.scala 143:103:@23240.4]
  wire [6:0] _T_76347; // @[Modules.scala 143:103:@23244.4]
  wire [5:0] _T_76348; // @[Modules.scala 143:103:@23245.4]
  wire [5:0] _T_76349; // @[Modules.scala 143:103:@23246.4]
  wire [5:0] _GEN_516; // @[Modules.scala 143:103:@23250.4]
  wire [6:0] _T_76354; // @[Modules.scala 143:103:@23250.4]
  wire [5:0] _T_76355; // @[Modules.scala 143:103:@23251.4]
  wire [5:0] _T_76356; // @[Modules.scala 143:103:@23252.4]
  wire [6:0] _T_76368; // @[Modules.scala 143:103:@23262.4]
  wire [5:0] _T_76369; // @[Modules.scala 143:103:@23263.4]
  wire [5:0] _T_76370; // @[Modules.scala 143:103:@23264.4]
  wire [6:0] _T_76466; // @[Modules.scala 143:103:@23346.4]
  wire [5:0] _T_76467; // @[Modules.scala 143:103:@23347.4]
  wire [5:0] _T_76468; // @[Modules.scala 143:103:@23348.4]
  wire [5:0] _GEN_518; // @[Modules.scala 143:103:@23418.4]
  wire [6:0] _T_76550; // @[Modules.scala 143:103:@23418.4]
  wire [5:0] _T_76551; // @[Modules.scala 143:103:@23419.4]
  wire [5:0] _T_76552; // @[Modules.scala 143:103:@23420.4]
  wire [5:0] _GEN_519; // @[Modules.scala 143:103:@23436.4]
  wire [6:0] _T_76571; // @[Modules.scala 143:103:@23436.4]
  wire [5:0] _T_76572; // @[Modules.scala 143:103:@23437.4]
  wire [5:0] _T_76573; // @[Modules.scala 143:103:@23438.4]
  wire [6:0] _T_76606; // @[Modules.scala 143:103:@23466.4]
  wire [5:0] _T_76607; // @[Modules.scala 143:103:@23467.4]
  wire [5:0] _T_76608; // @[Modules.scala 143:103:@23468.4]
  wire [5:0] _GEN_521; // @[Modules.scala 143:103:@23496.4]
  wire [6:0] _T_76641; // @[Modules.scala 143:103:@23496.4]
  wire [5:0] _T_76642; // @[Modules.scala 143:103:@23497.4]
  wire [5:0] _T_76643; // @[Modules.scala 143:103:@23498.4]
  wire [6:0] _T_76648; // @[Modules.scala 143:103:@23502.4]
  wire [5:0] _T_76649; // @[Modules.scala 143:103:@23503.4]
  wire [5:0] _T_76650; // @[Modules.scala 143:103:@23504.4]
  wire [5:0] _GEN_523; // @[Modules.scala 143:103:@23520.4]
  wire [6:0] _T_76669; // @[Modules.scala 143:103:@23520.4]
  wire [5:0] _T_76670; // @[Modules.scala 143:103:@23521.4]
  wire [5:0] _T_76671; // @[Modules.scala 143:103:@23522.4]
  wire [4:0] _T_76696; // @[Modules.scala 144:80:@23543.4]
  wire [5:0] _T_76697; // @[Modules.scala 143:103:@23544.4]
  wire [4:0] _T_76698; // @[Modules.scala 143:103:@23545.4]
  wire [4:0] _T_76699; // @[Modules.scala 143:103:@23546.4]
  wire [4:0] _T_76778; // @[Modules.scala 143:74:@23614.4]
  wire [5:0] _T_76781; // @[Modules.scala 143:103:@23616.4]
  wire [4:0] _T_76782; // @[Modules.scala 143:103:@23617.4]
  wire [4:0] _T_76783; // @[Modules.scala 143:103:@23618.4]
  wire [4:0] _T_76787; // @[Modules.scala 144:80:@23621.4]
  wire [5:0] _T_76788; // @[Modules.scala 143:103:@23622.4]
  wire [4:0] _T_76789; // @[Modules.scala 143:103:@23623.4]
  wire [4:0] _T_76790; // @[Modules.scala 143:103:@23624.4]
  wire [6:0] _T_76809; // @[Modules.scala 143:103:@23640.4]
  wire [5:0] _T_76810; // @[Modules.scala 143:103:@23641.4]
  wire [5:0] _T_76811; // @[Modules.scala 143:103:@23642.4]
  wire [6:0] _T_76816; // @[Modules.scala 143:103:@23646.4]
  wire [5:0] _T_76817; // @[Modules.scala 143:103:@23647.4]
  wire [5:0] _T_76818; // @[Modules.scala 143:103:@23648.4]
  wire [6:0] _T_76823; // @[Modules.scala 143:103:@23652.4]
  wire [5:0] _T_76824; // @[Modules.scala 143:103:@23653.4]
  wire [5:0] _T_76825; // @[Modules.scala 143:103:@23654.4]
  wire [5:0] _GEN_528; // @[Modules.scala 143:103:@23658.4]
  wire [6:0] _T_76830; // @[Modules.scala 143:103:@23658.4]
  wire [5:0] _T_76831; // @[Modules.scala 143:103:@23659.4]
  wire [5:0] _T_76832; // @[Modules.scala 143:103:@23660.4]
  wire [5:0] _GEN_529; // @[Modules.scala 143:103:@23688.4]
  wire [6:0] _T_76865; // @[Modules.scala 143:103:@23688.4]
  wire [5:0] _T_76866; // @[Modules.scala 143:103:@23689.4]
  wire [5:0] _T_76867; // @[Modules.scala 143:103:@23690.4]
  wire [5:0] _T_76872; // @[Modules.scala 143:103:@23694.4]
  wire [4:0] _T_76873; // @[Modules.scala 143:103:@23695.4]
  wire [4:0] _T_76874; // @[Modules.scala 143:103:@23696.4]
  wire [5:0] _T_76879; // @[Modules.scala 143:103:@23700.4]
  wire [4:0] _T_76880; // @[Modules.scala 143:103:@23701.4]
  wire [4:0] _T_76881; // @[Modules.scala 143:103:@23702.4]
  wire [5:0] _T_76900; // @[Modules.scala 143:103:@23718.4]
  wire [4:0] _T_76901; // @[Modules.scala 143:103:@23719.4]
  wire [4:0] _T_76902; // @[Modules.scala 143:103:@23720.4]
  wire [5:0] _T_76914; // @[Modules.scala 143:103:@23730.4]
  wire [4:0] _T_76915; // @[Modules.scala 143:103:@23731.4]
  wire [4:0] _T_76916; // @[Modules.scala 143:103:@23732.4]
  wire [5:0] _T_76921; // @[Modules.scala 143:103:@23736.4]
  wire [4:0] _T_76922; // @[Modules.scala 143:103:@23737.4]
  wire [4:0] _T_76923; // @[Modules.scala 143:103:@23738.4]
  wire [5:0] _T_76942; // @[Modules.scala 143:103:@23754.4]
  wire [4:0] _T_76943; // @[Modules.scala 143:103:@23755.4]
  wire [4:0] _T_76944; // @[Modules.scala 143:103:@23756.4]
  wire [5:0] _T_76963; // @[Modules.scala 143:103:@23772.4]
  wire [4:0] _T_76964; // @[Modules.scala 143:103:@23773.4]
  wire [4:0] _T_76965; // @[Modules.scala 143:103:@23774.4]
  wire [6:0] _T_76998; // @[Modules.scala 143:103:@23802.4]
  wire [5:0] _T_76999; // @[Modules.scala 143:103:@23803.4]
  wire [5:0] _T_77000; // @[Modules.scala 143:103:@23804.4]
  wire [6:0] _T_77005; // @[Modules.scala 143:103:@23808.4]
  wire [5:0] _T_77006; // @[Modules.scala 143:103:@23809.4]
  wire [5:0] _T_77007; // @[Modules.scala 143:103:@23810.4]
  wire [5:0] _GEN_533; // @[Modules.scala 143:103:@23880.4]
  wire [6:0] _T_77089; // @[Modules.scala 143:103:@23880.4]
  wire [5:0] _T_77090; // @[Modules.scala 143:103:@23881.4]
  wire [5:0] _T_77091; // @[Modules.scala 143:103:@23882.4]
  wire [5:0] _T_77103; // @[Modules.scala 143:103:@23892.4]
  wire [4:0] _T_77104; // @[Modules.scala 143:103:@23893.4]
  wire [4:0] _T_77105; // @[Modules.scala 143:103:@23894.4]
  wire [5:0] _T_77152; // @[Modules.scala 143:103:@23934.4]
  wire [4:0] _T_77153; // @[Modules.scala 143:103:@23935.4]
  wire [4:0] _T_77154; // @[Modules.scala 143:103:@23936.4]
  wire [5:0] _T_77166; // @[Modules.scala 143:103:@23946.4]
  wire [4:0] _T_77167; // @[Modules.scala 143:103:@23947.4]
  wire [4:0] _T_77168; // @[Modules.scala 143:103:@23948.4]
  wire [6:0] _T_77187; // @[Modules.scala 143:103:@23964.4]
  wire [5:0] _T_77188; // @[Modules.scala 143:103:@23965.4]
  wire [5:0] _T_77189; // @[Modules.scala 143:103:@23966.4]
  wire [5:0] _T_77194; // @[Modules.scala 143:103:@23970.4]
  wire [4:0] _T_77195; // @[Modules.scala 143:103:@23971.4]
  wire [4:0] _T_77196; // @[Modules.scala 143:103:@23972.4]
  wire [6:0] _T_77215; // @[Modules.scala 143:103:@23988.4]
  wire [5:0] _T_77216; // @[Modules.scala 143:103:@23989.4]
  wire [5:0] _T_77217; // @[Modules.scala 143:103:@23990.4]
  wire [6:0] _T_77222; // @[Modules.scala 143:103:@23994.4]
  wire [5:0] _T_77223; // @[Modules.scala 143:103:@23995.4]
  wire [5:0] _T_77224; // @[Modules.scala 143:103:@23996.4]
  wire [6:0] _T_77229; // @[Modules.scala 143:103:@24000.4]
  wire [5:0] _T_77230; // @[Modules.scala 143:103:@24001.4]
  wire [5:0] _T_77231; // @[Modules.scala 143:103:@24002.4]
  wire [5:0] _T_77243; // @[Modules.scala 143:103:@24012.4]
  wire [4:0] _T_77244; // @[Modules.scala 143:103:@24013.4]
  wire [4:0] _T_77245; // @[Modules.scala 143:103:@24014.4]
  wire [6:0] _T_77250; // @[Modules.scala 143:103:@24018.4]
  wire [5:0] _T_77251; // @[Modules.scala 143:103:@24019.4]
  wire [5:0] _T_77252; // @[Modules.scala 143:103:@24020.4]
  wire [5:0] _T_77257; // @[Modules.scala 143:103:@24024.4]
  wire [4:0] _T_77258; // @[Modules.scala 143:103:@24025.4]
  wire [4:0] _T_77259; // @[Modules.scala 143:103:@24026.4]
  wire [5:0] _GEN_537; // @[Modules.scala 143:103:@24030.4]
  wire [6:0] _T_77264; // @[Modules.scala 143:103:@24030.4]
  wire [5:0] _T_77265; // @[Modules.scala 143:103:@24031.4]
  wire [5:0] _T_77266; // @[Modules.scala 143:103:@24032.4]
  wire [6:0] _T_77278; // @[Modules.scala 143:103:@24042.4]
  wire [5:0] _T_77279; // @[Modules.scala 143:103:@24043.4]
  wire [5:0] _T_77280; // @[Modules.scala 143:103:@24044.4]
  wire [6:0] _T_77327; // @[Modules.scala 143:103:@24084.4]
  wire [5:0] _T_77328; // @[Modules.scala 143:103:@24085.4]
  wire [5:0] _T_77329; // @[Modules.scala 143:103:@24086.4]
  wire [5:0] _T_77334; // @[Modules.scala 143:103:@24090.4]
  wire [4:0] _T_77335; // @[Modules.scala 143:103:@24091.4]
  wire [4:0] _T_77336; // @[Modules.scala 143:103:@24092.4]
  wire [6:0] _T_77355; // @[Modules.scala 143:103:@24108.4]
  wire [5:0] _T_77356; // @[Modules.scala 143:103:@24109.4]
  wire [5:0] _T_77357; // @[Modules.scala 143:103:@24110.4]
  wire [5:0] _T_77382; // @[Modules.scala 144:80:@24131.4]
  wire [6:0] _T_77383; // @[Modules.scala 143:103:@24132.4]
  wire [5:0] _T_77384; // @[Modules.scala 143:103:@24133.4]
  wire [5:0] _T_77385; // @[Modules.scala 143:103:@24134.4]
  wire [6:0] _T_77390; // @[Modules.scala 143:103:@24138.4]
  wire [5:0] _T_77391; // @[Modules.scala 143:103:@24139.4]
  wire [5:0] _T_77392; // @[Modules.scala 143:103:@24140.4]
  wire [6:0] _T_77397; // @[Modules.scala 143:103:@24144.4]
  wire [5:0] _T_77398; // @[Modules.scala 143:103:@24145.4]
  wire [5:0] _T_77399; // @[Modules.scala 143:103:@24146.4]
  wire [6:0] _T_77404; // @[Modules.scala 143:103:@24150.4]
  wire [5:0] _T_77405; // @[Modules.scala 143:103:@24151.4]
  wire [5:0] _T_77406; // @[Modules.scala 143:103:@24152.4]
  wire [5:0] _GEN_540; // @[Modules.scala 143:103:@24156.4]
  wire [6:0] _T_77411; // @[Modules.scala 143:103:@24156.4]
  wire [5:0] _T_77412; // @[Modules.scala 143:103:@24157.4]
  wire [5:0] _T_77413; // @[Modules.scala 143:103:@24158.4]
  wire [5:0] _T_77418; // @[Modules.scala 143:103:@24162.4]
  wire [4:0] _T_77419; // @[Modules.scala 143:103:@24163.4]
  wire [4:0] _T_77420; // @[Modules.scala 143:103:@24164.4]
  wire [6:0] _T_77425; // @[Modules.scala 143:103:@24168.4]
  wire [5:0] _T_77426; // @[Modules.scala 143:103:@24169.4]
  wire [5:0] _T_77427; // @[Modules.scala 143:103:@24170.4]
  wire [6:0] _T_77432; // @[Modules.scala 143:103:@24174.4]
  wire [5:0] _T_77433; // @[Modules.scala 143:103:@24175.4]
  wire [5:0] _T_77434; // @[Modules.scala 143:103:@24176.4]
  wire [5:0] _T_77446; // @[Modules.scala 143:103:@24186.4]
  wire [4:0] _T_77447; // @[Modules.scala 143:103:@24187.4]
  wire [4:0] _T_77448; // @[Modules.scala 143:103:@24188.4]
  wire [5:0] _GEN_542; // @[Modules.scala 143:103:@24198.4]
  wire [6:0] _T_77460; // @[Modules.scala 143:103:@24198.4]
  wire [5:0] _T_77461; // @[Modules.scala 143:103:@24199.4]
  wire [5:0] _T_77462; // @[Modules.scala 143:103:@24200.4]
  wire [5:0] _T_77464; // @[Modules.scala 143:74:@24202.4]
  wire [6:0] _T_77467; // @[Modules.scala 143:103:@24204.4]
  wire [5:0] _T_77468; // @[Modules.scala 143:103:@24205.4]
  wire [5:0] _T_77469; // @[Modules.scala 143:103:@24206.4]
  wire [6:0] _T_77481; // @[Modules.scala 143:103:@24216.4]
  wire [5:0] _T_77482; // @[Modules.scala 143:103:@24217.4]
  wire [5:0] _T_77483; // @[Modules.scala 143:103:@24218.4]
  wire [5:0] _GEN_545; // @[Modules.scala 143:103:@24222.4]
  wire [6:0] _T_77488; // @[Modules.scala 143:103:@24222.4]
  wire [5:0] _T_77489; // @[Modules.scala 143:103:@24223.4]
  wire [5:0] _T_77490; // @[Modules.scala 143:103:@24224.4]
  wire [6:0] _T_77495; // @[Modules.scala 143:103:@24228.4]
  wire [5:0] _T_77496; // @[Modules.scala 143:103:@24229.4]
  wire [5:0] _T_77497; // @[Modules.scala 143:103:@24230.4]
  wire [5:0] _T_77516; // @[Modules.scala 143:103:@24246.4]
  wire [4:0] _T_77517; // @[Modules.scala 143:103:@24247.4]
  wire [4:0] _T_77518; // @[Modules.scala 143:103:@24248.4]
  wire [5:0] _GEN_547; // @[Modules.scala 143:103:@24252.4]
  wire [6:0] _T_77523; // @[Modules.scala 143:103:@24252.4]
  wire [5:0] _T_77524; // @[Modules.scala 143:103:@24253.4]
  wire [5:0] _T_77525; // @[Modules.scala 143:103:@24254.4]
  wire [5:0] _T_77544; // @[Modules.scala 143:103:@24270.4]
  wire [4:0] _T_77545; // @[Modules.scala 143:103:@24271.4]
  wire [4:0] _T_77546; // @[Modules.scala 143:103:@24272.4]
  wire [5:0] _GEN_549; // @[Modules.scala 143:103:@24276.4]
  wire [6:0] _T_77551; // @[Modules.scala 143:103:@24276.4]
  wire [5:0] _T_77552; // @[Modules.scala 143:103:@24277.4]
  wire [5:0] _T_77553; // @[Modules.scala 143:103:@24278.4]
  wire [6:0] _T_77558; // @[Modules.scala 143:103:@24282.4]
  wire [5:0] _T_77559; // @[Modules.scala 143:103:@24283.4]
  wire [5:0] _T_77560; // @[Modules.scala 143:103:@24284.4]
  wire [5:0] _GEN_551; // @[Modules.scala 143:103:@24306.4]
  wire [6:0] _T_77586; // @[Modules.scala 143:103:@24306.4]
  wire [5:0] _T_77587; // @[Modules.scala 143:103:@24307.4]
  wire [5:0] _T_77588; // @[Modules.scala 143:103:@24308.4]
  wire [5:0] _T_77600; // @[Modules.scala 143:103:@24318.4]
  wire [4:0] _T_77601; // @[Modules.scala 143:103:@24319.4]
  wire [4:0] _T_77602; // @[Modules.scala 143:103:@24320.4]
  wire [6:0] _T_77607; // @[Modules.scala 143:103:@24324.4]
  wire [5:0] _T_77608; // @[Modules.scala 143:103:@24325.4]
  wire [5:0] _T_77609; // @[Modules.scala 143:103:@24326.4]
  wire [6:0] _T_77642; // @[Modules.scala 143:103:@24354.4]
  wire [5:0] _T_77643; // @[Modules.scala 143:103:@24355.4]
  wire [5:0] _T_77644; // @[Modules.scala 143:103:@24356.4]
  wire [5:0] _T_77649; // @[Modules.scala 143:103:@24360.4]
  wire [4:0] _T_77650; // @[Modules.scala 143:103:@24361.4]
  wire [4:0] _T_77651; // @[Modules.scala 143:103:@24362.4]
  wire [6:0] _T_77670; // @[Modules.scala 143:103:@24378.4]
  wire [5:0] _T_77671; // @[Modules.scala 143:103:@24379.4]
  wire [5:0] _T_77672; // @[Modules.scala 143:103:@24380.4]
  wire [6:0] _T_77677; // @[Modules.scala 143:103:@24384.4]
  wire [5:0] _T_77678; // @[Modules.scala 143:103:@24385.4]
  wire [5:0] _T_77679; // @[Modules.scala 143:103:@24386.4]
  wire [6:0] _T_77712; // @[Modules.scala 143:103:@24414.4]
  wire [5:0] _T_77713; // @[Modules.scala 143:103:@24415.4]
  wire [5:0] _T_77714; // @[Modules.scala 143:103:@24416.4]
  wire [6:0] _T_77726; // @[Modules.scala 143:103:@24426.4]
  wire [5:0] _T_77727; // @[Modules.scala 143:103:@24427.4]
  wire [5:0] _T_77728; // @[Modules.scala 143:103:@24428.4]
  wire [5:0] _T_77733; // @[Modules.scala 143:103:@24432.4]
  wire [4:0] _T_77734; // @[Modules.scala 143:103:@24433.4]
  wire [4:0] _T_77735; // @[Modules.scala 143:103:@24434.4]
  wire [6:0] _T_77740; // @[Modules.scala 143:103:@24438.4]
  wire [5:0] _T_77741; // @[Modules.scala 143:103:@24439.4]
  wire [5:0] _T_77742; // @[Modules.scala 143:103:@24440.4]
  wire [5:0] _GEN_558; // @[Modules.scala 143:103:@24444.4]
  wire [6:0] _T_77747; // @[Modules.scala 143:103:@24444.4]
  wire [5:0] _T_77748; // @[Modules.scala 143:103:@24445.4]
  wire [5:0] _T_77749; // @[Modules.scala 143:103:@24446.4]
  wire [6:0] _T_77789; // @[Modules.scala 143:103:@24480.4]
  wire [5:0] _T_77790; // @[Modules.scala 143:103:@24481.4]
  wire [5:0] _T_77791; // @[Modules.scala 143:103:@24482.4]
  wire [4:0] _T_77802; // @[Modules.scala 144:80:@24491.4]
  wire [5:0] _T_77803; // @[Modules.scala 143:103:@24492.4]
  wire [4:0] _T_77804; // @[Modules.scala 143:103:@24493.4]
  wire [4:0] _T_77805; // @[Modules.scala 143:103:@24494.4]
  wire [5:0] _GEN_559; // @[Modules.scala 143:103:@24504.4]
  wire [6:0] _T_77817; // @[Modules.scala 143:103:@24504.4]
  wire [5:0] _T_77818; // @[Modules.scala 143:103:@24505.4]
  wire [5:0] _T_77819; // @[Modules.scala 143:103:@24506.4]
  wire [6:0] _T_77838; // @[Modules.scala 143:103:@24522.4]
  wire [5:0] _T_77839; // @[Modules.scala 143:103:@24523.4]
  wire [5:0] _T_77840; // @[Modules.scala 143:103:@24524.4]
  wire [5:0] _GEN_561; // @[Modules.scala 143:103:@24534.4]
  wire [6:0] _T_77852; // @[Modules.scala 143:103:@24534.4]
  wire [5:0] _T_77853; // @[Modules.scala 143:103:@24535.4]
  wire [5:0] _T_77854; // @[Modules.scala 143:103:@24536.4]
  wire [5:0] _GEN_562; // @[Modules.scala 143:103:@24540.4]
  wire [6:0] _T_77859; // @[Modules.scala 143:103:@24540.4]
  wire [5:0] _T_77860; // @[Modules.scala 143:103:@24541.4]
  wire [5:0] _T_77861; // @[Modules.scala 143:103:@24542.4]
  wire [6:0] _T_77866; // @[Modules.scala 143:103:@24546.4]
  wire [5:0] _T_77867; // @[Modules.scala 143:103:@24547.4]
  wire [5:0] _T_77868; // @[Modules.scala 143:103:@24548.4]
  wire [5:0] _GEN_564; // @[Modules.scala 143:103:@24552.4]
  wire [6:0] _T_77873; // @[Modules.scala 143:103:@24552.4]
  wire [5:0] _T_77874; // @[Modules.scala 143:103:@24553.4]
  wire [5:0] _T_77875; // @[Modules.scala 143:103:@24554.4]
  wire [6:0] _T_77887; // @[Modules.scala 143:103:@24564.4]
  wire [5:0] _T_77888; // @[Modules.scala 143:103:@24565.4]
  wire [5:0] _T_77889; // @[Modules.scala 143:103:@24566.4]
  wire [6:0] _T_77915; // @[Modules.scala 143:103:@24588.4]
  wire [5:0] _T_77916; // @[Modules.scala 143:103:@24589.4]
  wire [5:0] _T_77917; // @[Modules.scala 143:103:@24590.4]
  wire [6:0] _T_77922; // @[Modules.scala 143:103:@24594.4]
  wire [5:0] _T_77923; // @[Modules.scala 143:103:@24595.4]
  wire [5:0] _T_77924; // @[Modules.scala 143:103:@24596.4]
  wire [13:0] buffer_7_0; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77925; // @[Modules.scala 166:64:@24598.4]
  wire [13:0] _T_77926; // @[Modules.scala 166:64:@24599.4]
  wire [13:0] buffer_7_309; // @[Modules.scala 166:64:@24600.4]
  wire [14:0] _T_77928; // @[Modules.scala 166:64:@24602.4]
  wire [13:0] _T_77929; // @[Modules.scala 166:64:@24603.4]
  wire [13:0] buffer_7_310; // @[Modules.scala 166:64:@24604.4]
  wire [13:0] buffer_7_4; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77931; // @[Modules.scala 166:64:@24606.4]
  wire [13:0] _T_77932; // @[Modules.scala 166:64:@24607.4]
  wire [13:0] buffer_7_311; // @[Modules.scala 166:64:@24608.4]
  wire [14:0] _T_77934; // @[Modules.scala 166:64:@24610.4]
  wire [13:0] _T_77935; // @[Modules.scala 166:64:@24611.4]
  wire [13:0] buffer_7_312; // @[Modules.scala 166:64:@24612.4]
  wire [13:0] buffer_7_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77937; // @[Modules.scala 166:64:@24614.4]
  wire [13:0] _T_77938; // @[Modules.scala 166:64:@24615.4]
  wire [13:0] buffer_7_313; // @[Modules.scala 166:64:@24616.4]
  wire [13:0] buffer_7_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77943; // @[Modules.scala 166:64:@24622.4]
  wire [13:0] _T_77944; // @[Modules.scala 166:64:@24623.4]
  wire [13:0] buffer_7_315; // @[Modules.scala 166:64:@24624.4]
  wire [14:0] _T_77946; // @[Modules.scala 166:64:@24626.4]
  wire [13:0] _T_77947; // @[Modules.scala 166:64:@24627.4]
  wire [13:0] buffer_7_316; // @[Modules.scala 166:64:@24628.4]
  wire [14:0] _T_77949; // @[Modules.scala 166:64:@24630.4]
  wire [13:0] _T_77950; // @[Modules.scala 166:64:@24631.4]
  wire [13:0] buffer_7_317; // @[Modules.scala 166:64:@24632.4]
  wire [14:0] _T_77952; // @[Modules.scala 166:64:@24634.4]
  wire [13:0] _T_77953; // @[Modules.scala 166:64:@24635.4]
  wire [13:0] buffer_7_318; // @[Modules.scala 166:64:@24636.4]
  wire [13:0] buffer_7_20; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77955; // @[Modules.scala 166:64:@24638.4]
  wire [13:0] _T_77956; // @[Modules.scala 166:64:@24639.4]
  wire [13:0] buffer_7_319; // @[Modules.scala 166:64:@24640.4]
  wire [13:0] buffer_7_22; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77958; // @[Modules.scala 166:64:@24642.4]
  wire [13:0] _T_77959; // @[Modules.scala 166:64:@24643.4]
  wire [13:0] buffer_7_320; // @[Modules.scala 166:64:@24644.4]
  wire [13:0] buffer_7_24; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77961; // @[Modules.scala 166:64:@24646.4]
  wire [13:0] _T_77962; // @[Modules.scala 166:64:@24647.4]
  wire [13:0] buffer_7_321; // @[Modules.scala 166:64:@24648.4]
  wire [14:0] _T_77967; // @[Modules.scala 166:64:@24654.4]
  wire [13:0] _T_77968; // @[Modules.scala 166:64:@24655.4]
  wire [13:0] buffer_7_323; // @[Modules.scala 166:64:@24656.4]
  wire [14:0] _T_77970; // @[Modules.scala 166:64:@24658.4]
  wire [13:0] _T_77971; // @[Modules.scala 166:64:@24659.4]
  wire [13:0] buffer_7_324; // @[Modules.scala 166:64:@24660.4]
  wire [13:0] buffer_7_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77973; // @[Modules.scala 166:64:@24662.4]
  wire [13:0] _T_77974; // @[Modules.scala 166:64:@24663.4]
  wire [13:0] buffer_7_325; // @[Modules.scala 166:64:@24664.4]
  wire [13:0] buffer_7_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77976; // @[Modules.scala 166:64:@24666.4]
  wire [13:0] _T_77977; // @[Modules.scala 166:64:@24667.4]
  wire [13:0] buffer_7_326; // @[Modules.scala 166:64:@24668.4]
  wire [14:0] _T_77979; // @[Modules.scala 166:64:@24670.4]
  wire [13:0] _T_77980; // @[Modules.scala 166:64:@24671.4]
  wire [13:0] buffer_7_327; // @[Modules.scala 166:64:@24672.4]
  wire [13:0] buffer_7_38; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77982; // @[Modules.scala 166:64:@24674.4]
  wire [13:0] _T_77983; // @[Modules.scala 166:64:@24675.4]
  wire [13:0] buffer_7_328; // @[Modules.scala 166:64:@24676.4]
  wire [13:0] buffer_7_40; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77985; // @[Modules.scala 166:64:@24678.4]
  wire [13:0] _T_77986; // @[Modules.scala 166:64:@24679.4]
  wire [13:0] buffer_7_329; // @[Modules.scala 166:64:@24680.4]
  wire [13:0] buffer_7_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77988; // @[Modules.scala 166:64:@24682.4]
  wire [13:0] _T_77989; // @[Modules.scala 166:64:@24683.4]
  wire [13:0] buffer_7_330; // @[Modules.scala 166:64:@24684.4]
  wire [13:0] buffer_7_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77991; // @[Modules.scala 166:64:@24686.4]
  wire [13:0] _T_77992; // @[Modules.scala 166:64:@24687.4]
  wire [13:0] buffer_7_331; // @[Modules.scala 166:64:@24688.4]
  wire [13:0] buffer_7_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_77997; // @[Modules.scala 166:64:@24694.4]
  wire [13:0] _T_77998; // @[Modules.scala 166:64:@24695.4]
  wire [13:0] buffer_7_333; // @[Modules.scala 166:64:@24696.4]
  wire [13:0] buffer_7_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78000; // @[Modules.scala 166:64:@24698.4]
  wire [13:0] _T_78001; // @[Modules.scala 166:64:@24699.4]
  wire [13:0] buffer_7_334; // @[Modules.scala 166:64:@24700.4]
  wire [13:0] buffer_7_52; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78003; // @[Modules.scala 166:64:@24702.4]
  wire [13:0] _T_78004; // @[Modules.scala 166:64:@24703.4]
  wire [13:0] buffer_7_335; // @[Modules.scala 166:64:@24704.4]
  wire [13:0] buffer_7_54; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78006; // @[Modules.scala 166:64:@24706.4]
  wire [13:0] _T_78007; // @[Modules.scala 166:64:@24707.4]
  wire [13:0] buffer_7_336; // @[Modules.scala 166:64:@24708.4]
  wire [13:0] buffer_7_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78009; // @[Modules.scala 166:64:@24710.4]
  wire [13:0] _T_78010; // @[Modules.scala 166:64:@24711.4]
  wire [13:0] buffer_7_337; // @[Modules.scala 166:64:@24712.4]
  wire [14:0] _T_78012; // @[Modules.scala 166:64:@24714.4]
  wire [13:0] _T_78013; // @[Modules.scala 166:64:@24715.4]
  wire [13:0] buffer_7_338; // @[Modules.scala 166:64:@24716.4]
  wire [13:0] buffer_7_60; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78015; // @[Modules.scala 166:64:@24718.4]
  wire [13:0] _T_78016; // @[Modules.scala 166:64:@24719.4]
  wire [13:0] buffer_7_339; // @[Modules.scala 166:64:@24720.4]
  wire [13:0] buffer_7_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78018; // @[Modules.scala 166:64:@24722.4]
  wire [13:0] _T_78019; // @[Modules.scala 166:64:@24723.4]
  wire [13:0] buffer_7_340; // @[Modules.scala 166:64:@24724.4]
  wire [14:0] _T_78021; // @[Modules.scala 166:64:@24726.4]
  wire [13:0] _T_78022; // @[Modules.scala 166:64:@24727.4]
  wire [13:0] buffer_7_341; // @[Modules.scala 166:64:@24728.4]
  wire [13:0] buffer_7_66; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78024; // @[Modules.scala 166:64:@24730.4]
  wire [13:0] _T_78025; // @[Modules.scala 166:64:@24731.4]
  wire [13:0] buffer_7_342; // @[Modules.scala 166:64:@24732.4]
  wire [13:0] buffer_7_68; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78027; // @[Modules.scala 166:64:@24734.4]
  wire [13:0] _T_78028; // @[Modules.scala 166:64:@24735.4]
  wire [13:0] buffer_7_343; // @[Modules.scala 166:64:@24736.4]
  wire [14:0] _T_78030; // @[Modules.scala 166:64:@24738.4]
  wire [13:0] _T_78031; // @[Modules.scala 166:64:@24739.4]
  wire [13:0] buffer_7_344; // @[Modules.scala 166:64:@24740.4]
  wire [14:0] _T_78033; // @[Modules.scala 166:64:@24742.4]
  wire [13:0] _T_78034; // @[Modules.scala 166:64:@24743.4]
  wire [13:0] buffer_7_345; // @[Modules.scala 166:64:@24744.4]
  wire [13:0] buffer_7_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78036; // @[Modules.scala 166:64:@24746.4]
  wire [13:0] _T_78037; // @[Modules.scala 166:64:@24747.4]
  wire [13:0] buffer_7_346; // @[Modules.scala 166:64:@24748.4]
  wire [13:0] buffer_7_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78039; // @[Modules.scala 166:64:@24750.4]
  wire [13:0] _T_78040; // @[Modules.scala 166:64:@24751.4]
  wire [13:0] buffer_7_347; // @[Modules.scala 166:64:@24752.4]
  wire [13:0] buffer_7_82; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_83; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78048; // @[Modules.scala 166:64:@24762.4]
  wire [13:0] _T_78049; // @[Modules.scala 166:64:@24763.4]
  wire [13:0] buffer_7_350; // @[Modules.scala 166:64:@24764.4]
  wire [13:0] buffer_7_84; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78051; // @[Modules.scala 166:64:@24766.4]
  wire [13:0] _T_78052; // @[Modules.scala 166:64:@24767.4]
  wire [13:0] buffer_7_351; // @[Modules.scala 166:64:@24768.4]
  wire [13:0] buffer_7_86; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78054; // @[Modules.scala 166:64:@24770.4]
  wire [13:0] _T_78055; // @[Modules.scala 166:64:@24771.4]
  wire [13:0] buffer_7_352; // @[Modules.scala 166:64:@24772.4]
  wire [14:0] _T_78057; // @[Modules.scala 166:64:@24774.4]
  wire [13:0] _T_78058; // @[Modules.scala 166:64:@24775.4]
  wire [13:0] buffer_7_353; // @[Modules.scala 166:64:@24776.4]
  wire [14:0] _T_78060; // @[Modules.scala 166:64:@24778.4]
  wire [13:0] _T_78061; // @[Modules.scala 166:64:@24779.4]
  wire [13:0] buffer_7_354; // @[Modules.scala 166:64:@24780.4]
  wire [14:0] _T_78063; // @[Modules.scala 166:64:@24782.4]
  wire [13:0] _T_78064; // @[Modules.scala 166:64:@24783.4]
  wire [13:0] buffer_7_355; // @[Modules.scala 166:64:@24784.4]
  wire [14:0] _T_78066; // @[Modules.scala 166:64:@24786.4]
  wire [13:0] _T_78067; // @[Modules.scala 166:64:@24787.4]
  wire [13:0] buffer_7_356; // @[Modules.scala 166:64:@24788.4]
  wire [14:0] _T_78069; // @[Modules.scala 166:64:@24790.4]
  wire [13:0] _T_78070; // @[Modules.scala 166:64:@24791.4]
  wire [13:0] buffer_7_357; // @[Modules.scala 166:64:@24792.4]
  wire [13:0] buffer_7_100; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78075; // @[Modules.scala 166:64:@24798.4]
  wire [13:0] _T_78076; // @[Modules.scala 166:64:@24799.4]
  wire [13:0] buffer_7_359; // @[Modules.scala 166:64:@24800.4]
  wire [14:0] _T_78078; // @[Modules.scala 166:64:@24802.4]
  wire [13:0] _T_78079; // @[Modules.scala 166:64:@24803.4]
  wire [13:0] buffer_7_360; // @[Modules.scala 166:64:@24804.4]
  wire [14:0] _T_78081; // @[Modules.scala 166:64:@24806.4]
  wire [13:0] _T_78082; // @[Modules.scala 166:64:@24807.4]
  wire [13:0] buffer_7_361; // @[Modules.scala 166:64:@24808.4]
  wire [14:0] _T_78084; // @[Modules.scala 166:64:@24810.4]
  wire [13:0] _T_78085; // @[Modules.scala 166:64:@24811.4]
  wire [13:0] buffer_7_362; // @[Modules.scala 166:64:@24812.4]
  wire [13:0] buffer_7_112; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78093; // @[Modules.scala 166:64:@24822.4]
  wire [13:0] _T_78094; // @[Modules.scala 166:64:@24823.4]
  wire [13:0] buffer_7_365; // @[Modules.scala 166:64:@24824.4]
  wire [13:0] buffer_7_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78096; // @[Modules.scala 166:64:@24826.4]
  wire [13:0] _T_78097; // @[Modules.scala 166:64:@24827.4]
  wire [13:0] buffer_7_366; // @[Modules.scala 166:64:@24828.4]
  wire [14:0] _T_78099; // @[Modules.scala 166:64:@24830.4]
  wire [13:0] _T_78100; // @[Modules.scala 166:64:@24831.4]
  wire [13:0] buffer_7_367; // @[Modules.scala 166:64:@24832.4]
  wire [14:0] _T_78102; // @[Modules.scala 166:64:@24834.4]
  wire [13:0] _T_78103; // @[Modules.scala 166:64:@24835.4]
  wire [13:0] buffer_7_368; // @[Modules.scala 166:64:@24836.4]
  wire [13:0] buffer_7_120; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78105; // @[Modules.scala 166:64:@24838.4]
  wire [13:0] _T_78106; // @[Modules.scala 166:64:@24839.4]
  wire [13:0] buffer_7_369; // @[Modules.scala 166:64:@24840.4]
  wire [14:0] _T_78108; // @[Modules.scala 166:64:@24842.4]
  wire [13:0] _T_78109; // @[Modules.scala 166:64:@24843.4]
  wire [13:0] buffer_7_370; // @[Modules.scala 166:64:@24844.4]
  wire [13:0] buffer_7_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78111; // @[Modules.scala 166:64:@24846.4]
  wire [13:0] _T_78112; // @[Modules.scala 166:64:@24847.4]
  wire [13:0] buffer_7_371; // @[Modules.scala 166:64:@24848.4]
  wire [13:0] buffer_7_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78114; // @[Modules.scala 166:64:@24850.4]
  wire [13:0] _T_78115; // @[Modules.scala 166:64:@24851.4]
  wire [13:0] buffer_7_372; // @[Modules.scala 166:64:@24852.4]
  wire [13:0] buffer_7_129; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78117; // @[Modules.scala 166:64:@24854.4]
  wire [13:0] _T_78118; // @[Modules.scala 166:64:@24855.4]
  wire [13:0] buffer_7_373; // @[Modules.scala 166:64:@24856.4]
  wire [13:0] buffer_7_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78123; // @[Modules.scala 166:64:@24862.4]
  wire [13:0] _T_78124; // @[Modules.scala 166:64:@24863.4]
  wire [13:0] buffer_7_375; // @[Modules.scala 166:64:@24864.4]
  wire [14:0] _T_78126; // @[Modules.scala 166:64:@24866.4]
  wire [13:0] _T_78127; // @[Modules.scala 166:64:@24867.4]
  wire [13:0] buffer_7_376; // @[Modules.scala 166:64:@24868.4]
  wire [14:0] _T_78129; // @[Modules.scala 166:64:@24870.4]
  wire [13:0] _T_78130; // @[Modules.scala 166:64:@24871.4]
  wire [13:0] buffer_7_377; // @[Modules.scala 166:64:@24872.4]
  wire [14:0] _T_78132; // @[Modules.scala 166:64:@24874.4]
  wire [13:0] _T_78133; // @[Modules.scala 166:64:@24875.4]
  wire [13:0] buffer_7_378; // @[Modules.scala 166:64:@24876.4]
  wire [14:0] _T_78135; // @[Modules.scala 166:64:@24878.4]
  wire [13:0] _T_78136; // @[Modules.scala 166:64:@24879.4]
  wire [13:0] buffer_7_379; // @[Modules.scala 166:64:@24880.4]
  wire [14:0] _T_78138; // @[Modules.scala 166:64:@24882.4]
  wire [13:0] _T_78139; // @[Modules.scala 166:64:@24883.4]
  wire [13:0] buffer_7_380; // @[Modules.scala 166:64:@24884.4]
  wire [13:0] buffer_7_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78141; // @[Modules.scala 166:64:@24886.4]
  wire [13:0] _T_78142; // @[Modules.scala 166:64:@24887.4]
  wire [13:0] buffer_7_381; // @[Modules.scala 166:64:@24888.4]
  wire [13:0] buffer_7_146; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78144; // @[Modules.scala 166:64:@24890.4]
  wire [13:0] _T_78145; // @[Modules.scala 166:64:@24891.4]
  wire [13:0] buffer_7_382; // @[Modules.scala 166:64:@24892.4]
  wire [13:0] buffer_7_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78147; // @[Modules.scala 166:64:@24894.4]
  wire [13:0] _T_78148; // @[Modules.scala 166:64:@24895.4]
  wire [13:0] buffer_7_383; // @[Modules.scala 166:64:@24896.4]
  wire [13:0] buffer_7_150; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78150; // @[Modules.scala 166:64:@24898.4]
  wire [13:0] _T_78151; // @[Modules.scala 166:64:@24899.4]
  wire [13:0] buffer_7_384; // @[Modules.scala 166:64:@24900.4]
  wire [13:0] buffer_7_152; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78153; // @[Modules.scala 166:64:@24902.4]
  wire [13:0] _T_78154; // @[Modules.scala 166:64:@24903.4]
  wire [13:0] buffer_7_385; // @[Modules.scala 166:64:@24904.4]
  wire [13:0] buffer_7_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78159; // @[Modules.scala 166:64:@24910.4]
  wire [13:0] _T_78160; // @[Modules.scala 166:64:@24911.4]
  wire [13:0] buffer_7_387; // @[Modules.scala 166:64:@24912.4]
  wire [13:0] buffer_7_158; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78162; // @[Modules.scala 166:64:@24914.4]
  wire [13:0] _T_78163; // @[Modules.scala 166:64:@24915.4]
  wire [13:0] buffer_7_388; // @[Modules.scala 166:64:@24916.4]
  wire [14:0] _T_78165; // @[Modules.scala 166:64:@24918.4]
  wire [13:0] _T_78166; // @[Modules.scala 166:64:@24919.4]
  wire [13:0] buffer_7_389; // @[Modules.scala 166:64:@24920.4]
  wire [13:0] buffer_7_162; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78168; // @[Modules.scala 166:64:@24922.4]
  wire [13:0] _T_78169; // @[Modules.scala 166:64:@24923.4]
  wire [13:0] buffer_7_390; // @[Modules.scala 166:64:@24924.4]
  wire [13:0] buffer_7_164; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78171; // @[Modules.scala 166:64:@24926.4]
  wire [13:0] _T_78172; // @[Modules.scala 166:64:@24927.4]
  wire [13:0] buffer_7_391; // @[Modules.scala 166:64:@24928.4]
  wire [14:0] _T_78174; // @[Modules.scala 166:64:@24930.4]
  wire [13:0] _T_78175; // @[Modules.scala 166:64:@24931.4]
  wire [13:0] buffer_7_392; // @[Modules.scala 166:64:@24932.4]
  wire [13:0] buffer_7_168; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78177; // @[Modules.scala 166:64:@24934.4]
  wire [13:0] _T_78178; // @[Modules.scala 166:64:@24935.4]
  wire [13:0] buffer_7_393; // @[Modules.scala 166:64:@24936.4]
  wire [13:0] buffer_7_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78180; // @[Modules.scala 166:64:@24938.4]
  wire [13:0] _T_78181; // @[Modules.scala 166:64:@24939.4]
  wire [13:0] buffer_7_394; // @[Modules.scala 166:64:@24940.4]
  wire [14:0] _T_78183; // @[Modules.scala 166:64:@24942.4]
  wire [13:0] _T_78184; // @[Modules.scala 166:64:@24943.4]
  wire [13:0] buffer_7_395; // @[Modules.scala 166:64:@24944.4]
  wire [14:0] _T_78186; // @[Modules.scala 166:64:@24946.4]
  wire [13:0] _T_78187; // @[Modules.scala 166:64:@24947.4]
  wire [13:0] buffer_7_396; // @[Modules.scala 166:64:@24948.4]
  wire [13:0] buffer_7_176; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78189; // @[Modules.scala 166:64:@24950.4]
  wire [13:0] _T_78190; // @[Modules.scala 166:64:@24951.4]
  wire [13:0] buffer_7_397; // @[Modules.scala 166:64:@24952.4]
  wire [14:0] _T_78192; // @[Modules.scala 166:64:@24954.4]
  wire [13:0] _T_78193; // @[Modules.scala 166:64:@24955.4]
  wire [13:0] buffer_7_398; // @[Modules.scala 166:64:@24956.4]
  wire [14:0] _T_78198; // @[Modules.scala 166:64:@24962.4]
  wire [13:0] _T_78199; // @[Modules.scala 166:64:@24963.4]
  wire [13:0] buffer_7_400; // @[Modules.scala 166:64:@24964.4]
  wire [14:0] _T_78201; // @[Modules.scala 166:64:@24966.4]
  wire [13:0] _T_78202; // @[Modules.scala 166:64:@24967.4]
  wire [13:0] buffer_7_401; // @[Modules.scala 166:64:@24968.4]
  wire [14:0] _T_78204; // @[Modules.scala 166:64:@24970.4]
  wire [13:0] _T_78205; // @[Modules.scala 166:64:@24971.4]
  wire [13:0] buffer_7_402; // @[Modules.scala 166:64:@24972.4]
  wire [13:0] buffer_7_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78207; // @[Modules.scala 166:64:@24974.4]
  wire [13:0] _T_78208; // @[Modules.scala 166:64:@24975.4]
  wire [13:0] buffer_7_403; // @[Modules.scala 166:64:@24976.4]
  wire [13:0] buffer_7_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78210; // @[Modules.scala 166:64:@24978.4]
  wire [13:0] _T_78211; // @[Modules.scala 166:64:@24979.4]
  wire [13:0] buffer_7_404; // @[Modules.scala 166:64:@24980.4]
  wire [14:0] _T_78213; // @[Modules.scala 166:64:@24982.4]
  wire [13:0] _T_78214; // @[Modules.scala 166:64:@24983.4]
  wire [13:0] buffer_7_405; // @[Modules.scala 166:64:@24984.4]
  wire [14:0] _T_78216; // @[Modules.scala 166:64:@24986.4]
  wire [13:0] _T_78217; // @[Modules.scala 166:64:@24987.4]
  wire [13:0] buffer_7_406; // @[Modules.scala 166:64:@24988.4]
  wire [13:0] buffer_7_198; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78222; // @[Modules.scala 166:64:@24994.4]
  wire [13:0] _T_78223; // @[Modules.scala 166:64:@24995.4]
  wire [13:0] buffer_7_408; // @[Modules.scala 166:64:@24996.4]
  wire [13:0] buffer_7_200; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78225; // @[Modules.scala 166:64:@24998.4]
  wire [13:0] _T_78226; // @[Modules.scala 166:64:@24999.4]
  wire [13:0] buffer_7_409; // @[Modules.scala 166:64:@25000.4]
  wire [13:0] buffer_7_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78228; // @[Modules.scala 166:64:@25002.4]
  wire [13:0] _T_78229; // @[Modules.scala 166:64:@25003.4]
  wire [13:0] buffer_7_410; // @[Modules.scala 166:64:@25004.4]
  wire [13:0] buffer_7_204; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78231; // @[Modules.scala 166:64:@25006.4]
  wire [13:0] _T_78232; // @[Modules.scala 166:64:@25007.4]
  wire [13:0] buffer_7_411; // @[Modules.scala 166:64:@25008.4]
  wire [13:0] buffer_7_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78234; // @[Modules.scala 166:64:@25010.4]
  wire [13:0] _T_78235; // @[Modules.scala 166:64:@25011.4]
  wire [13:0] buffer_7_412; // @[Modules.scala 166:64:@25012.4]
  wire [13:0] buffer_7_208; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_209; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78237; // @[Modules.scala 166:64:@25014.4]
  wire [13:0] _T_78238; // @[Modules.scala 166:64:@25015.4]
  wire [13:0] buffer_7_413; // @[Modules.scala 166:64:@25016.4]
  wire [13:0] buffer_7_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78240; // @[Modules.scala 166:64:@25018.4]
  wire [13:0] _T_78241; // @[Modules.scala 166:64:@25019.4]
  wire [13:0] buffer_7_414; // @[Modules.scala 166:64:@25020.4]
  wire [13:0] buffer_7_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78243; // @[Modules.scala 166:64:@25022.4]
  wire [13:0] _T_78244; // @[Modules.scala 166:64:@25023.4]
  wire [13:0] buffer_7_415; // @[Modules.scala 166:64:@25024.4]
  wire [13:0] buffer_7_214; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78246; // @[Modules.scala 166:64:@25026.4]
  wire [13:0] _T_78247; // @[Modules.scala 166:64:@25027.4]
  wire [13:0] buffer_7_416; // @[Modules.scala 166:64:@25028.4]
  wire [13:0] buffer_7_216; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78249; // @[Modules.scala 166:64:@25030.4]
  wire [13:0] _T_78250; // @[Modules.scala 166:64:@25031.4]
  wire [13:0] buffer_7_417; // @[Modules.scala 166:64:@25032.4]
  wire [14:0] _T_78252; // @[Modules.scala 166:64:@25034.4]
  wire [13:0] _T_78253; // @[Modules.scala 166:64:@25035.4]
  wire [13:0] buffer_7_418; // @[Modules.scala 166:64:@25036.4]
  wire [14:0] _T_78255; // @[Modules.scala 166:64:@25038.4]
  wire [13:0] _T_78256; // @[Modules.scala 166:64:@25039.4]
  wire [13:0] buffer_7_419; // @[Modules.scala 166:64:@25040.4]
  wire [13:0] buffer_7_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78258; // @[Modules.scala 166:64:@25042.4]
  wire [13:0] _T_78259; // @[Modules.scala 166:64:@25043.4]
  wire [13:0] buffer_7_420; // @[Modules.scala 166:64:@25044.4]
  wire [13:0] buffer_7_224; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78261; // @[Modules.scala 166:64:@25046.4]
  wire [13:0] _T_78262; // @[Modules.scala 166:64:@25047.4]
  wire [13:0] buffer_7_421; // @[Modules.scala 166:64:@25048.4]
  wire [13:0] buffer_7_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78264; // @[Modules.scala 166:64:@25050.4]
  wire [13:0] _T_78265; // @[Modules.scala 166:64:@25051.4]
  wire [13:0] buffer_7_422; // @[Modules.scala 166:64:@25052.4]
  wire [14:0] _T_78267; // @[Modules.scala 166:64:@25054.4]
  wire [13:0] _T_78268; // @[Modules.scala 166:64:@25055.4]
  wire [13:0] buffer_7_423; // @[Modules.scala 166:64:@25056.4]
  wire [13:0] buffer_7_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78270; // @[Modules.scala 166:64:@25058.4]
  wire [13:0] _T_78271; // @[Modules.scala 166:64:@25059.4]
  wire [13:0] buffer_7_424; // @[Modules.scala 166:64:@25060.4]
  wire [13:0] buffer_7_232; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78273; // @[Modules.scala 166:64:@25062.4]
  wire [13:0] _T_78274; // @[Modules.scala 166:64:@25063.4]
  wire [13:0] buffer_7_425; // @[Modules.scala 166:64:@25064.4]
  wire [13:0] buffer_7_234; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78276; // @[Modules.scala 166:64:@25066.4]
  wire [13:0] _T_78277; // @[Modules.scala 166:64:@25067.4]
  wire [13:0] buffer_7_426; // @[Modules.scala 166:64:@25068.4]
  wire [13:0] buffer_7_236; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78279; // @[Modules.scala 166:64:@25070.4]
  wire [13:0] _T_78280; // @[Modules.scala 166:64:@25071.4]
  wire [13:0] buffer_7_427; // @[Modules.scala 166:64:@25072.4]
  wire [13:0] buffer_7_238; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78282; // @[Modules.scala 166:64:@25074.4]
  wire [13:0] _T_78283; // @[Modules.scala 166:64:@25075.4]
  wire [13:0] buffer_7_428; // @[Modules.scala 166:64:@25076.4]
  wire [13:0] buffer_7_240; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78285; // @[Modules.scala 166:64:@25078.4]
  wire [13:0] _T_78286; // @[Modules.scala 166:64:@25079.4]
  wire [13:0] buffer_7_429; // @[Modules.scala 166:64:@25080.4]
  wire [13:0] buffer_7_242; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78288; // @[Modules.scala 166:64:@25082.4]
  wire [13:0] _T_78289; // @[Modules.scala 166:64:@25083.4]
  wire [13:0] buffer_7_430; // @[Modules.scala 166:64:@25084.4]
  wire [13:0] buffer_7_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78291; // @[Modules.scala 166:64:@25086.4]
  wire [13:0] _T_78292; // @[Modules.scala 166:64:@25087.4]
  wire [13:0] buffer_7_431; // @[Modules.scala 166:64:@25088.4]
  wire [13:0] buffer_7_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78294; // @[Modules.scala 166:64:@25090.4]
  wire [13:0] _T_78295; // @[Modules.scala 166:64:@25091.4]
  wire [13:0] buffer_7_432; // @[Modules.scala 166:64:@25092.4]
  wire [13:0] buffer_7_250; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78300; // @[Modules.scala 166:64:@25098.4]
  wire [13:0] _T_78301; // @[Modules.scala 166:64:@25099.4]
  wire [13:0] buffer_7_434; // @[Modules.scala 166:64:@25100.4]
  wire [14:0] _T_78303; // @[Modules.scala 166:64:@25102.4]
  wire [13:0] _T_78304; // @[Modules.scala 166:64:@25103.4]
  wire [13:0] buffer_7_435; // @[Modules.scala 166:64:@25104.4]
  wire [13:0] buffer_7_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78306; // @[Modules.scala 166:64:@25106.4]
  wire [13:0] _T_78307; // @[Modules.scala 166:64:@25107.4]
  wire [13:0] buffer_7_436; // @[Modules.scala 166:64:@25108.4]
  wire [13:0] buffer_7_256; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78309; // @[Modules.scala 166:64:@25110.4]
  wire [13:0] _T_78310; // @[Modules.scala 166:64:@25111.4]
  wire [13:0] buffer_7_437; // @[Modules.scala 166:64:@25112.4]
  wire [14:0] _T_78312; // @[Modules.scala 166:64:@25114.4]
  wire [13:0] _T_78313; // @[Modules.scala 166:64:@25115.4]
  wire [13:0] buffer_7_438; // @[Modules.scala 166:64:@25116.4]
  wire [13:0] buffer_7_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78315; // @[Modules.scala 166:64:@25118.4]
  wire [13:0] _T_78316; // @[Modules.scala 166:64:@25119.4]
  wire [13:0] buffer_7_439; // @[Modules.scala 166:64:@25120.4]
  wire [13:0] buffer_7_262; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78318; // @[Modules.scala 166:64:@25122.4]
  wire [13:0] _T_78319; // @[Modules.scala 166:64:@25123.4]
  wire [13:0] buffer_7_440; // @[Modules.scala 166:64:@25124.4]
  wire [14:0] _T_78324; // @[Modules.scala 166:64:@25130.4]
  wire [13:0] _T_78325; // @[Modules.scala 166:64:@25131.4]
  wire [13:0] buffer_7_442; // @[Modules.scala 166:64:@25132.4]
  wire [13:0] buffer_7_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78327; // @[Modules.scala 166:64:@25134.4]
  wire [13:0] _T_78328; // @[Modules.scala 166:64:@25135.4]
  wire [13:0] buffer_7_443; // @[Modules.scala 166:64:@25136.4]
  wire [14:0] _T_78330; // @[Modules.scala 166:64:@25138.4]
  wire [13:0] _T_78331; // @[Modules.scala 166:64:@25139.4]
  wire [13:0] buffer_7_444; // @[Modules.scala 166:64:@25140.4]
  wire [13:0] buffer_7_272; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78333; // @[Modules.scala 166:64:@25142.4]
  wire [13:0] _T_78334; // @[Modules.scala 166:64:@25143.4]
  wire [13:0] buffer_7_445; // @[Modules.scala 166:64:@25144.4]
  wire [13:0] buffer_7_278; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78342; // @[Modules.scala 166:64:@25154.4]
  wire [13:0] _T_78343; // @[Modules.scala 166:64:@25155.4]
  wire [13:0] buffer_7_448; // @[Modules.scala 166:64:@25156.4]
  wire [13:0] buffer_7_280; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78345; // @[Modules.scala 166:64:@25158.4]
  wire [13:0] _T_78346; // @[Modules.scala 166:64:@25159.4]
  wire [13:0] buffer_7_449; // @[Modules.scala 166:64:@25160.4]
  wire [13:0] buffer_7_282; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_283; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78348; // @[Modules.scala 166:64:@25162.4]
  wire [13:0] _T_78349; // @[Modules.scala 166:64:@25163.4]
  wire [13:0] buffer_7_450; // @[Modules.scala 166:64:@25164.4]
  wire [14:0] _T_78351; // @[Modules.scala 166:64:@25166.4]
  wire [13:0] _T_78352; // @[Modules.scala 166:64:@25167.4]
  wire [13:0] buffer_7_451; // @[Modules.scala 166:64:@25168.4]
  wire [14:0] _T_78354; // @[Modules.scala 166:64:@25170.4]
  wire [13:0] _T_78355; // @[Modules.scala 166:64:@25171.4]
  wire [13:0] buffer_7_452; // @[Modules.scala 166:64:@25172.4]
  wire [13:0] buffer_7_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78357; // @[Modules.scala 166:64:@25174.4]
  wire [13:0] _T_78358; // @[Modules.scala 166:64:@25175.4]
  wire [13:0] buffer_7_453; // @[Modules.scala 166:64:@25176.4]
  wire [13:0] buffer_7_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78360; // @[Modules.scala 166:64:@25178.4]
  wire [13:0] _T_78361; // @[Modules.scala 166:64:@25179.4]
  wire [13:0] buffer_7_454; // @[Modules.scala 166:64:@25180.4]
  wire [13:0] buffer_7_293; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78363; // @[Modules.scala 166:64:@25182.4]
  wire [13:0] _T_78364; // @[Modules.scala 166:64:@25183.4]
  wire [13:0] buffer_7_455; // @[Modules.scala 166:64:@25184.4]
  wire [14:0] _T_78366; // @[Modules.scala 166:64:@25186.4]
  wire [13:0] _T_78367; // @[Modules.scala 166:64:@25187.4]
  wire [13:0] buffer_7_456; // @[Modules.scala 166:64:@25188.4]
  wire [13:0] buffer_7_296; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78369; // @[Modules.scala 166:64:@25190.4]
  wire [13:0] _T_78370; // @[Modules.scala 166:64:@25191.4]
  wire [13:0] buffer_7_457; // @[Modules.scala 166:64:@25192.4]
  wire [13:0] buffer_7_298; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78372; // @[Modules.scala 166:64:@25194.4]
  wire [13:0] _T_78373; // @[Modules.scala 166:64:@25195.4]
  wire [13:0] buffer_7_458; // @[Modules.scala 166:64:@25196.4]
  wire [13:0] buffer_7_300; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_7_301; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78375; // @[Modules.scala 166:64:@25198.4]
  wire [13:0] _T_78376; // @[Modules.scala 166:64:@25199.4]
  wire [13:0] buffer_7_459; // @[Modules.scala 166:64:@25200.4]
  wire [13:0] buffer_7_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78378; // @[Modules.scala 166:64:@25202.4]
  wire [13:0] _T_78379; // @[Modules.scala 166:64:@25203.4]
  wire [13:0] buffer_7_460; // @[Modules.scala 166:64:@25204.4]
  wire [13:0] buffer_7_307; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78384; // @[Modules.scala 166:64:@25210.4]
  wire [13:0] _T_78385; // @[Modules.scala 166:64:@25211.4]
  wire [13:0] buffer_7_462; // @[Modules.scala 166:64:@25212.4]
  wire [14:0] _T_78387; // @[Modules.scala 160:64:@25214.4]
  wire [13:0] _T_78388; // @[Modules.scala 160:64:@25215.4]
  wire [13:0] buffer_7_463; // @[Modules.scala 160:64:@25216.4]
  wire [14:0] _T_78390; // @[Modules.scala 160:64:@25218.4]
  wire [13:0] _T_78391; // @[Modules.scala 160:64:@25219.4]
  wire [13:0] buffer_7_464; // @[Modules.scala 160:64:@25220.4]
  wire [14:0] _T_78393; // @[Modules.scala 160:64:@25222.4]
  wire [13:0] _T_78394; // @[Modules.scala 160:64:@25223.4]
  wire [13:0] buffer_7_465; // @[Modules.scala 160:64:@25224.4]
  wire [14:0] _T_78396; // @[Modules.scala 160:64:@25226.4]
  wire [13:0] _T_78397; // @[Modules.scala 160:64:@25227.4]
  wire [13:0] buffer_7_466; // @[Modules.scala 160:64:@25228.4]
  wire [14:0] _T_78399; // @[Modules.scala 160:64:@25230.4]
  wire [13:0] _T_78400; // @[Modules.scala 160:64:@25231.4]
  wire [13:0] buffer_7_467; // @[Modules.scala 160:64:@25232.4]
  wire [14:0] _T_78402; // @[Modules.scala 160:64:@25234.4]
  wire [13:0] _T_78403; // @[Modules.scala 160:64:@25235.4]
  wire [13:0] buffer_7_468; // @[Modules.scala 160:64:@25236.4]
  wire [14:0] _T_78405; // @[Modules.scala 160:64:@25238.4]
  wire [13:0] _T_78406; // @[Modules.scala 160:64:@25239.4]
  wire [13:0] buffer_7_469; // @[Modules.scala 160:64:@25240.4]
  wire [14:0] _T_78408; // @[Modules.scala 160:64:@25242.4]
  wire [13:0] _T_78409; // @[Modules.scala 160:64:@25243.4]
  wire [13:0] buffer_7_470; // @[Modules.scala 160:64:@25244.4]
  wire [14:0] _T_78411; // @[Modules.scala 160:64:@25246.4]
  wire [13:0] _T_78412; // @[Modules.scala 160:64:@25247.4]
  wire [13:0] buffer_7_471; // @[Modules.scala 160:64:@25248.4]
  wire [14:0] _T_78414; // @[Modules.scala 160:64:@25250.4]
  wire [13:0] _T_78415; // @[Modules.scala 160:64:@25251.4]
  wire [13:0] buffer_7_472; // @[Modules.scala 160:64:@25252.4]
  wire [14:0] _T_78417; // @[Modules.scala 160:64:@25254.4]
  wire [13:0] _T_78418; // @[Modules.scala 160:64:@25255.4]
  wire [13:0] buffer_7_473; // @[Modules.scala 160:64:@25256.4]
  wire [14:0] _T_78420; // @[Modules.scala 160:64:@25258.4]
  wire [13:0] _T_78421; // @[Modules.scala 160:64:@25259.4]
  wire [13:0] buffer_7_474; // @[Modules.scala 160:64:@25260.4]
  wire [14:0] _T_78423; // @[Modules.scala 160:64:@25262.4]
  wire [13:0] _T_78424; // @[Modules.scala 160:64:@25263.4]
  wire [13:0] buffer_7_475; // @[Modules.scala 160:64:@25264.4]
  wire [14:0] _T_78426; // @[Modules.scala 160:64:@25266.4]
  wire [13:0] _T_78427; // @[Modules.scala 160:64:@25267.4]
  wire [13:0] buffer_7_476; // @[Modules.scala 160:64:@25268.4]
  wire [14:0] _T_78429; // @[Modules.scala 160:64:@25270.4]
  wire [13:0] _T_78430; // @[Modules.scala 160:64:@25271.4]
  wire [13:0] buffer_7_477; // @[Modules.scala 160:64:@25272.4]
  wire [14:0] _T_78432; // @[Modules.scala 160:64:@25274.4]
  wire [13:0] _T_78433; // @[Modules.scala 160:64:@25275.4]
  wire [13:0] buffer_7_478; // @[Modules.scala 160:64:@25276.4]
  wire [14:0] _T_78435; // @[Modules.scala 160:64:@25278.4]
  wire [13:0] _T_78436; // @[Modules.scala 160:64:@25279.4]
  wire [13:0] buffer_7_479; // @[Modules.scala 160:64:@25280.4]
  wire [14:0] _T_78438; // @[Modules.scala 160:64:@25282.4]
  wire [13:0] _T_78439; // @[Modules.scala 160:64:@25283.4]
  wire [13:0] buffer_7_480; // @[Modules.scala 160:64:@25284.4]
  wire [14:0] _T_78441; // @[Modules.scala 160:64:@25286.4]
  wire [13:0] _T_78442; // @[Modules.scala 160:64:@25287.4]
  wire [13:0] buffer_7_481; // @[Modules.scala 160:64:@25288.4]
  wire [14:0] _T_78444; // @[Modules.scala 160:64:@25290.4]
  wire [13:0] _T_78445; // @[Modules.scala 160:64:@25291.4]
  wire [13:0] buffer_7_482; // @[Modules.scala 160:64:@25292.4]
  wire [14:0] _T_78447; // @[Modules.scala 160:64:@25294.4]
  wire [13:0] _T_78448; // @[Modules.scala 160:64:@25295.4]
  wire [13:0] buffer_7_483; // @[Modules.scala 160:64:@25296.4]
  wire [14:0] _T_78450; // @[Modules.scala 160:64:@25298.4]
  wire [13:0] _T_78451; // @[Modules.scala 160:64:@25299.4]
  wire [13:0] buffer_7_484; // @[Modules.scala 160:64:@25300.4]
  wire [14:0] _T_78453; // @[Modules.scala 160:64:@25302.4]
  wire [13:0] _T_78454; // @[Modules.scala 160:64:@25303.4]
  wire [13:0] buffer_7_485; // @[Modules.scala 160:64:@25304.4]
  wire [14:0] _T_78456; // @[Modules.scala 160:64:@25306.4]
  wire [13:0] _T_78457; // @[Modules.scala 160:64:@25307.4]
  wire [13:0] buffer_7_486; // @[Modules.scala 160:64:@25308.4]
  wire [14:0] _T_78459; // @[Modules.scala 160:64:@25310.4]
  wire [13:0] _T_78460; // @[Modules.scala 160:64:@25311.4]
  wire [13:0] buffer_7_487; // @[Modules.scala 160:64:@25312.4]
  wire [14:0] _T_78462; // @[Modules.scala 160:64:@25314.4]
  wire [13:0] _T_78463; // @[Modules.scala 160:64:@25315.4]
  wire [13:0] buffer_7_488; // @[Modules.scala 160:64:@25316.4]
  wire [14:0] _T_78465; // @[Modules.scala 160:64:@25318.4]
  wire [13:0] _T_78466; // @[Modules.scala 160:64:@25319.4]
  wire [13:0] buffer_7_489; // @[Modules.scala 160:64:@25320.4]
  wire [14:0] _T_78468; // @[Modules.scala 160:64:@25322.4]
  wire [13:0] _T_78469; // @[Modules.scala 160:64:@25323.4]
  wire [13:0] buffer_7_490; // @[Modules.scala 160:64:@25324.4]
  wire [14:0] _T_78471; // @[Modules.scala 160:64:@25326.4]
  wire [13:0] _T_78472; // @[Modules.scala 160:64:@25327.4]
  wire [13:0] buffer_7_491; // @[Modules.scala 160:64:@25328.4]
  wire [14:0] _T_78474; // @[Modules.scala 160:64:@25330.4]
  wire [13:0] _T_78475; // @[Modules.scala 160:64:@25331.4]
  wire [13:0] buffer_7_492; // @[Modules.scala 160:64:@25332.4]
  wire [14:0] _T_78477; // @[Modules.scala 160:64:@25334.4]
  wire [13:0] _T_78478; // @[Modules.scala 160:64:@25335.4]
  wire [13:0] buffer_7_493; // @[Modules.scala 160:64:@25336.4]
  wire [14:0] _T_78480; // @[Modules.scala 160:64:@25338.4]
  wire [13:0] _T_78481; // @[Modules.scala 160:64:@25339.4]
  wire [13:0] buffer_7_494; // @[Modules.scala 160:64:@25340.4]
  wire [14:0] _T_78483; // @[Modules.scala 160:64:@25342.4]
  wire [13:0] _T_78484; // @[Modules.scala 160:64:@25343.4]
  wire [13:0] buffer_7_495; // @[Modules.scala 160:64:@25344.4]
  wire [14:0] _T_78486; // @[Modules.scala 160:64:@25346.4]
  wire [13:0] _T_78487; // @[Modules.scala 160:64:@25347.4]
  wire [13:0] buffer_7_496; // @[Modules.scala 160:64:@25348.4]
  wire [14:0] _T_78489; // @[Modules.scala 160:64:@25350.4]
  wire [13:0] _T_78490; // @[Modules.scala 160:64:@25351.4]
  wire [13:0] buffer_7_497; // @[Modules.scala 160:64:@25352.4]
  wire [14:0] _T_78492; // @[Modules.scala 160:64:@25354.4]
  wire [13:0] _T_78493; // @[Modules.scala 160:64:@25355.4]
  wire [13:0] buffer_7_498; // @[Modules.scala 160:64:@25356.4]
  wire [14:0] _T_78495; // @[Modules.scala 160:64:@25358.4]
  wire [13:0] _T_78496; // @[Modules.scala 160:64:@25359.4]
  wire [13:0] buffer_7_499; // @[Modules.scala 160:64:@25360.4]
  wire [14:0] _T_78498; // @[Modules.scala 160:64:@25362.4]
  wire [13:0] _T_78499; // @[Modules.scala 160:64:@25363.4]
  wire [13:0] buffer_7_500; // @[Modules.scala 160:64:@25364.4]
  wire [14:0] _T_78501; // @[Modules.scala 160:64:@25366.4]
  wire [13:0] _T_78502; // @[Modules.scala 160:64:@25367.4]
  wire [13:0] buffer_7_501; // @[Modules.scala 160:64:@25368.4]
  wire [14:0] _T_78504; // @[Modules.scala 160:64:@25370.4]
  wire [13:0] _T_78505; // @[Modules.scala 160:64:@25371.4]
  wire [13:0] buffer_7_502; // @[Modules.scala 160:64:@25372.4]
  wire [14:0] _T_78507; // @[Modules.scala 160:64:@25374.4]
  wire [13:0] _T_78508; // @[Modules.scala 160:64:@25375.4]
  wire [13:0] buffer_7_503; // @[Modules.scala 160:64:@25376.4]
  wire [14:0] _T_78510; // @[Modules.scala 160:64:@25378.4]
  wire [13:0] _T_78511; // @[Modules.scala 160:64:@25379.4]
  wire [13:0] buffer_7_504; // @[Modules.scala 160:64:@25380.4]
  wire [14:0] _T_78513; // @[Modules.scala 160:64:@25382.4]
  wire [13:0] _T_78514; // @[Modules.scala 160:64:@25383.4]
  wire [13:0] buffer_7_505; // @[Modules.scala 160:64:@25384.4]
  wire [14:0] _T_78516; // @[Modules.scala 160:64:@25386.4]
  wire [13:0] _T_78517; // @[Modules.scala 160:64:@25387.4]
  wire [13:0] buffer_7_506; // @[Modules.scala 160:64:@25388.4]
  wire [14:0] _T_78519; // @[Modules.scala 160:64:@25390.4]
  wire [13:0] _T_78520; // @[Modules.scala 160:64:@25391.4]
  wire [13:0] buffer_7_507; // @[Modules.scala 160:64:@25392.4]
  wire [14:0] _T_78522; // @[Modules.scala 160:64:@25394.4]
  wire [13:0] _T_78523; // @[Modules.scala 160:64:@25395.4]
  wire [13:0] buffer_7_508; // @[Modules.scala 160:64:@25396.4]
  wire [14:0] _T_78525; // @[Modules.scala 160:64:@25398.4]
  wire [13:0] _T_78526; // @[Modules.scala 160:64:@25399.4]
  wire [13:0] buffer_7_509; // @[Modules.scala 160:64:@25400.4]
  wire [14:0] _T_78528; // @[Modules.scala 160:64:@25402.4]
  wire [13:0] _T_78529; // @[Modules.scala 160:64:@25403.4]
  wire [13:0] buffer_7_510; // @[Modules.scala 160:64:@25404.4]
  wire [14:0] _T_78531; // @[Modules.scala 160:64:@25406.4]
  wire [13:0] _T_78532; // @[Modules.scala 160:64:@25407.4]
  wire [13:0] buffer_7_511; // @[Modules.scala 160:64:@25408.4]
  wire [14:0] _T_78534; // @[Modules.scala 160:64:@25410.4]
  wire [13:0] _T_78535; // @[Modules.scala 160:64:@25411.4]
  wire [13:0] buffer_7_512; // @[Modules.scala 160:64:@25412.4]
  wire [14:0] _T_78537; // @[Modules.scala 160:64:@25414.4]
  wire [13:0] _T_78538; // @[Modules.scala 160:64:@25415.4]
  wire [13:0] buffer_7_513; // @[Modules.scala 160:64:@25416.4]
  wire [14:0] _T_78540; // @[Modules.scala 160:64:@25418.4]
  wire [13:0] _T_78541; // @[Modules.scala 160:64:@25419.4]
  wire [13:0] buffer_7_514; // @[Modules.scala 160:64:@25420.4]
  wire [14:0] _T_78543; // @[Modules.scala 160:64:@25422.4]
  wire [13:0] _T_78544; // @[Modules.scala 160:64:@25423.4]
  wire [13:0] buffer_7_515; // @[Modules.scala 160:64:@25424.4]
  wire [14:0] _T_78546; // @[Modules.scala 160:64:@25426.4]
  wire [13:0] _T_78547; // @[Modules.scala 160:64:@25427.4]
  wire [13:0] buffer_7_516; // @[Modules.scala 160:64:@25428.4]
  wire [14:0] _T_78549; // @[Modules.scala 160:64:@25430.4]
  wire [13:0] _T_78550; // @[Modules.scala 160:64:@25431.4]
  wire [13:0] buffer_7_517; // @[Modules.scala 160:64:@25432.4]
  wire [14:0] _T_78552; // @[Modules.scala 160:64:@25434.4]
  wire [13:0] _T_78553; // @[Modules.scala 160:64:@25435.4]
  wire [13:0] buffer_7_518; // @[Modules.scala 160:64:@25436.4]
  wire [14:0] _T_78555; // @[Modules.scala 160:64:@25438.4]
  wire [13:0] _T_78556; // @[Modules.scala 160:64:@25439.4]
  wire [13:0] buffer_7_519; // @[Modules.scala 160:64:@25440.4]
  wire [14:0] _T_78558; // @[Modules.scala 160:64:@25442.4]
  wire [13:0] _T_78559; // @[Modules.scala 160:64:@25443.4]
  wire [13:0] buffer_7_520; // @[Modules.scala 160:64:@25444.4]
  wire [14:0] _T_78561; // @[Modules.scala 160:64:@25446.4]
  wire [13:0] _T_78562; // @[Modules.scala 160:64:@25447.4]
  wire [13:0] buffer_7_521; // @[Modules.scala 160:64:@25448.4]
  wire [14:0] _T_78564; // @[Modules.scala 160:64:@25450.4]
  wire [13:0] _T_78565; // @[Modules.scala 160:64:@25451.4]
  wire [13:0] buffer_7_522; // @[Modules.scala 160:64:@25452.4]
  wire [14:0] _T_78567; // @[Modules.scala 160:64:@25454.4]
  wire [13:0] _T_78568; // @[Modules.scala 160:64:@25455.4]
  wire [13:0] buffer_7_523; // @[Modules.scala 160:64:@25456.4]
  wire [14:0] _T_78570; // @[Modules.scala 160:64:@25458.4]
  wire [13:0] _T_78571; // @[Modules.scala 160:64:@25459.4]
  wire [13:0] buffer_7_524; // @[Modules.scala 160:64:@25460.4]
  wire [14:0] _T_78573; // @[Modules.scala 160:64:@25462.4]
  wire [13:0] _T_78574; // @[Modules.scala 160:64:@25463.4]
  wire [13:0] buffer_7_525; // @[Modules.scala 160:64:@25464.4]
  wire [14:0] _T_78576; // @[Modules.scala 160:64:@25466.4]
  wire [13:0] _T_78577; // @[Modules.scala 160:64:@25467.4]
  wire [13:0] buffer_7_526; // @[Modules.scala 160:64:@25468.4]
  wire [14:0] _T_78579; // @[Modules.scala 160:64:@25470.4]
  wire [13:0] _T_78580; // @[Modules.scala 160:64:@25471.4]
  wire [13:0] buffer_7_527; // @[Modules.scala 160:64:@25472.4]
  wire [14:0] _T_78582; // @[Modules.scala 160:64:@25474.4]
  wire [13:0] _T_78583; // @[Modules.scala 160:64:@25475.4]
  wire [13:0] buffer_7_528; // @[Modules.scala 160:64:@25476.4]
  wire [14:0] _T_78585; // @[Modules.scala 160:64:@25478.4]
  wire [13:0] _T_78586; // @[Modules.scala 160:64:@25479.4]
  wire [13:0] buffer_7_529; // @[Modules.scala 160:64:@25480.4]
  wire [14:0] _T_78588; // @[Modules.scala 160:64:@25482.4]
  wire [13:0] _T_78589; // @[Modules.scala 160:64:@25483.4]
  wire [13:0] buffer_7_530; // @[Modules.scala 160:64:@25484.4]
  wire [14:0] _T_78591; // @[Modules.scala 160:64:@25486.4]
  wire [13:0] _T_78592; // @[Modules.scala 160:64:@25487.4]
  wire [13:0] buffer_7_531; // @[Modules.scala 160:64:@25488.4]
  wire [14:0] _T_78594; // @[Modules.scala 160:64:@25490.4]
  wire [13:0] _T_78595; // @[Modules.scala 160:64:@25491.4]
  wire [13:0] buffer_7_532; // @[Modules.scala 160:64:@25492.4]
  wire [14:0] _T_78597; // @[Modules.scala 160:64:@25494.4]
  wire [13:0] _T_78598; // @[Modules.scala 160:64:@25495.4]
  wire [13:0] buffer_7_533; // @[Modules.scala 160:64:@25496.4]
  wire [14:0] _T_78600; // @[Modules.scala 160:64:@25498.4]
  wire [13:0] _T_78601; // @[Modules.scala 160:64:@25499.4]
  wire [13:0] buffer_7_534; // @[Modules.scala 160:64:@25500.4]
  wire [14:0] _T_78603; // @[Modules.scala 160:64:@25502.4]
  wire [13:0] _T_78604; // @[Modules.scala 160:64:@25503.4]
  wire [13:0] buffer_7_535; // @[Modules.scala 160:64:@25504.4]
  wire [14:0] _T_78606; // @[Modules.scala 160:64:@25506.4]
  wire [13:0] _T_78607; // @[Modules.scala 160:64:@25507.4]
  wire [13:0] buffer_7_536; // @[Modules.scala 160:64:@25508.4]
  wire [14:0] _T_78609; // @[Modules.scala 160:64:@25510.4]
  wire [13:0] _T_78610; // @[Modules.scala 160:64:@25511.4]
  wire [13:0] buffer_7_537; // @[Modules.scala 160:64:@25512.4]
  wire [14:0] _T_78612; // @[Modules.scala 160:64:@25514.4]
  wire [13:0] _T_78613; // @[Modules.scala 160:64:@25515.4]
  wire [13:0] buffer_7_538; // @[Modules.scala 160:64:@25516.4]
  wire [14:0] _T_78615; // @[Modules.scala 160:64:@25518.4]
  wire [13:0] _T_78616; // @[Modules.scala 160:64:@25519.4]
  wire [13:0] buffer_7_539; // @[Modules.scala 160:64:@25520.4]
  wire [14:0] _T_78618; // @[Modules.scala 166:64:@25522.4]
  wire [13:0] _T_78619; // @[Modules.scala 166:64:@25523.4]
  wire [13:0] buffer_7_540; // @[Modules.scala 166:64:@25524.4]
  wire [14:0] _T_78621; // @[Modules.scala 166:64:@25526.4]
  wire [13:0] _T_78622; // @[Modules.scala 166:64:@25527.4]
  wire [13:0] buffer_7_541; // @[Modules.scala 166:64:@25528.4]
  wire [14:0] _T_78624; // @[Modules.scala 166:64:@25530.4]
  wire [13:0] _T_78625; // @[Modules.scala 166:64:@25531.4]
  wire [13:0] buffer_7_542; // @[Modules.scala 166:64:@25532.4]
  wire [14:0] _T_78627; // @[Modules.scala 166:64:@25534.4]
  wire [13:0] _T_78628; // @[Modules.scala 166:64:@25535.4]
  wire [13:0] buffer_7_543; // @[Modules.scala 166:64:@25536.4]
  wire [14:0] _T_78630; // @[Modules.scala 166:64:@25538.4]
  wire [13:0] _T_78631; // @[Modules.scala 166:64:@25539.4]
  wire [13:0] buffer_7_544; // @[Modules.scala 166:64:@25540.4]
  wire [14:0] _T_78633; // @[Modules.scala 166:64:@25542.4]
  wire [13:0] _T_78634; // @[Modules.scala 166:64:@25543.4]
  wire [13:0] buffer_7_545; // @[Modules.scala 166:64:@25544.4]
  wire [14:0] _T_78636; // @[Modules.scala 166:64:@25546.4]
  wire [13:0] _T_78637; // @[Modules.scala 166:64:@25547.4]
  wire [13:0] buffer_7_546; // @[Modules.scala 166:64:@25548.4]
  wire [14:0] _T_78639; // @[Modules.scala 166:64:@25550.4]
  wire [13:0] _T_78640; // @[Modules.scala 166:64:@25551.4]
  wire [13:0] buffer_7_547; // @[Modules.scala 166:64:@25552.4]
  wire [14:0] _T_78642; // @[Modules.scala 166:64:@25554.4]
  wire [13:0] _T_78643; // @[Modules.scala 166:64:@25555.4]
  wire [13:0] buffer_7_548; // @[Modules.scala 166:64:@25556.4]
  wire [14:0] _T_78645; // @[Modules.scala 166:64:@25558.4]
  wire [13:0] _T_78646; // @[Modules.scala 166:64:@25559.4]
  wire [13:0] buffer_7_549; // @[Modules.scala 166:64:@25560.4]
  wire [14:0] _T_78648; // @[Modules.scala 166:64:@25562.4]
  wire [13:0] _T_78649; // @[Modules.scala 166:64:@25563.4]
  wire [13:0] buffer_7_550; // @[Modules.scala 166:64:@25564.4]
  wire [14:0] _T_78651; // @[Modules.scala 166:64:@25566.4]
  wire [13:0] _T_78652; // @[Modules.scala 166:64:@25567.4]
  wire [13:0] buffer_7_551; // @[Modules.scala 166:64:@25568.4]
  wire [14:0] _T_78654; // @[Modules.scala 166:64:@25570.4]
  wire [13:0] _T_78655; // @[Modules.scala 166:64:@25571.4]
  wire [13:0] buffer_7_552; // @[Modules.scala 166:64:@25572.4]
  wire [14:0] _T_78657; // @[Modules.scala 166:64:@25574.4]
  wire [13:0] _T_78658; // @[Modules.scala 166:64:@25575.4]
  wire [13:0] buffer_7_553; // @[Modules.scala 166:64:@25576.4]
  wire [14:0] _T_78660; // @[Modules.scala 166:64:@25578.4]
  wire [13:0] _T_78661; // @[Modules.scala 166:64:@25579.4]
  wire [13:0] buffer_7_554; // @[Modules.scala 166:64:@25580.4]
  wire [14:0] _T_78663; // @[Modules.scala 166:64:@25582.4]
  wire [13:0] _T_78664; // @[Modules.scala 166:64:@25583.4]
  wire [13:0] buffer_7_555; // @[Modules.scala 166:64:@25584.4]
  wire [14:0] _T_78666; // @[Modules.scala 166:64:@25586.4]
  wire [13:0] _T_78667; // @[Modules.scala 166:64:@25587.4]
  wire [13:0] buffer_7_556; // @[Modules.scala 166:64:@25588.4]
  wire [14:0] _T_78669; // @[Modules.scala 166:64:@25590.4]
  wire [13:0] _T_78670; // @[Modules.scala 166:64:@25591.4]
  wire [13:0] buffer_7_557; // @[Modules.scala 166:64:@25592.4]
  wire [14:0] _T_78672; // @[Modules.scala 166:64:@25594.4]
  wire [13:0] _T_78673; // @[Modules.scala 166:64:@25595.4]
  wire [13:0] buffer_7_558; // @[Modules.scala 166:64:@25596.4]
  wire [14:0] _T_78675; // @[Modules.scala 166:64:@25598.4]
  wire [13:0] _T_78676; // @[Modules.scala 166:64:@25599.4]
  wire [13:0] buffer_7_559; // @[Modules.scala 166:64:@25600.4]
  wire [14:0] _T_78678; // @[Modules.scala 166:64:@25602.4]
  wire [13:0] _T_78679; // @[Modules.scala 166:64:@25603.4]
  wire [13:0] buffer_7_560; // @[Modules.scala 166:64:@25604.4]
  wire [14:0] _T_78681; // @[Modules.scala 166:64:@25606.4]
  wire [13:0] _T_78682; // @[Modules.scala 166:64:@25607.4]
  wire [13:0] buffer_7_561; // @[Modules.scala 166:64:@25608.4]
  wire [14:0] _T_78684; // @[Modules.scala 166:64:@25610.4]
  wire [13:0] _T_78685; // @[Modules.scala 166:64:@25611.4]
  wire [13:0] buffer_7_562; // @[Modules.scala 166:64:@25612.4]
  wire [14:0] _T_78687; // @[Modules.scala 166:64:@25614.4]
  wire [13:0] _T_78688; // @[Modules.scala 166:64:@25615.4]
  wire [13:0] buffer_7_563; // @[Modules.scala 166:64:@25616.4]
  wire [14:0] _T_78690; // @[Modules.scala 166:64:@25618.4]
  wire [13:0] _T_78691; // @[Modules.scala 166:64:@25619.4]
  wire [13:0] buffer_7_564; // @[Modules.scala 166:64:@25620.4]
  wire [14:0] _T_78693; // @[Modules.scala 166:64:@25622.4]
  wire [13:0] _T_78694; // @[Modules.scala 166:64:@25623.4]
  wire [13:0] buffer_7_565; // @[Modules.scala 166:64:@25624.4]
  wire [14:0] _T_78696; // @[Modules.scala 166:64:@25626.4]
  wire [13:0] _T_78697; // @[Modules.scala 166:64:@25627.4]
  wire [13:0] buffer_7_566; // @[Modules.scala 166:64:@25628.4]
  wire [14:0] _T_78699; // @[Modules.scala 166:64:@25630.4]
  wire [13:0] _T_78700; // @[Modules.scala 166:64:@25631.4]
  wire [13:0] buffer_7_567; // @[Modules.scala 166:64:@25632.4]
  wire [14:0] _T_78702; // @[Modules.scala 166:64:@25634.4]
  wire [13:0] _T_78703; // @[Modules.scala 166:64:@25635.4]
  wire [13:0] buffer_7_568; // @[Modules.scala 166:64:@25636.4]
  wire [14:0] _T_78705; // @[Modules.scala 166:64:@25638.4]
  wire [13:0] _T_78706; // @[Modules.scala 166:64:@25639.4]
  wire [13:0] buffer_7_569; // @[Modules.scala 166:64:@25640.4]
  wire [14:0] _T_78708; // @[Modules.scala 166:64:@25642.4]
  wire [13:0] _T_78709; // @[Modules.scala 166:64:@25643.4]
  wire [13:0] buffer_7_570; // @[Modules.scala 166:64:@25644.4]
  wire [14:0] _T_78711; // @[Modules.scala 166:64:@25646.4]
  wire [13:0] _T_78712; // @[Modules.scala 166:64:@25647.4]
  wire [13:0] buffer_7_571; // @[Modules.scala 166:64:@25648.4]
  wire [14:0] _T_78714; // @[Modules.scala 166:64:@25650.4]
  wire [13:0] _T_78715; // @[Modules.scala 166:64:@25651.4]
  wire [13:0] buffer_7_572; // @[Modules.scala 166:64:@25652.4]
  wire [14:0] _T_78717; // @[Modules.scala 166:64:@25654.4]
  wire [13:0] _T_78718; // @[Modules.scala 166:64:@25655.4]
  wire [13:0] buffer_7_573; // @[Modules.scala 166:64:@25656.4]
  wire [14:0] _T_78720; // @[Modules.scala 166:64:@25658.4]
  wire [13:0] _T_78721; // @[Modules.scala 166:64:@25659.4]
  wire [13:0] buffer_7_574; // @[Modules.scala 166:64:@25660.4]
  wire [14:0] _T_78723; // @[Modules.scala 166:64:@25662.4]
  wire [13:0] _T_78724; // @[Modules.scala 166:64:@25663.4]
  wire [13:0] buffer_7_575; // @[Modules.scala 166:64:@25664.4]
  wire [14:0] _T_78726; // @[Modules.scala 166:64:@25666.4]
  wire [13:0] _T_78727; // @[Modules.scala 166:64:@25667.4]
  wire [13:0] buffer_7_576; // @[Modules.scala 166:64:@25668.4]
  wire [14:0] _T_78729; // @[Modules.scala 166:64:@25670.4]
  wire [13:0] _T_78730; // @[Modules.scala 166:64:@25671.4]
  wire [13:0] buffer_7_577; // @[Modules.scala 166:64:@25672.4]
  wire [13:0] buffer_7_308; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_78732; // @[Modules.scala 172:66:@25674.4]
  wire [13:0] _T_78733; // @[Modules.scala 172:66:@25675.4]
  wire [13:0] buffer_7_578; // @[Modules.scala 172:66:@25676.4]
  wire [14:0] _T_78735; // @[Modules.scala 166:64:@25678.4]
  wire [13:0] _T_78736; // @[Modules.scala 166:64:@25679.4]
  wire [13:0] buffer_7_579; // @[Modules.scala 166:64:@25680.4]
  wire [14:0] _T_78738; // @[Modules.scala 166:64:@25682.4]
  wire [13:0] _T_78739; // @[Modules.scala 166:64:@25683.4]
  wire [13:0] buffer_7_580; // @[Modules.scala 166:64:@25684.4]
  wire [14:0] _T_78741; // @[Modules.scala 166:64:@25686.4]
  wire [13:0] _T_78742; // @[Modules.scala 166:64:@25687.4]
  wire [13:0] buffer_7_581; // @[Modules.scala 166:64:@25688.4]
  wire [14:0] _T_78744; // @[Modules.scala 166:64:@25690.4]
  wire [13:0] _T_78745; // @[Modules.scala 166:64:@25691.4]
  wire [13:0] buffer_7_582; // @[Modules.scala 166:64:@25692.4]
  wire [14:0] _T_78747; // @[Modules.scala 166:64:@25694.4]
  wire [13:0] _T_78748; // @[Modules.scala 166:64:@25695.4]
  wire [13:0] buffer_7_583; // @[Modules.scala 166:64:@25696.4]
  wire [14:0] _T_78750; // @[Modules.scala 166:64:@25698.4]
  wire [13:0] _T_78751; // @[Modules.scala 166:64:@25699.4]
  wire [13:0] buffer_7_584; // @[Modules.scala 166:64:@25700.4]
  wire [14:0] _T_78753; // @[Modules.scala 166:64:@25702.4]
  wire [13:0] _T_78754; // @[Modules.scala 166:64:@25703.4]
  wire [13:0] buffer_7_585; // @[Modules.scala 166:64:@25704.4]
  wire [14:0] _T_78756; // @[Modules.scala 166:64:@25706.4]
  wire [13:0] _T_78757; // @[Modules.scala 166:64:@25707.4]
  wire [13:0] buffer_7_586; // @[Modules.scala 166:64:@25708.4]
  wire [14:0] _T_78759; // @[Modules.scala 166:64:@25710.4]
  wire [13:0] _T_78760; // @[Modules.scala 166:64:@25711.4]
  wire [13:0] buffer_7_587; // @[Modules.scala 166:64:@25712.4]
  wire [14:0] _T_78762; // @[Modules.scala 166:64:@25714.4]
  wire [13:0] _T_78763; // @[Modules.scala 166:64:@25715.4]
  wire [13:0] buffer_7_588; // @[Modules.scala 166:64:@25716.4]
  wire [14:0] _T_78765; // @[Modules.scala 166:64:@25718.4]
  wire [13:0] _T_78766; // @[Modules.scala 166:64:@25719.4]
  wire [13:0] buffer_7_589; // @[Modules.scala 166:64:@25720.4]
  wire [14:0] _T_78768; // @[Modules.scala 166:64:@25722.4]
  wire [13:0] _T_78769; // @[Modules.scala 166:64:@25723.4]
  wire [13:0] buffer_7_590; // @[Modules.scala 166:64:@25724.4]
  wire [14:0] _T_78771; // @[Modules.scala 166:64:@25726.4]
  wire [13:0] _T_78772; // @[Modules.scala 166:64:@25727.4]
  wire [13:0] buffer_7_591; // @[Modules.scala 166:64:@25728.4]
  wire [14:0] _T_78774; // @[Modules.scala 166:64:@25730.4]
  wire [13:0] _T_78775; // @[Modules.scala 166:64:@25731.4]
  wire [13:0] buffer_7_592; // @[Modules.scala 166:64:@25732.4]
  wire [14:0] _T_78777; // @[Modules.scala 166:64:@25734.4]
  wire [13:0] _T_78778; // @[Modules.scala 166:64:@25735.4]
  wire [13:0] buffer_7_593; // @[Modules.scala 166:64:@25736.4]
  wire [14:0] _T_78780; // @[Modules.scala 166:64:@25738.4]
  wire [13:0] _T_78781; // @[Modules.scala 166:64:@25739.4]
  wire [13:0] buffer_7_594; // @[Modules.scala 166:64:@25740.4]
  wire [14:0] _T_78783; // @[Modules.scala 166:64:@25742.4]
  wire [13:0] _T_78784; // @[Modules.scala 166:64:@25743.4]
  wire [13:0] buffer_7_595; // @[Modules.scala 166:64:@25744.4]
  wire [14:0] _T_78786; // @[Modules.scala 166:64:@25746.4]
  wire [13:0] _T_78787; // @[Modules.scala 166:64:@25747.4]
  wire [13:0] buffer_7_596; // @[Modules.scala 166:64:@25748.4]
  wire [14:0] _T_78789; // @[Modules.scala 166:64:@25750.4]
  wire [13:0] _T_78790; // @[Modules.scala 166:64:@25751.4]
  wire [13:0] buffer_7_597; // @[Modules.scala 166:64:@25752.4]
  wire [14:0] _T_78792; // @[Modules.scala 166:64:@25754.4]
  wire [13:0] _T_78793; // @[Modules.scala 166:64:@25755.4]
  wire [13:0] buffer_7_598; // @[Modules.scala 166:64:@25756.4]
  wire [14:0] _T_78795; // @[Modules.scala 166:64:@25758.4]
  wire [13:0] _T_78796; // @[Modules.scala 166:64:@25759.4]
  wire [13:0] buffer_7_599; // @[Modules.scala 166:64:@25760.4]
  wire [14:0] _T_78798; // @[Modules.scala 166:64:@25762.4]
  wire [13:0] _T_78799; // @[Modules.scala 166:64:@25763.4]
  wire [13:0] buffer_7_600; // @[Modules.scala 166:64:@25764.4]
  wire [14:0] _T_78801; // @[Modules.scala 166:64:@25766.4]
  wire [13:0] _T_78802; // @[Modules.scala 166:64:@25767.4]
  wire [13:0] buffer_7_601; // @[Modules.scala 166:64:@25768.4]
  wire [14:0] _T_78804; // @[Modules.scala 166:64:@25770.4]
  wire [13:0] _T_78805; // @[Modules.scala 166:64:@25771.4]
  wire [13:0] buffer_7_602; // @[Modules.scala 166:64:@25772.4]
  wire [14:0] _T_78807; // @[Modules.scala 166:64:@25774.4]
  wire [13:0] _T_78808; // @[Modules.scala 166:64:@25775.4]
  wire [13:0] buffer_7_603; // @[Modules.scala 166:64:@25776.4]
  wire [14:0] _T_78810; // @[Modules.scala 166:64:@25778.4]
  wire [13:0] _T_78811; // @[Modules.scala 166:64:@25779.4]
  wire [13:0] buffer_7_604; // @[Modules.scala 166:64:@25780.4]
  wire [14:0] _T_78813; // @[Modules.scala 166:64:@25782.4]
  wire [13:0] _T_78814; // @[Modules.scala 166:64:@25783.4]
  wire [13:0] buffer_7_605; // @[Modules.scala 166:64:@25784.4]
  wire [14:0] _T_78816; // @[Modules.scala 166:64:@25786.4]
  wire [13:0] _T_78817; // @[Modules.scala 166:64:@25787.4]
  wire [13:0] buffer_7_606; // @[Modules.scala 166:64:@25788.4]
  wire [14:0] _T_78819; // @[Modules.scala 172:66:@25790.4]
  wire [13:0] _T_78820; // @[Modules.scala 172:66:@25791.4]
  wire [13:0] buffer_7_607; // @[Modules.scala 172:66:@25792.4]
  wire [14:0] _T_78822; // @[Modules.scala 160:64:@25794.4]
  wire [13:0] _T_78823; // @[Modules.scala 160:64:@25795.4]
  wire [13:0] buffer_7_608; // @[Modules.scala 160:64:@25796.4]
  wire [14:0] _T_78825; // @[Modules.scala 160:64:@25798.4]
  wire [13:0] _T_78826; // @[Modules.scala 160:64:@25799.4]
  wire [13:0] buffer_7_609; // @[Modules.scala 160:64:@25800.4]
  wire [14:0] _T_78828; // @[Modules.scala 160:64:@25802.4]
  wire [13:0] _T_78829; // @[Modules.scala 160:64:@25803.4]
  wire [13:0] buffer_7_610; // @[Modules.scala 160:64:@25804.4]
  wire [14:0] _T_78831; // @[Modules.scala 160:64:@25806.4]
  wire [13:0] _T_78832; // @[Modules.scala 160:64:@25807.4]
  wire [13:0] buffer_7_611; // @[Modules.scala 160:64:@25808.4]
  wire [14:0] _T_78834; // @[Modules.scala 160:64:@25810.4]
  wire [13:0] _T_78835; // @[Modules.scala 160:64:@25811.4]
  wire [13:0] buffer_7_612; // @[Modules.scala 160:64:@25812.4]
  wire [14:0] _T_78837; // @[Modules.scala 166:64:@25814.4]
  wire [13:0] _T_78838; // @[Modules.scala 166:64:@25815.4]
  wire [13:0] buffer_7_613; // @[Modules.scala 166:64:@25816.4]
  wire [14:0] _T_78840; // @[Modules.scala 166:64:@25818.4]
  wire [13:0] _T_78841; // @[Modules.scala 166:64:@25819.4]
  wire [13:0] buffer_7_614; // @[Modules.scala 166:64:@25820.4]
  wire [14:0] _T_78843; // @[Modules.scala 160:64:@25822.4]
  wire [13:0] _T_78844; // @[Modules.scala 160:64:@25823.4]
  wire [13:0] buffer_7_615; // @[Modules.scala 160:64:@25824.4]
  wire [14:0] _T_78846; // @[Modules.scala 172:66:@25826.4]
  wire [13:0] _T_78847; // @[Modules.scala 172:66:@25827.4]
  wire [13:0] buffer_7_616; // @[Modules.scala 172:66:@25828.4]
  wire [5:0] _T_78864; // @[Modules.scala 143:74:@26009.4]
  wire [5:0] _T_78866; // @[Modules.scala 144:80:@26010.4]
  wire [6:0] _T_78867; // @[Modules.scala 143:103:@26011.4]
  wire [5:0] _T_78868; // @[Modules.scala 143:103:@26012.4]
  wire [5:0] _T_78869; // @[Modules.scala 143:103:@26013.4]
  wire [5:0] _GEN_566; // @[Modules.scala 143:103:@26029.4]
  wire [6:0] _T_78888; // @[Modules.scala 143:103:@26029.4]
  wire [5:0] _T_78889; // @[Modules.scala 143:103:@26030.4]
  wire [5:0] _T_78890; // @[Modules.scala 143:103:@26031.4]
  wire [5:0] _T_78909; // @[Modules.scala 143:103:@26047.4]
  wire [4:0] _T_78910; // @[Modules.scala 143:103:@26048.4]
  wire [4:0] _T_78911; // @[Modules.scala 143:103:@26049.4]
  wire [5:0] _GEN_568; // @[Modules.scala 143:103:@26071.4]
  wire [6:0] _T_78937; // @[Modules.scala 143:103:@26071.4]
  wire [5:0] _T_78938; // @[Modules.scala 143:103:@26072.4]
  wire [5:0] _T_78939; // @[Modules.scala 143:103:@26073.4]
  wire [5:0] _GEN_570; // @[Modules.scala 143:103:@26131.4]
  wire [6:0] _T_79007; // @[Modules.scala 143:103:@26131.4]
  wire [5:0] _T_79008; // @[Modules.scala 143:103:@26132.4]
  wire [5:0] _T_79009; // @[Modules.scala 143:103:@26133.4]
  wire [5:0] _GEN_571; // @[Modules.scala 143:103:@26143.4]
  wire [6:0] _T_79021; // @[Modules.scala 143:103:@26143.4]
  wire [5:0] _T_79022; // @[Modules.scala 143:103:@26144.4]
  wire [5:0] _T_79023; // @[Modules.scala 143:103:@26145.4]
  wire [5:0] _T_79091; // @[Modules.scala 143:103:@26203.4]
  wire [4:0] _T_79092; // @[Modules.scala 143:103:@26204.4]
  wire [4:0] _T_79093; // @[Modules.scala 143:103:@26205.4]
  wire [6:0] _T_79098; // @[Modules.scala 143:103:@26209.4]
  wire [5:0] _T_79099; // @[Modules.scala 143:103:@26210.4]
  wire [5:0] _T_79100; // @[Modules.scala 143:103:@26211.4]
  wire [6:0] _T_79105; // @[Modules.scala 143:103:@26215.4]
  wire [5:0] _T_79106; // @[Modules.scala 143:103:@26216.4]
  wire [5:0] _T_79107; // @[Modules.scala 143:103:@26217.4]
  wire [5:0] _GEN_575; // @[Modules.scala 143:103:@26239.4]
  wire [6:0] _T_79133; // @[Modules.scala 143:103:@26239.4]
  wire [5:0] _T_79134; // @[Modules.scala 143:103:@26240.4]
  wire [5:0] _T_79135; // @[Modules.scala 143:103:@26241.4]
  wire [6:0] _T_79140; // @[Modules.scala 143:103:@26245.4]
  wire [5:0] _T_79141; // @[Modules.scala 143:103:@26246.4]
  wire [5:0] _T_79142; // @[Modules.scala 143:103:@26247.4]
  wire [5:0] _GEN_578; // @[Modules.scala 143:103:@26275.4]
  wire [6:0] _T_79175; // @[Modules.scala 143:103:@26275.4]
  wire [5:0] _T_79176; // @[Modules.scala 143:103:@26276.4]
  wire [5:0] _T_79177; // @[Modules.scala 143:103:@26277.4]
  wire [5:0] _GEN_579; // @[Modules.scala 143:103:@26281.4]
  wire [6:0] _T_79182; // @[Modules.scala 143:103:@26281.4]
  wire [5:0] _T_79183; // @[Modules.scala 143:103:@26282.4]
  wire [5:0] _T_79184; // @[Modules.scala 143:103:@26283.4]
  wire [6:0] _T_79189; // @[Modules.scala 143:103:@26287.4]
  wire [5:0] _T_79190; // @[Modules.scala 143:103:@26288.4]
  wire [5:0] _T_79191; // @[Modules.scala 143:103:@26289.4]
  wire [6:0] _T_79196; // @[Modules.scala 143:103:@26293.4]
  wire [5:0] _T_79197; // @[Modules.scala 143:103:@26294.4]
  wire [5:0] _T_79198; // @[Modules.scala 143:103:@26295.4]
  wire [5:0] _T_79238; // @[Modules.scala 143:103:@26329.4]
  wire [4:0] _T_79239; // @[Modules.scala 143:103:@26330.4]
  wire [4:0] _T_79240; // @[Modules.scala 143:103:@26331.4]
  wire [6:0] _T_79245; // @[Modules.scala 143:103:@26335.4]
  wire [5:0] _T_79246; // @[Modules.scala 143:103:@26336.4]
  wire [5:0] _T_79247; // @[Modules.scala 143:103:@26337.4]
  wire [6:0] _T_79266; // @[Modules.scala 143:103:@26353.4]
  wire [5:0] _T_79267; // @[Modules.scala 143:103:@26354.4]
  wire [5:0] _T_79268; // @[Modules.scala 143:103:@26355.4]
  wire [6:0] _T_79273; // @[Modules.scala 143:103:@26359.4]
  wire [5:0] _T_79274; // @[Modules.scala 143:103:@26360.4]
  wire [5:0] _T_79275; // @[Modules.scala 143:103:@26361.4]
  wire [6:0] _T_79280; // @[Modules.scala 143:103:@26365.4]
  wire [5:0] _T_79281; // @[Modules.scala 143:103:@26366.4]
  wire [5:0] _T_79282; // @[Modules.scala 143:103:@26367.4]
  wire [6:0] _T_79287; // @[Modules.scala 143:103:@26371.4]
  wire [5:0] _T_79288; // @[Modules.scala 143:103:@26372.4]
  wire [5:0] _T_79289; // @[Modules.scala 143:103:@26373.4]
  wire [6:0] _T_79294; // @[Modules.scala 143:103:@26377.4]
  wire [5:0] _T_79295; // @[Modules.scala 143:103:@26378.4]
  wire [5:0] _T_79296; // @[Modules.scala 143:103:@26379.4]
  wire [6:0] _T_79301; // @[Modules.scala 143:103:@26383.4]
  wire [5:0] _T_79302; // @[Modules.scala 143:103:@26384.4]
  wire [5:0] _T_79303; // @[Modules.scala 143:103:@26385.4]
  wire [5:0] _GEN_587; // @[Modules.scala 143:103:@26395.4]
  wire [6:0] _T_79315; // @[Modules.scala 143:103:@26395.4]
  wire [5:0] _T_79316; // @[Modules.scala 143:103:@26396.4]
  wire [5:0] _T_79317; // @[Modules.scala 143:103:@26397.4]
  wire [5:0] _GEN_588; // @[Modules.scala 143:103:@26401.4]
  wire [6:0] _T_79322; // @[Modules.scala 143:103:@26401.4]
  wire [5:0] _T_79323; // @[Modules.scala 143:103:@26402.4]
  wire [5:0] _T_79324; // @[Modules.scala 143:103:@26403.4]
  wire [5:0] _GEN_589; // @[Modules.scala 143:103:@26413.4]
  wire [6:0] _T_79336; // @[Modules.scala 143:103:@26413.4]
  wire [5:0] _T_79337; // @[Modules.scala 143:103:@26414.4]
  wire [5:0] _T_79338; // @[Modules.scala 143:103:@26415.4]
  wire [6:0] _T_79343; // @[Modules.scala 143:103:@26419.4]
  wire [5:0] _T_79344; // @[Modules.scala 143:103:@26420.4]
  wire [5:0] _T_79345; // @[Modules.scala 143:103:@26421.4]
  wire [6:0] _T_79350; // @[Modules.scala 143:103:@26425.4]
  wire [5:0] _T_79351; // @[Modules.scala 143:103:@26426.4]
  wire [5:0] _T_79352; // @[Modules.scala 143:103:@26427.4]
  wire [5:0] _T_79371; // @[Modules.scala 143:103:@26443.4]
  wire [4:0] _T_79372; // @[Modules.scala 143:103:@26444.4]
  wire [4:0] _T_79373; // @[Modules.scala 143:103:@26445.4]
  wire [5:0] _GEN_590; // @[Modules.scala 143:103:@26455.4]
  wire [6:0] _T_79385; // @[Modules.scala 143:103:@26455.4]
  wire [5:0] _T_79386; // @[Modules.scala 143:103:@26456.4]
  wire [5:0] _T_79387; // @[Modules.scala 143:103:@26457.4]
  wire [6:0] _T_79392; // @[Modules.scala 143:103:@26461.4]
  wire [5:0] _T_79393; // @[Modules.scala 143:103:@26462.4]
  wire [5:0] _T_79394; // @[Modules.scala 143:103:@26463.4]
  wire [6:0] _T_79399; // @[Modules.scala 143:103:@26467.4]
  wire [5:0] _T_79400; // @[Modules.scala 143:103:@26468.4]
  wire [5:0] _T_79401; // @[Modules.scala 143:103:@26469.4]
  wire [6:0] _T_79406; // @[Modules.scala 143:103:@26473.4]
  wire [5:0] _T_79407; // @[Modules.scala 143:103:@26474.4]
  wire [5:0] _T_79408; // @[Modules.scala 143:103:@26475.4]
  wire [5:0] _T_79413; // @[Modules.scala 143:103:@26479.4]
  wire [4:0] _T_79414; // @[Modules.scala 143:103:@26480.4]
  wire [4:0] _T_79415; // @[Modules.scala 143:103:@26481.4]
  wire [6:0] _T_79420; // @[Modules.scala 143:103:@26485.4]
  wire [5:0] _T_79421; // @[Modules.scala 143:103:@26486.4]
  wire [5:0] _T_79422; // @[Modules.scala 143:103:@26487.4]
  wire [5:0] _GEN_592; // @[Modules.scala 143:103:@26491.4]
  wire [6:0] _T_79427; // @[Modules.scala 143:103:@26491.4]
  wire [5:0] _T_79428; // @[Modules.scala 143:103:@26492.4]
  wire [5:0] _T_79429; // @[Modules.scala 143:103:@26493.4]
  wire [6:0] _T_79448; // @[Modules.scala 143:103:@26509.4]
  wire [5:0] _T_79449; // @[Modules.scala 143:103:@26510.4]
  wire [5:0] _T_79450; // @[Modules.scala 143:103:@26511.4]
  wire [5:0] _T_79455; // @[Modules.scala 143:103:@26515.4]
  wire [4:0] _T_79456; // @[Modules.scala 143:103:@26516.4]
  wire [4:0] _T_79457; // @[Modules.scala 143:103:@26517.4]
  wire [5:0] _GEN_593; // @[Modules.scala 143:103:@26521.4]
  wire [6:0] _T_79462; // @[Modules.scala 143:103:@26521.4]
  wire [5:0] _T_79463; // @[Modules.scala 143:103:@26522.4]
  wire [5:0] _T_79464; // @[Modules.scala 143:103:@26523.4]
  wire [6:0] _T_79476; // @[Modules.scala 143:103:@26533.4]
  wire [5:0] _T_79477; // @[Modules.scala 143:103:@26534.4]
  wire [5:0] _T_79478; // @[Modules.scala 143:103:@26535.4]
  wire [6:0] _T_79497; // @[Modules.scala 143:103:@26551.4]
  wire [5:0] _T_79498; // @[Modules.scala 143:103:@26552.4]
  wire [5:0] _T_79499; // @[Modules.scala 143:103:@26553.4]
  wire [5:0] _GEN_595; // @[Modules.scala 143:103:@26563.4]
  wire [6:0] _T_79511; // @[Modules.scala 143:103:@26563.4]
  wire [5:0] _T_79512; // @[Modules.scala 143:103:@26564.4]
  wire [5:0] _T_79513; // @[Modules.scala 143:103:@26565.4]
  wire [6:0] _T_79518; // @[Modules.scala 143:103:@26569.4]
  wire [5:0] _T_79519; // @[Modules.scala 143:103:@26570.4]
  wire [5:0] _T_79520; // @[Modules.scala 143:103:@26571.4]
  wire [5:0] _GEN_596; // @[Modules.scala 143:103:@26599.4]
  wire [6:0] _T_79553; // @[Modules.scala 143:103:@26599.4]
  wire [5:0] _T_79554; // @[Modules.scala 143:103:@26600.4]
  wire [5:0] _T_79555; // @[Modules.scala 143:103:@26601.4]
  wire [6:0] _T_79560; // @[Modules.scala 143:103:@26605.4]
  wire [5:0] _T_79561; // @[Modules.scala 143:103:@26606.4]
  wire [5:0] _T_79562; // @[Modules.scala 143:103:@26607.4]
  wire [6:0] _T_79602; // @[Modules.scala 143:103:@26641.4]
  wire [5:0] _T_79603; // @[Modules.scala 143:103:@26642.4]
  wire [5:0] _T_79604; // @[Modules.scala 143:103:@26643.4]
  wire [5:0] _T_79609; // @[Modules.scala 143:103:@26647.4]
  wire [4:0] _T_79610; // @[Modules.scala 143:103:@26648.4]
  wire [4:0] _T_79611; // @[Modules.scala 143:103:@26649.4]
  wire [6:0] _T_79623; // @[Modules.scala 143:103:@26659.4]
  wire [5:0] _T_79624; // @[Modules.scala 143:103:@26660.4]
  wire [5:0] _T_79625; // @[Modules.scala 143:103:@26661.4]
  wire [6:0] _T_79630; // @[Modules.scala 143:103:@26665.4]
  wire [5:0] _T_79631; // @[Modules.scala 143:103:@26666.4]
  wire [5:0] _T_79632; // @[Modules.scala 143:103:@26667.4]
  wire [5:0] _GEN_598; // @[Modules.scala 143:103:@26671.4]
  wire [6:0] _T_79637; // @[Modules.scala 143:103:@26671.4]
  wire [5:0] _T_79638; // @[Modules.scala 143:103:@26672.4]
  wire [5:0] _T_79639; // @[Modules.scala 143:103:@26673.4]
  wire [6:0] _T_79721; // @[Modules.scala 143:103:@26743.4]
  wire [5:0] _T_79722; // @[Modules.scala 143:103:@26744.4]
  wire [5:0] _T_79723; // @[Modules.scala 143:103:@26745.4]
  wire [5:0] _T_79784; // @[Modules.scala 143:103:@26797.4]
  wire [4:0] _T_79785; // @[Modules.scala 143:103:@26798.4]
  wire [4:0] _T_79786; // @[Modules.scala 143:103:@26799.4]
  wire [6:0] _T_79896; // @[Modules.scala 143:103:@26893.4]
  wire [5:0] _T_79897; // @[Modules.scala 143:103:@26894.4]
  wire [5:0] _T_79898; // @[Modules.scala 143:103:@26895.4]
  wire [6:0] _T_79903; // @[Modules.scala 143:103:@26899.4]
  wire [5:0] _T_79904; // @[Modules.scala 143:103:@26900.4]
  wire [5:0] _T_79905; // @[Modules.scala 143:103:@26901.4]
  wire [6:0] _T_79924; // @[Modules.scala 143:103:@26917.4]
  wire [5:0] _T_79925; // @[Modules.scala 143:103:@26918.4]
  wire [5:0] _T_79926; // @[Modules.scala 143:103:@26919.4]
  wire [6:0] _T_79938; // @[Modules.scala 143:103:@26929.4]
  wire [5:0] _T_79939; // @[Modules.scala 143:103:@26930.4]
  wire [5:0] _T_79940; // @[Modules.scala 143:103:@26931.4]
  wire [6:0] _T_79945; // @[Modules.scala 143:103:@26935.4]
  wire [5:0] _T_79946; // @[Modules.scala 143:103:@26936.4]
  wire [5:0] _T_79947; // @[Modules.scala 143:103:@26937.4]
  wire [6:0] _T_79952; // @[Modules.scala 143:103:@26941.4]
  wire [5:0] _T_79953; // @[Modules.scala 143:103:@26942.4]
  wire [5:0] _T_79954; // @[Modules.scala 143:103:@26943.4]
  wire [5:0] _T_79966; // @[Modules.scala 143:103:@26953.4]
  wire [4:0] _T_79967; // @[Modules.scala 143:103:@26954.4]
  wire [4:0] _T_79968; // @[Modules.scala 143:103:@26955.4]
  wire [6:0] _T_79973; // @[Modules.scala 143:103:@26959.4]
  wire [5:0] _T_79974; // @[Modules.scala 143:103:@26960.4]
  wire [5:0] _T_79975; // @[Modules.scala 143:103:@26961.4]
  wire [5:0] _GEN_607; // @[Modules.scala 143:103:@26989.4]
  wire [6:0] _T_80008; // @[Modules.scala 143:103:@26989.4]
  wire [5:0] _T_80009; // @[Modules.scala 143:103:@26990.4]
  wire [5:0] _T_80010; // @[Modules.scala 143:103:@26991.4]
  wire [6:0] _T_80022; // @[Modules.scala 143:103:@27001.4]
  wire [5:0] _T_80023; // @[Modules.scala 143:103:@27002.4]
  wire [5:0] _T_80024; // @[Modules.scala 143:103:@27003.4]
  wire [5:0] _T_80050; // @[Modules.scala 143:103:@27025.4]
  wire [4:0] _T_80051; // @[Modules.scala 143:103:@27026.4]
  wire [4:0] _T_80052; // @[Modules.scala 143:103:@27027.4]
  wire [6:0] _T_80064; // @[Modules.scala 143:103:@27037.4]
  wire [5:0] _T_80065; // @[Modules.scala 143:103:@27038.4]
  wire [5:0] _T_80066; // @[Modules.scala 143:103:@27039.4]
  wire [5:0] _T_80085; // @[Modules.scala 143:103:@27055.4]
  wire [4:0] _T_80086; // @[Modules.scala 143:103:@27056.4]
  wire [4:0] _T_80087; // @[Modules.scala 143:103:@27057.4]
  wire [5:0] _T_80092; // @[Modules.scala 143:103:@27061.4]
  wire [4:0] _T_80093; // @[Modules.scala 143:103:@27062.4]
  wire [4:0] _T_80094; // @[Modules.scala 143:103:@27063.4]
  wire [6:0] _T_80113; // @[Modules.scala 143:103:@27079.4]
  wire [5:0] _T_80114; // @[Modules.scala 143:103:@27080.4]
  wire [5:0] _T_80115; // @[Modules.scala 143:103:@27081.4]
  wire [6:0] _T_80120; // @[Modules.scala 143:103:@27085.4]
  wire [5:0] _T_80121; // @[Modules.scala 143:103:@27086.4]
  wire [5:0] _T_80122; // @[Modules.scala 143:103:@27087.4]
  wire [5:0] _T_80169; // @[Modules.scala 143:103:@27127.4]
  wire [4:0] _T_80170; // @[Modules.scala 143:103:@27128.4]
  wire [4:0] _T_80171; // @[Modules.scala 143:103:@27129.4]
  wire [5:0] _T_80176; // @[Modules.scala 143:103:@27133.4]
  wire [4:0] _T_80177; // @[Modules.scala 143:103:@27134.4]
  wire [4:0] _T_80178; // @[Modules.scala 143:103:@27135.4]
  wire [5:0] _T_80183; // @[Modules.scala 143:103:@27139.4]
  wire [4:0] _T_80184; // @[Modules.scala 143:103:@27140.4]
  wire [4:0] _T_80185; // @[Modules.scala 143:103:@27141.4]
  wire [5:0] _GEN_610; // @[Modules.scala 143:103:@27145.4]
  wire [6:0] _T_80190; // @[Modules.scala 143:103:@27145.4]
  wire [5:0] _T_80191; // @[Modules.scala 143:103:@27146.4]
  wire [5:0] _T_80192; // @[Modules.scala 143:103:@27147.4]
  wire [5:0] _T_80232; // @[Modules.scala 143:103:@27181.4]
  wire [4:0] _T_80233; // @[Modules.scala 143:103:@27182.4]
  wire [4:0] _T_80234; // @[Modules.scala 143:103:@27183.4]
  wire [6:0] _T_80239; // @[Modules.scala 143:103:@27187.4]
  wire [5:0] _T_80240; // @[Modules.scala 143:103:@27188.4]
  wire [5:0] _T_80241; // @[Modules.scala 143:103:@27189.4]
  wire [6:0] _T_80246; // @[Modules.scala 143:103:@27193.4]
  wire [5:0] _T_80247; // @[Modules.scala 143:103:@27194.4]
  wire [5:0] _T_80248; // @[Modules.scala 143:103:@27195.4]
  wire [5:0] _T_80274; // @[Modules.scala 143:103:@27217.4]
  wire [4:0] _T_80275; // @[Modules.scala 143:103:@27218.4]
  wire [4:0] _T_80276; // @[Modules.scala 143:103:@27219.4]
  wire [5:0] _T_80281; // @[Modules.scala 143:103:@27223.4]
  wire [4:0] _T_80282; // @[Modules.scala 143:103:@27224.4]
  wire [4:0] _T_80283; // @[Modules.scala 143:103:@27225.4]
  wire [5:0] _T_80288; // @[Modules.scala 143:103:@27229.4]
  wire [4:0] _T_80289; // @[Modules.scala 143:103:@27230.4]
  wire [4:0] _T_80290; // @[Modules.scala 143:103:@27231.4]
  wire [4:0] _T_80301; // @[Modules.scala 144:80:@27240.4]
  wire [5:0] _T_80302; // @[Modules.scala 143:103:@27241.4]
  wire [4:0] _T_80303; // @[Modules.scala 143:103:@27242.4]
  wire [4:0] _T_80304; // @[Modules.scala 143:103:@27243.4]
  wire [5:0] _T_80309; // @[Modules.scala 143:103:@27247.4]
  wire [4:0] _T_80310; // @[Modules.scala 143:103:@27248.4]
  wire [4:0] _T_80311; // @[Modules.scala 143:103:@27249.4]
  wire [5:0] _T_80323; // @[Modules.scala 143:103:@27259.4]
  wire [4:0] _T_80324; // @[Modules.scala 143:103:@27260.4]
  wire [4:0] _T_80325; // @[Modules.scala 143:103:@27261.4]
  wire [6:0] _T_80330; // @[Modules.scala 143:103:@27265.4]
  wire [5:0] _T_80331; // @[Modules.scala 143:103:@27266.4]
  wire [5:0] _T_80332; // @[Modules.scala 143:103:@27267.4]
  wire [5:0] _GEN_612; // @[Modules.scala 143:103:@27277.4]
  wire [6:0] _T_80344; // @[Modules.scala 143:103:@27277.4]
  wire [5:0] _T_80345; // @[Modules.scala 143:103:@27278.4]
  wire [5:0] _T_80346; // @[Modules.scala 143:103:@27279.4]
  wire [5:0] _T_80372; // @[Modules.scala 143:103:@27301.4]
  wire [4:0] _T_80373; // @[Modules.scala 143:103:@27302.4]
  wire [4:0] _T_80374; // @[Modules.scala 143:103:@27303.4]
  wire [5:0] _T_80379; // @[Modules.scala 143:103:@27307.4]
  wire [4:0] _T_80380; // @[Modules.scala 143:103:@27308.4]
  wire [4:0] _T_80381; // @[Modules.scala 143:103:@27309.4]
  wire [5:0] _T_80386; // @[Modules.scala 143:103:@27313.4]
  wire [4:0] _T_80387; // @[Modules.scala 143:103:@27314.4]
  wire [4:0] _T_80388; // @[Modules.scala 143:103:@27315.4]
  wire [5:0] _T_80407; // @[Modules.scala 143:103:@27331.4]
  wire [4:0] _T_80408; // @[Modules.scala 143:103:@27332.4]
  wire [4:0] _T_80409; // @[Modules.scala 143:103:@27333.4]
  wire [6:0] _T_80414; // @[Modules.scala 143:103:@27337.4]
  wire [5:0] _T_80415; // @[Modules.scala 143:103:@27338.4]
  wire [5:0] _T_80416; // @[Modules.scala 143:103:@27339.4]
  wire [6:0] _T_80435; // @[Modules.scala 143:103:@27355.4]
  wire [5:0] _T_80436; // @[Modules.scala 143:103:@27356.4]
  wire [5:0] _T_80437; // @[Modules.scala 143:103:@27357.4]
  wire [6:0] _T_80442; // @[Modules.scala 143:103:@27361.4]
  wire [5:0] _T_80443; // @[Modules.scala 143:103:@27362.4]
  wire [5:0] _T_80444; // @[Modules.scala 143:103:@27363.4]
  wire [5:0] _T_80470; // @[Modules.scala 143:103:@27385.4]
  wire [4:0] _T_80471; // @[Modules.scala 143:103:@27386.4]
  wire [4:0] _T_80472; // @[Modules.scala 143:103:@27387.4]
  wire [5:0] _T_80491; // @[Modules.scala 143:103:@27403.4]
  wire [4:0] _T_80492; // @[Modules.scala 143:103:@27404.4]
  wire [4:0] _T_80493; // @[Modules.scala 143:103:@27405.4]
  wire [5:0] _T_80498; // @[Modules.scala 143:103:@27409.4]
  wire [4:0] _T_80499; // @[Modules.scala 143:103:@27410.4]
  wire [4:0] _T_80500; // @[Modules.scala 143:103:@27411.4]
  wire [6:0] _T_80505; // @[Modules.scala 143:103:@27415.4]
  wire [5:0] _T_80506; // @[Modules.scala 143:103:@27416.4]
  wire [5:0] _T_80507; // @[Modules.scala 143:103:@27417.4]
  wire [5:0] _GEN_616; // @[Modules.scala 143:103:@27433.4]
  wire [6:0] _T_80526; // @[Modules.scala 143:103:@27433.4]
  wire [5:0] _T_80527; // @[Modules.scala 143:103:@27434.4]
  wire [5:0] _T_80528; // @[Modules.scala 143:103:@27435.4]
  wire [6:0] _T_80596; // @[Modules.scala 143:103:@27493.4]
  wire [5:0] _T_80597; // @[Modules.scala 143:103:@27494.4]
  wire [5:0] _T_80598; // @[Modules.scala 143:103:@27495.4]
  wire [5:0] _GEN_617; // @[Modules.scala 143:103:@27499.4]
  wire [6:0] _T_80603; // @[Modules.scala 143:103:@27499.4]
  wire [5:0] _T_80604; // @[Modules.scala 143:103:@27500.4]
  wire [5:0] _T_80605; // @[Modules.scala 143:103:@27501.4]
  wire [6:0] _T_80617; // @[Modules.scala 143:103:@27511.4]
  wire [5:0] _T_80618; // @[Modules.scala 143:103:@27512.4]
  wire [5:0] _T_80619; // @[Modules.scala 143:103:@27513.4]
  wire [6:0] _T_80624; // @[Modules.scala 143:103:@27517.4]
  wire [5:0] _T_80625; // @[Modules.scala 143:103:@27518.4]
  wire [5:0] _T_80626; // @[Modules.scala 143:103:@27519.4]
  wire [5:0] _T_80652; // @[Modules.scala 143:103:@27541.4]
  wire [4:0] _T_80653; // @[Modules.scala 143:103:@27542.4]
  wire [4:0] _T_80654; // @[Modules.scala 143:103:@27543.4]
  wire [6:0] _T_80659; // @[Modules.scala 143:103:@27547.4]
  wire [5:0] _T_80660; // @[Modules.scala 143:103:@27548.4]
  wire [5:0] _T_80661; // @[Modules.scala 143:103:@27549.4]
  wire [6:0] _T_80673; // @[Modules.scala 143:103:@27559.4]
  wire [5:0] _T_80674; // @[Modules.scala 143:103:@27560.4]
  wire [5:0] _T_80675; // @[Modules.scala 143:103:@27561.4]
  wire [6:0] _T_80680; // @[Modules.scala 143:103:@27565.4]
  wire [5:0] _T_80681; // @[Modules.scala 143:103:@27566.4]
  wire [5:0] _T_80682; // @[Modules.scala 143:103:@27567.4]
  wire [6:0] _T_80708; // @[Modules.scala 143:103:@27589.4]
  wire [5:0] _T_80709; // @[Modules.scala 143:103:@27590.4]
  wire [5:0] _T_80710; // @[Modules.scala 143:103:@27591.4]
  wire [6:0] _T_80715; // @[Modules.scala 143:103:@27595.4]
  wire [5:0] _T_80716; // @[Modules.scala 143:103:@27596.4]
  wire [5:0] _T_80717; // @[Modules.scala 143:103:@27597.4]
  wire [6:0] _T_80799; // @[Modules.scala 143:103:@27667.4]
  wire [5:0] _T_80800; // @[Modules.scala 143:103:@27668.4]
  wire [5:0] _T_80801; // @[Modules.scala 143:103:@27669.4]
  wire [6:0] _T_80883; // @[Modules.scala 143:103:@27739.4]
  wire [5:0] _T_80884; // @[Modules.scala 143:103:@27740.4]
  wire [5:0] _T_80885; // @[Modules.scala 143:103:@27741.4]
  wire [5:0] _GEN_627; // @[Modules.scala 143:103:@27745.4]
  wire [6:0] _T_80890; // @[Modules.scala 143:103:@27745.4]
  wire [5:0] _T_80891; // @[Modules.scala 143:103:@27746.4]
  wire [5:0] _T_80892; // @[Modules.scala 143:103:@27747.4]
  wire [5:0] _T_80943; // @[Modules.scala 143:74:@27791.4]
  wire [5:0] _T_80945; // @[Modules.scala 144:80:@27792.4]
  wire [6:0] _T_80946; // @[Modules.scala 143:103:@27793.4]
  wire [5:0] _T_80947; // @[Modules.scala 143:103:@27794.4]
  wire [5:0] _T_80948; // @[Modules.scala 143:103:@27795.4]
  wire [6:0] _T_80953; // @[Modules.scala 143:103:@27799.4]
  wire [5:0] _T_80954; // @[Modules.scala 143:103:@27800.4]
  wire [5:0] _T_80955; // @[Modules.scala 143:103:@27801.4]
  wire [5:0] _GEN_630; // @[Modules.scala 143:103:@27823.4]
  wire [6:0] _T_80981; // @[Modules.scala 143:103:@27823.4]
  wire [5:0] _T_80982; // @[Modules.scala 143:103:@27824.4]
  wire [5:0] _T_80983; // @[Modules.scala 143:103:@27825.4]
  wire [5:0] _GEN_631; // @[Modules.scala 143:103:@27835.4]
  wire [6:0] _T_80995; // @[Modules.scala 143:103:@27835.4]
  wire [5:0] _T_80996; // @[Modules.scala 143:103:@27836.4]
  wire [5:0] _T_80997; // @[Modules.scala 143:103:@27837.4]
  wire [13:0] buffer_8_2; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81015; // @[Modules.scala 166:64:@27855.4]
  wire [13:0] _T_81016; // @[Modules.scala 166:64:@27856.4]
  wire [13:0] buffer_8_310; // @[Modules.scala 166:64:@27857.4]
  wire [13:0] buffer_8_5; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81018; // @[Modules.scala 166:64:@27859.4]
  wire [13:0] _T_81019; // @[Modules.scala 166:64:@27860.4]
  wire [13:0] buffer_8_311; // @[Modules.scala 166:64:@27861.4]
  wire [14:0] _T_81021; // @[Modules.scala 166:64:@27863.4]
  wire [13:0] _T_81022; // @[Modules.scala 166:64:@27864.4]
  wire [13:0] buffer_8_312; // @[Modules.scala 166:64:@27865.4]
  wire [13:0] buffer_8_8; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81024; // @[Modules.scala 166:64:@27867.4]
  wire [13:0] _T_81025; // @[Modules.scala 166:64:@27868.4]
  wire [13:0] buffer_8_313; // @[Modules.scala 166:64:@27869.4]
  wire [14:0] _T_81027; // @[Modules.scala 166:64:@27871.4]
  wire [13:0] _T_81028; // @[Modules.scala 166:64:@27872.4]
  wire [13:0] buffer_8_314; // @[Modules.scala 166:64:@27873.4]
  wire [13:0] buffer_8_12; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81030; // @[Modules.scala 166:64:@27875.4]
  wire [13:0] _T_81031; // @[Modules.scala 166:64:@27876.4]
  wire [13:0] buffer_8_315; // @[Modules.scala 166:64:@27877.4]
  wire [14:0] _T_81033; // @[Modules.scala 166:64:@27879.4]
  wire [13:0] _T_81034; // @[Modules.scala 166:64:@27880.4]
  wire [13:0] buffer_8_316; // @[Modules.scala 166:64:@27881.4]
  wire [13:0] buffer_8_22; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81045; // @[Modules.scala 166:64:@27895.4]
  wire [13:0] _T_81046; // @[Modules.scala 166:64:@27896.4]
  wire [13:0] buffer_8_320; // @[Modules.scala 166:64:@27897.4]
  wire [13:0] buffer_8_24; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81048; // @[Modules.scala 166:64:@27899.4]
  wire [13:0] _T_81049; // @[Modules.scala 166:64:@27900.4]
  wire [13:0] buffer_8_321; // @[Modules.scala 166:64:@27901.4]
  wire [13:0] buffer_8_34; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81063; // @[Modules.scala 166:64:@27919.4]
  wire [13:0] _T_81064; // @[Modules.scala 166:64:@27920.4]
  wire [13:0] buffer_8_326; // @[Modules.scala 166:64:@27921.4]
  wire [13:0] buffer_8_36; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81066; // @[Modules.scala 166:64:@27923.4]
  wire [13:0] _T_81067; // @[Modules.scala 166:64:@27924.4]
  wire [13:0] buffer_8_327; // @[Modules.scala 166:64:@27925.4]
  wire [14:0] _T_81069; // @[Modules.scala 166:64:@27927.4]
  wire [13:0] _T_81070; // @[Modules.scala 166:64:@27928.4]
  wire [13:0] buffer_8_328; // @[Modules.scala 166:64:@27929.4]
  wire [13:0] buffer_8_40; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81072; // @[Modules.scala 166:64:@27931.4]
  wire [13:0] _T_81073; // @[Modules.scala 166:64:@27932.4]
  wire [13:0] buffer_8_329; // @[Modules.scala 166:64:@27933.4]
  wire [14:0] _T_81075; // @[Modules.scala 166:64:@27935.4]
  wire [13:0] _T_81076; // @[Modules.scala 166:64:@27936.4]
  wire [13:0] buffer_8_330; // @[Modules.scala 166:64:@27937.4]
  wire [13:0] buffer_8_46; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_47; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81081; // @[Modules.scala 166:64:@27943.4]
  wire [13:0] _T_81082; // @[Modules.scala 166:64:@27944.4]
  wire [13:0] buffer_8_332; // @[Modules.scala 166:64:@27945.4]
  wire [13:0] buffer_8_48; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81084; // @[Modules.scala 166:64:@27947.4]
  wire [13:0] _T_81085; // @[Modules.scala 166:64:@27948.4]
  wire [13:0] buffer_8_333; // @[Modules.scala 166:64:@27949.4]
  wire [14:0] _T_81087; // @[Modules.scala 166:64:@27951.4]
  wire [13:0] _T_81088; // @[Modules.scala 166:64:@27952.4]
  wire [13:0] buffer_8_334; // @[Modules.scala 166:64:@27953.4]
  wire [14:0] _T_81090; // @[Modules.scala 166:64:@27955.4]
  wire [13:0] _T_81091; // @[Modules.scala 166:64:@27956.4]
  wire [13:0] buffer_8_335; // @[Modules.scala 166:64:@27957.4]
  wire [13:0] buffer_8_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81093; // @[Modules.scala 166:64:@27959.4]
  wire [13:0] _T_81094; // @[Modules.scala 166:64:@27960.4]
  wire [13:0] buffer_8_336; // @[Modules.scala 166:64:@27961.4]
  wire [13:0] buffer_8_56; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81096; // @[Modules.scala 166:64:@27963.4]
  wire [13:0] _T_81097; // @[Modules.scala 166:64:@27964.4]
  wire [13:0] buffer_8_337; // @[Modules.scala 166:64:@27965.4]
  wire [13:0] buffer_8_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81099; // @[Modules.scala 166:64:@27967.4]
  wire [13:0] _T_81100; // @[Modules.scala 166:64:@27968.4]
  wire [13:0] buffer_8_338; // @[Modules.scala 166:64:@27969.4]
  wire [13:0] buffer_8_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81102; // @[Modules.scala 166:64:@27971.4]
  wire [13:0] _T_81103; // @[Modules.scala 166:64:@27972.4]
  wire [13:0] buffer_8_339; // @[Modules.scala 166:64:@27973.4]
  wire [13:0] buffer_8_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81105; // @[Modules.scala 166:64:@27975.4]
  wire [13:0] _T_81106; // @[Modules.scala 166:64:@27976.4]
  wire [13:0] buffer_8_340; // @[Modules.scala 166:64:@27977.4]
  wire [13:0] buffer_8_64; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81108; // @[Modules.scala 166:64:@27979.4]
  wire [13:0] _T_81109; // @[Modules.scala 166:64:@27980.4]
  wire [13:0] buffer_8_341; // @[Modules.scala 166:64:@27981.4]
  wire [13:0] buffer_8_66; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81111; // @[Modules.scala 166:64:@27983.4]
  wire [13:0] _T_81112; // @[Modules.scala 166:64:@27984.4]
  wire [13:0] buffer_8_342; // @[Modules.scala 166:64:@27985.4]
  wire [13:0] buffer_8_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81114; // @[Modules.scala 166:64:@27987.4]
  wire [13:0] _T_81115; // @[Modules.scala 166:64:@27988.4]
  wire [13:0] buffer_8_343; // @[Modules.scala 166:64:@27989.4]
  wire [13:0] buffer_8_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81117; // @[Modules.scala 166:64:@27991.4]
  wire [13:0] _T_81118; // @[Modules.scala 166:64:@27992.4]
  wire [13:0] buffer_8_344; // @[Modules.scala 166:64:@27993.4]
  wire [13:0] buffer_8_74; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81123; // @[Modules.scala 166:64:@27999.4]
  wire [13:0] _T_81124; // @[Modules.scala 166:64:@28000.4]
  wire [13:0] buffer_8_346; // @[Modules.scala 166:64:@28001.4]
  wire [13:0] buffer_8_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81126; // @[Modules.scala 166:64:@28003.4]
  wire [13:0] _T_81127; // @[Modules.scala 166:64:@28004.4]
  wire [13:0] buffer_8_347; // @[Modules.scala 166:64:@28005.4]
  wire [13:0] buffer_8_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81129; // @[Modules.scala 166:64:@28007.4]
  wire [13:0] _T_81130; // @[Modules.scala 166:64:@28008.4]
  wire [13:0] buffer_8_348; // @[Modules.scala 166:64:@28009.4]
  wire [13:0] buffer_8_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81132; // @[Modules.scala 166:64:@28011.4]
  wire [13:0] _T_81133; // @[Modules.scala 166:64:@28012.4]
  wire [13:0] buffer_8_349; // @[Modules.scala 166:64:@28013.4]
  wire [13:0] buffer_8_82; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81135; // @[Modules.scala 166:64:@28015.4]
  wire [13:0] _T_81136; // @[Modules.scala 166:64:@28016.4]
  wire [13:0] buffer_8_350; // @[Modules.scala 166:64:@28017.4]
  wire [13:0] buffer_8_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81138; // @[Modules.scala 166:64:@28019.4]
  wire [13:0] _T_81139; // @[Modules.scala 166:64:@28020.4]
  wire [13:0] buffer_8_351; // @[Modules.scala 166:64:@28021.4]
  wire [13:0] buffer_8_86; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_87; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81141; // @[Modules.scala 166:64:@28023.4]
  wire [13:0] _T_81142; // @[Modules.scala 166:64:@28024.4]
  wire [13:0] buffer_8_352; // @[Modules.scala 166:64:@28025.4]
  wire [13:0] buffer_8_89; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81144; // @[Modules.scala 166:64:@28027.4]
  wire [13:0] _T_81145; // @[Modules.scala 166:64:@28028.4]
  wire [13:0] buffer_8_353; // @[Modules.scala 166:64:@28029.4]
  wire [13:0] buffer_8_92; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81150; // @[Modules.scala 166:64:@28035.4]
  wire [13:0] _T_81151; // @[Modules.scala 166:64:@28036.4]
  wire [13:0] buffer_8_355; // @[Modules.scala 166:64:@28037.4]
  wire [13:0] buffer_8_94; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81153; // @[Modules.scala 166:64:@28039.4]
  wire [13:0] _T_81154; // @[Modules.scala 166:64:@28040.4]
  wire [13:0] buffer_8_356; // @[Modules.scala 166:64:@28041.4]
  wire [14:0] _T_81159; // @[Modules.scala 166:64:@28047.4]
  wire [13:0] _T_81160; // @[Modules.scala 166:64:@28048.4]
  wire [13:0] buffer_8_358; // @[Modules.scala 166:64:@28049.4]
  wire [13:0] buffer_8_100; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_101; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81162; // @[Modules.scala 166:64:@28051.4]
  wire [13:0] _T_81163; // @[Modules.scala 166:64:@28052.4]
  wire [13:0] buffer_8_359; // @[Modules.scala 166:64:@28053.4]
  wire [14:0] _T_81165; // @[Modules.scala 166:64:@28055.4]
  wire [13:0] _T_81166; // @[Modules.scala 166:64:@28056.4]
  wire [13:0] buffer_8_360; // @[Modules.scala 166:64:@28057.4]
  wire [14:0] _T_81168; // @[Modules.scala 166:64:@28059.4]
  wire [13:0] _T_81169; // @[Modules.scala 166:64:@28060.4]
  wire [13:0] buffer_8_361; // @[Modules.scala 166:64:@28061.4]
  wire [13:0] buffer_8_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81171; // @[Modules.scala 166:64:@28063.4]
  wire [13:0] _T_81172; // @[Modules.scala 166:64:@28064.4]
  wire [13:0] buffer_8_362; // @[Modules.scala 166:64:@28065.4]
  wire [13:0] buffer_8_108; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81174; // @[Modules.scala 166:64:@28067.4]
  wire [13:0] _T_81175; // @[Modules.scala 166:64:@28068.4]
  wire [13:0] buffer_8_363; // @[Modules.scala 166:64:@28069.4]
  wire [13:0] buffer_8_110; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_111; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81177; // @[Modules.scala 166:64:@28071.4]
  wire [13:0] _T_81178; // @[Modules.scala 166:64:@28072.4]
  wire [13:0] buffer_8_364; // @[Modules.scala 166:64:@28073.4]
  wire [13:0] buffer_8_112; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81180; // @[Modules.scala 166:64:@28075.4]
  wire [13:0] _T_81181; // @[Modules.scala 166:64:@28076.4]
  wire [13:0] buffer_8_365; // @[Modules.scala 166:64:@28077.4]
  wire [14:0] _T_81183; // @[Modules.scala 166:64:@28079.4]
  wire [13:0] _T_81184; // @[Modules.scala 166:64:@28080.4]
  wire [13:0] buffer_8_366; // @[Modules.scala 166:64:@28081.4]
  wire [14:0] _T_81186; // @[Modules.scala 166:64:@28083.4]
  wire [13:0] _T_81187; // @[Modules.scala 166:64:@28084.4]
  wire [13:0] buffer_8_367; // @[Modules.scala 166:64:@28085.4]
  wire [14:0] _T_81189; // @[Modules.scala 166:64:@28087.4]
  wire [13:0] _T_81190; // @[Modules.scala 166:64:@28088.4]
  wire [13:0] buffer_8_368; // @[Modules.scala 166:64:@28089.4]
  wire [14:0] _T_81195; // @[Modules.scala 166:64:@28095.4]
  wire [13:0] _T_81196; // @[Modules.scala 166:64:@28096.4]
  wire [13:0] buffer_8_370; // @[Modules.scala 166:64:@28097.4]
  wire [13:0] buffer_8_124; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81198; // @[Modules.scala 166:64:@28099.4]
  wire [13:0] _T_81199; // @[Modules.scala 166:64:@28100.4]
  wire [13:0] buffer_8_371; // @[Modules.scala 166:64:@28101.4]
  wire [14:0] _T_81201; // @[Modules.scala 166:64:@28103.4]
  wire [13:0] _T_81202; // @[Modules.scala 166:64:@28104.4]
  wire [13:0] buffer_8_372; // @[Modules.scala 166:64:@28105.4]
  wire [14:0] _T_81207; // @[Modules.scala 166:64:@28111.4]
  wire [13:0] _T_81208; // @[Modules.scala 166:64:@28112.4]
  wire [13:0] buffer_8_374; // @[Modules.scala 166:64:@28113.4]
  wire [13:0] buffer_8_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81210; // @[Modules.scala 166:64:@28115.4]
  wire [13:0] _T_81211; // @[Modules.scala 166:64:@28116.4]
  wire [13:0] buffer_8_375; // @[Modules.scala 166:64:@28117.4]
  wire [14:0] _T_81219; // @[Modules.scala 166:64:@28127.4]
  wire [13:0] _T_81220; // @[Modules.scala 166:64:@28128.4]
  wire [13:0] buffer_8_378; // @[Modules.scala 166:64:@28129.4]
  wire [14:0] _T_81222; // @[Modules.scala 166:64:@28131.4]
  wire [13:0] _T_81223; // @[Modules.scala 166:64:@28132.4]
  wire [13:0] buffer_8_379; // @[Modules.scala 166:64:@28133.4]
  wire [14:0] _T_81225; // @[Modules.scala 166:64:@28135.4]
  wire [13:0] _T_81226; // @[Modules.scala 166:64:@28136.4]
  wire [13:0] buffer_8_380; // @[Modules.scala 166:64:@28137.4]
  wire [14:0] _T_81228; // @[Modules.scala 166:64:@28139.4]
  wire [13:0] _T_81229; // @[Modules.scala 166:64:@28140.4]
  wire [13:0] buffer_8_381; // @[Modules.scala 166:64:@28141.4]
  wire [14:0] _T_81231; // @[Modules.scala 166:64:@28143.4]
  wire [13:0] _T_81232; // @[Modules.scala 166:64:@28144.4]
  wire [13:0] buffer_8_382; // @[Modules.scala 166:64:@28145.4]
  wire [13:0] buffer_8_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81234; // @[Modules.scala 166:64:@28147.4]
  wire [13:0] _T_81235; // @[Modules.scala 166:64:@28148.4]
  wire [13:0] buffer_8_383; // @[Modules.scala 166:64:@28149.4]
  wire [13:0] buffer_8_150; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81237; // @[Modules.scala 166:64:@28151.4]
  wire [13:0] _T_81238; // @[Modules.scala 166:64:@28152.4]
  wire [13:0] buffer_8_384; // @[Modules.scala 166:64:@28153.4]
  wire [13:0] buffer_8_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81240; // @[Modules.scala 166:64:@28155.4]
  wire [13:0] _T_81241; // @[Modules.scala 166:64:@28156.4]
  wire [13:0] buffer_8_385; // @[Modules.scala 166:64:@28157.4]
  wire [13:0] buffer_8_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81243; // @[Modules.scala 166:64:@28159.4]
  wire [13:0] _T_81244; // @[Modules.scala 166:64:@28160.4]
  wire [13:0] buffer_8_386; // @[Modules.scala 166:64:@28161.4]
  wire [13:0] buffer_8_156; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81246; // @[Modules.scala 166:64:@28163.4]
  wire [13:0] _T_81247; // @[Modules.scala 166:64:@28164.4]
  wire [13:0] buffer_8_387; // @[Modules.scala 166:64:@28165.4]
  wire [13:0] buffer_8_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81249; // @[Modules.scala 166:64:@28167.4]
  wire [13:0] _T_81250; // @[Modules.scala 166:64:@28168.4]
  wire [13:0] buffer_8_388; // @[Modules.scala 166:64:@28169.4]
  wire [13:0] buffer_8_160; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81252; // @[Modules.scala 166:64:@28171.4]
  wire [13:0] _T_81253; // @[Modules.scala 166:64:@28172.4]
  wire [13:0] buffer_8_389; // @[Modules.scala 166:64:@28173.4]
  wire [13:0] buffer_8_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81258; // @[Modules.scala 166:64:@28179.4]
  wire [13:0] _T_81259; // @[Modules.scala 166:64:@28180.4]
  wire [13:0] buffer_8_391; // @[Modules.scala 166:64:@28181.4]
  wire [13:0] buffer_8_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81261; // @[Modules.scala 166:64:@28183.4]
  wire [13:0] _T_81262; // @[Modules.scala 166:64:@28184.4]
  wire [13:0] buffer_8_392; // @[Modules.scala 166:64:@28185.4]
  wire [14:0] _T_81264; // @[Modules.scala 166:64:@28187.4]
  wire [13:0] _T_81265; // @[Modules.scala 166:64:@28188.4]
  wire [13:0] buffer_8_393; // @[Modules.scala 166:64:@28189.4]
  wire [13:0] buffer_8_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81267; // @[Modules.scala 166:64:@28191.4]
  wire [13:0] _T_81268; // @[Modules.scala 166:64:@28192.4]
  wire [13:0] buffer_8_394; // @[Modules.scala 166:64:@28193.4]
  wire [13:0] buffer_8_173; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81270; // @[Modules.scala 166:64:@28195.4]
  wire [13:0] _T_81271; // @[Modules.scala 166:64:@28196.4]
  wire [13:0] buffer_8_395; // @[Modules.scala 166:64:@28197.4]
  wire [14:0] _T_81273; // @[Modules.scala 166:64:@28199.4]
  wire [13:0] _T_81274; // @[Modules.scala 166:64:@28200.4]
  wire [13:0] buffer_8_396; // @[Modules.scala 166:64:@28201.4]
  wire [13:0] buffer_8_176; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81276; // @[Modules.scala 166:64:@28203.4]
  wire [13:0] _T_81277; // @[Modules.scala 166:64:@28204.4]
  wire [13:0] buffer_8_397; // @[Modules.scala 166:64:@28205.4]
  wire [13:0] buffer_8_180; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81282; // @[Modules.scala 166:64:@28211.4]
  wire [13:0] _T_81283; // @[Modules.scala 166:64:@28212.4]
  wire [13:0] buffer_8_399; // @[Modules.scala 166:64:@28213.4]
  wire [14:0] _T_81291; // @[Modules.scala 166:64:@28223.4]
  wire [13:0] _T_81292; // @[Modules.scala 166:64:@28224.4]
  wire [13:0] buffer_8_402; // @[Modules.scala 166:64:@28225.4]
  wire [13:0] buffer_8_188; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81294; // @[Modules.scala 166:64:@28227.4]
  wire [13:0] _T_81295; // @[Modules.scala 166:64:@28228.4]
  wire [13:0] buffer_8_403; // @[Modules.scala 166:64:@28229.4]
  wire [13:0] buffer_8_190; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81297; // @[Modules.scala 166:64:@28231.4]
  wire [13:0] _T_81298; // @[Modules.scala 166:64:@28232.4]
  wire [13:0] buffer_8_404; // @[Modules.scala 166:64:@28233.4]
  wire [14:0] _T_81300; // @[Modules.scala 166:64:@28235.4]
  wire [13:0] _T_81301; // @[Modules.scala 166:64:@28236.4]
  wire [13:0] buffer_8_405; // @[Modules.scala 166:64:@28237.4]
  wire [14:0] _T_81303; // @[Modules.scala 166:64:@28239.4]
  wire [13:0] _T_81304; // @[Modules.scala 166:64:@28240.4]
  wire [13:0] buffer_8_406; // @[Modules.scala 166:64:@28241.4]
  wire [13:0] buffer_8_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81306; // @[Modules.scala 166:64:@28243.4]
  wire [13:0] _T_81307; // @[Modules.scala 166:64:@28244.4]
  wire [13:0] buffer_8_407; // @[Modules.scala 166:64:@28245.4]
  wire [13:0] buffer_8_198; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81309; // @[Modules.scala 166:64:@28247.4]
  wire [13:0] _T_81310; // @[Modules.scala 166:64:@28248.4]
  wire [13:0] buffer_8_408; // @[Modules.scala 166:64:@28249.4]
  wire [14:0] _T_81312; // @[Modules.scala 166:64:@28251.4]
  wire [13:0] _T_81313; // @[Modules.scala 166:64:@28252.4]
  wire [13:0] buffer_8_409; // @[Modules.scala 166:64:@28253.4]
  wire [13:0] buffer_8_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81315; // @[Modules.scala 166:64:@28255.4]
  wire [13:0] _T_81316; // @[Modules.scala 166:64:@28256.4]
  wire [13:0] buffer_8_410; // @[Modules.scala 166:64:@28257.4]
  wire [13:0] buffer_8_204; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81318; // @[Modules.scala 166:64:@28259.4]
  wire [13:0] _T_81319; // @[Modules.scala 166:64:@28260.4]
  wire [13:0] buffer_8_411; // @[Modules.scala 166:64:@28261.4]
  wire [13:0] buffer_8_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81321; // @[Modules.scala 166:64:@28263.4]
  wire [13:0] _T_81322; // @[Modules.scala 166:64:@28264.4]
  wire [13:0] buffer_8_412; // @[Modules.scala 166:64:@28265.4]
  wire [13:0] buffer_8_208; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81324; // @[Modules.scala 166:64:@28267.4]
  wire [13:0] _T_81325; // @[Modules.scala 166:64:@28268.4]
  wire [13:0] buffer_8_413; // @[Modules.scala 166:64:@28269.4]
  wire [13:0] buffer_8_210; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81327; // @[Modules.scala 166:64:@28271.4]
  wire [13:0] _T_81328; // @[Modules.scala 166:64:@28272.4]
  wire [13:0] buffer_8_414; // @[Modules.scala 166:64:@28273.4]
  wire [13:0] buffer_8_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81330; // @[Modules.scala 166:64:@28275.4]
  wire [13:0] _T_81331; // @[Modules.scala 166:64:@28276.4]
  wire [13:0] buffer_8_415; // @[Modules.scala 166:64:@28277.4]
  wire [13:0] buffer_8_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81336; // @[Modules.scala 166:64:@28283.4]
  wire [13:0] _T_81337; // @[Modules.scala 166:64:@28284.4]
  wire [13:0] buffer_8_417; // @[Modules.scala 166:64:@28285.4]
  wire [13:0] buffer_8_218; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81339; // @[Modules.scala 166:64:@28287.4]
  wire [13:0] _T_81340; // @[Modules.scala 166:64:@28288.4]
  wire [13:0] buffer_8_418; // @[Modules.scala 166:64:@28289.4]
  wire [13:0] buffer_8_222; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81345; // @[Modules.scala 166:64:@28295.4]
  wire [13:0] _T_81346; // @[Modules.scala 166:64:@28296.4]
  wire [13:0] buffer_8_420; // @[Modules.scala 166:64:@28297.4]
  wire [14:0] _T_81348; // @[Modules.scala 166:64:@28299.4]
  wire [13:0] _T_81349; // @[Modules.scala 166:64:@28300.4]
  wire [13:0] buffer_8_421; // @[Modules.scala 166:64:@28301.4]
  wire [13:0] buffer_8_226; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81351; // @[Modules.scala 166:64:@28303.4]
  wire [13:0] _T_81352; // @[Modules.scala 166:64:@28304.4]
  wire [13:0] buffer_8_422; // @[Modules.scala 166:64:@28305.4]
  wire [14:0] _T_81354; // @[Modules.scala 166:64:@28307.4]
  wire [13:0] _T_81355; // @[Modules.scala 166:64:@28308.4]
  wire [13:0] buffer_8_423; // @[Modules.scala 166:64:@28309.4]
  wire [13:0] buffer_8_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81357; // @[Modules.scala 166:64:@28311.4]
  wire [13:0] _T_81358; // @[Modules.scala 166:64:@28312.4]
  wire [13:0] buffer_8_424; // @[Modules.scala 166:64:@28313.4]
  wire [14:0] _T_81360; // @[Modules.scala 166:64:@28315.4]
  wire [13:0] _T_81361; // @[Modules.scala 166:64:@28316.4]
  wire [13:0] buffer_8_425; // @[Modules.scala 166:64:@28317.4]
  wire [13:0] buffer_8_234; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81363; // @[Modules.scala 166:64:@28319.4]
  wire [13:0] _T_81364; // @[Modules.scala 166:64:@28320.4]
  wire [13:0] buffer_8_426; // @[Modules.scala 166:64:@28321.4]
  wire [13:0] buffer_8_236; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81366; // @[Modules.scala 166:64:@28323.4]
  wire [13:0] _T_81367; // @[Modules.scala 166:64:@28324.4]
  wire [13:0] buffer_8_427; // @[Modules.scala 166:64:@28325.4]
  wire [13:0] buffer_8_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81369; // @[Modules.scala 166:64:@28327.4]
  wire [13:0] _T_81370; // @[Modules.scala 166:64:@28328.4]
  wire [13:0] buffer_8_428; // @[Modules.scala 166:64:@28329.4]
  wire [14:0] _T_81372; // @[Modules.scala 166:64:@28331.4]
  wire [13:0] _T_81373; // @[Modules.scala 166:64:@28332.4]
  wire [13:0] buffer_8_429; // @[Modules.scala 166:64:@28333.4]
  wire [14:0] _T_81375; // @[Modules.scala 166:64:@28335.4]
  wire [13:0] _T_81376; // @[Modules.scala 166:64:@28336.4]
  wire [13:0] buffer_8_430; // @[Modules.scala 166:64:@28337.4]
  wire [14:0] _T_81381; // @[Modules.scala 166:64:@28343.4]
  wire [13:0] _T_81382; // @[Modules.scala 166:64:@28344.4]
  wire [13:0] buffer_8_432; // @[Modules.scala 166:64:@28345.4]
  wire [13:0] buffer_8_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81384; // @[Modules.scala 166:64:@28347.4]
  wire [13:0] _T_81385; // @[Modules.scala 166:64:@28348.4]
  wire [13:0] buffer_8_433; // @[Modules.scala 166:64:@28349.4]
  wire [13:0] buffer_8_250; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81387; // @[Modules.scala 166:64:@28351.4]
  wire [13:0] _T_81388; // @[Modules.scala 166:64:@28352.4]
  wire [13:0] buffer_8_434; // @[Modules.scala 166:64:@28353.4]
  wire [13:0] buffer_8_252; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81390; // @[Modules.scala 166:64:@28355.4]
  wire [13:0] _T_81391; // @[Modules.scala 166:64:@28356.4]
  wire [13:0] buffer_8_435; // @[Modules.scala 166:64:@28357.4]
  wire [14:0] _T_81393; // @[Modules.scala 166:64:@28359.4]
  wire [13:0] _T_81394; // @[Modules.scala 166:64:@28360.4]
  wire [13:0] buffer_8_436; // @[Modules.scala 166:64:@28361.4]
  wire [13:0] buffer_8_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81396; // @[Modules.scala 166:64:@28363.4]
  wire [13:0] _T_81397; // @[Modules.scala 166:64:@28364.4]
  wire [13:0] buffer_8_437; // @[Modules.scala 166:64:@28365.4]
  wire [13:0] buffer_8_258; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81399; // @[Modules.scala 166:64:@28367.4]
  wire [13:0] _T_81400; // @[Modules.scala 166:64:@28368.4]
  wire [13:0] buffer_8_438; // @[Modules.scala 166:64:@28369.4]
  wire [13:0] buffer_8_260; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_261; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81402; // @[Modules.scala 166:64:@28371.4]
  wire [13:0] _T_81403; // @[Modules.scala 166:64:@28372.4]
  wire [13:0] buffer_8_439; // @[Modules.scala 166:64:@28373.4]
  wire [14:0] _T_81405; // @[Modules.scala 166:64:@28375.4]
  wire [13:0] _T_81406; // @[Modules.scala 166:64:@28376.4]
  wire [13:0] buffer_8_440; // @[Modules.scala 166:64:@28377.4]
  wire [13:0] buffer_8_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81408; // @[Modules.scala 166:64:@28379.4]
  wire [13:0] _T_81409; // @[Modules.scala 166:64:@28380.4]
  wire [13:0] buffer_8_441; // @[Modules.scala 166:64:@28381.4]
  wire [13:0] buffer_8_266; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81411; // @[Modules.scala 166:64:@28383.4]
  wire [13:0] _T_81412; // @[Modules.scala 166:64:@28384.4]
  wire [13:0] buffer_8_442; // @[Modules.scala 166:64:@28385.4]
  wire [14:0] _T_81414; // @[Modules.scala 166:64:@28387.4]
  wire [13:0] _T_81415; // @[Modules.scala 166:64:@28388.4]
  wire [13:0] buffer_8_443; // @[Modules.scala 166:64:@28389.4]
  wire [14:0] _T_81417; // @[Modules.scala 166:64:@28391.4]
  wire [13:0] _T_81418; // @[Modules.scala 166:64:@28392.4]
  wire [13:0] buffer_8_444; // @[Modules.scala 166:64:@28393.4]
  wire [14:0] _T_81426; // @[Modules.scala 166:64:@28403.4]
  wire [13:0] _T_81427; // @[Modules.scala 166:64:@28404.4]
  wire [13:0] buffer_8_447; // @[Modules.scala 166:64:@28405.4]
  wire [13:0] buffer_8_278; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81429; // @[Modules.scala 166:64:@28407.4]
  wire [13:0] _T_81430; // @[Modules.scala 166:64:@28408.4]
  wire [13:0] buffer_8_448; // @[Modules.scala 166:64:@28409.4]
  wire [14:0] _T_81444; // @[Modules.scala 166:64:@28427.4]
  wire [13:0] _T_81445; // @[Modules.scala 166:64:@28428.4]
  wire [13:0] buffer_8_453; // @[Modules.scala 166:64:@28429.4]
  wire [13:0] buffer_8_290; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_8_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81447; // @[Modules.scala 166:64:@28431.4]
  wire [13:0] _T_81448; // @[Modules.scala 166:64:@28432.4]
  wire [13:0] buffer_8_454; // @[Modules.scala 166:64:@28433.4]
  wire [14:0] _T_81453; // @[Modules.scala 166:64:@28439.4]
  wire [13:0] _T_81454; // @[Modules.scala 166:64:@28440.4]
  wire [13:0] buffer_8_456; // @[Modules.scala 166:64:@28441.4]
  wire [14:0] _T_81456; // @[Modules.scala 166:64:@28443.4]
  wire [13:0] _T_81457; // @[Modules.scala 166:64:@28444.4]
  wire [13:0] buffer_8_457; // @[Modules.scala 166:64:@28445.4]
  wire [13:0] buffer_8_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81459; // @[Modules.scala 166:64:@28447.4]
  wire [13:0] _T_81460; // @[Modules.scala 166:64:@28448.4]
  wire [13:0] buffer_8_458; // @[Modules.scala 166:64:@28449.4]
  wire [13:0] buffer_8_300; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81462; // @[Modules.scala 166:64:@28451.4]
  wire [13:0] _T_81463; // @[Modules.scala 166:64:@28452.4]
  wire [13:0] buffer_8_459; // @[Modules.scala 166:64:@28453.4]
  wire [13:0] buffer_8_304; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81468; // @[Modules.scala 166:64:@28459.4]
  wire [13:0] _T_81469; // @[Modules.scala 166:64:@28460.4]
  wire [13:0] buffer_8_461; // @[Modules.scala 166:64:@28461.4]
  wire [13:0] buffer_8_306; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_81471; // @[Modules.scala 166:64:@28463.4]
  wire [13:0] _T_81472; // @[Modules.scala 166:64:@28464.4]
  wire [13:0] buffer_8_462; // @[Modules.scala 166:64:@28465.4]
  wire [14:0] _T_81474; // @[Modules.scala 160:64:@28467.4]
  wire [13:0] _T_81475; // @[Modules.scala 160:64:@28468.4]
  wire [13:0] buffer_8_463; // @[Modules.scala 160:64:@28469.4]
  wire [14:0] _T_81477; // @[Modules.scala 160:64:@28471.4]
  wire [13:0] _T_81478; // @[Modules.scala 160:64:@28472.4]
  wire [13:0] buffer_8_464; // @[Modules.scala 160:64:@28473.4]
  wire [14:0] _T_81480; // @[Modules.scala 160:64:@28475.4]
  wire [13:0] _T_81481; // @[Modules.scala 160:64:@28476.4]
  wire [13:0] buffer_8_465; // @[Modules.scala 160:64:@28477.4]
  wire [14:0] _T_81483; // @[Modules.scala 160:64:@28479.4]
  wire [13:0] _T_81484; // @[Modules.scala 160:64:@28480.4]
  wire [13:0] buffer_8_466; // @[Modules.scala 160:64:@28481.4]
  wire [14:0] _T_81486; // @[Modules.scala 160:64:@28483.4]
  wire [13:0] _T_81487; // @[Modules.scala 160:64:@28484.4]
  wire [13:0] buffer_8_467; // @[Modules.scala 160:64:@28485.4]
  wire [14:0] _T_81489; // @[Modules.scala 160:64:@28487.4]
  wire [13:0] _T_81490; // @[Modules.scala 160:64:@28488.4]
  wire [13:0] buffer_8_468; // @[Modules.scala 160:64:@28489.4]
  wire [14:0] _T_81492; // @[Modules.scala 160:64:@28491.4]
  wire [13:0] _T_81493; // @[Modules.scala 160:64:@28492.4]
  wire [13:0] buffer_8_469; // @[Modules.scala 160:64:@28493.4]
  wire [14:0] _T_81495; // @[Modules.scala 160:64:@28495.4]
  wire [13:0] _T_81496; // @[Modules.scala 160:64:@28496.4]
  wire [13:0] buffer_8_470; // @[Modules.scala 160:64:@28497.4]
  wire [14:0] _T_81498; // @[Modules.scala 160:64:@28499.4]
  wire [13:0] _T_81499; // @[Modules.scala 160:64:@28500.4]
  wire [13:0] buffer_8_471; // @[Modules.scala 160:64:@28501.4]
  wire [14:0] _T_81501; // @[Modules.scala 160:64:@28503.4]
  wire [13:0] _T_81502; // @[Modules.scala 160:64:@28504.4]
  wire [13:0] buffer_8_472; // @[Modules.scala 160:64:@28505.4]
  wire [14:0] _T_81504; // @[Modules.scala 160:64:@28507.4]
  wire [13:0] _T_81505; // @[Modules.scala 160:64:@28508.4]
  wire [13:0] buffer_8_473; // @[Modules.scala 160:64:@28509.4]
  wire [14:0] _T_81507; // @[Modules.scala 160:64:@28511.4]
  wire [13:0] _T_81508; // @[Modules.scala 160:64:@28512.4]
  wire [13:0] buffer_8_474; // @[Modules.scala 160:64:@28513.4]
  wire [14:0] _T_81510; // @[Modules.scala 160:64:@28515.4]
  wire [13:0] _T_81511; // @[Modules.scala 160:64:@28516.4]
  wire [13:0] buffer_8_475; // @[Modules.scala 160:64:@28517.4]
  wire [14:0] _T_81513; // @[Modules.scala 160:64:@28519.4]
  wire [13:0] _T_81514; // @[Modules.scala 160:64:@28520.4]
  wire [13:0] buffer_8_476; // @[Modules.scala 160:64:@28521.4]
  wire [14:0] _T_81516; // @[Modules.scala 160:64:@28523.4]
  wire [13:0] _T_81517; // @[Modules.scala 160:64:@28524.4]
  wire [13:0] buffer_8_477; // @[Modules.scala 160:64:@28525.4]
  wire [14:0] _T_81519; // @[Modules.scala 160:64:@28527.4]
  wire [13:0] _T_81520; // @[Modules.scala 160:64:@28528.4]
  wire [13:0] buffer_8_478; // @[Modules.scala 160:64:@28529.4]
  wire [14:0] _T_81522; // @[Modules.scala 160:64:@28531.4]
  wire [13:0] _T_81523; // @[Modules.scala 160:64:@28532.4]
  wire [13:0] buffer_8_479; // @[Modules.scala 160:64:@28533.4]
  wire [14:0] _T_81525; // @[Modules.scala 160:64:@28535.4]
  wire [13:0] _T_81526; // @[Modules.scala 160:64:@28536.4]
  wire [13:0] buffer_8_480; // @[Modules.scala 160:64:@28537.4]
  wire [14:0] _T_81528; // @[Modules.scala 160:64:@28539.4]
  wire [13:0] _T_81529; // @[Modules.scala 160:64:@28540.4]
  wire [13:0] buffer_8_481; // @[Modules.scala 160:64:@28541.4]
  wire [14:0] _T_81531; // @[Modules.scala 160:64:@28543.4]
  wire [13:0] _T_81532; // @[Modules.scala 160:64:@28544.4]
  wire [13:0] buffer_8_482; // @[Modules.scala 160:64:@28545.4]
  wire [14:0] _T_81534; // @[Modules.scala 160:64:@28547.4]
  wire [13:0] _T_81535; // @[Modules.scala 160:64:@28548.4]
  wire [13:0] buffer_8_483; // @[Modules.scala 160:64:@28549.4]
  wire [14:0] _T_81537; // @[Modules.scala 160:64:@28551.4]
  wire [13:0] _T_81538; // @[Modules.scala 160:64:@28552.4]
  wire [13:0] buffer_8_484; // @[Modules.scala 160:64:@28553.4]
  wire [14:0] _T_81540; // @[Modules.scala 160:64:@28555.4]
  wire [13:0] _T_81541; // @[Modules.scala 160:64:@28556.4]
  wire [13:0] buffer_8_485; // @[Modules.scala 160:64:@28557.4]
  wire [14:0] _T_81543; // @[Modules.scala 160:64:@28559.4]
  wire [13:0] _T_81544; // @[Modules.scala 160:64:@28560.4]
  wire [13:0] buffer_8_486; // @[Modules.scala 160:64:@28561.4]
  wire [14:0] _T_81546; // @[Modules.scala 160:64:@28563.4]
  wire [13:0] _T_81547; // @[Modules.scala 160:64:@28564.4]
  wire [13:0] buffer_8_487; // @[Modules.scala 160:64:@28565.4]
  wire [14:0] _T_81549; // @[Modules.scala 160:64:@28567.4]
  wire [13:0] _T_81550; // @[Modules.scala 160:64:@28568.4]
  wire [13:0] buffer_8_488; // @[Modules.scala 160:64:@28569.4]
  wire [14:0] _T_81552; // @[Modules.scala 160:64:@28571.4]
  wire [13:0] _T_81553; // @[Modules.scala 160:64:@28572.4]
  wire [13:0] buffer_8_489; // @[Modules.scala 160:64:@28573.4]
  wire [14:0] _T_81555; // @[Modules.scala 160:64:@28575.4]
  wire [13:0] _T_81556; // @[Modules.scala 160:64:@28576.4]
  wire [13:0] buffer_8_490; // @[Modules.scala 160:64:@28577.4]
  wire [14:0] _T_81558; // @[Modules.scala 160:64:@28579.4]
  wire [13:0] _T_81559; // @[Modules.scala 160:64:@28580.4]
  wire [13:0] buffer_8_491; // @[Modules.scala 160:64:@28581.4]
  wire [14:0] _T_81561; // @[Modules.scala 160:64:@28583.4]
  wire [13:0] _T_81562; // @[Modules.scala 160:64:@28584.4]
  wire [13:0] buffer_8_492; // @[Modules.scala 160:64:@28585.4]
  wire [14:0] _T_81564; // @[Modules.scala 160:64:@28587.4]
  wire [13:0] _T_81565; // @[Modules.scala 160:64:@28588.4]
  wire [13:0] buffer_8_493; // @[Modules.scala 160:64:@28589.4]
  wire [14:0] _T_81567; // @[Modules.scala 160:64:@28591.4]
  wire [13:0] _T_81568; // @[Modules.scala 160:64:@28592.4]
  wire [13:0] buffer_8_494; // @[Modules.scala 160:64:@28593.4]
  wire [14:0] _T_81570; // @[Modules.scala 160:64:@28595.4]
  wire [13:0] _T_81571; // @[Modules.scala 160:64:@28596.4]
  wire [13:0] buffer_8_495; // @[Modules.scala 160:64:@28597.4]
  wire [14:0] _T_81573; // @[Modules.scala 160:64:@28599.4]
  wire [13:0] _T_81574; // @[Modules.scala 160:64:@28600.4]
  wire [13:0] buffer_8_496; // @[Modules.scala 160:64:@28601.4]
  wire [14:0] _T_81576; // @[Modules.scala 160:64:@28603.4]
  wire [13:0] _T_81577; // @[Modules.scala 160:64:@28604.4]
  wire [13:0] buffer_8_497; // @[Modules.scala 160:64:@28605.4]
  wire [14:0] _T_81579; // @[Modules.scala 160:64:@28607.4]
  wire [13:0] _T_81580; // @[Modules.scala 160:64:@28608.4]
  wire [13:0] buffer_8_498; // @[Modules.scala 160:64:@28609.4]
  wire [14:0] _T_81582; // @[Modules.scala 160:64:@28611.4]
  wire [13:0] _T_81583; // @[Modules.scala 160:64:@28612.4]
  wire [13:0] buffer_8_499; // @[Modules.scala 160:64:@28613.4]
  wire [14:0] _T_81585; // @[Modules.scala 160:64:@28615.4]
  wire [13:0] _T_81586; // @[Modules.scala 160:64:@28616.4]
  wire [13:0] buffer_8_500; // @[Modules.scala 160:64:@28617.4]
  wire [14:0] _T_81588; // @[Modules.scala 160:64:@28619.4]
  wire [13:0] _T_81589; // @[Modules.scala 160:64:@28620.4]
  wire [13:0] buffer_8_501; // @[Modules.scala 160:64:@28621.4]
  wire [14:0] _T_81591; // @[Modules.scala 160:64:@28623.4]
  wire [13:0] _T_81592; // @[Modules.scala 160:64:@28624.4]
  wire [13:0] buffer_8_502; // @[Modules.scala 160:64:@28625.4]
  wire [14:0] _T_81594; // @[Modules.scala 160:64:@28627.4]
  wire [13:0] _T_81595; // @[Modules.scala 160:64:@28628.4]
  wire [13:0] buffer_8_503; // @[Modules.scala 160:64:@28629.4]
  wire [14:0] _T_81597; // @[Modules.scala 160:64:@28631.4]
  wire [13:0] _T_81598; // @[Modules.scala 160:64:@28632.4]
  wire [13:0] buffer_8_504; // @[Modules.scala 160:64:@28633.4]
  wire [14:0] _T_81600; // @[Modules.scala 160:64:@28635.4]
  wire [13:0] _T_81601; // @[Modules.scala 160:64:@28636.4]
  wire [13:0] buffer_8_505; // @[Modules.scala 160:64:@28637.4]
  wire [14:0] _T_81603; // @[Modules.scala 160:64:@28639.4]
  wire [13:0] _T_81604; // @[Modules.scala 160:64:@28640.4]
  wire [13:0] buffer_8_506; // @[Modules.scala 160:64:@28641.4]
  wire [14:0] _T_81606; // @[Modules.scala 160:64:@28643.4]
  wire [13:0] _T_81607; // @[Modules.scala 160:64:@28644.4]
  wire [13:0] buffer_8_507; // @[Modules.scala 160:64:@28645.4]
  wire [14:0] _T_81609; // @[Modules.scala 160:64:@28647.4]
  wire [13:0] _T_81610; // @[Modules.scala 160:64:@28648.4]
  wire [13:0] buffer_8_508; // @[Modules.scala 160:64:@28649.4]
  wire [14:0] _T_81612; // @[Modules.scala 160:64:@28651.4]
  wire [13:0] _T_81613; // @[Modules.scala 160:64:@28652.4]
  wire [13:0] buffer_8_509; // @[Modules.scala 160:64:@28653.4]
  wire [14:0] _T_81615; // @[Modules.scala 160:64:@28655.4]
  wire [13:0] _T_81616; // @[Modules.scala 160:64:@28656.4]
  wire [13:0] buffer_8_510; // @[Modules.scala 160:64:@28657.4]
  wire [14:0] _T_81618; // @[Modules.scala 160:64:@28659.4]
  wire [13:0] _T_81619; // @[Modules.scala 160:64:@28660.4]
  wire [13:0] buffer_8_511; // @[Modules.scala 160:64:@28661.4]
  wire [14:0] _T_81621; // @[Modules.scala 160:64:@28663.4]
  wire [13:0] _T_81622; // @[Modules.scala 160:64:@28664.4]
  wire [13:0] buffer_8_512; // @[Modules.scala 160:64:@28665.4]
  wire [14:0] _T_81624; // @[Modules.scala 160:64:@28667.4]
  wire [13:0] _T_81625; // @[Modules.scala 160:64:@28668.4]
  wire [13:0] buffer_8_513; // @[Modules.scala 160:64:@28669.4]
  wire [14:0] _T_81627; // @[Modules.scala 160:64:@28671.4]
  wire [13:0] _T_81628; // @[Modules.scala 160:64:@28672.4]
  wire [13:0] buffer_8_514; // @[Modules.scala 160:64:@28673.4]
  wire [14:0] _T_81630; // @[Modules.scala 160:64:@28675.4]
  wire [13:0] _T_81631; // @[Modules.scala 160:64:@28676.4]
  wire [13:0] buffer_8_515; // @[Modules.scala 160:64:@28677.4]
  wire [14:0] _T_81633; // @[Modules.scala 160:64:@28679.4]
  wire [13:0] _T_81634; // @[Modules.scala 160:64:@28680.4]
  wire [13:0] buffer_8_516; // @[Modules.scala 160:64:@28681.4]
  wire [14:0] _T_81636; // @[Modules.scala 160:64:@28683.4]
  wire [13:0] _T_81637; // @[Modules.scala 160:64:@28684.4]
  wire [13:0] buffer_8_517; // @[Modules.scala 160:64:@28685.4]
  wire [14:0] _T_81639; // @[Modules.scala 160:64:@28687.4]
  wire [13:0] _T_81640; // @[Modules.scala 160:64:@28688.4]
  wire [13:0] buffer_8_518; // @[Modules.scala 160:64:@28689.4]
  wire [14:0] _T_81642; // @[Modules.scala 160:64:@28691.4]
  wire [13:0] _T_81643; // @[Modules.scala 160:64:@28692.4]
  wire [13:0] buffer_8_519; // @[Modules.scala 160:64:@28693.4]
  wire [14:0] _T_81645; // @[Modules.scala 160:64:@28695.4]
  wire [13:0] _T_81646; // @[Modules.scala 160:64:@28696.4]
  wire [13:0] buffer_8_520; // @[Modules.scala 160:64:@28697.4]
  wire [14:0] _T_81648; // @[Modules.scala 160:64:@28699.4]
  wire [13:0] _T_81649; // @[Modules.scala 160:64:@28700.4]
  wire [13:0] buffer_8_521; // @[Modules.scala 160:64:@28701.4]
  wire [14:0] _T_81651; // @[Modules.scala 160:64:@28703.4]
  wire [13:0] _T_81652; // @[Modules.scala 160:64:@28704.4]
  wire [13:0] buffer_8_522; // @[Modules.scala 160:64:@28705.4]
  wire [14:0] _T_81654; // @[Modules.scala 160:64:@28707.4]
  wire [13:0] _T_81655; // @[Modules.scala 160:64:@28708.4]
  wire [13:0] buffer_8_523; // @[Modules.scala 160:64:@28709.4]
  wire [14:0] _T_81657; // @[Modules.scala 160:64:@28711.4]
  wire [13:0] _T_81658; // @[Modules.scala 160:64:@28712.4]
  wire [13:0] buffer_8_524; // @[Modules.scala 160:64:@28713.4]
  wire [14:0] _T_81660; // @[Modules.scala 160:64:@28715.4]
  wire [13:0] _T_81661; // @[Modules.scala 160:64:@28716.4]
  wire [13:0] buffer_8_525; // @[Modules.scala 160:64:@28717.4]
  wire [14:0] _T_81663; // @[Modules.scala 160:64:@28719.4]
  wire [13:0] _T_81664; // @[Modules.scala 160:64:@28720.4]
  wire [13:0] buffer_8_526; // @[Modules.scala 160:64:@28721.4]
  wire [14:0] _T_81666; // @[Modules.scala 160:64:@28723.4]
  wire [13:0] _T_81667; // @[Modules.scala 160:64:@28724.4]
  wire [13:0] buffer_8_527; // @[Modules.scala 160:64:@28725.4]
  wire [14:0] _T_81669; // @[Modules.scala 160:64:@28727.4]
  wire [13:0] _T_81670; // @[Modules.scala 160:64:@28728.4]
  wire [13:0] buffer_8_528; // @[Modules.scala 160:64:@28729.4]
  wire [14:0] _T_81672; // @[Modules.scala 160:64:@28731.4]
  wire [13:0] _T_81673; // @[Modules.scala 160:64:@28732.4]
  wire [13:0] buffer_8_529; // @[Modules.scala 160:64:@28733.4]
  wire [14:0] _T_81675; // @[Modules.scala 160:64:@28735.4]
  wire [13:0] _T_81676; // @[Modules.scala 160:64:@28736.4]
  wire [13:0] buffer_8_530; // @[Modules.scala 160:64:@28737.4]
  wire [14:0] _T_81681; // @[Modules.scala 160:64:@28743.4]
  wire [13:0] _T_81682; // @[Modules.scala 160:64:@28744.4]
  wire [13:0] buffer_8_532; // @[Modules.scala 160:64:@28745.4]
  wire [14:0] _T_81684; // @[Modules.scala 160:64:@28747.4]
  wire [13:0] _T_81685; // @[Modules.scala 160:64:@28748.4]
  wire [13:0] buffer_8_533; // @[Modules.scala 160:64:@28749.4]
  wire [14:0] _T_81687; // @[Modules.scala 160:64:@28751.4]
  wire [13:0] _T_81688; // @[Modules.scala 160:64:@28752.4]
  wire [13:0] buffer_8_534; // @[Modules.scala 160:64:@28753.4]
  wire [14:0] _T_81690; // @[Modules.scala 160:64:@28755.4]
  wire [13:0] _T_81691; // @[Modules.scala 160:64:@28756.4]
  wire [13:0] buffer_8_535; // @[Modules.scala 160:64:@28757.4]
  wire [14:0] _T_81693; // @[Modules.scala 160:64:@28759.4]
  wire [13:0] _T_81694; // @[Modules.scala 160:64:@28760.4]
  wire [13:0] buffer_8_536; // @[Modules.scala 160:64:@28761.4]
  wire [14:0] _T_81696; // @[Modules.scala 160:64:@28763.4]
  wire [13:0] _T_81697; // @[Modules.scala 160:64:@28764.4]
  wire [13:0] buffer_8_537; // @[Modules.scala 160:64:@28765.4]
  wire [14:0] _T_81699; // @[Modules.scala 160:64:@28767.4]
  wire [13:0] _T_81700; // @[Modules.scala 160:64:@28768.4]
  wire [13:0] buffer_8_538; // @[Modules.scala 160:64:@28769.4]
  wire [14:0] _T_81702; // @[Modules.scala 160:64:@28771.4]
  wire [13:0] _T_81703; // @[Modules.scala 160:64:@28772.4]
  wire [13:0] buffer_8_539; // @[Modules.scala 160:64:@28773.4]
  wire [14:0] _T_81705; // @[Modules.scala 166:64:@28775.4]
  wire [13:0] _T_81706; // @[Modules.scala 166:64:@28776.4]
  wire [13:0] buffer_8_540; // @[Modules.scala 166:64:@28777.4]
  wire [14:0] _T_81708; // @[Modules.scala 166:64:@28779.4]
  wire [13:0] _T_81709; // @[Modules.scala 166:64:@28780.4]
  wire [13:0] buffer_8_541; // @[Modules.scala 166:64:@28781.4]
  wire [14:0] _T_81711; // @[Modules.scala 166:64:@28783.4]
  wire [13:0] _T_81712; // @[Modules.scala 166:64:@28784.4]
  wire [13:0] buffer_8_542; // @[Modules.scala 166:64:@28785.4]
  wire [14:0] _T_81714; // @[Modules.scala 166:64:@28787.4]
  wire [13:0] _T_81715; // @[Modules.scala 166:64:@28788.4]
  wire [13:0] buffer_8_543; // @[Modules.scala 166:64:@28789.4]
  wire [14:0] _T_81717; // @[Modules.scala 166:64:@28791.4]
  wire [13:0] _T_81718; // @[Modules.scala 166:64:@28792.4]
  wire [13:0] buffer_8_544; // @[Modules.scala 166:64:@28793.4]
  wire [14:0] _T_81720; // @[Modules.scala 166:64:@28795.4]
  wire [13:0] _T_81721; // @[Modules.scala 166:64:@28796.4]
  wire [13:0] buffer_8_545; // @[Modules.scala 166:64:@28797.4]
  wire [14:0] _T_81723; // @[Modules.scala 166:64:@28799.4]
  wire [13:0] _T_81724; // @[Modules.scala 166:64:@28800.4]
  wire [13:0] buffer_8_546; // @[Modules.scala 166:64:@28801.4]
  wire [14:0] _T_81726; // @[Modules.scala 166:64:@28803.4]
  wire [13:0] _T_81727; // @[Modules.scala 166:64:@28804.4]
  wire [13:0] buffer_8_547; // @[Modules.scala 166:64:@28805.4]
  wire [14:0] _T_81729; // @[Modules.scala 166:64:@28807.4]
  wire [13:0] _T_81730; // @[Modules.scala 166:64:@28808.4]
  wire [13:0] buffer_8_548; // @[Modules.scala 166:64:@28809.4]
  wire [14:0] _T_81732; // @[Modules.scala 166:64:@28811.4]
  wire [13:0] _T_81733; // @[Modules.scala 166:64:@28812.4]
  wire [13:0] buffer_8_549; // @[Modules.scala 166:64:@28813.4]
  wire [14:0] _T_81735; // @[Modules.scala 166:64:@28815.4]
  wire [13:0] _T_81736; // @[Modules.scala 166:64:@28816.4]
  wire [13:0] buffer_8_550; // @[Modules.scala 166:64:@28817.4]
  wire [14:0] _T_81738; // @[Modules.scala 166:64:@28819.4]
  wire [13:0] _T_81739; // @[Modules.scala 166:64:@28820.4]
  wire [13:0] buffer_8_551; // @[Modules.scala 166:64:@28821.4]
  wire [14:0] _T_81741; // @[Modules.scala 166:64:@28823.4]
  wire [13:0] _T_81742; // @[Modules.scala 166:64:@28824.4]
  wire [13:0] buffer_8_552; // @[Modules.scala 166:64:@28825.4]
  wire [14:0] _T_81744; // @[Modules.scala 166:64:@28827.4]
  wire [13:0] _T_81745; // @[Modules.scala 166:64:@28828.4]
  wire [13:0] buffer_8_553; // @[Modules.scala 166:64:@28829.4]
  wire [14:0] _T_81747; // @[Modules.scala 166:64:@28831.4]
  wire [13:0] _T_81748; // @[Modules.scala 166:64:@28832.4]
  wire [13:0] buffer_8_554; // @[Modules.scala 166:64:@28833.4]
  wire [14:0] _T_81750; // @[Modules.scala 166:64:@28835.4]
  wire [13:0] _T_81751; // @[Modules.scala 166:64:@28836.4]
  wire [13:0] buffer_8_555; // @[Modules.scala 166:64:@28837.4]
  wire [14:0] _T_81753; // @[Modules.scala 166:64:@28839.4]
  wire [13:0] _T_81754; // @[Modules.scala 166:64:@28840.4]
  wire [13:0] buffer_8_556; // @[Modules.scala 166:64:@28841.4]
  wire [14:0] _T_81756; // @[Modules.scala 166:64:@28843.4]
  wire [13:0] _T_81757; // @[Modules.scala 166:64:@28844.4]
  wire [13:0] buffer_8_557; // @[Modules.scala 166:64:@28845.4]
  wire [14:0] _T_81759; // @[Modules.scala 166:64:@28847.4]
  wire [13:0] _T_81760; // @[Modules.scala 166:64:@28848.4]
  wire [13:0] buffer_8_558; // @[Modules.scala 166:64:@28849.4]
  wire [14:0] _T_81762; // @[Modules.scala 166:64:@28851.4]
  wire [13:0] _T_81763; // @[Modules.scala 166:64:@28852.4]
  wire [13:0] buffer_8_559; // @[Modules.scala 166:64:@28853.4]
  wire [14:0] _T_81765; // @[Modules.scala 166:64:@28855.4]
  wire [13:0] _T_81766; // @[Modules.scala 166:64:@28856.4]
  wire [13:0] buffer_8_560; // @[Modules.scala 166:64:@28857.4]
  wire [14:0] _T_81768; // @[Modules.scala 166:64:@28859.4]
  wire [13:0] _T_81769; // @[Modules.scala 166:64:@28860.4]
  wire [13:0] buffer_8_561; // @[Modules.scala 166:64:@28861.4]
  wire [14:0] _T_81771; // @[Modules.scala 166:64:@28863.4]
  wire [13:0] _T_81772; // @[Modules.scala 166:64:@28864.4]
  wire [13:0] buffer_8_562; // @[Modules.scala 166:64:@28865.4]
  wire [14:0] _T_81774; // @[Modules.scala 166:64:@28867.4]
  wire [13:0] _T_81775; // @[Modules.scala 166:64:@28868.4]
  wire [13:0] buffer_8_563; // @[Modules.scala 166:64:@28869.4]
  wire [14:0] _T_81777; // @[Modules.scala 166:64:@28871.4]
  wire [13:0] _T_81778; // @[Modules.scala 166:64:@28872.4]
  wire [13:0] buffer_8_564; // @[Modules.scala 166:64:@28873.4]
  wire [14:0] _T_81780; // @[Modules.scala 166:64:@28875.4]
  wire [13:0] _T_81781; // @[Modules.scala 166:64:@28876.4]
  wire [13:0] buffer_8_565; // @[Modules.scala 166:64:@28877.4]
  wire [14:0] _T_81783; // @[Modules.scala 166:64:@28879.4]
  wire [13:0] _T_81784; // @[Modules.scala 166:64:@28880.4]
  wire [13:0] buffer_8_566; // @[Modules.scala 166:64:@28881.4]
  wire [14:0] _T_81786; // @[Modules.scala 166:64:@28883.4]
  wire [13:0] _T_81787; // @[Modules.scala 166:64:@28884.4]
  wire [13:0] buffer_8_567; // @[Modules.scala 166:64:@28885.4]
  wire [14:0] _T_81789; // @[Modules.scala 166:64:@28887.4]
  wire [13:0] _T_81790; // @[Modules.scala 166:64:@28888.4]
  wire [13:0] buffer_8_568; // @[Modules.scala 166:64:@28889.4]
  wire [14:0] _T_81792; // @[Modules.scala 166:64:@28891.4]
  wire [13:0] _T_81793; // @[Modules.scala 166:64:@28892.4]
  wire [13:0] buffer_8_569; // @[Modules.scala 166:64:@28893.4]
  wire [14:0] _T_81795; // @[Modules.scala 166:64:@28895.4]
  wire [13:0] _T_81796; // @[Modules.scala 166:64:@28896.4]
  wire [13:0] buffer_8_570; // @[Modules.scala 166:64:@28897.4]
  wire [14:0] _T_81798; // @[Modules.scala 166:64:@28899.4]
  wire [13:0] _T_81799; // @[Modules.scala 166:64:@28900.4]
  wire [13:0] buffer_8_571; // @[Modules.scala 166:64:@28901.4]
  wire [14:0] _T_81801; // @[Modules.scala 166:64:@28903.4]
  wire [13:0] _T_81802; // @[Modules.scala 166:64:@28904.4]
  wire [13:0] buffer_8_572; // @[Modules.scala 166:64:@28905.4]
  wire [14:0] _T_81804; // @[Modules.scala 166:64:@28907.4]
  wire [13:0] _T_81805; // @[Modules.scala 166:64:@28908.4]
  wire [13:0] buffer_8_573; // @[Modules.scala 166:64:@28909.4]
  wire [14:0] _T_81807; // @[Modules.scala 166:64:@28911.4]
  wire [13:0] _T_81808; // @[Modules.scala 166:64:@28912.4]
  wire [13:0] buffer_8_574; // @[Modules.scala 166:64:@28913.4]
  wire [14:0] _T_81810; // @[Modules.scala 166:64:@28915.4]
  wire [13:0] _T_81811; // @[Modules.scala 166:64:@28916.4]
  wire [13:0] buffer_8_575; // @[Modules.scala 166:64:@28917.4]
  wire [14:0] _T_81813; // @[Modules.scala 166:64:@28919.4]
  wire [13:0] _T_81814; // @[Modules.scala 166:64:@28920.4]
  wire [13:0] buffer_8_576; // @[Modules.scala 166:64:@28921.4]
  wire [14:0] _T_81816; // @[Modules.scala 166:64:@28923.4]
  wire [13:0] _T_81817; // @[Modules.scala 166:64:@28924.4]
  wire [13:0] buffer_8_577; // @[Modules.scala 166:64:@28925.4]
  wire [14:0] _T_81819; // @[Modules.scala 172:66:@28927.4]
  wire [13:0] _T_81820; // @[Modules.scala 172:66:@28928.4]
  wire [13:0] buffer_8_578; // @[Modules.scala 172:66:@28929.4]
  wire [14:0] _T_81822; // @[Modules.scala 166:64:@28931.4]
  wire [13:0] _T_81823; // @[Modules.scala 166:64:@28932.4]
  wire [13:0] buffer_8_579; // @[Modules.scala 166:64:@28933.4]
  wire [14:0] _T_81825; // @[Modules.scala 166:64:@28935.4]
  wire [13:0] _T_81826; // @[Modules.scala 166:64:@28936.4]
  wire [13:0] buffer_8_580; // @[Modules.scala 166:64:@28937.4]
  wire [14:0] _T_81828; // @[Modules.scala 166:64:@28939.4]
  wire [13:0] _T_81829; // @[Modules.scala 166:64:@28940.4]
  wire [13:0] buffer_8_581; // @[Modules.scala 166:64:@28941.4]
  wire [14:0] _T_81831; // @[Modules.scala 166:64:@28943.4]
  wire [13:0] _T_81832; // @[Modules.scala 166:64:@28944.4]
  wire [13:0] buffer_8_582; // @[Modules.scala 166:64:@28945.4]
  wire [14:0] _T_81834; // @[Modules.scala 166:64:@28947.4]
  wire [13:0] _T_81835; // @[Modules.scala 166:64:@28948.4]
  wire [13:0] buffer_8_583; // @[Modules.scala 166:64:@28949.4]
  wire [14:0] _T_81837; // @[Modules.scala 166:64:@28951.4]
  wire [13:0] _T_81838; // @[Modules.scala 166:64:@28952.4]
  wire [13:0] buffer_8_584; // @[Modules.scala 166:64:@28953.4]
  wire [14:0] _T_81840; // @[Modules.scala 166:64:@28955.4]
  wire [13:0] _T_81841; // @[Modules.scala 166:64:@28956.4]
  wire [13:0] buffer_8_585; // @[Modules.scala 166:64:@28957.4]
  wire [14:0] _T_81843; // @[Modules.scala 166:64:@28959.4]
  wire [13:0] _T_81844; // @[Modules.scala 166:64:@28960.4]
  wire [13:0] buffer_8_586; // @[Modules.scala 166:64:@28961.4]
  wire [14:0] _T_81846; // @[Modules.scala 166:64:@28963.4]
  wire [13:0] _T_81847; // @[Modules.scala 166:64:@28964.4]
  wire [13:0] buffer_8_587; // @[Modules.scala 166:64:@28965.4]
  wire [14:0] _T_81849; // @[Modules.scala 166:64:@28967.4]
  wire [13:0] _T_81850; // @[Modules.scala 166:64:@28968.4]
  wire [13:0] buffer_8_588; // @[Modules.scala 166:64:@28969.4]
  wire [14:0] _T_81852; // @[Modules.scala 166:64:@28971.4]
  wire [13:0] _T_81853; // @[Modules.scala 166:64:@28972.4]
  wire [13:0] buffer_8_589; // @[Modules.scala 166:64:@28973.4]
  wire [14:0] _T_81855; // @[Modules.scala 166:64:@28975.4]
  wire [13:0] _T_81856; // @[Modules.scala 166:64:@28976.4]
  wire [13:0] buffer_8_590; // @[Modules.scala 166:64:@28977.4]
  wire [14:0] _T_81858; // @[Modules.scala 166:64:@28979.4]
  wire [13:0] _T_81859; // @[Modules.scala 166:64:@28980.4]
  wire [13:0] buffer_8_591; // @[Modules.scala 166:64:@28981.4]
  wire [14:0] _T_81861; // @[Modules.scala 166:64:@28983.4]
  wire [13:0] _T_81862; // @[Modules.scala 166:64:@28984.4]
  wire [13:0] buffer_8_592; // @[Modules.scala 166:64:@28985.4]
  wire [14:0] _T_81864; // @[Modules.scala 166:64:@28987.4]
  wire [13:0] _T_81865; // @[Modules.scala 166:64:@28988.4]
  wire [13:0] buffer_8_593; // @[Modules.scala 166:64:@28989.4]
  wire [14:0] _T_81867; // @[Modules.scala 166:64:@28991.4]
  wire [13:0] _T_81868; // @[Modules.scala 166:64:@28992.4]
  wire [13:0] buffer_8_594; // @[Modules.scala 166:64:@28993.4]
  wire [14:0] _T_81870; // @[Modules.scala 166:64:@28995.4]
  wire [13:0] _T_81871; // @[Modules.scala 166:64:@28996.4]
  wire [13:0] buffer_8_595; // @[Modules.scala 166:64:@28997.4]
  wire [14:0] _T_81873; // @[Modules.scala 166:64:@28999.4]
  wire [13:0] _T_81874; // @[Modules.scala 166:64:@29000.4]
  wire [13:0] buffer_8_596; // @[Modules.scala 166:64:@29001.4]
  wire [14:0] _T_81876; // @[Modules.scala 166:64:@29003.4]
  wire [13:0] _T_81877; // @[Modules.scala 166:64:@29004.4]
  wire [13:0] buffer_8_597; // @[Modules.scala 166:64:@29005.4]
  wire [14:0] _T_81879; // @[Modules.scala 166:64:@29007.4]
  wire [13:0] _T_81880; // @[Modules.scala 166:64:@29008.4]
  wire [13:0] buffer_8_598; // @[Modules.scala 166:64:@29009.4]
  wire [14:0] _T_81882; // @[Modules.scala 166:64:@29011.4]
  wire [13:0] _T_81883; // @[Modules.scala 166:64:@29012.4]
  wire [13:0] buffer_8_599; // @[Modules.scala 166:64:@29013.4]
  wire [14:0] _T_81885; // @[Modules.scala 166:64:@29015.4]
  wire [13:0] _T_81886; // @[Modules.scala 166:64:@29016.4]
  wire [13:0] buffer_8_600; // @[Modules.scala 166:64:@29017.4]
  wire [14:0] _T_81888; // @[Modules.scala 166:64:@29019.4]
  wire [13:0] _T_81889; // @[Modules.scala 166:64:@29020.4]
  wire [13:0] buffer_8_601; // @[Modules.scala 166:64:@29021.4]
  wire [14:0] _T_81891; // @[Modules.scala 166:64:@29023.4]
  wire [13:0] _T_81892; // @[Modules.scala 166:64:@29024.4]
  wire [13:0] buffer_8_602; // @[Modules.scala 166:64:@29025.4]
  wire [14:0] _T_81894; // @[Modules.scala 166:64:@29027.4]
  wire [13:0] _T_81895; // @[Modules.scala 166:64:@29028.4]
  wire [13:0] buffer_8_603; // @[Modules.scala 166:64:@29029.4]
  wire [14:0] _T_81897; // @[Modules.scala 166:64:@29031.4]
  wire [13:0] _T_81898; // @[Modules.scala 166:64:@29032.4]
  wire [13:0] buffer_8_604; // @[Modules.scala 166:64:@29033.4]
  wire [14:0] _T_81900; // @[Modules.scala 166:64:@29035.4]
  wire [13:0] _T_81901; // @[Modules.scala 166:64:@29036.4]
  wire [13:0] buffer_8_605; // @[Modules.scala 166:64:@29037.4]
  wire [14:0] _T_81903; // @[Modules.scala 166:64:@29039.4]
  wire [13:0] _T_81904; // @[Modules.scala 166:64:@29040.4]
  wire [13:0] buffer_8_606; // @[Modules.scala 166:64:@29041.4]
  wire [14:0] _T_81906; // @[Modules.scala 172:66:@29043.4]
  wire [13:0] _T_81907; // @[Modules.scala 172:66:@29044.4]
  wire [13:0] buffer_8_607; // @[Modules.scala 172:66:@29045.4]
  wire [14:0] _T_81909; // @[Modules.scala 160:64:@29047.4]
  wire [13:0] _T_81910; // @[Modules.scala 160:64:@29048.4]
  wire [13:0] buffer_8_608; // @[Modules.scala 160:64:@29049.4]
  wire [14:0] _T_81912; // @[Modules.scala 160:64:@29051.4]
  wire [13:0] _T_81913; // @[Modules.scala 160:64:@29052.4]
  wire [13:0] buffer_8_609; // @[Modules.scala 160:64:@29053.4]
  wire [14:0] _T_81915; // @[Modules.scala 160:64:@29055.4]
  wire [13:0] _T_81916; // @[Modules.scala 160:64:@29056.4]
  wire [13:0] buffer_8_610; // @[Modules.scala 160:64:@29057.4]
  wire [14:0] _T_81918; // @[Modules.scala 160:64:@29059.4]
  wire [13:0] _T_81919; // @[Modules.scala 160:64:@29060.4]
  wire [13:0] buffer_8_611; // @[Modules.scala 160:64:@29061.4]
  wire [14:0] _T_81921; // @[Modules.scala 160:64:@29063.4]
  wire [13:0] _T_81922; // @[Modules.scala 160:64:@29064.4]
  wire [13:0] buffer_8_612; // @[Modules.scala 160:64:@29065.4]
  wire [14:0] _T_81924; // @[Modules.scala 166:64:@29067.4]
  wire [13:0] _T_81925; // @[Modules.scala 166:64:@29068.4]
  wire [13:0] buffer_8_613; // @[Modules.scala 166:64:@29069.4]
  wire [14:0] _T_81927; // @[Modules.scala 166:64:@29071.4]
  wire [13:0] _T_81928; // @[Modules.scala 166:64:@29072.4]
  wire [13:0] buffer_8_614; // @[Modules.scala 166:64:@29073.4]
  wire [14:0] _T_81930; // @[Modules.scala 160:64:@29075.4]
  wire [13:0] _T_81931; // @[Modules.scala 160:64:@29076.4]
  wire [13:0] buffer_8_615; // @[Modules.scala 160:64:@29077.4]
  wire [14:0] _T_81933; // @[Modules.scala 172:66:@29079.4]
  wire [13:0] _T_81934; // @[Modules.scala 172:66:@29080.4]
  wire [13:0] buffer_8_616; // @[Modules.scala 172:66:@29081.4]
  wire [5:0] _GEN_633; // @[Modules.scala 143:103:@29270.4]
  wire [6:0] _T_81961; // @[Modules.scala 143:103:@29270.4]
  wire [5:0] _T_81962; // @[Modules.scala 143:103:@29271.4]
  wire [5:0] _T_81963; // @[Modules.scala 143:103:@29272.4]
  wire [6:0] _T_81982; // @[Modules.scala 143:103:@29288.4]
  wire [5:0] _T_81983; // @[Modules.scala 143:103:@29289.4]
  wire [5:0] _T_81984; // @[Modules.scala 143:103:@29290.4]
  wire [6:0] _T_81989; // @[Modules.scala 143:103:@29294.4]
  wire [5:0] _T_81990; // @[Modules.scala 143:103:@29295.4]
  wire [5:0] _T_81991; // @[Modules.scala 143:103:@29296.4]
  wire [6:0] _T_81996; // @[Modules.scala 143:103:@29300.4]
  wire [5:0] _T_81997; // @[Modules.scala 143:103:@29301.4]
  wire [5:0] _T_81998; // @[Modules.scala 143:103:@29302.4]
  wire [6:0] _T_82010; // @[Modules.scala 143:103:@29312.4]
  wire [5:0] _T_82011; // @[Modules.scala 143:103:@29313.4]
  wire [5:0] _T_82012; // @[Modules.scala 143:103:@29314.4]
  wire [6:0] _T_82038; // @[Modules.scala 143:103:@29336.4]
  wire [5:0] _T_82039; // @[Modules.scala 143:103:@29337.4]
  wire [5:0] _T_82040; // @[Modules.scala 143:103:@29338.4]
  wire [6:0] _T_82094; // @[Modules.scala 143:103:@29384.4]
  wire [5:0] _T_82095; // @[Modules.scala 143:103:@29385.4]
  wire [5:0] _T_82096; // @[Modules.scala 143:103:@29386.4]
  wire [6:0] _T_82143; // @[Modules.scala 143:103:@29426.4]
  wire [5:0] _T_82144; // @[Modules.scala 143:103:@29427.4]
  wire [5:0] _T_82145; // @[Modules.scala 143:103:@29428.4]
  wire [6:0] _T_82199; // @[Modules.scala 143:103:@29474.4]
  wire [5:0] _T_82200; // @[Modules.scala 143:103:@29475.4]
  wire [5:0] _T_82201; // @[Modules.scala 143:103:@29476.4]
  wire [5:0] _GEN_637; // @[Modules.scala 143:103:@29480.4]
  wire [6:0] _T_82206; // @[Modules.scala 143:103:@29480.4]
  wire [5:0] _T_82207; // @[Modules.scala 143:103:@29481.4]
  wire [5:0] _T_82208; // @[Modules.scala 143:103:@29482.4]
  wire [5:0] _T_82227; // @[Modules.scala 143:103:@29498.4]
  wire [4:0] _T_82228; // @[Modules.scala 143:103:@29499.4]
  wire [4:0] _T_82229; // @[Modules.scala 143:103:@29500.4]
  wire [6:0] _T_82234; // @[Modules.scala 143:103:@29504.4]
  wire [5:0] _T_82235; // @[Modules.scala 143:103:@29505.4]
  wire [5:0] _T_82236; // @[Modules.scala 143:103:@29506.4]
  wire [5:0] _GEN_639; // @[Modules.scala 143:103:@29510.4]
  wire [6:0] _T_82241; // @[Modules.scala 143:103:@29510.4]
  wire [5:0] _T_82242; // @[Modules.scala 143:103:@29511.4]
  wire [5:0] _T_82243; // @[Modules.scala 143:103:@29512.4]
  wire [6:0] _T_82262; // @[Modules.scala 143:103:@29528.4]
  wire [5:0] _T_82263; // @[Modules.scala 143:103:@29529.4]
  wire [5:0] _T_82264; // @[Modules.scala 143:103:@29530.4]
  wire [5:0] _GEN_642; // @[Modules.scala 143:103:@29558.4]
  wire [6:0] _T_82297; // @[Modules.scala 143:103:@29558.4]
  wire [5:0] _T_82298; // @[Modules.scala 143:103:@29559.4]
  wire [5:0] _T_82299; // @[Modules.scala 143:103:@29560.4]
  wire [6:0] _T_82325; // @[Modules.scala 143:103:@29582.4]
  wire [5:0] _T_82326; // @[Modules.scala 143:103:@29583.4]
  wire [5:0] _T_82327; // @[Modules.scala 143:103:@29584.4]
  wire [6:0] _T_82353; // @[Modules.scala 143:103:@29606.4]
  wire [5:0] _T_82354; // @[Modules.scala 143:103:@29607.4]
  wire [5:0] _T_82355; // @[Modules.scala 143:103:@29608.4]
  wire [6:0] _T_82360; // @[Modules.scala 143:103:@29612.4]
  wire [5:0] _T_82361; // @[Modules.scala 143:103:@29613.4]
  wire [5:0] _T_82362; // @[Modules.scala 143:103:@29614.4]
  wire [6:0] _T_82381; // @[Modules.scala 143:103:@29630.4]
  wire [5:0] _T_82382; // @[Modules.scala 143:103:@29631.4]
  wire [5:0] _T_82383; // @[Modules.scala 143:103:@29632.4]
  wire [5:0] _GEN_646; // @[Modules.scala 143:103:@29678.4]
  wire [6:0] _T_82437; // @[Modules.scala 143:103:@29678.4]
  wire [5:0] _T_82438; // @[Modules.scala 143:103:@29679.4]
  wire [5:0] _T_82439; // @[Modules.scala 143:103:@29680.4]
  wire [6:0] _T_82451; // @[Modules.scala 143:103:@29690.4]
  wire [5:0] _T_82452; // @[Modules.scala 143:103:@29691.4]
  wire [5:0] _T_82453; // @[Modules.scala 143:103:@29692.4]
  wire [6:0] _T_82458; // @[Modules.scala 143:103:@29696.4]
  wire [5:0] _T_82459; // @[Modules.scala 143:103:@29697.4]
  wire [5:0] _T_82460; // @[Modules.scala 143:103:@29698.4]
  wire [6:0] _T_82465; // @[Modules.scala 143:103:@29702.4]
  wire [5:0] _T_82466; // @[Modules.scala 143:103:@29703.4]
  wire [5:0] _T_82467; // @[Modules.scala 143:103:@29704.4]
  wire [5:0] _T_82479; // @[Modules.scala 143:103:@29714.4]
  wire [4:0] _T_82480; // @[Modules.scala 143:103:@29715.4]
  wire [4:0] _T_82481; // @[Modules.scala 143:103:@29716.4]
  wire [6:0] _T_82486; // @[Modules.scala 143:103:@29720.4]
  wire [5:0] _T_82487; // @[Modules.scala 143:103:@29721.4]
  wire [5:0] _T_82488; // @[Modules.scala 143:103:@29722.4]
  wire [5:0] _T_82528; // @[Modules.scala 143:103:@29756.4]
  wire [4:0] _T_82529; // @[Modules.scala 143:103:@29757.4]
  wire [4:0] _T_82530; // @[Modules.scala 143:103:@29758.4]
  wire [5:0] _T_82535; // @[Modules.scala 143:103:@29762.4]
  wire [4:0] _T_82536; // @[Modules.scala 143:103:@29763.4]
  wire [4:0] _T_82537; // @[Modules.scala 143:103:@29764.4]
  wire [5:0] _T_82542; // @[Modules.scala 143:103:@29768.4]
  wire [4:0] _T_82543; // @[Modules.scala 143:103:@29769.4]
  wire [4:0] _T_82544; // @[Modules.scala 143:103:@29770.4]
  wire [6:0] _T_82570; // @[Modules.scala 143:103:@29792.4]
  wire [5:0] _T_82571; // @[Modules.scala 143:103:@29793.4]
  wire [5:0] _T_82572; // @[Modules.scala 143:103:@29794.4]
  wire [5:0] _GEN_652; // @[Modules.scala 143:103:@29798.4]
  wire [6:0] _T_82577; // @[Modules.scala 143:103:@29798.4]
  wire [5:0] _T_82578; // @[Modules.scala 143:103:@29799.4]
  wire [5:0] _T_82579; // @[Modules.scala 143:103:@29800.4]
  wire [5:0] _T_82619; // @[Modules.scala 143:103:@29834.4]
  wire [4:0] _T_82620; // @[Modules.scala 143:103:@29835.4]
  wire [4:0] _T_82621; // @[Modules.scala 143:103:@29836.4]
  wire [5:0] _T_82654; // @[Modules.scala 143:103:@29864.4]
  wire [4:0] _T_82655; // @[Modules.scala 143:103:@29865.4]
  wire [4:0] _T_82656; // @[Modules.scala 143:103:@29866.4]
  wire [5:0] _T_82661; // @[Modules.scala 143:103:@29870.4]
  wire [4:0] _T_82662; // @[Modules.scala 143:103:@29871.4]
  wire [4:0] _T_82663; // @[Modules.scala 143:103:@29872.4]
  wire [5:0] _T_82668; // @[Modules.scala 143:103:@29876.4]
  wire [4:0] _T_82669; // @[Modules.scala 143:103:@29877.4]
  wire [4:0] _T_82670; // @[Modules.scala 143:103:@29878.4]
  wire [5:0] _GEN_654; // @[Modules.scala 143:103:@29894.4]
  wire [6:0] _T_82689; // @[Modules.scala 143:103:@29894.4]
  wire [5:0] _T_82690; // @[Modules.scala 143:103:@29895.4]
  wire [5:0] _T_82691; // @[Modules.scala 143:103:@29896.4]
  wire [5:0] _T_82731; // @[Modules.scala 143:103:@29930.4]
  wire [4:0] _T_82732; // @[Modules.scala 143:103:@29931.4]
  wire [4:0] _T_82733; // @[Modules.scala 143:103:@29932.4]
  wire [5:0] _GEN_655; // @[Modules.scala 143:103:@29936.4]
  wire [6:0] _T_82738; // @[Modules.scala 143:103:@29936.4]
  wire [5:0] _T_82739; // @[Modules.scala 143:103:@29937.4]
  wire [5:0] _T_82740; // @[Modules.scala 143:103:@29938.4]
  wire [6:0] _T_82780; // @[Modules.scala 143:103:@29972.4]
  wire [5:0] _T_82781; // @[Modules.scala 143:103:@29973.4]
  wire [5:0] _T_82782; // @[Modules.scala 143:103:@29974.4]
  wire [5:0] _T_82787; // @[Modules.scala 143:103:@29978.4]
  wire [4:0] _T_82788; // @[Modules.scala 143:103:@29979.4]
  wire [4:0] _T_82789; // @[Modules.scala 143:103:@29980.4]
  wire [5:0] _GEN_657; // @[Modules.scala 143:103:@29990.4]
  wire [6:0] _T_82801; // @[Modules.scala 143:103:@29990.4]
  wire [5:0] _T_82802; // @[Modules.scala 143:103:@29991.4]
  wire [5:0] _T_82803; // @[Modules.scala 143:103:@29992.4]
  wire [5:0] _GEN_658; // @[Modules.scala 143:103:@29996.4]
  wire [6:0] _T_82808; // @[Modules.scala 143:103:@29996.4]
  wire [5:0] _T_82809; // @[Modules.scala 143:103:@29997.4]
  wire [5:0] _T_82810; // @[Modules.scala 143:103:@29998.4]
  wire [6:0] _T_82815; // @[Modules.scala 143:103:@30002.4]
  wire [5:0] _T_82816; // @[Modules.scala 143:103:@30003.4]
  wire [5:0] _T_82817; // @[Modules.scala 143:103:@30004.4]
  wire [5:0] _T_82829; // @[Modules.scala 143:103:@30014.4]
  wire [4:0] _T_82830; // @[Modules.scala 143:103:@30015.4]
  wire [4:0] _T_82831; // @[Modules.scala 143:103:@30016.4]
  wire [5:0] _T_82836; // @[Modules.scala 143:103:@30020.4]
  wire [4:0] _T_82837; // @[Modules.scala 143:103:@30021.4]
  wire [4:0] _T_82838; // @[Modules.scala 143:103:@30022.4]
  wire [5:0] _T_82878; // @[Modules.scala 143:103:@30056.4]
  wire [4:0] _T_82879; // @[Modules.scala 143:103:@30057.4]
  wire [4:0] _T_82880; // @[Modules.scala 143:103:@30058.4]
  wire [6:0] _T_82885; // @[Modules.scala 143:103:@30062.4]
  wire [5:0] _T_82886; // @[Modules.scala 143:103:@30063.4]
  wire [5:0] _T_82887; // @[Modules.scala 143:103:@30064.4]
  wire [6:0] _T_82920; // @[Modules.scala 143:103:@30092.4]
  wire [5:0] _T_82921; // @[Modules.scala 143:103:@30093.4]
  wire [5:0] _T_82922; // @[Modules.scala 143:103:@30094.4]
  wire [5:0] _T_82927; // @[Modules.scala 143:103:@30098.4]
  wire [4:0] _T_82928; // @[Modules.scala 143:103:@30099.4]
  wire [4:0] _T_82929; // @[Modules.scala 143:103:@30100.4]
  wire [5:0] _T_82934; // @[Modules.scala 143:103:@30104.4]
  wire [4:0] _T_82935; // @[Modules.scala 143:103:@30105.4]
  wire [4:0] _T_82936; // @[Modules.scala 143:103:@30106.4]
  wire [5:0] _T_82962; // @[Modules.scala 143:103:@30128.4]
  wire [4:0] _T_82963; // @[Modules.scala 143:103:@30129.4]
  wire [4:0] _T_82964; // @[Modules.scala 143:103:@30130.4]
  wire [6:0] _T_83011; // @[Modules.scala 143:103:@30170.4]
  wire [5:0] _T_83012; // @[Modules.scala 143:103:@30171.4]
  wire [5:0] _T_83013; // @[Modules.scala 143:103:@30172.4]
  wire [5:0] _T_83018; // @[Modules.scala 143:103:@30176.4]
  wire [4:0] _T_83019; // @[Modules.scala 143:103:@30177.4]
  wire [4:0] _T_83020; // @[Modules.scala 143:103:@30178.4]
  wire [5:0] _T_83039; // @[Modules.scala 143:103:@30194.4]
  wire [4:0] _T_83040; // @[Modules.scala 143:103:@30195.4]
  wire [4:0] _T_83041; // @[Modules.scala 143:103:@30196.4]
  wire [6:0] _T_83088; // @[Modules.scala 143:103:@30236.4]
  wire [5:0] _T_83089; // @[Modules.scala 143:103:@30237.4]
  wire [5:0] _T_83090; // @[Modules.scala 143:103:@30238.4]
  wire [6:0] _T_83095; // @[Modules.scala 143:103:@30242.4]
  wire [5:0] _T_83096; // @[Modules.scala 143:103:@30243.4]
  wire [5:0] _T_83097; // @[Modules.scala 143:103:@30244.4]
  wire [6:0] _T_83102; // @[Modules.scala 143:103:@30248.4]
  wire [5:0] _T_83103; // @[Modules.scala 143:103:@30249.4]
  wire [5:0] _T_83104; // @[Modules.scala 143:103:@30250.4]
  wire [5:0] _T_83116; // @[Modules.scala 143:103:@30260.4]
  wire [4:0] _T_83117; // @[Modules.scala 143:103:@30261.4]
  wire [4:0] _T_83118; // @[Modules.scala 143:103:@30262.4]
  wire [6:0] _T_83123; // @[Modules.scala 143:103:@30266.4]
  wire [5:0] _T_83124; // @[Modules.scala 143:103:@30267.4]
  wire [5:0] _T_83125; // @[Modules.scala 143:103:@30268.4]
  wire [6:0] _T_83144; // @[Modules.scala 143:103:@30284.4]
  wire [5:0] _T_83145; // @[Modules.scala 143:103:@30285.4]
  wire [5:0] _T_83146; // @[Modules.scala 143:103:@30286.4]
  wire [6:0] _T_83151; // @[Modules.scala 143:103:@30290.4]
  wire [5:0] _T_83152; // @[Modules.scala 143:103:@30291.4]
  wire [5:0] _T_83153; // @[Modules.scala 143:103:@30292.4]
  wire [6:0] _T_83165; // @[Modules.scala 143:103:@30302.4]
  wire [5:0] _T_83166; // @[Modules.scala 143:103:@30303.4]
  wire [5:0] _T_83167; // @[Modules.scala 143:103:@30304.4]
  wire [6:0] _T_83179; // @[Modules.scala 143:103:@30314.4]
  wire [5:0] _T_83180; // @[Modules.scala 143:103:@30315.4]
  wire [5:0] _T_83181; // @[Modules.scala 143:103:@30316.4]
  wire [5:0] _T_83183; // @[Modules.scala 143:74:@30318.4]
  wire [6:0] _T_83186; // @[Modules.scala 143:103:@30320.4]
  wire [5:0] _T_83187; // @[Modules.scala 143:103:@30321.4]
  wire [5:0] _T_83188; // @[Modules.scala 143:103:@30322.4]
  wire [5:0] _GEN_664; // @[Modules.scala 143:103:@30326.4]
  wire [6:0] _T_83193; // @[Modules.scala 143:103:@30326.4]
  wire [5:0] _T_83194; // @[Modules.scala 143:103:@30327.4]
  wire [5:0] _T_83195; // @[Modules.scala 143:103:@30328.4]
  wire [6:0] _T_83207; // @[Modules.scala 143:103:@30338.4]
  wire [5:0] _T_83208; // @[Modules.scala 143:103:@30339.4]
  wire [5:0] _T_83209; // @[Modules.scala 143:103:@30340.4]
  wire [5:0] _GEN_665; // @[Modules.scala 143:103:@30344.4]
  wire [6:0] _T_83214; // @[Modules.scala 143:103:@30344.4]
  wire [5:0] _T_83215; // @[Modules.scala 143:103:@30345.4]
  wire [5:0] _T_83216; // @[Modules.scala 143:103:@30346.4]
  wire [6:0] _T_83256; // @[Modules.scala 143:103:@30380.4]
  wire [5:0] _T_83257; // @[Modules.scala 143:103:@30381.4]
  wire [5:0] _T_83258; // @[Modules.scala 143:103:@30382.4]
  wire [5:0] _T_83284; // @[Modules.scala 143:103:@30404.4]
  wire [4:0] _T_83285; // @[Modules.scala 143:103:@30405.4]
  wire [4:0] _T_83286; // @[Modules.scala 143:103:@30406.4]
  wire [6:0] _T_83340; // @[Modules.scala 143:103:@30452.4]
  wire [5:0] _T_83341; // @[Modules.scala 143:103:@30453.4]
  wire [5:0] _T_83342; // @[Modules.scala 143:103:@30454.4]
  wire [6:0] _T_83347; // @[Modules.scala 143:103:@30458.4]
  wire [5:0] _T_83348; // @[Modules.scala 143:103:@30459.4]
  wire [5:0] _T_83349; // @[Modules.scala 143:103:@30460.4]
  wire [6:0] _T_83354; // @[Modules.scala 143:103:@30464.4]
  wire [5:0] _T_83355; // @[Modules.scala 143:103:@30465.4]
  wire [5:0] _T_83356; // @[Modules.scala 143:103:@30466.4]
  wire [5:0] _GEN_668; // @[Modules.scala 143:103:@30470.4]
  wire [6:0] _T_83361; // @[Modules.scala 143:103:@30470.4]
  wire [5:0] _T_83362; // @[Modules.scala 143:103:@30471.4]
  wire [5:0] _T_83363; // @[Modules.scala 143:103:@30472.4]
  wire [5:0] _T_83375; // @[Modules.scala 143:103:@30482.4]
  wire [4:0] _T_83376; // @[Modules.scala 143:103:@30483.4]
  wire [4:0] _T_83377; // @[Modules.scala 143:103:@30484.4]
  wire [5:0] _GEN_669; // @[Modules.scala 143:103:@30494.4]
  wire [6:0] _T_83389; // @[Modules.scala 143:103:@30494.4]
  wire [5:0] _T_83390; // @[Modules.scala 143:103:@30495.4]
  wire [5:0] _T_83391; // @[Modules.scala 143:103:@30496.4]
  wire [6:0] _T_83438; // @[Modules.scala 143:103:@30536.4]
  wire [5:0] _T_83439; // @[Modules.scala 143:103:@30537.4]
  wire [5:0] _T_83440; // @[Modules.scala 143:103:@30538.4]
  wire [5:0] _GEN_672; // @[Modules.scala 143:103:@30542.4]
  wire [6:0] _T_83445; // @[Modules.scala 143:103:@30542.4]
  wire [5:0] _T_83446; // @[Modules.scala 143:103:@30543.4]
  wire [5:0] _T_83447; // @[Modules.scala 143:103:@30544.4]
  wire [5:0] _GEN_673; // @[Modules.scala 143:103:@30566.4]
  wire [6:0] _T_83473; // @[Modules.scala 143:103:@30566.4]
  wire [5:0] _T_83474; // @[Modules.scala 143:103:@30567.4]
  wire [5:0] _T_83475; // @[Modules.scala 143:103:@30568.4]
  wire [6:0] _T_83501; // @[Modules.scala 143:103:@30590.4]
  wire [5:0] _T_83502; // @[Modules.scala 143:103:@30591.4]
  wire [5:0] _T_83503; // @[Modules.scala 143:103:@30592.4]
  wire [6:0] _T_83508; // @[Modules.scala 143:103:@30596.4]
  wire [5:0] _T_83509; // @[Modules.scala 143:103:@30597.4]
  wire [5:0] _T_83510; // @[Modules.scala 143:103:@30598.4]
  wire [6:0] _T_83515; // @[Modules.scala 143:103:@30602.4]
  wire [5:0] _T_83516; // @[Modules.scala 143:103:@30603.4]
  wire [5:0] _T_83517; // @[Modules.scala 143:103:@30604.4]
  wire [5:0] _T_83543; // @[Modules.scala 143:103:@30626.4]
  wire [4:0] _T_83544; // @[Modules.scala 143:103:@30627.4]
  wire [4:0] _T_83545; // @[Modules.scala 143:103:@30628.4]
  wire [6:0] _T_83550; // @[Modules.scala 143:103:@30632.4]
  wire [5:0] _T_83551; // @[Modules.scala 143:103:@30633.4]
  wire [5:0] _T_83552; // @[Modules.scala 143:103:@30634.4]
  wire [5:0] _GEN_676; // @[Modules.scala 143:103:@30638.4]
  wire [6:0] _T_83557; // @[Modules.scala 143:103:@30638.4]
  wire [5:0] _T_83558; // @[Modules.scala 143:103:@30639.4]
  wire [5:0] _T_83559; // @[Modules.scala 143:103:@30640.4]
  wire [6:0] _T_83585; // @[Modules.scala 143:103:@30662.4]
  wire [5:0] _T_83586; // @[Modules.scala 143:103:@30663.4]
  wire [5:0] _T_83587; // @[Modules.scala 143:103:@30664.4]
  wire [5:0] _T_83599; // @[Modules.scala 143:103:@30674.4]
  wire [4:0] _T_83600; // @[Modules.scala 143:103:@30675.4]
  wire [4:0] _T_83601; // @[Modules.scala 143:103:@30676.4]
  wire [6:0] _T_83606; // @[Modules.scala 143:103:@30680.4]
  wire [5:0] _T_83607; // @[Modules.scala 143:103:@30681.4]
  wire [5:0] _T_83608; // @[Modules.scala 143:103:@30682.4]
  wire [5:0] _GEN_679; // @[Modules.scala 143:103:@30698.4]
  wire [6:0] _T_83627; // @[Modules.scala 143:103:@30698.4]
  wire [5:0] _T_83628; // @[Modules.scala 143:103:@30699.4]
  wire [5:0] _T_83629; // @[Modules.scala 143:103:@30700.4]
  wire [6:0] _T_83634; // @[Modules.scala 143:103:@30704.4]
  wire [5:0] _T_83635; // @[Modules.scala 143:103:@30705.4]
  wire [5:0] _T_83636; // @[Modules.scala 143:103:@30706.4]
  wire [6:0] _T_83641; // @[Modules.scala 143:103:@30710.4]
  wire [5:0] _T_83642; // @[Modules.scala 143:103:@30711.4]
  wire [5:0] _T_83643; // @[Modules.scala 143:103:@30712.4]
  wire [6:0] _T_83655; // @[Modules.scala 143:103:@30722.4]
  wire [5:0] _T_83656; // @[Modules.scala 143:103:@30723.4]
  wire [5:0] _T_83657; // @[Modules.scala 143:103:@30724.4]
  wire [6:0] _T_83662; // @[Modules.scala 143:103:@30728.4]
  wire [5:0] _T_83663; // @[Modules.scala 143:103:@30729.4]
  wire [5:0] _T_83664; // @[Modules.scala 143:103:@30730.4]
  wire [6:0] _T_83669; // @[Modules.scala 143:103:@30734.4]
  wire [5:0] _T_83670; // @[Modules.scala 143:103:@30735.4]
  wire [5:0] _T_83671; // @[Modules.scala 143:103:@30736.4]
  wire [5:0] _T_83676; // @[Modules.scala 143:103:@30740.4]
  wire [4:0] _T_83677; // @[Modules.scala 143:103:@30741.4]
  wire [4:0] _T_83678; // @[Modules.scala 143:103:@30742.4]
  wire [6:0] _T_83697; // @[Modules.scala 143:103:@30758.4]
  wire [5:0] _T_83698; // @[Modules.scala 143:103:@30759.4]
  wire [5:0] _T_83699; // @[Modules.scala 143:103:@30760.4]
  wire [5:0] _T_83753; // @[Modules.scala 143:103:@30806.4]
  wire [4:0] _T_83754; // @[Modules.scala 143:103:@30807.4]
  wire [4:0] _T_83755; // @[Modules.scala 143:103:@30808.4]
  wire [6:0] _T_83760; // @[Modules.scala 143:103:@30812.4]
  wire [5:0] _T_83761; // @[Modules.scala 143:103:@30813.4]
  wire [5:0] _T_83762; // @[Modules.scala 143:103:@30814.4]
  wire [6:0] _T_83781; // @[Modules.scala 143:103:@30830.4]
  wire [5:0] _T_83782; // @[Modules.scala 143:103:@30831.4]
  wire [5:0] _T_83783; // @[Modules.scala 143:103:@30832.4]
  wire [5:0] _GEN_686; // @[Modules.scala 143:103:@30854.4]
  wire [6:0] _T_83809; // @[Modules.scala 143:103:@30854.4]
  wire [5:0] _T_83810; // @[Modules.scala 143:103:@30855.4]
  wire [5:0] _T_83811; // @[Modules.scala 143:103:@30856.4]
  wire [6:0] _T_83816; // @[Modules.scala 143:103:@30860.4]
  wire [5:0] _T_83817; // @[Modules.scala 143:103:@30861.4]
  wire [5:0] _T_83818; // @[Modules.scala 143:103:@30862.4]
  wire [6:0] _T_83837; // @[Modules.scala 143:103:@30878.4]
  wire [5:0] _T_83838; // @[Modules.scala 143:103:@30879.4]
  wire [5:0] _T_83839; // @[Modules.scala 143:103:@30880.4]
  wire [6:0] _T_83858; // @[Modules.scala 143:103:@30896.4]
  wire [5:0] _T_83859; // @[Modules.scala 143:103:@30897.4]
  wire [5:0] _T_83860; // @[Modules.scala 143:103:@30898.4]
  wire [6:0] _T_83865; // @[Modules.scala 143:103:@30902.4]
  wire [5:0] _T_83866; // @[Modules.scala 143:103:@30903.4]
  wire [5:0] _T_83867; // @[Modules.scala 143:103:@30904.4]
  wire [5:0] _GEN_689; // @[Modules.scala 143:103:@30908.4]
  wire [6:0] _T_83872; // @[Modules.scala 143:103:@30908.4]
  wire [5:0] _T_83873; // @[Modules.scala 143:103:@30909.4]
  wire [5:0] _T_83874; // @[Modules.scala 143:103:@30910.4]
  wire [5:0] _GEN_690; // @[Modules.scala 143:103:@30920.4]
  wire [6:0] _T_83886; // @[Modules.scala 143:103:@30920.4]
  wire [5:0] _T_83887; // @[Modules.scala 143:103:@30921.4]
  wire [5:0] _T_83888; // @[Modules.scala 143:103:@30922.4]
  wire [5:0] _T_83900; // @[Modules.scala 143:103:@30932.4]
  wire [4:0] _T_83901; // @[Modules.scala 143:103:@30933.4]
  wire [4:0] _T_83902; // @[Modules.scala 143:103:@30934.4]
  wire [6:0] _T_83907; // @[Modules.scala 143:103:@30938.4]
  wire [5:0] _T_83908; // @[Modules.scala 143:103:@30939.4]
  wire [5:0] _T_83909; // @[Modules.scala 143:103:@30940.4]
  wire [6:0] _T_83984; // @[Modules.scala 143:103:@31004.4]
  wire [5:0] _T_83985; // @[Modules.scala 143:103:@31005.4]
  wire [5:0] _T_83986; // @[Modules.scala 143:103:@31006.4]
  wire [5:0] _T_84012; // @[Modules.scala 143:103:@31028.4]
  wire [4:0] _T_84013; // @[Modules.scala 143:103:@31029.4]
  wire [4:0] _T_84014; // @[Modules.scala 143:103:@31030.4]
  wire [5:0] _T_84019; // @[Modules.scala 143:103:@31034.4]
  wire [4:0] _T_84020; // @[Modules.scala 143:103:@31035.4]
  wire [4:0] _T_84021; // @[Modules.scala 143:103:@31036.4]
  wire [5:0] _T_84026; // @[Modules.scala 143:103:@31040.4]
  wire [4:0] _T_84027; // @[Modules.scala 143:103:@31041.4]
  wire [4:0] _T_84028; // @[Modules.scala 143:103:@31042.4]
  wire [5:0] _T_84033; // @[Modules.scala 143:103:@31046.4]
  wire [4:0] _T_84034; // @[Modules.scala 143:103:@31047.4]
  wire [4:0] _T_84035; // @[Modules.scala 143:103:@31048.4]
  wire [5:0] _T_84040; // @[Modules.scala 143:103:@31052.4]
  wire [4:0] _T_84041; // @[Modules.scala 143:103:@31053.4]
  wire [4:0] _T_84042; // @[Modules.scala 143:103:@31054.4]
  wire [5:0] _T_84047; // @[Modules.scala 143:103:@31058.4]
  wire [4:0] _T_84048; // @[Modules.scala 143:103:@31059.4]
  wire [4:0] _T_84049; // @[Modules.scala 143:103:@31060.4]
  wire [5:0] _T_84075; // @[Modules.scala 143:103:@31082.4]
  wire [4:0] _T_84076; // @[Modules.scala 143:103:@31083.4]
  wire [4:0] _T_84077; // @[Modules.scala 143:103:@31084.4]
  wire [5:0] _T_84089; // @[Modules.scala 143:103:@31094.4]
  wire [4:0] _T_84090; // @[Modules.scala 143:103:@31095.4]
  wire [4:0] _T_84091; // @[Modules.scala 143:103:@31096.4]
  wire [5:0] _T_84103; // @[Modules.scala 143:103:@31106.4]
  wire [4:0] _T_84104; // @[Modules.scala 143:103:@31107.4]
  wire [4:0] _T_84105; // @[Modules.scala 143:103:@31108.4]
  wire [5:0] _T_84110; // @[Modules.scala 143:103:@31112.4]
  wire [4:0] _T_84111; // @[Modules.scala 143:103:@31113.4]
  wire [4:0] _T_84112; // @[Modules.scala 143:103:@31114.4]
  wire [5:0] _T_84117; // @[Modules.scala 143:103:@31118.4]
  wire [4:0] _T_84118; // @[Modules.scala 143:103:@31119.4]
  wire [4:0] _T_84119; // @[Modules.scala 143:103:@31120.4]
  wire [5:0] _GEN_693; // @[Modules.scala 143:103:@31124.4]
  wire [6:0] _T_84124; // @[Modules.scala 143:103:@31124.4]
  wire [5:0] _T_84125; // @[Modules.scala 143:103:@31125.4]
  wire [5:0] _T_84126; // @[Modules.scala 143:103:@31126.4]
  wire [5:0] _T_84131; // @[Modules.scala 143:103:@31130.4]
  wire [4:0] _T_84132; // @[Modules.scala 143:103:@31131.4]
  wire [4:0] _T_84133; // @[Modules.scala 143:103:@31132.4]
  wire [13:0] buffer_9_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84137; // @[Modules.scala 160:64:@31138.4]
  wire [13:0] _T_84138; // @[Modules.scala 160:64:@31139.4]
  wire [13:0] buffer_9_315; // @[Modules.scala 160:64:@31140.4]
  wire [13:0] buffer_9_6; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_7; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84143; // @[Modules.scala 160:64:@31146.4]
  wire [13:0] _T_84144; // @[Modules.scala 160:64:@31147.4]
  wire [13:0] buffer_9_317; // @[Modules.scala 160:64:@31148.4]
  wire [13:0] buffer_9_8; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84146; // @[Modules.scala 160:64:@31150.4]
  wire [13:0] _T_84147; // @[Modules.scala 160:64:@31151.4]
  wire [13:0] buffer_9_318; // @[Modules.scala 160:64:@31152.4]
  wire [13:0] buffer_9_10; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84149; // @[Modules.scala 160:64:@31154.4]
  wire [13:0] _T_84150; // @[Modules.scala 160:64:@31155.4]
  wire [13:0] buffer_9_319; // @[Modules.scala 160:64:@31156.4]
  wire [14:0] _T_84152; // @[Modules.scala 160:64:@31158.4]
  wire [13:0] _T_84153; // @[Modules.scala 160:64:@31159.4]
  wire [13:0] buffer_9_320; // @[Modules.scala 160:64:@31160.4]
  wire [13:0] buffer_9_14; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84155; // @[Modules.scala 160:64:@31162.4]
  wire [13:0] _T_84156; // @[Modules.scala 160:64:@31163.4]
  wire [13:0] buffer_9_321; // @[Modules.scala 160:64:@31164.4]
  wire [14:0] _T_84158; // @[Modules.scala 160:64:@31166.4]
  wire [13:0] _T_84159; // @[Modules.scala 160:64:@31167.4]
  wire [13:0] buffer_9_322; // @[Modules.scala 160:64:@31168.4]
  wire [14:0] _T_84161; // @[Modules.scala 160:64:@31170.4]
  wire [13:0] _T_84162; // @[Modules.scala 160:64:@31171.4]
  wire [13:0] buffer_9_323; // @[Modules.scala 160:64:@31172.4]
  wire [14:0] _T_84164; // @[Modules.scala 160:64:@31174.4]
  wire [13:0] _T_84165; // @[Modules.scala 160:64:@31175.4]
  wire [13:0] buffer_9_324; // @[Modules.scala 160:64:@31176.4]
  wire [13:0] buffer_9_22; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84167; // @[Modules.scala 160:64:@31178.4]
  wire [13:0] _T_84168; // @[Modules.scala 160:64:@31179.4]
  wire [13:0] buffer_9_325; // @[Modules.scala 160:64:@31180.4]
  wire [14:0] _T_84170; // @[Modules.scala 160:64:@31182.4]
  wire [13:0] _T_84171; // @[Modules.scala 160:64:@31183.4]
  wire [13:0] buffer_9_326; // @[Modules.scala 160:64:@31184.4]
  wire [14:0] _T_84173; // @[Modules.scala 160:64:@31186.4]
  wire [13:0] _T_84174; // @[Modules.scala 160:64:@31187.4]
  wire [13:0] buffer_9_327; // @[Modules.scala 160:64:@31188.4]
  wire [13:0] buffer_9_29; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84176; // @[Modules.scala 160:64:@31190.4]
  wire [13:0] _T_84177; // @[Modules.scala 160:64:@31191.4]
  wire [13:0] buffer_9_328; // @[Modules.scala 160:64:@31192.4]
  wire [14:0] _T_84179; // @[Modules.scala 160:64:@31194.4]
  wire [13:0] _T_84180; // @[Modules.scala 160:64:@31195.4]
  wire [13:0] buffer_9_329; // @[Modules.scala 160:64:@31196.4]
  wire [14:0] _T_84182; // @[Modules.scala 160:64:@31198.4]
  wire [13:0] _T_84183; // @[Modules.scala 160:64:@31199.4]
  wire [13:0] buffer_9_330; // @[Modules.scala 160:64:@31200.4]
  wire [14:0] _T_84185; // @[Modules.scala 160:64:@31202.4]
  wire [13:0] _T_84186; // @[Modules.scala 160:64:@31203.4]
  wire [13:0] buffer_9_331; // @[Modules.scala 160:64:@31204.4]
  wire [13:0] buffer_9_37; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84188; // @[Modules.scala 160:64:@31206.4]
  wire [13:0] _T_84189; // @[Modules.scala 160:64:@31207.4]
  wire [13:0] buffer_9_332; // @[Modules.scala 160:64:@31208.4]
  wire [13:0] buffer_9_38; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84191; // @[Modules.scala 160:64:@31210.4]
  wire [13:0] _T_84192; // @[Modules.scala 160:64:@31211.4]
  wire [13:0] buffer_9_333; // @[Modules.scala 160:64:@31212.4]
  wire [13:0] buffer_9_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84194; // @[Modules.scala 160:64:@31214.4]
  wire [13:0] _T_84195; // @[Modules.scala 160:64:@31215.4]
  wire [13:0] buffer_9_334; // @[Modules.scala 160:64:@31216.4]
  wire [13:0] buffer_9_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84197; // @[Modules.scala 160:64:@31218.4]
  wire [13:0] _T_84198; // @[Modules.scala 160:64:@31219.4]
  wire [13:0] buffer_9_335; // @[Modules.scala 160:64:@31220.4]
  wire [13:0] buffer_9_46; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84203; // @[Modules.scala 160:64:@31226.4]
  wire [13:0] _T_84204; // @[Modules.scala 160:64:@31227.4]
  wire [13:0] buffer_9_337; // @[Modules.scala 160:64:@31228.4]
  wire [14:0] _T_84206; // @[Modules.scala 160:64:@31230.4]
  wire [13:0] _T_84207; // @[Modules.scala 160:64:@31231.4]
  wire [13:0] buffer_9_338; // @[Modules.scala 160:64:@31232.4]
  wire [13:0] buffer_9_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84209; // @[Modules.scala 160:64:@31234.4]
  wire [13:0] _T_84210; // @[Modules.scala 160:64:@31235.4]
  wire [13:0] buffer_9_339; // @[Modules.scala 160:64:@31236.4]
  wire [13:0] buffer_9_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84215; // @[Modules.scala 160:64:@31242.4]
  wire [13:0] _T_84216; // @[Modules.scala 160:64:@31243.4]
  wire [13:0] buffer_9_341; // @[Modules.scala 160:64:@31244.4]
  wire [13:0] buffer_9_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84221; // @[Modules.scala 160:64:@31250.4]
  wire [13:0] _T_84222; // @[Modules.scala 160:64:@31251.4]
  wire [13:0] buffer_9_343; // @[Modules.scala 160:64:@31252.4]
  wire [13:0] buffer_9_60; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84224; // @[Modules.scala 160:64:@31254.4]
  wire [13:0] _T_84225; // @[Modules.scala 160:64:@31255.4]
  wire [13:0] buffer_9_344; // @[Modules.scala 160:64:@31256.4]
  wire [13:0] buffer_9_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84227; // @[Modules.scala 160:64:@31258.4]
  wire [13:0] _T_84228; // @[Modules.scala 160:64:@31259.4]
  wire [13:0] buffer_9_345; // @[Modules.scala 160:64:@31260.4]
  wire [13:0] buffer_9_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84239; // @[Modules.scala 160:64:@31274.4]
  wire [13:0] _T_84240; // @[Modules.scala 160:64:@31275.4]
  wire [13:0] buffer_9_349; // @[Modules.scala 160:64:@31276.4]
  wire [13:0] buffer_9_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84242; // @[Modules.scala 160:64:@31278.4]
  wire [13:0] _T_84243; // @[Modules.scala 160:64:@31279.4]
  wire [13:0] buffer_9_350; // @[Modules.scala 160:64:@31280.4]
  wire [13:0] buffer_9_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84245; // @[Modules.scala 160:64:@31282.4]
  wire [13:0] _T_84246; // @[Modules.scala 160:64:@31283.4]
  wire [13:0] buffer_9_351; // @[Modules.scala 160:64:@31284.4]
  wire [13:0] buffer_9_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84248; // @[Modules.scala 160:64:@31286.4]
  wire [13:0] _T_84249; // @[Modules.scala 160:64:@31287.4]
  wire [13:0] buffer_9_352; // @[Modules.scala 160:64:@31288.4]
  wire [13:0] buffer_9_78; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84251; // @[Modules.scala 160:64:@31290.4]
  wire [13:0] _T_84252; // @[Modules.scala 160:64:@31291.4]
  wire [13:0] buffer_9_353; // @[Modules.scala 160:64:@31292.4]
  wire [14:0] _T_84254; // @[Modules.scala 160:64:@31294.4]
  wire [13:0] _T_84255; // @[Modules.scala 160:64:@31295.4]
  wire [13:0] buffer_9_354; // @[Modules.scala 160:64:@31296.4]
  wire [13:0] buffer_9_84; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84260; // @[Modules.scala 160:64:@31302.4]
  wire [13:0] _T_84261; // @[Modules.scala 160:64:@31303.4]
  wire [13:0] buffer_9_356; // @[Modules.scala 160:64:@31304.4]
  wire [13:0] buffer_9_86; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84263; // @[Modules.scala 160:64:@31306.4]
  wire [13:0] _T_84264; // @[Modules.scala 160:64:@31307.4]
  wire [13:0] buffer_9_357; // @[Modules.scala 160:64:@31308.4]
  wire [14:0] _T_84266; // @[Modules.scala 160:64:@31310.4]
  wire [13:0] _T_84267; // @[Modules.scala 160:64:@31311.4]
  wire [13:0] buffer_9_358; // @[Modules.scala 160:64:@31312.4]
  wire [13:0] buffer_9_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84269; // @[Modules.scala 160:64:@31314.4]
  wire [13:0] _T_84270; // @[Modules.scala 160:64:@31315.4]
  wire [13:0] buffer_9_359; // @[Modules.scala 160:64:@31316.4]
  wire [13:0] buffer_9_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84278; // @[Modules.scala 160:64:@31326.4]
  wire [13:0] _T_84279; // @[Modules.scala 160:64:@31327.4]
  wire [13:0] buffer_9_362; // @[Modules.scala 160:64:@31328.4]
  wire [14:0] _T_84281; // @[Modules.scala 160:64:@31330.4]
  wire [13:0] _T_84282; // @[Modules.scala 160:64:@31331.4]
  wire [13:0] buffer_9_363; // @[Modules.scala 160:64:@31332.4]
  wire [13:0] buffer_9_102; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_103; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84287; // @[Modules.scala 160:64:@31338.4]
  wire [13:0] _T_84288; // @[Modules.scala 160:64:@31339.4]
  wire [13:0] buffer_9_365; // @[Modules.scala 160:64:@31340.4]
  wire [13:0] buffer_9_104; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84290; // @[Modules.scala 160:64:@31342.4]
  wire [13:0] _T_84291; // @[Modules.scala 160:64:@31343.4]
  wire [13:0] buffer_9_366; // @[Modules.scala 160:64:@31344.4]
  wire [13:0] buffer_9_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84293; // @[Modules.scala 160:64:@31346.4]
  wire [13:0] _T_84294; // @[Modules.scala 160:64:@31347.4]
  wire [13:0] buffer_9_367; // @[Modules.scala 160:64:@31348.4]
  wire [14:0] _T_84296; // @[Modules.scala 160:64:@31350.4]
  wire [13:0] _T_84297; // @[Modules.scala 160:64:@31351.4]
  wire [13:0] buffer_9_368; // @[Modules.scala 160:64:@31352.4]
  wire [14:0] _T_84299; // @[Modules.scala 160:64:@31354.4]
  wire [13:0] _T_84300; // @[Modules.scala 160:64:@31355.4]
  wire [13:0] buffer_9_369; // @[Modules.scala 160:64:@31356.4]
  wire [13:0] buffer_9_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84302; // @[Modules.scala 160:64:@31358.4]
  wire [13:0] _T_84303; // @[Modules.scala 160:64:@31359.4]
  wire [13:0] buffer_9_370; // @[Modules.scala 160:64:@31360.4]
  wire [13:0] buffer_9_114; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84305; // @[Modules.scala 160:64:@31362.4]
  wire [13:0] _T_84306; // @[Modules.scala 160:64:@31363.4]
  wire [13:0] buffer_9_371; // @[Modules.scala 160:64:@31364.4]
  wire [14:0] _T_84308; // @[Modules.scala 160:64:@31366.4]
  wire [13:0] _T_84309; // @[Modules.scala 160:64:@31367.4]
  wire [13:0] buffer_9_372; // @[Modules.scala 160:64:@31368.4]
  wire [14:0] _T_84311; // @[Modules.scala 160:64:@31370.4]
  wire [13:0] _T_84312; // @[Modules.scala 160:64:@31371.4]
  wire [13:0] buffer_9_373; // @[Modules.scala 160:64:@31372.4]
  wire [13:0] buffer_9_120; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84314; // @[Modules.scala 160:64:@31374.4]
  wire [13:0] _T_84315; // @[Modules.scala 160:64:@31375.4]
  wire [13:0] buffer_9_374; // @[Modules.scala 160:64:@31376.4]
  wire [13:0] buffer_9_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84317; // @[Modules.scala 160:64:@31378.4]
  wire [13:0] _T_84318; // @[Modules.scala 160:64:@31379.4]
  wire [13:0] buffer_9_375; // @[Modules.scala 160:64:@31380.4]
  wire [13:0] buffer_9_124; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84320; // @[Modules.scala 160:64:@31382.4]
  wire [13:0] _T_84321; // @[Modules.scala 160:64:@31383.4]
  wire [13:0] buffer_9_376; // @[Modules.scala 160:64:@31384.4]
  wire [13:0] buffer_9_127; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84323; // @[Modules.scala 160:64:@31386.4]
  wire [13:0] _T_84324; // @[Modules.scala 160:64:@31387.4]
  wire [13:0] buffer_9_377; // @[Modules.scala 160:64:@31388.4]
  wire [13:0] buffer_9_128; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84326; // @[Modules.scala 160:64:@31390.4]
  wire [13:0] _T_84327; // @[Modules.scala 160:64:@31391.4]
  wire [13:0] buffer_9_378; // @[Modules.scala 160:64:@31392.4]
  wire [14:0] _T_84329; // @[Modules.scala 160:64:@31394.4]
  wire [13:0] _T_84330; // @[Modules.scala 160:64:@31395.4]
  wire [13:0] buffer_9_379; // @[Modules.scala 160:64:@31396.4]
  wire [14:0] _T_84332; // @[Modules.scala 160:64:@31398.4]
  wire [13:0] _T_84333; // @[Modules.scala 160:64:@31399.4]
  wire [13:0] buffer_9_380; // @[Modules.scala 160:64:@31400.4]
  wire [13:0] buffer_9_134; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84335; // @[Modules.scala 160:64:@31402.4]
  wire [13:0] _T_84336; // @[Modules.scala 160:64:@31403.4]
  wire [13:0] buffer_9_381; // @[Modules.scala 160:64:@31404.4]
  wire [13:0] buffer_9_140; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_141; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84344; // @[Modules.scala 160:64:@31414.4]
  wire [13:0] _T_84345; // @[Modules.scala 160:64:@31415.4]
  wire [13:0] buffer_9_384; // @[Modules.scala 160:64:@31416.4]
  wire [13:0] buffer_9_142; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84347; // @[Modules.scala 160:64:@31418.4]
  wire [13:0] _T_84348; // @[Modules.scala 160:64:@31419.4]
  wire [13:0] buffer_9_385; // @[Modules.scala 160:64:@31420.4]
  wire [14:0] _T_84350; // @[Modules.scala 160:64:@31422.4]
  wire [13:0] _T_84351; // @[Modules.scala 160:64:@31423.4]
  wire [13:0] buffer_9_386; // @[Modules.scala 160:64:@31424.4]
  wire [13:0] buffer_9_146; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84353; // @[Modules.scala 160:64:@31426.4]
  wire [13:0] _T_84354; // @[Modules.scala 160:64:@31427.4]
  wire [13:0] buffer_9_387; // @[Modules.scala 160:64:@31428.4]
  wire [14:0] _T_84356; // @[Modules.scala 160:64:@31430.4]
  wire [13:0] _T_84357; // @[Modules.scala 160:64:@31431.4]
  wire [13:0] buffer_9_388; // @[Modules.scala 160:64:@31432.4]
  wire [13:0] buffer_9_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84362; // @[Modules.scala 160:64:@31438.4]
  wire [13:0] _T_84363; // @[Modules.scala 160:64:@31439.4]
  wire [13:0] buffer_9_390; // @[Modules.scala 160:64:@31440.4]
  wire [13:0] buffer_9_154; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84365; // @[Modules.scala 160:64:@31442.4]
  wire [13:0] _T_84366; // @[Modules.scala 160:64:@31443.4]
  wire [13:0] buffer_9_391; // @[Modules.scala 160:64:@31444.4]
  wire [13:0] buffer_9_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84368; // @[Modules.scala 160:64:@31446.4]
  wire [13:0] _T_84369; // @[Modules.scala 160:64:@31447.4]
  wire [13:0] buffer_9_392; // @[Modules.scala 160:64:@31448.4]
  wire [14:0] _T_84371; // @[Modules.scala 160:64:@31450.4]
  wire [13:0] _T_84372; // @[Modules.scala 160:64:@31451.4]
  wire [13:0] buffer_9_393; // @[Modules.scala 160:64:@31452.4]
  wire [13:0] buffer_9_164; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_165; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84380; // @[Modules.scala 160:64:@31462.4]
  wire [13:0] _T_84381; // @[Modules.scala 160:64:@31463.4]
  wire [13:0] buffer_9_396; // @[Modules.scala 160:64:@31464.4]
  wire [13:0] buffer_9_166; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84383; // @[Modules.scala 160:64:@31466.4]
  wire [13:0] _T_84384; // @[Modules.scala 160:64:@31467.4]
  wire [13:0] buffer_9_397; // @[Modules.scala 160:64:@31468.4]
  wire [13:0] buffer_9_168; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84386; // @[Modules.scala 160:64:@31470.4]
  wire [13:0] _T_84387; // @[Modules.scala 160:64:@31471.4]
  wire [13:0] buffer_9_398; // @[Modules.scala 160:64:@31472.4]
  wire [14:0] _T_84389; // @[Modules.scala 160:64:@31474.4]
  wire [13:0] _T_84390; // @[Modules.scala 160:64:@31475.4]
  wire [13:0] buffer_9_399; // @[Modules.scala 160:64:@31476.4]
  wire [13:0] buffer_9_172; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_173; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84392; // @[Modules.scala 160:64:@31478.4]
  wire [13:0] _T_84393; // @[Modules.scala 160:64:@31479.4]
  wire [13:0] buffer_9_400; // @[Modules.scala 160:64:@31480.4]
  wire [13:0] buffer_9_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84395; // @[Modules.scala 160:64:@31482.4]
  wire [13:0] _T_84396; // @[Modules.scala 160:64:@31483.4]
  wire [13:0] buffer_9_401; // @[Modules.scala 160:64:@31484.4]
  wire [13:0] buffer_9_177; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84398; // @[Modules.scala 160:64:@31486.4]
  wire [13:0] _T_84399; // @[Modules.scala 160:64:@31487.4]
  wire [13:0] buffer_9_402; // @[Modules.scala 160:64:@31488.4]
  wire [13:0] buffer_9_178; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_179; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84401; // @[Modules.scala 160:64:@31490.4]
  wire [13:0] _T_84402; // @[Modules.scala 160:64:@31491.4]
  wire [13:0] buffer_9_403; // @[Modules.scala 160:64:@31492.4]
  wire [13:0] buffer_9_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84404; // @[Modules.scala 160:64:@31494.4]
  wire [13:0] _T_84405; // @[Modules.scala 160:64:@31495.4]
  wire [13:0] buffer_9_404; // @[Modules.scala 160:64:@31496.4]
  wire [13:0] buffer_9_182; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84407; // @[Modules.scala 160:64:@31498.4]
  wire [13:0] _T_84408; // @[Modules.scala 160:64:@31499.4]
  wire [13:0] buffer_9_405; // @[Modules.scala 160:64:@31500.4]
  wire [14:0] _T_84410; // @[Modules.scala 160:64:@31502.4]
  wire [13:0] _T_84411; // @[Modules.scala 160:64:@31503.4]
  wire [13:0] buffer_9_406; // @[Modules.scala 160:64:@31504.4]
  wire [14:0] _T_84413; // @[Modules.scala 160:64:@31506.4]
  wire [13:0] _T_84414; // @[Modules.scala 160:64:@31507.4]
  wire [13:0] buffer_9_407; // @[Modules.scala 160:64:@31508.4]
  wire [13:0] buffer_9_188; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84416; // @[Modules.scala 160:64:@31510.4]
  wire [13:0] _T_84417; // @[Modules.scala 160:64:@31511.4]
  wire [13:0] buffer_9_408; // @[Modules.scala 160:64:@31512.4]
  wire [14:0] _T_84419; // @[Modules.scala 160:64:@31514.4]
  wire [13:0] _T_84420; // @[Modules.scala 160:64:@31515.4]
  wire [13:0] buffer_9_409; // @[Modules.scala 160:64:@31516.4]
  wire [13:0] buffer_9_192; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84422; // @[Modules.scala 160:64:@31518.4]
  wire [13:0] _T_84423; // @[Modules.scala 160:64:@31519.4]
  wire [13:0] buffer_9_410; // @[Modules.scala 160:64:@31520.4]
  wire [13:0] buffer_9_200; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84434; // @[Modules.scala 160:64:@31534.4]
  wire [13:0] _T_84435; // @[Modules.scala 160:64:@31535.4]
  wire [13:0] buffer_9_414; // @[Modules.scala 160:64:@31536.4]
  wire [13:0] buffer_9_202; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_203; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84437; // @[Modules.scala 160:64:@31538.4]
  wire [13:0] _T_84438; // @[Modules.scala 160:64:@31539.4]
  wire [13:0] buffer_9_415; // @[Modules.scala 160:64:@31540.4]
  wire [13:0] buffer_9_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84440; // @[Modules.scala 160:64:@31542.4]
  wire [13:0] _T_84441; // @[Modules.scala 160:64:@31543.4]
  wire [13:0] buffer_9_416; // @[Modules.scala 160:64:@31544.4]
  wire [13:0] buffer_9_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84443; // @[Modules.scala 160:64:@31546.4]
  wire [13:0] _T_84444; // @[Modules.scala 160:64:@31547.4]
  wire [13:0] buffer_9_417; // @[Modules.scala 160:64:@31548.4]
  wire [14:0] _T_84446; // @[Modules.scala 160:64:@31550.4]
  wire [13:0] _T_84447; // @[Modules.scala 160:64:@31551.4]
  wire [13:0] buffer_9_418; // @[Modules.scala 160:64:@31552.4]
  wire [14:0] _T_84452; // @[Modules.scala 160:64:@31558.4]
  wire [13:0] _T_84453; // @[Modules.scala 160:64:@31559.4]
  wire [13:0] buffer_9_420; // @[Modules.scala 160:64:@31560.4]
  wire [13:0] buffer_9_214; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84455; // @[Modules.scala 160:64:@31562.4]
  wire [13:0] _T_84456; // @[Modules.scala 160:64:@31563.4]
  wire [13:0] buffer_9_421; // @[Modules.scala 160:64:@31564.4]
  wire [14:0] _T_84458; // @[Modules.scala 160:64:@31566.4]
  wire [13:0] _T_84459; // @[Modules.scala 160:64:@31567.4]
  wire [13:0] buffer_9_422; // @[Modules.scala 160:64:@31568.4]
  wire [13:0] buffer_9_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84461; // @[Modules.scala 160:64:@31570.4]
  wire [13:0] _T_84462; // @[Modules.scala 160:64:@31571.4]
  wire [13:0] buffer_9_423; // @[Modules.scala 160:64:@31572.4]
  wire [13:0] buffer_9_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84467; // @[Modules.scala 160:64:@31578.4]
  wire [13:0] _T_84468; // @[Modules.scala 160:64:@31579.4]
  wire [13:0] buffer_9_425; // @[Modules.scala 160:64:@31580.4]
  wire [13:0] buffer_9_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84470; // @[Modules.scala 160:64:@31582.4]
  wire [13:0] _T_84471; // @[Modules.scala 160:64:@31583.4]
  wire [13:0] buffer_9_426; // @[Modules.scala 160:64:@31584.4]
  wire [14:0] _T_84473; // @[Modules.scala 160:64:@31586.4]
  wire [13:0] _T_84474; // @[Modules.scala 160:64:@31587.4]
  wire [13:0] buffer_9_427; // @[Modules.scala 160:64:@31588.4]
  wire [13:0] buffer_9_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84476; // @[Modules.scala 160:64:@31590.4]
  wire [13:0] _T_84477; // @[Modules.scala 160:64:@31591.4]
  wire [13:0] buffer_9_428; // @[Modules.scala 160:64:@31592.4]
  wire [13:0] buffer_9_230; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84479; // @[Modules.scala 160:64:@31594.4]
  wire [13:0] _T_84480; // @[Modules.scala 160:64:@31595.4]
  wire [13:0] buffer_9_429; // @[Modules.scala 160:64:@31596.4]
  wire [14:0] _T_84482; // @[Modules.scala 160:64:@31598.4]
  wire [13:0] _T_84483; // @[Modules.scala 160:64:@31599.4]
  wire [13:0] buffer_9_430; // @[Modules.scala 160:64:@31600.4]
  wire [13:0] buffer_9_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84485; // @[Modules.scala 160:64:@31602.4]
  wire [13:0] _T_84486; // @[Modules.scala 160:64:@31603.4]
  wire [13:0] buffer_9_431; // @[Modules.scala 160:64:@31604.4]
  wire [13:0] buffer_9_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84488; // @[Modules.scala 160:64:@31606.4]
  wire [13:0] _T_84489; // @[Modules.scala 160:64:@31607.4]
  wire [13:0] buffer_9_432; // @[Modules.scala 160:64:@31608.4]
  wire [13:0] buffer_9_238; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84491; // @[Modules.scala 160:64:@31610.4]
  wire [13:0] _T_84492; // @[Modules.scala 160:64:@31611.4]
  wire [13:0] buffer_9_433; // @[Modules.scala 160:64:@31612.4]
  wire [13:0] buffer_9_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84494; // @[Modules.scala 160:64:@31614.4]
  wire [13:0] _T_84495; // @[Modules.scala 160:64:@31615.4]
  wire [13:0] buffer_9_434; // @[Modules.scala 160:64:@31616.4]
  wire [13:0] buffer_9_242; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84497; // @[Modules.scala 160:64:@31618.4]
  wire [13:0] _T_84498; // @[Modules.scala 160:64:@31619.4]
  wire [13:0] buffer_9_435; // @[Modules.scala 160:64:@31620.4]
  wire [13:0] buffer_9_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84500; // @[Modules.scala 160:64:@31622.4]
  wire [13:0] _T_84501; // @[Modules.scala 160:64:@31623.4]
  wire [13:0] buffer_9_436; // @[Modules.scala 160:64:@31624.4]
  wire [13:0] buffer_9_246; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_247; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84503; // @[Modules.scala 160:64:@31626.4]
  wire [13:0] _T_84504; // @[Modules.scala 160:64:@31627.4]
  wire [13:0] buffer_9_437; // @[Modules.scala 160:64:@31628.4]
  wire [13:0] buffer_9_248; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84506; // @[Modules.scala 160:64:@31630.4]
  wire [13:0] _T_84507; // @[Modules.scala 160:64:@31631.4]
  wire [13:0] buffer_9_438; // @[Modules.scala 160:64:@31632.4]
  wire [13:0] buffer_9_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84509; // @[Modules.scala 160:64:@31634.4]
  wire [13:0] _T_84510; // @[Modules.scala 160:64:@31635.4]
  wire [13:0] buffer_9_439; // @[Modules.scala 160:64:@31636.4]
  wire [14:0] _T_84512; // @[Modules.scala 160:64:@31638.4]
  wire [13:0] _T_84513; // @[Modules.scala 160:64:@31639.4]
  wire [13:0] buffer_9_440; // @[Modules.scala 160:64:@31640.4]
  wire [14:0] _T_84518; // @[Modules.scala 160:64:@31646.4]
  wire [13:0] _T_84519; // @[Modules.scala 160:64:@31647.4]
  wire [13:0] buffer_9_442; // @[Modules.scala 160:64:@31648.4]
  wire [13:0] buffer_9_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84521; // @[Modules.scala 160:64:@31650.4]
  wire [13:0] _T_84522; // @[Modules.scala 160:64:@31651.4]
  wire [13:0] buffer_9_443; // @[Modules.scala 160:64:@31652.4]
  wire [13:0] buffer_9_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84524; // @[Modules.scala 160:64:@31654.4]
  wire [13:0] _T_84525; // @[Modules.scala 160:64:@31655.4]
  wire [13:0] buffer_9_444; // @[Modules.scala 160:64:@31656.4]
  wire [13:0] buffer_9_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84527; // @[Modules.scala 160:64:@31658.4]
  wire [13:0] _T_84528; // @[Modules.scala 160:64:@31659.4]
  wire [13:0] buffer_9_445; // @[Modules.scala 160:64:@31660.4]
  wire [14:0] _T_84530; // @[Modules.scala 160:64:@31662.4]
  wire [13:0] _T_84531; // @[Modules.scala 160:64:@31663.4]
  wire [13:0] buffer_9_446; // @[Modules.scala 160:64:@31664.4]
  wire [13:0] buffer_9_267; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84533; // @[Modules.scala 160:64:@31666.4]
  wire [13:0] _T_84534; // @[Modules.scala 160:64:@31667.4]
  wire [13:0] buffer_9_447; // @[Modules.scala 160:64:@31668.4]
  wire [13:0] buffer_9_268; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84536; // @[Modules.scala 160:64:@31670.4]
  wire [13:0] _T_84537; // @[Modules.scala 160:64:@31671.4]
  wire [13:0] buffer_9_448; // @[Modules.scala 160:64:@31672.4]
  wire [13:0] buffer_9_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84539; // @[Modules.scala 160:64:@31674.4]
  wire [13:0] _T_84540; // @[Modules.scala 160:64:@31675.4]
  wire [13:0] buffer_9_449; // @[Modules.scala 160:64:@31676.4]
  wire [14:0] _T_84542; // @[Modules.scala 160:64:@31678.4]
  wire [13:0] _T_84543; // @[Modules.scala 160:64:@31679.4]
  wire [13:0] buffer_9_450; // @[Modules.scala 160:64:@31680.4]
  wire [13:0] buffer_9_274; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_275; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84545; // @[Modules.scala 160:64:@31682.4]
  wire [13:0] _T_84546; // @[Modules.scala 160:64:@31683.4]
  wire [13:0] buffer_9_451; // @[Modules.scala 160:64:@31684.4]
  wire [13:0] buffer_9_276; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84548; // @[Modules.scala 160:64:@31686.4]
  wire [13:0] _T_84549; // @[Modules.scala 160:64:@31687.4]
  wire [13:0] buffer_9_452; // @[Modules.scala 160:64:@31688.4]
  wire [13:0] buffer_9_278; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84551; // @[Modules.scala 160:64:@31690.4]
  wire [13:0] _T_84552; // @[Modules.scala 160:64:@31691.4]
  wire [13:0] buffer_9_453; // @[Modules.scala 160:64:@31692.4]
  wire [13:0] buffer_9_280; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84554; // @[Modules.scala 160:64:@31694.4]
  wire [13:0] _T_84555; // @[Modules.scala 160:64:@31695.4]
  wire [13:0] buffer_9_454; // @[Modules.scala 160:64:@31696.4]
  wire [14:0] _T_84569; // @[Modules.scala 160:64:@31714.4]
  wire [13:0] _T_84570; // @[Modules.scala 160:64:@31715.4]
  wire [13:0] buffer_9_459; // @[Modules.scala 160:64:@31716.4]
  wire [13:0] buffer_9_292; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84572; // @[Modules.scala 160:64:@31718.4]
  wire [13:0] _T_84573; // @[Modules.scala 160:64:@31719.4]
  wire [13:0] buffer_9_460; // @[Modules.scala 160:64:@31720.4]
  wire [13:0] buffer_9_296; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_297; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84578; // @[Modules.scala 160:64:@31726.4]
  wire [13:0] _T_84579; // @[Modules.scala 160:64:@31727.4]
  wire [13:0] buffer_9_462; // @[Modules.scala 160:64:@31728.4]
  wire [13:0] buffer_9_298; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84581; // @[Modules.scala 160:64:@31730.4]
  wire [13:0] _T_84582; // @[Modules.scala 160:64:@31731.4]
  wire [13:0] buffer_9_463; // @[Modules.scala 160:64:@31732.4]
  wire [13:0] buffer_9_300; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_301; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84584; // @[Modules.scala 160:64:@31734.4]
  wire [13:0] _T_84585; // @[Modules.scala 160:64:@31735.4]
  wire [13:0] buffer_9_464; // @[Modules.scala 160:64:@31736.4]
  wire [14:0] _T_84587; // @[Modules.scala 160:64:@31738.4]
  wire [13:0] _T_84588; // @[Modules.scala 160:64:@31739.4]
  wire [13:0] buffer_9_465; // @[Modules.scala 160:64:@31740.4]
  wire [13:0] buffer_9_305; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84590; // @[Modules.scala 160:64:@31742.4]
  wire [13:0] _T_84591; // @[Modules.scala 160:64:@31743.4]
  wire [13:0] buffer_9_466; // @[Modules.scala 160:64:@31744.4]
  wire [13:0] buffer_9_307; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84593; // @[Modules.scala 160:64:@31746.4]
  wire [13:0] _T_84594; // @[Modules.scala 160:64:@31747.4]
  wire [13:0] buffer_9_467; // @[Modules.scala 160:64:@31748.4]
  wire [13:0] buffer_9_309; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84596; // @[Modules.scala 160:64:@31750.4]
  wire [13:0] _T_84597; // @[Modules.scala 160:64:@31751.4]
  wire [13:0] buffer_9_468; // @[Modules.scala 160:64:@31752.4]
  wire [13:0] buffer_9_310; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_311; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84599; // @[Modules.scala 160:64:@31754.4]
  wire [13:0] _T_84600; // @[Modules.scala 160:64:@31755.4]
  wire [13:0] buffer_9_469; // @[Modules.scala 160:64:@31756.4]
  wire [13:0] buffer_9_312; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_9_313; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_84602; // @[Modules.scala 160:64:@31758.4]
  wire [13:0] _T_84603; // @[Modules.scala 160:64:@31759.4]
  wire [13:0] buffer_9_470; // @[Modules.scala 160:64:@31760.4]
  wire [14:0] _T_84605; // @[Modules.scala 166:64:@31762.4]
  wire [13:0] _T_84606; // @[Modules.scala 166:64:@31763.4]
  wire [13:0] buffer_9_471; // @[Modules.scala 166:64:@31764.4]
  wire [14:0] _T_84608; // @[Modules.scala 166:64:@31766.4]
  wire [13:0] _T_84609; // @[Modules.scala 166:64:@31767.4]
  wire [13:0] buffer_9_472; // @[Modules.scala 166:64:@31768.4]
  wire [14:0] _T_84611; // @[Modules.scala 166:64:@31770.4]
  wire [13:0] _T_84612; // @[Modules.scala 166:64:@31771.4]
  wire [13:0] buffer_9_473; // @[Modules.scala 166:64:@31772.4]
  wire [14:0] _T_84614; // @[Modules.scala 166:64:@31774.4]
  wire [13:0] _T_84615; // @[Modules.scala 166:64:@31775.4]
  wire [13:0] buffer_9_474; // @[Modules.scala 166:64:@31776.4]
  wire [14:0] _T_84617; // @[Modules.scala 166:64:@31778.4]
  wire [13:0] _T_84618; // @[Modules.scala 166:64:@31779.4]
  wire [13:0] buffer_9_475; // @[Modules.scala 166:64:@31780.4]
  wire [14:0] _T_84620; // @[Modules.scala 166:64:@31782.4]
  wire [13:0] _T_84621; // @[Modules.scala 166:64:@31783.4]
  wire [13:0] buffer_9_476; // @[Modules.scala 166:64:@31784.4]
  wire [14:0] _T_84623; // @[Modules.scala 166:64:@31786.4]
  wire [13:0] _T_84624; // @[Modules.scala 166:64:@31787.4]
  wire [13:0] buffer_9_477; // @[Modules.scala 166:64:@31788.4]
  wire [14:0] _T_84626; // @[Modules.scala 166:64:@31790.4]
  wire [13:0] _T_84627; // @[Modules.scala 166:64:@31791.4]
  wire [13:0] buffer_9_478; // @[Modules.scala 166:64:@31792.4]
  wire [14:0] _T_84629; // @[Modules.scala 166:64:@31794.4]
  wire [13:0] _T_84630; // @[Modules.scala 166:64:@31795.4]
  wire [13:0] buffer_9_479; // @[Modules.scala 166:64:@31796.4]
  wire [14:0] _T_84632; // @[Modules.scala 166:64:@31798.4]
  wire [13:0] _T_84633; // @[Modules.scala 166:64:@31799.4]
  wire [13:0] buffer_9_480; // @[Modules.scala 166:64:@31800.4]
  wire [14:0] _T_84635; // @[Modules.scala 166:64:@31802.4]
  wire [13:0] _T_84636; // @[Modules.scala 166:64:@31803.4]
  wire [13:0] buffer_9_481; // @[Modules.scala 166:64:@31804.4]
  wire [14:0] _T_84638; // @[Modules.scala 166:64:@31806.4]
  wire [13:0] _T_84639; // @[Modules.scala 166:64:@31807.4]
  wire [13:0] buffer_9_482; // @[Modules.scala 166:64:@31808.4]
  wire [14:0] _T_84641; // @[Modules.scala 166:64:@31810.4]
  wire [13:0] _T_84642; // @[Modules.scala 166:64:@31811.4]
  wire [13:0] buffer_9_483; // @[Modules.scala 166:64:@31812.4]
  wire [14:0] _T_84644; // @[Modules.scala 166:64:@31814.4]
  wire [13:0] _T_84645; // @[Modules.scala 166:64:@31815.4]
  wire [13:0] buffer_9_484; // @[Modules.scala 166:64:@31816.4]
  wire [14:0] _T_84647; // @[Modules.scala 166:64:@31818.4]
  wire [13:0] _T_84648; // @[Modules.scala 166:64:@31819.4]
  wire [13:0] buffer_9_485; // @[Modules.scala 166:64:@31820.4]
  wire [14:0] _T_84650; // @[Modules.scala 166:64:@31822.4]
  wire [13:0] _T_84651; // @[Modules.scala 166:64:@31823.4]
  wire [13:0] buffer_9_486; // @[Modules.scala 166:64:@31824.4]
  wire [14:0] _T_84656; // @[Modules.scala 166:64:@31830.4]
  wire [13:0] _T_84657; // @[Modules.scala 166:64:@31831.4]
  wire [13:0] buffer_9_488; // @[Modules.scala 166:64:@31832.4]
  wire [14:0] _T_84659; // @[Modules.scala 166:64:@31834.4]
  wire [13:0] _T_84660; // @[Modules.scala 166:64:@31835.4]
  wire [13:0] buffer_9_489; // @[Modules.scala 166:64:@31836.4]
  wire [14:0] _T_84662; // @[Modules.scala 166:64:@31838.4]
  wire [13:0] _T_84663; // @[Modules.scala 166:64:@31839.4]
  wire [13:0] buffer_9_490; // @[Modules.scala 166:64:@31840.4]
  wire [14:0] _T_84665; // @[Modules.scala 166:64:@31842.4]
  wire [13:0] _T_84666; // @[Modules.scala 166:64:@31843.4]
  wire [13:0] buffer_9_491; // @[Modules.scala 166:64:@31844.4]
  wire [14:0] _T_84668; // @[Modules.scala 166:64:@31846.4]
  wire [13:0] _T_84669; // @[Modules.scala 166:64:@31847.4]
  wire [13:0] buffer_9_492; // @[Modules.scala 166:64:@31848.4]
  wire [14:0] _T_84671; // @[Modules.scala 166:64:@31850.4]
  wire [13:0] _T_84672; // @[Modules.scala 166:64:@31851.4]
  wire [13:0] buffer_9_493; // @[Modules.scala 166:64:@31852.4]
  wire [14:0] _T_84674; // @[Modules.scala 166:64:@31854.4]
  wire [13:0] _T_84675; // @[Modules.scala 166:64:@31855.4]
  wire [13:0] buffer_9_494; // @[Modules.scala 166:64:@31856.4]
  wire [14:0] _T_84677; // @[Modules.scala 166:64:@31858.4]
  wire [13:0] _T_84678; // @[Modules.scala 166:64:@31859.4]
  wire [13:0] buffer_9_495; // @[Modules.scala 166:64:@31860.4]
  wire [14:0] _T_84680; // @[Modules.scala 166:64:@31862.4]
  wire [13:0] _T_84681; // @[Modules.scala 166:64:@31863.4]
  wire [13:0] buffer_9_496; // @[Modules.scala 166:64:@31864.4]
  wire [14:0] _T_84683; // @[Modules.scala 166:64:@31866.4]
  wire [13:0] _T_84684; // @[Modules.scala 166:64:@31867.4]
  wire [13:0] buffer_9_497; // @[Modules.scala 166:64:@31868.4]
  wire [14:0] _T_84686; // @[Modules.scala 166:64:@31870.4]
  wire [13:0] _T_84687; // @[Modules.scala 166:64:@31871.4]
  wire [13:0] buffer_9_498; // @[Modules.scala 166:64:@31872.4]
  wire [14:0] _T_84689; // @[Modules.scala 166:64:@31874.4]
  wire [13:0] _T_84690; // @[Modules.scala 166:64:@31875.4]
  wire [13:0] buffer_9_499; // @[Modules.scala 166:64:@31876.4]
  wire [14:0] _T_84692; // @[Modules.scala 166:64:@31878.4]
  wire [13:0] _T_84693; // @[Modules.scala 166:64:@31879.4]
  wire [13:0] buffer_9_500; // @[Modules.scala 166:64:@31880.4]
  wire [14:0] _T_84695; // @[Modules.scala 166:64:@31882.4]
  wire [13:0] _T_84696; // @[Modules.scala 166:64:@31883.4]
  wire [13:0] buffer_9_501; // @[Modules.scala 166:64:@31884.4]
  wire [14:0] _T_84698; // @[Modules.scala 166:64:@31886.4]
  wire [13:0] _T_84699; // @[Modules.scala 166:64:@31887.4]
  wire [13:0] buffer_9_502; // @[Modules.scala 166:64:@31888.4]
  wire [14:0] _T_84701; // @[Modules.scala 166:64:@31890.4]
  wire [13:0] _T_84702; // @[Modules.scala 166:64:@31891.4]
  wire [13:0] buffer_9_503; // @[Modules.scala 166:64:@31892.4]
  wire [14:0] _T_84704; // @[Modules.scala 166:64:@31894.4]
  wire [13:0] _T_84705; // @[Modules.scala 166:64:@31895.4]
  wire [13:0] buffer_9_504; // @[Modules.scala 166:64:@31896.4]
  wire [14:0] _T_84710; // @[Modules.scala 166:64:@31902.4]
  wire [13:0] _T_84711; // @[Modules.scala 166:64:@31903.4]
  wire [13:0] buffer_9_506; // @[Modules.scala 166:64:@31904.4]
  wire [14:0] _T_84713; // @[Modules.scala 166:64:@31906.4]
  wire [13:0] _T_84714; // @[Modules.scala 166:64:@31907.4]
  wire [13:0] buffer_9_507; // @[Modules.scala 166:64:@31908.4]
  wire [14:0] _T_84716; // @[Modules.scala 166:64:@31910.4]
  wire [13:0] _T_84717; // @[Modules.scala 166:64:@31911.4]
  wire [13:0] buffer_9_508; // @[Modules.scala 166:64:@31912.4]
  wire [14:0] _T_84719; // @[Modules.scala 166:64:@31914.4]
  wire [13:0] _T_84720; // @[Modules.scala 166:64:@31915.4]
  wire [13:0] buffer_9_509; // @[Modules.scala 166:64:@31916.4]
  wire [14:0] _T_84722; // @[Modules.scala 166:64:@31918.4]
  wire [13:0] _T_84723; // @[Modules.scala 166:64:@31919.4]
  wire [13:0] buffer_9_510; // @[Modules.scala 166:64:@31920.4]
  wire [14:0] _T_84728; // @[Modules.scala 166:64:@31926.4]
  wire [13:0] _T_84729; // @[Modules.scala 166:64:@31927.4]
  wire [13:0] buffer_9_512; // @[Modules.scala 166:64:@31928.4]
  wire [14:0] _T_84731; // @[Modules.scala 166:64:@31930.4]
  wire [13:0] _T_84732; // @[Modules.scala 166:64:@31931.4]
  wire [13:0] buffer_9_513; // @[Modules.scala 166:64:@31932.4]
  wire [14:0] _T_84734; // @[Modules.scala 166:64:@31934.4]
  wire [13:0] _T_84735; // @[Modules.scala 166:64:@31935.4]
  wire [13:0] buffer_9_514; // @[Modules.scala 166:64:@31936.4]
  wire [14:0] _T_84737; // @[Modules.scala 166:64:@31938.4]
  wire [13:0] _T_84738; // @[Modules.scala 166:64:@31939.4]
  wire [13:0] buffer_9_515; // @[Modules.scala 166:64:@31940.4]
  wire [14:0] _T_84740; // @[Modules.scala 166:64:@31942.4]
  wire [13:0] _T_84741; // @[Modules.scala 166:64:@31943.4]
  wire [13:0] buffer_9_516; // @[Modules.scala 166:64:@31944.4]
  wire [14:0] _T_84743; // @[Modules.scala 166:64:@31946.4]
  wire [13:0] _T_84744; // @[Modules.scala 166:64:@31947.4]
  wire [13:0] buffer_9_517; // @[Modules.scala 166:64:@31948.4]
  wire [14:0] _T_84746; // @[Modules.scala 166:64:@31950.4]
  wire [13:0] _T_84747; // @[Modules.scala 166:64:@31951.4]
  wire [13:0] buffer_9_518; // @[Modules.scala 166:64:@31952.4]
  wire [14:0] _T_84749; // @[Modules.scala 166:64:@31954.4]
  wire [13:0] _T_84750; // @[Modules.scala 166:64:@31955.4]
  wire [13:0] buffer_9_519; // @[Modules.scala 166:64:@31956.4]
  wire [14:0] _T_84755; // @[Modules.scala 166:64:@31962.4]
  wire [13:0] _T_84756; // @[Modules.scala 166:64:@31963.4]
  wire [13:0] buffer_9_521; // @[Modules.scala 166:64:@31964.4]
  wire [14:0] _T_84758; // @[Modules.scala 166:64:@31966.4]
  wire [13:0] _T_84759; // @[Modules.scala 166:64:@31967.4]
  wire [13:0] buffer_9_522; // @[Modules.scala 166:64:@31968.4]
  wire [14:0] _T_84761; // @[Modules.scala 166:64:@31970.4]
  wire [13:0] _T_84762; // @[Modules.scala 166:64:@31971.4]
  wire [13:0] buffer_9_523; // @[Modules.scala 166:64:@31972.4]
  wire [14:0] _T_84764; // @[Modules.scala 166:64:@31974.4]
  wire [13:0] _T_84765; // @[Modules.scala 166:64:@31975.4]
  wire [13:0] buffer_9_524; // @[Modules.scala 166:64:@31976.4]
  wire [14:0] _T_84767; // @[Modules.scala 166:64:@31978.4]
  wire [13:0] _T_84768; // @[Modules.scala 166:64:@31979.4]
  wire [13:0] buffer_9_525; // @[Modules.scala 166:64:@31980.4]
  wire [14:0] _T_84770; // @[Modules.scala 166:64:@31982.4]
  wire [13:0] _T_84771; // @[Modules.scala 166:64:@31983.4]
  wire [13:0] buffer_9_526; // @[Modules.scala 166:64:@31984.4]
  wire [14:0] _T_84773; // @[Modules.scala 166:64:@31986.4]
  wire [13:0] _T_84774; // @[Modules.scala 166:64:@31987.4]
  wire [13:0] buffer_9_527; // @[Modules.scala 166:64:@31988.4]
  wire [14:0] _T_84776; // @[Modules.scala 166:64:@31990.4]
  wire [13:0] _T_84777; // @[Modules.scala 166:64:@31991.4]
  wire [13:0] buffer_9_528; // @[Modules.scala 166:64:@31992.4]
  wire [14:0] _T_84779; // @[Modules.scala 166:64:@31994.4]
  wire [13:0] _T_84780; // @[Modules.scala 166:64:@31995.4]
  wire [13:0] buffer_9_529; // @[Modules.scala 166:64:@31996.4]
  wire [14:0] _T_84782; // @[Modules.scala 166:64:@31998.4]
  wire [13:0] _T_84783; // @[Modules.scala 166:64:@31999.4]
  wire [13:0] buffer_9_530; // @[Modules.scala 166:64:@32000.4]
  wire [14:0] _T_84785; // @[Modules.scala 166:64:@32002.4]
  wire [13:0] _T_84786; // @[Modules.scala 166:64:@32003.4]
  wire [13:0] buffer_9_531; // @[Modules.scala 166:64:@32004.4]
  wire [14:0] _T_84788; // @[Modules.scala 166:64:@32006.4]
  wire [13:0] _T_84789; // @[Modules.scala 166:64:@32007.4]
  wire [13:0] buffer_9_532; // @[Modules.scala 166:64:@32008.4]
  wire [14:0] _T_84791; // @[Modules.scala 166:64:@32010.4]
  wire [13:0] _T_84792; // @[Modules.scala 166:64:@32011.4]
  wire [13:0] buffer_9_533; // @[Modules.scala 166:64:@32012.4]
  wire [14:0] _T_84794; // @[Modules.scala 166:64:@32014.4]
  wire [13:0] _T_84795; // @[Modules.scala 166:64:@32015.4]
  wire [13:0] buffer_9_534; // @[Modules.scala 166:64:@32016.4]
  wire [14:0] _T_84797; // @[Modules.scala 166:64:@32018.4]
  wire [13:0] _T_84798; // @[Modules.scala 166:64:@32019.4]
  wire [13:0] buffer_9_535; // @[Modules.scala 166:64:@32020.4]
  wire [14:0] _T_84800; // @[Modules.scala 166:64:@32022.4]
  wire [13:0] _T_84801; // @[Modules.scala 166:64:@32023.4]
  wire [13:0] buffer_9_536; // @[Modules.scala 166:64:@32024.4]
  wire [14:0] _T_84803; // @[Modules.scala 166:64:@32026.4]
  wire [13:0] _T_84804; // @[Modules.scala 166:64:@32027.4]
  wire [13:0] buffer_9_537; // @[Modules.scala 166:64:@32028.4]
  wire [14:0] _T_84806; // @[Modules.scala 166:64:@32030.4]
  wire [13:0] _T_84807; // @[Modules.scala 166:64:@32031.4]
  wire [13:0] buffer_9_538; // @[Modules.scala 166:64:@32032.4]
  wire [14:0] _T_84809; // @[Modules.scala 166:64:@32034.4]
  wire [13:0] _T_84810; // @[Modules.scala 166:64:@32035.4]
  wire [13:0] buffer_9_539; // @[Modules.scala 166:64:@32036.4]
  wire [14:0] _T_84812; // @[Modules.scala 166:64:@32038.4]
  wire [13:0] _T_84813; // @[Modules.scala 166:64:@32039.4]
  wire [13:0] buffer_9_540; // @[Modules.scala 166:64:@32040.4]
  wire [14:0] _T_84815; // @[Modules.scala 166:64:@32042.4]
  wire [13:0] _T_84816; // @[Modules.scala 166:64:@32043.4]
  wire [13:0] buffer_9_541; // @[Modules.scala 166:64:@32044.4]
  wire [14:0] _T_84821; // @[Modules.scala 166:64:@32050.4]
  wire [13:0] _T_84822; // @[Modules.scala 166:64:@32051.4]
  wire [13:0] buffer_9_543; // @[Modules.scala 166:64:@32052.4]
  wire [14:0] _T_84824; // @[Modules.scala 166:64:@32054.4]
  wire [13:0] _T_84825; // @[Modules.scala 166:64:@32055.4]
  wire [13:0] buffer_9_544; // @[Modules.scala 166:64:@32056.4]
  wire [14:0] _T_84827; // @[Modules.scala 166:64:@32058.4]
  wire [13:0] _T_84828; // @[Modules.scala 166:64:@32059.4]
  wire [13:0] buffer_9_545; // @[Modules.scala 166:64:@32060.4]
  wire [14:0] _T_84830; // @[Modules.scala 166:64:@32062.4]
  wire [13:0] _T_84831; // @[Modules.scala 166:64:@32063.4]
  wire [13:0] buffer_9_546; // @[Modules.scala 166:64:@32064.4]
  wire [14:0] _T_84833; // @[Modules.scala 166:64:@32066.4]
  wire [13:0] _T_84834; // @[Modules.scala 166:64:@32067.4]
  wire [13:0] buffer_9_547; // @[Modules.scala 166:64:@32068.4]
  wire [14:0] _T_84836; // @[Modules.scala 166:64:@32070.4]
  wire [13:0] _T_84837; // @[Modules.scala 166:64:@32071.4]
  wire [13:0] buffer_9_548; // @[Modules.scala 166:64:@32072.4]
  wire [14:0] _T_84839; // @[Modules.scala 160:64:@32074.4]
  wire [13:0] _T_84840; // @[Modules.scala 160:64:@32075.4]
  wire [13:0] buffer_9_549; // @[Modules.scala 160:64:@32076.4]
  wire [14:0] _T_84842; // @[Modules.scala 160:64:@32078.4]
  wire [13:0] _T_84843; // @[Modules.scala 160:64:@32079.4]
  wire [13:0] buffer_9_550; // @[Modules.scala 160:64:@32080.4]
  wire [14:0] _T_84845; // @[Modules.scala 160:64:@32082.4]
  wire [13:0] _T_84846; // @[Modules.scala 160:64:@32083.4]
  wire [13:0] buffer_9_551; // @[Modules.scala 160:64:@32084.4]
  wire [14:0] _T_84848; // @[Modules.scala 160:64:@32086.4]
  wire [13:0] _T_84849; // @[Modules.scala 160:64:@32087.4]
  wire [13:0] buffer_9_552; // @[Modules.scala 160:64:@32088.4]
  wire [14:0] _T_84851; // @[Modules.scala 160:64:@32090.4]
  wire [13:0] _T_84852; // @[Modules.scala 160:64:@32091.4]
  wire [13:0] buffer_9_553; // @[Modules.scala 160:64:@32092.4]
  wire [14:0] _T_84854; // @[Modules.scala 160:64:@32094.4]
  wire [13:0] _T_84855; // @[Modules.scala 160:64:@32095.4]
  wire [13:0] buffer_9_554; // @[Modules.scala 160:64:@32096.4]
  wire [14:0] _T_84857; // @[Modules.scala 160:64:@32098.4]
  wire [13:0] _T_84858; // @[Modules.scala 160:64:@32099.4]
  wire [13:0] buffer_9_555; // @[Modules.scala 160:64:@32100.4]
  wire [14:0] _T_84860; // @[Modules.scala 160:64:@32102.4]
  wire [13:0] _T_84861; // @[Modules.scala 160:64:@32103.4]
  wire [13:0] buffer_9_556; // @[Modules.scala 160:64:@32104.4]
  wire [14:0] _T_84863; // @[Modules.scala 160:64:@32106.4]
  wire [13:0] _T_84864; // @[Modules.scala 160:64:@32107.4]
  wire [13:0] buffer_9_557; // @[Modules.scala 160:64:@32108.4]
  wire [14:0] _T_84866; // @[Modules.scala 160:64:@32110.4]
  wire [13:0] _T_84867; // @[Modules.scala 160:64:@32111.4]
  wire [13:0] buffer_9_558; // @[Modules.scala 160:64:@32112.4]
  wire [14:0] _T_84869; // @[Modules.scala 160:64:@32114.4]
  wire [13:0] _T_84870; // @[Modules.scala 160:64:@32115.4]
  wire [13:0] buffer_9_559; // @[Modules.scala 160:64:@32116.4]
  wire [14:0] _T_84872; // @[Modules.scala 160:64:@32118.4]
  wire [13:0] _T_84873; // @[Modules.scala 160:64:@32119.4]
  wire [13:0] buffer_9_560; // @[Modules.scala 160:64:@32120.4]
  wire [14:0] _T_84875; // @[Modules.scala 160:64:@32122.4]
  wire [13:0] _T_84876; // @[Modules.scala 160:64:@32123.4]
  wire [13:0] buffer_9_561; // @[Modules.scala 160:64:@32124.4]
  wire [14:0] _T_84878; // @[Modules.scala 160:64:@32126.4]
  wire [13:0] _T_84879; // @[Modules.scala 160:64:@32127.4]
  wire [13:0] buffer_9_562; // @[Modules.scala 160:64:@32128.4]
  wire [14:0] _T_84881; // @[Modules.scala 160:64:@32130.4]
  wire [13:0] _T_84882; // @[Modules.scala 160:64:@32131.4]
  wire [13:0] buffer_9_563; // @[Modules.scala 160:64:@32132.4]
  wire [14:0] _T_84884; // @[Modules.scala 160:64:@32134.4]
  wire [13:0] _T_84885; // @[Modules.scala 160:64:@32135.4]
  wire [13:0] buffer_9_564; // @[Modules.scala 160:64:@32136.4]
  wire [14:0] _T_84887; // @[Modules.scala 160:64:@32138.4]
  wire [13:0] _T_84888; // @[Modules.scala 160:64:@32139.4]
  wire [13:0] buffer_9_565; // @[Modules.scala 160:64:@32140.4]
  wire [14:0] _T_84890; // @[Modules.scala 160:64:@32142.4]
  wire [13:0] _T_84891; // @[Modules.scala 160:64:@32143.4]
  wire [13:0] buffer_9_566; // @[Modules.scala 160:64:@32144.4]
  wire [14:0] _T_84893; // @[Modules.scala 160:64:@32146.4]
  wire [13:0] _T_84894; // @[Modules.scala 160:64:@32147.4]
  wire [13:0] buffer_9_567; // @[Modules.scala 160:64:@32148.4]
  wire [14:0] _T_84896; // @[Modules.scala 160:64:@32150.4]
  wire [13:0] _T_84897; // @[Modules.scala 160:64:@32151.4]
  wire [13:0] buffer_9_568; // @[Modules.scala 160:64:@32152.4]
  wire [14:0] _T_84899; // @[Modules.scala 160:64:@32154.4]
  wire [13:0] _T_84900; // @[Modules.scala 160:64:@32155.4]
  wire [13:0] buffer_9_569; // @[Modules.scala 160:64:@32156.4]
  wire [14:0] _T_84902; // @[Modules.scala 160:64:@32158.4]
  wire [13:0] _T_84903; // @[Modules.scala 160:64:@32159.4]
  wire [13:0] buffer_9_570; // @[Modules.scala 160:64:@32160.4]
  wire [14:0] _T_84905; // @[Modules.scala 160:64:@32162.4]
  wire [13:0] _T_84906; // @[Modules.scala 160:64:@32163.4]
  wire [13:0] buffer_9_571; // @[Modules.scala 160:64:@32164.4]
  wire [14:0] _T_84908; // @[Modules.scala 160:64:@32166.4]
  wire [13:0] _T_84909; // @[Modules.scala 160:64:@32167.4]
  wire [13:0] buffer_9_572; // @[Modules.scala 160:64:@32168.4]
  wire [14:0] _T_84911; // @[Modules.scala 160:64:@32170.4]
  wire [13:0] _T_84912; // @[Modules.scala 160:64:@32171.4]
  wire [13:0] buffer_9_573; // @[Modules.scala 160:64:@32172.4]
  wire [14:0] _T_84914; // @[Modules.scala 160:64:@32174.4]
  wire [13:0] _T_84915; // @[Modules.scala 160:64:@32175.4]
  wire [13:0] buffer_9_574; // @[Modules.scala 160:64:@32176.4]
  wire [14:0] _T_84917; // @[Modules.scala 160:64:@32178.4]
  wire [13:0] _T_84918; // @[Modules.scala 160:64:@32179.4]
  wire [13:0] buffer_9_575; // @[Modules.scala 160:64:@32180.4]
  wire [14:0] _T_84920; // @[Modules.scala 160:64:@32182.4]
  wire [13:0] _T_84921; // @[Modules.scala 160:64:@32183.4]
  wire [13:0] buffer_9_576; // @[Modules.scala 160:64:@32184.4]
  wire [14:0] _T_84923; // @[Modules.scala 160:64:@32186.4]
  wire [13:0] _T_84924; // @[Modules.scala 160:64:@32187.4]
  wire [13:0] buffer_9_577; // @[Modules.scala 160:64:@32188.4]
  wire [14:0] _T_84926; // @[Modules.scala 160:64:@32190.4]
  wire [13:0] _T_84927; // @[Modules.scala 160:64:@32191.4]
  wire [13:0] buffer_9_578; // @[Modules.scala 160:64:@32192.4]
  wire [14:0] _T_84929; // @[Modules.scala 160:64:@32194.4]
  wire [13:0] _T_84930; // @[Modules.scala 160:64:@32195.4]
  wire [13:0] buffer_9_579; // @[Modules.scala 160:64:@32196.4]
  wire [14:0] _T_84932; // @[Modules.scala 160:64:@32198.4]
  wire [13:0] _T_84933; // @[Modules.scala 160:64:@32199.4]
  wire [13:0] buffer_9_580; // @[Modules.scala 160:64:@32200.4]
  wire [14:0] _T_84935; // @[Modules.scala 160:64:@32202.4]
  wire [13:0] _T_84936; // @[Modules.scala 160:64:@32203.4]
  wire [13:0] buffer_9_581; // @[Modules.scala 160:64:@32204.4]
  wire [14:0] _T_84938; // @[Modules.scala 160:64:@32206.4]
  wire [13:0] _T_84939; // @[Modules.scala 160:64:@32207.4]
  wire [13:0] buffer_9_582; // @[Modules.scala 160:64:@32208.4]
  wire [14:0] _T_84941; // @[Modules.scala 160:64:@32210.4]
  wire [13:0] _T_84942; // @[Modules.scala 160:64:@32211.4]
  wire [13:0] buffer_9_583; // @[Modules.scala 160:64:@32212.4]
  wire [14:0] _T_84944; // @[Modules.scala 160:64:@32214.4]
  wire [13:0] _T_84945; // @[Modules.scala 160:64:@32215.4]
  wire [13:0] buffer_9_584; // @[Modules.scala 160:64:@32216.4]
  wire [14:0] _T_84947; // @[Modules.scala 160:64:@32218.4]
  wire [13:0] _T_84948; // @[Modules.scala 160:64:@32219.4]
  wire [13:0] buffer_9_585; // @[Modules.scala 160:64:@32220.4]
  wire [14:0] _T_84950; // @[Modules.scala 160:64:@32222.4]
  wire [13:0] _T_84951; // @[Modules.scala 160:64:@32223.4]
  wire [13:0] buffer_9_586; // @[Modules.scala 160:64:@32224.4]
  wire [14:0] _T_84953; // @[Modules.scala 160:64:@32226.4]
  wire [13:0] _T_84954; // @[Modules.scala 160:64:@32227.4]
  wire [13:0] buffer_9_587; // @[Modules.scala 160:64:@32228.4]
  wire [14:0] _T_84956; // @[Modules.scala 166:64:@32230.4]
  wire [13:0] _T_84957; // @[Modules.scala 166:64:@32231.4]
  wire [13:0] buffer_9_588; // @[Modules.scala 166:64:@32232.4]
  wire [14:0] _T_84959; // @[Modules.scala 166:64:@32234.4]
  wire [13:0] _T_84960; // @[Modules.scala 166:64:@32235.4]
  wire [13:0] buffer_9_589; // @[Modules.scala 166:64:@32236.4]
  wire [14:0] _T_84962; // @[Modules.scala 166:64:@32238.4]
  wire [13:0] _T_84963; // @[Modules.scala 166:64:@32239.4]
  wire [13:0] buffer_9_590; // @[Modules.scala 166:64:@32240.4]
  wire [14:0] _T_84965; // @[Modules.scala 166:64:@32242.4]
  wire [13:0] _T_84966; // @[Modules.scala 166:64:@32243.4]
  wire [13:0] buffer_9_591; // @[Modules.scala 166:64:@32244.4]
  wire [14:0] _T_84968; // @[Modules.scala 166:64:@32246.4]
  wire [13:0] _T_84969; // @[Modules.scala 166:64:@32247.4]
  wire [13:0] buffer_9_592; // @[Modules.scala 166:64:@32248.4]
  wire [14:0] _T_84971; // @[Modules.scala 166:64:@32250.4]
  wire [13:0] _T_84972; // @[Modules.scala 166:64:@32251.4]
  wire [13:0] buffer_9_593; // @[Modules.scala 166:64:@32252.4]
  wire [14:0] _T_84974; // @[Modules.scala 166:64:@32254.4]
  wire [13:0] _T_84975; // @[Modules.scala 166:64:@32255.4]
  wire [13:0] buffer_9_594; // @[Modules.scala 166:64:@32256.4]
  wire [14:0] _T_84977; // @[Modules.scala 166:64:@32258.4]
  wire [13:0] _T_84978; // @[Modules.scala 166:64:@32259.4]
  wire [13:0] buffer_9_595; // @[Modules.scala 166:64:@32260.4]
  wire [14:0] _T_84980; // @[Modules.scala 166:64:@32262.4]
  wire [13:0] _T_84981; // @[Modules.scala 166:64:@32263.4]
  wire [13:0] buffer_9_596; // @[Modules.scala 166:64:@32264.4]
  wire [14:0] _T_84983; // @[Modules.scala 166:64:@32266.4]
  wire [13:0] _T_84984; // @[Modules.scala 166:64:@32267.4]
  wire [13:0] buffer_9_597; // @[Modules.scala 166:64:@32268.4]
  wire [14:0] _T_84986; // @[Modules.scala 166:64:@32270.4]
  wire [13:0] _T_84987; // @[Modules.scala 166:64:@32271.4]
  wire [13:0] buffer_9_598; // @[Modules.scala 166:64:@32272.4]
  wire [14:0] _T_84989; // @[Modules.scala 166:64:@32274.4]
  wire [13:0] _T_84990; // @[Modules.scala 166:64:@32275.4]
  wire [13:0] buffer_9_599; // @[Modules.scala 166:64:@32276.4]
  wire [14:0] _T_84992; // @[Modules.scala 166:64:@32278.4]
  wire [13:0] _T_84993; // @[Modules.scala 166:64:@32279.4]
  wire [13:0] buffer_9_600; // @[Modules.scala 166:64:@32280.4]
  wire [14:0] _T_84995; // @[Modules.scala 166:64:@32282.4]
  wire [13:0] _T_84996; // @[Modules.scala 166:64:@32283.4]
  wire [13:0] buffer_9_601; // @[Modules.scala 166:64:@32284.4]
  wire [14:0] _T_84998; // @[Modules.scala 166:64:@32286.4]
  wire [13:0] _T_84999; // @[Modules.scala 166:64:@32287.4]
  wire [13:0] buffer_9_602; // @[Modules.scala 166:64:@32288.4]
  wire [14:0] _T_85001; // @[Modules.scala 166:64:@32290.4]
  wire [13:0] _T_85002; // @[Modules.scala 166:64:@32291.4]
  wire [13:0] buffer_9_603; // @[Modules.scala 166:64:@32292.4]
  wire [14:0] _T_85004; // @[Modules.scala 166:64:@32294.4]
  wire [13:0] _T_85005; // @[Modules.scala 166:64:@32295.4]
  wire [13:0] buffer_9_604; // @[Modules.scala 166:64:@32296.4]
  wire [14:0] _T_85007; // @[Modules.scala 166:64:@32298.4]
  wire [13:0] _T_85008; // @[Modules.scala 166:64:@32299.4]
  wire [13:0] buffer_9_605; // @[Modules.scala 166:64:@32300.4]
  wire [14:0] _T_85010; // @[Modules.scala 166:64:@32302.4]
  wire [13:0] _T_85011; // @[Modules.scala 166:64:@32303.4]
  wire [13:0] buffer_9_606; // @[Modules.scala 166:64:@32304.4]
  wire [14:0] _T_85013; // @[Modules.scala 172:66:@32306.4]
  wire [13:0] _T_85014; // @[Modules.scala 172:66:@32307.4]
  wire [13:0] buffer_9_607; // @[Modules.scala 172:66:@32308.4]
  wire [14:0] _T_85016; // @[Modules.scala 160:64:@32310.4]
  wire [13:0] _T_85017; // @[Modules.scala 160:64:@32311.4]
  wire [13:0] buffer_9_608; // @[Modules.scala 160:64:@32312.4]
  wire [14:0] _T_85019; // @[Modules.scala 160:64:@32314.4]
  wire [13:0] _T_85020; // @[Modules.scala 160:64:@32315.4]
  wire [13:0] buffer_9_609; // @[Modules.scala 160:64:@32316.4]
  wire [14:0] _T_85022; // @[Modules.scala 160:64:@32318.4]
  wire [13:0] _T_85023; // @[Modules.scala 160:64:@32319.4]
  wire [13:0] buffer_9_610; // @[Modules.scala 160:64:@32320.4]
  wire [14:0] _T_85025; // @[Modules.scala 160:64:@32322.4]
  wire [13:0] _T_85026; // @[Modules.scala 160:64:@32323.4]
  wire [13:0] buffer_9_611; // @[Modules.scala 160:64:@32324.4]
  wire [14:0] _T_85028; // @[Modules.scala 160:64:@32326.4]
  wire [13:0] _T_85029; // @[Modules.scala 160:64:@32327.4]
  wire [13:0] buffer_9_612; // @[Modules.scala 160:64:@32328.4]
  wire [14:0] _T_85031; // @[Modules.scala 160:64:@32330.4]
  wire [13:0] _T_85032; // @[Modules.scala 160:64:@32331.4]
  wire [13:0] buffer_9_613; // @[Modules.scala 160:64:@32332.4]
  wire [14:0] _T_85034; // @[Modules.scala 160:64:@32334.4]
  wire [13:0] _T_85035; // @[Modules.scala 160:64:@32335.4]
  wire [13:0] buffer_9_614; // @[Modules.scala 160:64:@32336.4]
  wire [14:0] _T_85037; // @[Modules.scala 160:64:@32338.4]
  wire [13:0] _T_85038; // @[Modules.scala 160:64:@32339.4]
  wire [13:0] buffer_9_615; // @[Modules.scala 160:64:@32340.4]
  wire [14:0] _T_85040; // @[Modules.scala 160:64:@32342.4]
  wire [13:0] _T_85041; // @[Modules.scala 160:64:@32343.4]
  wire [13:0] buffer_9_616; // @[Modules.scala 160:64:@32344.4]
  wire [14:0] _T_85043; // @[Modules.scala 160:64:@32346.4]
  wire [13:0] _T_85044; // @[Modules.scala 160:64:@32347.4]
  wire [13:0] buffer_9_617; // @[Modules.scala 160:64:@32348.4]
  wire [14:0] _T_85046; // @[Modules.scala 160:64:@32350.4]
  wire [13:0] _T_85047; // @[Modules.scala 160:64:@32351.4]
  wire [13:0] buffer_9_618; // @[Modules.scala 160:64:@32352.4]
  wire [14:0] _T_85049; // @[Modules.scala 160:64:@32354.4]
  wire [13:0] _T_85050; // @[Modules.scala 160:64:@32355.4]
  wire [13:0] buffer_9_619; // @[Modules.scala 160:64:@32356.4]
  wire [14:0] _T_85052; // @[Modules.scala 160:64:@32358.4]
  wire [13:0] _T_85053; // @[Modules.scala 160:64:@32359.4]
  wire [13:0] buffer_9_620; // @[Modules.scala 160:64:@32360.4]
  wire [14:0] _T_85055; // @[Modules.scala 160:64:@32362.4]
  wire [13:0] _T_85056; // @[Modules.scala 160:64:@32363.4]
  wire [13:0] buffer_9_621; // @[Modules.scala 160:64:@32364.4]
  wire [14:0] _T_85058; // @[Modules.scala 160:64:@32366.4]
  wire [13:0] _T_85059; // @[Modules.scala 160:64:@32367.4]
  wire [13:0] buffer_9_622; // @[Modules.scala 160:64:@32368.4]
  wire [14:0] _T_85061; // @[Modules.scala 166:64:@32370.4]
  wire [13:0] _T_85062; // @[Modules.scala 166:64:@32371.4]
  wire [13:0] buffer_9_623; // @[Modules.scala 166:64:@32372.4]
  wire [14:0] _T_85064; // @[Modules.scala 166:64:@32374.4]
  wire [13:0] _T_85065; // @[Modules.scala 166:64:@32375.4]
  wire [13:0] buffer_9_624; // @[Modules.scala 166:64:@32376.4]
  wire [14:0] _T_85067; // @[Modules.scala 160:64:@32378.4]
  wire [13:0] _T_85068; // @[Modules.scala 160:64:@32379.4]
  wire [13:0] buffer_9_625; // @[Modules.scala 160:64:@32380.4]
  wire [14:0] _T_85070; // @[Modules.scala 172:66:@32382.4]
  wire [13:0] _T_85071; // @[Modules.scala 172:66:@32383.4]
  wire [13:0] buffer_9_626; // @[Modules.scala 172:66:@32384.4]
  wire [5:0] _GEN_694; // @[Modules.scala 150:103:@32545.4]
  wire [6:0] _T_85077; // @[Modules.scala 150:103:@32545.4]
  wire [5:0] _T_85078; // @[Modules.scala 150:103:@32546.4]
  wire [5:0] _T_85079; // @[Modules.scala 150:103:@32547.4]
  wire [5:0] _T_85084; // @[Modules.scala 150:103:@32551.4]
  wire [4:0] _T_85085; // @[Modules.scala 150:103:@32552.4]
  wire [4:0] _T_85086; // @[Modules.scala 150:103:@32553.4]
  wire [5:0] _GEN_695; // @[Modules.scala 150:103:@32557.4]
  wire [6:0] _T_85091; // @[Modules.scala 150:103:@32557.4]
  wire [5:0] _T_85092; // @[Modules.scala 150:103:@32558.4]
  wire [5:0] _T_85093; // @[Modules.scala 150:103:@32559.4]
  wire [6:0] _T_85098; // @[Modules.scala 150:103:@32563.4]
  wire [5:0] _T_85099; // @[Modules.scala 150:103:@32564.4]
  wire [5:0] _T_85100; // @[Modules.scala 150:103:@32565.4]
  wire [5:0] _GEN_696; // @[Modules.scala 150:103:@32599.4]
  wire [6:0] _T_85140; // @[Modules.scala 150:103:@32599.4]
  wire [5:0] _T_85141; // @[Modules.scala 150:103:@32600.4]
  wire [5:0] _T_85142; // @[Modules.scala 150:103:@32601.4]
  wire [5:0] _T_85154; // @[Modules.scala 150:103:@32611.4]
  wire [4:0] _T_85155; // @[Modules.scala 150:103:@32612.4]
  wire [4:0] _T_85156; // @[Modules.scala 150:103:@32613.4]
  wire [5:0] _T_85231; // @[Modules.scala 150:103:@32677.4]
  wire [4:0] _T_85232; // @[Modules.scala 150:103:@32678.4]
  wire [4:0] _T_85233; // @[Modules.scala 150:103:@32679.4]
  wire [6:0] _T_85252; // @[Modules.scala 150:103:@32695.4]
  wire [5:0] _T_85253; // @[Modules.scala 150:103:@32696.4]
  wire [5:0] _T_85254; // @[Modules.scala 150:103:@32697.4]
  wire [6:0] _T_85266; // @[Modules.scala 150:103:@32707.4]
  wire [5:0] _T_85267; // @[Modules.scala 150:103:@32708.4]
  wire [5:0] _T_85268; // @[Modules.scala 150:103:@32709.4]
  wire [5:0] _T_85322; // @[Modules.scala 150:103:@32755.4]
  wire [4:0] _T_85323; // @[Modules.scala 150:103:@32756.4]
  wire [4:0] _T_85324; // @[Modules.scala 150:103:@32757.4]
  wire [6:0] _T_85329; // @[Modules.scala 150:103:@32761.4]
  wire [5:0] _T_85330; // @[Modules.scala 150:103:@32762.4]
  wire [5:0] _T_85331; // @[Modules.scala 150:103:@32763.4]
  wire [6:0] _T_85357; // @[Modules.scala 150:103:@32785.4]
  wire [5:0] _T_85358; // @[Modules.scala 150:103:@32786.4]
  wire [5:0] _T_85359; // @[Modules.scala 150:103:@32787.4]
  wire [5:0] _T_85371; // @[Modules.scala 150:103:@32797.4]
  wire [4:0] _T_85372; // @[Modules.scala 150:103:@32798.4]
  wire [4:0] _T_85373; // @[Modules.scala 150:103:@32799.4]
  wire [5:0] _T_85378; // @[Modules.scala 150:103:@32803.4]
  wire [4:0] _T_85379; // @[Modules.scala 150:103:@32804.4]
  wire [4:0] _T_85380; // @[Modules.scala 150:103:@32805.4]
  wire [6:0] _T_85399; // @[Modules.scala 150:103:@32821.4]
  wire [5:0] _T_85400; // @[Modules.scala 150:103:@32822.4]
  wire [5:0] _T_85401; // @[Modules.scala 150:103:@32823.4]
  wire [5:0] _T_85406; // @[Modules.scala 150:103:@32827.4]
  wire [4:0] _T_85407; // @[Modules.scala 150:103:@32828.4]
  wire [4:0] _T_85408; // @[Modules.scala 150:103:@32829.4]
  wire [5:0] _T_85413; // @[Modules.scala 150:103:@32833.4]
  wire [4:0] _T_85414; // @[Modules.scala 150:103:@32834.4]
  wire [4:0] _T_85415; // @[Modules.scala 150:103:@32835.4]
  wire [5:0] _GEN_701; // @[Modules.scala 150:103:@32839.4]
  wire [6:0] _T_85420; // @[Modules.scala 150:103:@32839.4]
  wire [5:0] _T_85421; // @[Modules.scala 150:103:@32840.4]
  wire [5:0] _T_85422; // @[Modules.scala 150:103:@32841.4]
  wire [6:0] _T_85434; // @[Modules.scala 150:103:@32851.4]
  wire [5:0] _T_85435; // @[Modules.scala 150:103:@32852.4]
  wire [5:0] _T_85436; // @[Modules.scala 150:103:@32853.4]
  wire [6:0] _T_85469; // @[Modules.scala 150:103:@32881.4]
  wire [5:0] _T_85470; // @[Modules.scala 150:103:@32882.4]
  wire [5:0] _T_85471; // @[Modules.scala 150:103:@32883.4]
  wire [6:0] _T_85476; // @[Modules.scala 150:103:@32887.4]
  wire [5:0] _T_85477; // @[Modules.scala 150:103:@32888.4]
  wire [5:0] _T_85478; // @[Modules.scala 150:103:@32889.4]
  wire [5:0] _T_85490; // @[Modules.scala 150:103:@32899.4]
  wire [4:0] _T_85491; // @[Modules.scala 150:103:@32900.4]
  wire [4:0] _T_85492; // @[Modules.scala 150:103:@32901.4]
  wire [5:0] _GEN_703; // @[Modules.scala 150:103:@32923.4]
  wire [6:0] _T_85518; // @[Modules.scala 150:103:@32923.4]
  wire [5:0] _T_85519; // @[Modules.scala 150:103:@32924.4]
  wire [5:0] _T_85520; // @[Modules.scala 150:103:@32925.4]
  wire [5:0] _T_85525; // @[Modules.scala 150:103:@32929.4]
  wire [4:0] _T_85526; // @[Modules.scala 150:103:@32930.4]
  wire [4:0] _T_85527; // @[Modules.scala 150:103:@32931.4]
  wire [5:0] _T_85539; // @[Modules.scala 150:103:@32941.4]
  wire [4:0] _T_85540; // @[Modules.scala 150:103:@32942.4]
  wire [4:0] _T_85541; // @[Modules.scala 150:103:@32943.4]
  wire [5:0] _GEN_704; // @[Modules.scala 150:103:@32947.4]
  wire [6:0] _T_85546; // @[Modules.scala 150:103:@32947.4]
  wire [5:0] _T_85547; // @[Modules.scala 150:103:@32948.4]
  wire [5:0] _T_85548; // @[Modules.scala 150:103:@32949.4]
  wire [5:0] _GEN_705; // @[Modules.scala 150:103:@32953.4]
  wire [6:0] _T_85553; // @[Modules.scala 150:103:@32953.4]
  wire [5:0] _T_85554; // @[Modules.scala 150:103:@32954.4]
  wire [5:0] _T_85555; // @[Modules.scala 150:103:@32955.4]
  wire [5:0] _T_85588; // @[Modules.scala 150:103:@32983.4]
  wire [4:0] _T_85589; // @[Modules.scala 150:103:@32984.4]
  wire [4:0] _T_85590; // @[Modules.scala 150:103:@32985.4]
  wire [6:0] _T_85609; // @[Modules.scala 150:103:@33001.4]
  wire [5:0] _T_85610; // @[Modules.scala 150:103:@33002.4]
  wire [5:0] _T_85611; // @[Modules.scala 150:103:@33003.4]
  wire [5:0] _T_85616; // @[Modules.scala 150:103:@33007.4]
  wire [4:0] _T_85617; // @[Modules.scala 150:103:@33008.4]
  wire [4:0] _T_85618; // @[Modules.scala 150:103:@33009.4]
  wire [5:0] _T_85637; // @[Modules.scala 150:103:@33025.4]
  wire [4:0] _T_85638; // @[Modules.scala 150:103:@33026.4]
  wire [4:0] _T_85639; // @[Modules.scala 150:103:@33027.4]
  wire [5:0] _GEN_707; // @[Modules.scala 150:103:@33049.4]
  wire [6:0] _T_85665; // @[Modules.scala 150:103:@33049.4]
  wire [5:0] _T_85666; // @[Modules.scala 150:103:@33050.4]
  wire [5:0] _T_85667; // @[Modules.scala 150:103:@33051.4]
  wire [5:0] _GEN_709; // @[Modules.scala 150:103:@33073.4]
  wire [6:0] _T_85693; // @[Modules.scala 150:103:@33073.4]
  wire [5:0] _T_85694; // @[Modules.scala 150:103:@33074.4]
  wire [5:0] _T_85695; // @[Modules.scala 150:103:@33075.4]
  wire [5:0] _T_85707; // @[Modules.scala 150:103:@33085.4]
  wire [4:0] _T_85708; // @[Modules.scala 150:103:@33086.4]
  wire [4:0] _T_85709; // @[Modules.scala 150:103:@33087.4]
  wire [6:0] _T_85714; // @[Modules.scala 150:103:@33091.4]
  wire [5:0] _T_85715; // @[Modules.scala 150:103:@33092.4]
  wire [5:0] _T_85716; // @[Modules.scala 150:103:@33093.4]
  wire [6:0] _T_85728; // @[Modules.scala 150:103:@33103.4]
  wire [5:0] _T_85729; // @[Modules.scala 150:103:@33104.4]
  wire [5:0] _T_85730; // @[Modules.scala 150:103:@33105.4]
  wire [5:0] _T_85777; // @[Modules.scala 150:103:@33145.4]
  wire [4:0] _T_85778; // @[Modules.scala 150:103:@33146.4]
  wire [4:0] _T_85779; // @[Modules.scala 150:103:@33147.4]
  wire [6:0] _T_85805; // @[Modules.scala 150:103:@33169.4]
  wire [5:0] _T_85806; // @[Modules.scala 150:103:@33170.4]
  wire [5:0] _T_85807; // @[Modules.scala 150:103:@33171.4]
  wire [6:0] _T_85819; // @[Modules.scala 150:103:@33181.4]
  wire [5:0] _T_85820; // @[Modules.scala 150:103:@33182.4]
  wire [5:0] _T_85821; // @[Modules.scala 150:103:@33183.4]
  wire [5:0] _T_85840; // @[Modules.scala 150:103:@33199.4]
  wire [4:0] _T_85841; // @[Modules.scala 150:103:@33200.4]
  wire [4:0] _T_85842; // @[Modules.scala 150:103:@33201.4]
  wire [5:0] _T_85868; // @[Modules.scala 150:103:@33223.4]
  wire [4:0] _T_85869; // @[Modules.scala 150:103:@33224.4]
  wire [4:0] _T_85870; // @[Modules.scala 150:103:@33225.4]
  wire [5:0] _T_85875; // @[Modules.scala 150:103:@33229.4]
  wire [4:0] _T_85876; // @[Modules.scala 150:103:@33230.4]
  wire [4:0] _T_85877; // @[Modules.scala 150:103:@33231.4]
  wire [5:0] _T_85882; // @[Modules.scala 150:103:@33235.4]
  wire [4:0] _T_85883; // @[Modules.scala 150:103:@33236.4]
  wire [4:0] _T_85884; // @[Modules.scala 150:103:@33237.4]
  wire [6:0] _T_85924; // @[Modules.scala 150:103:@33271.4]
  wire [5:0] _T_85925; // @[Modules.scala 150:103:@33272.4]
  wire [5:0] _T_85926; // @[Modules.scala 150:103:@33273.4]
  wire [6:0] _T_85938; // @[Modules.scala 150:103:@33283.4]
  wire [5:0] _T_85939; // @[Modules.scala 150:103:@33284.4]
  wire [5:0] _T_85940; // @[Modules.scala 150:103:@33285.4]
  wire [6:0] _T_85987; // @[Modules.scala 150:103:@33325.4]
  wire [5:0] _T_85988; // @[Modules.scala 150:103:@33326.4]
  wire [5:0] _T_85989; // @[Modules.scala 150:103:@33327.4]
  wire [5:0] _GEN_719; // @[Modules.scala 150:103:@33337.4]
  wire [6:0] _T_86001; // @[Modules.scala 150:103:@33337.4]
  wire [5:0] _T_86002; // @[Modules.scala 150:103:@33338.4]
  wire [5:0] _T_86003; // @[Modules.scala 150:103:@33339.4]
  wire [6:0] _T_86015; // @[Modules.scala 150:103:@33349.4]
  wire [5:0] _T_86016; // @[Modules.scala 150:103:@33350.4]
  wire [5:0] _T_86017; // @[Modules.scala 150:103:@33351.4]
  wire [6:0] _T_86036; // @[Modules.scala 150:103:@33367.4]
  wire [5:0] _T_86037; // @[Modules.scala 150:103:@33368.4]
  wire [5:0] _T_86038; // @[Modules.scala 150:103:@33369.4]
  wire [6:0] _T_86106; // @[Modules.scala 150:103:@33427.4]
  wire [5:0] _T_86107; // @[Modules.scala 150:103:@33428.4]
  wire [5:0] _T_86108; // @[Modules.scala 150:103:@33429.4]
  wire [6:0] _T_86127; // @[Modules.scala 150:103:@33445.4]
  wire [5:0] _T_86128; // @[Modules.scala 150:103:@33446.4]
  wire [5:0] _T_86129; // @[Modules.scala 150:103:@33447.4]
  wire [6:0] _T_86134; // @[Modules.scala 150:103:@33451.4]
  wire [5:0] _T_86135; // @[Modules.scala 150:103:@33452.4]
  wire [5:0] _T_86136; // @[Modules.scala 150:103:@33453.4]
  wire [5:0] _T_86155; // @[Modules.scala 150:103:@33469.4]
  wire [4:0] _T_86156; // @[Modules.scala 150:103:@33470.4]
  wire [4:0] _T_86157; // @[Modules.scala 150:103:@33471.4]
  wire [5:0] _T_86204; // @[Modules.scala 150:103:@33511.4]
  wire [4:0] _T_86205; // @[Modules.scala 150:103:@33512.4]
  wire [4:0] _T_86206; // @[Modules.scala 150:103:@33513.4]
  wire [6:0] _T_86225; // @[Modules.scala 150:103:@33529.4]
  wire [5:0] _T_86226; // @[Modules.scala 150:103:@33530.4]
  wire [5:0] _T_86227; // @[Modules.scala 150:103:@33531.4]
  wire [5:0] _GEN_726; // @[Modules.scala 150:103:@33565.4]
  wire [6:0] _T_86267; // @[Modules.scala 150:103:@33565.4]
  wire [5:0] _T_86268; // @[Modules.scala 150:103:@33566.4]
  wire [5:0] _T_86269; // @[Modules.scala 150:103:@33567.4]
  wire [6:0] _T_86274; // @[Modules.scala 150:103:@33571.4]
  wire [5:0] _T_86275; // @[Modules.scala 150:103:@33572.4]
  wire [5:0] _T_86276; // @[Modules.scala 150:103:@33573.4]
  wire [5:0] _GEN_729; // @[Modules.scala 150:103:@33619.4]
  wire [6:0] _T_86330; // @[Modules.scala 150:103:@33619.4]
  wire [5:0] _T_86331; // @[Modules.scala 150:103:@33620.4]
  wire [5:0] _T_86332; // @[Modules.scala 150:103:@33621.4]
  wire [6:0] _T_86344; // @[Modules.scala 150:103:@33631.4]
  wire [5:0] _T_86345; // @[Modules.scala 150:103:@33632.4]
  wire [5:0] _T_86346; // @[Modules.scala 150:103:@33633.4]
  wire [5:0] _GEN_731; // @[Modules.scala 150:103:@33637.4]
  wire [6:0] _T_86351; // @[Modules.scala 150:103:@33637.4]
  wire [5:0] _T_86352; // @[Modules.scala 150:103:@33638.4]
  wire [5:0] _T_86353; // @[Modules.scala 150:103:@33639.4]
  wire [5:0] _GEN_732; // @[Modules.scala 150:103:@33655.4]
  wire [6:0] _T_86372; // @[Modules.scala 150:103:@33655.4]
  wire [5:0] _T_86373; // @[Modules.scala 150:103:@33656.4]
  wire [5:0] _T_86374; // @[Modules.scala 150:103:@33657.4]
  wire [5:0] _T_86379; // @[Modules.scala 150:103:@33661.4]
  wire [4:0] _T_86380; // @[Modules.scala 150:103:@33662.4]
  wire [4:0] _T_86381; // @[Modules.scala 150:103:@33663.4]
  wire [5:0] _T_86386; // @[Modules.scala 150:103:@33667.4]
  wire [4:0] _T_86387; // @[Modules.scala 150:103:@33668.4]
  wire [4:0] _T_86388; // @[Modules.scala 150:103:@33669.4]
  wire [5:0] _T_86393; // @[Modules.scala 150:103:@33673.4]
  wire [4:0] _T_86394; // @[Modules.scala 150:103:@33674.4]
  wire [4:0] _T_86395; // @[Modules.scala 150:103:@33675.4]
  wire [6:0] _T_86414; // @[Modules.scala 150:103:@33691.4]
  wire [5:0] _T_86415; // @[Modules.scala 150:103:@33692.4]
  wire [5:0] _T_86416; // @[Modules.scala 150:103:@33693.4]
  wire [6:0] _T_86456; // @[Modules.scala 150:103:@33727.4]
  wire [5:0] _T_86457; // @[Modules.scala 150:103:@33728.4]
  wire [5:0] _T_86458; // @[Modules.scala 150:103:@33729.4]
  wire [5:0] _T_86463; // @[Modules.scala 150:103:@33733.4]
  wire [4:0] _T_86464; // @[Modules.scala 150:103:@33734.4]
  wire [4:0] _T_86465; // @[Modules.scala 150:103:@33735.4]
  wire [5:0] _T_86470; // @[Modules.scala 150:103:@33739.4]
  wire [4:0] _T_86471; // @[Modules.scala 150:103:@33740.4]
  wire [4:0] _T_86472; // @[Modules.scala 150:103:@33741.4]
  wire [6:0] _T_86484; // @[Modules.scala 150:103:@33751.4]
  wire [5:0] _T_86485; // @[Modules.scala 150:103:@33752.4]
  wire [5:0] _T_86486; // @[Modules.scala 150:103:@33753.4]
  wire [5:0] _T_86491; // @[Modules.scala 150:103:@33757.4]
  wire [4:0] _T_86492; // @[Modules.scala 150:103:@33758.4]
  wire [4:0] _T_86493; // @[Modules.scala 150:103:@33759.4]
  wire [5:0] _T_86568; // @[Modules.scala 150:103:@33823.4]
  wire [4:0] _T_86569; // @[Modules.scala 150:103:@33824.4]
  wire [4:0] _T_86570; // @[Modules.scala 150:103:@33825.4]
  wire [5:0] _GEN_738; // @[Modules.scala 150:103:@33859.4]
  wire [6:0] _T_86610; // @[Modules.scala 150:103:@33859.4]
  wire [5:0] _T_86611; // @[Modules.scala 150:103:@33860.4]
  wire [5:0] _T_86612; // @[Modules.scala 150:103:@33861.4]
  wire [5:0] _GEN_739; // @[Modules.scala 150:103:@33871.4]
  wire [6:0] _T_86624; // @[Modules.scala 150:103:@33871.4]
  wire [5:0] _T_86625; // @[Modules.scala 150:103:@33872.4]
  wire [5:0] _T_86626; // @[Modules.scala 150:103:@33873.4]
  wire [6:0] _T_86659; // @[Modules.scala 150:103:@33901.4]
  wire [5:0] _T_86660; // @[Modules.scala 150:103:@33902.4]
  wire [5:0] _T_86661; // @[Modules.scala 150:103:@33903.4]
  wire [5:0] _GEN_742; // @[Modules.scala 150:103:@33919.4]
  wire [6:0] _T_86680; // @[Modules.scala 150:103:@33919.4]
  wire [5:0] _T_86681; // @[Modules.scala 150:103:@33920.4]
  wire [5:0] _T_86682; // @[Modules.scala 150:103:@33921.4]
  wire [5:0] _T_86687; // @[Modules.scala 150:103:@33925.4]
  wire [4:0] _T_86688; // @[Modules.scala 150:103:@33926.4]
  wire [4:0] _T_86689; // @[Modules.scala 150:103:@33927.4]
  wire [6:0] _T_86694; // @[Modules.scala 150:103:@33931.4]
  wire [5:0] _T_86695; // @[Modules.scala 150:103:@33932.4]
  wire [5:0] _T_86696; // @[Modules.scala 150:103:@33933.4]
  wire [6:0] _T_86708; // @[Modules.scala 150:103:@33943.4]
  wire [5:0] _T_86709; // @[Modules.scala 150:103:@33944.4]
  wire [5:0] _T_86710; // @[Modules.scala 150:103:@33945.4]
  wire [6:0] _T_86736; // @[Modules.scala 150:103:@33967.4]
  wire [5:0] _T_86737; // @[Modules.scala 150:103:@33968.4]
  wire [5:0] _T_86738; // @[Modules.scala 150:103:@33969.4]
  wire [5:0] _T_86757; // @[Modules.scala 150:103:@33985.4]
  wire [4:0] _T_86758; // @[Modules.scala 150:103:@33986.4]
  wire [4:0] _T_86759; // @[Modules.scala 150:103:@33987.4]
  wire [6:0] _T_86764; // @[Modules.scala 150:103:@33991.4]
  wire [5:0] _T_86765; // @[Modules.scala 150:103:@33992.4]
  wire [5:0] _T_86766; // @[Modules.scala 150:103:@33993.4]
  wire [6:0] _T_86785; // @[Modules.scala 150:103:@34009.4]
  wire [5:0] _T_86786; // @[Modules.scala 150:103:@34010.4]
  wire [5:0] _T_86787; // @[Modules.scala 150:103:@34011.4]
  wire [6:0] _T_86834; // @[Modules.scala 150:103:@34051.4]
  wire [5:0] _T_86835; // @[Modules.scala 150:103:@34052.4]
  wire [5:0] _T_86836; // @[Modules.scala 150:103:@34053.4]
  wire [5:0] _T_86841; // @[Modules.scala 150:103:@34057.4]
  wire [4:0] _T_86842; // @[Modules.scala 150:103:@34058.4]
  wire [4:0] _T_86843; // @[Modules.scala 150:103:@34059.4]
  wire [6:0] _T_86862; // @[Modules.scala 150:103:@34075.4]
  wire [5:0] _T_86863; // @[Modules.scala 150:103:@34076.4]
  wire [5:0] _T_86864; // @[Modules.scala 150:103:@34077.4]
  wire [5:0] _T_86869; // @[Modules.scala 150:103:@34081.4]
  wire [4:0] _T_86870; // @[Modules.scala 150:103:@34082.4]
  wire [4:0] _T_86871; // @[Modules.scala 150:103:@34083.4]
  wire [5:0] _T_86883; // @[Modules.scala 150:103:@34093.4]
  wire [4:0] _T_86884; // @[Modules.scala 150:103:@34094.4]
  wire [4:0] _T_86885; // @[Modules.scala 150:103:@34095.4]
  wire [5:0] _GEN_749; // @[Modules.scala 150:103:@34117.4]
  wire [6:0] _T_86911; // @[Modules.scala 150:103:@34117.4]
  wire [5:0] _T_86912; // @[Modules.scala 150:103:@34118.4]
  wire [5:0] _T_86913; // @[Modules.scala 150:103:@34119.4]
  wire [6:0] _T_86918; // @[Modules.scala 150:103:@34123.4]
  wire [5:0] _T_86919; // @[Modules.scala 150:103:@34124.4]
  wire [5:0] _T_86920; // @[Modules.scala 150:103:@34125.4]
  wire [6:0] _T_86974; // @[Modules.scala 150:103:@34171.4]
  wire [5:0] _T_86975; // @[Modules.scala 150:103:@34172.4]
  wire [5:0] _T_86976; // @[Modules.scala 150:103:@34173.4]
  wire [6:0] _T_86981; // @[Modules.scala 150:103:@34177.4]
  wire [5:0] _T_86982; // @[Modules.scala 150:103:@34178.4]
  wire [5:0] _T_86983; // @[Modules.scala 150:103:@34179.4]
  wire [6:0] _T_87009; // @[Modules.scala 150:103:@34201.4]
  wire [5:0] _T_87010; // @[Modules.scala 150:103:@34202.4]
  wire [5:0] _T_87011; // @[Modules.scala 150:103:@34203.4]
  wire [6:0] _T_87016; // @[Modules.scala 150:103:@34207.4]
  wire [5:0] _T_87017; // @[Modules.scala 150:103:@34208.4]
  wire [5:0] _T_87018; // @[Modules.scala 150:103:@34209.4]
  wire [5:0] _T_87023; // @[Modules.scala 150:103:@34213.4]
  wire [4:0] _T_87024; // @[Modules.scala 150:103:@34214.4]
  wire [4:0] _T_87025; // @[Modules.scala 150:103:@34215.4]
  wire [5:0] _GEN_753; // @[Modules.scala 150:103:@34267.4]
  wire [6:0] _T_87086; // @[Modules.scala 150:103:@34267.4]
  wire [5:0] _T_87087; // @[Modules.scala 150:103:@34268.4]
  wire [5:0] _T_87088; // @[Modules.scala 150:103:@34269.4]
  wire [5:0] _GEN_756; // @[Modules.scala 150:103:@34291.4]
  wire [6:0] _T_87114; // @[Modules.scala 150:103:@34291.4]
  wire [5:0] _T_87115; // @[Modules.scala 150:103:@34292.4]
  wire [5:0] _T_87116; // @[Modules.scala 150:103:@34293.4]
  wire [5:0] _GEN_757; // @[Modules.scala 150:103:@34297.4]
  wire [6:0] _T_87121; // @[Modules.scala 150:103:@34297.4]
  wire [5:0] _T_87122; // @[Modules.scala 150:103:@34298.4]
  wire [5:0] _T_87123; // @[Modules.scala 150:103:@34299.4]
  wire [5:0] _T_87163; // @[Modules.scala 150:103:@34333.4]
  wire [4:0] _T_87164; // @[Modules.scala 150:103:@34334.4]
  wire [4:0] _T_87165; // @[Modules.scala 150:103:@34335.4]
  wire [6:0] _T_87170; // @[Modules.scala 150:103:@34339.4]
  wire [5:0] _T_87171; // @[Modules.scala 150:103:@34340.4]
  wire [5:0] _T_87172; // @[Modules.scala 150:103:@34341.4]
  wire [5:0] _GEN_759; // @[Modules.scala 150:103:@34345.4]
  wire [6:0] _T_87177; // @[Modules.scala 150:103:@34345.4]
  wire [5:0] _T_87178; // @[Modules.scala 150:103:@34346.4]
  wire [5:0] _T_87179; // @[Modules.scala 150:103:@34347.4]
  wire [13:0] buffer_10_0; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87224; // @[Modules.scala 160:64:@34387.4]
  wire [13:0] _T_87225; // @[Modules.scala 160:64:@34388.4]
  wire [13:0] buffer_10_308; // @[Modules.scala 160:64:@34389.4]
  wire [13:0] buffer_10_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87227; // @[Modules.scala 160:64:@34391.4]
  wire [13:0] _T_87228; // @[Modules.scala 160:64:@34392.4]
  wire [13:0] buffer_10_309; // @[Modules.scala 160:64:@34393.4]
  wire [14:0] _T_87233; // @[Modules.scala 160:64:@34399.4]
  wire [13:0] _T_87234; // @[Modules.scala 160:64:@34400.4]
  wire [13:0] buffer_10_311; // @[Modules.scala 160:64:@34401.4]
  wire [13:0] buffer_10_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87236; // @[Modules.scala 160:64:@34403.4]
  wire [13:0] _T_87237; // @[Modules.scala 160:64:@34404.4]
  wire [13:0] buffer_10_312; // @[Modules.scala 160:64:@34405.4]
  wire [13:0] buffer_10_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87239; // @[Modules.scala 160:64:@34407.4]
  wire [13:0] _T_87240; // @[Modules.scala 160:64:@34408.4]
  wire [13:0] buffer_10_313; // @[Modules.scala 160:64:@34409.4]
  wire [14:0] _T_87254; // @[Modules.scala 160:64:@34427.4]
  wire [13:0] _T_87255; // @[Modules.scala 160:64:@34428.4]
  wire [13:0] buffer_10_318; // @[Modules.scala 160:64:@34429.4]
  wire [13:0] buffer_10_22; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87257; // @[Modules.scala 160:64:@34431.4]
  wire [13:0] _T_87258; // @[Modules.scala 160:64:@34432.4]
  wire [13:0] buffer_10_319; // @[Modules.scala 160:64:@34433.4]
  wire [13:0] buffer_10_25; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87260; // @[Modules.scala 160:64:@34435.4]
  wire [13:0] _T_87261; // @[Modules.scala 160:64:@34436.4]
  wire [13:0] buffer_10_320; // @[Modules.scala 160:64:@34437.4]
  wire [13:0] buffer_10_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87263; // @[Modules.scala 160:64:@34439.4]
  wire [13:0] _T_87264; // @[Modules.scala 160:64:@34440.4]
  wire [13:0] buffer_10_321; // @[Modules.scala 160:64:@34441.4]
  wire [14:0] _T_87266; // @[Modules.scala 160:64:@34443.4]
  wire [13:0] _T_87267; // @[Modules.scala 160:64:@34444.4]
  wire [13:0] buffer_10_322; // @[Modules.scala 160:64:@34445.4]
  wire [14:0] _T_87272; // @[Modules.scala 160:64:@34451.4]
  wire [13:0] _T_87273; // @[Modules.scala 160:64:@34452.4]
  wire [13:0] buffer_10_324; // @[Modules.scala 160:64:@34453.4]
  wire [13:0] buffer_10_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87275; // @[Modules.scala 160:64:@34455.4]
  wire [13:0] _T_87276; // @[Modules.scala 160:64:@34456.4]
  wire [13:0] buffer_10_325; // @[Modules.scala 160:64:@34457.4]
  wire [13:0] buffer_10_36; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87278; // @[Modules.scala 160:64:@34459.4]
  wire [13:0] _T_87279; // @[Modules.scala 160:64:@34460.4]
  wire [13:0] buffer_10_326; // @[Modules.scala 160:64:@34461.4]
  wire [14:0] _T_87281; // @[Modules.scala 160:64:@34463.4]
  wire [13:0] _T_87282; // @[Modules.scala 160:64:@34464.4]
  wire [13:0] buffer_10_327; // @[Modules.scala 160:64:@34465.4]
  wire [13:0] buffer_10_40; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87284; // @[Modules.scala 160:64:@34467.4]
  wire [13:0] _T_87285; // @[Modules.scala 160:64:@34468.4]
  wire [13:0] buffer_10_328; // @[Modules.scala 160:64:@34469.4]
  wire [13:0] buffer_10_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87287; // @[Modules.scala 160:64:@34471.4]
  wire [13:0] _T_87288; // @[Modules.scala 160:64:@34472.4]
  wire [13:0] buffer_10_329; // @[Modules.scala 160:64:@34473.4]
  wire [13:0] buffer_10_46; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_47; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87293; // @[Modules.scala 160:64:@34479.4]
  wire [13:0] _T_87294; // @[Modules.scala 160:64:@34480.4]
  wire [13:0] buffer_10_331; // @[Modules.scala 160:64:@34481.4]
  wire [13:0] buffer_10_48; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87296; // @[Modules.scala 160:64:@34483.4]
  wire [13:0] _T_87297; // @[Modules.scala 160:64:@34484.4]
  wire [13:0] buffer_10_332; // @[Modules.scala 160:64:@34485.4]
  wire [13:0] buffer_10_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87299; // @[Modules.scala 160:64:@34487.4]
  wire [13:0] _T_87300; // @[Modules.scala 160:64:@34488.4]
  wire [13:0] buffer_10_333; // @[Modules.scala 160:64:@34489.4]
  wire [13:0] buffer_10_56; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87308; // @[Modules.scala 160:64:@34499.4]
  wire [13:0] _T_87309; // @[Modules.scala 160:64:@34500.4]
  wire [13:0] buffer_10_336; // @[Modules.scala 160:64:@34501.4]
  wire [13:0] buffer_10_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87311; // @[Modules.scala 160:64:@34503.4]
  wire [13:0] _T_87312; // @[Modules.scala 160:64:@34504.4]
  wire [13:0] buffer_10_337; // @[Modules.scala 160:64:@34505.4]
  wire [14:0] _T_87314; // @[Modules.scala 160:64:@34507.4]
  wire [13:0] _T_87315; // @[Modules.scala 160:64:@34508.4]
  wire [13:0] buffer_10_338; // @[Modules.scala 160:64:@34509.4]
  wire [13:0] buffer_10_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87317; // @[Modules.scala 160:64:@34511.4]
  wire [13:0] _T_87318; // @[Modules.scala 160:64:@34512.4]
  wire [13:0] buffer_10_339; // @[Modules.scala 160:64:@34513.4]
  wire [13:0] buffer_10_64; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87320; // @[Modules.scala 160:64:@34515.4]
  wire [13:0] _T_87321; // @[Modules.scala 160:64:@34516.4]
  wire [13:0] buffer_10_340; // @[Modules.scala 160:64:@34517.4]
  wire [13:0] buffer_10_66; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87323; // @[Modules.scala 160:64:@34519.4]
  wire [13:0] _T_87324; // @[Modules.scala 160:64:@34520.4]
  wire [13:0] buffer_10_341; // @[Modules.scala 160:64:@34521.4]
  wire [13:0] buffer_10_68; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87326; // @[Modules.scala 160:64:@34523.4]
  wire [13:0] _T_87327; // @[Modules.scala 160:64:@34524.4]
  wire [13:0] buffer_10_342; // @[Modules.scala 160:64:@34525.4]
  wire [14:0] _T_87329; // @[Modules.scala 160:64:@34527.4]
  wire [13:0] _T_87330; // @[Modules.scala 160:64:@34528.4]
  wire [13:0] buffer_10_343; // @[Modules.scala 160:64:@34529.4]
  wire [13:0] buffer_10_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87332; // @[Modules.scala 160:64:@34531.4]
  wire [13:0] _T_87333; // @[Modules.scala 160:64:@34532.4]
  wire [13:0] buffer_10_344; // @[Modules.scala 160:64:@34533.4]
  wire [13:0] buffer_10_76; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87338; // @[Modules.scala 160:64:@34539.4]
  wire [13:0] _T_87339; // @[Modules.scala 160:64:@34540.4]
  wire [13:0] buffer_10_346; // @[Modules.scala 160:64:@34541.4]
  wire [14:0] _T_87341; // @[Modules.scala 160:64:@34543.4]
  wire [13:0] _T_87342; // @[Modules.scala 160:64:@34544.4]
  wire [13:0] buffer_10_347; // @[Modules.scala 160:64:@34545.4]
  wire [13:0] buffer_10_80; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87344; // @[Modules.scala 160:64:@34547.4]
  wire [13:0] _T_87345; // @[Modules.scala 160:64:@34548.4]
  wire [13:0] buffer_10_348; // @[Modules.scala 160:64:@34549.4]
  wire [13:0] buffer_10_84; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87350; // @[Modules.scala 160:64:@34555.4]
  wire [13:0] _T_87351; // @[Modules.scala 160:64:@34556.4]
  wire [13:0] buffer_10_350; // @[Modules.scala 160:64:@34557.4]
  wire [14:0] _T_87353; // @[Modules.scala 160:64:@34559.4]
  wire [13:0] _T_87354; // @[Modules.scala 160:64:@34560.4]
  wire [13:0] buffer_10_351; // @[Modules.scala 160:64:@34561.4]
  wire [13:0] buffer_10_88; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87356; // @[Modules.scala 160:64:@34563.4]
  wire [13:0] _T_87357; // @[Modules.scala 160:64:@34564.4]
  wire [13:0] buffer_10_352; // @[Modules.scala 160:64:@34565.4]
  wire [13:0] buffer_10_90; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87359; // @[Modules.scala 160:64:@34567.4]
  wire [13:0] _T_87360; // @[Modules.scala 160:64:@34568.4]
  wire [13:0] buffer_10_353; // @[Modules.scala 160:64:@34569.4]
  wire [13:0] buffer_10_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87362; // @[Modules.scala 160:64:@34571.4]
  wire [13:0] _T_87363; // @[Modules.scala 160:64:@34572.4]
  wire [13:0] buffer_10_354; // @[Modules.scala 160:64:@34573.4]
  wire [14:0] _T_87365; // @[Modules.scala 160:64:@34575.4]
  wire [13:0] _T_87366; // @[Modules.scala 160:64:@34576.4]
  wire [13:0] buffer_10_355; // @[Modules.scala 160:64:@34577.4]
  wire [14:0] _T_87371; // @[Modules.scala 160:64:@34583.4]
  wire [13:0] _T_87372; // @[Modules.scala 160:64:@34584.4]
  wire [13:0] buffer_10_357; // @[Modules.scala 160:64:@34585.4]
  wire [13:0] buffer_10_100; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87374; // @[Modules.scala 160:64:@34587.4]
  wire [13:0] _T_87375; // @[Modules.scala 160:64:@34588.4]
  wire [13:0] buffer_10_358; // @[Modules.scala 160:64:@34589.4]
  wire [13:0] buffer_10_104; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87380; // @[Modules.scala 160:64:@34595.4]
  wire [13:0] _T_87381; // @[Modules.scala 160:64:@34596.4]
  wire [13:0] buffer_10_360; // @[Modules.scala 160:64:@34597.4]
  wire [13:0] buffer_10_106; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87383; // @[Modules.scala 160:64:@34599.4]
  wire [13:0] _T_87384; // @[Modules.scala 160:64:@34600.4]
  wire [13:0] buffer_10_361; // @[Modules.scala 160:64:@34601.4]
  wire [13:0] buffer_10_109; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87386; // @[Modules.scala 160:64:@34603.4]
  wire [13:0] _T_87387; // @[Modules.scala 160:64:@34604.4]
  wire [13:0] buffer_10_362; // @[Modules.scala 160:64:@34605.4]
  wire [14:0] _T_87389; // @[Modules.scala 160:64:@34607.4]
  wire [13:0] _T_87390; // @[Modules.scala 160:64:@34608.4]
  wire [13:0] buffer_10_363; // @[Modules.scala 160:64:@34609.4]
  wire [13:0] buffer_10_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87392; // @[Modules.scala 160:64:@34611.4]
  wire [13:0] _T_87393; // @[Modules.scala 160:64:@34612.4]
  wire [13:0] buffer_10_364; // @[Modules.scala 160:64:@34613.4]
  wire [13:0] buffer_10_114; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87395; // @[Modules.scala 160:64:@34615.4]
  wire [13:0] _T_87396; // @[Modules.scala 160:64:@34616.4]
  wire [13:0] buffer_10_365; // @[Modules.scala 160:64:@34617.4]
  wire [14:0] _T_87398; // @[Modules.scala 160:64:@34619.4]
  wire [13:0] _T_87399; // @[Modules.scala 160:64:@34620.4]
  wire [13:0] buffer_10_366; // @[Modules.scala 160:64:@34621.4]
  wire [14:0] _T_87401; // @[Modules.scala 160:64:@34623.4]
  wire [13:0] _T_87402; // @[Modules.scala 160:64:@34624.4]
  wire [13:0] buffer_10_367; // @[Modules.scala 160:64:@34625.4]
  wire [13:0] buffer_10_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87404; // @[Modules.scala 160:64:@34627.4]
  wire [13:0] _T_87405; // @[Modules.scala 160:64:@34628.4]
  wire [13:0] buffer_10_368; // @[Modules.scala 160:64:@34629.4]
  wire [13:0] buffer_10_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87407; // @[Modules.scala 160:64:@34631.4]
  wire [13:0] _T_87408; // @[Modules.scala 160:64:@34632.4]
  wire [13:0] buffer_10_369; // @[Modules.scala 160:64:@34633.4]
  wire [14:0] _T_87410; // @[Modules.scala 160:64:@34635.4]
  wire [13:0] _T_87411; // @[Modules.scala 160:64:@34636.4]
  wire [13:0] buffer_10_370; // @[Modules.scala 160:64:@34637.4]
  wire [14:0] _T_87413; // @[Modules.scala 160:64:@34639.4]
  wire [13:0] _T_87414; // @[Modules.scala 160:64:@34640.4]
  wire [13:0] buffer_10_371; // @[Modules.scala 160:64:@34641.4]
  wire [13:0] buffer_10_130; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87419; // @[Modules.scala 160:64:@34647.4]
  wire [13:0] _T_87420; // @[Modules.scala 160:64:@34648.4]
  wire [13:0] buffer_10_373; // @[Modules.scala 160:64:@34649.4]
  wire [13:0] buffer_10_132; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87422; // @[Modules.scala 160:64:@34651.4]
  wire [13:0] _T_87423; // @[Modules.scala 160:64:@34652.4]
  wire [13:0] buffer_10_374; // @[Modules.scala 160:64:@34653.4]
  wire [13:0] buffer_10_134; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87425; // @[Modules.scala 160:64:@34655.4]
  wire [13:0] _T_87426; // @[Modules.scala 160:64:@34656.4]
  wire [13:0] buffer_10_375; // @[Modules.scala 160:64:@34657.4]
  wire [13:0] buffer_10_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87428; // @[Modules.scala 160:64:@34659.4]
  wire [13:0] _T_87429; // @[Modules.scala 160:64:@34660.4]
  wire [13:0] buffer_10_376; // @[Modules.scala 160:64:@34661.4]
  wire [14:0] _T_87434; // @[Modules.scala 160:64:@34667.4]
  wire [13:0] _T_87435; // @[Modules.scala 160:64:@34668.4]
  wire [13:0] buffer_10_378; // @[Modules.scala 160:64:@34669.4]
  wire [14:0] _T_87440; // @[Modules.scala 160:64:@34675.4]
  wire [13:0] _T_87441; // @[Modules.scala 160:64:@34676.4]
  wire [13:0] buffer_10_380; // @[Modules.scala 160:64:@34677.4]
  wire [13:0] buffer_10_147; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87443; // @[Modules.scala 160:64:@34679.4]
  wire [13:0] _T_87444; // @[Modules.scala 160:64:@34680.4]
  wire [13:0] buffer_10_381; // @[Modules.scala 160:64:@34681.4]
  wire [13:0] buffer_10_150; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_151; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87449; // @[Modules.scala 160:64:@34687.4]
  wire [13:0] _T_87450; // @[Modules.scala 160:64:@34688.4]
  wire [13:0] buffer_10_383; // @[Modules.scala 160:64:@34689.4]
  wire [13:0] buffer_10_154; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87455; // @[Modules.scala 160:64:@34695.4]
  wire [13:0] _T_87456; // @[Modules.scala 160:64:@34696.4]
  wire [13:0] buffer_10_385; // @[Modules.scala 160:64:@34697.4]
  wire [14:0] _T_87461; // @[Modules.scala 160:64:@34703.4]
  wire [13:0] _T_87462; // @[Modules.scala 160:64:@34704.4]
  wire [13:0] buffer_10_387; // @[Modules.scala 160:64:@34705.4]
  wire [13:0] buffer_10_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87464; // @[Modules.scala 160:64:@34707.4]
  wire [13:0] _T_87465; // @[Modules.scala 160:64:@34708.4]
  wire [13:0] buffer_10_388; // @[Modules.scala 160:64:@34709.4]
  wire [13:0] buffer_10_164; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87470; // @[Modules.scala 160:64:@34715.4]
  wire [13:0] _T_87471; // @[Modules.scala 160:64:@34716.4]
  wire [13:0] buffer_10_390; // @[Modules.scala 160:64:@34717.4]
  wire [14:0] _T_87473; // @[Modules.scala 160:64:@34719.4]
  wire [13:0] _T_87474; // @[Modules.scala 160:64:@34720.4]
  wire [13:0] buffer_10_391; // @[Modules.scala 160:64:@34721.4]
  wire [14:0] _T_87476; // @[Modules.scala 160:64:@34723.4]
  wire [13:0] _T_87477; // @[Modules.scala 160:64:@34724.4]
  wire [13:0] buffer_10_392; // @[Modules.scala 160:64:@34725.4]
  wire [13:0] buffer_10_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87479; // @[Modules.scala 160:64:@34727.4]
  wire [13:0] _T_87480; // @[Modules.scala 160:64:@34728.4]
  wire [13:0] buffer_10_393; // @[Modules.scala 160:64:@34729.4]
  wire [14:0] _T_87482; // @[Modules.scala 160:64:@34731.4]
  wire [13:0] _T_87483; // @[Modules.scala 160:64:@34732.4]
  wire [13:0] buffer_10_394; // @[Modules.scala 160:64:@34733.4]
  wire [14:0] _T_87488; // @[Modules.scala 160:64:@34739.4]
  wire [13:0] _T_87489; // @[Modules.scala 160:64:@34740.4]
  wire [13:0] buffer_10_396; // @[Modules.scala 160:64:@34741.4]
  wire [13:0] buffer_10_179; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87491; // @[Modules.scala 160:64:@34743.4]
  wire [13:0] _T_87492; // @[Modules.scala 160:64:@34744.4]
  wire [13:0] buffer_10_397; // @[Modules.scala 160:64:@34745.4]
  wire [13:0] buffer_10_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87494; // @[Modules.scala 160:64:@34747.4]
  wire [13:0] _T_87495; // @[Modules.scala 160:64:@34748.4]
  wire [13:0] buffer_10_398; // @[Modules.scala 160:64:@34749.4]
  wire [13:0] buffer_10_182; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87497; // @[Modules.scala 160:64:@34751.4]
  wire [13:0] _T_87498; // @[Modules.scala 160:64:@34752.4]
  wire [13:0] buffer_10_399; // @[Modules.scala 160:64:@34753.4]
  wire [13:0] buffer_10_185; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87500; // @[Modules.scala 160:64:@34755.4]
  wire [13:0] _T_87501; // @[Modules.scala 160:64:@34756.4]
  wire [13:0] buffer_10_400; // @[Modules.scala 160:64:@34757.4]
  wire [13:0] buffer_10_186; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_187; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87503; // @[Modules.scala 160:64:@34759.4]
  wire [13:0] _T_87504; // @[Modules.scala 160:64:@34760.4]
  wire [13:0] buffer_10_401; // @[Modules.scala 160:64:@34761.4]
  wire [13:0] buffer_10_188; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87506; // @[Modules.scala 160:64:@34763.4]
  wire [13:0] _T_87507; // @[Modules.scala 160:64:@34764.4]
  wire [13:0] buffer_10_402; // @[Modules.scala 160:64:@34765.4]
  wire [13:0] buffer_10_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87509; // @[Modules.scala 160:64:@34767.4]
  wire [13:0] _T_87510; // @[Modules.scala 160:64:@34768.4]
  wire [13:0] buffer_10_403; // @[Modules.scala 160:64:@34769.4]
  wire [14:0] _T_87512; // @[Modules.scala 160:64:@34771.4]
  wire [13:0] _T_87513; // @[Modules.scala 160:64:@34772.4]
  wire [13:0] buffer_10_404; // @[Modules.scala 160:64:@34773.4]
  wire [14:0] _T_87515; // @[Modules.scala 160:64:@34775.4]
  wire [13:0] _T_87516; // @[Modules.scala 160:64:@34776.4]
  wire [13:0] buffer_10_405; // @[Modules.scala 160:64:@34777.4]
  wire [13:0] buffer_10_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87518; // @[Modules.scala 160:64:@34779.4]
  wire [13:0] _T_87519; // @[Modules.scala 160:64:@34780.4]
  wire [13:0] buffer_10_406; // @[Modules.scala 160:64:@34781.4]
  wire [13:0] buffer_10_198; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87521; // @[Modules.scala 160:64:@34783.4]
  wire [13:0] _T_87522; // @[Modules.scala 160:64:@34784.4]
  wire [13:0] buffer_10_407; // @[Modules.scala 160:64:@34785.4]
  wire [13:0] buffer_10_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87524; // @[Modules.scala 160:64:@34787.4]
  wire [13:0] _T_87525; // @[Modules.scala 160:64:@34788.4]
  wire [13:0] buffer_10_408; // @[Modules.scala 160:64:@34789.4]
  wire [13:0] buffer_10_202; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87527; // @[Modules.scala 160:64:@34791.4]
  wire [13:0] _T_87528; // @[Modules.scala 160:64:@34792.4]
  wire [13:0] buffer_10_409; // @[Modules.scala 160:64:@34793.4]
  wire [14:0] _T_87530; // @[Modules.scala 160:64:@34795.4]
  wire [13:0] _T_87531; // @[Modules.scala 160:64:@34796.4]
  wire [13:0] buffer_10_410; // @[Modules.scala 160:64:@34797.4]
  wire [14:0] _T_87533; // @[Modules.scala 160:64:@34799.4]
  wire [13:0] _T_87534; // @[Modules.scala 160:64:@34800.4]
  wire [13:0] buffer_10_411; // @[Modules.scala 160:64:@34801.4]
  wire [14:0] _T_87536; // @[Modules.scala 160:64:@34803.4]
  wire [13:0] _T_87537; // @[Modules.scala 160:64:@34804.4]
  wire [13:0] buffer_10_412; // @[Modules.scala 160:64:@34805.4]
  wire [13:0] buffer_10_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87542; // @[Modules.scala 160:64:@34811.4]
  wire [13:0] _T_87543; // @[Modules.scala 160:64:@34812.4]
  wire [13:0] buffer_10_414; // @[Modules.scala 160:64:@34813.4]
  wire [13:0] buffer_10_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87551; // @[Modules.scala 160:64:@34823.4]
  wire [13:0] _T_87552; // @[Modules.scala 160:64:@34824.4]
  wire [13:0] buffer_10_417; // @[Modules.scala 160:64:@34825.4]
  wire [13:0] buffer_10_221; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87554; // @[Modules.scala 160:64:@34827.4]
  wire [13:0] _T_87555; // @[Modules.scala 160:64:@34828.4]
  wire [13:0] buffer_10_418; // @[Modules.scala 160:64:@34829.4]
  wire [13:0] buffer_10_226; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87563; // @[Modules.scala 160:64:@34839.4]
  wire [13:0] _T_87564; // @[Modules.scala 160:64:@34840.4]
  wire [13:0] buffer_10_421; // @[Modules.scala 160:64:@34841.4]
  wire [13:0] buffer_10_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87566; // @[Modules.scala 160:64:@34843.4]
  wire [13:0] _T_87567; // @[Modules.scala 160:64:@34844.4]
  wire [13:0] buffer_10_422; // @[Modules.scala 160:64:@34845.4]
  wire [13:0] buffer_10_230; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87569; // @[Modules.scala 160:64:@34847.4]
  wire [13:0] _T_87570; // @[Modules.scala 160:64:@34848.4]
  wire [13:0] buffer_10_423; // @[Modules.scala 160:64:@34849.4]
  wire [13:0] buffer_10_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87572; // @[Modules.scala 160:64:@34851.4]
  wire [13:0] _T_87573; // @[Modules.scala 160:64:@34852.4]
  wire [13:0] buffer_10_424; // @[Modules.scala 160:64:@34853.4]
  wire [14:0] _T_87575; // @[Modules.scala 160:64:@34855.4]
  wire [13:0] _T_87576; // @[Modules.scala 160:64:@34856.4]
  wire [13:0] buffer_10_425; // @[Modules.scala 160:64:@34857.4]
  wire [13:0] buffer_10_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87578; // @[Modules.scala 160:64:@34859.4]
  wire [13:0] _T_87579; // @[Modules.scala 160:64:@34860.4]
  wire [13:0] buffer_10_426; // @[Modules.scala 160:64:@34861.4]
  wire [14:0] _T_87581; // @[Modules.scala 160:64:@34863.4]
  wire [13:0] _T_87582; // @[Modules.scala 160:64:@34864.4]
  wire [13:0] buffer_10_427; // @[Modules.scala 160:64:@34865.4]
  wire [13:0] buffer_10_240; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87584; // @[Modules.scala 160:64:@34867.4]
  wire [13:0] _T_87585; // @[Modules.scala 160:64:@34868.4]
  wire [13:0] buffer_10_428; // @[Modules.scala 160:64:@34869.4]
  wire [14:0] _T_87587; // @[Modules.scala 160:64:@34871.4]
  wire [13:0] _T_87588; // @[Modules.scala 160:64:@34872.4]
  wire [13:0] buffer_10_429; // @[Modules.scala 160:64:@34873.4]
  wire [13:0] buffer_10_244; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87590; // @[Modules.scala 160:64:@34875.4]
  wire [13:0] _T_87591; // @[Modules.scala 160:64:@34876.4]
  wire [13:0] buffer_10_430; // @[Modules.scala 160:64:@34877.4]
  wire [14:0] _T_87593; // @[Modules.scala 160:64:@34879.4]
  wire [13:0] _T_87594; // @[Modules.scala 160:64:@34880.4]
  wire [13:0] buffer_10_431; // @[Modules.scala 160:64:@34881.4]
  wire [13:0] buffer_10_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87599; // @[Modules.scala 160:64:@34887.4]
  wire [13:0] _T_87600; // @[Modules.scala 160:64:@34888.4]
  wire [13:0] buffer_10_433; // @[Modules.scala 160:64:@34889.4]
  wire [13:0] buffer_10_252; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87602; // @[Modules.scala 160:64:@34891.4]
  wire [13:0] _T_87603; // @[Modules.scala 160:64:@34892.4]
  wire [13:0] buffer_10_434; // @[Modules.scala 160:64:@34893.4]
  wire [13:0] buffer_10_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87605; // @[Modules.scala 160:64:@34895.4]
  wire [13:0] _T_87606; // @[Modules.scala 160:64:@34896.4]
  wire [13:0] buffer_10_435; // @[Modules.scala 160:64:@34897.4]
  wire [13:0] buffer_10_256; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87608; // @[Modules.scala 160:64:@34899.4]
  wire [13:0] _T_87609; // @[Modules.scala 160:64:@34900.4]
  wire [13:0] buffer_10_436; // @[Modules.scala 160:64:@34901.4]
  wire [13:0] buffer_10_258; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87611; // @[Modules.scala 160:64:@34903.4]
  wire [13:0] _T_87612; // @[Modules.scala 160:64:@34904.4]
  wire [13:0] buffer_10_437; // @[Modules.scala 160:64:@34905.4]
  wire [13:0] buffer_10_262; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87617; // @[Modules.scala 160:64:@34911.4]
  wire [13:0] _T_87618; // @[Modules.scala 160:64:@34912.4]
  wire [13:0] buffer_10_439; // @[Modules.scala 160:64:@34913.4]
  wire [14:0] _T_87620; // @[Modules.scala 160:64:@34915.4]
  wire [13:0] _T_87621; // @[Modules.scala 160:64:@34916.4]
  wire [13:0] buffer_10_440; // @[Modules.scala 160:64:@34917.4]
  wire [13:0] buffer_10_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87629; // @[Modules.scala 160:64:@34927.4]
  wire [13:0] _T_87630; // @[Modules.scala 160:64:@34928.4]
  wire [13:0] buffer_10_443; // @[Modules.scala 160:64:@34929.4]
  wire [13:0] buffer_10_272; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87632; // @[Modules.scala 160:64:@34931.4]
  wire [13:0] _T_87633; // @[Modules.scala 160:64:@34932.4]
  wire [13:0] buffer_10_444; // @[Modules.scala 160:64:@34933.4]
  wire [14:0] _T_87635; // @[Modules.scala 160:64:@34935.4]
  wire [13:0] _T_87636; // @[Modules.scala 160:64:@34936.4]
  wire [13:0] buffer_10_445; // @[Modules.scala 160:64:@34937.4]
  wire [13:0] buffer_10_276; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_277; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87638; // @[Modules.scala 160:64:@34939.4]
  wire [13:0] _T_87639; // @[Modules.scala 160:64:@34940.4]
  wire [13:0] buffer_10_446; // @[Modules.scala 160:64:@34941.4]
  wire [13:0] buffer_10_278; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87641; // @[Modules.scala 160:64:@34943.4]
  wire [13:0] _T_87642; // @[Modules.scala 160:64:@34944.4]
  wire [13:0] buffer_10_447; // @[Modules.scala 160:64:@34945.4]
  wire [14:0] _T_87644; // @[Modules.scala 160:64:@34947.4]
  wire [13:0] _T_87645; // @[Modules.scala 160:64:@34948.4]
  wire [13:0] buffer_10_448; // @[Modules.scala 160:64:@34949.4]
  wire [13:0] buffer_10_287; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87653; // @[Modules.scala 160:64:@34959.4]
  wire [13:0] _T_87654; // @[Modules.scala 160:64:@34960.4]
  wire [13:0] buffer_10_451; // @[Modules.scala 160:64:@34961.4]
  wire [14:0] _T_87656; // @[Modules.scala 160:64:@34963.4]
  wire [13:0] _T_87657; // @[Modules.scala 160:64:@34964.4]
  wire [13:0] buffer_10_452; // @[Modules.scala 160:64:@34965.4]
  wire [13:0] buffer_10_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87659; // @[Modules.scala 160:64:@34967.4]
  wire [13:0] _T_87660; // @[Modules.scala 160:64:@34968.4]
  wire [13:0] buffer_10_453; // @[Modules.scala 160:64:@34969.4]
  wire [13:0] buffer_10_292; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87662; // @[Modules.scala 160:64:@34971.4]
  wire [13:0] _T_87663; // @[Modules.scala 160:64:@34972.4]
  wire [13:0] buffer_10_454; // @[Modules.scala 160:64:@34973.4]
  wire [14:0] _T_87665; // @[Modules.scala 160:64:@34975.4]
  wire [13:0] _T_87666; // @[Modules.scala 160:64:@34976.4]
  wire [13:0] buffer_10_455; // @[Modules.scala 160:64:@34977.4]
  wire [14:0] _T_87668; // @[Modules.scala 160:64:@34979.4]
  wire [13:0] _T_87669; // @[Modules.scala 160:64:@34980.4]
  wire [13:0] buffer_10_456; // @[Modules.scala 160:64:@34981.4]
  wire [13:0] buffer_10_298; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_10_299; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87671; // @[Modules.scala 160:64:@34983.4]
  wire [13:0] _T_87672; // @[Modules.scala 160:64:@34984.4]
  wire [13:0] buffer_10_457; // @[Modules.scala 160:64:@34985.4]
  wire [13:0] buffer_10_300; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_87674; // @[Modules.scala 160:64:@34987.4]
  wire [13:0] _T_87675; // @[Modules.scala 160:64:@34988.4]
  wire [13:0] buffer_10_458; // @[Modules.scala 160:64:@34989.4]
  wire [14:0] _T_87677; // @[Modules.scala 160:64:@34991.4]
  wire [13:0] _T_87678; // @[Modules.scala 160:64:@34992.4]
  wire [13:0] buffer_10_459; // @[Modules.scala 160:64:@34993.4]
  wire [14:0] _T_87686; // @[Modules.scala 160:64:@35003.4]
  wire [13:0] _T_87687; // @[Modules.scala 160:64:@35004.4]
  wire [13:0] buffer_10_462; // @[Modules.scala 160:64:@35005.4]
  wire [14:0] _T_87689; // @[Modules.scala 160:64:@35007.4]
  wire [13:0] _T_87690; // @[Modules.scala 160:64:@35008.4]
  wire [13:0] buffer_10_463; // @[Modules.scala 160:64:@35009.4]
  wire [14:0] _T_87692; // @[Modules.scala 160:64:@35011.4]
  wire [13:0] _T_87693; // @[Modules.scala 160:64:@35012.4]
  wire [13:0] buffer_10_464; // @[Modules.scala 160:64:@35013.4]
  wire [14:0] _T_87701; // @[Modules.scala 160:64:@35023.4]
  wire [13:0] _T_87702; // @[Modules.scala 160:64:@35024.4]
  wire [13:0] buffer_10_467; // @[Modules.scala 160:64:@35025.4]
  wire [14:0] _T_87704; // @[Modules.scala 160:64:@35027.4]
  wire [13:0] _T_87705; // @[Modules.scala 160:64:@35028.4]
  wire [13:0] buffer_10_468; // @[Modules.scala 160:64:@35029.4]
  wire [14:0] _T_87707; // @[Modules.scala 160:64:@35031.4]
  wire [13:0] _T_87708; // @[Modules.scala 160:64:@35032.4]
  wire [13:0] buffer_10_469; // @[Modules.scala 160:64:@35033.4]
  wire [14:0] _T_87710; // @[Modules.scala 160:64:@35035.4]
  wire [13:0] _T_87711; // @[Modules.scala 160:64:@35036.4]
  wire [13:0] buffer_10_470; // @[Modules.scala 160:64:@35037.4]
  wire [14:0] _T_87713; // @[Modules.scala 160:64:@35039.4]
  wire [13:0] _T_87714; // @[Modules.scala 160:64:@35040.4]
  wire [13:0] buffer_10_471; // @[Modules.scala 160:64:@35041.4]
  wire [14:0] _T_87716; // @[Modules.scala 160:64:@35043.4]
  wire [13:0] _T_87717; // @[Modules.scala 160:64:@35044.4]
  wire [13:0] buffer_10_472; // @[Modules.scala 160:64:@35045.4]
  wire [14:0] _T_87719; // @[Modules.scala 160:64:@35047.4]
  wire [13:0] _T_87720; // @[Modules.scala 160:64:@35048.4]
  wire [13:0] buffer_10_473; // @[Modules.scala 160:64:@35049.4]
  wire [14:0] _T_87722; // @[Modules.scala 160:64:@35051.4]
  wire [13:0] _T_87723; // @[Modules.scala 160:64:@35052.4]
  wire [13:0] buffer_10_474; // @[Modules.scala 160:64:@35053.4]
  wire [14:0] _T_87728; // @[Modules.scala 160:64:@35059.4]
  wire [13:0] _T_87729; // @[Modules.scala 160:64:@35060.4]
  wire [13:0] buffer_10_476; // @[Modules.scala 160:64:@35061.4]
  wire [14:0] _T_87731; // @[Modules.scala 160:64:@35063.4]
  wire [13:0] _T_87732; // @[Modules.scala 160:64:@35064.4]
  wire [13:0] buffer_10_477; // @[Modules.scala 160:64:@35065.4]
  wire [14:0] _T_87734; // @[Modules.scala 160:64:@35067.4]
  wire [13:0] _T_87735; // @[Modules.scala 160:64:@35068.4]
  wire [13:0] buffer_10_478; // @[Modules.scala 160:64:@35069.4]
  wire [14:0] _T_87737; // @[Modules.scala 160:64:@35071.4]
  wire [13:0] _T_87738; // @[Modules.scala 160:64:@35072.4]
  wire [13:0] buffer_10_479; // @[Modules.scala 160:64:@35073.4]
  wire [14:0] _T_87740; // @[Modules.scala 160:64:@35075.4]
  wire [13:0] _T_87741; // @[Modules.scala 160:64:@35076.4]
  wire [13:0] buffer_10_480; // @[Modules.scala 160:64:@35077.4]
  wire [14:0] _T_87743; // @[Modules.scala 160:64:@35079.4]
  wire [13:0] _T_87744; // @[Modules.scala 160:64:@35080.4]
  wire [13:0] buffer_10_481; // @[Modules.scala 160:64:@35081.4]
  wire [14:0] _T_87746; // @[Modules.scala 160:64:@35083.4]
  wire [13:0] _T_87747; // @[Modules.scala 160:64:@35084.4]
  wire [13:0] buffer_10_482; // @[Modules.scala 160:64:@35085.4]
  wire [14:0] _T_87749; // @[Modules.scala 160:64:@35087.4]
  wire [13:0] _T_87750; // @[Modules.scala 160:64:@35088.4]
  wire [13:0] buffer_10_483; // @[Modules.scala 160:64:@35089.4]
  wire [14:0] _T_87752; // @[Modules.scala 160:64:@35091.4]
  wire [13:0] _T_87753; // @[Modules.scala 160:64:@35092.4]
  wire [13:0] buffer_10_484; // @[Modules.scala 160:64:@35093.4]
  wire [14:0] _T_87755; // @[Modules.scala 160:64:@35095.4]
  wire [13:0] _T_87756; // @[Modules.scala 160:64:@35096.4]
  wire [13:0] buffer_10_485; // @[Modules.scala 160:64:@35097.4]
  wire [14:0] _T_87758; // @[Modules.scala 160:64:@35099.4]
  wire [13:0] _T_87759; // @[Modules.scala 160:64:@35100.4]
  wire [13:0] buffer_10_486; // @[Modules.scala 160:64:@35101.4]
  wire [14:0] _T_87761; // @[Modules.scala 160:64:@35103.4]
  wire [13:0] _T_87762; // @[Modules.scala 160:64:@35104.4]
  wire [13:0] buffer_10_487; // @[Modules.scala 160:64:@35105.4]
  wire [14:0] _T_87764; // @[Modules.scala 160:64:@35107.4]
  wire [13:0] _T_87765; // @[Modules.scala 160:64:@35108.4]
  wire [13:0] buffer_10_488; // @[Modules.scala 160:64:@35109.4]
  wire [14:0] _T_87767; // @[Modules.scala 160:64:@35111.4]
  wire [13:0] _T_87768; // @[Modules.scala 160:64:@35112.4]
  wire [13:0] buffer_10_489; // @[Modules.scala 160:64:@35113.4]
  wire [14:0] _T_87770; // @[Modules.scala 160:64:@35115.4]
  wire [13:0] _T_87771; // @[Modules.scala 160:64:@35116.4]
  wire [13:0] buffer_10_490; // @[Modules.scala 160:64:@35117.4]
  wire [14:0] _T_87773; // @[Modules.scala 160:64:@35119.4]
  wire [13:0] _T_87774; // @[Modules.scala 160:64:@35120.4]
  wire [13:0] buffer_10_491; // @[Modules.scala 160:64:@35121.4]
  wire [14:0] _T_87776; // @[Modules.scala 160:64:@35123.4]
  wire [13:0] _T_87777; // @[Modules.scala 160:64:@35124.4]
  wire [13:0] buffer_10_492; // @[Modules.scala 160:64:@35125.4]
  wire [14:0] _T_87779; // @[Modules.scala 160:64:@35127.4]
  wire [13:0] _T_87780; // @[Modules.scala 160:64:@35128.4]
  wire [13:0] buffer_10_493; // @[Modules.scala 160:64:@35129.4]
  wire [14:0] _T_87782; // @[Modules.scala 160:64:@35131.4]
  wire [13:0] _T_87783; // @[Modules.scala 160:64:@35132.4]
  wire [13:0] buffer_10_494; // @[Modules.scala 160:64:@35133.4]
  wire [14:0] _T_87785; // @[Modules.scala 160:64:@35135.4]
  wire [13:0] _T_87786; // @[Modules.scala 160:64:@35136.4]
  wire [13:0] buffer_10_495; // @[Modules.scala 160:64:@35137.4]
  wire [14:0] _T_87788; // @[Modules.scala 160:64:@35139.4]
  wire [13:0] _T_87789; // @[Modules.scala 160:64:@35140.4]
  wire [13:0] buffer_10_496; // @[Modules.scala 160:64:@35141.4]
  wire [14:0] _T_87791; // @[Modules.scala 160:64:@35143.4]
  wire [13:0] _T_87792; // @[Modules.scala 160:64:@35144.4]
  wire [13:0] buffer_10_497; // @[Modules.scala 160:64:@35145.4]
  wire [14:0] _T_87794; // @[Modules.scala 160:64:@35147.4]
  wire [13:0] _T_87795; // @[Modules.scala 160:64:@35148.4]
  wire [13:0] buffer_10_498; // @[Modules.scala 160:64:@35149.4]
  wire [14:0] _T_87797; // @[Modules.scala 160:64:@35151.4]
  wire [13:0] _T_87798; // @[Modules.scala 160:64:@35152.4]
  wire [13:0] buffer_10_499; // @[Modules.scala 160:64:@35153.4]
  wire [14:0] _T_87800; // @[Modules.scala 160:64:@35155.4]
  wire [13:0] _T_87801; // @[Modules.scala 160:64:@35156.4]
  wire [13:0] buffer_10_500; // @[Modules.scala 160:64:@35157.4]
  wire [14:0] _T_87803; // @[Modules.scala 160:64:@35159.4]
  wire [13:0] _T_87804; // @[Modules.scala 160:64:@35160.4]
  wire [13:0] buffer_10_501; // @[Modules.scala 160:64:@35161.4]
  wire [14:0] _T_87806; // @[Modules.scala 160:64:@35163.4]
  wire [13:0] _T_87807; // @[Modules.scala 160:64:@35164.4]
  wire [13:0] buffer_10_502; // @[Modules.scala 160:64:@35165.4]
  wire [14:0] _T_87809; // @[Modules.scala 160:64:@35167.4]
  wire [13:0] _T_87810; // @[Modules.scala 160:64:@35168.4]
  wire [13:0] buffer_10_503; // @[Modules.scala 160:64:@35169.4]
  wire [14:0] _T_87812; // @[Modules.scala 160:64:@35171.4]
  wire [13:0] _T_87813; // @[Modules.scala 160:64:@35172.4]
  wire [13:0] buffer_10_504; // @[Modules.scala 160:64:@35173.4]
  wire [14:0] _T_87815; // @[Modules.scala 160:64:@35175.4]
  wire [13:0] _T_87816; // @[Modules.scala 160:64:@35176.4]
  wire [13:0] buffer_10_505; // @[Modules.scala 160:64:@35177.4]
  wire [14:0] _T_87818; // @[Modules.scala 160:64:@35179.4]
  wire [13:0] _T_87819; // @[Modules.scala 160:64:@35180.4]
  wire [13:0] buffer_10_506; // @[Modules.scala 160:64:@35181.4]
  wire [14:0] _T_87821; // @[Modules.scala 160:64:@35183.4]
  wire [13:0] _T_87822; // @[Modules.scala 160:64:@35184.4]
  wire [13:0] buffer_10_507; // @[Modules.scala 160:64:@35185.4]
  wire [14:0] _T_87824; // @[Modules.scala 160:64:@35187.4]
  wire [13:0] _T_87825; // @[Modules.scala 160:64:@35188.4]
  wire [13:0] buffer_10_508; // @[Modules.scala 160:64:@35189.4]
  wire [14:0] _T_87827; // @[Modules.scala 160:64:@35191.4]
  wire [13:0] _T_87828; // @[Modules.scala 160:64:@35192.4]
  wire [13:0] buffer_10_509; // @[Modules.scala 160:64:@35193.4]
  wire [14:0] _T_87830; // @[Modules.scala 160:64:@35195.4]
  wire [13:0] _T_87831; // @[Modules.scala 160:64:@35196.4]
  wire [13:0] buffer_10_510; // @[Modules.scala 160:64:@35197.4]
  wire [14:0] _T_87833; // @[Modules.scala 160:64:@35199.4]
  wire [13:0] _T_87834; // @[Modules.scala 160:64:@35200.4]
  wire [13:0] buffer_10_511; // @[Modules.scala 160:64:@35201.4]
  wire [14:0] _T_87836; // @[Modules.scala 160:64:@35203.4]
  wire [13:0] _T_87837; // @[Modules.scala 160:64:@35204.4]
  wire [13:0] buffer_10_512; // @[Modules.scala 160:64:@35205.4]
  wire [14:0] _T_87839; // @[Modules.scala 160:64:@35207.4]
  wire [13:0] _T_87840; // @[Modules.scala 160:64:@35208.4]
  wire [13:0] buffer_10_513; // @[Modules.scala 160:64:@35209.4]
  wire [14:0] _T_87842; // @[Modules.scala 160:64:@35211.4]
  wire [13:0] _T_87843; // @[Modules.scala 160:64:@35212.4]
  wire [13:0] buffer_10_514; // @[Modules.scala 160:64:@35213.4]
  wire [14:0] _T_87845; // @[Modules.scala 160:64:@35215.4]
  wire [13:0] _T_87846; // @[Modules.scala 160:64:@35216.4]
  wire [13:0] buffer_10_515; // @[Modules.scala 160:64:@35217.4]
  wire [14:0] _T_87848; // @[Modules.scala 160:64:@35219.4]
  wire [13:0] _T_87849; // @[Modules.scala 160:64:@35220.4]
  wire [13:0] buffer_10_516; // @[Modules.scala 160:64:@35221.4]
  wire [14:0] _T_87851; // @[Modules.scala 160:64:@35223.4]
  wire [13:0] _T_87852; // @[Modules.scala 160:64:@35224.4]
  wire [13:0] buffer_10_517; // @[Modules.scala 160:64:@35225.4]
  wire [14:0] _T_87854; // @[Modules.scala 160:64:@35227.4]
  wire [13:0] _T_87855; // @[Modules.scala 160:64:@35228.4]
  wire [13:0] buffer_10_518; // @[Modules.scala 160:64:@35229.4]
  wire [14:0] _T_87857; // @[Modules.scala 160:64:@35231.4]
  wire [13:0] _T_87858; // @[Modules.scala 160:64:@35232.4]
  wire [13:0] buffer_10_519; // @[Modules.scala 160:64:@35233.4]
  wire [14:0] _T_87860; // @[Modules.scala 160:64:@35235.4]
  wire [13:0] _T_87861; // @[Modules.scala 160:64:@35236.4]
  wire [13:0] buffer_10_520; // @[Modules.scala 160:64:@35237.4]
  wire [14:0] _T_87863; // @[Modules.scala 160:64:@35239.4]
  wire [13:0] _T_87864; // @[Modules.scala 160:64:@35240.4]
  wire [13:0] buffer_10_521; // @[Modules.scala 160:64:@35241.4]
  wire [14:0] _T_87866; // @[Modules.scala 160:64:@35243.4]
  wire [13:0] _T_87867; // @[Modules.scala 160:64:@35244.4]
  wire [13:0] buffer_10_522; // @[Modules.scala 160:64:@35245.4]
  wire [14:0] _T_87869; // @[Modules.scala 160:64:@35247.4]
  wire [13:0] _T_87870; // @[Modules.scala 160:64:@35248.4]
  wire [13:0] buffer_10_523; // @[Modules.scala 160:64:@35249.4]
  wire [14:0] _T_87872; // @[Modules.scala 160:64:@35251.4]
  wire [13:0] _T_87873; // @[Modules.scala 160:64:@35252.4]
  wire [13:0] buffer_10_524; // @[Modules.scala 160:64:@35253.4]
  wire [14:0] _T_87875; // @[Modules.scala 160:64:@35255.4]
  wire [13:0] _T_87876; // @[Modules.scala 160:64:@35256.4]
  wire [13:0] buffer_10_525; // @[Modules.scala 160:64:@35257.4]
  wire [14:0] _T_87878; // @[Modules.scala 160:64:@35259.4]
  wire [13:0] _T_87879; // @[Modules.scala 160:64:@35260.4]
  wire [13:0] buffer_10_526; // @[Modules.scala 160:64:@35261.4]
  wire [14:0] _T_87881; // @[Modules.scala 160:64:@35263.4]
  wire [13:0] _T_87882; // @[Modules.scala 160:64:@35264.4]
  wire [13:0] buffer_10_527; // @[Modules.scala 160:64:@35265.4]
  wire [14:0] _T_87884; // @[Modules.scala 160:64:@35267.4]
  wire [13:0] _T_87885; // @[Modules.scala 160:64:@35268.4]
  wire [13:0] buffer_10_528; // @[Modules.scala 160:64:@35269.4]
  wire [14:0] _T_87887; // @[Modules.scala 160:64:@35271.4]
  wire [13:0] _T_87888; // @[Modules.scala 160:64:@35272.4]
  wire [13:0] buffer_10_529; // @[Modules.scala 160:64:@35273.4]
  wire [14:0] _T_87890; // @[Modules.scala 160:64:@35275.4]
  wire [13:0] _T_87891; // @[Modules.scala 160:64:@35276.4]
  wire [13:0] buffer_10_530; // @[Modules.scala 160:64:@35277.4]
  wire [14:0] _T_87893; // @[Modules.scala 160:64:@35279.4]
  wire [13:0] _T_87894; // @[Modules.scala 160:64:@35280.4]
  wire [13:0] buffer_10_531; // @[Modules.scala 160:64:@35281.4]
  wire [14:0] _T_87896; // @[Modules.scala 160:64:@35283.4]
  wire [13:0] _T_87897; // @[Modules.scala 160:64:@35284.4]
  wire [13:0] buffer_10_532; // @[Modules.scala 160:64:@35285.4]
  wire [14:0] _T_87899; // @[Modules.scala 160:64:@35287.4]
  wire [13:0] _T_87900; // @[Modules.scala 160:64:@35288.4]
  wire [13:0] buffer_10_533; // @[Modules.scala 160:64:@35289.4]
  wire [14:0] _T_87902; // @[Modules.scala 160:64:@35291.4]
  wire [13:0] _T_87903; // @[Modules.scala 160:64:@35292.4]
  wire [13:0] buffer_10_534; // @[Modules.scala 160:64:@35293.4]
  wire [14:0] _T_87905; // @[Modules.scala 160:64:@35295.4]
  wire [13:0] _T_87906; // @[Modules.scala 160:64:@35296.4]
  wire [13:0] buffer_10_535; // @[Modules.scala 160:64:@35297.4]
  wire [14:0] _T_87908; // @[Modules.scala 160:64:@35299.4]
  wire [13:0] _T_87909; // @[Modules.scala 160:64:@35300.4]
  wire [13:0] buffer_10_536; // @[Modules.scala 160:64:@35301.4]
  wire [14:0] _T_87911; // @[Modules.scala 160:64:@35303.4]
  wire [13:0] _T_87912; // @[Modules.scala 160:64:@35304.4]
  wire [13:0] buffer_10_537; // @[Modules.scala 160:64:@35305.4]
  wire [14:0] _T_87917; // @[Modules.scala 166:64:@35311.4]
  wire [13:0] _T_87918; // @[Modules.scala 166:64:@35312.4]
  wire [13:0] buffer_10_539; // @[Modules.scala 166:64:@35313.4]
  wire [14:0] _T_87920; // @[Modules.scala 166:64:@35315.4]
  wire [13:0] _T_87921; // @[Modules.scala 166:64:@35316.4]
  wire [13:0] buffer_10_540; // @[Modules.scala 166:64:@35317.4]
  wire [14:0] _T_87923; // @[Modules.scala 166:64:@35319.4]
  wire [13:0] _T_87924; // @[Modules.scala 166:64:@35320.4]
  wire [13:0] buffer_10_541; // @[Modules.scala 166:64:@35321.4]
  wire [14:0] _T_87926; // @[Modules.scala 166:64:@35323.4]
  wire [13:0] _T_87927; // @[Modules.scala 166:64:@35324.4]
  wire [13:0] buffer_10_542; // @[Modules.scala 166:64:@35325.4]
  wire [14:0] _T_87929; // @[Modules.scala 166:64:@35327.4]
  wire [13:0] _T_87930; // @[Modules.scala 166:64:@35328.4]
  wire [13:0] buffer_10_543; // @[Modules.scala 166:64:@35329.4]
  wire [14:0] _T_87932; // @[Modules.scala 166:64:@35331.4]
  wire [13:0] _T_87933; // @[Modules.scala 166:64:@35332.4]
  wire [13:0] buffer_10_544; // @[Modules.scala 166:64:@35333.4]
  wire [14:0] _T_87935; // @[Modules.scala 166:64:@35335.4]
  wire [13:0] _T_87936; // @[Modules.scala 166:64:@35336.4]
  wire [13:0] buffer_10_545; // @[Modules.scala 166:64:@35337.4]
  wire [14:0] _T_87938; // @[Modules.scala 166:64:@35339.4]
  wire [13:0] _T_87939; // @[Modules.scala 166:64:@35340.4]
  wire [13:0] buffer_10_546; // @[Modules.scala 166:64:@35341.4]
  wire [14:0] _T_87941; // @[Modules.scala 166:64:@35343.4]
  wire [13:0] _T_87942; // @[Modules.scala 166:64:@35344.4]
  wire [13:0] buffer_10_547; // @[Modules.scala 166:64:@35345.4]
  wire [14:0] _T_87944; // @[Modules.scala 166:64:@35347.4]
  wire [13:0] _T_87945; // @[Modules.scala 166:64:@35348.4]
  wire [13:0] buffer_10_548; // @[Modules.scala 166:64:@35349.4]
  wire [14:0] _T_87947; // @[Modules.scala 166:64:@35351.4]
  wire [13:0] _T_87948; // @[Modules.scala 166:64:@35352.4]
  wire [13:0] buffer_10_549; // @[Modules.scala 166:64:@35353.4]
  wire [14:0] _T_87950; // @[Modules.scala 166:64:@35355.4]
  wire [13:0] _T_87951; // @[Modules.scala 166:64:@35356.4]
  wire [13:0] buffer_10_550; // @[Modules.scala 166:64:@35357.4]
  wire [14:0] _T_87953; // @[Modules.scala 166:64:@35359.4]
  wire [13:0] _T_87954; // @[Modules.scala 166:64:@35360.4]
  wire [13:0] buffer_10_551; // @[Modules.scala 166:64:@35361.4]
  wire [14:0] _T_87956; // @[Modules.scala 166:64:@35363.4]
  wire [13:0] _T_87957; // @[Modules.scala 166:64:@35364.4]
  wire [13:0] buffer_10_552; // @[Modules.scala 166:64:@35365.4]
  wire [14:0] _T_87959; // @[Modules.scala 166:64:@35367.4]
  wire [13:0] _T_87960; // @[Modules.scala 166:64:@35368.4]
  wire [13:0] buffer_10_553; // @[Modules.scala 166:64:@35369.4]
  wire [14:0] _T_87962; // @[Modules.scala 166:64:@35371.4]
  wire [13:0] _T_87963; // @[Modules.scala 166:64:@35372.4]
  wire [13:0] buffer_10_554; // @[Modules.scala 166:64:@35373.4]
  wire [14:0] _T_87965; // @[Modules.scala 166:64:@35375.4]
  wire [13:0] _T_87966; // @[Modules.scala 166:64:@35376.4]
  wire [13:0] buffer_10_555; // @[Modules.scala 166:64:@35377.4]
  wire [14:0] _T_87968; // @[Modules.scala 166:64:@35379.4]
  wire [13:0] _T_87969; // @[Modules.scala 166:64:@35380.4]
  wire [13:0] buffer_10_556; // @[Modules.scala 166:64:@35381.4]
  wire [14:0] _T_87971; // @[Modules.scala 166:64:@35383.4]
  wire [13:0] _T_87972; // @[Modules.scala 166:64:@35384.4]
  wire [13:0] buffer_10_557; // @[Modules.scala 166:64:@35385.4]
  wire [14:0] _T_87974; // @[Modules.scala 166:64:@35387.4]
  wire [13:0] _T_87975; // @[Modules.scala 166:64:@35388.4]
  wire [13:0] buffer_10_558; // @[Modules.scala 166:64:@35389.4]
  wire [14:0] _T_87977; // @[Modules.scala 166:64:@35391.4]
  wire [13:0] _T_87978; // @[Modules.scala 166:64:@35392.4]
  wire [13:0] buffer_10_559; // @[Modules.scala 166:64:@35393.4]
  wire [14:0] _T_87980; // @[Modules.scala 166:64:@35395.4]
  wire [13:0] _T_87981; // @[Modules.scala 166:64:@35396.4]
  wire [13:0] buffer_10_560; // @[Modules.scala 166:64:@35397.4]
  wire [14:0] _T_87983; // @[Modules.scala 166:64:@35399.4]
  wire [13:0] _T_87984; // @[Modules.scala 166:64:@35400.4]
  wire [13:0] buffer_10_561; // @[Modules.scala 166:64:@35401.4]
  wire [14:0] _T_87986; // @[Modules.scala 166:64:@35403.4]
  wire [13:0] _T_87987; // @[Modules.scala 166:64:@35404.4]
  wire [13:0] buffer_10_562; // @[Modules.scala 166:64:@35405.4]
  wire [14:0] _T_87989; // @[Modules.scala 166:64:@35407.4]
  wire [13:0] _T_87990; // @[Modules.scala 166:64:@35408.4]
  wire [13:0] buffer_10_563; // @[Modules.scala 166:64:@35409.4]
  wire [14:0] _T_87992; // @[Modules.scala 166:64:@35411.4]
  wire [13:0] _T_87993; // @[Modules.scala 166:64:@35412.4]
  wire [13:0] buffer_10_564; // @[Modules.scala 166:64:@35413.4]
  wire [14:0] _T_87995; // @[Modules.scala 166:64:@35415.4]
  wire [13:0] _T_87996; // @[Modules.scala 166:64:@35416.4]
  wire [13:0] buffer_10_565; // @[Modules.scala 166:64:@35417.4]
  wire [14:0] _T_87998; // @[Modules.scala 166:64:@35419.4]
  wire [13:0] _T_87999; // @[Modules.scala 166:64:@35420.4]
  wire [13:0] buffer_10_566; // @[Modules.scala 166:64:@35421.4]
  wire [14:0] _T_88001; // @[Modules.scala 166:64:@35423.4]
  wire [13:0] _T_88002; // @[Modules.scala 166:64:@35424.4]
  wire [13:0] buffer_10_567; // @[Modules.scala 166:64:@35425.4]
  wire [14:0] _T_88004; // @[Modules.scala 166:64:@35427.4]
  wire [13:0] _T_88005; // @[Modules.scala 166:64:@35428.4]
  wire [13:0] buffer_10_568; // @[Modules.scala 166:64:@35429.4]
  wire [14:0] _T_88007; // @[Modules.scala 166:64:@35431.4]
  wire [13:0] _T_88008; // @[Modules.scala 166:64:@35432.4]
  wire [13:0] buffer_10_569; // @[Modules.scala 166:64:@35433.4]
  wire [14:0] _T_88010; // @[Modules.scala 166:64:@35435.4]
  wire [13:0] _T_88011; // @[Modules.scala 166:64:@35436.4]
  wire [13:0] buffer_10_570; // @[Modules.scala 166:64:@35437.4]
  wire [14:0] _T_88013; // @[Modules.scala 166:64:@35439.4]
  wire [13:0] _T_88014; // @[Modules.scala 166:64:@35440.4]
  wire [13:0] buffer_10_571; // @[Modules.scala 166:64:@35441.4]
  wire [14:0] _T_88016; // @[Modules.scala 166:64:@35443.4]
  wire [13:0] _T_88017; // @[Modules.scala 166:64:@35444.4]
  wire [13:0] buffer_10_572; // @[Modules.scala 166:64:@35445.4]
  wire [14:0] _T_88019; // @[Modules.scala 166:64:@35447.4]
  wire [13:0] _T_88020; // @[Modules.scala 166:64:@35448.4]
  wire [13:0] buffer_10_573; // @[Modules.scala 166:64:@35449.4]
  wire [14:0] _T_88022; // @[Modules.scala 166:64:@35451.4]
  wire [13:0] _T_88023; // @[Modules.scala 166:64:@35452.4]
  wire [13:0] buffer_10_574; // @[Modules.scala 166:64:@35453.4]
  wire [14:0] _T_88025; // @[Modules.scala 166:64:@35455.4]
  wire [13:0] _T_88026; // @[Modules.scala 166:64:@35456.4]
  wire [13:0] buffer_10_575; // @[Modules.scala 166:64:@35457.4]
  wire [14:0] _T_88028; // @[Modules.scala 166:64:@35459.4]
  wire [13:0] _T_88029; // @[Modules.scala 166:64:@35460.4]
  wire [13:0] buffer_10_576; // @[Modules.scala 166:64:@35461.4]
  wire [14:0] _T_88031; // @[Modules.scala 160:64:@35463.4]
  wire [13:0] _T_88032; // @[Modules.scala 160:64:@35464.4]
  wire [13:0] buffer_10_577; // @[Modules.scala 160:64:@35465.4]
  wire [14:0] _T_88034; // @[Modules.scala 160:64:@35467.4]
  wire [13:0] _T_88035; // @[Modules.scala 160:64:@35468.4]
  wire [13:0] buffer_10_578; // @[Modules.scala 160:64:@35469.4]
  wire [14:0] _T_88037; // @[Modules.scala 160:64:@35471.4]
  wire [13:0] _T_88038; // @[Modules.scala 160:64:@35472.4]
  wire [13:0] buffer_10_579; // @[Modules.scala 160:64:@35473.4]
  wire [14:0] _T_88040; // @[Modules.scala 160:64:@35475.4]
  wire [13:0] _T_88041; // @[Modules.scala 160:64:@35476.4]
  wire [13:0] buffer_10_580; // @[Modules.scala 160:64:@35477.4]
  wire [14:0] _T_88043; // @[Modules.scala 160:64:@35479.4]
  wire [13:0] _T_88044; // @[Modules.scala 160:64:@35480.4]
  wire [13:0] buffer_10_581; // @[Modules.scala 160:64:@35481.4]
  wire [14:0] _T_88046; // @[Modules.scala 160:64:@35483.4]
  wire [13:0] _T_88047; // @[Modules.scala 160:64:@35484.4]
  wire [13:0] buffer_10_582; // @[Modules.scala 160:64:@35485.4]
  wire [14:0] _T_88049; // @[Modules.scala 160:64:@35487.4]
  wire [13:0] _T_88050; // @[Modules.scala 160:64:@35488.4]
  wire [13:0] buffer_10_583; // @[Modules.scala 160:64:@35489.4]
  wire [14:0] _T_88052; // @[Modules.scala 160:64:@35491.4]
  wire [13:0] _T_88053; // @[Modules.scala 160:64:@35492.4]
  wire [13:0] buffer_10_584; // @[Modules.scala 160:64:@35493.4]
  wire [14:0] _T_88055; // @[Modules.scala 160:64:@35495.4]
  wire [13:0] _T_88056; // @[Modules.scala 160:64:@35496.4]
  wire [13:0] buffer_10_585; // @[Modules.scala 160:64:@35497.4]
  wire [14:0] _T_88058; // @[Modules.scala 160:64:@35499.4]
  wire [13:0] _T_88059; // @[Modules.scala 160:64:@35500.4]
  wire [13:0] buffer_10_586; // @[Modules.scala 160:64:@35501.4]
  wire [14:0] _T_88061; // @[Modules.scala 160:64:@35503.4]
  wire [13:0] _T_88062; // @[Modules.scala 160:64:@35504.4]
  wire [13:0] buffer_10_587; // @[Modules.scala 160:64:@35505.4]
  wire [14:0] _T_88064; // @[Modules.scala 160:64:@35507.4]
  wire [13:0] _T_88065; // @[Modules.scala 160:64:@35508.4]
  wire [13:0] buffer_10_588; // @[Modules.scala 160:64:@35509.4]
  wire [14:0] _T_88067; // @[Modules.scala 160:64:@35511.4]
  wire [13:0] _T_88068; // @[Modules.scala 160:64:@35512.4]
  wire [13:0] buffer_10_589; // @[Modules.scala 160:64:@35513.4]
  wire [14:0] _T_88070; // @[Modules.scala 160:64:@35515.4]
  wire [13:0] _T_88071; // @[Modules.scala 160:64:@35516.4]
  wire [13:0] buffer_10_590; // @[Modules.scala 160:64:@35517.4]
  wire [14:0] _T_88073; // @[Modules.scala 160:64:@35519.4]
  wire [13:0] _T_88074; // @[Modules.scala 160:64:@35520.4]
  wire [13:0] buffer_10_591; // @[Modules.scala 160:64:@35521.4]
  wire [14:0] _T_88076; // @[Modules.scala 160:64:@35523.4]
  wire [13:0] _T_88077; // @[Modules.scala 160:64:@35524.4]
  wire [13:0] buffer_10_592; // @[Modules.scala 160:64:@35525.4]
  wire [14:0] _T_88079; // @[Modules.scala 160:64:@35527.4]
  wire [13:0] _T_88080; // @[Modules.scala 160:64:@35528.4]
  wire [13:0] buffer_10_593; // @[Modules.scala 160:64:@35529.4]
  wire [14:0] _T_88082; // @[Modules.scala 160:64:@35531.4]
  wire [13:0] _T_88083; // @[Modules.scala 160:64:@35532.4]
  wire [13:0] buffer_10_594; // @[Modules.scala 160:64:@35533.4]
  wire [14:0] _T_88085; // @[Modules.scala 160:64:@35535.4]
  wire [13:0] _T_88086; // @[Modules.scala 160:64:@35536.4]
  wire [13:0] buffer_10_595; // @[Modules.scala 160:64:@35537.4]
  wire [14:0] _T_88088; // @[Modules.scala 166:64:@35539.4]
  wire [13:0] _T_88089; // @[Modules.scala 166:64:@35540.4]
  wire [13:0] buffer_10_596; // @[Modules.scala 166:64:@35541.4]
  wire [14:0] _T_88091; // @[Modules.scala 166:64:@35543.4]
  wire [13:0] _T_88092; // @[Modules.scala 166:64:@35544.4]
  wire [13:0] buffer_10_597; // @[Modules.scala 166:64:@35545.4]
  wire [14:0] _T_88094; // @[Modules.scala 166:64:@35547.4]
  wire [13:0] _T_88095; // @[Modules.scala 166:64:@35548.4]
  wire [13:0] buffer_10_598; // @[Modules.scala 166:64:@35549.4]
  wire [14:0] _T_88097; // @[Modules.scala 166:64:@35551.4]
  wire [13:0] _T_88098; // @[Modules.scala 166:64:@35552.4]
  wire [13:0] buffer_10_599; // @[Modules.scala 166:64:@35553.4]
  wire [14:0] _T_88100; // @[Modules.scala 166:64:@35555.4]
  wire [13:0] _T_88101; // @[Modules.scala 166:64:@35556.4]
  wire [13:0] buffer_10_600; // @[Modules.scala 166:64:@35557.4]
  wire [14:0] _T_88103; // @[Modules.scala 166:64:@35559.4]
  wire [13:0] _T_88104; // @[Modules.scala 166:64:@35560.4]
  wire [13:0] buffer_10_601; // @[Modules.scala 166:64:@35561.4]
  wire [14:0] _T_88106; // @[Modules.scala 166:64:@35563.4]
  wire [13:0] _T_88107; // @[Modules.scala 166:64:@35564.4]
  wire [13:0] buffer_10_602; // @[Modules.scala 166:64:@35565.4]
  wire [14:0] _T_88109; // @[Modules.scala 166:64:@35567.4]
  wire [13:0] _T_88110; // @[Modules.scala 166:64:@35568.4]
  wire [13:0] buffer_10_603; // @[Modules.scala 166:64:@35569.4]
  wire [14:0] _T_88112; // @[Modules.scala 166:64:@35571.4]
  wire [13:0] _T_88113; // @[Modules.scala 166:64:@35572.4]
  wire [13:0] buffer_10_604; // @[Modules.scala 166:64:@35573.4]
  wire [14:0] _T_88115; // @[Modules.scala 172:66:@35575.4]
  wire [13:0] _T_88116; // @[Modules.scala 172:66:@35576.4]
  wire [13:0] buffer_10_605; // @[Modules.scala 172:66:@35577.4]
  wire [14:0] _T_88118; // @[Modules.scala 160:64:@35579.4]
  wire [13:0] _T_88119; // @[Modules.scala 160:64:@35580.4]
  wire [13:0] buffer_10_606; // @[Modules.scala 160:64:@35581.4]
  wire [14:0] _T_88121; // @[Modules.scala 160:64:@35583.4]
  wire [13:0] _T_88122; // @[Modules.scala 160:64:@35584.4]
  wire [13:0] buffer_10_607; // @[Modules.scala 160:64:@35585.4]
  wire [14:0] _T_88124; // @[Modules.scala 160:64:@35587.4]
  wire [13:0] _T_88125; // @[Modules.scala 160:64:@35588.4]
  wire [13:0] buffer_10_608; // @[Modules.scala 160:64:@35589.4]
  wire [14:0] _T_88127; // @[Modules.scala 160:64:@35591.4]
  wire [13:0] _T_88128; // @[Modules.scala 160:64:@35592.4]
  wire [13:0] buffer_10_609; // @[Modules.scala 160:64:@35593.4]
  wire [14:0] _T_88130; // @[Modules.scala 160:64:@35595.4]
  wire [13:0] _T_88131; // @[Modules.scala 160:64:@35596.4]
  wire [13:0] buffer_10_610; // @[Modules.scala 160:64:@35597.4]
  wire [14:0] _T_88133; // @[Modules.scala 166:64:@35599.4]
  wire [13:0] _T_88134; // @[Modules.scala 166:64:@35600.4]
  wire [13:0] buffer_10_611; // @[Modules.scala 166:64:@35601.4]
  wire [14:0] _T_88136; // @[Modules.scala 166:64:@35603.4]
  wire [13:0] _T_88137; // @[Modules.scala 166:64:@35604.4]
  wire [13:0] buffer_10_612; // @[Modules.scala 166:64:@35605.4]
  wire [14:0] _T_88139; // @[Modules.scala 160:64:@35607.4]
  wire [13:0] _T_88140; // @[Modules.scala 160:64:@35608.4]
  wire [13:0] buffer_10_613; // @[Modules.scala 160:64:@35609.4]
  wire [14:0] _T_88142; // @[Modules.scala 172:66:@35611.4]
  wire [13:0] _T_88143; // @[Modules.scala 172:66:@35612.4]
  wire [13:0] buffer_10_614; // @[Modules.scala 172:66:@35613.4]
  wire [5:0] _T_88146; // @[Modules.scala 150:74:@35784.4]
  wire [6:0] _T_88149; // @[Modules.scala 150:103:@35786.4]
  wire [5:0] _T_88150; // @[Modules.scala 150:103:@35787.4]
  wire [5:0] _T_88151; // @[Modules.scala 150:103:@35788.4]
  wire [6:0] _T_88156; // @[Modules.scala 150:103:@35792.4]
  wire [5:0] _T_88157; // @[Modules.scala 150:103:@35793.4]
  wire [5:0] _T_88158; // @[Modules.scala 150:103:@35794.4]
  wire [6:0] _T_88163; // @[Modules.scala 150:103:@35798.4]
  wire [5:0] _T_88164; // @[Modules.scala 150:103:@35799.4]
  wire [5:0] _T_88165; // @[Modules.scala 150:103:@35800.4]
  wire [6:0] _T_88170; // @[Modules.scala 150:103:@35804.4]
  wire [5:0] _T_88171; // @[Modules.scala 150:103:@35805.4]
  wire [5:0] _T_88172; // @[Modules.scala 150:103:@35806.4]
  wire [6:0] _T_88205; // @[Modules.scala 150:103:@35834.4]
  wire [5:0] _T_88206; // @[Modules.scala 150:103:@35835.4]
  wire [5:0] _T_88207; // @[Modules.scala 150:103:@35836.4]
  wire [6:0] _T_88226; // @[Modules.scala 150:103:@35852.4]
  wire [5:0] _T_88227; // @[Modules.scala 150:103:@35853.4]
  wire [5:0] _T_88228; // @[Modules.scala 150:103:@35854.4]
  wire [5:0] _T_88302; // @[Modules.scala 151:80:@35917.4]
  wire [6:0] _T_88303; // @[Modules.scala 150:103:@35918.4]
  wire [5:0] _T_88304; // @[Modules.scala 150:103:@35919.4]
  wire [5:0] _T_88305; // @[Modules.scala 150:103:@35920.4]
  wire [6:0] _T_88387; // @[Modules.scala 150:103:@35990.4]
  wire [5:0] _T_88388; // @[Modules.scala 150:103:@35991.4]
  wire [5:0] _T_88389; // @[Modules.scala 150:103:@35992.4]
  wire [5:0] _GEN_766; // @[Modules.scala 150:103:@36038.4]
  wire [6:0] _T_88443; // @[Modules.scala 150:103:@36038.4]
  wire [5:0] _T_88444; // @[Modules.scala 150:103:@36039.4]
  wire [5:0] _T_88445; // @[Modules.scala 150:103:@36040.4]
  wire [6:0] _T_88457; // @[Modules.scala 150:103:@36050.4]
  wire [5:0] _T_88458; // @[Modules.scala 150:103:@36051.4]
  wire [5:0] _T_88459; // @[Modules.scala 150:103:@36052.4]
  wire [5:0] _T_88463; // @[Modules.scala 151:80:@36055.4]
  wire [6:0] _T_88464; // @[Modules.scala 150:103:@36056.4]
  wire [5:0] _T_88465; // @[Modules.scala 150:103:@36057.4]
  wire [5:0] _T_88466; // @[Modules.scala 150:103:@36058.4]
  wire [6:0] _T_88485; // @[Modules.scala 150:103:@36074.4]
  wire [5:0] _T_88486; // @[Modules.scala 150:103:@36075.4]
  wire [5:0] _T_88487; // @[Modules.scala 150:103:@36076.4]
  wire [6:0] _T_88541; // @[Modules.scala 150:103:@36122.4]
  wire [5:0] _T_88542; // @[Modules.scala 150:103:@36123.4]
  wire [5:0] _T_88543; // @[Modules.scala 150:103:@36124.4]
  wire [6:0] _T_88562; // @[Modules.scala 150:103:@36140.4]
  wire [5:0] _T_88563; // @[Modules.scala 150:103:@36141.4]
  wire [5:0] _T_88564; // @[Modules.scala 150:103:@36142.4]
  wire [5:0] _T_88580; // @[Modules.scala 150:74:@36156.4]
  wire [6:0] _T_88583; // @[Modules.scala 150:103:@36158.4]
  wire [5:0] _T_88584; // @[Modules.scala 150:103:@36159.4]
  wire [5:0] _T_88585; // @[Modules.scala 150:103:@36160.4]
  wire [5:0] _T_88590; // @[Modules.scala 150:103:@36164.4]
  wire [4:0] _T_88591; // @[Modules.scala 150:103:@36165.4]
  wire [4:0] _T_88592; // @[Modules.scala 150:103:@36166.4]
  wire [6:0] _T_88597; // @[Modules.scala 150:103:@36170.4]
  wire [5:0] _T_88598; // @[Modules.scala 150:103:@36171.4]
  wire [5:0] _T_88599; // @[Modules.scala 150:103:@36172.4]
  wire [5:0] _T_88604; // @[Modules.scala 150:103:@36176.4]
  wire [4:0] _T_88605; // @[Modules.scala 150:103:@36177.4]
  wire [4:0] _T_88606; // @[Modules.scala 150:103:@36178.4]
  wire [5:0] _GEN_776; // @[Modules.scala 150:103:@36188.4]
  wire [6:0] _T_88618; // @[Modules.scala 150:103:@36188.4]
  wire [5:0] _T_88619; // @[Modules.scala 150:103:@36189.4]
  wire [5:0] _T_88620; // @[Modules.scala 150:103:@36190.4]
  wire [6:0] _T_88639; // @[Modules.scala 150:103:@36206.4]
  wire [5:0] _T_88640; // @[Modules.scala 150:103:@36207.4]
  wire [5:0] _T_88641; // @[Modules.scala 150:103:@36208.4]
  wire [6:0] _T_88653; // @[Modules.scala 150:103:@36218.4]
  wire [5:0] _T_88654; // @[Modules.scala 150:103:@36219.4]
  wire [5:0] _T_88655; // @[Modules.scala 150:103:@36220.4]
  wire [5:0] _T_88681; // @[Modules.scala 150:103:@36242.4]
  wire [4:0] _T_88682; // @[Modules.scala 150:103:@36243.4]
  wire [4:0] _T_88683; // @[Modules.scala 150:103:@36244.4]
  wire [5:0] _GEN_777; // @[Modules.scala 150:103:@36254.4]
  wire [6:0] _T_88695; // @[Modules.scala 150:103:@36254.4]
  wire [5:0] _T_88696; // @[Modules.scala 150:103:@36255.4]
  wire [5:0] _T_88697; // @[Modules.scala 150:103:@36256.4]
  wire [6:0] _T_88702; // @[Modules.scala 150:103:@36260.4]
  wire [5:0] _T_88703; // @[Modules.scala 150:103:@36261.4]
  wire [5:0] _T_88704; // @[Modules.scala 150:103:@36262.4]
  wire [6:0] _T_88709; // @[Modules.scala 150:103:@36266.4]
  wire [5:0] _T_88710; // @[Modules.scala 150:103:@36267.4]
  wire [5:0] _T_88711; // @[Modules.scala 150:103:@36268.4]
  wire [6:0] _T_88716; // @[Modules.scala 150:103:@36272.4]
  wire [5:0] _T_88717; // @[Modules.scala 150:103:@36273.4]
  wire [5:0] _T_88718; // @[Modules.scala 150:103:@36274.4]
  wire [5:0] _GEN_779; // @[Modules.scala 150:103:@36284.4]
  wire [6:0] _T_88730; // @[Modules.scala 150:103:@36284.4]
  wire [5:0] _T_88731; // @[Modules.scala 150:103:@36285.4]
  wire [5:0] _T_88732; // @[Modules.scala 150:103:@36286.4]
  wire [5:0] _T_88765; // @[Modules.scala 150:103:@36314.4]
  wire [4:0] _T_88766; // @[Modules.scala 150:103:@36315.4]
  wire [4:0] _T_88767; // @[Modules.scala 150:103:@36316.4]
  wire [5:0] _GEN_781; // @[Modules.scala 150:103:@36332.4]
  wire [6:0] _T_88786; // @[Modules.scala 150:103:@36332.4]
  wire [5:0] _T_88787; // @[Modules.scala 150:103:@36333.4]
  wire [5:0] _T_88788; // @[Modules.scala 150:103:@36334.4]
  wire [5:0] _GEN_782; // @[Modules.scala 150:103:@36344.4]
  wire [6:0] _T_88800; // @[Modules.scala 150:103:@36344.4]
  wire [5:0] _T_88801; // @[Modules.scala 150:103:@36345.4]
  wire [5:0] _T_88802; // @[Modules.scala 150:103:@36346.4]
  wire [5:0] _T_88814; // @[Modules.scala 150:103:@36356.4]
  wire [4:0] _T_88815; // @[Modules.scala 150:103:@36357.4]
  wire [4:0] _T_88816; // @[Modules.scala 150:103:@36358.4]
  wire [5:0] _T_88835; // @[Modules.scala 150:103:@36374.4]
  wire [4:0] _T_88836; // @[Modules.scala 150:103:@36375.4]
  wire [4:0] _T_88837; // @[Modules.scala 150:103:@36376.4]
  wire [5:0] _GEN_783; // @[Modules.scala 150:103:@36392.4]
  wire [6:0] _T_88856; // @[Modules.scala 150:103:@36392.4]
  wire [5:0] _T_88857; // @[Modules.scala 150:103:@36393.4]
  wire [5:0] _T_88858; // @[Modules.scala 150:103:@36394.4]
  wire [5:0] _T_88940; // @[Modules.scala 150:103:@36464.4]
  wire [4:0] _T_88941; // @[Modules.scala 150:103:@36465.4]
  wire [4:0] _T_88942; // @[Modules.scala 150:103:@36466.4]
  wire [6:0] _T_88975; // @[Modules.scala 150:103:@36494.4]
  wire [5:0] _T_88976; // @[Modules.scala 150:103:@36495.4]
  wire [5:0] _T_88977; // @[Modules.scala 150:103:@36496.4]
  wire [5:0] _GEN_787; // @[Modules.scala 150:103:@36500.4]
  wire [6:0] _T_88982; // @[Modules.scala 150:103:@36500.4]
  wire [5:0] _T_88983; // @[Modules.scala 150:103:@36501.4]
  wire [5:0] _T_88984; // @[Modules.scala 150:103:@36502.4]
  wire [6:0] _T_89045; // @[Modules.scala 150:103:@36554.4]
  wire [5:0] _T_89046; // @[Modules.scala 150:103:@36555.4]
  wire [5:0] _T_89047; // @[Modules.scala 150:103:@36556.4]
  wire [6:0] _T_89052; // @[Modules.scala 150:103:@36560.4]
  wire [5:0] _T_89053; // @[Modules.scala 150:103:@36561.4]
  wire [5:0] _T_89054; // @[Modules.scala 150:103:@36562.4]
  wire [6:0] _T_89066; // @[Modules.scala 150:103:@36572.4]
  wire [5:0] _T_89067; // @[Modules.scala 150:103:@36573.4]
  wire [5:0] _T_89068; // @[Modules.scala 150:103:@36574.4]
  wire [6:0] _T_89073; // @[Modules.scala 150:103:@36578.4]
  wire [5:0] _T_89074; // @[Modules.scala 150:103:@36579.4]
  wire [5:0] _T_89075; // @[Modules.scala 150:103:@36580.4]
  wire [5:0] _T_89101; // @[Modules.scala 150:103:@36602.4]
  wire [4:0] _T_89102; // @[Modules.scala 150:103:@36603.4]
  wire [4:0] _T_89103; // @[Modules.scala 150:103:@36604.4]
  wire [5:0] _GEN_792; // @[Modules.scala 150:103:@36608.4]
  wire [6:0] _T_89108; // @[Modules.scala 150:103:@36608.4]
  wire [5:0] _T_89109; // @[Modules.scala 150:103:@36609.4]
  wire [5:0] _T_89110; // @[Modules.scala 150:103:@36610.4]
  wire [5:0] _T_89164; // @[Modules.scala 150:103:@36656.4]
  wire [4:0] _T_89165; // @[Modules.scala 150:103:@36657.4]
  wire [4:0] _T_89166; // @[Modules.scala 150:103:@36658.4]
  wire [6:0] _T_89220; // @[Modules.scala 150:103:@36704.4]
  wire [5:0] _T_89221; // @[Modules.scala 150:103:@36705.4]
  wire [5:0] _T_89222; // @[Modules.scala 150:103:@36706.4]
  wire [6:0] _T_89241; // @[Modules.scala 150:103:@36722.4]
  wire [5:0] _T_89242; // @[Modules.scala 150:103:@36723.4]
  wire [5:0] _T_89243; // @[Modules.scala 150:103:@36724.4]
  wire [6:0] _T_89248; // @[Modules.scala 150:103:@36728.4]
  wire [5:0] _T_89249; // @[Modules.scala 150:103:@36729.4]
  wire [5:0] _T_89250; // @[Modules.scala 150:103:@36730.4]
  wire [6:0] _T_89262; // @[Modules.scala 150:103:@36740.4]
  wire [5:0] _T_89263; // @[Modules.scala 150:103:@36741.4]
  wire [5:0] _T_89264; // @[Modules.scala 150:103:@36742.4]
  wire [6:0] _T_89276; // @[Modules.scala 150:103:@36752.4]
  wire [5:0] _T_89277; // @[Modules.scala 150:103:@36753.4]
  wire [5:0] _T_89278; // @[Modules.scala 150:103:@36754.4]
  wire [6:0] _T_89283; // @[Modules.scala 150:103:@36758.4]
  wire [5:0] _T_89284; // @[Modules.scala 150:103:@36759.4]
  wire [5:0] _T_89285; // @[Modules.scala 150:103:@36760.4]
  wire [6:0] _T_89332; // @[Modules.scala 150:103:@36800.4]
  wire [5:0] _T_89333; // @[Modules.scala 150:103:@36801.4]
  wire [5:0] _T_89334; // @[Modules.scala 150:103:@36802.4]
  wire [6:0] _T_89339; // @[Modules.scala 150:103:@36806.4]
  wire [5:0] _T_89340; // @[Modules.scala 150:103:@36807.4]
  wire [5:0] _T_89341; // @[Modules.scala 150:103:@36808.4]
  wire [5:0] _T_89345; // @[Modules.scala 151:80:@36811.4]
  wire [6:0] _T_89346; // @[Modules.scala 150:103:@36812.4]
  wire [5:0] _T_89347; // @[Modules.scala 150:103:@36813.4]
  wire [5:0] _T_89348; // @[Modules.scala 150:103:@36814.4]
  wire [6:0] _T_89381; // @[Modules.scala 150:103:@36842.4]
  wire [5:0] _T_89382; // @[Modules.scala 150:103:@36843.4]
  wire [5:0] _T_89383; // @[Modules.scala 150:103:@36844.4]
  wire [6:0] _T_89451; // @[Modules.scala 150:103:@36902.4]
  wire [5:0] _T_89452; // @[Modules.scala 150:103:@36903.4]
  wire [5:0] _T_89453; // @[Modules.scala 150:103:@36904.4]
  wire [6:0] _T_89486; // @[Modules.scala 150:103:@36932.4]
  wire [5:0] _T_89487; // @[Modules.scala 150:103:@36933.4]
  wire [5:0] _T_89488; // @[Modules.scala 150:103:@36934.4]
  wire [6:0] _T_89514; // @[Modules.scala 150:103:@36956.4]
  wire [5:0] _T_89515; // @[Modules.scala 150:103:@36957.4]
  wire [5:0] _T_89516; // @[Modules.scala 150:103:@36958.4]
  wire [6:0] _T_89521; // @[Modules.scala 150:103:@36962.4]
  wire [5:0] _T_89522; // @[Modules.scala 150:103:@36963.4]
  wire [5:0] _T_89523; // @[Modules.scala 150:103:@36964.4]
  wire [6:0] _T_89542; // @[Modules.scala 150:103:@36980.4]
  wire [5:0] _T_89543; // @[Modules.scala 150:103:@36981.4]
  wire [5:0] _T_89544; // @[Modules.scala 150:103:@36982.4]
  wire [5:0] _T_89556; // @[Modules.scala 150:103:@36992.4]
  wire [4:0] _T_89557; // @[Modules.scala 150:103:@36993.4]
  wire [4:0] _T_89558; // @[Modules.scala 150:103:@36994.4]
  wire [6:0] _T_89563; // @[Modules.scala 150:103:@36998.4]
  wire [5:0] _T_89564; // @[Modules.scala 150:103:@36999.4]
  wire [5:0] _T_89565; // @[Modules.scala 150:103:@37000.4]
  wire [6:0] _T_89577; // @[Modules.scala 150:103:@37010.4]
  wire [5:0] _T_89578; // @[Modules.scala 150:103:@37011.4]
  wire [5:0] _T_89579; // @[Modules.scala 150:103:@37012.4]
  wire [5:0] _T_89584; // @[Modules.scala 150:103:@37016.4]
  wire [4:0] _T_89585; // @[Modules.scala 150:103:@37017.4]
  wire [4:0] _T_89586; // @[Modules.scala 150:103:@37018.4]
  wire [6:0] _T_89598; // @[Modules.scala 150:103:@37028.4]
  wire [5:0] _T_89599; // @[Modules.scala 150:103:@37029.4]
  wire [5:0] _T_89600; // @[Modules.scala 150:103:@37030.4]
  wire [6:0] _T_89605; // @[Modules.scala 150:103:@37034.4]
  wire [5:0] _T_89606; // @[Modules.scala 150:103:@37035.4]
  wire [5:0] _T_89607; // @[Modules.scala 150:103:@37036.4]
  wire [5:0] _T_89633; // @[Modules.scala 150:103:@37058.4]
  wire [4:0] _T_89634; // @[Modules.scala 150:103:@37059.4]
  wire [4:0] _T_89635; // @[Modules.scala 150:103:@37060.4]
  wire [5:0] _T_89640; // @[Modules.scala 150:103:@37064.4]
  wire [4:0] _T_89641; // @[Modules.scala 150:103:@37065.4]
  wire [4:0] _T_89642; // @[Modules.scala 150:103:@37066.4]
  wire [5:0] _GEN_814; // @[Modules.scala 150:103:@37100.4]
  wire [6:0] _T_89682; // @[Modules.scala 150:103:@37100.4]
  wire [5:0] _T_89683; // @[Modules.scala 150:103:@37101.4]
  wire [5:0] _T_89684; // @[Modules.scala 150:103:@37102.4]
  wire [5:0] _T_89710; // @[Modules.scala 150:103:@37124.4]
  wire [4:0] _T_89711; // @[Modules.scala 150:103:@37125.4]
  wire [4:0] _T_89712; // @[Modules.scala 150:103:@37126.4]
  wire [6:0] _T_89766; // @[Modules.scala 150:103:@37172.4]
  wire [5:0] _T_89767; // @[Modules.scala 150:103:@37173.4]
  wire [5:0] _T_89768; // @[Modules.scala 150:103:@37174.4]
  wire [5:0] _T_89773; // @[Modules.scala 150:103:@37178.4]
  wire [4:0] _T_89774; // @[Modules.scala 150:103:@37179.4]
  wire [4:0] _T_89775; // @[Modules.scala 150:103:@37180.4]
  wire [5:0] _T_89780; // @[Modules.scala 150:103:@37184.4]
  wire [4:0] _T_89781; // @[Modules.scala 150:103:@37185.4]
  wire [4:0] _T_89782; // @[Modules.scala 150:103:@37186.4]
  wire [5:0] _T_89794; // @[Modules.scala 150:103:@37196.4]
  wire [4:0] _T_89795; // @[Modules.scala 150:103:@37197.4]
  wire [4:0] _T_89796; // @[Modules.scala 150:103:@37198.4]
  wire [6:0] _T_89801; // @[Modules.scala 150:103:@37202.4]
  wire [5:0] _T_89802; // @[Modules.scala 150:103:@37203.4]
  wire [5:0] _T_89803; // @[Modules.scala 150:103:@37204.4]
  wire [6:0] _T_89808; // @[Modules.scala 150:103:@37208.4]
  wire [5:0] _T_89809; // @[Modules.scala 150:103:@37209.4]
  wire [5:0] _T_89810; // @[Modules.scala 150:103:@37210.4]
  wire [6:0] _T_89815; // @[Modules.scala 150:103:@37214.4]
  wire [5:0] _T_89816; // @[Modules.scala 150:103:@37215.4]
  wire [5:0] _T_89817; // @[Modules.scala 150:103:@37216.4]
  wire [6:0] _T_89836; // @[Modules.scala 150:103:@37232.4]
  wire [5:0] _T_89837; // @[Modules.scala 150:103:@37233.4]
  wire [5:0] _T_89838; // @[Modules.scala 150:103:@37234.4]
  wire [5:0] _T_89843; // @[Modules.scala 150:103:@37238.4]
  wire [4:0] _T_89844; // @[Modules.scala 150:103:@37239.4]
  wire [4:0] _T_89845; // @[Modules.scala 150:103:@37240.4]
  wire [5:0] _GEN_818; // @[Modules.scala 150:103:@37250.4]
  wire [6:0] _T_89857; // @[Modules.scala 150:103:@37250.4]
  wire [5:0] _T_89858; // @[Modules.scala 150:103:@37251.4]
  wire [5:0] _T_89859; // @[Modules.scala 150:103:@37252.4]
  wire [5:0] _GEN_819; // @[Modules.scala 150:103:@37274.4]
  wire [6:0] _T_89885; // @[Modules.scala 150:103:@37274.4]
  wire [5:0] _T_89886; // @[Modules.scala 150:103:@37275.4]
  wire [5:0] _T_89887; // @[Modules.scala 150:103:@37276.4]
  wire [6:0] _T_89927; // @[Modules.scala 150:103:@37310.4]
  wire [5:0] _T_89928; // @[Modules.scala 150:103:@37311.4]
  wire [5:0] _T_89929; // @[Modules.scala 150:103:@37312.4]
  wire [5:0] _GEN_821; // @[Modules.scala 150:103:@37322.4]
  wire [6:0] _T_89941; // @[Modules.scala 150:103:@37322.4]
  wire [5:0] _T_89942; // @[Modules.scala 150:103:@37323.4]
  wire [5:0] _T_89943; // @[Modules.scala 150:103:@37324.4]
  wire [5:0] _T_89947; // @[Modules.scala 151:80:@37327.4]
  wire [5:0] _GEN_822; // @[Modules.scala 150:103:@37328.4]
  wire [6:0] _T_89948; // @[Modules.scala 150:103:@37328.4]
  wire [5:0] _T_89949; // @[Modules.scala 150:103:@37329.4]
  wire [5:0] _T_89950; // @[Modules.scala 150:103:@37330.4]
  wire [5:0] _T_89983; // @[Modules.scala 150:103:@37358.4]
  wire [4:0] _T_89984; // @[Modules.scala 150:103:@37359.4]
  wire [4:0] _T_89985; // @[Modules.scala 150:103:@37360.4]
  wire [6:0] _T_90018; // @[Modules.scala 150:103:@37388.4]
  wire [5:0] _T_90019; // @[Modules.scala 150:103:@37389.4]
  wire [5:0] _T_90020; // @[Modules.scala 150:103:@37390.4]
  wire [6:0] _T_90025; // @[Modules.scala 150:103:@37394.4]
  wire [5:0] _T_90026; // @[Modules.scala 150:103:@37395.4]
  wire [5:0] _T_90027; // @[Modules.scala 150:103:@37396.4]
  wire [6:0] _T_90032; // @[Modules.scala 150:103:@37400.4]
  wire [5:0] _T_90033; // @[Modules.scala 150:103:@37401.4]
  wire [5:0] _T_90034; // @[Modules.scala 150:103:@37402.4]
  wire [5:0] _T_90039; // @[Modules.scala 150:103:@37406.4]
  wire [4:0] _T_90040; // @[Modules.scala 150:103:@37407.4]
  wire [4:0] _T_90041; // @[Modules.scala 150:103:@37408.4]
  wire [5:0] _T_90046; // @[Modules.scala 150:103:@37412.4]
  wire [4:0] _T_90047; // @[Modules.scala 150:103:@37413.4]
  wire [4:0] _T_90048; // @[Modules.scala 150:103:@37414.4]
  wire [5:0] _T_90053; // @[Modules.scala 150:103:@37418.4]
  wire [4:0] _T_90054; // @[Modules.scala 150:103:@37419.4]
  wire [4:0] _T_90055; // @[Modules.scala 150:103:@37420.4]
  wire [5:0] _GEN_828; // @[Modules.scala 150:103:@37430.4]
  wire [6:0] _T_90067; // @[Modules.scala 150:103:@37430.4]
  wire [5:0] _T_90068; // @[Modules.scala 150:103:@37431.4]
  wire [5:0] _T_90069; // @[Modules.scala 150:103:@37432.4]
  wire [5:0] _T_90116; // @[Modules.scala 150:103:@37472.4]
  wire [4:0] _T_90117; // @[Modules.scala 150:103:@37473.4]
  wire [4:0] _T_90118; // @[Modules.scala 150:103:@37474.4]
  wire [6:0] _T_90172; // @[Modules.scala 150:103:@37520.4]
  wire [5:0] _T_90173; // @[Modules.scala 150:103:@37521.4]
  wire [5:0] _T_90174; // @[Modules.scala 150:103:@37522.4]
  wire [5:0] _GEN_831; // @[Modules.scala 150:103:@37532.4]
  wire [6:0] _T_90186; // @[Modules.scala 150:103:@37532.4]
  wire [5:0] _T_90187; // @[Modules.scala 150:103:@37533.4]
  wire [5:0] _T_90188; // @[Modules.scala 150:103:@37534.4]
  wire [5:0] _T_90214; // @[Modules.scala 150:103:@37556.4]
  wire [4:0] _T_90215; // @[Modules.scala 150:103:@37557.4]
  wire [4:0] _T_90216; // @[Modules.scala 150:103:@37558.4]
  wire [13:0] buffer_11_0; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90233; // @[Modules.scala 166:64:@37574.4]
  wire [13:0] _T_90234; // @[Modules.scala 166:64:@37575.4]
  wire [13:0] buffer_11_299; // @[Modules.scala 166:64:@37576.4]
  wire [13:0] buffer_11_2; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_3; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90236; // @[Modules.scala 166:64:@37578.4]
  wire [13:0] _T_90237; // @[Modules.scala 166:64:@37579.4]
  wire [13:0] buffer_11_300; // @[Modules.scala 166:64:@37580.4]
  wire [14:0] _T_90239; // @[Modules.scala 166:64:@37582.4]
  wire [13:0] _T_90240; // @[Modules.scala 166:64:@37583.4]
  wire [13:0] buffer_11_301; // @[Modules.scala 166:64:@37584.4]
  wire [14:0] _T_90242; // @[Modules.scala 166:64:@37586.4]
  wire [13:0] _T_90243; // @[Modules.scala 166:64:@37587.4]
  wire [13:0] buffer_11_302; // @[Modules.scala 166:64:@37588.4]
  wire [13:0] buffer_11_8; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90245; // @[Modules.scala 166:64:@37590.4]
  wire [13:0] _T_90246; // @[Modules.scala 166:64:@37591.4]
  wire [13:0] buffer_11_303; // @[Modules.scala 166:64:@37592.4]
  wire [13:0] buffer_11_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90248; // @[Modules.scala 166:64:@37594.4]
  wire [13:0] _T_90249; // @[Modules.scala 166:64:@37595.4]
  wire [13:0] buffer_11_304; // @[Modules.scala 166:64:@37596.4]
  wire [14:0] _T_90263; // @[Modules.scala 166:64:@37614.4]
  wire [13:0] _T_90264; // @[Modules.scala 166:64:@37615.4]
  wire [13:0] buffer_11_309; // @[Modules.scala 166:64:@37616.4]
  wire [13:0] buffer_11_22; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90266; // @[Modules.scala 166:64:@37618.4]
  wire [13:0] _T_90267; // @[Modules.scala 166:64:@37619.4]
  wire [13:0] buffer_11_310; // @[Modules.scala 166:64:@37620.4]
  wire [14:0] _T_90269; // @[Modules.scala 166:64:@37622.4]
  wire [13:0] _T_90270; // @[Modules.scala 166:64:@37623.4]
  wire [13:0] buffer_11_311; // @[Modules.scala 166:64:@37624.4]
  wire [14:0] _T_90272; // @[Modules.scala 166:64:@37626.4]
  wire [13:0] _T_90273; // @[Modules.scala 166:64:@37627.4]
  wire [13:0] buffer_11_312; // @[Modules.scala 166:64:@37628.4]
  wire [14:0] _T_90275; // @[Modules.scala 166:64:@37630.4]
  wire [13:0] _T_90276; // @[Modules.scala 166:64:@37631.4]
  wire [13:0] buffer_11_313; // @[Modules.scala 166:64:@37632.4]
  wire [13:0] buffer_11_34; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90284; // @[Modules.scala 166:64:@37642.4]
  wire [13:0] _T_90285; // @[Modules.scala 166:64:@37643.4]
  wire [13:0] buffer_11_316; // @[Modules.scala 166:64:@37644.4]
  wire [14:0] _T_90287; // @[Modules.scala 166:64:@37646.4]
  wire [13:0] _T_90288; // @[Modules.scala 166:64:@37647.4]
  wire [13:0] buffer_11_317; // @[Modules.scala 166:64:@37648.4]
  wire [14:0] _T_90290; // @[Modules.scala 166:64:@37650.4]
  wire [13:0] _T_90291; // @[Modules.scala 166:64:@37651.4]
  wire [13:0] buffer_11_318; // @[Modules.scala 166:64:@37652.4]
  wire [14:0] _T_90293; // @[Modules.scala 166:64:@37654.4]
  wire [13:0] _T_90294; // @[Modules.scala 166:64:@37655.4]
  wire [13:0] buffer_11_319; // @[Modules.scala 166:64:@37656.4]
  wire [13:0] buffer_11_42; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90296; // @[Modules.scala 166:64:@37658.4]
  wire [13:0] _T_90297; // @[Modules.scala 166:64:@37659.4]
  wire [13:0] buffer_11_320; // @[Modules.scala 166:64:@37660.4]
  wire [13:0] buffer_11_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90299; // @[Modules.scala 166:64:@37662.4]
  wire [13:0] _T_90300; // @[Modules.scala 166:64:@37663.4]
  wire [13:0] buffer_11_321; // @[Modules.scala 166:64:@37664.4]
  wire [14:0] _T_90302; // @[Modules.scala 166:64:@37666.4]
  wire [13:0] _T_90303; // @[Modules.scala 166:64:@37667.4]
  wire [13:0] buffer_11_322; // @[Modules.scala 166:64:@37668.4]
  wire [13:0] buffer_11_48; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90305; // @[Modules.scala 166:64:@37670.4]
  wire [13:0] _T_90306; // @[Modules.scala 166:64:@37671.4]
  wire [13:0] buffer_11_323; // @[Modules.scala 166:64:@37672.4]
  wire [14:0] _T_90308; // @[Modules.scala 166:64:@37674.4]
  wire [13:0] _T_90309; // @[Modules.scala 166:64:@37675.4]
  wire [13:0] buffer_11_324; // @[Modules.scala 166:64:@37676.4]
  wire [14:0] _T_90311; // @[Modules.scala 166:64:@37678.4]
  wire [13:0] _T_90312; // @[Modules.scala 166:64:@37679.4]
  wire [13:0] buffer_11_325; // @[Modules.scala 166:64:@37680.4]
  wire [14:0] _T_90314; // @[Modules.scala 166:64:@37682.4]
  wire [13:0] _T_90315; // @[Modules.scala 166:64:@37683.4]
  wire [13:0] buffer_11_326; // @[Modules.scala 166:64:@37684.4]
  wire [13:0] buffer_11_56; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90317; // @[Modules.scala 166:64:@37686.4]
  wire [13:0] _T_90318; // @[Modules.scala 166:64:@37687.4]
  wire [13:0] buffer_11_327; // @[Modules.scala 166:64:@37688.4]
  wire [13:0] buffer_11_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90320; // @[Modules.scala 166:64:@37690.4]
  wire [13:0] _T_90321; // @[Modules.scala 166:64:@37691.4]
  wire [13:0] buffer_11_328; // @[Modules.scala 166:64:@37692.4]
  wire [14:0] _T_90323; // @[Modules.scala 166:64:@37694.4]
  wire [13:0] _T_90324; // @[Modules.scala 166:64:@37695.4]
  wire [13:0] buffer_11_329; // @[Modules.scala 166:64:@37696.4]
  wire [13:0] buffer_11_62; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90326; // @[Modules.scala 166:64:@37698.4]
  wire [13:0] _T_90327; // @[Modules.scala 166:64:@37699.4]
  wire [13:0] buffer_11_330; // @[Modules.scala 166:64:@37700.4]
  wire [13:0] buffer_11_64; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_65; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90329; // @[Modules.scala 166:64:@37702.4]
  wire [13:0] _T_90330; // @[Modules.scala 166:64:@37703.4]
  wire [13:0] buffer_11_331; // @[Modules.scala 166:64:@37704.4]
  wire [13:0] buffer_11_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90332; // @[Modules.scala 166:64:@37706.4]
  wire [13:0] _T_90333; // @[Modules.scala 166:64:@37707.4]
  wire [13:0] buffer_11_332; // @[Modules.scala 166:64:@37708.4]
  wire [13:0] buffer_11_70; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90338; // @[Modules.scala 166:64:@37714.4]
  wire [13:0] _T_90339; // @[Modules.scala 166:64:@37715.4]
  wire [13:0] buffer_11_334; // @[Modules.scala 166:64:@37716.4]
  wire [13:0] buffer_11_72; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90341; // @[Modules.scala 166:64:@37718.4]
  wire [13:0] _T_90342; // @[Modules.scala 166:64:@37719.4]
  wire [13:0] buffer_11_335; // @[Modules.scala 166:64:@37720.4]
  wire [14:0] _T_90344; // @[Modules.scala 166:64:@37722.4]
  wire [13:0] _T_90345; // @[Modules.scala 166:64:@37723.4]
  wire [13:0] buffer_11_336; // @[Modules.scala 166:64:@37724.4]
  wire [13:0] buffer_11_76; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90347; // @[Modules.scala 166:64:@37726.4]
  wire [13:0] _T_90348; // @[Modules.scala 166:64:@37727.4]
  wire [13:0] buffer_11_337; // @[Modules.scala 166:64:@37728.4]
  wire [13:0] buffer_11_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90350; // @[Modules.scala 166:64:@37730.4]
  wire [13:0] _T_90351; // @[Modules.scala 166:64:@37731.4]
  wire [13:0] buffer_11_338; // @[Modules.scala 166:64:@37732.4]
  wire [13:0] buffer_11_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90353; // @[Modules.scala 166:64:@37734.4]
  wire [13:0] _T_90354; // @[Modules.scala 166:64:@37735.4]
  wire [13:0] buffer_11_339; // @[Modules.scala 166:64:@37736.4]
  wire [13:0] buffer_11_83; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90356; // @[Modules.scala 166:64:@37738.4]
  wire [13:0] _T_90357; // @[Modules.scala 166:64:@37739.4]
  wire [13:0] buffer_11_340; // @[Modules.scala 166:64:@37740.4]
  wire [14:0] _T_90359; // @[Modules.scala 166:64:@37742.4]
  wire [13:0] _T_90360; // @[Modules.scala 166:64:@37743.4]
  wire [13:0] buffer_11_341; // @[Modules.scala 166:64:@37744.4]
  wire [13:0] buffer_11_88; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90365; // @[Modules.scala 166:64:@37750.4]
  wire [13:0] _T_90366; // @[Modules.scala 166:64:@37751.4]
  wire [13:0] buffer_11_343; // @[Modules.scala 166:64:@37752.4]
  wire [13:0] buffer_11_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90368; // @[Modules.scala 166:64:@37754.4]
  wire [13:0] _T_90369; // @[Modules.scala 166:64:@37755.4]
  wire [13:0] buffer_11_344; // @[Modules.scala 166:64:@37756.4]
  wire [13:0] buffer_11_93; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90371; // @[Modules.scala 166:64:@37758.4]
  wire [13:0] _T_90372; // @[Modules.scala 166:64:@37759.4]
  wire [13:0] buffer_11_345; // @[Modules.scala 166:64:@37760.4]
  wire [13:0] buffer_11_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90374; // @[Modules.scala 166:64:@37762.4]
  wire [13:0] _T_90375; // @[Modules.scala 166:64:@37763.4]
  wire [13:0] buffer_11_346; // @[Modules.scala 166:64:@37764.4]
  wire [13:0] buffer_11_98; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90380; // @[Modules.scala 166:64:@37770.4]
  wire [13:0] _T_90381; // @[Modules.scala 166:64:@37771.4]
  wire [13:0] buffer_11_348; // @[Modules.scala 166:64:@37772.4]
  wire [13:0] buffer_11_101; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90383; // @[Modules.scala 166:64:@37774.4]
  wire [13:0] _T_90384; // @[Modules.scala 166:64:@37775.4]
  wire [13:0] buffer_11_349; // @[Modules.scala 166:64:@37776.4]
  wire [14:0] _T_90386; // @[Modules.scala 166:64:@37778.4]
  wire [13:0] _T_90387; // @[Modules.scala 166:64:@37779.4]
  wire [13:0] buffer_11_350; // @[Modules.scala 166:64:@37780.4]
  wire [14:0] _T_90389; // @[Modules.scala 166:64:@37782.4]
  wire [13:0] _T_90390; // @[Modules.scala 166:64:@37783.4]
  wire [13:0] buffer_11_351; // @[Modules.scala 166:64:@37784.4]
  wire [14:0] _T_90392; // @[Modules.scala 166:64:@37786.4]
  wire [13:0] _T_90393; // @[Modules.scala 166:64:@37787.4]
  wire [13:0] buffer_11_352; // @[Modules.scala 166:64:@37788.4]
  wire [14:0] _T_90395; // @[Modules.scala 166:64:@37790.4]
  wire [13:0] _T_90396; // @[Modules.scala 166:64:@37791.4]
  wire [13:0] buffer_11_353; // @[Modules.scala 166:64:@37792.4]
  wire [13:0] buffer_11_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90401; // @[Modules.scala 166:64:@37798.4]
  wire [13:0] _T_90402; // @[Modules.scala 166:64:@37799.4]
  wire [13:0] buffer_11_355; // @[Modules.scala 166:64:@37800.4]
  wire [14:0] _T_90404; // @[Modules.scala 166:64:@37802.4]
  wire [13:0] _T_90405; // @[Modules.scala 166:64:@37803.4]
  wire [13:0] buffer_11_356; // @[Modules.scala 166:64:@37804.4]
  wire [14:0] _T_90407; // @[Modules.scala 166:64:@37806.4]
  wire [13:0] _T_90408; // @[Modules.scala 166:64:@37807.4]
  wire [13:0] buffer_11_357; // @[Modules.scala 166:64:@37808.4]
  wire [13:0] buffer_11_118; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_119; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90410; // @[Modules.scala 166:64:@37810.4]
  wire [13:0] _T_90411; // @[Modules.scala 166:64:@37811.4]
  wire [13:0] buffer_11_358; // @[Modules.scala 166:64:@37812.4]
  wire [14:0] _T_90413; // @[Modules.scala 166:64:@37814.4]
  wire [13:0] _T_90414; // @[Modules.scala 166:64:@37815.4]
  wire [13:0] buffer_11_359; // @[Modules.scala 166:64:@37816.4]
  wire [14:0] _T_90419; // @[Modules.scala 166:64:@37822.4]
  wire [13:0] _T_90420; // @[Modules.scala 166:64:@37823.4]
  wire [13:0] buffer_11_361; // @[Modules.scala 166:64:@37824.4]
  wire [14:0] _T_90422; // @[Modules.scala 166:64:@37826.4]
  wire [13:0] _T_90423; // @[Modules.scala 166:64:@37827.4]
  wire [13:0] buffer_11_362; // @[Modules.scala 166:64:@37828.4]
  wire [13:0] buffer_11_128; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_129; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90425; // @[Modules.scala 166:64:@37830.4]
  wire [13:0] _T_90426; // @[Modules.scala 166:64:@37831.4]
  wire [13:0] buffer_11_363; // @[Modules.scala 166:64:@37832.4]
  wire [13:0] buffer_11_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90428; // @[Modules.scala 166:64:@37834.4]
  wire [13:0] _T_90429; // @[Modules.scala 166:64:@37835.4]
  wire [13:0] buffer_11_364; // @[Modules.scala 166:64:@37836.4]
  wire [13:0] buffer_11_132; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90431; // @[Modules.scala 166:64:@37838.4]
  wire [13:0] _T_90432; // @[Modules.scala 166:64:@37839.4]
  wire [13:0] buffer_11_365; // @[Modules.scala 166:64:@37840.4]
  wire [14:0] _T_90434; // @[Modules.scala 166:64:@37842.4]
  wire [13:0] _T_90435; // @[Modules.scala 166:64:@37843.4]
  wire [13:0] buffer_11_366; // @[Modules.scala 166:64:@37844.4]
  wire [13:0] buffer_11_136; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_137; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90437; // @[Modules.scala 166:64:@37846.4]
  wire [13:0] _T_90438; // @[Modules.scala 166:64:@37847.4]
  wire [13:0] buffer_11_367; // @[Modules.scala 166:64:@37848.4]
  wire [14:0] _T_90443; // @[Modules.scala 166:64:@37854.4]
  wire [13:0] _T_90444; // @[Modules.scala 166:64:@37855.4]
  wire [13:0] buffer_11_369; // @[Modules.scala 166:64:@37856.4]
  wire [13:0] buffer_11_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90449; // @[Modules.scala 166:64:@37862.4]
  wire [13:0] _T_90450; // @[Modules.scala 166:64:@37863.4]
  wire [13:0] buffer_11_371; // @[Modules.scala 166:64:@37864.4]
  wire [14:0] _T_90455; // @[Modules.scala 166:64:@37870.4]
  wire [13:0] _T_90456; // @[Modules.scala 166:64:@37871.4]
  wire [13:0] buffer_11_373; // @[Modules.scala 166:64:@37872.4]
  wire [13:0] buffer_11_153; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90461; // @[Modules.scala 166:64:@37878.4]
  wire [13:0] _T_90462; // @[Modules.scala 166:64:@37879.4]
  wire [13:0] buffer_11_375; // @[Modules.scala 166:64:@37880.4]
  wire [13:0] buffer_11_156; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_157; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90467; // @[Modules.scala 166:64:@37886.4]
  wire [13:0] _T_90468; // @[Modules.scala 166:64:@37887.4]
  wire [13:0] buffer_11_377; // @[Modules.scala 166:64:@37888.4]
  wire [13:0] buffer_11_159; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90470; // @[Modules.scala 166:64:@37890.4]
  wire [13:0] _T_90471; // @[Modules.scala 166:64:@37891.4]
  wire [13:0] buffer_11_378; // @[Modules.scala 166:64:@37892.4]
  wire [13:0] buffer_11_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90473; // @[Modules.scala 166:64:@37894.4]
  wire [13:0] _T_90474; // @[Modules.scala 166:64:@37895.4]
  wire [13:0] buffer_11_379; // @[Modules.scala 166:64:@37896.4]
  wire [13:0] buffer_11_162; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90476; // @[Modules.scala 166:64:@37898.4]
  wire [13:0] _T_90477; // @[Modules.scala 166:64:@37899.4]
  wire [13:0] buffer_11_380; // @[Modules.scala 166:64:@37900.4]
  wire [14:0] _T_90479; // @[Modules.scala 166:64:@37902.4]
  wire [13:0] _T_90480; // @[Modules.scala 166:64:@37903.4]
  wire [13:0] buffer_11_381; // @[Modules.scala 166:64:@37904.4]
  wire [13:0] buffer_11_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90485; // @[Modules.scala 166:64:@37910.4]
  wire [13:0] _T_90486; // @[Modules.scala 166:64:@37911.4]
  wire [13:0] buffer_11_383; // @[Modules.scala 166:64:@37912.4]
  wire [13:0] buffer_11_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90488; // @[Modules.scala 166:64:@37914.4]
  wire [13:0] _T_90489; // @[Modules.scala 166:64:@37915.4]
  wire [13:0] buffer_11_384; // @[Modules.scala 166:64:@37916.4]
  wire [14:0] _T_90491; // @[Modules.scala 166:64:@37918.4]
  wire [13:0] _T_90492; // @[Modules.scala 166:64:@37919.4]
  wire [13:0] buffer_11_385; // @[Modules.scala 166:64:@37920.4]
  wire [14:0] _T_90494; // @[Modules.scala 166:64:@37922.4]
  wire [13:0] _T_90495; // @[Modules.scala 166:64:@37923.4]
  wire [13:0] buffer_11_386; // @[Modules.scala 166:64:@37924.4]
  wire [13:0] buffer_11_176; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90497; // @[Modules.scala 166:64:@37926.4]
  wire [13:0] _T_90498; // @[Modules.scala 166:64:@37927.4]
  wire [13:0] buffer_11_387; // @[Modules.scala 166:64:@37928.4]
  wire [14:0] _T_90503; // @[Modules.scala 166:64:@37934.4]
  wire [13:0] _T_90504; // @[Modules.scala 166:64:@37935.4]
  wire [13:0] buffer_11_389; // @[Modules.scala 166:64:@37936.4]
  wire [14:0] _T_90509; // @[Modules.scala 166:64:@37942.4]
  wire [13:0] _T_90510; // @[Modules.scala 166:64:@37943.4]
  wire [13:0] buffer_11_391; // @[Modules.scala 166:64:@37944.4]
  wire [13:0] buffer_11_186; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90512; // @[Modules.scala 166:64:@37946.4]
  wire [13:0] _T_90513; // @[Modules.scala 166:64:@37947.4]
  wire [13:0] buffer_11_392; // @[Modules.scala 166:64:@37948.4]
  wire [14:0] _T_90515; // @[Modules.scala 166:64:@37950.4]
  wire [13:0] _T_90516; // @[Modules.scala 166:64:@37951.4]
  wire [13:0] buffer_11_393; // @[Modules.scala 166:64:@37952.4]
  wire [13:0] buffer_11_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90518; // @[Modules.scala 166:64:@37954.4]
  wire [13:0] _T_90519; // @[Modules.scala 166:64:@37955.4]
  wire [13:0] buffer_11_394; // @[Modules.scala 166:64:@37956.4]
  wire [13:0] buffer_11_195; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90524; // @[Modules.scala 166:64:@37962.4]
  wire [13:0] _T_90525; // @[Modules.scala 166:64:@37963.4]
  wire [13:0] buffer_11_396; // @[Modules.scala 166:64:@37964.4]
  wire [13:0] buffer_11_196; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90527; // @[Modules.scala 166:64:@37966.4]
  wire [13:0] _T_90528; // @[Modules.scala 166:64:@37967.4]
  wire [13:0] buffer_11_397; // @[Modules.scala 166:64:@37968.4]
  wire [13:0] buffer_11_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90530; // @[Modules.scala 166:64:@37970.4]
  wire [13:0] _T_90531; // @[Modules.scala 166:64:@37971.4]
  wire [13:0] buffer_11_398; // @[Modules.scala 166:64:@37972.4]
  wire [13:0] buffer_11_201; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90533; // @[Modules.scala 166:64:@37974.4]
  wire [13:0] _T_90534; // @[Modules.scala 166:64:@37975.4]
  wire [13:0] buffer_11_399; // @[Modules.scala 166:64:@37976.4]
  wire [13:0] buffer_11_202; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90536; // @[Modules.scala 166:64:@37978.4]
  wire [13:0] _T_90537; // @[Modules.scala 166:64:@37979.4]
  wire [13:0] buffer_11_400; // @[Modules.scala 166:64:@37980.4]
  wire [13:0] buffer_11_204; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90539; // @[Modules.scala 166:64:@37982.4]
  wire [13:0] _T_90540; // @[Modules.scala 166:64:@37983.4]
  wire [13:0] buffer_11_401; // @[Modules.scala 166:64:@37984.4]
  wire [13:0] buffer_11_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90542; // @[Modules.scala 166:64:@37986.4]
  wire [13:0] _T_90543; // @[Modules.scala 166:64:@37987.4]
  wire [13:0] buffer_11_402; // @[Modules.scala 166:64:@37988.4]
  wire [13:0] buffer_11_208; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90545; // @[Modules.scala 166:64:@37990.4]
  wire [13:0] _T_90546; // @[Modules.scala 166:64:@37991.4]
  wire [13:0] buffer_11_403; // @[Modules.scala 166:64:@37992.4]
  wire [13:0] buffer_11_212; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_213; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90551; // @[Modules.scala 166:64:@37998.4]
  wire [13:0] _T_90552; // @[Modules.scala 166:64:@37999.4]
  wire [13:0] buffer_11_405; // @[Modules.scala 166:64:@38000.4]
  wire [13:0] buffer_11_219; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90560; // @[Modules.scala 166:64:@38010.4]
  wire [13:0] _T_90561; // @[Modules.scala 166:64:@38011.4]
  wire [13:0] buffer_11_408; // @[Modules.scala 166:64:@38012.4]
  wire [14:0] _T_90563; // @[Modules.scala 166:64:@38014.4]
  wire [13:0] _T_90564; // @[Modules.scala 166:64:@38015.4]
  wire [13:0] buffer_11_409; // @[Modules.scala 166:64:@38016.4]
  wire [13:0] buffer_11_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90566; // @[Modules.scala 166:64:@38018.4]
  wire [13:0] _T_90567; // @[Modules.scala 166:64:@38019.4]
  wire [13:0] buffer_11_410; // @[Modules.scala 166:64:@38020.4]
  wire [14:0] _T_90569; // @[Modules.scala 166:64:@38022.4]
  wire [13:0] _T_90570; // @[Modules.scala 166:64:@38023.4]
  wire [13:0] buffer_11_411; // @[Modules.scala 166:64:@38024.4]
  wire [14:0] _T_90572; // @[Modules.scala 166:64:@38026.4]
  wire [13:0] _T_90573; // @[Modules.scala 166:64:@38027.4]
  wire [13:0] buffer_11_412; // @[Modules.scala 166:64:@38028.4]
  wire [14:0] _T_90575; // @[Modules.scala 166:64:@38030.4]
  wire [13:0] _T_90576; // @[Modules.scala 166:64:@38031.4]
  wire [13:0] buffer_11_413; // @[Modules.scala 166:64:@38032.4]
  wire [13:0] buffer_11_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90578; // @[Modules.scala 166:64:@38034.4]
  wire [13:0] _T_90579; // @[Modules.scala 166:64:@38035.4]
  wire [13:0] buffer_11_414; // @[Modules.scala 166:64:@38036.4]
  wire [13:0] buffer_11_232; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_233; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90581; // @[Modules.scala 166:64:@38038.4]
  wire [13:0] _T_90582; // @[Modules.scala 166:64:@38039.4]
  wire [13:0] buffer_11_415; // @[Modules.scala 166:64:@38040.4]
  wire [13:0] buffer_11_235; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90584; // @[Modules.scala 166:64:@38042.4]
  wire [13:0] _T_90585; // @[Modules.scala 166:64:@38043.4]
  wire [13:0] buffer_11_416; // @[Modules.scala 166:64:@38044.4]
  wire [13:0] buffer_11_236; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90587; // @[Modules.scala 166:64:@38046.4]
  wire [13:0] _T_90588; // @[Modules.scala 166:64:@38047.4]
  wire [13:0] buffer_11_417; // @[Modules.scala 166:64:@38048.4]
  wire [13:0] buffer_11_238; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90590; // @[Modules.scala 166:64:@38050.4]
  wire [13:0] _T_90591; // @[Modules.scala 166:64:@38051.4]
  wire [13:0] buffer_11_418; // @[Modules.scala 166:64:@38052.4]
  wire [13:0] buffer_11_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90593; // @[Modules.scala 166:64:@38054.4]
  wire [13:0] _T_90594; // @[Modules.scala 166:64:@38055.4]
  wire [13:0] buffer_11_419; // @[Modules.scala 166:64:@38056.4]
  wire [13:0] buffer_11_242; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90596; // @[Modules.scala 166:64:@38058.4]
  wire [13:0] _T_90597; // @[Modules.scala 166:64:@38059.4]
  wire [13:0] buffer_11_420; // @[Modules.scala 166:64:@38060.4]
  wire [13:0] buffer_11_244; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90599; // @[Modules.scala 166:64:@38062.4]
  wire [13:0] _T_90600; // @[Modules.scala 166:64:@38063.4]
  wire [13:0] buffer_11_421; // @[Modules.scala 166:64:@38064.4]
  wire [14:0] _T_90602; // @[Modules.scala 166:64:@38066.4]
  wire [13:0] _T_90603; // @[Modules.scala 166:64:@38067.4]
  wire [13:0] buffer_11_422; // @[Modules.scala 166:64:@38068.4]
  wire [13:0] buffer_11_248; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90605; // @[Modules.scala 166:64:@38070.4]
  wire [13:0] _T_90606; // @[Modules.scala 166:64:@38071.4]
  wire [13:0] buffer_11_423; // @[Modules.scala 166:64:@38072.4]
  wire [14:0] _T_90608; // @[Modules.scala 166:64:@38074.4]
  wire [13:0] _T_90609; // @[Modules.scala 166:64:@38075.4]
  wire [13:0] buffer_11_424; // @[Modules.scala 166:64:@38076.4]
  wire [14:0] _T_90611; // @[Modules.scala 166:64:@38078.4]
  wire [13:0] _T_90612; // @[Modules.scala 166:64:@38079.4]
  wire [13:0] buffer_11_425; // @[Modules.scala 166:64:@38080.4]
  wire [13:0] buffer_11_254; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90614; // @[Modules.scala 166:64:@38082.4]
  wire [13:0] _T_90615; // @[Modules.scala 166:64:@38083.4]
  wire [13:0] buffer_11_426; // @[Modules.scala 166:64:@38084.4]
  wire [13:0] buffer_11_256; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90617; // @[Modules.scala 166:64:@38086.4]
  wire [13:0] _T_90618; // @[Modules.scala 166:64:@38087.4]
  wire [13:0] buffer_11_427; // @[Modules.scala 166:64:@38088.4]
  wire [14:0] _T_90620; // @[Modules.scala 166:64:@38090.4]
  wire [13:0] _T_90621; // @[Modules.scala 166:64:@38091.4]
  wire [13:0] buffer_11_428; // @[Modules.scala 166:64:@38092.4]
  wire [13:0] buffer_11_262; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90626; // @[Modules.scala 166:64:@38098.4]
  wire [13:0] _T_90627; // @[Modules.scala 166:64:@38099.4]
  wire [13:0] buffer_11_430; // @[Modules.scala 166:64:@38100.4]
  wire [13:0] buffer_11_267; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90632; // @[Modules.scala 166:64:@38106.4]
  wire [13:0] _T_90633; // @[Modules.scala 166:64:@38107.4]
  wire [13:0] buffer_11_432; // @[Modules.scala 166:64:@38108.4]
  wire [13:0] buffer_11_268; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90635; // @[Modules.scala 166:64:@38110.4]
  wire [13:0] _T_90636; // @[Modules.scala 166:64:@38111.4]
  wire [13:0] buffer_11_433; // @[Modules.scala 166:64:@38112.4]
  wire [13:0] buffer_11_270; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_11_271; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90638; // @[Modules.scala 166:64:@38114.4]
  wire [13:0] _T_90639; // @[Modules.scala 166:64:@38115.4]
  wire [13:0] buffer_11_434; // @[Modules.scala 166:64:@38116.4]
  wire [13:0] buffer_11_272; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90641; // @[Modules.scala 166:64:@38118.4]
  wire [13:0] _T_90642; // @[Modules.scala 166:64:@38119.4]
  wire [13:0] buffer_11_435; // @[Modules.scala 166:64:@38120.4]
  wire [13:0] buffer_11_274; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90644; // @[Modules.scala 166:64:@38122.4]
  wire [13:0] _T_90645; // @[Modules.scala 166:64:@38123.4]
  wire [13:0] buffer_11_436; // @[Modules.scala 166:64:@38124.4]
  wire [14:0] _T_90650; // @[Modules.scala 166:64:@38130.4]
  wire [13:0] _T_90651; // @[Modules.scala 166:64:@38131.4]
  wire [13:0] buffer_11_438; // @[Modules.scala 166:64:@38132.4]
  wire [13:0] buffer_11_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90653; // @[Modules.scala 166:64:@38134.4]
  wire [13:0] _T_90654; // @[Modules.scala 166:64:@38135.4]
  wire [13:0] buffer_11_439; // @[Modules.scala 166:64:@38136.4]
  wire [14:0] _T_90659; // @[Modules.scala 166:64:@38142.4]
  wire [13:0] _T_90660; // @[Modules.scala 166:64:@38143.4]
  wire [13:0] buffer_11_441; // @[Modules.scala 166:64:@38144.4]
  wire [13:0] buffer_11_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90665; // @[Modules.scala 166:64:@38150.4]
  wire [13:0] _T_90666; // @[Modules.scala 166:64:@38151.4]
  wire [13:0] buffer_11_443; // @[Modules.scala 166:64:@38152.4]
  wire [13:0] buffer_11_291; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90668; // @[Modules.scala 166:64:@38154.4]
  wire [13:0] _T_90669; // @[Modules.scala 166:64:@38155.4]
  wire [13:0] buffer_11_444; // @[Modules.scala 166:64:@38156.4]
  wire [14:0] _T_90671; // @[Modules.scala 166:64:@38158.4]
  wire [13:0] _T_90672; // @[Modules.scala 166:64:@38159.4]
  wire [13:0] buffer_11_445; // @[Modules.scala 166:64:@38160.4]
  wire [13:0] buffer_11_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90674; // @[Modules.scala 166:64:@38162.4]
  wire [13:0] _T_90675; // @[Modules.scala 166:64:@38163.4]
  wire [13:0] buffer_11_446; // @[Modules.scala 166:64:@38164.4]
  wire [14:0] _T_90677; // @[Modules.scala 166:64:@38166.4]
  wire [13:0] _T_90678; // @[Modules.scala 166:64:@38167.4]
  wire [13:0] buffer_11_447; // @[Modules.scala 166:64:@38168.4]
  wire [14:0] _T_90680; // @[Modules.scala 166:64:@38170.4]
  wire [13:0] _T_90681; // @[Modules.scala 166:64:@38171.4]
  wire [13:0] buffer_11_448; // @[Modules.scala 166:64:@38172.4]
  wire [14:0] _T_90683; // @[Modules.scala 166:64:@38174.4]
  wire [13:0] _T_90684; // @[Modules.scala 166:64:@38175.4]
  wire [13:0] buffer_11_449; // @[Modules.scala 166:64:@38176.4]
  wire [14:0] _T_90686; // @[Modules.scala 166:64:@38178.4]
  wire [13:0] _T_90687; // @[Modules.scala 166:64:@38179.4]
  wire [13:0] buffer_11_450; // @[Modules.scala 166:64:@38180.4]
  wire [14:0] _T_90689; // @[Modules.scala 166:64:@38182.4]
  wire [13:0] _T_90690; // @[Modules.scala 166:64:@38183.4]
  wire [13:0] buffer_11_451; // @[Modules.scala 166:64:@38184.4]
  wire [14:0] _T_90695; // @[Modules.scala 166:64:@38190.4]
  wire [13:0] _T_90696; // @[Modules.scala 166:64:@38191.4]
  wire [13:0] buffer_11_453; // @[Modules.scala 166:64:@38192.4]
  wire [14:0] _T_90698; // @[Modules.scala 166:64:@38194.4]
  wire [13:0] _T_90699; // @[Modules.scala 166:64:@38195.4]
  wire [13:0] buffer_11_454; // @[Modules.scala 166:64:@38196.4]
  wire [14:0] _T_90701; // @[Modules.scala 166:64:@38198.4]
  wire [13:0] _T_90702; // @[Modules.scala 166:64:@38199.4]
  wire [13:0] buffer_11_455; // @[Modules.scala 166:64:@38200.4]
  wire [14:0] _T_90704; // @[Modules.scala 166:64:@38202.4]
  wire [13:0] _T_90705; // @[Modules.scala 166:64:@38203.4]
  wire [13:0] buffer_11_456; // @[Modules.scala 166:64:@38204.4]
  wire [14:0] _T_90707; // @[Modules.scala 166:64:@38206.4]
  wire [13:0] _T_90708; // @[Modules.scala 166:64:@38207.4]
  wire [13:0] buffer_11_457; // @[Modules.scala 166:64:@38208.4]
  wire [14:0] _T_90710; // @[Modules.scala 166:64:@38210.4]
  wire [13:0] _T_90711; // @[Modules.scala 166:64:@38211.4]
  wire [13:0] buffer_11_458; // @[Modules.scala 166:64:@38212.4]
  wire [14:0] _T_90713; // @[Modules.scala 166:64:@38214.4]
  wire [13:0] _T_90714; // @[Modules.scala 166:64:@38215.4]
  wire [13:0] buffer_11_459; // @[Modules.scala 166:64:@38216.4]
  wire [14:0] _T_90716; // @[Modules.scala 166:64:@38218.4]
  wire [13:0] _T_90717; // @[Modules.scala 166:64:@38219.4]
  wire [13:0] buffer_11_460; // @[Modules.scala 166:64:@38220.4]
  wire [14:0] _T_90719; // @[Modules.scala 166:64:@38222.4]
  wire [13:0] _T_90720; // @[Modules.scala 166:64:@38223.4]
  wire [13:0] buffer_11_461; // @[Modules.scala 166:64:@38224.4]
  wire [14:0] _T_90722; // @[Modules.scala 166:64:@38226.4]
  wire [13:0] _T_90723; // @[Modules.scala 166:64:@38227.4]
  wire [13:0] buffer_11_462; // @[Modules.scala 166:64:@38228.4]
  wire [14:0] _T_90725; // @[Modules.scala 166:64:@38230.4]
  wire [13:0] _T_90726; // @[Modules.scala 166:64:@38231.4]
  wire [13:0] buffer_11_463; // @[Modules.scala 166:64:@38232.4]
  wire [14:0] _T_90728; // @[Modules.scala 166:64:@38234.4]
  wire [13:0] _T_90729; // @[Modules.scala 166:64:@38235.4]
  wire [13:0] buffer_11_464; // @[Modules.scala 166:64:@38236.4]
  wire [14:0] _T_90731; // @[Modules.scala 166:64:@38238.4]
  wire [13:0] _T_90732; // @[Modules.scala 166:64:@38239.4]
  wire [13:0] buffer_11_465; // @[Modules.scala 166:64:@38240.4]
  wire [14:0] _T_90734; // @[Modules.scala 166:64:@38242.4]
  wire [13:0] _T_90735; // @[Modules.scala 166:64:@38243.4]
  wire [13:0] buffer_11_466; // @[Modules.scala 166:64:@38244.4]
  wire [14:0] _T_90737; // @[Modules.scala 166:64:@38246.4]
  wire [13:0] _T_90738; // @[Modules.scala 166:64:@38247.4]
  wire [13:0] buffer_11_467; // @[Modules.scala 166:64:@38248.4]
  wire [14:0] _T_90740; // @[Modules.scala 166:64:@38250.4]
  wire [13:0] _T_90741; // @[Modules.scala 166:64:@38251.4]
  wire [13:0] buffer_11_468; // @[Modules.scala 166:64:@38252.4]
  wire [14:0] _T_90743; // @[Modules.scala 166:64:@38254.4]
  wire [13:0] _T_90744; // @[Modules.scala 166:64:@38255.4]
  wire [13:0] buffer_11_469; // @[Modules.scala 166:64:@38256.4]
  wire [14:0] _T_90746; // @[Modules.scala 166:64:@38258.4]
  wire [13:0] _T_90747; // @[Modules.scala 166:64:@38259.4]
  wire [13:0] buffer_11_470; // @[Modules.scala 166:64:@38260.4]
  wire [14:0] _T_90749; // @[Modules.scala 166:64:@38262.4]
  wire [13:0] _T_90750; // @[Modules.scala 166:64:@38263.4]
  wire [13:0] buffer_11_471; // @[Modules.scala 166:64:@38264.4]
  wire [14:0] _T_90752; // @[Modules.scala 166:64:@38266.4]
  wire [13:0] _T_90753; // @[Modules.scala 166:64:@38267.4]
  wire [13:0] buffer_11_472; // @[Modules.scala 166:64:@38268.4]
  wire [14:0] _T_90755; // @[Modules.scala 166:64:@38270.4]
  wire [13:0] _T_90756; // @[Modules.scala 166:64:@38271.4]
  wire [13:0] buffer_11_473; // @[Modules.scala 166:64:@38272.4]
  wire [14:0] _T_90758; // @[Modules.scala 166:64:@38274.4]
  wire [13:0] _T_90759; // @[Modules.scala 166:64:@38275.4]
  wire [13:0] buffer_11_474; // @[Modules.scala 166:64:@38276.4]
  wire [14:0] _T_90761; // @[Modules.scala 166:64:@38278.4]
  wire [13:0] _T_90762; // @[Modules.scala 166:64:@38279.4]
  wire [13:0] buffer_11_475; // @[Modules.scala 166:64:@38280.4]
  wire [14:0] _T_90764; // @[Modules.scala 166:64:@38282.4]
  wire [13:0] _T_90765; // @[Modules.scala 166:64:@38283.4]
  wire [13:0] buffer_11_476; // @[Modules.scala 166:64:@38284.4]
  wire [14:0] _T_90767; // @[Modules.scala 166:64:@38286.4]
  wire [13:0] _T_90768; // @[Modules.scala 166:64:@38287.4]
  wire [13:0] buffer_11_477; // @[Modules.scala 166:64:@38288.4]
  wire [14:0] _T_90770; // @[Modules.scala 166:64:@38290.4]
  wire [13:0] _T_90771; // @[Modules.scala 166:64:@38291.4]
  wire [13:0] buffer_11_478; // @[Modules.scala 166:64:@38292.4]
  wire [14:0] _T_90773; // @[Modules.scala 166:64:@38294.4]
  wire [13:0] _T_90774; // @[Modules.scala 166:64:@38295.4]
  wire [13:0] buffer_11_479; // @[Modules.scala 166:64:@38296.4]
  wire [14:0] _T_90776; // @[Modules.scala 166:64:@38298.4]
  wire [13:0] _T_90777; // @[Modules.scala 166:64:@38299.4]
  wire [13:0] buffer_11_480; // @[Modules.scala 166:64:@38300.4]
  wire [14:0] _T_90779; // @[Modules.scala 166:64:@38302.4]
  wire [13:0] _T_90780; // @[Modules.scala 166:64:@38303.4]
  wire [13:0] buffer_11_481; // @[Modules.scala 166:64:@38304.4]
  wire [14:0] _T_90782; // @[Modules.scala 166:64:@38306.4]
  wire [13:0] _T_90783; // @[Modules.scala 166:64:@38307.4]
  wire [13:0] buffer_11_482; // @[Modules.scala 166:64:@38308.4]
  wire [14:0] _T_90785; // @[Modules.scala 166:64:@38310.4]
  wire [13:0] _T_90786; // @[Modules.scala 166:64:@38311.4]
  wire [13:0] buffer_11_483; // @[Modules.scala 166:64:@38312.4]
  wire [14:0] _T_90788; // @[Modules.scala 166:64:@38314.4]
  wire [13:0] _T_90789; // @[Modules.scala 166:64:@38315.4]
  wire [13:0] buffer_11_484; // @[Modules.scala 166:64:@38316.4]
  wire [14:0] _T_90791; // @[Modules.scala 166:64:@38318.4]
  wire [13:0] _T_90792; // @[Modules.scala 166:64:@38319.4]
  wire [13:0] buffer_11_485; // @[Modules.scala 166:64:@38320.4]
  wire [14:0] _T_90794; // @[Modules.scala 166:64:@38322.4]
  wire [13:0] _T_90795; // @[Modules.scala 166:64:@38323.4]
  wire [13:0] buffer_11_486; // @[Modules.scala 166:64:@38324.4]
  wire [14:0] _T_90797; // @[Modules.scala 166:64:@38326.4]
  wire [13:0] _T_90798; // @[Modules.scala 166:64:@38327.4]
  wire [13:0] buffer_11_487; // @[Modules.scala 166:64:@38328.4]
  wire [14:0] _T_90800; // @[Modules.scala 166:64:@38330.4]
  wire [13:0] _T_90801; // @[Modules.scala 166:64:@38331.4]
  wire [13:0] buffer_11_488; // @[Modules.scala 166:64:@38332.4]
  wire [14:0] _T_90803; // @[Modules.scala 166:64:@38334.4]
  wire [13:0] _T_90804; // @[Modules.scala 166:64:@38335.4]
  wire [13:0] buffer_11_489; // @[Modules.scala 166:64:@38336.4]
  wire [14:0] _T_90806; // @[Modules.scala 166:64:@38338.4]
  wire [13:0] _T_90807; // @[Modules.scala 166:64:@38339.4]
  wire [13:0] buffer_11_490; // @[Modules.scala 166:64:@38340.4]
  wire [14:0] _T_90809; // @[Modules.scala 166:64:@38342.4]
  wire [13:0] _T_90810; // @[Modules.scala 166:64:@38343.4]
  wire [13:0] buffer_11_491; // @[Modules.scala 166:64:@38344.4]
  wire [14:0] _T_90812; // @[Modules.scala 166:64:@38346.4]
  wire [13:0] _T_90813; // @[Modules.scala 166:64:@38347.4]
  wire [13:0] buffer_11_492; // @[Modules.scala 166:64:@38348.4]
  wire [14:0] _T_90815; // @[Modules.scala 166:64:@38350.4]
  wire [13:0] _T_90816; // @[Modules.scala 166:64:@38351.4]
  wire [13:0] buffer_11_493; // @[Modules.scala 166:64:@38352.4]
  wire [14:0] _T_90818; // @[Modules.scala 166:64:@38354.4]
  wire [13:0] _T_90819; // @[Modules.scala 166:64:@38355.4]
  wire [13:0] buffer_11_494; // @[Modules.scala 166:64:@38356.4]
  wire [14:0] _T_90821; // @[Modules.scala 166:64:@38358.4]
  wire [13:0] _T_90822; // @[Modules.scala 166:64:@38359.4]
  wire [13:0] buffer_11_495; // @[Modules.scala 166:64:@38360.4]
  wire [14:0] _T_90824; // @[Modules.scala 166:64:@38362.4]
  wire [13:0] _T_90825; // @[Modules.scala 166:64:@38363.4]
  wire [13:0] buffer_11_496; // @[Modules.scala 166:64:@38364.4]
  wire [14:0] _T_90827; // @[Modules.scala 166:64:@38366.4]
  wire [13:0] _T_90828; // @[Modules.scala 166:64:@38367.4]
  wire [13:0] buffer_11_497; // @[Modules.scala 166:64:@38368.4]
  wire [14:0] _T_90830; // @[Modules.scala 166:64:@38370.4]
  wire [13:0] _T_90831; // @[Modules.scala 166:64:@38371.4]
  wire [13:0] buffer_11_498; // @[Modules.scala 166:64:@38372.4]
  wire [14:0] _T_90833; // @[Modules.scala 166:64:@38374.4]
  wire [13:0] _T_90834; // @[Modules.scala 166:64:@38375.4]
  wire [13:0] buffer_11_499; // @[Modules.scala 166:64:@38376.4]
  wire [14:0] _T_90836; // @[Modules.scala 166:64:@38378.4]
  wire [13:0] _T_90837; // @[Modules.scala 166:64:@38379.4]
  wire [13:0] buffer_11_500; // @[Modules.scala 166:64:@38380.4]
  wire [14:0] _T_90839; // @[Modules.scala 166:64:@38382.4]
  wire [13:0] _T_90840; // @[Modules.scala 166:64:@38383.4]
  wire [13:0] buffer_11_501; // @[Modules.scala 166:64:@38384.4]
  wire [14:0] _T_90842; // @[Modules.scala 166:64:@38386.4]
  wire [13:0] _T_90843; // @[Modules.scala 166:64:@38387.4]
  wire [13:0] buffer_11_502; // @[Modules.scala 166:64:@38388.4]
  wire [14:0] _T_90845; // @[Modules.scala 166:64:@38390.4]
  wire [13:0] _T_90846; // @[Modules.scala 166:64:@38391.4]
  wire [13:0] buffer_11_503; // @[Modules.scala 166:64:@38392.4]
  wire [14:0] _T_90848; // @[Modules.scala 166:64:@38394.4]
  wire [13:0] _T_90849; // @[Modules.scala 166:64:@38395.4]
  wire [13:0] buffer_11_504; // @[Modules.scala 166:64:@38396.4]
  wire [14:0] _T_90851; // @[Modules.scala 166:64:@38398.4]
  wire [13:0] _T_90852; // @[Modules.scala 166:64:@38399.4]
  wire [13:0] buffer_11_505; // @[Modules.scala 166:64:@38400.4]
  wire [14:0] _T_90854; // @[Modules.scala 166:64:@38402.4]
  wire [13:0] _T_90855; // @[Modules.scala 166:64:@38403.4]
  wire [13:0] buffer_11_506; // @[Modules.scala 166:64:@38404.4]
  wire [14:0] _T_90857; // @[Modules.scala 166:64:@38406.4]
  wire [13:0] _T_90858; // @[Modules.scala 166:64:@38407.4]
  wire [13:0] buffer_11_507; // @[Modules.scala 166:64:@38408.4]
  wire [14:0] _T_90860; // @[Modules.scala 166:64:@38410.4]
  wire [13:0] _T_90861; // @[Modules.scala 166:64:@38411.4]
  wire [13:0] buffer_11_508; // @[Modules.scala 166:64:@38412.4]
  wire [14:0] _T_90863; // @[Modules.scala 166:64:@38414.4]
  wire [13:0] _T_90864; // @[Modules.scala 166:64:@38415.4]
  wire [13:0] buffer_11_509; // @[Modules.scala 166:64:@38416.4]
  wire [14:0] _T_90866; // @[Modules.scala 166:64:@38418.4]
  wire [13:0] _T_90867; // @[Modules.scala 166:64:@38419.4]
  wire [13:0] buffer_11_510; // @[Modules.scala 166:64:@38420.4]
  wire [14:0] _T_90869; // @[Modules.scala 166:64:@38422.4]
  wire [13:0] _T_90870; // @[Modules.scala 166:64:@38423.4]
  wire [13:0] buffer_11_511; // @[Modules.scala 166:64:@38424.4]
  wire [14:0] _T_90872; // @[Modules.scala 166:64:@38426.4]
  wire [13:0] _T_90873; // @[Modules.scala 166:64:@38427.4]
  wire [13:0] buffer_11_512; // @[Modules.scala 166:64:@38428.4]
  wire [14:0] _T_90875; // @[Modules.scala 166:64:@38430.4]
  wire [13:0] _T_90876; // @[Modules.scala 166:64:@38431.4]
  wire [13:0] buffer_11_513; // @[Modules.scala 166:64:@38432.4]
  wire [14:0] _T_90878; // @[Modules.scala 166:64:@38434.4]
  wire [13:0] _T_90879; // @[Modules.scala 166:64:@38435.4]
  wire [13:0] buffer_11_514; // @[Modules.scala 166:64:@38436.4]
  wire [14:0] _T_90881; // @[Modules.scala 166:64:@38438.4]
  wire [13:0] _T_90882; // @[Modules.scala 166:64:@38439.4]
  wire [13:0] buffer_11_515; // @[Modules.scala 166:64:@38440.4]
  wire [14:0] _T_90884; // @[Modules.scala 166:64:@38442.4]
  wire [13:0] _T_90885; // @[Modules.scala 166:64:@38443.4]
  wire [13:0] buffer_11_516; // @[Modules.scala 166:64:@38444.4]
  wire [14:0] _T_90887; // @[Modules.scala 166:64:@38446.4]
  wire [13:0] _T_90888; // @[Modules.scala 166:64:@38447.4]
  wire [13:0] buffer_11_517; // @[Modules.scala 166:64:@38448.4]
  wire [14:0] _T_90890; // @[Modules.scala 166:64:@38450.4]
  wire [13:0] _T_90891; // @[Modules.scala 166:64:@38451.4]
  wire [13:0] buffer_11_518; // @[Modules.scala 166:64:@38452.4]
  wire [14:0] _T_90893; // @[Modules.scala 166:64:@38454.4]
  wire [13:0] _T_90894; // @[Modules.scala 166:64:@38455.4]
  wire [13:0] buffer_11_519; // @[Modules.scala 166:64:@38456.4]
  wire [14:0] _T_90896; // @[Modules.scala 166:64:@38458.4]
  wire [13:0] _T_90897; // @[Modules.scala 166:64:@38459.4]
  wire [13:0] buffer_11_520; // @[Modules.scala 166:64:@38460.4]
  wire [14:0] _T_90899; // @[Modules.scala 166:64:@38462.4]
  wire [13:0] _T_90900; // @[Modules.scala 166:64:@38463.4]
  wire [13:0] buffer_11_521; // @[Modules.scala 166:64:@38464.4]
  wire [13:0] buffer_11_298; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_90902; // @[Modules.scala 172:66:@38466.4]
  wire [13:0] _T_90903; // @[Modules.scala 172:66:@38467.4]
  wire [13:0] buffer_11_522; // @[Modules.scala 172:66:@38468.4]
  wire [14:0] _T_90905; // @[Modules.scala 166:64:@38470.4]
  wire [13:0] _T_90906; // @[Modules.scala 166:64:@38471.4]
  wire [13:0] buffer_11_523; // @[Modules.scala 166:64:@38472.4]
  wire [14:0] _T_90908; // @[Modules.scala 166:64:@38474.4]
  wire [13:0] _T_90909; // @[Modules.scala 166:64:@38475.4]
  wire [13:0] buffer_11_524; // @[Modules.scala 166:64:@38476.4]
  wire [14:0] _T_90911; // @[Modules.scala 166:64:@38478.4]
  wire [13:0] _T_90912; // @[Modules.scala 166:64:@38479.4]
  wire [13:0] buffer_11_525; // @[Modules.scala 166:64:@38480.4]
  wire [14:0] _T_90914; // @[Modules.scala 166:64:@38482.4]
  wire [13:0] _T_90915; // @[Modules.scala 166:64:@38483.4]
  wire [13:0] buffer_11_526; // @[Modules.scala 166:64:@38484.4]
  wire [14:0] _T_90917; // @[Modules.scala 166:64:@38486.4]
  wire [13:0] _T_90918; // @[Modules.scala 166:64:@38487.4]
  wire [13:0] buffer_11_527; // @[Modules.scala 166:64:@38488.4]
  wire [14:0] _T_90920; // @[Modules.scala 166:64:@38490.4]
  wire [13:0] _T_90921; // @[Modules.scala 166:64:@38491.4]
  wire [13:0] buffer_11_528; // @[Modules.scala 166:64:@38492.4]
  wire [14:0] _T_90923; // @[Modules.scala 166:64:@38494.4]
  wire [13:0] _T_90924; // @[Modules.scala 166:64:@38495.4]
  wire [13:0] buffer_11_529; // @[Modules.scala 166:64:@38496.4]
  wire [14:0] _T_90926; // @[Modules.scala 166:64:@38498.4]
  wire [13:0] _T_90927; // @[Modules.scala 166:64:@38499.4]
  wire [13:0] buffer_11_530; // @[Modules.scala 166:64:@38500.4]
  wire [14:0] _T_90929; // @[Modules.scala 166:64:@38502.4]
  wire [13:0] _T_90930; // @[Modules.scala 166:64:@38503.4]
  wire [13:0] buffer_11_531; // @[Modules.scala 166:64:@38504.4]
  wire [14:0] _T_90932; // @[Modules.scala 166:64:@38506.4]
  wire [13:0] _T_90933; // @[Modules.scala 166:64:@38507.4]
  wire [13:0] buffer_11_532; // @[Modules.scala 166:64:@38508.4]
  wire [14:0] _T_90935; // @[Modules.scala 166:64:@38510.4]
  wire [13:0] _T_90936; // @[Modules.scala 166:64:@38511.4]
  wire [13:0] buffer_11_533; // @[Modules.scala 166:64:@38512.4]
  wire [14:0] _T_90938; // @[Modules.scala 166:64:@38514.4]
  wire [13:0] _T_90939; // @[Modules.scala 166:64:@38515.4]
  wire [13:0] buffer_11_534; // @[Modules.scala 166:64:@38516.4]
  wire [14:0] _T_90941; // @[Modules.scala 166:64:@38518.4]
  wire [13:0] _T_90942; // @[Modules.scala 166:64:@38519.4]
  wire [13:0] buffer_11_535; // @[Modules.scala 166:64:@38520.4]
  wire [14:0] _T_90944; // @[Modules.scala 166:64:@38522.4]
  wire [13:0] _T_90945; // @[Modules.scala 166:64:@38523.4]
  wire [13:0] buffer_11_536; // @[Modules.scala 166:64:@38524.4]
  wire [14:0] _T_90947; // @[Modules.scala 166:64:@38526.4]
  wire [13:0] _T_90948; // @[Modules.scala 166:64:@38527.4]
  wire [13:0] buffer_11_537; // @[Modules.scala 166:64:@38528.4]
  wire [14:0] _T_90950; // @[Modules.scala 166:64:@38530.4]
  wire [13:0] _T_90951; // @[Modules.scala 166:64:@38531.4]
  wire [13:0] buffer_11_538; // @[Modules.scala 166:64:@38532.4]
  wire [14:0] _T_90953; // @[Modules.scala 166:64:@38534.4]
  wire [13:0] _T_90954; // @[Modules.scala 166:64:@38535.4]
  wire [13:0] buffer_11_539; // @[Modules.scala 166:64:@38536.4]
  wire [14:0] _T_90956; // @[Modules.scala 166:64:@38538.4]
  wire [13:0] _T_90957; // @[Modules.scala 166:64:@38539.4]
  wire [13:0] buffer_11_540; // @[Modules.scala 166:64:@38540.4]
  wire [14:0] _T_90959; // @[Modules.scala 166:64:@38542.4]
  wire [13:0] _T_90960; // @[Modules.scala 166:64:@38543.4]
  wire [13:0] buffer_11_541; // @[Modules.scala 166:64:@38544.4]
  wire [14:0] _T_90962; // @[Modules.scala 166:64:@38546.4]
  wire [13:0] _T_90963; // @[Modules.scala 166:64:@38547.4]
  wire [13:0] buffer_11_542; // @[Modules.scala 166:64:@38548.4]
  wire [14:0] _T_90965; // @[Modules.scala 166:64:@38550.4]
  wire [13:0] _T_90966; // @[Modules.scala 166:64:@38551.4]
  wire [13:0] buffer_11_543; // @[Modules.scala 166:64:@38552.4]
  wire [14:0] _T_90968; // @[Modules.scala 166:64:@38554.4]
  wire [13:0] _T_90969; // @[Modules.scala 166:64:@38555.4]
  wire [13:0] buffer_11_544; // @[Modules.scala 166:64:@38556.4]
  wire [14:0] _T_90971; // @[Modules.scala 166:64:@38558.4]
  wire [13:0] _T_90972; // @[Modules.scala 166:64:@38559.4]
  wire [13:0] buffer_11_545; // @[Modules.scala 166:64:@38560.4]
  wire [14:0] _T_90974; // @[Modules.scala 166:64:@38562.4]
  wire [13:0] _T_90975; // @[Modules.scala 166:64:@38563.4]
  wire [13:0] buffer_11_546; // @[Modules.scala 166:64:@38564.4]
  wire [14:0] _T_90977; // @[Modules.scala 166:64:@38566.4]
  wire [13:0] _T_90978; // @[Modules.scala 166:64:@38567.4]
  wire [13:0] buffer_11_547; // @[Modules.scala 166:64:@38568.4]
  wire [14:0] _T_90980; // @[Modules.scala 166:64:@38570.4]
  wire [13:0] _T_90981; // @[Modules.scala 166:64:@38571.4]
  wire [13:0] buffer_11_548; // @[Modules.scala 166:64:@38572.4]
  wire [14:0] _T_90983; // @[Modules.scala 166:64:@38574.4]
  wire [13:0] _T_90984; // @[Modules.scala 166:64:@38575.4]
  wire [13:0] buffer_11_549; // @[Modules.scala 166:64:@38576.4]
  wire [14:0] _T_90986; // @[Modules.scala 166:64:@38578.4]
  wire [13:0] _T_90987; // @[Modules.scala 166:64:@38579.4]
  wire [13:0] buffer_11_550; // @[Modules.scala 166:64:@38580.4]
  wire [14:0] _T_90989; // @[Modules.scala 166:64:@38582.4]
  wire [13:0] _T_90990; // @[Modules.scala 166:64:@38583.4]
  wire [13:0] buffer_11_551; // @[Modules.scala 166:64:@38584.4]
  wire [14:0] _T_90992; // @[Modules.scala 166:64:@38586.4]
  wire [13:0] _T_90993; // @[Modules.scala 166:64:@38587.4]
  wire [13:0] buffer_11_552; // @[Modules.scala 166:64:@38588.4]
  wire [14:0] _T_90995; // @[Modules.scala 166:64:@38590.4]
  wire [13:0] _T_90996; // @[Modules.scala 166:64:@38591.4]
  wire [13:0] buffer_11_553; // @[Modules.scala 166:64:@38592.4]
  wire [14:0] _T_90998; // @[Modules.scala 166:64:@38594.4]
  wire [13:0] _T_90999; // @[Modules.scala 166:64:@38595.4]
  wire [13:0] buffer_11_554; // @[Modules.scala 166:64:@38596.4]
  wire [14:0] _T_91001; // @[Modules.scala 166:64:@38598.4]
  wire [13:0] _T_91002; // @[Modules.scala 166:64:@38599.4]
  wire [13:0] buffer_11_555; // @[Modules.scala 166:64:@38600.4]
  wire [14:0] _T_91004; // @[Modules.scala 166:64:@38602.4]
  wire [13:0] _T_91005; // @[Modules.scala 166:64:@38603.4]
  wire [13:0] buffer_11_556; // @[Modules.scala 166:64:@38604.4]
  wire [14:0] _T_91007; // @[Modules.scala 166:64:@38606.4]
  wire [13:0] _T_91008; // @[Modules.scala 166:64:@38607.4]
  wire [13:0] buffer_11_557; // @[Modules.scala 166:64:@38608.4]
  wire [14:0] _T_91010; // @[Modules.scala 166:64:@38610.4]
  wire [13:0] _T_91011; // @[Modules.scala 166:64:@38611.4]
  wire [13:0] buffer_11_558; // @[Modules.scala 166:64:@38612.4]
  wire [14:0] _T_91013; // @[Modules.scala 166:64:@38614.4]
  wire [13:0] _T_91014; // @[Modules.scala 166:64:@38615.4]
  wire [13:0] buffer_11_559; // @[Modules.scala 166:64:@38616.4]
  wire [14:0] _T_91016; // @[Modules.scala 166:64:@38618.4]
  wire [13:0] _T_91017; // @[Modules.scala 166:64:@38619.4]
  wire [13:0] buffer_11_560; // @[Modules.scala 166:64:@38620.4]
  wire [14:0] _T_91019; // @[Modules.scala 166:64:@38622.4]
  wire [13:0] _T_91020; // @[Modules.scala 166:64:@38623.4]
  wire [13:0] buffer_11_561; // @[Modules.scala 166:64:@38624.4]
  wire [14:0] _T_91022; // @[Modules.scala 166:64:@38626.4]
  wire [13:0] _T_91023; // @[Modules.scala 166:64:@38627.4]
  wire [13:0] buffer_11_562; // @[Modules.scala 166:64:@38628.4]
  wire [14:0] _T_91025; // @[Modules.scala 166:64:@38630.4]
  wire [13:0] _T_91026; // @[Modules.scala 166:64:@38631.4]
  wire [13:0] buffer_11_563; // @[Modules.scala 166:64:@38632.4]
  wire [14:0] _T_91028; // @[Modules.scala 166:64:@38634.4]
  wire [13:0] _T_91029; // @[Modules.scala 166:64:@38635.4]
  wire [13:0] buffer_11_564; // @[Modules.scala 166:64:@38636.4]
  wire [14:0] _T_91031; // @[Modules.scala 166:64:@38638.4]
  wire [13:0] _T_91032; // @[Modules.scala 166:64:@38639.4]
  wire [13:0] buffer_11_565; // @[Modules.scala 166:64:@38640.4]
  wire [14:0] _T_91034; // @[Modules.scala 166:64:@38642.4]
  wire [13:0] _T_91035; // @[Modules.scala 166:64:@38643.4]
  wire [13:0] buffer_11_566; // @[Modules.scala 166:64:@38644.4]
  wire [14:0] _T_91037; // @[Modules.scala 166:64:@38646.4]
  wire [13:0] _T_91038; // @[Modules.scala 166:64:@38647.4]
  wire [13:0] buffer_11_567; // @[Modules.scala 166:64:@38648.4]
  wire [14:0] _T_91040; // @[Modules.scala 166:64:@38650.4]
  wire [13:0] _T_91041; // @[Modules.scala 166:64:@38651.4]
  wire [13:0] buffer_11_568; // @[Modules.scala 166:64:@38652.4]
  wire [14:0] _T_91043; // @[Modules.scala 166:64:@38654.4]
  wire [13:0] _T_91044; // @[Modules.scala 166:64:@38655.4]
  wire [13:0] buffer_11_569; // @[Modules.scala 166:64:@38656.4]
  wire [14:0] _T_91046; // @[Modules.scala 166:64:@38658.4]
  wire [13:0] _T_91047; // @[Modules.scala 166:64:@38659.4]
  wire [13:0] buffer_11_570; // @[Modules.scala 166:64:@38660.4]
  wire [14:0] _T_91049; // @[Modules.scala 166:64:@38662.4]
  wire [13:0] _T_91050; // @[Modules.scala 166:64:@38663.4]
  wire [13:0] buffer_11_571; // @[Modules.scala 166:64:@38664.4]
  wire [14:0] _T_91052; // @[Modules.scala 166:64:@38666.4]
  wire [13:0] _T_91053; // @[Modules.scala 166:64:@38667.4]
  wire [13:0] buffer_11_572; // @[Modules.scala 166:64:@38668.4]
  wire [14:0] _T_91055; // @[Modules.scala 166:64:@38670.4]
  wire [13:0] _T_91056; // @[Modules.scala 166:64:@38671.4]
  wire [13:0] buffer_11_573; // @[Modules.scala 166:64:@38672.4]
  wire [14:0] _T_91058; // @[Modules.scala 166:64:@38674.4]
  wire [13:0] _T_91059; // @[Modules.scala 166:64:@38675.4]
  wire [13:0] buffer_11_574; // @[Modules.scala 166:64:@38676.4]
  wire [14:0] _T_91061; // @[Modules.scala 166:64:@38678.4]
  wire [13:0] _T_91062; // @[Modules.scala 166:64:@38679.4]
  wire [13:0] buffer_11_575; // @[Modules.scala 166:64:@38680.4]
  wire [14:0] _T_91064; // @[Modules.scala 166:64:@38682.4]
  wire [13:0] _T_91065; // @[Modules.scala 166:64:@38683.4]
  wire [13:0] buffer_11_576; // @[Modules.scala 166:64:@38684.4]
  wire [14:0] _T_91067; // @[Modules.scala 166:64:@38686.4]
  wire [13:0] _T_91068; // @[Modules.scala 166:64:@38687.4]
  wire [13:0] buffer_11_577; // @[Modules.scala 166:64:@38688.4]
  wire [14:0] _T_91070; // @[Modules.scala 172:66:@38690.4]
  wire [13:0] _T_91071; // @[Modules.scala 172:66:@38691.4]
  wire [13:0] buffer_11_578; // @[Modules.scala 172:66:@38692.4]
  wire [14:0] _T_91073; // @[Modules.scala 166:64:@38694.4]
  wire [13:0] _T_91074; // @[Modules.scala 166:64:@38695.4]
  wire [13:0] buffer_11_579; // @[Modules.scala 166:64:@38696.4]
  wire [14:0] _T_91076; // @[Modules.scala 166:64:@38698.4]
  wire [13:0] _T_91077; // @[Modules.scala 166:64:@38699.4]
  wire [13:0] buffer_11_580; // @[Modules.scala 166:64:@38700.4]
  wire [14:0] _T_91079; // @[Modules.scala 166:64:@38702.4]
  wire [13:0] _T_91080; // @[Modules.scala 166:64:@38703.4]
  wire [13:0] buffer_11_581; // @[Modules.scala 166:64:@38704.4]
  wire [14:0] _T_91082; // @[Modules.scala 166:64:@38706.4]
  wire [13:0] _T_91083; // @[Modules.scala 166:64:@38707.4]
  wire [13:0] buffer_11_582; // @[Modules.scala 166:64:@38708.4]
  wire [14:0] _T_91085; // @[Modules.scala 166:64:@38710.4]
  wire [13:0] _T_91086; // @[Modules.scala 166:64:@38711.4]
  wire [13:0] buffer_11_583; // @[Modules.scala 166:64:@38712.4]
  wire [14:0] _T_91088; // @[Modules.scala 166:64:@38714.4]
  wire [13:0] _T_91089; // @[Modules.scala 166:64:@38715.4]
  wire [13:0] buffer_11_584; // @[Modules.scala 166:64:@38716.4]
  wire [14:0] _T_91091; // @[Modules.scala 166:64:@38718.4]
  wire [13:0] _T_91092; // @[Modules.scala 166:64:@38719.4]
  wire [13:0] buffer_11_585; // @[Modules.scala 166:64:@38720.4]
  wire [14:0] _T_91094; // @[Modules.scala 166:64:@38722.4]
  wire [13:0] _T_91095; // @[Modules.scala 166:64:@38723.4]
  wire [13:0] buffer_11_586; // @[Modules.scala 166:64:@38724.4]
  wire [14:0] _T_91097; // @[Modules.scala 166:64:@38726.4]
  wire [13:0] _T_91098; // @[Modules.scala 166:64:@38727.4]
  wire [13:0] buffer_11_587; // @[Modules.scala 166:64:@38728.4]
  wire [14:0] _T_91100; // @[Modules.scala 166:64:@38730.4]
  wire [13:0] _T_91101; // @[Modules.scala 166:64:@38731.4]
  wire [13:0] buffer_11_588; // @[Modules.scala 166:64:@38732.4]
  wire [14:0] _T_91103; // @[Modules.scala 166:64:@38734.4]
  wire [13:0] _T_91104; // @[Modules.scala 166:64:@38735.4]
  wire [13:0] buffer_11_589; // @[Modules.scala 166:64:@38736.4]
  wire [14:0] _T_91106; // @[Modules.scala 166:64:@38738.4]
  wire [13:0] _T_91107; // @[Modules.scala 166:64:@38739.4]
  wire [13:0] buffer_11_590; // @[Modules.scala 166:64:@38740.4]
  wire [14:0] _T_91109; // @[Modules.scala 166:64:@38742.4]
  wire [13:0] _T_91110; // @[Modules.scala 166:64:@38743.4]
  wire [13:0] buffer_11_591; // @[Modules.scala 166:64:@38744.4]
  wire [14:0] _T_91112; // @[Modules.scala 172:66:@38746.4]
  wire [13:0] _T_91113; // @[Modules.scala 172:66:@38747.4]
  wire [13:0] buffer_11_592; // @[Modules.scala 172:66:@38748.4]
  wire [14:0] _T_91115; // @[Modules.scala 166:64:@38750.4]
  wire [13:0] _T_91116; // @[Modules.scala 166:64:@38751.4]
  wire [13:0] buffer_11_593; // @[Modules.scala 166:64:@38752.4]
  wire [14:0] _T_91118; // @[Modules.scala 166:64:@38754.4]
  wire [13:0] _T_91119; // @[Modules.scala 166:64:@38755.4]
  wire [13:0] buffer_11_594; // @[Modules.scala 166:64:@38756.4]
  wire [14:0] _T_91121; // @[Modules.scala 160:64:@38758.4]
  wire [13:0] _T_91122; // @[Modules.scala 160:64:@38759.4]
  wire [13:0] buffer_11_595; // @[Modules.scala 160:64:@38760.4]
  wire [14:0] _T_91124; // @[Modules.scala 172:66:@38762.4]
  wire [13:0] _T_91125; // @[Modules.scala 172:66:@38763.4]
  wire [13:0] buffer_11_596; // @[Modules.scala 172:66:@38764.4]
  wire [5:0] _T_91128; // @[Modules.scala 143:74:@38953.4]
  wire [5:0] _GEN_832; // @[Modules.scala 143:103:@38955.4]
  wire [6:0] _T_91131; // @[Modules.scala 143:103:@38955.4]
  wire [5:0] _T_91132; // @[Modules.scala 143:103:@38956.4]
  wire [5:0] _T_91133; // @[Modules.scala 143:103:@38957.4]
  wire [5:0] _GEN_833; // @[Modules.scala 143:103:@38961.4]
  wire [6:0] _T_91138; // @[Modules.scala 143:103:@38961.4]
  wire [5:0] _T_91139; // @[Modules.scala 143:103:@38962.4]
  wire [5:0] _T_91140; // @[Modules.scala 143:103:@38963.4]
  wire [6:0] _T_91166; // @[Modules.scala 143:103:@38985.4]
  wire [5:0] _T_91167; // @[Modules.scala 143:103:@38986.4]
  wire [5:0] _T_91168; // @[Modules.scala 143:103:@38987.4]
  wire [5:0] _GEN_834; // @[Modules.scala 143:103:@39009.4]
  wire [6:0] _T_91194; // @[Modules.scala 143:103:@39009.4]
  wire [5:0] _T_91195; // @[Modules.scala 143:103:@39010.4]
  wire [5:0] _T_91196; // @[Modules.scala 143:103:@39011.4]
  wire [5:0] _T_91207; // @[Modules.scala 144:80:@39020.4]
  wire [6:0] _T_91208; // @[Modules.scala 143:103:@39021.4]
  wire [5:0] _T_91209; // @[Modules.scala 143:103:@39022.4]
  wire [5:0] _T_91210; // @[Modules.scala 143:103:@39023.4]
  wire [5:0] _T_91222; // @[Modules.scala 143:103:@39033.4]
  wire [4:0] _T_91223; // @[Modules.scala 143:103:@39034.4]
  wire [4:0] _T_91224; // @[Modules.scala 143:103:@39035.4]
  wire [5:0] _GEN_835; // @[Modules.scala 143:103:@39039.4]
  wire [6:0] _T_91229; // @[Modules.scala 143:103:@39039.4]
  wire [5:0] _T_91230; // @[Modules.scala 143:103:@39040.4]
  wire [5:0] _T_91231; // @[Modules.scala 143:103:@39041.4]
  wire [5:0] _GEN_836; // @[Modules.scala 143:103:@39045.4]
  wire [6:0] _T_91236; // @[Modules.scala 143:103:@39045.4]
  wire [5:0] _T_91237; // @[Modules.scala 143:103:@39046.4]
  wire [5:0] _T_91238; // @[Modules.scala 143:103:@39047.4]
  wire [5:0] _GEN_837; // @[Modules.scala 143:103:@39051.4]
  wire [6:0] _T_91243; // @[Modules.scala 143:103:@39051.4]
  wire [5:0] _T_91244; // @[Modules.scala 143:103:@39052.4]
  wire [5:0] _T_91245; // @[Modules.scala 143:103:@39053.4]
  wire [5:0] _GEN_838; // @[Modules.scala 143:103:@39057.4]
  wire [6:0] _T_91250; // @[Modules.scala 143:103:@39057.4]
  wire [5:0] _T_91251; // @[Modules.scala 143:103:@39058.4]
  wire [5:0] _T_91252; // @[Modules.scala 143:103:@39059.4]
  wire [5:0] _T_91320; // @[Modules.scala 143:103:@39117.4]
  wire [4:0] _T_91321; // @[Modules.scala 143:103:@39118.4]
  wire [4:0] _T_91322; // @[Modules.scala 143:103:@39119.4]
  wire [6:0] _T_91362; // @[Modules.scala 143:103:@39153.4]
  wire [5:0] _T_91363; // @[Modules.scala 143:103:@39154.4]
  wire [5:0] _T_91364; // @[Modules.scala 143:103:@39155.4]
  wire [5:0] _GEN_843; // @[Modules.scala 143:103:@39165.4]
  wire [6:0] _T_91376; // @[Modules.scala 143:103:@39165.4]
  wire [5:0] _T_91377; // @[Modules.scala 143:103:@39166.4]
  wire [5:0] _T_91378; // @[Modules.scala 143:103:@39167.4]
  wire [5:0] _T_91383; // @[Modules.scala 143:103:@39171.4]
  wire [4:0] _T_91384; // @[Modules.scala 143:103:@39172.4]
  wire [4:0] _T_91385; // @[Modules.scala 143:103:@39173.4]
  wire [6:0] _T_91397; // @[Modules.scala 143:103:@39183.4]
  wire [5:0] _T_91398; // @[Modules.scala 143:103:@39184.4]
  wire [5:0] _T_91399; // @[Modules.scala 143:103:@39185.4]
  wire [6:0] _T_91418; // @[Modules.scala 143:103:@39201.4]
  wire [5:0] _T_91419; // @[Modules.scala 143:103:@39202.4]
  wire [5:0] _T_91420; // @[Modules.scala 143:103:@39203.4]
  wire [6:0] _T_91432; // @[Modules.scala 143:103:@39213.4]
  wire [5:0] _T_91433; // @[Modules.scala 143:103:@39214.4]
  wire [5:0] _T_91434; // @[Modules.scala 143:103:@39215.4]
  wire [5:0] _T_91439; // @[Modules.scala 143:103:@39219.4]
  wire [4:0] _T_91440; // @[Modules.scala 143:103:@39220.4]
  wire [4:0] _T_91441; // @[Modules.scala 143:103:@39221.4]
  wire [5:0] _GEN_845; // @[Modules.scala 143:103:@39225.4]
  wire [6:0] _T_91446; // @[Modules.scala 143:103:@39225.4]
  wire [5:0] _T_91447; // @[Modules.scala 143:103:@39226.4]
  wire [5:0] _T_91448; // @[Modules.scala 143:103:@39227.4]
  wire [6:0] _T_91453; // @[Modules.scala 143:103:@39231.4]
  wire [5:0] _T_91454; // @[Modules.scala 143:103:@39232.4]
  wire [5:0] _T_91455; // @[Modules.scala 143:103:@39233.4]
  wire [6:0] _T_91481; // @[Modules.scala 143:103:@39255.4]
  wire [5:0] _T_91482; // @[Modules.scala 143:103:@39256.4]
  wire [5:0] _T_91483; // @[Modules.scala 143:103:@39257.4]
  wire [6:0] _T_91488; // @[Modules.scala 143:103:@39261.4]
  wire [5:0] _T_91489; // @[Modules.scala 143:103:@39262.4]
  wire [5:0] _T_91490; // @[Modules.scala 143:103:@39263.4]
  wire [6:0] _T_91502; // @[Modules.scala 143:103:@39273.4]
  wire [5:0] _T_91503; // @[Modules.scala 143:103:@39274.4]
  wire [5:0] _T_91504; // @[Modules.scala 143:103:@39275.4]
  wire [6:0] _T_91530; // @[Modules.scala 143:103:@39297.4]
  wire [5:0] _T_91531; // @[Modules.scala 143:103:@39298.4]
  wire [5:0] _T_91532; // @[Modules.scala 143:103:@39299.4]
  wire [6:0] _T_91551; // @[Modules.scala 143:103:@39315.4]
  wire [5:0] _T_91552; // @[Modules.scala 143:103:@39316.4]
  wire [5:0] _T_91553; // @[Modules.scala 143:103:@39317.4]
  wire [6:0] _T_91558; // @[Modules.scala 143:103:@39321.4]
  wire [5:0] _T_91559; // @[Modules.scala 143:103:@39322.4]
  wire [5:0] _T_91560; // @[Modules.scala 143:103:@39323.4]
  wire [5:0] _GEN_850; // @[Modules.scala 143:103:@39327.4]
  wire [6:0] _T_91565; // @[Modules.scala 143:103:@39327.4]
  wire [5:0] _T_91566; // @[Modules.scala 143:103:@39328.4]
  wire [5:0] _T_91567; // @[Modules.scala 143:103:@39329.4]
  wire [6:0] _T_91600; // @[Modules.scala 143:103:@39357.4]
  wire [5:0] _T_91601; // @[Modules.scala 143:103:@39358.4]
  wire [5:0] _T_91602; // @[Modules.scala 143:103:@39359.4]
  wire [6:0] _T_91621; // @[Modules.scala 143:103:@39375.4]
  wire [5:0] _T_91622; // @[Modules.scala 143:103:@39376.4]
  wire [5:0] _T_91623; // @[Modules.scala 143:103:@39377.4]
  wire [5:0] _T_91642; // @[Modules.scala 143:103:@39393.4]
  wire [4:0] _T_91643; // @[Modules.scala 143:103:@39394.4]
  wire [4:0] _T_91644; // @[Modules.scala 143:103:@39395.4]
  wire [5:0] _GEN_854; // @[Modules.scala 143:103:@39399.4]
  wire [6:0] _T_91649; // @[Modules.scala 143:103:@39399.4]
  wire [5:0] _T_91650; // @[Modules.scala 143:103:@39400.4]
  wire [5:0] _T_91651; // @[Modules.scala 143:103:@39401.4]
  wire [5:0] _GEN_855; // @[Modules.scala 143:103:@39405.4]
  wire [6:0] _T_91656; // @[Modules.scala 143:103:@39405.4]
  wire [5:0] _T_91657; // @[Modules.scala 143:103:@39406.4]
  wire [5:0] _T_91658; // @[Modules.scala 143:103:@39407.4]
  wire [6:0] _T_91663; // @[Modules.scala 143:103:@39411.4]
  wire [5:0] _T_91664; // @[Modules.scala 143:103:@39412.4]
  wire [5:0] _T_91665; // @[Modules.scala 143:103:@39413.4]
  wire [6:0] _T_91698; // @[Modules.scala 143:103:@39441.4]
  wire [5:0] _T_91699; // @[Modules.scala 143:103:@39442.4]
  wire [5:0] _T_91700; // @[Modules.scala 143:103:@39443.4]
  wire [5:0] _GEN_858; // @[Modules.scala 143:103:@39483.4]
  wire [6:0] _T_91747; // @[Modules.scala 143:103:@39483.4]
  wire [5:0] _T_91748; // @[Modules.scala 143:103:@39484.4]
  wire [5:0] _T_91749; // @[Modules.scala 143:103:@39485.4]
  wire [6:0] _T_91768; // @[Modules.scala 143:103:@39501.4]
  wire [5:0] _T_91769; // @[Modules.scala 143:103:@39502.4]
  wire [5:0] _T_91770; // @[Modules.scala 143:103:@39503.4]
  wire [5:0] _T_91775; // @[Modules.scala 143:103:@39507.4]
  wire [4:0] _T_91776; // @[Modules.scala 143:103:@39508.4]
  wire [4:0] _T_91777; // @[Modules.scala 143:103:@39509.4]
  wire [5:0] _GEN_860; // @[Modules.scala 143:103:@39519.4]
  wire [6:0] _T_91789; // @[Modules.scala 143:103:@39519.4]
  wire [5:0] _T_91790; // @[Modules.scala 143:103:@39520.4]
  wire [5:0] _T_91791; // @[Modules.scala 143:103:@39521.4]
  wire [6:0] _T_91859; // @[Modules.scala 143:103:@39579.4]
  wire [5:0] _T_91860; // @[Modules.scala 143:103:@39580.4]
  wire [5:0] _T_91861; // @[Modules.scala 143:103:@39581.4]
  wire [6:0] _T_91866; // @[Modules.scala 143:103:@39585.4]
  wire [5:0] _T_91867; // @[Modules.scala 143:103:@39586.4]
  wire [5:0] _T_91868; // @[Modules.scala 143:103:@39587.4]
  wire [6:0] _T_91873; // @[Modules.scala 143:103:@39591.4]
  wire [5:0] _T_91874; // @[Modules.scala 143:103:@39592.4]
  wire [5:0] _T_91875; // @[Modules.scala 143:103:@39593.4]
  wire [5:0] _T_91950; // @[Modules.scala 143:103:@39657.4]
  wire [4:0] _T_91951; // @[Modules.scala 143:103:@39658.4]
  wire [4:0] _T_91952; // @[Modules.scala 143:103:@39659.4]
  wire [5:0] _T_91957; // @[Modules.scala 143:103:@39663.4]
  wire [4:0] _T_91958; // @[Modules.scala 143:103:@39664.4]
  wire [4:0] _T_91959; // @[Modules.scala 143:103:@39665.4]
  wire [5:0] _GEN_865; // @[Modules.scala 143:103:@39687.4]
  wire [6:0] _T_91985; // @[Modules.scala 143:103:@39687.4]
  wire [5:0] _T_91986; // @[Modules.scala 143:103:@39688.4]
  wire [5:0] _T_91987; // @[Modules.scala 143:103:@39689.4]
  wire [6:0] _T_92013; // @[Modules.scala 143:103:@39711.4]
  wire [5:0] _T_92014; // @[Modules.scala 143:103:@39712.4]
  wire [5:0] _T_92015; // @[Modules.scala 143:103:@39713.4]
  wire [5:0] _T_92027; // @[Modules.scala 143:103:@39723.4]
  wire [4:0] _T_92028; // @[Modules.scala 143:103:@39724.4]
  wire [4:0] _T_92029; // @[Modules.scala 143:103:@39725.4]
  wire [5:0] _T_92048; // @[Modules.scala 143:103:@39741.4]
  wire [4:0] _T_92049; // @[Modules.scala 143:103:@39742.4]
  wire [4:0] _T_92050; // @[Modules.scala 143:103:@39743.4]
  wire [5:0] _GEN_872; // @[Modules.scala 143:103:@39855.4]
  wire [6:0] _T_92181; // @[Modules.scala 143:103:@39855.4]
  wire [5:0] _T_92182; // @[Modules.scala 143:103:@39856.4]
  wire [5:0] _T_92183; // @[Modules.scala 143:103:@39857.4]
  wire [5:0] _T_92251; // @[Modules.scala 143:103:@39915.4]
  wire [4:0] _T_92252; // @[Modules.scala 143:103:@39916.4]
  wire [4:0] _T_92253; // @[Modules.scala 143:103:@39917.4]
  wire [5:0] _GEN_874; // @[Modules.scala 143:103:@39951.4]
  wire [6:0] _T_92293; // @[Modules.scala 143:103:@39951.4]
  wire [5:0] _T_92294; // @[Modules.scala 143:103:@39952.4]
  wire [5:0] _T_92295; // @[Modules.scala 143:103:@39953.4]
  wire [6:0] _T_92321; // @[Modules.scala 143:103:@39975.4]
  wire [5:0] _T_92322; // @[Modules.scala 143:103:@39976.4]
  wire [5:0] _T_92323; // @[Modules.scala 143:103:@39977.4]
  wire [5:0] _GEN_876; // @[Modules.scala 143:103:@39981.4]
  wire [6:0] _T_92328; // @[Modules.scala 143:103:@39981.4]
  wire [5:0] _T_92329; // @[Modules.scala 143:103:@39982.4]
  wire [5:0] _T_92330; // @[Modules.scala 143:103:@39983.4]
  wire [5:0] _T_92335; // @[Modules.scala 143:103:@39987.4]
  wire [4:0] _T_92336; // @[Modules.scala 143:103:@39988.4]
  wire [4:0] _T_92337; // @[Modules.scala 143:103:@39989.4]
  wire [5:0] _T_92349; // @[Modules.scala 143:103:@39999.4]
  wire [4:0] _T_92350; // @[Modules.scala 143:103:@40000.4]
  wire [4:0] _T_92351; // @[Modules.scala 143:103:@40001.4]
  wire [5:0] _GEN_878; // @[Modules.scala 143:103:@40023.4]
  wire [6:0] _T_92377; // @[Modules.scala 143:103:@40023.4]
  wire [5:0] _T_92378; // @[Modules.scala 143:103:@40024.4]
  wire [5:0] _T_92379; // @[Modules.scala 143:103:@40025.4]
  wire [5:0] _T_92405; // @[Modules.scala 143:103:@40047.4]
  wire [4:0] _T_92406; // @[Modules.scala 143:103:@40048.4]
  wire [4:0] _T_92407; // @[Modules.scala 143:103:@40049.4]
  wire [6:0] _T_92503; // @[Modules.scala 143:103:@40131.4]
  wire [5:0] _T_92504; // @[Modules.scala 143:103:@40132.4]
  wire [5:0] _T_92505; // @[Modules.scala 143:103:@40133.4]
  wire [6:0] _T_92510; // @[Modules.scala 143:103:@40137.4]
  wire [5:0] _T_92511; // @[Modules.scala 143:103:@40138.4]
  wire [5:0] _T_92512; // @[Modules.scala 143:103:@40139.4]
  wire [6:0] _T_92573; // @[Modules.scala 143:103:@40191.4]
  wire [5:0] _T_92574; // @[Modules.scala 143:103:@40192.4]
  wire [5:0] _T_92575; // @[Modules.scala 143:103:@40193.4]
  wire [6:0] _T_92580; // @[Modules.scala 143:103:@40197.4]
  wire [5:0] _T_92581; // @[Modules.scala 143:103:@40198.4]
  wire [5:0] _T_92582; // @[Modules.scala 143:103:@40199.4]
  wire [5:0] _GEN_884; // @[Modules.scala 143:103:@40203.4]
  wire [6:0] _T_92587; // @[Modules.scala 143:103:@40203.4]
  wire [5:0] _T_92588; // @[Modules.scala 143:103:@40204.4]
  wire [5:0] _T_92589; // @[Modules.scala 143:103:@40205.4]
  wire [6:0] _T_92636; // @[Modules.scala 143:103:@40245.4]
  wire [5:0] _T_92637; // @[Modules.scala 143:103:@40246.4]
  wire [5:0] _T_92638; // @[Modules.scala 143:103:@40247.4]
  wire [6:0] _T_92643; // @[Modules.scala 143:103:@40251.4]
  wire [5:0] _T_92644; // @[Modules.scala 143:103:@40252.4]
  wire [5:0] _T_92645; // @[Modules.scala 143:103:@40253.4]
  wire [5:0] _GEN_886; // @[Modules.scala 143:103:@40275.4]
  wire [6:0] _T_92671; // @[Modules.scala 143:103:@40275.4]
  wire [5:0] _T_92672; // @[Modules.scala 143:103:@40276.4]
  wire [5:0] _T_92673; // @[Modules.scala 143:103:@40277.4]
  wire [6:0] _T_92720; // @[Modules.scala 143:103:@40317.4]
  wire [5:0] _T_92721; // @[Modules.scala 143:103:@40318.4]
  wire [5:0] _T_92722; // @[Modules.scala 143:103:@40319.4]
  wire [6:0] _T_92727; // @[Modules.scala 143:103:@40323.4]
  wire [5:0] _T_92728; // @[Modules.scala 143:103:@40324.4]
  wire [5:0] _T_92729; // @[Modules.scala 143:103:@40325.4]
  wire [6:0] _T_92734; // @[Modules.scala 143:103:@40329.4]
  wire [5:0] _T_92735; // @[Modules.scala 143:103:@40330.4]
  wire [5:0] _T_92736; // @[Modules.scala 143:103:@40331.4]
  wire [5:0] _GEN_888; // @[Modules.scala 143:103:@40335.4]
  wire [6:0] _T_92741; // @[Modules.scala 143:103:@40335.4]
  wire [5:0] _T_92742; // @[Modules.scala 143:103:@40336.4]
  wire [5:0] _T_92743; // @[Modules.scala 143:103:@40337.4]
  wire [5:0] _GEN_889; // @[Modules.scala 143:103:@40341.4]
  wire [6:0] _T_92748; // @[Modules.scala 143:103:@40341.4]
  wire [5:0] _T_92749; // @[Modules.scala 143:103:@40342.4]
  wire [5:0] _T_92750; // @[Modules.scala 143:103:@40343.4]
  wire [5:0] _GEN_891; // @[Modules.scala 143:103:@40383.4]
  wire [6:0] _T_92797; // @[Modules.scala 143:103:@40383.4]
  wire [5:0] _T_92798; // @[Modules.scala 143:103:@40384.4]
  wire [5:0] _T_92799; // @[Modules.scala 143:103:@40385.4]
  wire [6:0] _T_92804; // @[Modules.scala 143:103:@40389.4]
  wire [5:0] _T_92805; // @[Modules.scala 143:103:@40390.4]
  wire [5:0] _T_92806; // @[Modules.scala 143:103:@40391.4]
  wire [6:0] _T_92811; // @[Modules.scala 143:103:@40395.4]
  wire [5:0] _T_92812; // @[Modules.scala 143:103:@40396.4]
  wire [5:0] _T_92813; // @[Modules.scala 143:103:@40397.4]
  wire [6:0] _T_92825; // @[Modules.scala 143:103:@40407.4]
  wire [5:0] _T_92826; // @[Modules.scala 143:103:@40408.4]
  wire [5:0] _T_92827; // @[Modules.scala 143:103:@40409.4]
  wire [6:0] _T_92846; // @[Modules.scala 143:103:@40425.4]
  wire [5:0] _T_92847; // @[Modules.scala 143:103:@40426.4]
  wire [5:0] _T_92848; // @[Modules.scala 143:103:@40427.4]
  wire [6:0] _T_92888; // @[Modules.scala 143:103:@40461.4]
  wire [5:0] _T_92889; // @[Modules.scala 143:103:@40462.4]
  wire [5:0] _T_92890; // @[Modules.scala 143:103:@40463.4]
  wire [6:0] _T_92902; // @[Modules.scala 143:103:@40473.4]
  wire [5:0] _T_92903; // @[Modules.scala 143:103:@40474.4]
  wire [5:0] _T_92904; // @[Modules.scala 143:103:@40475.4]
  wire [5:0] _T_92909; // @[Modules.scala 143:103:@40479.4]
  wire [4:0] _T_92910; // @[Modules.scala 143:103:@40480.4]
  wire [4:0] _T_92911; // @[Modules.scala 143:103:@40481.4]
  wire [5:0] _T_92916; // @[Modules.scala 143:103:@40485.4]
  wire [4:0] _T_92917; // @[Modules.scala 143:103:@40486.4]
  wire [4:0] _T_92918; // @[Modules.scala 143:103:@40487.4]
  wire [6:0] _T_92923; // @[Modules.scala 143:103:@40491.4]
  wire [5:0] _T_92924; // @[Modules.scala 143:103:@40492.4]
  wire [5:0] _T_92925; // @[Modules.scala 143:103:@40493.4]
  wire [6:0] _T_92958; // @[Modules.scala 143:103:@40521.4]
  wire [5:0] _T_92959; // @[Modules.scala 143:103:@40522.4]
  wire [5:0] _T_92960; // @[Modules.scala 143:103:@40523.4]
  wire [6:0] _T_92972; // @[Modules.scala 143:103:@40533.4]
  wire [5:0] _T_92973; // @[Modules.scala 143:103:@40534.4]
  wire [5:0] _T_92974; // @[Modules.scala 143:103:@40535.4]
  wire [6:0] _T_92993; // @[Modules.scala 143:103:@40551.4]
  wire [5:0] _T_92994; // @[Modules.scala 143:103:@40552.4]
  wire [5:0] _T_92995; // @[Modules.scala 143:103:@40553.4]
  wire [6:0] _T_93007; // @[Modules.scala 143:103:@40563.4]
  wire [5:0] _T_93008; // @[Modules.scala 143:103:@40564.4]
  wire [5:0] _T_93009; // @[Modules.scala 143:103:@40565.4]
  wire [5:0] _GEN_903; // @[Modules.scala 143:103:@40593.4]
  wire [6:0] _T_93042; // @[Modules.scala 143:103:@40593.4]
  wire [5:0] _T_93043; // @[Modules.scala 143:103:@40594.4]
  wire [5:0] _T_93044; // @[Modules.scala 143:103:@40595.4]
  wire [5:0] _GEN_904; // @[Modules.scala 143:103:@40611.4]
  wire [6:0] _T_93063; // @[Modules.scala 143:103:@40611.4]
  wire [5:0] _T_93064; // @[Modules.scala 143:103:@40612.4]
  wire [5:0] _T_93065; // @[Modules.scala 143:103:@40613.4]
  wire [5:0] _T_93077; // @[Modules.scala 143:103:@40623.4]
  wire [4:0] _T_93078; // @[Modules.scala 143:103:@40624.4]
  wire [4:0] _T_93079; // @[Modules.scala 143:103:@40625.4]
  wire [6:0] _T_93091; // @[Modules.scala 143:103:@40635.4]
  wire [5:0] _T_93092; // @[Modules.scala 143:103:@40636.4]
  wire [5:0] _T_93093; // @[Modules.scala 143:103:@40637.4]
  wire [5:0] _T_93154; // @[Modules.scala 143:103:@40689.4]
  wire [4:0] _T_93155; // @[Modules.scala 143:103:@40690.4]
  wire [4:0] _T_93156; // @[Modules.scala 143:103:@40691.4]
  wire [6:0] _T_93203; // @[Modules.scala 143:103:@40731.4]
  wire [5:0] _T_93204; // @[Modules.scala 143:103:@40732.4]
  wire [5:0] _T_93205; // @[Modules.scala 143:103:@40733.4]
  wire [13:0] buffer_12_0; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93213; // @[Modules.scala 160:64:@40741.4]
  wire [13:0] _T_93214; // @[Modules.scala 160:64:@40742.4]
  wire [13:0] buffer_12_298; // @[Modules.scala 160:64:@40743.4]
  wire [13:0] buffer_12_5; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93219; // @[Modules.scala 160:64:@40749.4]
  wire [13:0] _T_93220; // @[Modules.scala 160:64:@40750.4]
  wire [13:0] buffer_12_300; // @[Modules.scala 160:64:@40751.4]
  wire [13:0] buffer_12_9; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93225; // @[Modules.scala 160:64:@40757.4]
  wire [13:0] _T_93226; // @[Modules.scala 160:64:@40758.4]
  wire [13:0] buffer_12_302; // @[Modules.scala 160:64:@40759.4]
  wire [13:0] buffer_12_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93228; // @[Modules.scala 160:64:@40761.4]
  wire [13:0] _T_93229; // @[Modules.scala 160:64:@40762.4]
  wire [13:0] buffer_12_303; // @[Modules.scala 160:64:@40763.4]
  wire [13:0] buffer_12_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93231; // @[Modules.scala 160:64:@40765.4]
  wire [13:0] _T_93232; // @[Modules.scala 160:64:@40766.4]
  wire [13:0] buffer_12_304; // @[Modules.scala 160:64:@40767.4]
  wire [13:0] buffer_12_14; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_15; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93234; // @[Modules.scala 160:64:@40769.4]
  wire [13:0] _T_93235; // @[Modules.scala 160:64:@40770.4]
  wire [13:0] buffer_12_305; // @[Modules.scala 160:64:@40771.4]
  wire [13:0] buffer_12_16; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_17; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93237; // @[Modules.scala 160:64:@40773.4]
  wire [13:0] _T_93238; // @[Modules.scala 160:64:@40774.4]
  wire [13:0] buffer_12_306; // @[Modules.scala 160:64:@40775.4]
  wire [14:0] _T_93240; // @[Modules.scala 160:64:@40777.4]
  wire [13:0] _T_93241; // @[Modules.scala 160:64:@40778.4]
  wire [13:0] buffer_12_307; // @[Modules.scala 160:64:@40779.4]
  wire [14:0] _T_93243; // @[Modules.scala 160:64:@40781.4]
  wire [13:0] _T_93244; // @[Modules.scala 160:64:@40782.4]
  wire [13:0] buffer_12_308; // @[Modules.scala 160:64:@40783.4]
  wire [13:0] buffer_12_27; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93252; // @[Modules.scala 160:64:@40793.4]
  wire [13:0] _T_93253; // @[Modules.scala 160:64:@40794.4]
  wire [13:0] buffer_12_311; // @[Modules.scala 160:64:@40795.4]
  wire [14:0] _T_93255; // @[Modules.scala 160:64:@40797.4]
  wire [13:0] _T_93256; // @[Modules.scala 160:64:@40798.4]
  wire [13:0] buffer_12_312; // @[Modules.scala 160:64:@40799.4]
  wire [14:0] _T_93258; // @[Modules.scala 160:64:@40801.4]
  wire [13:0] _T_93259; // @[Modules.scala 160:64:@40802.4]
  wire [13:0] buffer_12_313; // @[Modules.scala 160:64:@40803.4]
  wire [13:0] buffer_12_33; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93261; // @[Modules.scala 160:64:@40805.4]
  wire [13:0] _T_93262; // @[Modules.scala 160:64:@40806.4]
  wire [13:0] buffer_12_314; // @[Modules.scala 160:64:@40807.4]
  wire [13:0] buffer_12_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93264; // @[Modules.scala 160:64:@40809.4]
  wire [13:0] _T_93265; // @[Modules.scala 160:64:@40810.4]
  wire [13:0] buffer_12_315; // @[Modules.scala 160:64:@40811.4]
  wire [13:0] buffer_12_36; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93267; // @[Modules.scala 160:64:@40813.4]
  wire [13:0] _T_93268; // @[Modules.scala 160:64:@40814.4]
  wire [13:0] buffer_12_316; // @[Modules.scala 160:64:@40815.4]
  wire [13:0] buffer_12_38; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93270; // @[Modules.scala 160:64:@40817.4]
  wire [13:0] _T_93271; // @[Modules.scala 160:64:@40818.4]
  wire [13:0] buffer_12_317; // @[Modules.scala 160:64:@40819.4]
  wire [13:0] buffer_12_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93273; // @[Modules.scala 160:64:@40821.4]
  wire [13:0] _T_93274; // @[Modules.scala 160:64:@40822.4]
  wire [13:0] buffer_12_318; // @[Modules.scala 160:64:@40823.4]
  wire [13:0] buffer_12_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93276; // @[Modules.scala 160:64:@40825.4]
  wire [13:0] _T_93277; // @[Modules.scala 160:64:@40826.4]
  wire [13:0] buffer_12_319; // @[Modules.scala 160:64:@40827.4]
  wire [13:0] buffer_12_44; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93279; // @[Modules.scala 160:64:@40829.4]
  wire [13:0] _T_93280; // @[Modules.scala 160:64:@40830.4]
  wire [13:0] buffer_12_320; // @[Modules.scala 160:64:@40831.4]
  wire [13:0] buffer_12_46; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93282; // @[Modules.scala 160:64:@40833.4]
  wire [13:0] _T_93283; // @[Modules.scala 160:64:@40834.4]
  wire [13:0] buffer_12_321; // @[Modules.scala 160:64:@40835.4]
  wire [14:0] _T_93285; // @[Modules.scala 160:64:@40837.4]
  wire [13:0] _T_93286; // @[Modules.scala 160:64:@40838.4]
  wire [13:0] buffer_12_322; // @[Modules.scala 160:64:@40839.4]
  wire [13:0] buffer_12_50; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_51; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93288; // @[Modules.scala 160:64:@40841.4]
  wire [13:0] _T_93289; // @[Modules.scala 160:64:@40842.4]
  wire [13:0] buffer_12_323; // @[Modules.scala 160:64:@40843.4]
  wire [13:0] buffer_12_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93291; // @[Modules.scala 160:64:@40845.4]
  wire [13:0] _T_93292; // @[Modules.scala 160:64:@40846.4]
  wire [13:0] buffer_12_324; // @[Modules.scala 160:64:@40847.4]
  wire [14:0] _T_93294; // @[Modules.scala 160:64:@40849.4]
  wire [13:0] _T_93295; // @[Modules.scala 160:64:@40850.4]
  wire [13:0] buffer_12_325; // @[Modules.scala 160:64:@40851.4]
  wire [13:0] buffer_12_57; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93297; // @[Modules.scala 160:64:@40853.4]
  wire [13:0] _T_93298; // @[Modules.scala 160:64:@40854.4]
  wire [13:0] buffer_12_326; // @[Modules.scala 160:64:@40855.4]
  wire [14:0] _T_93300; // @[Modules.scala 160:64:@40857.4]
  wire [13:0] _T_93301; // @[Modules.scala 160:64:@40858.4]
  wire [13:0] buffer_12_327; // @[Modules.scala 160:64:@40859.4]
  wire [13:0] buffer_12_60; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93303; // @[Modules.scala 160:64:@40861.4]
  wire [13:0] _T_93304; // @[Modules.scala 160:64:@40862.4]
  wire [13:0] buffer_12_328; // @[Modules.scala 160:64:@40863.4]
  wire [13:0] buffer_12_62; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93306; // @[Modules.scala 160:64:@40865.4]
  wire [13:0] _T_93307; // @[Modules.scala 160:64:@40866.4]
  wire [13:0] buffer_12_329; // @[Modules.scala 160:64:@40867.4]
  wire [14:0] _T_93309; // @[Modules.scala 160:64:@40869.4]
  wire [13:0] _T_93310; // @[Modules.scala 160:64:@40870.4]
  wire [13:0] buffer_12_330; // @[Modules.scala 160:64:@40871.4]
  wire [13:0] buffer_12_67; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93312; // @[Modules.scala 160:64:@40873.4]
  wire [13:0] _T_93313; // @[Modules.scala 160:64:@40874.4]
  wire [13:0] buffer_12_331; // @[Modules.scala 160:64:@40875.4]
  wire [13:0] buffer_12_70; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93318; // @[Modules.scala 160:64:@40881.4]
  wire [13:0] _T_93319; // @[Modules.scala 160:64:@40882.4]
  wire [13:0] buffer_12_333; // @[Modules.scala 160:64:@40883.4]
  wire [13:0] buffer_12_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93321; // @[Modules.scala 160:64:@40885.4]
  wire [13:0] _T_93322; // @[Modules.scala 160:64:@40886.4]
  wire [13:0] buffer_12_334; // @[Modules.scala 160:64:@40887.4]
  wire [13:0] buffer_12_74; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93324; // @[Modules.scala 160:64:@40889.4]
  wire [13:0] _T_93325; // @[Modules.scala 160:64:@40890.4]
  wire [13:0] buffer_12_335; // @[Modules.scala 160:64:@40891.4]
  wire [13:0] buffer_12_76; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93327; // @[Modules.scala 160:64:@40893.4]
  wire [13:0] _T_93328; // @[Modules.scala 160:64:@40894.4]
  wire [13:0] buffer_12_336; // @[Modules.scala 160:64:@40895.4]
  wire [13:0] buffer_12_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93333; // @[Modules.scala 160:64:@40901.4]
  wire [13:0] _T_93334; // @[Modules.scala 160:64:@40902.4]
  wire [13:0] buffer_12_338; // @[Modules.scala 160:64:@40903.4]
  wire [14:0] _T_93336; // @[Modules.scala 160:64:@40905.4]
  wire [13:0] _T_93337; // @[Modules.scala 160:64:@40906.4]
  wire [13:0] buffer_12_339; // @[Modules.scala 160:64:@40907.4]
  wire [14:0] _T_93339; // @[Modules.scala 160:64:@40909.4]
  wire [13:0] _T_93340; // @[Modules.scala 160:64:@40910.4]
  wire [13:0] buffer_12_340; // @[Modules.scala 160:64:@40911.4]
  wire [14:0] _T_93342; // @[Modules.scala 160:64:@40913.4]
  wire [13:0] _T_93343; // @[Modules.scala 160:64:@40914.4]
  wire [13:0] buffer_12_341; // @[Modules.scala 160:64:@40915.4]
  wire [13:0] buffer_12_88; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93345; // @[Modules.scala 160:64:@40917.4]
  wire [13:0] _T_93346; // @[Modules.scala 160:64:@40918.4]
  wire [13:0] buffer_12_342; // @[Modules.scala 160:64:@40919.4]
  wire [13:0] buffer_12_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93348; // @[Modules.scala 160:64:@40921.4]
  wire [13:0] _T_93349; // @[Modules.scala 160:64:@40922.4]
  wire [13:0] buffer_12_343; // @[Modules.scala 160:64:@40923.4]
  wire [13:0] buffer_12_92; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93351; // @[Modules.scala 160:64:@40925.4]
  wire [13:0] _T_93352; // @[Modules.scala 160:64:@40926.4]
  wire [13:0] buffer_12_344; // @[Modules.scala 160:64:@40927.4]
  wire [13:0] buffer_12_94; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93354; // @[Modules.scala 160:64:@40929.4]
  wire [13:0] _T_93355; // @[Modules.scala 160:64:@40930.4]
  wire [13:0] buffer_12_345; // @[Modules.scala 160:64:@40931.4]
  wire [14:0] _T_93357; // @[Modules.scala 160:64:@40933.4]
  wire [13:0] _T_93358; // @[Modules.scala 160:64:@40934.4]
  wire [13:0] buffer_12_346; // @[Modules.scala 160:64:@40935.4]
  wire [13:0] buffer_12_104; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93369; // @[Modules.scala 160:64:@40949.4]
  wire [13:0] _T_93370; // @[Modules.scala 160:64:@40950.4]
  wire [13:0] buffer_12_350; // @[Modules.scala 160:64:@40951.4]
  wire [13:0] buffer_12_106; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93372; // @[Modules.scala 160:64:@40953.4]
  wire [13:0] _T_93373; // @[Modules.scala 160:64:@40954.4]
  wire [13:0] buffer_12_351; // @[Modules.scala 160:64:@40955.4]
  wire [14:0] _T_93375; // @[Modules.scala 160:64:@40957.4]
  wire [13:0] _T_93376; // @[Modules.scala 160:64:@40958.4]
  wire [13:0] buffer_12_352; // @[Modules.scala 160:64:@40959.4]
  wire [13:0] buffer_12_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93387; // @[Modules.scala 160:64:@40973.4]
  wire [13:0] _T_93388; // @[Modules.scala 160:64:@40974.4]
  wire [13:0] buffer_12_356; // @[Modules.scala 160:64:@40975.4]
  wire [13:0] buffer_12_118; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93390; // @[Modules.scala 160:64:@40977.4]
  wire [13:0] _T_93391; // @[Modules.scala 160:64:@40978.4]
  wire [13:0] buffer_12_357; // @[Modules.scala 160:64:@40979.4]
  wire [13:0] buffer_12_122; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93396; // @[Modules.scala 160:64:@40985.4]
  wire [13:0] _T_93397; // @[Modules.scala 160:64:@40986.4]
  wire [13:0] buffer_12_359; // @[Modules.scala 160:64:@40987.4]
  wire [14:0] _T_93399; // @[Modules.scala 160:64:@40989.4]
  wire [13:0] _T_93400; // @[Modules.scala 160:64:@40990.4]
  wire [13:0] buffer_12_360; // @[Modules.scala 160:64:@40991.4]
  wire [13:0] buffer_12_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93402; // @[Modules.scala 160:64:@40993.4]
  wire [13:0] _T_93403; // @[Modules.scala 160:64:@40994.4]
  wire [13:0] buffer_12_361; // @[Modules.scala 160:64:@40995.4]
  wire [13:0] buffer_12_128; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93405; // @[Modules.scala 160:64:@40997.4]
  wire [13:0] _T_93406; // @[Modules.scala 160:64:@40998.4]
  wire [13:0] buffer_12_362; // @[Modules.scala 160:64:@40999.4]
  wire [13:0] buffer_12_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93408; // @[Modules.scala 160:64:@41001.4]
  wire [13:0] _T_93409; // @[Modules.scala 160:64:@41002.4]
  wire [13:0] buffer_12_363; // @[Modules.scala 160:64:@41003.4]
  wire [14:0] _T_93414; // @[Modules.scala 160:64:@41009.4]
  wire [13:0] _T_93415; // @[Modules.scala 160:64:@41010.4]
  wire [13:0] buffer_12_365; // @[Modules.scala 160:64:@41011.4]
  wire [14:0] _T_93417; // @[Modules.scala 160:64:@41013.4]
  wire [13:0] _T_93418; // @[Modules.scala 160:64:@41014.4]
  wire [13:0] buffer_12_366; // @[Modules.scala 160:64:@41015.4]
  wire [14:0] _T_93420; // @[Modules.scala 160:64:@41017.4]
  wire [13:0] _T_93421; // @[Modules.scala 160:64:@41018.4]
  wire [13:0] buffer_12_367; // @[Modules.scala 160:64:@41019.4]
  wire [14:0] _T_93426; // @[Modules.scala 160:64:@41025.4]
  wire [13:0] _T_93427; // @[Modules.scala 160:64:@41026.4]
  wire [13:0] buffer_12_369; // @[Modules.scala 160:64:@41027.4]
  wire [14:0] _T_93429; // @[Modules.scala 160:64:@41029.4]
  wire [13:0] _T_93430; // @[Modules.scala 160:64:@41030.4]
  wire [13:0] buffer_12_370; // @[Modules.scala 160:64:@41031.4]
  wire [14:0] _T_93432; // @[Modules.scala 160:64:@41033.4]
  wire [13:0] _T_93433; // @[Modules.scala 160:64:@41034.4]
  wire [13:0] buffer_12_371; // @[Modules.scala 160:64:@41035.4]
  wire [14:0] _T_93435; // @[Modules.scala 160:64:@41037.4]
  wire [13:0] _T_93436; // @[Modules.scala 160:64:@41038.4]
  wire [13:0] buffer_12_372; // @[Modules.scala 160:64:@41039.4]
  wire [13:0] buffer_12_150; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93438; // @[Modules.scala 160:64:@41041.4]
  wire [13:0] _T_93439; // @[Modules.scala 160:64:@41042.4]
  wire [13:0] buffer_12_373; // @[Modules.scala 160:64:@41043.4]
  wire [14:0] _T_93441; // @[Modules.scala 160:64:@41045.4]
  wire [13:0] _T_93442; // @[Modules.scala 160:64:@41046.4]
  wire [13:0] buffer_12_374; // @[Modules.scala 160:64:@41047.4]
  wire [14:0] _T_93444; // @[Modules.scala 160:64:@41049.4]
  wire [13:0] _T_93445; // @[Modules.scala 160:64:@41050.4]
  wire [13:0] buffer_12_375; // @[Modules.scala 160:64:@41051.4]
  wire [14:0] _T_93450; // @[Modules.scala 160:64:@41057.4]
  wire [13:0] _T_93451; // @[Modules.scala 160:64:@41058.4]
  wire [13:0] buffer_12_377; // @[Modules.scala 160:64:@41059.4]
  wire [13:0] buffer_12_160; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93453; // @[Modules.scala 160:64:@41061.4]
  wire [13:0] _T_93454; // @[Modules.scala 160:64:@41062.4]
  wire [13:0] buffer_12_378; // @[Modules.scala 160:64:@41063.4]
  wire [14:0] _T_93456; // @[Modules.scala 160:64:@41065.4]
  wire [13:0] _T_93457; // @[Modules.scala 160:64:@41066.4]
  wire [13:0] buffer_12_379; // @[Modules.scala 160:64:@41067.4]
  wire [14:0] _T_93459; // @[Modules.scala 160:64:@41069.4]
  wire [13:0] _T_93460; // @[Modules.scala 160:64:@41070.4]
  wire [13:0] buffer_12_380; // @[Modules.scala 160:64:@41071.4]
  wire [13:0] buffer_12_166; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93462; // @[Modules.scala 160:64:@41073.4]
  wire [13:0] _T_93463; // @[Modules.scala 160:64:@41074.4]
  wire [13:0] buffer_12_381; // @[Modules.scala 160:64:@41075.4]
  wire [14:0] _T_93465; // @[Modules.scala 160:64:@41077.4]
  wire [13:0] _T_93466; // @[Modules.scala 160:64:@41078.4]
  wire [13:0] buffer_12_382; // @[Modules.scala 160:64:@41079.4]
  wire [13:0] buffer_12_170; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93468; // @[Modules.scala 160:64:@41081.4]
  wire [13:0] _T_93469; // @[Modules.scala 160:64:@41082.4]
  wire [13:0] buffer_12_383; // @[Modules.scala 160:64:@41083.4]
  wire [13:0] buffer_12_172; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93471; // @[Modules.scala 160:64:@41085.4]
  wire [13:0] _T_93472; // @[Modules.scala 160:64:@41086.4]
  wire [13:0] buffer_12_384; // @[Modules.scala 160:64:@41087.4]
  wire [13:0] buffer_12_174; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93474; // @[Modules.scala 160:64:@41089.4]
  wire [13:0] _T_93475; // @[Modules.scala 160:64:@41090.4]
  wire [13:0] buffer_12_385; // @[Modules.scala 160:64:@41091.4]
  wire [14:0] _T_93477; // @[Modules.scala 160:64:@41093.4]
  wire [13:0] _T_93478; // @[Modules.scala 160:64:@41094.4]
  wire [13:0] buffer_12_386; // @[Modules.scala 160:64:@41095.4]
  wire [13:0] buffer_12_178; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93480; // @[Modules.scala 160:64:@41097.4]
  wire [13:0] _T_93481; // @[Modules.scala 160:64:@41098.4]
  wire [13:0] buffer_12_387; // @[Modules.scala 160:64:@41099.4]
  wire [14:0] _T_93483; // @[Modules.scala 160:64:@41101.4]
  wire [13:0] _T_93484; // @[Modules.scala 160:64:@41102.4]
  wire [13:0] buffer_12_388; // @[Modules.scala 160:64:@41103.4]
  wire [13:0] buffer_12_182; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93486; // @[Modules.scala 160:64:@41105.4]
  wire [13:0] _T_93487; // @[Modules.scala 160:64:@41106.4]
  wire [13:0] buffer_12_389; // @[Modules.scala 160:64:@41107.4]
  wire [14:0] _T_93489; // @[Modules.scala 160:64:@41109.4]
  wire [13:0] _T_93490; // @[Modules.scala 160:64:@41110.4]
  wire [13:0] buffer_12_390; // @[Modules.scala 160:64:@41111.4]
  wire [14:0] _T_93492; // @[Modules.scala 160:64:@41113.4]
  wire [13:0] _T_93493; // @[Modules.scala 160:64:@41114.4]
  wire [13:0] buffer_12_391; // @[Modules.scala 160:64:@41115.4]
  wire [14:0] _T_93495; // @[Modules.scala 160:64:@41117.4]
  wire [13:0] _T_93496; // @[Modules.scala 160:64:@41118.4]
  wire [13:0] buffer_12_392; // @[Modules.scala 160:64:@41119.4]
  wire [14:0] _T_93498; // @[Modules.scala 160:64:@41121.4]
  wire [13:0] _T_93499; // @[Modules.scala 160:64:@41122.4]
  wire [13:0] buffer_12_393; // @[Modules.scala 160:64:@41123.4]
  wire [14:0] _T_93504; // @[Modules.scala 160:64:@41129.4]
  wire [13:0] _T_93505; // @[Modules.scala 160:64:@41130.4]
  wire [13:0] buffer_12_395; // @[Modules.scala 160:64:@41131.4]
  wire [13:0] buffer_12_196; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93507; // @[Modules.scala 160:64:@41133.4]
  wire [13:0] _T_93508; // @[Modules.scala 160:64:@41134.4]
  wire [13:0] buffer_12_396; // @[Modules.scala 160:64:@41135.4]
  wire [14:0] _T_93510; // @[Modules.scala 160:64:@41137.4]
  wire [13:0] _T_93511; // @[Modules.scala 160:64:@41138.4]
  wire [13:0] buffer_12_397; // @[Modules.scala 160:64:@41139.4]
  wire [14:0] _T_93516; // @[Modules.scala 160:64:@41145.4]
  wire [13:0] _T_93517; // @[Modules.scala 160:64:@41146.4]
  wire [13:0] buffer_12_399; // @[Modules.scala 160:64:@41147.4]
  wire [14:0] _T_93519; // @[Modules.scala 160:64:@41149.4]
  wire [13:0] _T_93520; // @[Modules.scala 160:64:@41150.4]
  wire [13:0] buffer_12_400; // @[Modules.scala 160:64:@41151.4]
  wire [13:0] buffer_12_206; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_207; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93522; // @[Modules.scala 160:64:@41153.4]
  wire [13:0] _T_93523; // @[Modules.scala 160:64:@41154.4]
  wire [13:0] buffer_12_401; // @[Modules.scala 160:64:@41155.4]
  wire [13:0] buffer_12_208; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93525; // @[Modules.scala 160:64:@41157.4]
  wire [13:0] _T_93526; // @[Modules.scala 160:64:@41158.4]
  wire [13:0] buffer_12_402; // @[Modules.scala 160:64:@41159.4]
  wire [14:0] _T_93531; // @[Modules.scala 160:64:@41165.4]
  wire [13:0] _T_93532; // @[Modules.scala 160:64:@41166.4]
  wire [13:0] buffer_12_404; // @[Modules.scala 160:64:@41167.4]
  wire [13:0] buffer_12_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93534; // @[Modules.scala 160:64:@41169.4]
  wire [13:0] _T_93535; // @[Modules.scala 160:64:@41170.4]
  wire [13:0] buffer_12_405; // @[Modules.scala 160:64:@41171.4]
  wire [13:0] buffer_12_216; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93537; // @[Modules.scala 160:64:@41173.4]
  wire [13:0] _T_93538; // @[Modules.scala 160:64:@41174.4]
  wire [13:0] buffer_12_406; // @[Modules.scala 160:64:@41175.4]
  wire [13:0] buffer_12_220; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93543; // @[Modules.scala 160:64:@41181.4]
  wire [13:0] _T_93544; // @[Modules.scala 160:64:@41182.4]
  wire [13:0] buffer_12_408; // @[Modules.scala 160:64:@41183.4]
  wire [14:0] _T_93546; // @[Modules.scala 160:64:@41185.4]
  wire [13:0] _T_93547; // @[Modules.scala 160:64:@41186.4]
  wire [13:0] buffer_12_409; // @[Modules.scala 160:64:@41187.4]
  wire [13:0] buffer_12_227; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93552; // @[Modules.scala 160:64:@41193.4]
  wire [13:0] _T_93553; // @[Modules.scala 160:64:@41194.4]
  wire [13:0] buffer_12_411; // @[Modules.scala 160:64:@41195.4]
  wire [13:0] buffer_12_228; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93555; // @[Modules.scala 160:64:@41197.4]
  wire [13:0] _T_93556; // @[Modules.scala 160:64:@41198.4]
  wire [13:0] buffer_12_412; // @[Modules.scala 160:64:@41199.4]
  wire [13:0] buffer_12_230; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93558; // @[Modules.scala 160:64:@41201.4]
  wire [13:0] _T_93559; // @[Modules.scala 160:64:@41202.4]
  wire [13:0] buffer_12_413; // @[Modules.scala 160:64:@41203.4]
  wire [13:0] buffer_12_238; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93570; // @[Modules.scala 160:64:@41217.4]
  wire [13:0] _T_93571; // @[Modules.scala 160:64:@41218.4]
  wire [13:0] buffer_12_417; // @[Modules.scala 160:64:@41219.4]
  wire [13:0] buffer_12_240; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93573; // @[Modules.scala 160:64:@41221.4]
  wire [13:0] _T_93574; // @[Modules.scala 160:64:@41222.4]
  wire [13:0] buffer_12_418; // @[Modules.scala 160:64:@41223.4]
  wire [13:0] buffer_12_242; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93576; // @[Modules.scala 160:64:@41225.4]
  wire [13:0] _T_93577; // @[Modules.scala 160:64:@41226.4]
  wire [13:0] buffer_12_419; // @[Modules.scala 160:64:@41227.4]
  wire [13:0] buffer_12_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93579; // @[Modules.scala 160:64:@41229.4]
  wire [13:0] _T_93580; // @[Modules.scala 160:64:@41230.4]
  wire [13:0] buffer_12_420; // @[Modules.scala 160:64:@41231.4]
  wire [14:0] _T_93585; // @[Modules.scala 160:64:@41237.4]
  wire [13:0] _T_93586; // @[Modules.scala 160:64:@41238.4]
  wire [13:0] buffer_12_422; // @[Modules.scala 160:64:@41239.4]
  wire [13:0] buffer_12_251; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93588; // @[Modules.scala 160:64:@41241.4]
  wire [13:0] _T_93589; // @[Modules.scala 160:64:@41242.4]
  wire [13:0] buffer_12_423; // @[Modules.scala 160:64:@41243.4]
  wire [13:0] buffer_12_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93591; // @[Modules.scala 160:64:@41245.4]
  wire [13:0] _T_93592; // @[Modules.scala 160:64:@41246.4]
  wire [13:0] buffer_12_424; // @[Modules.scala 160:64:@41247.4]
  wire [13:0] buffer_12_254; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_12_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93594; // @[Modules.scala 160:64:@41249.4]
  wire [13:0] _T_93595; // @[Modules.scala 160:64:@41250.4]
  wire [13:0] buffer_12_425; // @[Modules.scala 160:64:@41251.4]
  wire [13:0] buffer_12_256; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93597; // @[Modules.scala 160:64:@41253.4]
  wire [13:0] _T_93598; // @[Modules.scala 160:64:@41254.4]
  wire [13:0] buffer_12_426; // @[Modules.scala 160:64:@41255.4]
  wire [13:0] buffer_12_261; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93603; // @[Modules.scala 160:64:@41261.4]
  wire [13:0] _T_93604; // @[Modules.scala 160:64:@41262.4]
  wire [13:0] buffer_12_428; // @[Modules.scala 160:64:@41263.4]
  wire [13:0] buffer_12_263; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93606; // @[Modules.scala 160:64:@41265.4]
  wire [13:0] _T_93607; // @[Modules.scala 160:64:@41266.4]
  wire [13:0] buffer_12_429; // @[Modules.scala 160:64:@41267.4]
  wire [14:0] _T_93609; // @[Modules.scala 160:64:@41269.4]
  wire [13:0] _T_93610; // @[Modules.scala 160:64:@41270.4]
  wire [13:0] buffer_12_430; // @[Modules.scala 160:64:@41271.4]
  wire [13:0] buffer_12_266; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93612; // @[Modules.scala 160:64:@41273.4]
  wire [13:0] _T_93613; // @[Modules.scala 160:64:@41274.4]
  wire [13:0] buffer_12_431; // @[Modules.scala 160:64:@41275.4]
  wire [13:0] buffer_12_268; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93615; // @[Modules.scala 160:64:@41277.4]
  wire [13:0] _T_93616; // @[Modules.scala 160:64:@41278.4]
  wire [13:0] buffer_12_432; // @[Modules.scala 160:64:@41279.4]
  wire [13:0] buffer_12_273; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93621; // @[Modules.scala 160:64:@41285.4]
  wire [13:0] _T_93622; // @[Modules.scala 160:64:@41286.4]
  wire [13:0] buffer_12_434; // @[Modules.scala 160:64:@41287.4]
  wire [14:0] _T_93624; // @[Modules.scala 160:64:@41289.4]
  wire [13:0] _T_93625; // @[Modules.scala 160:64:@41290.4]
  wire [13:0] buffer_12_435; // @[Modules.scala 160:64:@41291.4]
  wire [13:0] buffer_12_276; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93627; // @[Modules.scala 160:64:@41293.4]
  wire [13:0] _T_93628; // @[Modules.scala 160:64:@41294.4]
  wire [13:0] buffer_12_436; // @[Modules.scala 160:64:@41295.4]
  wire [13:0] buffer_12_278; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93630; // @[Modules.scala 160:64:@41297.4]
  wire [13:0] _T_93631; // @[Modules.scala 160:64:@41298.4]
  wire [13:0] buffer_12_437; // @[Modules.scala 160:64:@41299.4]
  wire [13:0] buffer_12_280; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93633; // @[Modules.scala 160:64:@41301.4]
  wire [13:0] _T_93634; // @[Modules.scala 160:64:@41302.4]
  wire [13:0] buffer_12_438; // @[Modules.scala 160:64:@41303.4]
  wire [13:0] buffer_12_289; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93645; // @[Modules.scala 160:64:@41317.4]
  wire [13:0] _T_93646; // @[Modules.scala 160:64:@41318.4]
  wire [13:0] buffer_12_442; // @[Modules.scala 160:64:@41319.4]
  wire [14:0] _T_93648; // @[Modules.scala 160:64:@41321.4]
  wire [13:0] _T_93649; // @[Modules.scala 160:64:@41322.4]
  wire [13:0] buffer_12_443; // @[Modules.scala 160:64:@41323.4]
  wire [13:0] buffer_12_296; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_93657; // @[Modules.scala 160:64:@41333.4]
  wire [13:0] _T_93658; // @[Modules.scala 160:64:@41334.4]
  wire [13:0] buffer_12_446; // @[Modules.scala 160:64:@41335.4]
  wire [14:0] _T_93660; // @[Modules.scala 166:64:@41337.4]
  wire [13:0] _T_93661; // @[Modules.scala 166:64:@41338.4]
  wire [13:0] buffer_12_447; // @[Modules.scala 166:64:@41339.4]
  wire [14:0] _T_93663; // @[Modules.scala 166:64:@41341.4]
  wire [13:0] _T_93664; // @[Modules.scala 166:64:@41342.4]
  wire [13:0] buffer_12_448; // @[Modules.scala 166:64:@41343.4]
  wire [14:0] _T_93666; // @[Modules.scala 166:64:@41345.4]
  wire [13:0] _T_93667; // @[Modules.scala 166:64:@41346.4]
  wire [13:0] buffer_12_449; // @[Modules.scala 166:64:@41347.4]
  wire [14:0] _T_93669; // @[Modules.scala 166:64:@41349.4]
  wire [13:0] _T_93670; // @[Modules.scala 166:64:@41350.4]
  wire [13:0] buffer_12_450; // @[Modules.scala 166:64:@41351.4]
  wire [14:0] _T_93672; // @[Modules.scala 166:64:@41353.4]
  wire [13:0] _T_93673; // @[Modules.scala 166:64:@41354.4]
  wire [13:0] buffer_12_451; // @[Modules.scala 166:64:@41355.4]
  wire [14:0] _T_93675; // @[Modules.scala 166:64:@41357.4]
  wire [13:0] _T_93676; // @[Modules.scala 166:64:@41358.4]
  wire [13:0] buffer_12_452; // @[Modules.scala 166:64:@41359.4]
  wire [14:0] _T_93678; // @[Modules.scala 166:64:@41361.4]
  wire [13:0] _T_93679; // @[Modules.scala 166:64:@41362.4]
  wire [13:0] buffer_12_453; // @[Modules.scala 166:64:@41363.4]
  wire [14:0] _T_93681; // @[Modules.scala 166:64:@41365.4]
  wire [13:0] _T_93682; // @[Modules.scala 166:64:@41366.4]
  wire [13:0] buffer_12_454; // @[Modules.scala 166:64:@41367.4]
  wire [14:0] _T_93684; // @[Modules.scala 166:64:@41369.4]
  wire [13:0] _T_93685; // @[Modules.scala 166:64:@41370.4]
  wire [13:0] buffer_12_455; // @[Modules.scala 166:64:@41371.4]
  wire [14:0] _T_93687; // @[Modules.scala 166:64:@41373.4]
  wire [13:0] _T_93688; // @[Modules.scala 166:64:@41374.4]
  wire [13:0] buffer_12_456; // @[Modules.scala 166:64:@41375.4]
  wire [14:0] _T_93690; // @[Modules.scala 166:64:@41377.4]
  wire [13:0] _T_93691; // @[Modules.scala 166:64:@41378.4]
  wire [13:0] buffer_12_457; // @[Modules.scala 166:64:@41379.4]
  wire [14:0] _T_93693; // @[Modules.scala 166:64:@41381.4]
  wire [13:0] _T_93694; // @[Modules.scala 166:64:@41382.4]
  wire [13:0] buffer_12_458; // @[Modules.scala 166:64:@41383.4]
  wire [14:0] _T_93696; // @[Modules.scala 166:64:@41385.4]
  wire [13:0] _T_93697; // @[Modules.scala 166:64:@41386.4]
  wire [13:0] buffer_12_459; // @[Modules.scala 166:64:@41387.4]
  wire [14:0] _T_93699; // @[Modules.scala 166:64:@41389.4]
  wire [13:0] _T_93700; // @[Modules.scala 166:64:@41390.4]
  wire [13:0] buffer_12_460; // @[Modules.scala 166:64:@41391.4]
  wire [14:0] _T_93702; // @[Modules.scala 166:64:@41393.4]
  wire [13:0] _T_93703; // @[Modules.scala 166:64:@41394.4]
  wire [13:0] buffer_12_461; // @[Modules.scala 166:64:@41395.4]
  wire [14:0] _T_93705; // @[Modules.scala 166:64:@41397.4]
  wire [13:0] _T_93706; // @[Modules.scala 166:64:@41398.4]
  wire [13:0] buffer_12_462; // @[Modules.scala 166:64:@41399.4]
  wire [14:0] _T_93708; // @[Modules.scala 166:64:@41401.4]
  wire [13:0] _T_93709; // @[Modules.scala 166:64:@41402.4]
  wire [13:0] buffer_12_463; // @[Modules.scala 166:64:@41403.4]
  wire [14:0] _T_93711; // @[Modules.scala 166:64:@41405.4]
  wire [13:0] _T_93712; // @[Modules.scala 166:64:@41406.4]
  wire [13:0] buffer_12_464; // @[Modules.scala 166:64:@41407.4]
  wire [14:0] _T_93714; // @[Modules.scala 166:64:@41409.4]
  wire [13:0] _T_93715; // @[Modules.scala 166:64:@41410.4]
  wire [13:0] buffer_12_465; // @[Modules.scala 166:64:@41411.4]
  wire [14:0] _T_93717; // @[Modules.scala 166:64:@41413.4]
  wire [13:0] _T_93718; // @[Modules.scala 166:64:@41414.4]
  wire [13:0] buffer_12_466; // @[Modules.scala 166:64:@41415.4]
  wire [14:0] _T_93720; // @[Modules.scala 166:64:@41417.4]
  wire [13:0] _T_93721; // @[Modules.scala 166:64:@41418.4]
  wire [13:0] buffer_12_467; // @[Modules.scala 166:64:@41419.4]
  wire [14:0] _T_93723; // @[Modules.scala 166:64:@41421.4]
  wire [13:0] _T_93724; // @[Modules.scala 166:64:@41422.4]
  wire [13:0] buffer_12_468; // @[Modules.scala 166:64:@41423.4]
  wire [14:0] _T_93726; // @[Modules.scala 166:64:@41425.4]
  wire [13:0] _T_93727; // @[Modules.scala 166:64:@41426.4]
  wire [13:0] buffer_12_469; // @[Modules.scala 166:64:@41427.4]
  wire [14:0] _T_93729; // @[Modules.scala 166:64:@41429.4]
  wire [13:0] _T_93730; // @[Modules.scala 166:64:@41430.4]
  wire [13:0] buffer_12_470; // @[Modules.scala 166:64:@41431.4]
  wire [14:0] _T_93732; // @[Modules.scala 166:64:@41433.4]
  wire [13:0] _T_93733; // @[Modules.scala 166:64:@41434.4]
  wire [13:0] buffer_12_471; // @[Modules.scala 166:64:@41435.4]
  wire [14:0] _T_93738; // @[Modules.scala 166:64:@41441.4]
  wire [13:0] _T_93739; // @[Modules.scala 166:64:@41442.4]
  wire [13:0] buffer_12_473; // @[Modules.scala 166:64:@41443.4]
  wire [14:0] _T_93741; // @[Modules.scala 166:64:@41445.4]
  wire [13:0] _T_93742; // @[Modules.scala 166:64:@41446.4]
  wire [13:0] buffer_12_474; // @[Modules.scala 166:64:@41447.4]
  wire [14:0] _T_93744; // @[Modules.scala 166:64:@41449.4]
  wire [13:0] _T_93745; // @[Modules.scala 166:64:@41450.4]
  wire [13:0] buffer_12_475; // @[Modules.scala 166:64:@41451.4]
  wire [14:0] _T_93747; // @[Modules.scala 166:64:@41453.4]
  wire [13:0] _T_93748; // @[Modules.scala 166:64:@41454.4]
  wire [13:0] buffer_12_476; // @[Modules.scala 166:64:@41455.4]
  wire [14:0] _T_93750; // @[Modules.scala 166:64:@41457.4]
  wire [13:0] _T_93751; // @[Modules.scala 166:64:@41458.4]
  wire [13:0] buffer_12_477; // @[Modules.scala 166:64:@41459.4]
  wire [14:0] _T_93753; // @[Modules.scala 166:64:@41461.4]
  wire [13:0] _T_93754; // @[Modules.scala 166:64:@41462.4]
  wire [13:0] buffer_12_478; // @[Modules.scala 166:64:@41463.4]
  wire [14:0] _T_93756; // @[Modules.scala 166:64:@41465.4]
  wire [13:0] _T_93757; // @[Modules.scala 166:64:@41466.4]
  wire [13:0] buffer_12_479; // @[Modules.scala 166:64:@41467.4]
  wire [14:0] _T_93759; // @[Modules.scala 166:64:@41469.4]
  wire [13:0] _T_93760; // @[Modules.scala 166:64:@41470.4]
  wire [13:0] buffer_12_480; // @[Modules.scala 166:64:@41471.4]
  wire [14:0] _T_93762; // @[Modules.scala 166:64:@41473.4]
  wire [13:0] _T_93763; // @[Modules.scala 166:64:@41474.4]
  wire [13:0] buffer_12_481; // @[Modules.scala 166:64:@41475.4]
  wire [14:0] _T_93765; // @[Modules.scala 166:64:@41477.4]
  wire [13:0] _T_93766; // @[Modules.scala 166:64:@41478.4]
  wire [13:0] buffer_12_482; // @[Modules.scala 166:64:@41479.4]
  wire [14:0] _T_93768; // @[Modules.scala 166:64:@41481.4]
  wire [13:0] _T_93769; // @[Modules.scala 166:64:@41482.4]
  wire [13:0] buffer_12_483; // @[Modules.scala 166:64:@41483.4]
  wire [14:0] _T_93771; // @[Modules.scala 166:64:@41485.4]
  wire [13:0] _T_93772; // @[Modules.scala 166:64:@41486.4]
  wire [13:0] buffer_12_484; // @[Modules.scala 166:64:@41487.4]
  wire [14:0] _T_93774; // @[Modules.scala 166:64:@41489.4]
  wire [13:0] _T_93775; // @[Modules.scala 166:64:@41490.4]
  wire [13:0] buffer_12_485; // @[Modules.scala 166:64:@41491.4]
  wire [14:0] _T_93777; // @[Modules.scala 166:64:@41493.4]
  wire [13:0] _T_93778; // @[Modules.scala 166:64:@41494.4]
  wire [13:0] buffer_12_486; // @[Modules.scala 166:64:@41495.4]
  wire [14:0] _T_93780; // @[Modules.scala 166:64:@41497.4]
  wire [13:0] _T_93781; // @[Modules.scala 166:64:@41498.4]
  wire [13:0] buffer_12_487; // @[Modules.scala 166:64:@41499.4]
  wire [14:0] _T_93783; // @[Modules.scala 166:64:@41501.4]
  wire [13:0] _T_93784; // @[Modules.scala 166:64:@41502.4]
  wire [13:0] buffer_12_488; // @[Modules.scala 166:64:@41503.4]
  wire [14:0] _T_93786; // @[Modules.scala 166:64:@41505.4]
  wire [13:0] _T_93787; // @[Modules.scala 166:64:@41506.4]
  wire [13:0] buffer_12_489; // @[Modules.scala 166:64:@41507.4]
  wire [14:0] _T_93789; // @[Modules.scala 166:64:@41509.4]
  wire [13:0] _T_93790; // @[Modules.scala 166:64:@41510.4]
  wire [13:0] buffer_12_490; // @[Modules.scala 166:64:@41511.4]
  wire [14:0] _T_93792; // @[Modules.scala 166:64:@41513.4]
  wire [13:0] _T_93793; // @[Modules.scala 166:64:@41514.4]
  wire [13:0] buffer_12_491; // @[Modules.scala 166:64:@41515.4]
  wire [14:0] _T_93795; // @[Modules.scala 166:64:@41517.4]
  wire [13:0] _T_93796; // @[Modules.scala 166:64:@41518.4]
  wire [13:0] buffer_12_492; // @[Modules.scala 166:64:@41519.4]
  wire [14:0] _T_93798; // @[Modules.scala 166:64:@41521.4]
  wire [13:0] _T_93799; // @[Modules.scala 166:64:@41522.4]
  wire [13:0] buffer_12_493; // @[Modules.scala 166:64:@41523.4]
  wire [14:0] _T_93801; // @[Modules.scala 166:64:@41525.4]
  wire [13:0] _T_93802; // @[Modules.scala 166:64:@41526.4]
  wire [13:0] buffer_12_494; // @[Modules.scala 166:64:@41527.4]
  wire [14:0] _T_93804; // @[Modules.scala 166:64:@41529.4]
  wire [13:0] _T_93805; // @[Modules.scala 166:64:@41530.4]
  wire [13:0] buffer_12_495; // @[Modules.scala 166:64:@41531.4]
  wire [14:0] _T_93807; // @[Modules.scala 166:64:@41533.4]
  wire [13:0] _T_93808; // @[Modules.scala 166:64:@41534.4]
  wire [13:0] buffer_12_496; // @[Modules.scala 166:64:@41535.4]
  wire [14:0] _T_93810; // @[Modules.scala 166:64:@41537.4]
  wire [13:0] _T_93811; // @[Modules.scala 166:64:@41538.4]
  wire [13:0] buffer_12_497; // @[Modules.scala 166:64:@41539.4]
  wire [14:0] _T_93813; // @[Modules.scala 166:64:@41541.4]
  wire [13:0] _T_93814; // @[Modules.scala 166:64:@41542.4]
  wire [13:0] buffer_12_498; // @[Modules.scala 166:64:@41543.4]
  wire [14:0] _T_93816; // @[Modules.scala 166:64:@41545.4]
  wire [13:0] _T_93817; // @[Modules.scala 166:64:@41546.4]
  wire [13:0] buffer_12_499; // @[Modules.scala 166:64:@41547.4]
  wire [14:0] _T_93819; // @[Modules.scala 166:64:@41549.4]
  wire [13:0] _T_93820; // @[Modules.scala 166:64:@41550.4]
  wire [13:0] buffer_12_500; // @[Modules.scala 166:64:@41551.4]
  wire [14:0] _T_93822; // @[Modules.scala 166:64:@41553.4]
  wire [13:0] _T_93823; // @[Modules.scala 166:64:@41554.4]
  wire [13:0] buffer_12_501; // @[Modules.scala 166:64:@41555.4]
  wire [14:0] _T_93825; // @[Modules.scala 166:64:@41557.4]
  wire [13:0] _T_93826; // @[Modules.scala 166:64:@41558.4]
  wire [13:0] buffer_12_502; // @[Modules.scala 166:64:@41559.4]
  wire [14:0] _T_93828; // @[Modules.scala 166:64:@41561.4]
  wire [13:0] _T_93829; // @[Modules.scala 166:64:@41562.4]
  wire [13:0] buffer_12_503; // @[Modules.scala 166:64:@41563.4]
  wire [14:0] _T_93831; // @[Modules.scala 166:64:@41565.4]
  wire [13:0] _T_93832; // @[Modules.scala 166:64:@41566.4]
  wire [13:0] buffer_12_504; // @[Modules.scala 166:64:@41567.4]
  wire [14:0] _T_93837; // @[Modules.scala 166:64:@41573.4]
  wire [13:0] _T_93838; // @[Modules.scala 166:64:@41574.4]
  wire [13:0] buffer_12_506; // @[Modules.scala 166:64:@41575.4]
  wire [14:0] _T_93840; // @[Modules.scala 166:64:@41577.4]
  wire [13:0] _T_93841; // @[Modules.scala 166:64:@41578.4]
  wire [13:0] buffer_12_507; // @[Modules.scala 166:64:@41579.4]
  wire [14:0] _T_93843; // @[Modules.scala 166:64:@41581.4]
  wire [13:0] _T_93844; // @[Modules.scala 166:64:@41582.4]
  wire [13:0] buffer_12_508; // @[Modules.scala 166:64:@41583.4]
  wire [14:0] _T_93846; // @[Modules.scala 166:64:@41585.4]
  wire [13:0] _T_93847; // @[Modules.scala 166:64:@41586.4]
  wire [13:0] buffer_12_509; // @[Modules.scala 166:64:@41587.4]
  wire [14:0] _T_93849; // @[Modules.scala 166:64:@41589.4]
  wire [13:0] _T_93850; // @[Modules.scala 166:64:@41590.4]
  wire [13:0] buffer_12_510; // @[Modules.scala 166:64:@41591.4]
  wire [14:0] _T_93852; // @[Modules.scala 166:64:@41593.4]
  wire [13:0] _T_93853; // @[Modules.scala 166:64:@41594.4]
  wire [13:0] buffer_12_511; // @[Modules.scala 166:64:@41595.4]
  wire [14:0] _T_93855; // @[Modules.scala 166:64:@41597.4]
  wire [13:0] _T_93856; // @[Modules.scala 166:64:@41598.4]
  wire [13:0] buffer_12_512; // @[Modules.scala 166:64:@41599.4]
  wire [14:0] _T_93858; // @[Modules.scala 166:64:@41601.4]
  wire [13:0] _T_93859; // @[Modules.scala 166:64:@41602.4]
  wire [13:0] buffer_12_513; // @[Modules.scala 166:64:@41603.4]
  wire [14:0] _T_93861; // @[Modules.scala 166:64:@41605.4]
  wire [13:0] _T_93862; // @[Modules.scala 166:64:@41606.4]
  wire [13:0] buffer_12_514; // @[Modules.scala 166:64:@41607.4]
  wire [14:0] _T_93864; // @[Modules.scala 166:64:@41609.4]
  wire [13:0] _T_93865; // @[Modules.scala 166:64:@41610.4]
  wire [13:0] buffer_12_515; // @[Modules.scala 166:64:@41611.4]
  wire [14:0] _T_93867; // @[Modules.scala 166:64:@41613.4]
  wire [13:0] _T_93868; // @[Modules.scala 166:64:@41614.4]
  wire [13:0] buffer_12_516; // @[Modules.scala 166:64:@41615.4]
  wire [14:0] _T_93870; // @[Modules.scala 166:64:@41617.4]
  wire [13:0] _T_93871; // @[Modules.scala 166:64:@41618.4]
  wire [13:0] buffer_12_517; // @[Modules.scala 166:64:@41619.4]
  wire [14:0] _T_93873; // @[Modules.scala 166:64:@41621.4]
  wire [13:0] _T_93874; // @[Modules.scala 166:64:@41622.4]
  wire [13:0] buffer_12_518; // @[Modules.scala 166:64:@41623.4]
  wire [14:0] _T_93876; // @[Modules.scala 166:64:@41625.4]
  wire [13:0] _T_93877; // @[Modules.scala 166:64:@41626.4]
  wire [13:0] buffer_12_519; // @[Modules.scala 166:64:@41627.4]
  wire [14:0] _T_93882; // @[Modules.scala 160:64:@41633.4]
  wire [13:0] _T_93883; // @[Modules.scala 160:64:@41634.4]
  wire [13:0] buffer_12_521; // @[Modules.scala 160:64:@41635.4]
  wire [14:0] _T_93885; // @[Modules.scala 160:64:@41637.4]
  wire [13:0] _T_93886; // @[Modules.scala 160:64:@41638.4]
  wire [13:0] buffer_12_522; // @[Modules.scala 160:64:@41639.4]
  wire [14:0] _T_93888; // @[Modules.scala 160:64:@41641.4]
  wire [13:0] _T_93889; // @[Modules.scala 160:64:@41642.4]
  wire [13:0] buffer_12_523; // @[Modules.scala 160:64:@41643.4]
  wire [14:0] _T_93891; // @[Modules.scala 160:64:@41645.4]
  wire [13:0] _T_93892; // @[Modules.scala 160:64:@41646.4]
  wire [13:0] buffer_12_524; // @[Modules.scala 160:64:@41647.4]
  wire [14:0] _T_93894; // @[Modules.scala 160:64:@41649.4]
  wire [13:0] _T_93895; // @[Modules.scala 160:64:@41650.4]
  wire [13:0] buffer_12_525; // @[Modules.scala 160:64:@41651.4]
  wire [14:0] _T_93897; // @[Modules.scala 160:64:@41653.4]
  wire [13:0] _T_93898; // @[Modules.scala 160:64:@41654.4]
  wire [13:0] buffer_12_526; // @[Modules.scala 160:64:@41655.4]
  wire [14:0] _T_93900; // @[Modules.scala 160:64:@41657.4]
  wire [13:0] _T_93901; // @[Modules.scala 160:64:@41658.4]
  wire [13:0] buffer_12_527; // @[Modules.scala 160:64:@41659.4]
  wire [14:0] _T_93903; // @[Modules.scala 160:64:@41661.4]
  wire [13:0] _T_93904; // @[Modules.scala 160:64:@41662.4]
  wire [13:0] buffer_12_528; // @[Modules.scala 160:64:@41663.4]
  wire [14:0] _T_93906; // @[Modules.scala 160:64:@41665.4]
  wire [13:0] _T_93907; // @[Modules.scala 160:64:@41666.4]
  wire [13:0] buffer_12_529; // @[Modules.scala 160:64:@41667.4]
  wire [14:0] _T_93909; // @[Modules.scala 160:64:@41669.4]
  wire [13:0] _T_93910; // @[Modules.scala 160:64:@41670.4]
  wire [13:0] buffer_12_530; // @[Modules.scala 160:64:@41671.4]
  wire [14:0] _T_93912; // @[Modules.scala 160:64:@41673.4]
  wire [13:0] _T_93913; // @[Modules.scala 160:64:@41674.4]
  wire [13:0] buffer_12_531; // @[Modules.scala 160:64:@41675.4]
  wire [14:0] _T_93915; // @[Modules.scala 160:64:@41677.4]
  wire [13:0] _T_93916; // @[Modules.scala 160:64:@41678.4]
  wire [13:0] buffer_12_532; // @[Modules.scala 160:64:@41679.4]
  wire [14:0] _T_93918; // @[Modules.scala 160:64:@41681.4]
  wire [13:0] _T_93919; // @[Modules.scala 160:64:@41682.4]
  wire [13:0] buffer_12_533; // @[Modules.scala 160:64:@41683.4]
  wire [14:0] _T_93921; // @[Modules.scala 160:64:@41685.4]
  wire [13:0] _T_93922; // @[Modules.scala 160:64:@41686.4]
  wire [13:0] buffer_12_534; // @[Modules.scala 160:64:@41687.4]
  wire [14:0] _T_93924; // @[Modules.scala 160:64:@41689.4]
  wire [13:0] _T_93925; // @[Modules.scala 160:64:@41690.4]
  wire [13:0] buffer_12_535; // @[Modules.scala 160:64:@41691.4]
  wire [14:0] _T_93927; // @[Modules.scala 160:64:@41693.4]
  wire [13:0] _T_93928; // @[Modules.scala 160:64:@41694.4]
  wire [13:0] buffer_12_536; // @[Modules.scala 160:64:@41695.4]
  wire [14:0] _T_93930; // @[Modules.scala 160:64:@41697.4]
  wire [13:0] _T_93931; // @[Modules.scala 160:64:@41698.4]
  wire [13:0] buffer_12_537; // @[Modules.scala 160:64:@41699.4]
  wire [14:0] _T_93933; // @[Modules.scala 160:64:@41701.4]
  wire [13:0] _T_93934; // @[Modules.scala 160:64:@41702.4]
  wire [13:0] buffer_12_538; // @[Modules.scala 160:64:@41703.4]
  wire [14:0] _T_93936; // @[Modules.scala 160:64:@41705.4]
  wire [13:0] _T_93937; // @[Modules.scala 160:64:@41706.4]
  wire [13:0] buffer_12_539; // @[Modules.scala 160:64:@41707.4]
  wire [14:0] _T_93939; // @[Modules.scala 160:64:@41709.4]
  wire [13:0] _T_93940; // @[Modules.scala 160:64:@41710.4]
  wire [13:0] buffer_12_540; // @[Modules.scala 160:64:@41711.4]
  wire [14:0] _T_93942; // @[Modules.scala 160:64:@41713.4]
  wire [13:0] _T_93943; // @[Modules.scala 160:64:@41714.4]
  wire [13:0] buffer_12_541; // @[Modules.scala 160:64:@41715.4]
  wire [14:0] _T_93945; // @[Modules.scala 160:64:@41717.4]
  wire [13:0] _T_93946; // @[Modules.scala 160:64:@41718.4]
  wire [13:0] buffer_12_542; // @[Modules.scala 160:64:@41719.4]
  wire [14:0] _T_93948; // @[Modules.scala 160:64:@41721.4]
  wire [13:0] _T_93949; // @[Modules.scala 160:64:@41722.4]
  wire [13:0] buffer_12_543; // @[Modules.scala 160:64:@41723.4]
  wire [14:0] _T_93951; // @[Modules.scala 160:64:@41725.4]
  wire [13:0] _T_93952; // @[Modules.scala 160:64:@41726.4]
  wire [13:0] buffer_12_544; // @[Modules.scala 160:64:@41727.4]
  wire [14:0] _T_93954; // @[Modules.scala 160:64:@41729.4]
  wire [13:0] _T_93955; // @[Modules.scala 160:64:@41730.4]
  wire [13:0] buffer_12_545; // @[Modules.scala 160:64:@41731.4]
  wire [14:0] _T_93957; // @[Modules.scala 160:64:@41733.4]
  wire [13:0] _T_93958; // @[Modules.scala 160:64:@41734.4]
  wire [13:0] buffer_12_546; // @[Modules.scala 160:64:@41735.4]
  wire [14:0] _T_93960; // @[Modules.scala 160:64:@41737.4]
  wire [13:0] _T_93961; // @[Modules.scala 160:64:@41738.4]
  wire [13:0] buffer_12_547; // @[Modules.scala 160:64:@41739.4]
  wire [14:0] _T_93963; // @[Modules.scala 160:64:@41741.4]
  wire [13:0] _T_93964; // @[Modules.scala 160:64:@41742.4]
  wire [13:0] buffer_12_548; // @[Modules.scala 160:64:@41743.4]
  wire [14:0] _T_93966; // @[Modules.scala 160:64:@41745.4]
  wire [13:0] _T_93967; // @[Modules.scala 160:64:@41746.4]
  wire [13:0] buffer_12_549; // @[Modules.scala 160:64:@41747.4]
  wire [14:0] _T_93969; // @[Modules.scala 160:64:@41749.4]
  wire [13:0] _T_93970; // @[Modules.scala 160:64:@41750.4]
  wire [13:0] buffer_12_550; // @[Modules.scala 160:64:@41751.4]
  wire [14:0] _T_93972; // @[Modules.scala 160:64:@41753.4]
  wire [13:0] _T_93973; // @[Modules.scala 160:64:@41754.4]
  wire [13:0] buffer_12_551; // @[Modules.scala 160:64:@41755.4]
  wire [14:0] _T_93975; // @[Modules.scala 160:64:@41757.4]
  wire [13:0] _T_93976; // @[Modules.scala 160:64:@41758.4]
  wire [13:0] buffer_12_552; // @[Modules.scala 160:64:@41759.4]
  wire [14:0] _T_93978; // @[Modules.scala 160:64:@41761.4]
  wire [13:0] _T_93979; // @[Modules.scala 160:64:@41762.4]
  wire [13:0] buffer_12_553; // @[Modules.scala 160:64:@41763.4]
  wire [14:0] _T_93981; // @[Modules.scala 160:64:@41765.4]
  wire [13:0] _T_93982; // @[Modules.scala 160:64:@41766.4]
  wire [13:0] buffer_12_554; // @[Modules.scala 160:64:@41767.4]
  wire [14:0] _T_93984; // @[Modules.scala 160:64:@41769.4]
  wire [13:0] _T_93985; // @[Modules.scala 160:64:@41770.4]
  wire [13:0] buffer_12_555; // @[Modules.scala 160:64:@41771.4]
  wire [14:0] _T_93987; // @[Modules.scala 160:64:@41773.4]
  wire [13:0] _T_93988; // @[Modules.scala 160:64:@41774.4]
  wire [13:0] buffer_12_556; // @[Modules.scala 160:64:@41775.4]
  wire [14:0] _T_93990; // @[Modules.scala 160:64:@41777.4]
  wire [13:0] _T_93991; // @[Modules.scala 160:64:@41778.4]
  wire [13:0] buffer_12_557; // @[Modules.scala 160:64:@41779.4]
  wire [14:0] _T_93993; // @[Modules.scala 166:64:@41781.4]
  wire [13:0] _T_93994; // @[Modules.scala 166:64:@41782.4]
  wire [13:0] buffer_12_558; // @[Modules.scala 166:64:@41783.4]
  wire [14:0] _T_93996; // @[Modules.scala 166:64:@41785.4]
  wire [13:0] _T_93997; // @[Modules.scala 166:64:@41786.4]
  wire [13:0] buffer_12_559; // @[Modules.scala 166:64:@41787.4]
  wire [14:0] _T_93999; // @[Modules.scala 166:64:@41789.4]
  wire [13:0] _T_94000; // @[Modules.scala 166:64:@41790.4]
  wire [13:0] buffer_12_560; // @[Modules.scala 166:64:@41791.4]
  wire [14:0] _T_94002; // @[Modules.scala 166:64:@41793.4]
  wire [13:0] _T_94003; // @[Modules.scala 166:64:@41794.4]
  wire [13:0] buffer_12_561; // @[Modules.scala 166:64:@41795.4]
  wire [14:0] _T_94005; // @[Modules.scala 166:64:@41797.4]
  wire [13:0] _T_94006; // @[Modules.scala 166:64:@41798.4]
  wire [13:0] buffer_12_562; // @[Modules.scala 166:64:@41799.4]
  wire [14:0] _T_94008; // @[Modules.scala 166:64:@41801.4]
  wire [13:0] _T_94009; // @[Modules.scala 166:64:@41802.4]
  wire [13:0] buffer_12_563; // @[Modules.scala 166:64:@41803.4]
  wire [14:0] _T_94011; // @[Modules.scala 166:64:@41805.4]
  wire [13:0] _T_94012; // @[Modules.scala 166:64:@41806.4]
  wire [13:0] buffer_12_564; // @[Modules.scala 166:64:@41807.4]
  wire [14:0] _T_94014; // @[Modules.scala 166:64:@41809.4]
  wire [13:0] _T_94015; // @[Modules.scala 166:64:@41810.4]
  wire [13:0] buffer_12_565; // @[Modules.scala 166:64:@41811.4]
  wire [14:0] _T_94017; // @[Modules.scala 166:64:@41813.4]
  wire [13:0] _T_94018; // @[Modules.scala 166:64:@41814.4]
  wire [13:0] buffer_12_566; // @[Modules.scala 166:64:@41815.4]
  wire [14:0] _T_94020; // @[Modules.scala 166:64:@41817.4]
  wire [13:0] _T_94021; // @[Modules.scala 166:64:@41818.4]
  wire [13:0] buffer_12_567; // @[Modules.scala 166:64:@41819.4]
  wire [14:0] _T_94023; // @[Modules.scala 166:64:@41821.4]
  wire [13:0] _T_94024; // @[Modules.scala 166:64:@41822.4]
  wire [13:0] buffer_12_568; // @[Modules.scala 166:64:@41823.4]
  wire [14:0] _T_94026; // @[Modules.scala 166:64:@41825.4]
  wire [13:0] _T_94027; // @[Modules.scala 166:64:@41826.4]
  wire [13:0] buffer_12_569; // @[Modules.scala 166:64:@41827.4]
  wire [14:0] _T_94029; // @[Modules.scala 166:64:@41829.4]
  wire [13:0] _T_94030; // @[Modules.scala 166:64:@41830.4]
  wire [13:0] buffer_12_570; // @[Modules.scala 166:64:@41831.4]
  wire [14:0] _T_94032; // @[Modules.scala 166:64:@41833.4]
  wire [13:0] _T_94033; // @[Modules.scala 166:64:@41834.4]
  wire [13:0] buffer_12_571; // @[Modules.scala 166:64:@41835.4]
  wire [14:0] _T_94035; // @[Modules.scala 166:64:@41837.4]
  wire [13:0] _T_94036; // @[Modules.scala 166:64:@41838.4]
  wire [13:0] buffer_12_572; // @[Modules.scala 166:64:@41839.4]
  wire [14:0] _T_94038; // @[Modules.scala 166:64:@41841.4]
  wire [13:0] _T_94039; // @[Modules.scala 166:64:@41842.4]
  wire [13:0] buffer_12_573; // @[Modules.scala 166:64:@41843.4]
  wire [14:0] _T_94041; // @[Modules.scala 166:64:@41845.4]
  wire [13:0] _T_94042; // @[Modules.scala 166:64:@41846.4]
  wire [13:0] buffer_12_574; // @[Modules.scala 166:64:@41847.4]
  wire [14:0] _T_94044; // @[Modules.scala 166:64:@41849.4]
  wire [13:0] _T_94045; // @[Modules.scala 166:64:@41850.4]
  wire [13:0] buffer_12_575; // @[Modules.scala 166:64:@41851.4]
  wire [14:0] _T_94047; // @[Modules.scala 172:66:@41853.4]
  wire [13:0] _T_94048; // @[Modules.scala 172:66:@41854.4]
  wire [13:0] buffer_12_576; // @[Modules.scala 172:66:@41855.4]
  wire [14:0] _T_94050; // @[Modules.scala 166:64:@41857.4]
  wire [13:0] _T_94051; // @[Modules.scala 166:64:@41858.4]
  wire [13:0] buffer_12_577; // @[Modules.scala 166:64:@41859.4]
  wire [14:0] _T_94053; // @[Modules.scala 166:64:@41861.4]
  wire [13:0] _T_94054; // @[Modules.scala 166:64:@41862.4]
  wire [13:0] buffer_12_578; // @[Modules.scala 166:64:@41863.4]
  wire [14:0] _T_94056; // @[Modules.scala 166:64:@41865.4]
  wire [13:0] _T_94057; // @[Modules.scala 166:64:@41866.4]
  wire [13:0] buffer_12_579; // @[Modules.scala 166:64:@41867.4]
  wire [14:0] _T_94059; // @[Modules.scala 166:64:@41869.4]
  wire [13:0] _T_94060; // @[Modules.scala 166:64:@41870.4]
  wire [13:0] buffer_12_580; // @[Modules.scala 166:64:@41871.4]
  wire [14:0] _T_94062; // @[Modules.scala 166:64:@41873.4]
  wire [13:0] _T_94063; // @[Modules.scala 166:64:@41874.4]
  wire [13:0] buffer_12_581; // @[Modules.scala 166:64:@41875.4]
  wire [14:0] _T_94065; // @[Modules.scala 166:64:@41877.4]
  wire [13:0] _T_94066; // @[Modules.scala 166:64:@41878.4]
  wire [13:0] buffer_12_582; // @[Modules.scala 166:64:@41879.4]
  wire [14:0] _T_94068; // @[Modules.scala 166:64:@41881.4]
  wire [13:0] _T_94069; // @[Modules.scala 166:64:@41882.4]
  wire [13:0] buffer_12_583; // @[Modules.scala 166:64:@41883.4]
  wire [14:0] _T_94071; // @[Modules.scala 166:64:@41885.4]
  wire [13:0] _T_94072; // @[Modules.scala 166:64:@41886.4]
  wire [13:0] buffer_12_584; // @[Modules.scala 166:64:@41887.4]
  wire [14:0] _T_94074; // @[Modules.scala 166:64:@41889.4]
  wire [13:0] _T_94075; // @[Modules.scala 166:64:@41890.4]
  wire [13:0] buffer_12_585; // @[Modules.scala 166:64:@41891.4]
  wire [14:0] _T_94077; // @[Modules.scala 166:64:@41893.4]
  wire [13:0] _T_94078; // @[Modules.scala 166:64:@41894.4]
  wire [13:0] buffer_12_586; // @[Modules.scala 166:64:@41895.4]
  wire [14:0] _T_94080; // @[Modules.scala 166:64:@41897.4]
  wire [13:0] _T_94081; // @[Modules.scala 166:64:@41898.4]
  wire [13:0] buffer_12_587; // @[Modules.scala 166:64:@41899.4]
  wire [14:0] _T_94083; // @[Modules.scala 166:64:@41901.4]
  wire [13:0] _T_94084; // @[Modules.scala 166:64:@41902.4]
  wire [13:0] buffer_12_588; // @[Modules.scala 166:64:@41903.4]
  wire [14:0] _T_94086; // @[Modules.scala 166:64:@41905.4]
  wire [13:0] _T_94087; // @[Modules.scala 166:64:@41906.4]
  wire [13:0] buffer_12_589; // @[Modules.scala 166:64:@41907.4]
  wire [14:0] _T_94089; // @[Modules.scala 172:66:@41909.4]
  wire [13:0] _T_94090; // @[Modules.scala 172:66:@41910.4]
  wire [13:0] buffer_12_590; // @[Modules.scala 172:66:@41911.4]
  wire [14:0] _T_94092; // @[Modules.scala 166:64:@41913.4]
  wire [13:0] _T_94093; // @[Modules.scala 166:64:@41914.4]
  wire [13:0] buffer_12_591; // @[Modules.scala 166:64:@41915.4]
  wire [14:0] _T_94095; // @[Modules.scala 166:64:@41917.4]
  wire [13:0] _T_94096; // @[Modules.scala 166:64:@41918.4]
  wire [13:0] buffer_12_592; // @[Modules.scala 166:64:@41919.4]
  wire [14:0] _T_94098; // @[Modules.scala 160:64:@41921.4]
  wire [13:0] _T_94099; // @[Modules.scala 160:64:@41922.4]
  wire [13:0] buffer_12_593; // @[Modules.scala 160:64:@41923.4]
  wire [14:0] _T_94101; // @[Modules.scala 172:66:@41925.4]
  wire [13:0] _T_94102; // @[Modules.scala 172:66:@41926.4]
  wire [13:0] buffer_12_594; // @[Modules.scala 172:66:@41927.4]
  wire [4:0] _T_94105; // @[Modules.scala 143:74:@42118.4]
  wire [5:0] _T_94108; // @[Modules.scala 143:103:@42120.4]
  wire [4:0] _T_94109; // @[Modules.scala 143:103:@42121.4]
  wire [4:0] _T_94110; // @[Modules.scala 143:103:@42122.4]
  wire [4:0] _T_94114; // @[Modules.scala 144:80:@42125.4]
  wire [5:0] _T_94115; // @[Modules.scala 143:103:@42126.4]
  wire [4:0] _T_94116; // @[Modules.scala 143:103:@42127.4]
  wire [4:0] _T_94117; // @[Modules.scala 143:103:@42128.4]
  wire [6:0] _T_94143; // @[Modules.scala 143:103:@42150.4]
  wire [5:0] _T_94144; // @[Modules.scala 143:103:@42151.4]
  wire [5:0] _T_94145; // @[Modules.scala 143:103:@42152.4]
  wire [6:0] _T_94150; // @[Modules.scala 143:103:@42156.4]
  wire [5:0] _T_94151; // @[Modules.scala 143:103:@42157.4]
  wire [5:0] _T_94152; // @[Modules.scala 143:103:@42158.4]
  wire [5:0] _T_94164; // @[Modules.scala 143:103:@42168.4]
  wire [4:0] _T_94165; // @[Modules.scala 143:103:@42169.4]
  wire [4:0] _T_94166; // @[Modules.scala 143:103:@42170.4]
  wire [6:0] _T_94178; // @[Modules.scala 143:103:@42180.4]
  wire [5:0] _T_94179; // @[Modules.scala 143:103:@42181.4]
  wire [5:0] _T_94180; // @[Modules.scala 143:103:@42182.4]
  wire [5:0] _T_94185; // @[Modules.scala 143:103:@42186.4]
  wire [4:0] _T_94186; // @[Modules.scala 143:103:@42187.4]
  wire [4:0] _T_94187; // @[Modules.scala 143:103:@42188.4]
  wire [5:0] _GEN_909; // @[Modules.scala 143:103:@42192.4]
  wire [6:0] _T_94192; // @[Modules.scala 143:103:@42192.4]
  wire [5:0] _T_94193; // @[Modules.scala 143:103:@42193.4]
  wire [5:0] _T_94194; // @[Modules.scala 143:103:@42194.4]
  wire [4:0] _T_94254; // @[Modules.scala 144:80:@42245.4]
  wire [5:0] _GEN_910; // @[Modules.scala 143:103:@42246.4]
  wire [6:0] _T_94255; // @[Modules.scala 143:103:@42246.4]
  wire [5:0] _T_94256; // @[Modules.scala 143:103:@42247.4]
  wire [5:0] _T_94257; // @[Modules.scala 143:103:@42248.4]
  wire [5:0] _GEN_911; // @[Modules.scala 143:103:@42258.4]
  wire [6:0] _T_94269; // @[Modules.scala 143:103:@42258.4]
  wire [5:0] _T_94270; // @[Modules.scala 143:103:@42259.4]
  wire [5:0] _T_94271; // @[Modules.scala 143:103:@42260.4]
  wire [6:0] _T_94360; // @[Modules.scala 143:103:@42336.4]
  wire [5:0] _T_94361; // @[Modules.scala 143:103:@42337.4]
  wire [5:0] _T_94362; // @[Modules.scala 143:103:@42338.4]
  wire [6:0] _T_94395; // @[Modules.scala 143:103:@42366.4]
  wire [5:0] _T_94396; // @[Modules.scala 143:103:@42367.4]
  wire [5:0] _T_94397; // @[Modules.scala 143:103:@42368.4]
  wire [6:0] _T_94402; // @[Modules.scala 143:103:@42372.4]
  wire [5:0] _T_94403; // @[Modules.scala 143:103:@42373.4]
  wire [5:0] _T_94404; // @[Modules.scala 143:103:@42374.4]
  wire [6:0] _T_94423; // @[Modules.scala 143:103:@42390.4]
  wire [5:0] _T_94424; // @[Modules.scala 143:103:@42391.4]
  wire [5:0] _T_94425; // @[Modules.scala 143:103:@42392.4]
  wire [6:0] _T_94444; // @[Modules.scala 143:103:@42408.4]
  wire [5:0] _T_94445; // @[Modules.scala 143:103:@42409.4]
  wire [5:0] _T_94446; // @[Modules.scala 143:103:@42410.4]
  wire [6:0] _T_94451; // @[Modules.scala 143:103:@42414.4]
  wire [5:0] _T_94452; // @[Modules.scala 143:103:@42415.4]
  wire [5:0] _T_94453; // @[Modules.scala 143:103:@42416.4]
  wire [5:0] _T_94493; // @[Modules.scala 143:103:@42450.4]
  wire [4:0] _T_94494; // @[Modules.scala 143:103:@42451.4]
  wire [4:0] _T_94495; // @[Modules.scala 143:103:@42452.4]
  wire [5:0] _GEN_916; // @[Modules.scala 143:103:@42486.4]
  wire [6:0] _T_94535; // @[Modules.scala 143:103:@42486.4]
  wire [5:0] _T_94536; // @[Modules.scala 143:103:@42487.4]
  wire [5:0] _T_94537; // @[Modules.scala 143:103:@42488.4]
  wire [5:0] _T_94563; // @[Modules.scala 143:103:@42510.4]
  wire [4:0] _T_94564; // @[Modules.scala 143:103:@42511.4]
  wire [4:0] _T_94565; // @[Modules.scala 143:103:@42512.4]
  wire [5:0] _GEN_918; // @[Modules.scala 143:103:@42558.4]
  wire [6:0] _T_94619; // @[Modules.scala 143:103:@42558.4]
  wire [5:0] _T_94620; // @[Modules.scala 143:103:@42559.4]
  wire [5:0] _T_94621; // @[Modules.scala 143:103:@42560.4]
  wire [5:0] _T_94626; // @[Modules.scala 143:103:@42564.4]
  wire [4:0] _T_94627; // @[Modules.scala 143:103:@42565.4]
  wire [4:0] _T_94628; // @[Modules.scala 143:103:@42566.4]
  wire [5:0] _T_94647; // @[Modules.scala 143:103:@42582.4]
  wire [4:0] _T_94648; // @[Modules.scala 143:103:@42583.4]
  wire [4:0] _T_94649; // @[Modules.scala 143:103:@42584.4]
  wire [5:0] _GEN_920; // @[Modules.scala 143:103:@42594.4]
  wire [6:0] _T_94661; // @[Modules.scala 143:103:@42594.4]
  wire [5:0] _T_94662; // @[Modules.scala 143:103:@42595.4]
  wire [5:0] _T_94663; // @[Modules.scala 143:103:@42596.4]
  wire [6:0] _T_94675; // @[Modules.scala 143:103:@42606.4]
  wire [5:0] _T_94676; // @[Modules.scala 143:103:@42607.4]
  wire [5:0] _T_94677; // @[Modules.scala 143:103:@42608.4]
  wire [5:0] _T_94696; // @[Modules.scala 143:103:@42624.4]
  wire [4:0] _T_94697; // @[Modules.scala 143:103:@42625.4]
  wire [4:0] _T_94698; // @[Modules.scala 143:103:@42626.4]
  wire [5:0] _T_94703; // @[Modules.scala 143:103:@42630.4]
  wire [4:0] _T_94704; // @[Modules.scala 143:103:@42631.4]
  wire [4:0] _T_94705; // @[Modules.scala 143:103:@42632.4]
  wire [5:0] _T_94717; // @[Modules.scala 143:103:@42642.4]
  wire [4:0] _T_94718; // @[Modules.scala 143:103:@42643.4]
  wire [4:0] _T_94719; // @[Modules.scala 143:103:@42644.4]
  wire [5:0] _GEN_923; // @[Modules.scala 143:103:@42648.4]
  wire [6:0] _T_94724; // @[Modules.scala 143:103:@42648.4]
  wire [5:0] _T_94725; // @[Modules.scala 143:103:@42649.4]
  wire [5:0] _T_94726; // @[Modules.scala 143:103:@42650.4]
  wire [5:0] _GEN_924; // @[Modules.scala 143:103:@42660.4]
  wire [6:0] _T_94738; // @[Modules.scala 143:103:@42660.4]
  wire [5:0] _T_94739; // @[Modules.scala 143:103:@42661.4]
  wire [5:0] _T_94740; // @[Modules.scala 143:103:@42662.4]
  wire [6:0] _T_94773; // @[Modules.scala 143:103:@42690.4]
  wire [5:0] _T_94774; // @[Modules.scala 143:103:@42691.4]
  wire [5:0] _T_94775; // @[Modules.scala 143:103:@42692.4]
  wire [5:0] _T_94780; // @[Modules.scala 143:103:@42696.4]
  wire [4:0] _T_94781; // @[Modules.scala 143:103:@42697.4]
  wire [4:0] _T_94782; // @[Modules.scala 143:103:@42698.4]
  wire [5:0] _GEN_927; // @[Modules.scala 143:103:@42738.4]
  wire [6:0] _T_94829; // @[Modules.scala 143:103:@42738.4]
  wire [5:0] _T_94830; // @[Modules.scala 143:103:@42739.4]
  wire [5:0] _T_94831; // @[Modules.scala 143:103:@42740.4]
  wire [5:0] _T_94836; // @[Modules.scala 143:103:@42744.4]
  wire [4:0] _T_94837; // @[Modules.scala 143:103:@42745.4]
  wire [4:0] _T_94838; // @[Modules.scala 143:103:@42746.4]
  wire [6:0] _T_94843; // @[Modules.scala 143:103:@42750.4]
  wire [5:0] _T_94844; // @[Modules.scala 143:103:@42751.4]
  wire [5:0] _T_94845; // @[Modules.scala 143:103:@42752.4]
  wire [6:0] _T_94850; // @[Modules.scala 143:103:@42756.4]
  wire [5:0] _T_94851; // @[Modules.scala 143:103:@42757.4]
  wire [5:0] _T_94852; // @[Modules.scala 143:103:@42758.4]
  wire [5:0] _GEN_928; // @[Modules.scala 143:103:@42762.4]
  wire [6:0] _T_94857; // @[Modules.scala 143:103:@42762.4]
  wire [5:0] _T_94858; // @[Modules.scala 143:103:@42763.4]
  wire [5:0] _T_94859; // @[Modules.scala 143:103:@42764.4]
  wire [5:0] _T_94864; // @[Modules.scala 143:103:@42768.4]
  wire [4:0] _T_94865; // @[Modules.scala 143:103:@42769.4]
  wire [4:0] _T_94866; // @[Modules.scala 143:103:@42770.4]
  wire [5:0] _GEN_929; // @[Modules.scala 143:103:@42792.4]
  wire [6:0] _T_94892; // @[Modules.scala 143:103:@42792.4]
  wire [5:0] _T_94893; // @[Modules.scala 143:103:@42793.4]
  wire [5:0] _T_94894; // @[Modules.scala 143:103:@42794.4]
  wire [6:0] _T_94899; // @[Modules.scala 143:103:@42798.4]
  wire [5:0] _T_94900; // @[Modules.scala 143:103:@42799.4]
  wire [5:0] _T_94901; // @[Modules.scala 143:103:@42800.4]
  wire [5:0] _GEN_930; // @[Modules.scala 143:103:@42810.4]
  wire [6:0] _T_94913; // @[Modules.scala 143:103:@42810.4]
  wire [5:0] _T_94914; // @[Modules.scala 143:103:@42811.4]
  wire [5:0] _T_94915; // @[Modules.scala 143:103:@42812.4]
  wire [6:0] _T_94920; // @[Modules.scala 143:103:@42816.4]
  wire [5:0] _T_94921; // @[Modules.scala 143:103:@42817.4]
  wire [5:0] _T_94922; // @[Modules.scala 143:103:@42818.4]
  wire [5:0] _T_94927; // @[Modules.scala 143:103:@42822.4]
  wire [4:0] _T_94928; // @[Modules.scala 143:103:@42823.4]
  wire [4:0] _T_94929; // @[Modules.scala 143:103:@42824.4]
  wire [5:0] _T_94955; // @[Modules.scala 143:103:@42846.4]
  wire [4:0] _T_94956; // @[Modules.scala 143:103:@42847.4]
  wire [4:0] _T_94957; // @[Modules.scala 143:103:@42848.4]
  wire [6:0] _T_94962; // @[Modules.scala 143:103:@42852.4]
  wire [5:0] _T_94963; // @[Modules.scala 143:103:@42853.4]
  wire [5:0] _T_94964; // @[Modules.scala 143:103:@42854.4]
  wire [6:0] _T_94976; // @[Modules.scala 143:103:@42864.4]
  wire [5:0] _T_94977; // @[Modules.scala 143:103:@42865.4]
  wire [5:0] _T_94978; // @[Modules.scala 143:103:@42866.4]
  wire [5:0] _GEN_934; // @[Modules.scala 143:103:@42876.4]
  wire [6:0] _T_94990; // @[Modules.scala 143:103:@42876.4]
  wire [5:0] _T_94991; // @[Modules.scala 143:103:@42877.4]
  wire [5:0] _T_94992; // @[Modules.scala 143:103:@42878.4]
  wire [6:0] _T_95032; // @[Modules.scala 143:103:@42912.4]
  wire [5:0] _T_95033; // @[Modules.scala 143:103:@42913.4]
  wire [5:0] _T_95034; // @[Modules.scala 143:103:@42914.4]
  wire [5:0] _T_95039; // @[Modules.scala 143:103:@42918.4]
  wire [4:0] _T_95040; // @[Modules.scala 143:103:@42919.4]
  wire [4:0] _T_95041; // @[Modules.scala 143:103:@42920.4]
  wire [5:0] _GEN_935; // @[Modules.scala 143:103:@42930.4]
  wire [6:0] _T_95053; // @[Modules.scala 143:103:@42930.4]
  wire [5:0] _T_95054; // @[Modules.scala 143:103:@42931.4]
  wire [5:0] _T_95055; // @[Modules.scala 143:103:@42932.4]
  wire [5:0] _GEN_936; // @[Modules.scala 143:103:@42948.4]
  wire [6:0] _T_95074; // @[Modules.scala 143:103:@42948.4]
  wire [5:0] _T_95075; // @[Modules.scala 143:103:@42949.4]
  wire [5:0] _T_95076; // @[Modules.scala 143:103:@42950.4]
  wire [6:0] _T_95102; // @[Modules.scala 143:103:@42972.4]
  wire [5:0] _T_95103; // @[Modules.scala 143:103:@42973.4]
  wire [5:0] _T_95104; // @[Modules.scala 143:103:@42974.4]
  wire [5:0] _GEN_938; // @[Modules.scala 143:103:@42990.4]
  wire [6:0] _T_95123; // @[Modules.scala 143:103:@42990.4]
  wire [5:0] _T_95124; // @[Modules.scala 143:103:@42991.4]
  wire [5:0] _T_95125; // @[Modules.scala 143:103:@42992.4]
  wire [5:0] _GEN_939; // @[Modules.scala 143:103:@42996.4]
  wire [6:0] _T_95130; // @[Modules.scala 143:103:@42996.4]
  wire [5:0] _T_95131; // @[Modules.scala 143:103:@42997.4]
  wire [5:0] _T_95132; // @[Modules.scala 143:103:@42998.4]
  wire [6:0] _T_95151; // @[Modules.scala 143:103:@43014.4]
  wire [5:0] _T_95152; // @[Modules.scala 143:103:@43015.4]
  wire [5:0] _T_95153; // @[Modules.scala 143:103:@43016.4]
  wire [5:0] _T_95172; // @[Modules.scala 143:103:@43032.4]
  wire [4:0] _T_95173; // @[Modules.scala 143:103:@43033.4]
  wire [4:0] _T_95174; // @[Modules.scala 143:103:@43034.4]
  wire [5:0] _T_95214; // @[Modules.scala 143:103:@43068.4]
  wire [4:0] _T_95215; // @[Modules.scala 143:103:@43069.4]
  wire [4:0] _T_95216; // @[Modules.scala 143:103:@43070.4]
  wire [5:0] _GEN_940; // @[Modules.scala 143:103:@43080.4]
  wire [6:0] _T_95228; // @[Modules.scala 143:103:@43080.4]
  wire [5:0] _T_95229; // @[Modules.scala 143:103:@43081.4]
  wire [5:0] _T_95230; // @[Modules.scala 143:103:@43082.4]
  wire [6:0] _T_95235; // @[Modules.scala 143:103:@43086.4]
  wire [5:0] _T_95236; // @[Modules.scala 143:103:@43087.4]
  wire [5:0] _T_95237; // @[Modules.scala 143:103:@43088.4]
  wire [6:0] _T_95242; // @[Modules.scala 143:103:@43092.4]
  wire [5:0] _T_95243; // @[Modules.scala 143:103:@43093.4]
  wire [5:0] _T_95244; // @[Modules.scala 143:103:@43094.4]
  wire [6:0] _T_95270; // @[Modules.scala 143:103:@43116.4]
  wire [5:0] _T_95271; // @[Modules.scala 143:103:@43117.4]
  wire [5:0] _T_95272; // @[Modules.scala 143:103:@43118.4]
  wire [6:0] _T_95277; // @[Modules.scala 143:103:@43122.4]
  wire [5:0] _T_95278; // @[Modules.scala 143:103:@43123.4]
  wire [5:0] _T_95279; // @[Modules.scala 143:103:@43124.4]
  wire [5:0] _GEN_942; // @[Modules.scala 143:103:@43146.4]
  wire [6:0] _T_95305; // @[Modules.scala 143:103:@43146.4]
  wire [5:0] _T_95306; // @[Modules.scala 143:103:@43147.4]
  wire [5:0] _T_95307; // @[Modules.scala 143:103:@43148.4]
  wire [5:0] _T_95312; // @[Modules.scala 143:103:@43152.4]
  wire [4:0] _T_95313; // @[Modules.scala 143:103:@43153.4]
  wire [4:0] _T_95314; // @[Modules.scala 143:103:@43154.4]
  wire [6:0] _T_95326; // @[Modules.scala 143:103:@43164.4]
  wire [5:0] _T_95327; // @[Modules.scala 143:103:@43165.4]
  wire [5:0] _T_95328; // @[Modules.scala 143:103:@43166.4]
  wire [6:0] _T_95375; // @[Modules.scala 143:103:@43206.4]
  wire [5:0] _T_95376; // @[Modules.scala 143:103:@43207.4]
  wire [5:0] _T_95377; // @[Modules.scala 143:103:@43208.4]
  wire [6:0] _T_95389; // @[Modules.scala 143:103:@43218.4]
  wire [5:0] _T_95390; // @[Modules.scala 143:103:@43219.4]
  wire [5:0] _T_95391; // @[Modules.scala 143:103:@43220.4]
  wire [6:0] _T_95410; // @[Modules.scala 143:103:@43236.4]
  wire [5:0] _T_95411; // @[Modules.scala 143:103:@43237.4]
  wire [5:0] _T_95412; // @[Modules.scala 143:103:@43238.4]
  wire [6:0] _T_95452; // @[Modules.scala 143:103:@43272.4]
  wire [5:0] _T_95453; // @[Modules.scala 143:103:@43273.4]
  wire [5:0] _T_95454; // @[Modules.scala 143:103:@43274.4]
  wire [5:0] _GEN_946; // @[Modules.scala 143:103:@43278.4]
  wire [6:0] _T_95459; // @[Modules.scala 143:103:@43278.4]
  wire [5:0] _T_95460; // @[Modules.scala 143:103:@43279.4]
  wire [5:0] _T_95461; // @[Modules.scala 143:103:@43280.4]
  wire [5:0] _T_95494; // @[Modules.scala 143:103:@43308.4]
  wire [4:0] _T_95495; // @[Modules.scala 143:103:@43309.4]
  wire [4:0] _T_95496; // @[Modules.scala 143:103:@43310.4]
  wire [6:0] _T_95508; // @[Modules.scala 143:103:@43320.4]
  wire [5:0] _T_95509; // @[Modules.scala 143:103:@43321.4]
  wire [5:0] _T_95510; // @[Modules.scala 143:103:@43322.4]
  wire [6:0] _T_95536; // @[Modules.scala 143:103:@43344.4]
  wire [5:0] _T_95537; // @[Modules.scala 143:103:@43345.4]
  wire [5:0] _T_95538; // @[Modules.scala 143:103:@43346.4]
  wire [5:0] _GEN_951; // @[Modules.scala 143:103:@43374.4]
  wire [6:0] _T_95571; // @[Modules.scala 143:103:@43374.4]
  wire [5:0] _T_95572; // @[Modules.scala 143:103:@43375.4]
  wire [5:0] _T_95573; // @[Modules.scala 143:103:@43376.4]
  wire [6:0] _T_95578; // @[Modules.scala 143:103:@43380.4]
  wire [5:0] _T_95579; // @[Modules.scala 143:103:@43381.4]
  wire [5:0] _T_95580; // @[Modules.scala 143:103:@43382.4]
  wire [6:0] _T_95585; // @[Modules.scala 143:103:@43386.4]
  wire [5:0] _T_95586; // @[Modules.scala 143:103:@43387.4]
  wire [5:0] _T_95587; // @[Modules.scala 143:103:@43388.4]
  wire [6:0] _T_95592; // @[Modules.scala 143:103:@43392.4]
  wire [5:0] _T_95593; // @[Modules.scala 143:103:@43393.4]
  wire [5:0] _T_95594; // @[Modules.scala 143:103:@43394.4]
  wire [6:0] _T_95620; // @[Modules.scala 143:103:@43416.4]
  wire [5:0] _T_95621; // @[Modules.scala 143:103:@43417.4]
  wire [5:0] _T_95622; // @[Modules.scala 143:103:@43418.4]
  wire [6:0] _T_95627; // @[Modules.scala 143:103:@43422.4]
  wire [5:0] _T_95628; // @[Modules.scala 143:103:@43423.4]
  wire [5:0] _T_95629; // @[Modules.scala 143:103:@43424.4]
  wire [6:0] _T_95704; // @[Modules.scala 143:103:@43488.4]
  wire [5:0] _T_95705; // @[Modules.scala 143:103:@43489.4]
  wire [5:0] _T_95706; // @[Modules.scala 143:103:@43490.4]
  wire [5:0] _GEN_957; // @[Modules.scala 143:103:@43524.4]
  wire [6:0] _T_95746; // @[Modules.scala 143:103:@43524.4]
  wire [5:0] _T_95747; // @[Modules.scala 143:103:@43525.4]
  wire [5:0] _T_95748; // @[Modules.scala 143:103:@43526.4]
  wire [6:0] _T_95781; // @[Modules.scala 143:103:@43554.4]
  wire [5:0] _T_95782; // @[Modules.scala 143:103:@43555.4]
  wire [5:0] _T_95783; // @[Modules.scala 143:103:@43556.4]
  wire [6:0] _T_95823; // @[Modules.scala 143:103:@43590.4]
  wire [5:0] _T_95824; // @[Modules.scala 143:103:@43591.4]
  wire [5:0] _T_95825; // @[Modules.scala 143:103:@43592.4]
  wire [6:0] _T_95844; // @[Modules.scala 143:103:@43608.4]
  wire [5:0] _T_95845; // @[Modules.scala 143:103:@43609.4]
  wire [5:0] _T_95846; // @[Modules.scala 143:103:@43610.4]
  wire [5:0] _GEN_964; // @[Modules.scala 143:103:@43614.4]
  wire [6:0] _T_95851; // @[Modules.scala 143:103:@43614.4]
  wire [5:0] _T_95852; // @[Modules.scala 143:103:@43615.4]
  wire [5:0] _T_95853; // @[Modules.scala 143:103:@43616.4]
  wire [5:0] _GEN_965; // @[Modules.scala 143:103:@43650.4]
  wire [6:0] _T_95893; // @[Modules.scala 143:103:@43650.4]
  wire [5:0] _T_95894; // @[Modules.scala 143:103:@43651.4]
  wire [5:0] _T_95895; // @[Modules.scala 143:103:@43652.4]
  wire [6:0] _T_95900; // @[Modules.scala 143:103:@43656.4]
  wire [5:0] _T_95901; // @[Modules.scala 143:103:@43657.4]
  wire [5:0] _T_95902; // @[Modules.scala 143:103:@43658.4]
  wire [6:0] _T_95907; // @[Modules.scala 143:103:@43662.4]
  wire [5:0] _T_95908; // @[Modules.scala 143:103:@43663.4]
  wire [5:0] _T_95909; // @[Modules.scala 143:103:@43664.4]
  wire [5:0] _GEN_966; // @[Modules.scala 143:103:@43674.4]
  wire [6:0] _T_95921; // @[Modules.scala 143:103:@43674.4]
  wire [5:0] _T_95922; // @[Modules.scala 143:103:@43675.4]
  wire [5:0] _T_95923; // @[Modules.scala 143:103:@43676.4]
  wire [5:0] _GEN_968; // @[Modules.scala 143:103:@43734.4]
  wire [6:0] _T_95991; // @[Modules.scala 143:103:@43734.4]
  wire [5:0] _T_95992; // @[Modules.scala 143:103:@43735.4]
  wire [5:0] _T_95993; // @[Modules.scala 143:103:@43736.4]
  wire [6:0] _T_95998; // @[Modules.scala 143:103:@43740.4]
  wire [5:0] _T_95999; // @[Modules.scala 143:103:@43741.4]
  wire [5:0] _T_96000; // @[Modules.scala 143:103:@43742.4]
  wire [5:0] _T_96075; // @[Modules.scala 143:103:@43806.4]
  wire [4:0] _T_96076; // @[Modules.scala 143:103:@43807.4]
  wire [4:0] _T_96077; // @[Modules.scala 143:103:@43808.4]
  wire [5:0] _T_96138; // @[Modules.scala 143:103:@43860.4]
  wire [4:0] _T_96139; // @[Modules.scala 143:103:@43861.4]
  wire [4:0] _T_96140; // @[Modules.scala 143:103:@43862.4]
  wire [6:0] _T_96215; // @[Modules.scala 143:103:@43926.4]
  wire [5:0] _T_96216; // @[Modules.scala 143:103:@43927.4]
  wire [5:0] _T_96217; // @[Modules.scala 143:103:@43928.4]
  wire [5:0] _GEN_974; // @[Modules.scala 143:103:@43938.4]
  wire [6:0] _T_96229; // @[Modules.scala 143:103:@43938.4]
  wire [5:0] _T_96230; // @[Modules.scala 143:103:@43939.4]
  wire [5:0] _T_96231; // @[Modules.scala 143:103:@43940.4]
  wire [13:0] buffer_13_0; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96253; // @[Modules.scala 166:64:@43960.4]
  wire [13:0] _T_96254; // @[Modules.scala 166:64:@43961.4]
  wire [13:0] buffer_13_307; // @[Modules.scala 166:64:@43962.4]
  wire [14:0] _T_96256; // @[Modules.scala 166:64:@43964.4]
  wire [13:0] _T_96257; // @[Modules.scala 166:64:@43965.4]
  wire [13:0] buffer_13_308; // @[Modules.scala 166:64:@43966.4]
  wire [13:0] buffer_13_5; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96259; // @[Modules.scala 166:64:@43968.4]
  wire [13:0] _T_96260; // @[Modules.scala 166:64:@43969.4]
  wire [13:0] buffer_13_309; // @[Modules.scala 166:64:@43970.4]
  wire [13:0] buffer_13_6; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96262; // @[Modules.scala 166:64:@43972.4]
  wire [13:0] _T_96263; // @[Modules.scala 166:64:@43973.4]
  wire [13:0] buffer_13_310; // @[Modules.scala 166:64:@43974.4]
  wire [13:0] buffer_13_8; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96265; // @[Modules.scala 166:64:@43976.4]
  wire [13:0] _T_96266; // @[Modules.scala 166:64:@43977.4]
  wire [13:0] buffer_13_311; // @[Modules.scala 166:64:@43978.4]
  wire [13:0] buffer_13_10; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_11; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96268; // @[Modules.scala 166:64:@43980.4]
  wire [13:0] _T_96269; // @[Modules.scala 166:64:@43981.4]
  wire [13:0] buffer_13_312; // @[Modules.scala 166:64:@43982.4]
  wire [13:0] buffer_13_12; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96271; // @[Modules.scala 166:64:@43984.4]
  wire [13:0] _T_96272; // @[Modules.scala 166:64:@43985.4]
  wire [13:0] buffer_13_313; // @[Modules.scala 166:64:@43986.4]
  wire [13:0] buffer_13_21; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96283; // @[Modules.scala 166:64:@44000.4]
  wire [13:0] _T_96284; // @[Modules.scala 166:64:@44001.4]
  wire [13:0] buffer_13_317; // @[Modules.scala 166:64:@44002.4]
  wire [13:0] buffer_13_23; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96286; // @[Modules.scala 166:64:@44004.4]
  wire [13:0] _T_96287; // @[Modules.scala 166:64:@44005.4]
  wire [13:0] buffer_13_318; // @[Modules.scala 166:64:@44006.4]
  wire [14:0] _T_96304; // @[Modules.scala 166:64:@44028.4]
  wire [13:0] _T_96305; // @[Modules.scala 166:64:@44029.4]
  wire [13:0] buffer_13_324; // @[Modules.scala 166:64:@44030.4]
  wire [13:0] buffer_13_36; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96307; // @[Modules.scala 166:64:@44032.4]
  wire [13:0] _T_96308; // @[Modules.scala 166:64:@44033.4]
  wire [13:0] buffer_13_325; // @[Modules.scala 166:64:@44034.4]
  wire [14:0] _T_96310; // @[Modules.scala 166:64:@44036.4]
  wire [13:0] _T_96311; // @[Modules.scala 166:64:@44037.4]
  wire [13:0] buffer_13_326; // @[Modules.scala 166:64:@44038.4]
  wire [13:0] buffer_13_41; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96313; // @[Modules.scala 166:64:@44040.4]
  wire [13:0] _T_96314; // @[Modules.scala 166:64:@44041.4]
  wire [13:0] buffer_13_327; // @[Modules.scala 166:64:@44042.4]
  wire [13:0] buffer_13_42; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96316; // @[Modules.scala 166:64:@44044.4]
  wire [13:0] _T_96317; // @[Modules.scala 166:64:@44045.4]
  wire [13:0] buffer_13_328; // @[Modules.scala 166:64:@44046.4]
  wire [13:0] buffer_13_45; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96319; // @[Modules.scala 166:64:@44048.4]
  wire [13:0] _T_96320; // @[Modules.scala 166:64:@44049.4]
  wire [13:0] buffer_13_329; // @[Modules.scala 166:64:@44050.4]
  wire [13:0] buffer_13_48; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96325; // @[Modules.scala 166:64:@44056.4]
  wire [13:0] _T_96326; // @[Modules.scala 166:64:@44057.4]
  wire [13:0] buffer_13_331; // @[Modules.scala 166:64:@44058.4]
  wire [14:0] _T_96331; // @[Modules.scala 166:64:@44064.4]
  wire [13:0] _T_96332; // @[Modules.scala 166:64:@44065.4]
  wire [13:0] buffer_13_333; // @[Modules.scala 166:64:@44066.4]
  wire [13:0] buffer_13_55; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96334; // @[Modules.scala 166:64:@44068.4]
  wire [13:0] _T_96335; // @[Modules.scala 166:64:@44069.4]
  wire [13:0] buffer_13_334; // @[Modules.scala 166:64:@44070.4]
  wire [14:0] _T_96337; // @[Modules.scala 166:64:@44072.4]
  wire [13:0] _T_96338; // @[Modules.scala 166:64:@44073.4]
  wire [13:0] buffer_13_335; // @[Modules.scala 166:64:@44074.4]
  wire [14:0] _T_96340; // @[Modules.scala 166:64:@44076.4]
  wire [13:0] _T_96341; // @[Modules.scala 166:64:@44077.4]
  wire [13:0] buffer_13_336; // @[Modules.scala 166:64:@44078.4]
  wire [13:0] buffer_13_61; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96343; // @[Modules.scala 166:64:@44080.4]
  wire [13:0] _T_96344; // @[Modules.scala 166:64:@44081.4]
  wire [13:0] buffer_13_337; // @[Modules.scala 166:64:@44082.4]
  wire [13:0] buffer_13_65; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96349; // @[Modules.scala 166:64:@44088.4]
  wire [13:0] _T_96350; // @[Modules.scala 166:64:@44089.4]
  wire [13:0] buffer_13_339; // @[Modules.scala 166:64:@44090.4]
  wire [14:0] _T_96352; // @[Modules.scala 166:64:@44092.4]
  wire [13:0] _T_96353; // @[Modules.scala 166:64:@44093.4]
  wire [13:0] buffer_13_340; // @[Modules.scala 166:64:@44094.4]
  wire [14:0] _T_96355; // @[Modules.scala 166:64:@44096.4]
  wire [13:0] _T_96356; // @[Modules.scala 166:64:@44097.4]
  wire [13:0] buffer_13_341; // @[Modules.scala 166:64:@44098.4]
  wire [14:0] _T_96358; // @[Modules.scala 166:64:@44100.4]
  wire [13:0] _T_96359; // @[Modules.scala 166:64:@44101.4]
  wire [13:0] buffer_13_342; // @[Modules.scala 166:64:@44102.4]
  wire [13:0] buffer_13_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96361; // @[Modules.scala 166:64:@44104.4]
  wire [13:0] _T_96362; // @[Modules.scala 166:64:@44105.4]
  wire [13:0] buffer_13_343; // @[Modules.scala 166:64:@44106.4]
  wire [13:0] buffer_13_74; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96364; // @[Modules.scala 166:64:@44108.4]
  wire [13:0] _T_96365; // @[Modules.scala 166:64:@44109.4]
  wire [13:0] buffer_13_344; // @[Modules.scala 166:64:@44110.4]
  wire [13:0] buffer_13_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96367; // @[Modules.scala 166:64:@44112.4]
  wire [13:0] _T_96368; // @[Modules.scala 166:64:@44113.4]
  wire [13:0] buffer_13_345; // @[Modules.scala 166:64:@44114.4]
  wire [13:0] buffer_13_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96370; // @[Modules.scala 166:64:@44116.4]
  wire [13:0] _T_96371; // @[Modules.scala 166:64:@44117.4]
  wire [13:0] buffer_13_346; // @[Modules.scala 166:64:@44118.4]
  wire [13:0] buffer_13_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96373; // @[Modules.scala 166:64:@44120.4]
  wire [13:0] _T_96374; // @[Modules.scala 166:64:@44121.4]
  wire [13:0] buffer_13_347; // @[Modules.scala 166:64:@44122.4]
  wire [13:0] buffer_13_84; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_85; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96379; // @[Modules.scala 166:64:@44128.4]
  wire [13:0] _T_96380; // @[Modules.scala 166:64:@44129.4]
  wire [13:0] buffer_13_349; // @[Modules.scala 166:64:@44130.4]
  wire [13:0] buffer_13_87; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96382; // @[Modules.scala 166:64:@44132.4]
  wire [13:0] _T_96383; // @[Modules.scala 166:64:@44133.4]
  wire [13:0] buffer_13_350; // @[Modules.scala 166:64:@44134.4]
  wire [13:0] buffer_13_88; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96385; // @[Modules.scala 166:64:@44136.4]
  wire [13:0] _T_96386; // @[Modules.scala 166:64:@44137.4]
  wire [13:0] buffer_13_351; // @[Modules.scala 166:64:@44138.4]
  wire [13:0] buffer_13_90; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96388; // @[Modules.scala 166:64:@44140.4]
  wire [13:0] _T_96389; // @[Modules.scala 166:64:@44141.4]
  wire [13:0] buffer_13_352; // @[Modules.scala 166:64:@44142.4]
  wire [14:0] _T_96391; // @[Modules.scala 166:64:@44144.4]
  wire [13:0] _T_96392; // @[Modules.scala 166:64:@44145.4]
  wire [13:0] buffer_13_353; // @[Modules.scala 166:64:@44146.4]
  wire [13:0] buffer_13_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96394; // @[Modules.scala 166:64:@44148.4]
  wire [13:0] _T_96395; // @[Modules.scala 166:64:@44149.4]
  wire [13:0] buffer_13_354; // @[Modules.scala 166:64:@44150.4]
  wire [13:0] buffer_13_96; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96397; // @[Modules.scala 166:64:@44152.4]
  wire [13:0] _T_96398; // @[Modules.scala 166:64:@44153.4]
  wire [13:0] buffer_13_355; // @[Modules.scala 166:64:@44154.4]
  wire [13:0] buffer_13_103; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96406; // @[Modules.scala 166:64:@44164.4]
  wire [13:0] _T_96407; // @[Modules.scala 166:64:@44165.4]
  wire [13:0] buffer_13_358; // @[Modules.scala 166:64:@44166.4]
  wire [13:0] buffer_13_104; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96409; // @[Modules.scala 166:64:@44168.4]
  wire [13:0] _T_96410; // @[Modules.scala 166:64:@44169.4]
  wire [13:0] buffer_13_359; // @[Modules.scala 166:64:@44170.4]
  wire [13:0] buffer_13_106; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_107; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96412; // @[Modules.scala 166:64:@44172.4]
  wire [13:0] _T_96413; // @[Modules.scala 166:64:@44173.4]
  wire [13:0] buffer_13_360; // @[Modules.scala 166:64:@44174.4]
  wire [13:0] buffer_13_108; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96415; // @[Modules.scala 166:64:@44176.4]
  wire [13:0] _T_96416; // @[Modules.scala 166:64:@44177.4]
  wire [13:0] buffer_13_361; // @[Modules.scala 166:64:@44178.4]
  wire [13:0] buffer_13_112; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_113; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96421; // @[Modules.scala 166:64:@44184.4]
  wire [13:0] _T_96422; // @[Modules.scala 166:64:@44185.4]
  wire [13:0] buffer_13_363; // @[Modules.scala 166:64:@44186.4]
  wire [13:0] buffer_13_115; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96424; // @[Modules.scala 166:64:@44188.4]
  wire [13:0] _T_96425; // @[Modules.scala 166:64:@44189.4]
  wire [13:0] buffer_13_364; // @[Modules.scala 166:64:@44190.4]
  wire [13:0] buffer_13_116; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_117; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96427; // @[Modules.scala 166:64:@44192.4]
  wire [13:0] _T_96428; // @[Modules.scala 166:64:@44193.4]
  wire [13:0] buffer_13_365; // @[Modules.scala 166:64:@44194.4]
  wire [13:0] buffer_13_121; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96433; // @[Modules.scala 166:64:@44200.4]
  wire [13:0] _T_96434; // @[Modules.scala 166:64:@44201.4]
  wire [13:0] buffer_13_367; // @[Modules.scala 166:64:@44202.4]
  wire [13:0] buffer_13_122; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96436; // @[Modules.scala 166:64:@44204.4]
  wire [13:0] _T_96437; // @[Modules.scala 166:64:@44205.4]
  wire [13:0] buffer_13_368; // @[Modules.scala 166:64:@44206.4]
  wire [13:0] buffer_13_124; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96439; // @[Modules.scala 166:64:@44208.4]
  wire [13:0] _T_96440; // @[Modules.scala 166:64:@44209.4]
  wire [13:0] buffer_13_369; // @[Modules.scala 166:64:@44210.4]
  wire [13:0] buffer_13_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96442; // @[Modules.scala 166:64:@44212.4]
  wire [13:0] _T_96443; // @[Modules.scala 166:64:@44213.4]
  wire [13:0] buffer_13_370; // @[Modules.scala 166:64:@44214.4]
  wire [14:0] _T_96445; // @[Modules.scala 166:64:@44216.4]
  wire [13:0] _T_96446; // @[Modules.scala 166:64:@44217.4]
  wire [13:0] buffer_13_371; // @[Modules.scala 166:64:@44218.4]
  wire [14:0] _T_96448; // @[Modules.scala 166:64:@44220.4]
  wire [13:0] _T_96449; // @[Modules.scala 166:64:@44221.4]
  wire [13:0] buffer_13_372; // @[Modules.scala 166:64:@44222.4]
  wire [13:0] buffer_13_132; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_133; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96451; // @[Modules.scala 166:64:@44224.4]
  wire [13:0] _T_96452; // @[Modules.scala 166:64:@44225.4]
  wire [13:0] buffer_13_373; // @[Modules.scala 166:64:@44226.4]
  wire [13:0] buffer_13_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96454; // @[Modules.scala 166:64:@44228.4]
  wire [13:0] _T_96455; // @[Modules.scala 166:64:@44229.4]
  wire [13:0] buffer_13_374; // @[Modules.scala 166:64:@44230.4]
  wire [14:0] _T_96457; // @[Modules.scala 166:64:@44232.4]
  wire [13:0] _T_96458; // @[Modules.scala 166:64:@44233.4]
  wire [13:0] buffer_13_375; // @[Modules.scala 166:64:@44234.4]
  wire [13:0] buffer_13_138; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96460; // @[Modules.scala 166:64:@44236.4]
  wire [13:0] _T_96461; // @[Modules.scala 166:64:@44237.4]
  wire [13:0] buffer_13_376; // @[Modules.scala 166:64:@44238.4]
  wire [13:0] buffer_13_142; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96466; // @[Modules.scala 166:64:@44244.4]
  wire [13:0] _T_96467; // @[Modules.scala 166:64:@44245.4]
  wire [13:0] buffer_13_378; // @[Modules.scala 166:64:@44246.4]
  wire [13:0] buffer_13_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96469; // @[Modules.scala 166:64:@44248.4]
  wire [13:0] _T_96470; // @[Modules.scala 166:64:@44249.4]
  wire [13:0] buffer_13_379; // @[Modules.scala 166:64:@44250.4]
  wire [13:0] buffer_13_146; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96472; // @[Modules.scala 166:64:@44252.4]
  wire [13:0] _T_96473; // @[Modules.scala 166:64:@44253.4]
  wire [13:0] buffer_13_380; // @[Modules.scala 166:64:@44254.4]
  wire [13:0] buffer_13_149; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96475; // @[Modules.scala 166:64:@44256.4]
  wire [13:0] _T_96476; // @[Modules.scala 166:64:@44257.4]
  wire [13:0] buffer_13_381; // @[Modules.scala 166:64:@44258.4]
  wire [14:0] _T_96478; // @[Modules.scala 166:64:@44260.4]
  wire [13:0] _T_96479; // @[Modules.scala 166:64:@44261.4]
  wire [13:0] buffer_13_382; // @[Modules.scala 166:64:@44262.4]
  wire [13:0] buffer_13_152; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96481; // @[Modules.scala 166:64:@44264.4]
  wire [13:0] _T_96482; // @[Modules.scala 166:64:@44265.4]
  wire [13:0] buffer_13_383; // @[Modules.scala 166:64:@44266.4]
  wire [14:0] _T_96484; // @[Modules.scala 166:64:@44268.4]
  wire [13:0] _T_96485; // @[Modules.scala 166:64:@44269.4]
  wire [13:0] buffer_13_384; // @[Modules.scala 166:64:@44270.4]
  wire [14:0] _T_96487; // @[Modules.scala 166:64:@44272.4]
  wire [13:0] _T_96488; // @[Modules.scala 166:64:@44273.4]
  wire [13:0] buffer_13_385; // @[Modules.scala 166:64:@44274.4]
  wire [13:0] buffer_13_158; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96490; // @[Modules.scala 166:64:@44276.4]
  wire [13:0] _T_96491; // @[Modules.scala 166:64:@44277.4]
  wire [13:0] buffer_13_386; // @[Modules.scala 166:64:@44278.4]
  wire [13:0] buffer_13_160; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96493; // @[Modules.scala 166:64:@44280.4]
  wire [13:0] _T_96494; // @[Modules.scala 166:64:@44281.4]
  wire [13:0] buffer_13_387; // @[Modules.scala 166:64:@44282.4]
  wire [13:0] buffer_13_162; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96496; // @[Modules.scala 166:64:@44284.4]
  wire [13:0] _T_96497; // @[Modules.scala 166:64:@44285.4]
  wire [13:0] buffer_13_388; // @[Modules.scala 166:64:@44286.4]
  wire [13:0] buffer_13_166; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96502; // @[Modules.scala 166:64:@44292.4]
  wire [13:0] _T_96503; // @[Modules.scala 166:64:@44293.4]
  wire [13:0] buffer_13_390; // @[Modules.scala 166:64:@44294.4]
  wire [13:0] buffer_13_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96508; // @[Modules.scala 166:64:@44300.4]
  wire [13:0] _T_96509; // @[Modules.scala 166:64:@44301.4]
  wire [13:0] buffer_13_392; // @[Modules.scala 166:64:@44302.4]
  wire [13:0] buffer_13_172; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96511; // @[Modules.scala 166:64:@44304.4]
  wire [13:0] _T_96512; // @[Modules.scala 166:64:@44305.4]
  wire [13:0] buffer_13_393; // @[Modules.scala 166:64:@44306.4]
  wire [13:0] buffer_13_174; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96514; // @[Modules.scala 166:64:@44308.4]
  wire [13:0] _T_96515; // @[Modules.scala 166:64:@44309.4]
  wire [13:0] buffer_13_394; // @[Modules.scala 166:64:@44310.4]
  wire [14:0] _T_96517; // @[Modules.scala 166:64:@44312.4]
  wire [13:0] _T_96518; // @[Modules.scala 166:64:@44313.4]
  wire [13:0] buffer_13_395; // @[Modules.scala 166:64:@44314.4]
  wire [14:0] _T_96520; // @[Modules.scala 166:64:@44316.4]
  wire [13:0] _T_96521; // @[Modules.scala 166:64:@44317.4]
  wire [13:0] buffer_13_396; // @[Modules.scala 166:64:@44318.4]
  wire [13:0] buffer_13_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96523; // @[Modules.scala 166:64:@44320.4]
  wire [13:0] _T_96524; // @[Modules.scala 166:64:@44321.4]
  wire [13:0] buffer_13_397; // @[Modules.scala 166:64:@44322.4]
  wire [13:0] buffer_13_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96526; // @[Modules.scala 166:64:@44324.4]
  wire [13:0] _T_96527; // @[Modules.scala 166:64:@44325.4]
  wire [13:0] buffer_13_398; // @[Modules.scala 166:64:@44326.4]
  wire [13:0] buffer_13_186; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96532; // @[Modules.scala 166:64:@44332.4]
  wire [13:0] _T_96533; // @[Modules.scala 166:64:@44333.4]
  wire [13:0] buffer_13_400; // @[Modules.scala 166:64:@44334.4]
  wire [13:0] buffer_13_192; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_193; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96541; // @[Modules.scala 166:64:@44344.4]
  wire [13:0] _T_96542; // @[Modules.scala 166:64:@44345.4]
  wire [13:0] buffer_13_403; // @[Modules.scala 166:64:@44346.4]
  wire [14:0] _T_96544; // @[Modules.scala 166:64:@44348.4]
  wire [13:0] _T_96545; // @[Modules.scala 166:64:@44349.4]
  wire [13:0] buffer_13_404; // @[Modules.scala 166:64:@44350.4]
  wire [13:0] buffer_13_198; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96550; // @[Modules.scala 166:64:@44356.4]
  wire [13:0] _T_96551; // @[Modules.scala 166:64:@44357.4]
  wire [13:0] buffer_13_406; // @[Modules.scala 166:64:@44358.4]
  wire [13:0] buffer_13_200; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96553; // @[Modules.scala 166:64:@44360.4]
  wire [13:0] _T_96554; // @[Modules.scala 166:64:@44361.4]
  wire [13:0] buffer_13_407; // @[Modules.scala 166:64:@44362.4]
  wire [13:0] buffer_13_204; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96559; // @[Modules.scala 166:64:@44368.4]
  wire [13:0] _T_96560; // @[Modules.scala 166:64:@44369.4]
  wire [13:0] buffer_13_409; // @[Modules.scala 166:64:@44370.4]
  wire [14:0] _T_96562; // @[Modules.scala 166:64:@44372.4]
  wire [13:0] _T_96563; // @[Modules.scala 166:64:@44373.4]
  wire [13:0] buffer_13_410; // @[Modules.scala 166:64:@44374.4]
  wire [13:0] buffer_13_209; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96565; // @[Modules.scala 166:64:@44376.4]
  wire [13:0] _T_96566; // @[Modules.scala 166:64:@44377.4]
  wire [13:0] buffer_13_411; // @[Modules.scala 166:64:@44378.4]
  wire [13:0] buffer_13_210; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_211; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96568; // @[Modules.scala 166:64:@44380.4]
  wire [13:0] _T_96569; // @[Modules.scala 166:64:@44381.4]
  wire [13:0] buffer_13_412; // @[Modules.scala 166:64:@44382.4]
  wire [13:0] buffer_13_212; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96571; // @[Modules.scala 166:64:@44384.4]
  wire [13:0] _T_96572; // @[Modules.scala 166:64:@44385.4]
  wire [13:0] buffer_13_413; // @[Modules.scala 166:64:@44386.4]
  wire [13:0] buffer_13_216; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_217; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96577; // @[Modules.scala 166:64:@44392.4]
  wire [13:0] _T_96578; // @[Modules.scala 166:64:@44393.4]
  wire [13:0] buffer_13_415; // @[Modules.scala 166:64:@44394.4]
  wire [14:0] _T_96580; // @[Modules.scala 166:64:@44396.4]
  wire [13:0] _T_96581; // @[Modules.scala 166:64:@44397.4]
  wire [13:0] buffer_13_416; // @[Modules.scala 166:64:@44398.4]
  wire [14:0] _T_96589; // @[Modules.scala 166:64:@44408.4]
  wire [13:0] _T_96590; // @[Modules.scala 166:64:@44409.4]
  wire [13:0] buffer_13_419; // @[Modules.scala 166:64:@44410.4]
  wire [14:0] _T_96592; // @[Modules.scala 166:64:@44412.4]
  wire [13:0] _T_96593; // @[Modules.scala 166:64:@44413.4]
  wire [13:0] buffer_13_420; // @[Modules.scala 166:64:@44414.4]
  wire [13:0] buffer_13_228; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96595; // @[Modules.scala 166:64:@44416.4]
  wire [13:0] _T_96596; // @[Modules.scala 166:64:@44417.4]
  wire [13:0] buffer_13_421; // @[Modules.scala 166:64:@44418.4]
  wire [14:0] _T_96598; // @[Modules.scala 166:64:@44420.4]
  wire [13:0] _T_96599; // @[Modules.scala 166:64:@44421.4]
  wire [13:0] buffer_13_422; // @[Modules.scala 166:64:@44422.4]
  wire [14:0] _T_96601; // @[Modules.scala 166:64:@44424.4]
  wire [13:0] _T_96602; // @[Modules.scala 166:64:@44425.4]
  wire [13:0] buffer_13_423; // @[Modules.scala 166:64:@44426.4]
  wire [13:0] buffer_13_234; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96604; // @[Modules.scala 166:64:@44428.4]
  wire [13:0] _T_96605; // @[Modules.scala 166:64:@44429.4]
  wire [13:0] buffer_13_424; // @[Modules.scala 166:64:@44430.4]
  wire [14:0] _T_96607; // @[Modules.scala 166:64:@44432.4]
  wire [13:0] _T_96608; // @[Modules.scala 166:64:@44433.4]
  wire [13:0] buffer_13_425; // @[Modules.scala 166:64:@44434.4]
  wire [13:0] buffer_13_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96610; // @[Modules.scala 166:64:@44436.4]
  wire [13:0] _T_96611; // @[Modules.scala 166:64:@44437.4]
  wire [13:0] buffer_13_426; // @[Modules.scala 166:64:@44438.4]
  wire [14:0] _T_96613; // @[Modules.scala 166:64:@44440.4]
  wire [13:0] _T_96614; // @[Modules.scala 166:64:@44441.4]
  wire [13:0] buffer_13_427; // @[Modules.scala 166:64:@44442.4]
  wire [13:0] buffer_13_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96619; // @[Modules.scala 166:64:@44448.4]
  wire [13:0] _T_96620; // @[Modules.scala 166:64:@44449.4]
  wire [13:0] buffer_13_429; // @[Modules.scala 166:64:@44450.4]
  wire [14:0] _T_96622; // @[Modules.scala 166:64:@44452.4]
  wire [13:0] _T_96623; // @[Modules.scala 166:64:@44453.4]
  wire [13:0] buffer_13_430; // @[Modules.scala 166:64:@44454.4]
  wire [13:0] buffer_13_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96625; // @[Modules.scala 166:64:@44456.4]
  wire [13:0] _T_96626; // @[Modules.scala 166:64:@44457.4]
  wire [13:0] buffer_13_431; // @[Modules.scala 166:64:@44458.4]
  wire [14:0] _T_96631; // @[Modules.scala 166:64:@44464.4]
  wire [13:0] _T_96632; // @[Modules.scala 166:64:@44465.4]
  wire [13:0] buffer_13_433; // @[Modules.scala 166:64:@44466.4]
  wire [13:0] buffer_13_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96634; // @[Modules.scala 166:64:@44468.4]
  wire [13:0] _T_96635; // @[Modules.scala 166:64:@44469.4]
  wire [13:0] buffer_13_434; // @[Modules.scala 166:64:@44470.4]
  wire [13:0] buffer_13_256; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_13_257; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96637; // @[Modules.scala 166:64:@44472.4]
  wire [13:0] _T_96638; // @[Modules.scala 166:64:@44473.4]
  wire [13:0] buffer_13_435; // @[Modules.scala 166:64:@44474.4]
  wire [13:0] buffer_13_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96640; // @[Modules.scala 166:64:@44476.4]
  wire [13:0] _T_96641; // @[Modules.scala 166:64:@44477.4]
  wire [13:0] buffer_13_436; // @[Modules.scala 166:64:@44478.4]
  wire [14:0] _T_96643; // @[Modules.scala 166:64:@44480.4]
  wire [13:0] _T_96644; // @[Modules.scala 166:64:@44481.4]
  wire [13:0] buffer_13_437; // @[Modules.scala 166:64:@44482.4]
  wire [14:0] _T_96652; // @[Modules.scala 166:64:@44492.4]
  wire [13:0] _T_96653; // @[Modules.scala 166:64:@44493.4]
  wire [13:0] buffer_13_440; // @[Modules.scala 166:64:@44494.4]
  wire [13:0] buffer_13_269; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96655; // @[Modules.scala 166:64:@44496.4]
  wire [13:0] _T_96656; // @[Modules.scala 166:64:@44497.4]
  wire [13:0] buffer_13_441; // @[Modules.scala 166:64:@44498.4]
  wire [13:0] buffer_13_270; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96658; // @[Modules.scala 166:64:@44500.4]
  wire [13:0] _T_96659; // @[Modules.scala 166:64:@44501.4]
  wire [13:0] buffer_13_442; // @[Modules.scala 166:64:@44502.4]
  wire [14:0] _T_96661; // @[Modules.scala 166:64:@44504.4]
  wire [13:0] _T_96662; // @[Modules.scala 166:64:@44505.4]
  wire [13:0] buffer_13_443; // @[Modules.scala 166:64:@44506.4]
  wire [14:0] _T_96664; // @[Modules.scala 166:64:@44508.4]
  wire [13:0] _T_96665; // @[Modules.scala 166:64:@44509.4]
  wire [13:0] buffer_13_444; // @[Modules.scala 166:64:@44510.4]
  wire [14:0] _T_96667; // @[Modules.scala 166:64:@44512.4]
  wire [13:0] _T_96668; // @[Modules.scala 166:64:@44513.4]
  wire [13:0] buffer_13_445; // @[Modules.scala 166:64:@44514.4]
  wire [14:0] _T_96670; // @[Modules.scala 166:64:@44516.4]
  wire [13:0] _T_96671; // @[Modules.scala 166:64:@44517.4]
  wire [13:0] buffer_13_446; // @[Modules.scala 166:64:@44518.4]
  wire [13:0] buffer_13_281; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96673; // @[Modules.scala 166:64:@44520.4]
  wire [13:0] _T_96674; // @[Modules.scala 166:64:@44521.4]
  wire [13:0] buffer_13_447; // @[Modules.scala 166:64:@44522.4]
  wire [14:0] _T_96685; // @[Modules.scala 166:64:@44536.4]
  wire [13:0] _T_96686; // @[Modules.scala 166:64:@44537.4]
  wire [13:0] buffer_13_451; // @[Modules.scala 166:64:@44538.4]
  wire [13:0] buffer_13_290; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96688; // @[Modules.scala 166:64:@44540.4]
  wire [13:0] _T_96689; // @[Modules.scala 166:64:@44541.4]
  wire [13:0] buffer_13_452; // @[Modules.scala 166:64:@44542.4]
  wire [14:0] _T_96691; // @[Modules.scala 166:64:@44544.4]
  wire [13:0] _T_96692; // @[Modules.scala 166:64:@44545.4]
  wire [13:0] buffer_13_453; // @[Modules.scala 166:64:@44546.4]
  wire [14:0] _T_96694; // @[Modules.scala 166:64:@44548.4]
  wire [13:0] _T_96695; // @[Modules.scala 166:64:@44549.4]
  wire [13:0] buffer_13_454; // @[Modules.scala 166:64:@44550.4]
  wire [14:0] _T_96697; // @[Modules.scala 166:64:@44552.4]
  wire [13:0] _T_96698; // @[Modules.scala 166:64:@44553.4]
  wire [13:0] buffer_13_455; // @[Modules.scala 166:64:@44554.4]
  wire [14:0] _T_96700; // @[Modules.scala 166:64:@44556.4]
  wire [13:0] _T_96701; // @[Modules.scala 166:64:@44557.4]
  wire [13:0] buffer_13_456; // @[Modules.scala 166:64:@44558.4]
  wire [13:0] buffer_13_301; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96703; // @[Modules.scala 166:64:@44560.4]
  wire [13:0] _T_96704; // @[Modules.scala 166:64:@44561.4]
  wire [13:0] buffer_13_457; // @[Modules.scala 166:64:@44562.4]
  wire [13:0] buffer_13_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_96706; // @[Modules.scala 166:64:@44564.4]
  wire [13:0] _T_96707; // @[Modules.scala 166:64:@44565.4]
  wire [13:0] buffer_13_458; // @[Modules.scala 166:64:@44566.4]
  wire [14:0] _T_96709; // @[Modules.scala 166:64:@44568.4]
  wire [13:0] _T_96710; // @[Modules.scala 166:64:@44569.4]
  wire [13:0] buffer_13_459; // @[Modules.scala 166:64:@44570.4]
  wire [14:0] _T_96712; // @[Modules.scala 166:64:@44572.4]
  wire [13:0] _T_96713; // @[Modules.scala 166:64:@44573.4]
  wire [13:0] buffer_13_460; // @[Modules.scala 166:64:@44574.4]
  wire [14:0] _T_96715; // @[Modules.scala 166:64:@44576.4]
  wire [13:0] _T_96716; // @[Modules.scala 166:64:@44577.4]
  wire [13:0] buffer_13_461; // @[Modules.scala 166:64:@44578.4]
  wire [14:0] _T_96718; // @[Modules.scala 166:64:@44580.4]
  wire [13:0] _T_96719; // @[Modules.scala 166:64:@44581.4]
  wire [13:0] buffer_13_462; // @[Modules.scala 166:64:@44582.4]
  wire [14:0] _T_96721; // @[Modules.scala 166:64:@44584.4]
  wire [13:0] _T_96722; // @[Modules.scala 166:64:@44585.4]
  wire [13:0] buffer_13_463; // @[Modules.scala 166:64:@44586.4]
  wire [14:0] _T_96724; // @[Modules.scala 166:64:@44588.4]
  wire [13:0] _T_96725; // @[Modules.scala 166:64:@44589.4]
  wire [13:0] buffer_13_464; // @[Modules.scala 166:64:@44590.4]
  wire [14:0] _T_96727; // @[Modules.scala 166:64:@44592.4]
  wire [13:0] _T_96728; // @[Modules.scala 166:64:@44593.4]
  wire [13:0] buffer_13_465; // @[Modules.scala 166:64:@44594.4]
  wire [14:0] _T_96736; // @[Modules.scala 166:64:@44604.4]
  wire [13:0] _T_96737; // @[Modules.scala 166:64:@44605.4]
  wire [13:0] buffer_13_468; // @[Modules.scala 166:64:@44606.4]
  wire [14:0] _T_96739; // @[Modules.scala 166:64:@44608.4]
  wire [13:0] _T_96740; // @[Modules.scala 166:64:@44609.4]
  wire [13:0] buffer_13_469; // @[Modules.scala 166:64:@44610.4]
  wire [14:0] _T_96742; // @[Modules.scala 166:64:@44612.4]
  wire [13:0] _T_96743; // @[Modules.scala 166:64:@44613.4]
  wire [13:0] buffer_13_470; // @[Modules.scala 166:64:@44614.4]
  wire [14:0] _T_96745; // @[Modules.scala 166:64:@44616.4]
  wire [13:0] _T_96746; // @[Modules.scala 166:64:@44617.4]
  wire [13:0] buffer_13_471; // @[Modules.scala 166:64:@44618.4]
  wire [14:0] _T_96748; // @[Modules.scala 166:64:@44620.4]
  wire [13:0] _T_96749; // @[Modules.scala 166:64:@44621.4]
  wire [13:0] buffer_13_472; // @[Modules.scala 166:64:@44622.4]
  wire [14:0] _T_96751; // @[Modules.scala 166:64:@44624.4]
  wire [13:0] _T_96752; // @[Modules.scala 166:64:@44625.4]
  wire [13:0] buffer_13_473; // @[Modules.scala 166:64:@44626.4]
  wire [14:0] _T_96754; // @[Modules.scala 166:64:@44628.4]
  wire [13:0] _T_96755; // @[Modules.scala 166:64:@44629.4]
  wire [13:0] buffer_13_474; // @[Modules.scala 166:64:@44630.4]
  wire [14:0] _T_96757; // @[Modules.scala 166:64:@44632.4]
  wire [13:0] _T_96758; // @[Modules.scala 166:64:@44633.4]
  wire [13:0] buffer_13_475; // @[Modules.scala 166:64:@44634.4]
  wire [14:0] _T_96760; // @[Modules.scala 166:64:@44636.4]
  wire [13:0] _T_96761; // @[Modules.scala 166:64:@44637.4]
  wire [13:0] buffer_13_476; // @[Modules.scala 166:64:@44638.4]
  wire [14:0] _T_96763; // @[Modules.scala 166:64:@44640.4]
  wire [13:0] _T_96764; // @[Modules.scala 166:64:@44641.4]
  wire [13:0] buffer_13_477; // @[Modules.scala 166:64:@44642.4]
  wire [14:0] _T_96766; // @[Modules.scala 166:64:@44644.4]
  wire [13:0] _T_96767; // @[Modules.scala 166:64:@44645.4]
  wire [13:0] buffer_13_478; // @[Modules.scala 166:64:@44646.4]
  wire [14:0] _T_96769; // @[Modules.scala 166:64:@44648.4]
  wire [13:0] _T_96770; // @[Modules.scala 166:64:@44649.4]
  wire [13:0] buffer_13_479; // @[Modules.scala 166:64:@44650.4]
  wire [14:0] _T_96772; // @[Modules.scala 166:64:@44652.4]
  wire [13:0] _T_96773; // @[Modules.scala 166:64:@44653.4]
  wire [13:0] buffer_13_480; // @[Modules.scala 166:64:@44654.4]
  wire [14:0] _T_96775; // @[Modules.scala 166:64:@44656.4]
  wire [13:0] _T_96776; // @[Modules.scala 166:64:@44657.4]
  wire [13:0] buffer_13_481; // @[Modules.scala 166:64:@44658.4]
  wire [14:0] _T_96778; // @[Modules.scala 166:64:@44660.4]
  wire [13:0] _T_96779; // @[Modules.scala 166:64:@44661.4]
  wire [13:0] buffer_13_482; // @[Modules.scala 166:64:@44662.4]
  wire [14:0] _T_96781; // @[Modules.scala 166:64:@44664.4]
  wire [13:0] _T_96782; // @[Modules.scala 166:64:@44665.4]
  wire [13:0] buffer_13_483; // @[Modules.scala 166:64:@44666.4]
  wire [14:0] _T_96784; // @[Modules.scala 166:64:@44668.4]
  wire [13:0] _T_96785; // @[Modules.scala 166:64:@44669.4]
  wire [13:0] buffer_13_484; // @[Modules.scala 166:64:@44670.4]
  wire [14:0] _T_96787; // @[Modules.scala 166:64:@44672.4]
  wire [13:0] _T_96788; // @[Modules.scala 166:64:@44673.4]
  wire [13:0] buffer_13_485; // @[Modules.scala 166:64:@44674.4]
  wire [14:0] _T_96790; // @[Modules.scala 166:64:@44676.4]
  wire [13:0] _T_96791; // @[Modules.scala 166:64:@44677.4]
  wire [13:0] buffer_13_486; // @[Modules.scala 166:64:@44678.4]
  wire [14:0] _T_96793; // @[Modules.scala 166:64:@44680.4]
  wire [13:0] _T_96794; // @[Modules.scala 166:64:@44681.4]
  wire [13:0] buffer_13_487; // @[Modules.scala 166:64:@44682.4]
  wire [14:0] _T_96796; // @[Modules.scala 166:64:@44684.4]
  wire [13:0] _T_96797; // @[Modules.scala 166:64:@44685.4]
  wire [13:0] buffer_13_488; // @[Modules.scala 166:64:@44686.4]
  wire [14:0] _T_96799; // @[Modules.scala 166:64:@44688.4]
  wire [13:0] _T_96800; // @[Modules.scala 166:64:@44689.4]
  wire [13:0] buffer_13_489; // @[Modules.scala 166:64:@44690.4]
  wire [14:0] _T_96802; // @[Modules.scala 166:64:@44692.4]
  wire [13:0] _T_96803; // @[Modules.scala 166:64:@44693.4]
  wire [13:0] buffer_13_490; // @[Modules.scala 166:64:@44694.4]
  wire [14:0] _T_96805; // @[Modules.scala 166:64:@44696.4]
  wire [13:0] _T_96806; // @[Modules.scala 166:64:@44697.4]
  wire [13:0] buffer_13_491; // @[Modules.scala 166:64:@44698.4]
  wire [14:0] _T_96808; // @[Modules.scala 166:64:@44700.4]
  wire [13:0] _T_96809; // @[Modules.scala 166:64:@44701.4]
  wire [13:0] buffer_13_492; // @[Modules.scala 166:64:@44702.4]
  wire [14:0] _T_96811; // @[Modules.scala 166:64:@44704.4]
  wire [13:0] _T_96812; // @[Modules.scala 166:64:@44705.4]
  wire [13:0] buffer_13_493; // @[Modules.scala 166:64:@44706.4]
  wire [14:0] _T_96814; // @[Modules.scala 166:64:@44708.4]
  wire [13:0] _T_96815; // @[Modules.scala 166:64:@44709.4]
  wire [13:0] buffer_13_494; // @[Modules.scala 166:64:@44710.4]
  wire [14:0] _T_96817; // @[Modules.scala 166:64:@44712.4]
  wire [13:0] _T_96818; // @[Modules.scala 166:64:@44713.4]
  wire [13:0] buffer_13_495; // @[Modules.scala 166:64:@44714.4]
  wire [14:0] _T_96820; // @[Modules.scala 166:64:@44716.4]
  wire [13:0] _T_96821; // @[Modules.scala 166:64:@44717.4]
  wire [13:0] buffer_13_496; // @[Modules.scala 166:64:@44718.4]
  wire [14:0] _T_96823; // @[Modules.scala 166:64:@44720.4]
  wire [13:0] _T_96824; // @[Modules.scala 166:64:@44721.4]
  wire [13:0] buffer_13_497; // @[Modules.scala 166:64:@44722.4]
  wire [14:0] _T_96826; // @[Modules.scala 166:64:@44724.4]
  wire [13:0] _T_96827; // @[Modules.scala 166:64:@44725.4]
  wire [13:0] buffer_13_498; // @[Modules.scala 166:64:@44726.4]
  wire [14:0] _T_96829; // @[Modules.scala 166:64:@44728.4]
  wire [13:0] _T_96830; // @[Modules.scala 166:64:@44729.4]
  wire [13:0] buffer_13_499; // @[Modules.scala 166:64:@44730.4]
  wire [14:0] _T_96832; // @[Modules.scala 166:64:@44732.4]
  wire [13:0] _T_96833; // @[Modules.scala 166:64:@44733.4]
  wire [13:0] buffer_13_500; // @[Modules.scala 166:64:@44734.4]
  wire [14:0] _T_96835; // @[Modules.scala 166:64:@44736.4]
  wire [13:0] _T_96836; // @[Modules.scala 166:64:@44737.4]
  wire [13:0] buffer_13_501; // @[Modules.scala 166:64:@44738.4]
  wire [14:0] _T_96838; // @[Modules.scala 166:64:@44740.4]
  wire [13:0] _T_96839; // @[Modules.scala 166:64:@44741.4]
  wire [13:0] buffer_13_502; // @[Modules.scala 166:64:@44742.4]
  wire [14:0] _T_96841; // @[Modules.scala 166:64:@44744.4]
  wire [13:0] _T_96842; // @[Modules.scala 166:64:@44745.4]
  wire [13:0] buffer_13_503; // @[Modules.scala 166:64:@44746.4]
  wire [14:0] _T_96844; // @[Modules.scala 166:64:@44748.4]
  wire [13:0] _T_96845; // @[Modules.scala 166:64:@44749.4]
  wire [13:0] buffer_13_504; // @[Modules.scala 166:64:@44750.4]
  wire [14:0] _T_96847; // @[Modules.scala 166:64:@44752.4]
  wire [13:0] _T_96848; // @[Modules.scala 166:64:@44753.4]
  wire [13:0] buffer_13_505; // @[Modules.scala 166:64:@44754.4]
  wire [14:0] _T_96850; // @[Modules.scala 166:64:@44756.4]
  wire [13:0] _T_96851; // @[Modules.scala 166:64:@44757.4]
  wire [13:0] buffer_13_506; // @[Modules.scala 166:64:@44758.4]
  wire [14:0] _T_96853; // @[Modules.scala 166:64:@44760.4]
  wire [13:0] _T_96854; // @[Modules.scala 166:64:@44761.4]
  wire [13:0] buffer_13_507; // @[Modules.scala 166:64:@44762.4]
  wire [14:0] _T_96856; // @[Modules.scala 166:64:@44764.4]
  wire [13:0] _T_96857; // @[Modules.scala 166:64:@44765.4]
  wire [13:0] buffer_13_508; // @[Modules.scala 166:64:@44766.4]
  wire [14:0] _T_96859; // @[Modules.scala 166:64:@44768.4]
  wire [13:0] _T_96860; // @[Modules.scala 166:64:@44769.4]
  wire [13:0] buffer_13_509; // @[Modules.scala 166:64:@44770.4]
  wire [14:0] _T_96862; // @[Modules.scala 166:64:@44772.4]
  wire [13:0] _T_96863; // @[Modules.scala 166:64:@44773.4]
  wire [13:0] buffer_13_510; // @[Modules.scala 166:64:@44774.4]
  wire [14:0] _T_96865; // @[Modules.scala 166:64:@44776.4]
  wire [13:0] _T_96866; // @[Modules.scala 166:64:@44777.4]
  wire [13:0] buffer_13_511; // @[Modules.scala 166:64:@44778.4]
  wire [14:0] _T_96868; // @[Modules.scala 166:64:@44780.4]
  wire [13:0] _T_96869; // @[Modules.scala 166:64:@44781.4]
  wire [13:0] buffer_13_512; // @[Modules.scala 166:64:@44782.4]
  wire [14:0] _T_96871; // @[Modules.scala 166:64:@44784.4]
  wire [13:0] _T_96872; // @[Modules.scala 166:64:@44785.4]
  wire [13:0] buffer_13_513; // @[Modules.scala 166:64:@44786.4]
  wire [14:0] _T_96874; // @[Modules.scala 166:64:@44788.4]
  wire [13:0] _T_96875; // @[Modules.scala 166:64:@44789.4]
  wire [13:0] buffer_13_514; // @[Modules.scala 166:64:@44790.4]
  wire [14:0] _T_96877; // @[Modules.scala 166:64:@44792.4]
  wire [13:0] _T_96878; // @[Modules.scala 166:64:@44793.4]
  wire [13:0] buffer_13_515; // @[Modules.scala 166:64:@44794.4]
  wire [14:0] _T_96880; // @[Modules.scala 166:64:@44796.4]
  wire [13:0] _T_96881; // @[Modules.scala 166:64:@44797.4]
  wire [13:0] buffer_13_516; // @[Modules.scala 166:64:@44798.4]
  wire [14:0] _T_96883; // @[Modules.scala 166:64:@44800.4]
  wire [13:0] _T_96884; // @[Modules.scala 166:64:@44801.4]
  wire [13:0] buffer_13_517; // @[Modules.scala 166:64:@44802.4]
  wire [14:0] _T_96886; // @[Modules.scala 166:64:@44804.4]
  wire [13:0] _T_96887; // @[Modules.scala 166:64:@44805.4]
  wire [13:0] buffer_13_518; // @[Modules.scala 166:64:@44806.4]
  wire [14:0] _T_96889; // @[Modules.scala 166:64:@44808.4]
  wire [13:0] _T_96890; // @[Modules.scala 166:64:@44809.4]
  wire [13:0] buffer_13_519; // @[Modules.scala 166:64:@44810.4]
  wire [14:0] _T_96892; // @[Modules.scala 166:64:@44812.4]
  wire [13:0] _T_96893; // @[Modules.scala 166:64:@44813.4]
  wire [13:0] buffer_13_520; // @[Modules.scala 166:64:@44814.4]
  wire [14:0] _T_96895; // @[Modules.scala 166:64:@44816.4]
  wire [13:0] _T_96896; // @[Modules.scala 166:64:@44817.4]
  wire [13:0] buffer_13_521; // @[Modules.scala 166:64:@44818.4]
  wire [14:0] _T_96898; // @[Modules.scala 166:64:@44820.4]
  wire [13:0] _T_96899; // @[Modules.scala 166:64:@44821.4]
  wire [13:0] buffer_13_522; // @[Modules.scala 166:64:@44822.4]
  wire [14:0] _T_96901; // @[Modules.scala 166:64:@44824.4]
  wire [13:0] _T_96902; // @[Modules.scala 166:64:@44825.4]
  wire [13:0] buffer_13_523; // @[Modules.scala 166:64:@44826.4]
  wire [14:0] _T_96904; // @[Modules.scala 166:64:@44828.4]
  wire [13:0] _T_96905; // @[Modules.scala 166:64:@44829.4]
  wire [13:0] buffer_13_524; // @[Modules.scala 166:64:@44830.4]
  wire [14:0] _T_96907; // @[Modules.scala 166:64:@44832.4]
  wire [13:0] _T_96908; // @[Modules.scala 166:64:@44833.4]
  wire [13:0] buffer_13_525; // @[Modules.scala 166:64:@44834.4]
  wire [14:0] _T_96910; // @[Modules.scala 166:64:@44836.4]
  wire [13:0] _T_96911; // @[Modules.scala 166:64:@44837.4]
  wire [13:0] buffer_13_526; // @[Modules.scala 166:64:@44838.4]
  wire [14:0] _T_96913; // @[Modules.scala 166:64:@44840.4]
  wire [13:0] _T_96914; // @[Modules.scala 166:64:@44841.4]
  wire [13:0] buffer_13_527; // @[Modules.scala 166:64:@44842.4]
  wire [14:0] _T_96916; // @[Modules.scala 166:64:@44844.4]
  wire [13:0] _T_96917; // @[Modules.scala 166:64:@44845.4]
  wire [13:0] buffer_13_528; // @[Modules.scala 166:64:@44846.4]
  wire [14:0] _T_96919; // @[Modules.scala 166:64:@44848.4]
  wire [13:0] _T_96920; // @[Modules.scala 166:64:@44849.4]
  wire [13:0] buffer_13_529; // @[Modules.scala 166:64:@44850.4]
  wire [14:0] _T_96922; // @[Modules.scala 166:64:@44852.4]
  wire [13:0] _T_96923; // @[Modules.scala 166:64:@44853.4]
  wire [13:0] buffer_13_530; // @[Modules.scala 166:64:@44854.4]
  wire [14:0] _T_96928; // @[Modules.scala 166:64:@44860.4]
  wire [13:0] _T_96929; // @[Modules.scala 166:64:@44861.4]
  wire [13:0] buffer_13_532; // @[Modules.scala 166:64:@44862.4]
  wire [14:0] _T_96931; // @[Modules.scala 166:64:@44864.4]
  wire [13:0] _T_96932; // @[Modules.scala 166:64:@44865.4]
  wire [13:0] buffer_13_533; // @[Modules.scala 166:64:@44866.4]
  wire [14:0] _T_96934; // @[Modules.scala 166:64:@44868.4]
  wire [13:0] _T_96935; // @[Modules.scala 166:64:@44869.4]
  wire [13:0] buffer_13_534; // @[Modules.scala 166:64:@44870.4]
  wire [14:0] _T_96937; // @[Modules.scala 166:64:@44872.4]
  wire [13:0] _T_96938; // @[Modules.scala 166:64:@44873.4]
  wire [13:0] buffer_13_535; // @[Modules.scala 166:64:@44874.4]
  wire [14:0] _T_96940; // @[Modules.scala 172:66:@44876.4]
  wire [13:0] _T_96941; // @[Modules.scala 172:66:@44877.4]
  wire [13:0] buffer_13_536; // @[Modules.scala 172:66:@44878.4]
  wire [14:0] _T_96943; // @[Modules.scala 166:64:@44880.4]
  wire [13:0] _T_96944; // @[Modules.scala 166:64:@44881.4]
  wire [13:0] buffer_13_537; // @[Modules.scala 166:64:@44882.4]
  wire [14:0] _T_96946; // @[Modules.scala 166:64:@44884.4]
  wire [13:0] _T_96947; // @[Modules.scala 166:64:@44885.4]
  wire [13:0] buffer_13_538; // @[Modules.scala 166:64:@44886.4]
  wire [14:0] _T_96949; // @[Modules.scala 166:64:@44888.4]
  wire [13:0] _T_96950; // @[Modules.scala 166:64:@44889.4]
  wire [13:0] buffer_13_539; // @[Modules.scala 166:64:@44890.4]
  wire [14:0] _T_96955; // @[Modules.scala 166:64:@44896.4]
  wire [13:0] _T_96956; // @[Modules.scala 166:64:@44897.4]
  wire [13:0] buffer_13_541; // @[Modules.scala 166:64:@44898.4]
  wire [14:0] _T_96958; // @[Modules.scala 166:64:@44900.4]
  wire [13:0] _T_96959; // @[Modules.scala 166:64:@44901.4]
  wire [13:0] buffer_13_542; // @[Modules.scala 166:64:@44902.4]
  wire [14:0] _T_96961; // @[Modules.scala 166:64:@44904.4]
  wire [13:0] _T_96962; // @[Modules.scala 166:64:@44905.4]
  wire [13:0] buffer_13_543; // @[Modules.scala 166:64:@44906.4]
  wire [14:0] _T_96964; // @[Modules.scala 166:64:@44908.4]
  wire [13:0] _T_96965; // @[Modules.scala 166:64:@44909.4]
  wire [13:0] buffer_13_544; // @[Modules.scala 166:64:@44910.4]
  wire [14:0] _T_96967; // @[Modules.scala 166:64:@44912.4]
  wire [13:0] _T_96968; // @[Modules.scala 166:64:@44913.4]
  wire [13:0] buffer_13_545; // @[Modules.scala 166:64:@44914.4]
  wire [14:0] _T_96970; // @[Modules.scala 166:64:@44916.4]
  wire [13:0] _T_96971; // @[Modules.scala 166:64:@44917.4]
  wire [13:0] buffer_13_546; // @[Modules.scala 166:64:@44918.4]
  wire [14:0] _T_96973; // @[Modules.scala 166:64:@44920.4]
  wire [13:0] _T_96974; // @[Modules.scala 166:64:@44921.4]
  wire [13:0] buffer_13_547; // @[Modules.scala 166:64:@44922.4]
  wire [14:0] _T_96976; // @[Modules.scala 166:64:@44924.4]
  wire [13:0] _T_96977; // @[Modules.scala 166:64:@44925.4]
  wire [13:0] buffer_13_548; // @[Modules.scala 166:64:@44926.4]
  wire [14:0] _T_96979; // @[Modules.scala 166:64:@44928.4]
  wire [13:0] _T_96980; // @[Modules.scala 166:64:@44929.4]
  wire [13:0] buffer_13_549; // @[Modules.scala 166:64:@44930.4]
  wire [14:0] _T_96982; // @[Modules.scala 166:64:@44932.4]
  wire [13:0] _T_96983; // @[Modules.scala 166:64:@44933.4]
  wire [13:0] buffer_13_550; // @[Modules.scala 166:64:@44934.4]
  wire [14:0] _T_96985; // @[Modules.scala 166:64:@44936.4]
  wire [13:0] _T_96986; // @[Modules.scala 166:64:@44937.4]
  wire [13:0] buffer_13_551; // @[Modules.scala 166:64:@44938.4]
  wire [14:0] _T_96988; // @[Modules.scala 166:64:@44940.4]
  wire [13:0] _T_96989; // @[Modules.scala 166:64:@44941.4]
  wire [13:0] buffer_13_552; // @[Modules.scala 166:64:@44942.4]
  wire [14:0] _T_96991; // @[Modules.scala 166:64:@44944.4]
  wire [13:0] _T_96992; // @[Modules.scala 166:64:@44945.4]
  wire [13:0] buffer_13_553; // @[Modules.scala 166:64:@44946.4]
  wire [14:0] _T_96994; // @[Modules.scala 166:64:@44948.4]
  wire [13:0] _T_96995; // @[Modules.scala 166:64:@44949.4]
  wire [13:0] buffer_13_554; // @[Modules.scala 166:64:@44950.4]
  wire [14:0] _T_96997; // @[Modules.scala 166:64:@44952.4]
  wire [13:0] _T_96998; // @[Modules.scala 166:64:@44953.4]
  wire [13:0] buffer_13_555; // @[Modules.scala 166:64:@44954.4]
  wire [14:0] _T_97000; // @[Modules.scala 166:64:@44956.4]
  wire [13:0] _T_97001; // @[Modules.scala 166:64:@44957.4]
  wire [13:0] buffer_13_556; // @[Modules.scala 166:64:@44958.4]
  wire [14:0] _T_97003; // @[Modules.scala 166:64:@44960.4]
  wire [13:0] _T_97004; // @[Modules.scala 166:64:@44961.4]
  wire [13:0] buffer_13_557; // @[Modules.scala 166:64:@44962.4]
  wire [14:0] _T_97006; // @[Modules.scala 166:64:@44964.4]
  wire [13:0] _T_97007; // @[Modules.scala 166:64:@44965.4]
  wire [13:0] buffer_13_558; // @[Modules.scala 166:64:@44966.4]
  wire [14:0] _T_97009; // @[Modules.scala 166:64:@44968.4]
  wire [13:0] _T_97010; // @[Modules.scala 166:64:@44969.4]
  wire [13:0] buffer_13_559; // @[Modules.scala 166:64:@44970.4]
  wire [14:0] _T_97012; // @[Modules.scala 166:64:@44972.4]
  wire [13:0] _T_97013; // @[Modules.scala 166:64:@44973.4]
  wire [13:0] buffer_13_560; // @[Modules.scala 166:64:@44974.4]
  wire [14:0] _T_97015; // @[Modules.scala 166:64:@44976.4]
  wire [13:0] _T_97016; // @[Modules.scala 166:64:@44977.4]
  wire [13:0] buffer_13_561; // @[Modules.scala 166:64:@44978.4]
  wire [14:0] _T_97018; // @[Modules.scala 166:64:@44980.4]
  wire [13:0] _T_97019; // @[Modules.scala 166:64:@44981.4]
  wire [13:0] buffer_13_562; // @[Modules.scala 166:64:@44982.4]
  wire [14:0] _T_97021; // @[Modules.scala 166:64:@44984.4]
  wire [13:0] _T_97022; // @[Modules.scala 166:64:@44985.4]
  wire [13:0] buffer_13_563; // @[Modules.scala 166:64:@44986.4]
  wire [14:0] _T_97024; // @[Modules.scala 166:64:@44988.4]
  wire [13:0] _T_97025; // @[Modules.scala 166:64:@44989.4]
  wire [13:0] buffer_13_564; // @[Modules.scala 166:64:@44990.4]
  wire [14:0] _T_97027; // @[Modules.scala 166:64:@44992.4]
  wire [13:0] _T_97028; // @[Modules.scala 166:64:@44993.4]
  wire [13:0] buffer_13_565; // @[Modules.scala 166:64:@44994.4]
  wire [14:0] _T_97030; // @[Modules.scala 166:64:@44996.4]
  wire [13:0] _T_97031; // @[Modules.scala 166:64:@44997.4]
  wire [13:0] buffer_13_566; // @[Modules.scala 166:64:@44998.4]
  wire [14:0] _T_97033; // @[Modules.scala 166:64:@45000.4]
  wire [13:0] _T_97034; // @[Modules.scala 166:64:@45001.4]
  wire [13:0] buffer_13_567; // @[Modules.scala 166:64:@45002.4]
  wire [14:0] _T_97036; // @[Modules.scala 166:64:@45004.4]
  wire [13:0] _T_97037; // @[Modules.scala 166:64:@45005.4]
  wire [13:0] buffer_13_568; // @[Modules.scala 166:64:@45006.4]
  wire [14:0] _T_97039; // @[Modules.scala 166:64:@45008.4]
  wire [13:0] _T_97040; // @[Modules.scala 166:64:@45009.4]
  wire [13:0] buffer_13_569; // @[Modules.scala 166:64:@45010.4]
  wire [14:0] _T_97042; // @[Modules.scala 166:64:@45012.4]
  wire [13:0] _T_97043; // @[Modules.scala 166:64:@45013.4]
  wire [13:0] buffer_13_570; // @[Modules.scala 166:64:@45014.4]
  wire [14:0] _T_97045; // @[Modules.scala 166:64:@45016.4]
  wire [13:0] _T_97046; // @[Modules.scala 166:64:@45017.4]
  wire [13:0] buffer_13_571; // @[Modules.scala 166:64:@45018.4]
  wire [14:0] _T_97048; // @[Modules.scala 166:64:@45020.4]
  wire [13:0] _T_97049; // @[Modules.scala 166:64:@45021.4]
  wire [13:0] buffer_13_572; // @[Modules.scala 166:64:@45022.4]
  wire [14:0] _T_97051; // @[Modules.scala 166:64:@45024.4]
  wire [13:0] _T_97052; // @[Modules.scala 166:64:@45025.4]
  wire [13:0] buffer_13_573; // @[Modules.scala 166:64:@45026.4]
  wire [14:0] _T_97054; // @[Modules.scala 166:64:@45028.4]
  wire [13:0] _T_97055; // @[Modules.scala 166:64:@45029.4]
  wire [13:0] buffer_13_574; // @[Modules.scala 166:64:@45030.4]
  wire [14:0] _T_97057; // @[Modules.scala 160:64:@45032.4]
  wire [13:0] _T_97058; // @[Modules.scala 160:64:@45033.4]
  wire [13:0] buffer_13_575; // @[Modules.scala 160:64:@45034.4]
  wire [14:0] _T_97060; // @[Modules.scala 160:64:@45036.4]
  wire [13:0] _T_97061; // @[Modules.scala 160:64:@45037.4]
  wire [13:0] buffer_13_576; // @[Modules.scala 160:64:@45038.4]
  wire [14:0] _T_97063; // @[Modules.scala 160:64:@45040.4]
  wire [13:0] _T_97064; // @[Modules.scala 160:64:@45041.4]
  wire [13:0] buffer_13_577; // @[Modules.scala 160:64:@45042.4]
  wire [14:0] _T_97066; // @[Modules.scala 160:64:@45044.4]
  wire [13:0] _T_97067; // @[Modules.scala 160:64:@45045.4]
  wire [13:0] buffer_13_578; // @[Modules.scala 160:64:@45046.4]
  wire [14:0] _T_97069; // @[Modules.scala 160:64:@45048.4]
  wire [13:0] _T_97070; // @[Modules.scala 160:64:@45049.4]
  wire [13:0] buffer_13_579; // @[Modules.scala 160:64:@45050.4]
  wire [14:0] _T_97072; // @[Modules.scala 160:64:@45052.4]
  wire [13:0] _T_97073; // @[Modules.scala 160:64:@45053.4]
  wire [13:0] buffer_13_580; // @[Modules.scala 160:64:@45054.4]
  wire [14:0] _T_97075; // @[Modules.scala 160:64:@45056.4]
  wire [13:0] _T_97076; // @[Modules.scala 160:64:@45057.4]
  wire [13:0] buffer_13_581; // @[Modules.scala 160:64:@45058.4]
  wire [14:0] _T_97078; // @[Modules.scala 160:64:@45060.4]
  wire [13:0] _T_97079; // @[Modules.scala 160:64:@45061.4]
  wire [13:0] buffer_13_582; // @[Modules.scala 160:64:@45062.4]
  wire [14:0] _T_97081; // @[Modules.scala 160:64:@45064.4]
  wire [13:0] _T_97082; // @[Modules.scala 160:64:@45065.4]
  wire [13:0] buffer_13_583; // @[Modules.scala 160:64:@45066.4]
  wire [14:0] _T_97084; // @[Modules.scala 160:64:@45068.4]
  wire [13:0] _T_97085; // @[Modules.scala 160:64:@45069.4]
  wire [13:0] buffer_13_584; // @[Modules.scala 160:64:@45070.4]
  wire [14:0] _T_97087; // @[Modules.scala 160:64:@45072.4]
  wire [13:0] _T_97088; // @[Modules.scala 160:64:@45073.4]
  wire [13:0] buffer_13_585; // @[Modules.scala 160:64:@45074.4]
  wire [14:0] _T_97090; // @[Modules.scala 160:64:@45076.4]
  wire [13:0] _T_97091; // @[Modules.scala 160:64:@45077.4]
  wire [13:0] buffer_13_586; // @[Modules.scala 160:64:@45078.4]
  wire [14:0] _T_97093; // @[Modules.scala 160:64:@45080.4]
  wire [13:0] _T_97094; // @[Modules.scala 160:64:@45081.4]
  wire [13:0] buffer_13_587; // @[Modules.scala 160:64:@45082.4]
  wire [14:0] _T_97096; // @[Modules.scala 160:64:@45084.4]
  wire [13:0] _T_97097; // @[Modules.scala 160:64:@45085.4]
  wire [13:0] buffer_13_588; // @[Modules.scala 160:64:@45086.4]
  wire [14:0] _T_97099; // @[Modules.scala 160:64:@45088.4]
  wire [13:0] _T_97100; // @[Modules.scala 160:64:@45089.4]
  wire [13:0] buffer_13_589; // @[Modules.scala 160:64:@45090.4]
  wire [14:0] _T_97102; // @[Modules.scala 160:64:@45092.4]
  wire [13:0] _T_97103; // @[Modules.scala 160:64:@45093.4]
  wire [13:0] buffer_13_590; // @[Modules.scala 160:64:@45094.4]
  wire [14:0] _T_97105; // @[Modules.scala 160:64:@45096.4]
  wire [13:0] _T_97106; // @[Modules.scala 160:64:@45097.4]
  wire [13:0] buffer_13_591; // @[Modules.scala 160:64:@45098.4]
  wire [14:0] _T_97108; // @[Modules.scala 160:64:@45100.4]
  wire [13:0] _T_97109; // @[Modules.scala 160:64:@45101.4]
  wire [13:0] buffer_13_592; // @[Modules.scala 160:64:@45102.4]
  wire [14:0] _T_97111; // @[Modules.scala 160:64:@45104.4]
  wire [13:0] _T_97112; // @[Modules.scala 160:64:@45105.4]
  wire [13:0] buffer_13_593; // @[Modules.scala 160:64:@45106.4]
  wire [14:0] _T_97114; // @[Modules.scala 166:64:@45108.4]
  wire [13:0] _T_97115; // @[Modules.scala 166:64:@45109.4]
  wire [13:0] buffer_13_594; // @[Modules.scala 166:64:@45110.4]
  wire [14:0] _T_97117; // @[Modules.scala 166:64:@45112.4]
  wire [13:0] _T_97118; // @[Modules.scala 166:64:@45113.4]
  wire [13:0] buffer_13_595; // @[Modules.scala 166:64:@45114.4]
  wire [14:0] _T_97120; // @[Modules.scala 166:64:@45116.4]
  wire [13:0] _T_97121; // @[Modules.scala 166:64:@45117.4]
  wire [13:0] buffer_13_596; // @[Modules.scala 166:64:@45118.4]
  wire [14:0] _T_97123; // @[Modules.scala 166:64:@45120.4]
  wire [13:0] _T_97124; // @[Modules.scala 166:64:@45121.4]
  wire [13:0] buffer_13_597; // @[Modules.scala 166:64:@45122.4]
  wire [14:0] _T_97126; // @[Modules.scala 166:64:@45124.4]
  wire [13:0] _T_97127; // @[Modules.scala 166:64:@45125.4]
  wire [13:0] buffer_13_598; // @[Modules.scala 166:64:@45126.4]
  wire [14:0] _T_97129; // @[Modules.scala 166:64:@45128.4]
  wire [13:0] _T_97130; // @[Modules.scala 166:64:@45129.4]
  wire [13:0] buffer_13_599; // @[Modules.scala 166:64:@45130.4]
  wire [14:0] _T_97132; // @[Modules.scala 166:64:@45132.4]
  wire [13:0] _T_97133; // @[Modules.scala 166:64:@45133.4]
  wire [13:0] buffer_13_600; // @[Modules.scala 166:64:@45134.4]
  wire [14:0] _T_97135; // @[Modules.scala 166:64:@45136.4]
  wire [13:0] _T_97136; // @[Modules.scala 166:64:@45137.4]
  wire [13:0] buffer_13_601; // @[Modules.scala 166:64:@45138.4]
  wire [14:0] _T_97138; // @[Modules.scala 166:64:@45140.4]
  wire [13:0] _T_97139; // @[Modules.scala 166:64:@45141.4]
  wire [13:0] buffer_13_602; // @[Modules.scala 166:64:@45142.4]
  wire [14:0] _T_97141; // @[Modules.scala 172:66:@45144.4]
  wire [13:0] _T_97142; // @[Modules.scala 172:66:@45145.4]
  wire [13:0] buffer_13_603; // @[Modules.scala 172:66:@45146.4]
  wire [14:0] _T_97144; // @[Modules.scala 160:64:@45148.4]
  wire [13:0] _T_97145; // @[Modules.scala 160:64:@45149.4]
  wire [13:0] buffer_13_604; // @[Modules.scala 160:64:@45150.4]
  wire [14:0] _T_97147; // @[Modules.scala 160:64:@45152.4]
  wire [13:0] _T_97148; // @[Modules.scala 160:64:@45153.4]
  wire [13:0] buffer_13_605; // @[Modules.scala 160:64:@45154.4]
  wire [14:0] _T_97150; // @[Modules.scala 160:64:@45156.4]
  wire [13:0] _T_97151; // @[Modules.scala 160:64:@45157.4]
  wire [13:0] buffer_13_606; // @[Modules.scala 160:64:@45158.4]
  wire [14:0] _T_97153; // @[Modules.scala 160:64:@45160.4]
  wire [13:0] _T_97154; // @[Modules.scala 160:64:@45161.4]
  wire [13:0] buffer_13_607; // @[Modules.scala 160:64:@45162.4]
  wire [14:0] _T_97156; // @[Modules.scala 160:64:@45164.4]
  wire [13:0] _T_97157; // @[Modules.scala 160:64:@45165.4]
  wire [13:0] buffer_13_608; // @[Modules.scala 160:64:@45166.4]
  wire [14:0] _T_97159; // @[Modules.scala 166:64:@45168.4]
  wire [13:0] _T_97160; // @[Modules.scala 166:64:@45169.4]
  wire [13:0] buffer_13_609; // @[Modules.scala 166:64:@45170.4]
  wire [14:0] _T_97162; // @[Modules.scala 166:64:@45172.4]
  wire [13:0] _T_97163; // @[Modules.scala 166:64:@45173.4]
  wire [13:0] buffer_13_610; // @[Modules.scala 166:64:@45174.4]
  wire [14:0] _T_97165; // @[Modules.scala 160:64:@45176.4]
  wire [13:0] _T_97166; // @[Modules.scala 160:64:@45177.4]
  wire [13:0] buffer_13_611; // @[Modules.scala 160:64:@45178.4]
  wire [14:0] _T_97168; // @[Modules.scala 172:66:@45180.4]
  wire [13:0] _T_97169; // @[Modules.scala 172:66:@45181.4]
  wire [13:0] buffer_13_612; // @[Modules.scala 172:66:@45182.4]
  wire [5:0] _GEN_976; // @[Modules.scala 143:103:@45363.4]
  wire [6:0] _T_97182; // @[Modules.scala 143:103:@45363.4]
  wire [5:0] _T_97183; // @[Modules.scala 143:103:@45364.4]
  wire [5:0] _T_97184; // @[Modules.scala 143:103:@45365.4]
  wire [5:0] _GEN_977; // @[Modules.scala 143:103:@45429.4]
  wire [6:0] _T_97259; // @[Modules.scala 143:103:@45429.4]
  wire [5:0] _T_97260; // @[Modules.scala 143:103:@45430.4]
  wire [5:0] _T_97261; // @[Modules.scala 143:103:@45431.4]
  wire [6:0] _T_97273; // @[Modules.scala 143:103:@45441.4]
  wire [5:0] _T_97274; // @[Modules.scala 143:103:@45442.4]
  wire [5:0] _T_97275; // @[Modules.scala 143:103:@45443.4]
  wire [6:0] _T_97280; // @[Modules.scala 143:103:@45447.4]
  wire [5:0] _T_97281; // @[Modules.scala 143:103:@45448.4]
  wire [5:0] _T_97282; // @[Modules.scala 143:103:@45449.4]
  wire [6:0] _T_97287; // @[Modules.scala 143:103:@45453.4]
  wire [5:0] _T_97288; // @[Modules.scala 143:103:@45454.4]
  wire [5:0] _T_97289; // @[Modules.scala 143:103:@45455.4]
  wire [6:0] _T_97294; // @[Modules.scala 143:103:@45459.4]
  wire [5:0] _T_97295; // @[Modules.scala 143:103:@45460.4]
  wire [5:0] _T_97296; // @[Modules.scala 143:103:@45461.4]
  wire [6:0] _T_97301; // @[Modules.scala 143:103:@45465.4]
  wire [5:0] _T_97302; // @[Modules.scala 143:103:@45466.4]
  wire [5:0] _T_97303; // @[Modules.scala 143:103:@45467.4]
  wire [6:0] _T_97308; // @[Modules.scala 143:103:@45471.4]
  wire [5:0] _T_97309; // @[Modules.scala 143:103:@45472.4]
  wire [5:0] _T_97310; // @[Modules.scala 143:103:@45473.4]
  wire [5:0] _GEN_978; // @[Modules.scala 143:103:@45501.4]
  wire [6:0] _T_97343; // @[Modules.scala 143:103:@45501.4]
  wire [5:0] _T_97344; // @[Modules.scala 143:103:@45502.4]
  wire [5:0] _T_97345; // @[Modules.scala 143:103:@45503.4]
  wire [5:0] _GEN_979; // @[Modules.scala 143:103:@45507.4]
  wire [6:0] _T_97350; // @[Modules.scala 143:103:@45507.4]
  wire [5:0] _T_97351; // @[Modules.scala 143:103:@45508.4]
  wire [5:0] _T_97352; // @[Modules.scala 143:103:@45509.4]
  wire [6:0] _T_97420; // @[Modules.scala 143:103:@45567.4]
  wire [5:0] _T_97421; // @[Modules.scala 143:103:@45568.4]
  wire [5:0] _T_97422; // @[Modules.scala 143:103:@45569.4]
  wire [5:0] _T_97441; // @[Modules.scala 143:103:@45585.4]
  wire [4:0] _T_97442; // @[Modules.scala 143:103:@45586.4]
  wire [4:0] _T_97443; // @[Modules.scala 143:103:@45587.4]
  wire [6:0] _T_97469; // @[Modules.scala 143:103:@45609.4]
  wire [5:0] _T_97470; // @[Modules.scala 143:103:@45610.4]
  wire [5:0] _T_97471; // @[Modules.scala 143:103:@45611.4]
  wire [5:0] _T_97476; // @[Modules.scala 143:103:@45615.4]
  wire [4:0] _T_97477; // @[Modules.scala 143:103:@45616.4]
  wire [4:0] _T_97478; // @[Modules.scala 143:103:@45617.4]
  wire [6:0] _T_97483; // @[Modules.scala 143:103:@45621.4]
  wire [5:0] _T_97484; // @[Modules.scala 143:103:@45622.4]
  wire [5:0] _T_97485; // @[Modules.scala 143:103:@45623.4]
  wire [6:0] _T_97518; // @[Modules.scala 143:103:@45651.4]
  wire [5:0] _T_97519; // @[Modules.scala 143:103:@45652.4]
  wire [5:0] _T_97520; // @[Modules.scala 143:103:@45653.4]
  wire [5:0] _GEN_990; // @[Modules.scala 143:103:@45705.4]
  wire [6:0] _T_97581; // @[Modules.scala 143:103:@45705.4]
  wire [5:0] _T_97582; // @[Modules.scala 143:103:@45706.4]
  wire [5:0] _T_97583; // @[Modules.scala 143:103:@45707.4]
  wire [5:0] _GEN_991; // @[Modules.scala 143:103:@45717.4]
  wire [6:0] _T_97595; // @[Modules.scala 143:103:@45717.4]
  wire [5:0] _T_97596; // @[Modules.scala 143:103:@45718.4]
  wire [5:0] _T_97597; // @[Modules.scala 143:103:@45719.4]
  wire [6:0] _T_97623; // @[Modules.scala 143:103:@45741.4]
  wire [5:0] _T_97624; // @[Modules.scala 143:103:@45742.4]
  wire [5:0] _T_97625; // @[Modules.scala 143:103:@45743.4]
  wire [6:0] _T_97630; // @[Modules.scala 143:103:@45747.4]
  wire [5:0] _T_97631; // @[Modules.scala 143:103:@45748.4]
  wire [5:0] _T_97632; // @[Modules.scala 143:103:@45749.4]
  wire [6:0] _T_97651; // @[Modules.scala 143:103:@45765.4]
  wire [5:0] _T_97652; // @[Modules.scala 143:103:@45766.4]
  wire [5:0] _T_97653; // @[Modules.scala 143:103:@45767.4]
  wire [6:0] _T_97658; // @[Modules.scala 143:103:@45771.4]
  wire [5:0] _T_97659; // @[Modules.scala 143:103:@45772.4]
  wire [5:0] _T_97660; // @[Modules.scala 143:103:@45773.4]
  wire [6:0] _T_97672; // @[Modules.scala 143:103:@45783.4]
  wire [5:0] _T_97673; // @[Modules.scala 143:103:@45784.4]
  wire [5:0] _T_97674; // @[Modules.scala 143:103:@45785.4]
  wire [6:0] _T_97686; // @[Modules.scala 143:103:@45795.4]
  wire [5:0] _T_97687; // @[Modules.scala 143:103:@45796.4]
  wire [5:0] _T_97688; // @[Modules.scala 143:103:@45797.4]
  wire [5:0] _GEN_997; // @[Modules.scala 143:103:@45807.4]
  wire [6:0] _T_97700; // @[Modules.scala 143:103:@45807.4]
  wire [5:0] _T_97701; // @[Modules.scala 143:103:@45808.4]
  wire [5:0] _T_97702; // @[Modules.scala 143:103:@45809.4]
  wire [6:0] _T_97721; // @[Modules.scala 143:103:@45825.4]
  wire [5:0] _T_97722; // @[Modules.scala 143:103:@45826.4]
  wire [5:0] _T_97723; // @[Modules.scala 143:103:@45827.4]
  wire [5:0] _GEN_999; // @[Modules.scala 143:103:@45831.4]
  wire [6:0] _T_97728; // @[Modules.scala 143:103:@45831.4]
  wire [5:0] _T_97729; // @[Modules.scala 143:103:@45832.4]
  wire [5:0] _T_97730; // @[Modules.scala 143:103:@45833.4]
  wire [5:0] _GEN_1000; // @[Modules.scala 143:103:@45879.4]
  wire [6:0] _T_97784; // @[Modules.scala 143:103:@45879.4]
  wire [5:0] _T_97785; // @[Modules.scala 143:103:@45880.4]
  wire [5:0] _T_97786; // @[Modules.scala 143:103:@45881.4]
  wire [5:0] _GEN_1001; // @[Modules.scala 143:103:@45885.4]
  wire [6:0] _T_97791; // @[Modules.scala 143:103:@45885.4]
  wire [5:0] _T_97792; // @[Modules.scala 143:103:@45886.4]
  wire [5:0] _T_97793; // @[Modules.scala 143:103:@45887.4]
  wire [5:0] _GEN_1002; // @[Modules.scala 143:103:@45909.4]
  wire [6:0] _T_97819; // @[Modules.scala 143:103:@45909.4]
  wire [5:0] _T_97820; // @[Modules.scala 143:103:@45910.4]
  wire [5:0] _T_97821; // @[Modules.scala 143:103:@45911.4]
  wire [5:0] _T_97847; // @[Modules.scala 143:103:@45933.4]
  wire [4:0] _T_97848; // @[Modules.scala 143:103:@45934.4]
  wire [4:0] _T_97849; // @[Modules.scala 143:103:@45935.4]
  wire [6:0] _T_97854; // @[Modules.scala 143:103:@45939.4]
  wire [5:0] _T_97855; // @[Modules.scala 143:103:@45940.4]
  wire [5:0] _T_97856; // @[Modules.scala 143:103:@45941.4]
  wire [5:0] _T_97861; // @[Modules.scala 143:103:@45945.4]
  wire [4:0] _T_97862; // @[Modules.scala 143:103:@45946.4]
  wire [4:0] _T_97863; // @[Modules.scala 143:103:@45947.4]
  wire [5:0] _T_97882; // @[Modules.scala 143:103:@45963.4]
  wire [4:0] _T_97883; // @[Modules.scala 143:103:@45964.4]
  wire [4:0] _T_97884; // @[Modules.scala 143:103:@45965.4]
  wire [5:0] _T_97910; // @[Modules.scala 143:103:@45987.4]
  wire [4:0] _T_97911; // @[Modules.scala 143:103:@45988.4]
  wire [4:0] _T_97912; // @[Modules.scala 143:103:@45989.4]
  wire [6:0] _T_97931; // @[Modules.scala 143:103:@46005.4]
  wire [5:0] _T_97932; // @[Modules.scala 143:103:@46006.4]
  wire [5:0] _T_97933; // @[Modules.scala 143:103:@46007.4]
  wire [5:0] _GEN_1006; // @[Modules.scala 143:103:@46029.4]
  wire [6:0] _T_97959; // @[Modules.scala 143:103:@46029.4]
  wire [5:0] _T_97960; // @[Modules.scala 143:103:@46030.4]
  wire [5:0] _T_97961; // @[Modules.scala 143:103:@46031.4]
  wire [6:0] _T_97987; // @[Modules.scala 143:103:@46053.4]
  wire [5:0] _T_97988; // @[Modules.scala 143:103:@46054.4]
  wire [5:0] _T_97989; // @[Modules.scala 143:103:@46055.4]
  wire [5:0] _GEN_1008; // @[Modules.scala 143:103:@46077.4]
  wire [6:0] _T_98015; // @[Modules.scala 143:103:@46077.4]
  wire [5:0] _T_98016; // @[Modules.scala 143:103:@46078.4]
  wire [5:0] _T_98017; // @[Modules.scala 143:103:@46079.4]
  wire [5:0] _T_98057; // @[Modules.scala 143:103:@46113.4]
  wire [4:0] _T_98058; // @[Modules.scala 143:103:@46114.4]
  wire [4:0] _T_98059; // @[Modules.scala 143:103:@46115.4]
  wire [5:0] _T_98085; // @[Modules.scala 143:103:@46137.4]
  wire [4:0] _T_98086; // @[Modules.scala 143:103:@46138.4]
  wire [4:0] _T_98087; // @[Modules.scala 143:103:@46139.4]
  wire [6:0] _T_98092; // @[Modules.scala 143:103:@46143.4]
  wire [5:0] _T_98093; // @[Modules.scala 143:103:@46144.4]
  wire [5:0] _T_98094; // @[Modules.scala 143:103:@46145.4]
  wire [6:0] _T_98099; // @[Modules.scala 143:103:@46149.4]
  wire [5:0] _T_98100; // @[Modules.scala 143:103:@46150.4]
  wire [5:0] _T_98101; // @[Modules.scala 143:103:@46151.4]
  wire [5:0] _T_98127; // @[Modules.scala 143:103:@46173.4]
  wire [4:0] _T_98128; // @[Modules.scala 143:103:@46174.4]
  wire [4:0] _T_98129; // @[Modules.scala 143:103:@46175.4]
  wire [5:0] _GEN_1013; // @[Modules.scala 143:103:@46197.4]
  wire [6:0] _T_98155; // @[Modules.scala 143:103:@46197.4]
  wire [5:0] _T_98156; // @[Modules.scala 143:103:@46198.4]
  wire [5:0] _T_98157; // @[Modules.scala 143:103:@46199.4]
  wire [5:0] _GEN_1014; // @[Modules.scala 143:103:@46209.4]
  wire [6:0] _T_98169; // @[Modules.scala 143:103:@46209.4]
  wire [5:0] _T_98170; // @[Modules.scala 143:103:@46210.4]
  wire [5:0] _T_98171; // @[Modules.scala 143:103:@46211.4]
  wire [5:0] _GEN_1015; // @[Modules.scala 143:103:@46215.4]
  wire [6:0] _T_98176; // @[Modules.scala 143:103:@46215.4]
  wire [5:0] _T_98177; // @[Modules.scala 143:103:@46216.4]
  wire [5:0] _T_98178; // @[Modules.scala 143:103:@46217.4]
  wire [6:0] _T_98183; // @[Modules.scala 143:103:@46221.4]
  wire [5:0] _T_98184; // @[Modules.scala 143:103:@46222.4]
  wire [5:0] _T_98185; // @[Modules.scala 143:103:@46223.4]
  wire [6:0] _T_98190; // @[Modules.scala 143:103:@46227.4]
  wire [5:0] _T_98191; // @[Modules.scala 143:103:@46228.4]
  wire [5:0] _T_98192; // @[Modules.scala 143:103:@46229.4]
  wire [5:0] _T_98211; // @[Modules.scala 143:103:@46245.4]
  wire [4:0] _T_98212; // @[Modules.scala 143:103:@46246.4]
  wire [4:0] _T_98213; // @[Modules.scala 143:103:@46247.4]
  wire [6:0] _T_98239; // @[Modules.scala 143:103:@46269.4]
  wire [5:0] _T_98240; // @[Modules.scala 143:103:@46270.4]
  wire [5:0] _T_98241; // @[Modules.scala 143:103:@46271.4]
  wire [6:0] _T_98260; // @[Modules.scala 143:103:@46287.4]
  wire [5:0] _T_98261; // @[Modules.scala 143:103:@46288.4]
  wire [5:0] _T_98262; // @[Modules.scala 143:103:@46289.4]
  wire [6:0] _T_98302; // @[Modules.scala 143:103:@46323.4]
  wire [5:0] _T_98303; // @[Modules.scala 143:103:@46324.4]
  wire [5:0] _T_98304; // @[Modules.scala 143:103:@46325.4]
  wire [6:0] _T_98309; // @[Modules.scala 143:103:@46329.4]
  wire [5:0] _T_98310; // @[Modules.scala 143:103:@46330.4]
  wire [5:0] _T_98311; // @[Modules.scala 143:103:@46331.4]
  wire [6:0] _T_98344; // @[Modules.scala 143:103:@46359.4]
  wire [5:0] _T_98345; // @[Modules.scala 143:103:@46360.4]
  wire [5:0] _T_98346; // @[Modules.scala 143:103:@46361.4]
  wire [6:0] _T_98358; // @[Modules.scala 143:103:@46371.4]
  wire [5:0] _T_98359; // @[Modules.scala 143:103:@46372.4]
  wire [5:0] _T_98360; // @[Modules.scala 143:103:@46373.4]
  wire [5:0] _T_98372; // @[Modules.scala 143:103:@46383.4]
  wire [4:0] _T_98373; // @[Modules.scala 143:103:@46384.4]
  wire [4:0] _T_98374; // @[Modules.scala 143:103:@46385.4]
  wire [5:0] _T_98393; // @[Modules.scala 143:103:@46401.4]
  wire [4:0] _T_98394; // @[Modules.scala 143:103:@46402.4]
  wire [4:0] _T_98395; // @[Modules.scala 143:103:@46403.4]
  wire [6:0] _T_98407; // @[Modules.scala 143:103:@46413.4]
  wire [5:0] _T_98408; // @[Modules.scala 143:103:@46414.4]
  wire [5:0] _T_98409; // @[Modules.scala 143:103:@46415.4]
  wire [6:0] _T_98421; // @[Modules.scala 143:103:@46425.4]
  wire [5:0] _T_98422; // @[Modules.scala 143:103:@46426.4]
  wire [5:0] _T_98423; // @[Modules.scala 143:103:@46427.4]
  wire [6:0] _T_98442; // @[Modules.scala 143:103:@46443.4]
  wire [5:0] _T_98443; // @[Modules.scala 143:103:@46444.4]
  wire [5:0] _T_98444; // @[Modules.scala 143:103:@46445.4]
  wire [6:0] _T_98449; // @[Modules.scala 143:103:@46449.4]
  wire [5:0] _T_98450; // @[Modules.scala 143:103:@46450.4]
  wire [5:0] _T_98451; // @[Modules.scala 143:103:@46451.4]
  wire [6:0] _T_98491; // @[Modules.scala 143:103:@46485.4]
  wire [5:0] _T_98492; // @[Modules.scala 143:103:@46486.4]
  wire [5:0] _T_98493; // @[Modules.scala 143:103:@46487.4]
  wire [6:0] _T_98498; // @[Modules.scala 143:103:@46491.4]
  wire [5:0] _T_98499; // @[Modules.scala 143:103:@46492.4]
  wire [5:0] _T_98500; // @[Modules.scala 143:103:@46493.4]
  wire [6:0] _T_98512; // @[Modules.scala 143:103:@46503.4]
  wire [5:0] _T_98513; // @[Modules.scala 143:103:@46504.4]
  wire [5:0] _T_98514; // @[Modules.scala 143:103:@46505.4]
  wire [6:0] _T_98533; // @[Modules.scala 143:103:@46521.4]
  wire [5:0] _T_98534; // @[Modules.scala 143:103:@46522.4]
  wire [5:0] _T_98535; // @[Modules.scala 143:103:@46523.4]
  wire [5:0] _GEN_1038; // @[Modules.scala 143:103:@46533.4]
  wire [6:0] _T_98547; // @[Modules.scala 143:103:@46533.4]
  wire [5:0] _T_98548; // @[Modules.scala 143:103:@46534.4]
  wire [5:0] _T_98549; // @[Modules.scala 143:103:@46535.4]
  wire [5:0] _GEN_1039; // @[Modules.scala 143:103:@46539.4]
  wire [6:0] _T_98554; // @[Modules.scala 143:103:@46539.4]
  wire [5:0] _T_98555; // @[Modules.scala 143:103:@46540.4]
  wire [5:0] _T_98556; // @[Modules.scala 143:103:@46541.4]
  wire [6:0] _T_98568; // @[Modules.scala 143:103:@46551.4]
  wire [5:0] _T_98569; // @[Modules.scala 143:103:@46552.4]
  wire [5:0] _T_98570; // @[Modules.scala 143:103:@46553.4]
  wire [6:0] _T_98610; // @[Modules.scala 143:103:@46587.4]
  wire [5:0] _T_98611; // @[Modules.scala 143:103:@46588.4]
  wire [5:0] _T_98612; // @[Modules.scala 143:103:@46589.4]
  wire [5:0] _T_98729; // @[Modules.scala 143:103:@46689.4]
  wire [4:0] _T_98730; // @[Modules.scala 143:103:@46690.4]
  wire [4:0] _T_98731; // @[Modules.scala 143:103:@46691.4]
  wire [6:0] _T_98743; // @[Modules.scala 143:103:@46701.4]
  wire [5:0] _T_98744; // @[Modules.scala 143:103:@46702.4]
  wire [5:0] _T_98745; // @[Modules.scala 143:103:@46703.4]
  wire [6:0] _T_98750; // @[Modules.scala 143:103:@46707.4]
  wire [5:0] _T_98751; // @[Modules.scala 143:103:@46708.4]
  wire [5:0] _T_98752; // @[Modules.scala 143:103:@46709.4]
  wire [6:0] _T_98757; // @[Modules.scala 143:103:@46713.4]
  wire [5:0] _T_98758; // @[Modules.scala 143:103:@46714.4]
  wire [5:0] _T_98759; // @[Modules.scala 143:103:@46715.4]
  wire [6:0] _T_98778; // @[Modules.scala 143:103:@46731.4]
  wire [5:0] _T_98779; // @[Modules.scala 143:103:@46732.4]
  wire [5:0] _T_98780; // @[Modules.scala 143:103:@46733.4]
  wire [5:0] _GEN_1045; // @[Modules.scala 143:103:@46743.4]
  wire [6:0] _T_98792; // @[Modules.scala 143:103:@46743.4]
  wire [5:0] _T_98793; // @[Modules.scala 143:103:@46744.4]
  wire [5:0] _T_98794; // @[Modules.scala 143:103:@46745.4]
  wire [6:0] _T_98799; // @[Modules.scala 143:103:@46749.4]
  wire [5:0] _T_98800; // @[Modules.scala 143:103:@46750.4]
  wire [5:0] _T_98801; // @[Modules.scala 143:103:@46751.4]
  wire [5:0] _T_98813; // @[Modules.scala 143:103:@46761.4]
  wire [4:0] _T_98814; // @[Modules.scala 143:103:@46762.4]
  wire [4:0] _T_98815; // @[Modules.scala 143:103:@46763.4]
  wire [6:0] _T_98834; // @[Modules.scala 143:103:@46779.4]
  wire [5:0] _T_98835; // @[Modules.scala 143:103:@46780.4]
  wire [5:0] _T_98836; // @[Modules.scala 143:103:@46781.4]
  wire [6:0] _T_98848; // @[Modules.scala 143:103:@46791.4]
  wire [5:0] _T_98849; // @[Modules.scala 143:103:@46792.4]
  wire [5:0] _T_98850; // @[Modules.scala 143:103:@46793.4]
  wire [6:0] _T_98855; // @[Modules.scala 143:103:@46797.4]
  wire [5:0] _T_98856; // @[Modules.scala 143:103:@46798.4]
  wire [5:0] _T_98857; // @[Modules.scala 143:103:@46799.4]
  wire [5:0] _GEN_1048; // @[Modules.scala 143:103:@46815.4]
  wire [6:0] _T_98876; // @[Modules.scala 143:103:@46815.4]
  wire [5:0] _T_98877; // @[Modules.scala 143:103:@46816.4]
  wire [5:0] _T_98878; // @[Modules.scala 143:103:@46817.4]
  wire [6:0] _T_98890; // @[Modules.scala 143:103:@46827.4]
  wire [5:0] _T_98891; // @[Modules.scala 143:103:@46828.4]
  wire [5:0] _T_98892; // @[Modules.scala 143:103:@46829.4]
  wire [6:0] _T_98925; // @[Modules.scala 143:103:@46857.4]
  wire [5:0] _T_98926; // @[Modules.scala 143:103:@46858.4]
  wire [5:0] _T_98927; // @[Modules.scala 143:103:@46859.4]
  wire [5:0] _GEN_1050; // @[Modules.scala 143:103:@46887.4]
  wire [6:0] _T_98960; // @[Modules.scala 143:103:@46887.4]
  wire [5:0] _T_98961; // @[Modules.scala 143:103:@46888.4]
  wire [5:0] _T_98962; // @[Modules.scala 143:103:@46889.4]
  wire [5:0] _GEN_1051; // @[Modules.scala 143:103:@46911.4]
  wire [6:0] _T_98988; // @[Modules.scala 143:103:@46911.4]
  wire [5:0] _T_98989; // @[Modules.scala 143:103:@46912.4]
  wire [5:0] _T_98990; // @[Modules.scala 143:103:@46913.4]
  wire [6:0] _T_99023; // @[Modules.scala 143:103:@46941.4]
  wire [5:0] _T_99024; // @[Modules.scala 143:103:@46942.4]
  wire [5:0] _T_99025; // @[Modules.scala 143:103:@46943.4]
  wire [5:0] _GEN_1053; // @[Modules.scala 143:103:@46947.4]
  wire [6:0] _T_99030; // @[Modules.scala 143:103:@46947.4]
  wire [5:0] _T_99031; // @[Modules.scala 143:103:@46948.4]
  wire [5:0] _T_99032; // @[Modules.scala 143:103:@46949.4]
  wire [5:0] _T_99044; // @[Modules.scala 143:103:@46959.4]
  wire [4:0] _T_99045; // @[Modules.scala 143:103:@46960.4]
  wire [4:0] _T_99046; // @[Modules.scala 143:103:@46961.4]
  wire [6:0] _T_99107; // @[Modules.scala 143:103:@47013.4]
  wire [5:0] _T_99108; // @[Modules.scala 143:103:@47014.4]
  wire [5:0] _T_99109; // @[Modules.scala 143:103:@47015.4]
  wire [6:0] _T_99128; // @[Modules.scala 143:103:@47031.4]
  wire [5:0] _T_99129; // @[Modules.scala 143:103:@47032.4]
  wire [5:0] _T_99130; // @[Modules.scala 143:103:@47033.4]
  wire [6:0] _T_99219; // @[Modules.scala 143:103:@47109.4]
  wire [5:0] _T_99220; // @[Modules.scala 143:103:@47110.4]
  wire [5:0] _T_99221; // @[Modules.scala 143:103:@47111.4]
  wire [6:0] _T_99233; // @[Modules.scala 143:103:@47121.4]
  wire [5:0] _T_99234; // @[Modules.scala 143:103:@47122.4]
  wire [5:0] _T_99235; // @[Modules.scala 143:103:@47123.4]
  wire [5:0] _GEN_1057; // @[Modules.scala 143:103:@47127.4]
  wire [6:0] _T_99240; // @[Modules.scala 143:103:@47127.4]
  wire [5:0] _T_99241; // @[Modules.scala 143:103:@47128.4]
  wire [5:0] _T_99242; // @[Modules.scala 143:103:@47129.4]
  wire [5:0] _T_99247; // @[Modules.scala 143:103:@47133.4]
  wire [4:0] _T_99248; // @[Modules.scala 143:103:@47134.4]
  wire [4:0] _T_99249; // @[Modules.scala 143:103:@47135.4]
  wire [5:0] _T_99275; // @[Modules.scala 143:103:@47157.4]
  wire [4:0] _T_99276; // @[Modules.scala 143:103:@47158.4]
  wire [4:0] _T_99277; // @[Modules.scala 143:103:@47159.4]
  wire [13:0] buffer_14_1; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99285; // @[Modules.scala 160:64:@47167.4]
  wire [13:0] _T_99286; // @[Modules.scala 160:64:@47168.4]
  wire [13:0] buffer_14_302; // @[Modules.scala 160:64:@47169.4]
  wire [14:0] _T_99288; // @[Modules.scala 160:64:@47171.4]
  wire [13:0] _T_99289; // @[Modules.scala 160:64:@47172.4]
  wire [13:0] buffer_14_303; // @[Modules.scala 160:64:@47173.4]
  wire [13:0] buffer_14_12; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99303; // @[Modules.scala 160:64:@47191.4]
  wire [13:0] _T_99304; // @[Modules.scala 160:64:@47192.4]
  wire [13:0] buffer_14_308; // @[Modules.scala 160:64:@47193.4]
  wire [13:0] buffer_14_14; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_15; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99306; // @[Modules.scala 160:64:@47195.4]
  wire [13:0] _T_99307; // @[Modules.scala 160:64:@47196.4]
  wire [13:0] buffer_14_309; // @[Modules.scala 160:64:@47197.4]
  wire [13:0] buffer_14_16; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_17; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99309; // @[Modules.scala 160:64:@47199.4]
  wire [13:0] _T_99310; // @[Modules.scala 160:64:@47200.4]
  wire [13:0] buffer_14_310; // @[Modules.scala 160:64:@47201.4]
  wire [13:0] buffer_14_18; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_19; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99312; // @[Modules.scala 160:64:@47203.4]
  wire [13:0] _T_99313; // @[Modules.scala 160:64:@47204.4]
  wire [13:0] buffer_14_311; // @[Modules.scala 160:64:@47205.4]
  wire [14:0] _T_99318; // @[Modules.scala 160:64:@47211.4]
  wire [13:0] _T_99319; // @[Modules.scala 160:64:@47212.4]
  wire [13:0] buffer_14_313; // @[Modules.scala 160:64:@47213.4]
  wire [13:0] buffer_14_24; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_25; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99321; // @[Modules.scala 160:64:@47215.4]
  wire [13:0] _T_99322; // @[Modules.scala 160:64:@47216.4]
  wire [13:0] buffer_14_314; // @[Modules.scala 160:64:@47217.4]
  wire [14:0] _T_99324; // @[Modules.scala 160:64:@47219.4]
  wire [13:0] _T_99325; // @[Modules.scala 160:64:@47220.4]
  wire [13:0] buffer_14_315; // @[Modules.scala 160:64:@47221.4]
  wire [14:0] _T_99327; // @[Modules.scala 160:64:@47223.4]
  wire [13:0] _T_99328; // @[Modules.scala 160:64:@47224.4]
  wire [13:0] buffer_14_316; // @[Modules.scala 160:64:@47225.4]
  wire [13:0] buffer_14_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99336; // @[Modules.scala 160:64:@47235.4]
  wire [13:0] _T_99337; // @[Modules.scala 160:64:@47236.4]
  wire [13:0] buffer_14_319; // @[Modules.scala 160:64:@47237.4]
  wire [14:0] _T_99339; // @[Modules.scala 160:64:@47239.4]
  wire [13:0] _T_99340; // @[Modules.scala 160:64:@47240.4]
  wire [13:0] buffer_14_320; // @[Modules.scala 160:64:@47241.4]
  wire [13:0] buffer_14_38; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99342; // @[Modules.scala 160:64:@47243.4]
  wire [13:0] _T_99343; // @[Modules.scala 160:64:@47244.4]
  wire [13:0] buffer_14_321; // @[Modules.scala 160:64:@47245.4]
  wire [14:0] _T_99345; // @[Modules.scala 160:64:@47247.4]
  wire [13:0] _T_99346; // @[Modules.scala 160:64:@47248.4]
  wire [13:0] buffer_14_322; // @[Modules.scala 160:64:@47249.4]
  wire [13:0] buffer_14_42; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_43; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99348; // @[Modules.scala 160:64:@47251.4]
  wire [13:0] _T_99349; // @[Modules.scala 160:64:@47252.4]
  wire [13:0] buffer_14_323; // @[Modules.scala 160:64:@47253.4]
  wire [13:0] buffer_14_44; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99351; // @[Modules.scala 160:64:@47255.4]
  wire [13:0] _T_99352; // @[Modules.scala 160:64:@47256.4]
  wire [13:0] buffer_14_324; // @[Modules.scala 160:64:@47257.4]
  wire [13:0] buffer_14_49; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99357; // @[Modules.scala 160:64:@47263.4]
  wire [13:0] _T_99358; // @[Modules.scala 160:64:@47264.4]
  wire [13:0] buffer_14_326; // @[Modules.scala 160:64:@47265.4]
  wire [14:0] _T_99366; // @[Modules.scala 160:64:@47275.4]
  wire [13:0] _T_99367; // @[Modules.scala 160:64:@47276.4]
  wire [13:0] buffer_14_329; // @[Modules.scala 160:64:@47277.4]
  wire [13:0] buffer_14_58; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99372; // @[Modules.scala 160:64:@47283.4]
  wire [13:0] _T_99373; // @[Modules.scala 160:64:@47284.4]
  wire [13:0] buffer_14_331; // @[Modules.scala 160:64:@47285.4]
  wire [13:0] buffer_14_60; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99375; // @[Modules.scala 160:64:@47287.4]
  wire [13:0] _T_99376; // @[Modules.scala 160:64:@47288.4]
  wire [13:0] buffer_14_332; // @[Modules.scala 160:64:@47289.4]
  wire [14:0] _T_99378; // @[Modules.scala 160:64:@47291.4]
  wire [13:0] _T_99379; // @[Modules.scala 160:64:@47292.4]
  wire [13:0] buffer_14_333; // @[Modules.scala 160:64:@47293.4]
  wire [13:0] buffer_14_64; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_65; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99381; // @[Modules.scala 160:64:@47295.4]
  wire [13:0] _T_99382; // @[Modules.scala 160:64:@47296.4]
  wire [13:0] buffer_14_334; // @[Modules.scala 160:64:@47297.4]
  wire [14:0] _T_99384; // @[Modules.scala 160:64:@47299.4]
  wire [13:0] _T_99385; // @[Modules.scala 160:64:@47300.4]
  wire [13:0] buffer_14_335; // @[Modules.scala 160:64:@47301.4]
  wire [13:0] buffer_14_68; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_69; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99387; // @[Modules.scala 160:64:@47303.4]
  wire [13:0] _T_99388; // @[Modules.scala 160:64:@47304.4]
  wire [13:0] buffer_14_336; // @[Modules.scala 160:64:@47305.4]
  wire [13:0] buffer_14_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99390; // @[Modules.scala 160:64:@47307.4]
  wire [13:0] _T_99391; // @[Modules.scala 160:64:@47308.4]
  wire [13:0] buffer_14_337; // @[Modules.scala 160:64:@47309.4]
  wire [13:0] buffer_14_73; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99393; // @[Modules.scala 160:64:@47311.4]
  wire [13:0] _T_99394; // @[Modules.scala 160:64:@47312.4]
  wire [13:0] buffer_14_338; // @[Modules.scala 160:64:@47313.4]
  wire [13:0] buffer_14_75; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99396; // @[Modules.scala 160:64:@47315.4]
  wire [13:0] _T_99397; // @[Modules.scala 160:64:@47316.4]
  wire [13:0] buffer_14_339; // @[Modules.scala 160:64:@47317.4]
  wire [14:0] _T_99399; // @[Modules.scala 160:64:@47319.4]
  wire [13:0] _T_99400; // @[Modules.scala 160:64:@47320.4]
  wire [13:0] buffer_14_340; // @[Modules.scala 160:64:@47321.4]
  wire [13:0] buffer_14_78; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99402; // @[Modules.scala 160:64:@47323.4]
  wire [13:0] _T_99403; // @[Modules.scala 160:64:@47324.4]
  wire [13:0] buffer_14_341; // @[Modules.scala 160:64:@47325.4]
  wire [14:0] _T_99405; // @[Modules.scala 160:64:@47327.4]
  wire [13:0] _T_99406; // @[Modules.scala 160:64:@47328.4]
  wire [13:0] buffer_14_342; // @[Modules.scala 160:64:@47329.4]
  wire [14:0] _T_99411; // @[Modules.scala 160:64:@47335.4]
  wire [13:0] _T_99412; // @[Modules.scala 160:64:@47336.4]
  wire [13:0] buffer_14_344; // @[Modules.scala 160:64:@47337.4]
  wire [13:0] buffer_14_87; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99414; // @[Modules.scala 160:64:@47339.4]
  wire [13:0] _T_99415; // @[Modules.scala 160:64:@47340.4]
  wire [13:0] buffer_14_345; // @[Modules.scala 160:64:@47341.4]
  wire [13:0] buffer_14_88; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99417; // @[Modules.scala 160:64:@47343.4]
  wire [13:0] _T_99418; // @[Modules.scala 160:64:@47344.4]
  wire [13:0] buffer_14_346; // @[Modules.scala 160:64:@47345.4]
  wire [13:0] buffer_14_92; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99423; // @[Modules.scala 160:64:@47351.4]
  wire [13:0] _T_99424; // @[Modules.scala 160:64:@47352.4]
  wire [13:0] buffer_14_348; // @[Modules.scala 160:64:@47353.4]
  wire [14:0] _T_99426; // @[Modules.scala 160:64:@47355.4]
  wire [13:0] _T_99427; // @[Modules.scala 160:64:@47356.4]
  wire [13:0] buffer_14_349; // @[Modules.scala 160:64:@47357.4]
  wire [13:0] buffer_14_96; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99429; // @[Modules.scala 160:64:@47359.4]
  wire [13:0] _T_99430; // @[Modules.scala 160:64:@47360.4]
  wire [13:0] buffer_14_350; // @[Modules.scala 160:64:@47361.4]
  wire [13:0] buffer_14_98; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99432; // @[Modules.scala 160:64:@47363.4]
  wire [13:0] _T_99433; // @[Modules.scala 160:64:@47364.4]
  wire [13:0] buffer_14_351; // @[Modules.scala 160:64:@47365.4]
  wire [13:0] buffer_14_101; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99435; // @[Modules.scala 160:64:@47367.4]
  wire [13:0] _T_99436; // @[Modules.scala 160:64:@47368.4]
  wire [13:0] buffer_14_352; // @[Modules.scala 160:64:@47369.4]
  wire [14:0] _T_99438; // @[Modules.scala 160:64:@47371.4]
  wire [13:0] _T_99439; // @[Modules.scala 160:64:@47372.4]
  wire [13:0] buffer_14_353; // @[Modules.scala 160:64:@47373.4]
  wire [13:0] buffer_14_105; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99441; // @[Modules.scala 160:64:@47375.4]
  wire [13:0] _T_99442; // @[Modules.scala 160:64:@47376.4]
  wire [13:0] buffer_14_354; // @[Modules.scala 160:64:@47377.4]
  wire [14:0] _T_99444; // @[Modules.scala 160:64:@47379.4]
  wire [13:0] _T_99445; // @[Modules.scala 160:64:@47380.4]
  wire [13:0] buffer_14_355; // @[Modules.scala 160:64:@47381.4]
  wire [13:0] buffer_14_108; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99447; // @[Modules.scala 160:64:@47383.4]
  wire [13:0] _T_99448; // @[Modules.scala 160:64:@47384.4]
  wire [13:0] buffer_14_356; // @[Modules.scala 160:64:@47385.4]
  wire [14:0] _T_99450; // @[Modules.scala 160:64:@47387.4]
  wire [13:0] _T_99451; // @[Modules.scala 160:64:@47388.4]
  wire [13:0] buffer_14_357; // @[Modules.scala 160:64:@47389.4]
  wire [13:0] buffer_14_112; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99453; // @[Modules.scala 160:64:@47391.4]
  wire [13:0] _T_99454; // @[Modules.scala 160:64:@47392.4]
  wire [13:0] buffer_14_358; // @[Modules.scala 160:64:@47393.4]
  wire [14:0] _T_99456; // @[Modules.scala 160:64:@47395.4]
  wire [13:0] _T_99457; // @[Modules.scala 160:64:@47396.4]
  wire [13:0] buffer_14_359; // @[Modules.scala 160:64:@47397.4]
  wire [13:0] buffer_14_116; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99459; // @[Modules.scala 160:64:@47399.4]
  wire [13:0] _T_99460; // @[Modules.scala 160:64:@47400.4]
  wire [13:0] buffer_14_360; // @[Modules.scala 160:64:@47401.4]
  wire [14:0] _T_99462; // @[Modules.scala 160:64:@47403.4]
  wire [13:0] _T_99463; // @[Modules.scala 160:64:@47404.4]
  wire [13:0] buffer_14_361; // @[Modules.scala 160:64:@47405.4]
  wire [13:0] buffer_14_120; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99465; // @[Modules.scala 160:64:@47407.4]
  wire [13:0] _T_99466; // @[Modules.scala 160:64:@47408.4]
  wire [13:0] buffer_14_362; // @[Modules.scala 160:64:@47409.4]
  wire [14:0] _T_99468; // @[Modules.scala 160:64:@47411.4]
  wire [13:0] _T_99469; // @[Modules.scala 160:64:@47412.4]
  wire [13:0] buffer_14_363; // @[Modules.scala 160:64:@47413.4]
  wire [14:0] _T_99471; // @[Modules.scala 160:64:@47415.4]
  wire [13:0] _T_99472; // @[Modules.scala 160:64:@47416.4]
  wire [13:0] buffer_14_364; // @[Modules.scala 160:64:@47417.4]
  wire [13:0] buffer_14_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99474; // @[Modules.scala 160:64:@47419.4]
  wire [13:0] _T_99475; // @[Modules.scala 160:64:@47420.4]
  wire [13:0] buffer_14_365; // @[Modules.scala 160:64:@47421.4]
  wire [13:0] buffer_14_130; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_131; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99480; // @[Modules.scala 160:64:@47427.4]
  wire [13:0] _T_99481; // @[Modules.scala 160:64:@47428.4]
  wire [13:0] buffer_14_367; // @[Modules.scala 160:64:@47429.4]
  wire [13:0] buffer_14_132; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99483; // @[Modules.scala 160:64:@47431.4]
  wire [13:0] _T_99484; // @[Modules.scala 160:64:@47432.4]
  wire [13:0] buffer_14_368; // @[Modules.scala 160:64:@47433.4]
  wire [14:0] _T_99486; // @[Modules.scala 160:64:@47435.4]
  wire [13:0] _T_99487; // @[Modules.scala 160:64:@47436.4]
  wire [13:0] buffer_14_369; // @[Modules.scala 160:64:@47437.4]
  wire [13:0] buffer_14_136; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99489; // @[Modules.scala 160:64:@47439.4]
  wire [13:0] _T_99490; // @[Modules.scala 160:64:@47440.4]
  wire [13:0] buffer_14_370; // @[Modules.scala 160:64:@47441.4]
  wire [14:0] _T_99492; // @[Modules.scala 160:64:@47443.4]
  wire [13:0] _T_99493; // @[Modules.scala 160:64:@47444.4]
  wire [13:0] buffer_14_371; // @[Modules.scala 160:64:@47445.4]
  wire [13:0] buffer_14_140; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99495; // @[Modules.scala 160:64:@47447.4]
  wire [13:0] _T_99496; // @[Modules.scala 160:64:@47448.4]
  wire [13:0] buffer_14_372; // @[Modules.scala 160:64:@47449.4]
  wire [13:0] buffer_14_142; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_143; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99498; // @[Modules.scala 160:64:@47451.4]
  wire [13:0] _T_99499; // @[Modules.scala 160:64:@47452.4]
  wire [13:0] buffer_14_373; // @[Modules.scala 160:64:@47453.4]
  wire [13:0] buffer_14_144; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_145; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99501; // @[Modules.scala 160:64:@47455.4]
  wire [13:0] _T_99502; // @[Modules.scala 160:64:@47456.4]
  wire [13:0] buffer_14_374; // @[Modules.scala 160:64:@47457.4]
  wire [13:0] buffer_14_148; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99507; // @[Modules.scala 160:64:@47463.4]
  wire [13:0] _T_99508; // @[Modules.scala 160:64:@47464.4]
  wire [13:0] buffer_14_376; // @[Modules.scala 160:64:@47465.4]
  wire [14:0] _T_99510; // @[Modules.scala 160:64:@47467.4]
  wire [13:0] _T_99511; // @[Modules.scala 160:64:@47468.4]
  wire [13:0] buffer_14_377; // @[Modules.scala 160:64:@47469.4]
  wire [13:0] buffer_14_152; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99513; // @[Modules.scala 160:64:@47471.4]
  wire [13:0] _T_99514; // @[Modules.scala 160:64:@47472.4]
  wire [13:0] buffer_14_378; // @[Modules.scala 160:64:@47473.4]
  wire [13:0] buffer_14_155; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99516; // @[Modules.scala 160:64:@47475.4]
  wire [13:0] _T_99517; // @[Modules.scala 160:64:@47476.4]
  wire [13:0] buffer_14_379; // @[Modules.scala 160:64:@47477.4]
  wire [14:0] _T_99519; // @[Modules.scala 160:64:@47479.4]
  wire [13:0] _T_99520; // @[Modules.scala 160:64:@47480.4]
  wire [13:0] buffer_14_380; // @[Modules.scala 160:64:@47481.4]
  wire [13:0] buffer_14_161; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99525; // @[Modules.scala 160:64:@47487.4]
  wire [13:0] _T_99526; // @[Modules.scala 160:64:@47488.4]
  wire [13:0] buffer_14_382; // @[Modules.scala 160:64:@47489.4]
  wire [13:0] buffer_14_162; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99528; // @[Modules.scala 160:64:@47491.4]
  wire [13:0] _T_99529; // @[Modules.scala 160:64:@47492.4]
  wire [13:0] buffer_14_383; // @[Modules.scala 160:64:@47493.4]
  wire [14:0] _T_99531; // @[Modules.scala 160:64:@47495.4]
  wire [13:0] _T_99532; // @[Modules.scala 160:64:@47496.4]
  wire [13:0] buffer_14_384; // @[Modules.scala 160:64:@47497.4]
  wire [13:0] buffer_14_167; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99534; // @[Modules.scala 160:64:@47499.4]
  wire [13:0] _T_99535; // @[Modules.scala 160:64:@47500.4]
  wire [13:0] buffer_14_385; // @[Modules.scala 160:64:@47501.4]
  wire [13:0] buffer_14_169; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99537; // @[Modules.scala 160:64:@47503.4]
  wire [13:0] _T_99538; // @[Modules.scala 160:64:@47504.4]
  wire [13:0] buffer_14_386; // @[Modules.scala 160:64:@47505.4]
  wire [13:0] buffer_14_171; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99540; // @[Modules.scala 160:64:@47507.4]
  wire [13:0] _T_99541; // @[Modules.scala 160:64:@47508.4]
  wire [13:0] buffer_14_387; // @[Modules.scala 160:64:@47509.4]
  wire [14:0] _T_99543; // @[Modules.scala 160:64:@47511.4]
  wire [13:0] _T_99544; // @[Modules.scala 160:64:@47512.4]
  wire [13:0] buffer_14_388; // @[Modules.scala 160:64:@47513.4]
  wire [13:0] buffer_14_174; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99546; // @[Modules.scala 160:64:@47515.4]
  wire [13:0] _T_99547; // @[Modules.scala 160:64:@47516.4]
  wire [13:0] buffer_14_389; // @[Modules.scala 160:64:@47517.4]
  wire [13:0] buffer_14_176; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99549; // @[Modules.scala 160:64:@47519.4]
  wire [13:0] _T_99550; // @[Modules.scala 160:64:@47520.4]
  wire [13:0] buffer_14_390; // @[Modules.scala 160:64:@47521.4]
  wire [13:0] buffer_14_178; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99552; // @[Modules.scala 160:64:@47523.4]
  wire [13:0] _T_99553; // @[Modules.scala 160:64:@47524.4]
  wire [13:0] buffer_14_391; // @[Modules.scala 160:64:@47525.4]
  wire [13:0] buffer_14_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99555; // @[Modules.scala 160:64:@47527.4]
  wire [13:0] _T_99556; // @[Modules.scala 160:64:@47528.4]
  wire [13:0] buffer_14_392; // @[Modules.scala 160:64:@47529.4]
  wire [13:0] buffer_14_182; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99558; // @[Modules.scala 160:64:@47531.4]
  wire [13:0] _T_99559; // @[Modules.scala 160:64:@47532.4]
  wire [13:0] buffer_14_393; // @[Modules.scala 160:64:@47533.4]
  wire [14:0] _T_99561; // @[Modules.scala 160:64:@47535.4]
  wire [13:0] _T_99562; // @[Modules.scala 160:64:@47536.4]
  wire [13:0] buffer_14_394; // @[Modules.scala 160:64:@47537.4]
  wire [14:0] _T_99564; // @[Modules.scala 160:64:@47539.4]
  wire [13:0] _T_99565; // @[Modules.scala 160:64:@47540.4]
  wire [13:0] buffer_14_395; // @[Modules.scala 160:64:@47541.4]
  wire [13:0] buffer_14_188; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_189; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99567; // @[Modules.scala 160:64:@47543.4]
  wire [13:0] _T_99568; // @[Modules.scala 160:64:@47544.4]
  wire [13:0] buffer_14_396; // @[Modules.scala 160:64:@47545.4]
  wire [13:0] buffer_14_191; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99570; // @[Modules.scala 160:64:@47547.4]
  wire [13:0] _T_99571; // @[Modules.scala 160:64:@47548.4]
  wire [13:0] buffer_14_397; // @[Modules.scala 160:64:@47549.4]
  wire [14:0] _T_99573; // @[Modules.scala 160:64:@47551.4]
  wire [13:0] _T_99574; // @[Modules.scala 160:64:@47552.4]
  wire [13:0] buffer_14_398; // @[Modules.scala 160:64:@47553.4]
  wire [13:0] buffer_14_194; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99576; // @[Modules.scala 160:64:@47555.4]
  wire [13:0] _T_99577; // @[Modules.scala 160:64:@47556.4]
  wire [13:0] buffer_14_399; // @[Modules.scala 160:64:@47557.4]
  wire [13:0] buffer_14_196; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_197; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99579; // @[Modules.scala 160:64:@47559.4]
  wire [13:0] _T_99580; // @[Modules.scala 160:64:@47560.4]
  wire [13:0] buffer_14_400; // @[Modules.scala 160:64:@47561.4]
  wire [13:0] buffer_14_199; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99582; // @[Modules.scala 160:64:@47563.4]
  wire [13:0] _T_99583; // @[Modules.scala 160:64:@47564.4]
  wire [13:0] buffer_14_401; // @[Modules.scala 160:64:@47565.4]
  wire [14:0] _T_99585; // @[Modules.scala 160:64:@47567.4]
  wire [13:0] _T_99586; // @[Modules.scala 160:64:@47568.4]
  wire [13:0] buffer_14_402; // @[Modules.scala 160:64:@47569.4]
  wire [14:0] _T_99588; // @[Modules.scala 160:64:@47571.4]
  wire [13:0] _T_99589; // @[Modules.scala 160:64:@47572.4]
  wire [13:0] buffer_14_403; // @[Modules.scala 160:64:@47573.4]
  wire [13:0] buffer_14_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99591; // @[Modules.scala 160:64:@47575.4]
  wire [13:0] _T_99592; // @[Modules.scala 160:64:@47576.4]
  wire [13:0] buffer_14_404; // @[Modules.scala 160:64:@47577.4]
  wire [14:0] _T_99594; // @[Modules.scala 160:64:@47579.4]
  wire [13:0] _T_99595; // @[Modules.scala 160:64:@47580.4]
  wire [13:0] buffer_14_405; // @[Modules.scala 160:64:@47581.4]
  wire [14:0] _T_99597; // @[Modules.scala 160:64:@47583.4]
  wire [13:0] _T_99598; // @[Modules.scala 160:64:@47584.4]
  wire [13:0] buffer_14_406; // @[Modules.scala 160:64:@47585.4]
  wire [14:0] _T_99612; // @[Modules.scala 160:64:@47603.4]
  wire [13:0] _T_99613; // @[Modules.scala 160:64:@47604.4]
  wire [13:0] buffer_14_411; // @[Modules.scala 160:64:@47605.4]
  wire [13:0] buffer_14_222; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99618; // @[Modules.scala 160:64:@47611.4]
  wire [13:0] _T_99619; // @[Modules.scala 160:64:@47612.4]
  wire [13:0] buffer_14_413; // @[Modules.scala 160:64:@47613.4]
  wire [13:0] buffer_14_224; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_225; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99621; // @[Modules.scala 160:64:@47615.4]
  wire [13:0] _T_99622; // @[Modules.scala 160:64:@47616.4]
  wire [13:0] buffer_14_414; // @[Modules.scala 160:64:@47617.4]
  wire [13:0] buffer_14_226; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99624; // @[Modules.scala 160:64:@47619.4]
  wire [13:0] _T_99625; // @[Modules.scala 160:64:@47620.4]
  wire [13:0] buffer_14_415; // @[Modules.scala 160:64:@47621.4]
  wire [13:0] buffer_14_229; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99627; // @[Modules.scala 160:64:@47623.4]
  wire [13:0] _T_99628; // @[Modules.scala 160:64:@47624.4]
  wire [13:0] buffer_14_416; // @[Modules.scala 160:64:@47625.4]
  wire [13:0] buffer_14_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99630; // @[Modules.scala 160:64:@47627.4]
  wire [13:0] _T_99631; // @[Modules.scala 160:64:@47628.4]
  wire [13:0] buffer_14_417; // @[Modules.scala 160:64:@47629.4]
  wire [13:0] buffer_14_232; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99633; // @[Modules.scala 160:64:@47631.4]
  wire [13:0] _T_99634; // @[Modules.scala 160:64:@47632.4]
  wire [13:0] buffer_14_418; // @[Modules.scala 160:64:@47633.4]
  wire [13:0] buffer_14_234; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99636; // @[Modules.scala 160:64:@47635.4]
  wire [13:0] _T_99637; // @[Modules.scala 160:64:@47636.4]
  wire [13:0] buffer_14_419; // @[Modules.scala 160:64:@47637.4]
  wire [13:0] buffer_14_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99639; // @[Modules.scala 160:64:@47639.4]
  wire [13:0] _T_99640; // @[Modules.scala 160:64:@47640.4]
  wire [13:0] buffer_14_420; // @[Modules.scala 160:64:@47641.4]
  wire [13:0] buffer_14_239; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99642; // @[Modules.scala 160:64:@47643.4]
  wire [13:0] _T_99643; // @[Modules.scala 160:64:@47644.4]
  wire [13:0] buffer_14_421; // @[Modules.scala 160:64:@47645.4]
  wire [13:0] buffer_14_240; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99645; // @[Modules.scala 160:64:@47647.4]
  wire [13:0] _T_99646; // @[Modules.scala 160:64:@47648.4]
  wire [13:0] buffer_14_422; // @[Modules.scala 160:64:@47649.4]
  wire [13:0] buffer_14_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99648; // @[Modules.scala 160:64:@47651.4]
  wire [13:0] _T_99649; // @[Modules.scala 160:64:@47652.4]
  wire [13:0] buffer_14_423; // @[Modules.scala 160:64:@47653.4]
  wire [13:0] buffer_14_245; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99651; // @[Modules.scala 160:64:@47655.4]
  wire [13:0] _T_99652; // @[Modules.scala 160:64:@47656.4]
  wire [13:0] buffer_14_424; // @[Modules.scala 160:64:@47657.4]
  wire [14:0] _T_99657; // @[Modules.scala 160:64:@47663.4]
  wire [13:0] _T_99658; // @[Modules.scala 160:64:@47664.4]
  wire [13:0] buffer_14_426; // @[Modules.scala 160:64:@47665.4]
  wire [13:0] buffer_14_250; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99660; // @[Modules.scala 160:64:@47667.4]
  wire [13:0] _T_99661; // @[Modules.scala 160:64:@47668.4]
  wire [13:0] buffer_14_427; // @[Modules.scala 160:64:@47669.4]
  wire [13:0] buffer_14_255; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99666; // @[Modules.scala 160:64:@47675.4]
  wire [13:0] _T_99667; // @[Modules.scala 160:64:@47676.4]
  wire [13:0] buffer_14_429; // @[Modules.scala 160:64:@47677.4]
  wire [14:0] _T_99669; // @[Modules.scala 160:64:@47679.4]
  wire [13:0] _T_99670; // @[Modules.scala 160:64:@47680.4]
  wire [13:0] buffer_14_430; // @[Modules.scala 160:64:@47681.4]
  wire [13:0] buffer_14_259; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99672; // @[Modules.scala 160:64:@47683.4]
  wire [13:0] _T_99673; // @[Modules.scala 160:64:@47684.4]
  wire [13:0] buffer_14_431; // @[Modules.scala 160:64:@47685.4]
  wire [14:0] _T_99678; // @[Modules.scala 160:64:@47691.4]
  wire [13:0] _T_99679; // @[Modules.scala 160:64:@47692.4]
  wire [13:0] buffer_14_433; // @[Modules.scala 160:64:@47693.4]
  wire [13:0] buffer_14_264; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_265; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99681; // @[Modules.scala 160:64:@47695.4]
  wire [13:0] _T_99682; // @[Modules.scala 160:64:@47696.4]
  wire [13:0] buffer_14_434; // @[Modules.scala 160:64:@47697.4]
  wire [13:0] buffer_14_267; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99684; // @[Modules.scala 160:64:@47699.4]
  wire [13:0] _T_99685; // @[Modules.scala 160:64:@47700.4]
  wire [13:0] buffer_14_435; // @[Modules.scala 160:64:@47701.4]
  wire [14:0] _T_99687; // @[Modules.scala 160:64:@47703.4]
  wire [13:0] _T_99688; // @[Modules.scala 160:64:@47704.4]
  wire [13:0] buffer_14_436; // @[Modules.scala 160:64:@47705.4]
  wire [14:0] _T_99696; // @[Modules.scala 160:64:@47715.4]
  wire [13:0] _T_99697; // @[Modules.scala 160:64:@47716.4]
  wire [13:0] buffer_14_439; // @[Modules.scala 160:64:@47717.4]
  wire [13:0] buffer_14_276; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99699; // @[Modules.scala 160:64:@47719.4]
  wire [13:0] _T_99700; // @[Modules.scala 160:64:@47720.4]
  wire [13:0] buffer_14_440; // @[Modules.scala 160:64:@47721.4]
  wire [13:0] buffer_14_279; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99702; // @[Modules.scala 160:64:@47723.4]
  wire [13:0] _T_99703; // @[Modules.scala 160:64:@47724.4]
  wire [13:0] buffer_14_441; // @[Modules.scala 160:64:@47725.4]
  wire [14:0] _T_99705; // @[Modules.scala 160:64:@47727.4]
  wire [13:0] _T_99706; // @[Modules.scala 160:64:@47728.4]
  wire [13:0] buffer_14_442; // @[Modules.scala 160:64:@47729.4]
  wire [14:0] _T_99708; // @[Modules.scala 160:64:@47731.4]
  wire [13:0] _T_99709; // @[Modules.scala 160:64:@47732.4]
  wire [13:0] buffer_14_443; // @[Modules.scala 160:64:@47733.4]
  wire [14:0] _T_99717; // @[Modules.scala 160:64:@47743.4]
  wire [13:0] _T_99718; // @[Modules.scala 160:64:@47744.4]
  wire [13:0] buffer_14_446; // @[Modules.scala 160:64:@47745.4]
  wire [13:0] buffer_14_292; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99723; // @[Modules.scala 160:64:@47751.4]
  wire [13:0] _T_99724; // @[Modules.scala 160:64:@47752.4]
  wire [13:0] buffer_14_448; // @[Modules.scala 160:64:@47753.4]
  wire [13:0] buffer_14_294; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_14_295; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99726; // @[Modules.scala 160:64:@47755.4]
  wire [13:0] _T_99727; // @[Modules.scala 160:64:@47756.4]
  wire [13:0] buffer_14_449; // @[Modules.scala 160:64:@47757.4]
  wire [13:0] buffer_14_296; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99729; // @[Modules.scala 160:64:@47759.4]
  wire [13:0] _T_99730; // @[Modules.scala 160:64:@47760.4]
  wire [13:0] buffer_14_450; // @[Modules.scala 160:64:@47761.4]
  wire [13:0] buffer_14_300; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_99735; // @[Modules.scala 160:64:@47767.4]
  wire [13:0] _T_99736; // @[Modules.scala 160:64:@47768.4]
  wire [13:0] buffer_14_452; // @[Modules.scala 160:64:@47769.4]
  wire [14:0] _T_99738; // @[Modules.scala 166:64:@47771.4]
  wire [13:0] _T_99739; // @[Modules.scala 166:64:@47772.4]
  wire [13:0] buffer_14_453; // @[Modules.scala 166:64:@47773.4]
  wire [14:0] _T_99747; // @[Modules.scala 166:64:@47783.4]
  wire [13:0] _T_99748; // @[Modules.scala 166:64:@47784.4]
  wire [13:0] buffer_14_456; // @[Modules.scala 166:64:@47785.4]
  wire [14:0] _T_99750; // @[Modules.scala 166:64:@47787.4]
  wire [13:0] _T_99751; // @[Modules.scala 166:64:@47788.4]
  wire [13:0] buffer_14_457; // @[Modules.scala 166:64:@47789.4]
  wire [14:0] _T_99753; // @[Modules.scala 166:64:@47791.4]
  wire [13:0] _T_99754; // @[Modules.scala 166:64:@47792.4]
  wire [13:0] buffer_14_458; // @[Modules.scala 166:64:@47793.4]
  wire [14:0] _T_99756; // @[Modules.scala 166:64:@47795.4]
  wire [13:0] _T_99757; // @[Modules.scala 166:64:@47796.4]
  wire [13:0] buffer_14_459; // @[Modules.scala 166:64:@47797.4]
  wire [14:0] _T_99759; // @[Modules.scala 166:64:@47799.4]
  wire [13:0] _T_99760; // @[Modules.scala 166:64:@47800.4]
  wire [13:0] buffer_14_460; // @[Modules.scala 166:64:@47801.4]
  wire [14:0] _T_99762; // @[Modules.scala 166:64:@47803.4]
  wire [13:0] _T_99763; // @[Modules.scala 166:64:@47804.4]
  wire [13:0] buffer_14_461; // @[Modules.scala 166:64:@47805.4]
  wire [14:0] _T_99765; // @[Modules.scala 166:64:@47807.4]
  wire [13:0] _T_99766; // @[Modules.scala 166:64:@47808.4]
  wire [13:0] buffer_14_462; // @[Modules.scala 166:64:@47809.4]
  wire [14:0] _T_99768; // @[Modules.scala 166:64:@47811.4]
  wire [13:0] _T_99769; // @[Modules.scala 166:64:@47812.4]
  wire [13:0] buffer_14_463; // @[Modules.scala 166:64:@47813.4]
  wire [14:0] _T_99771; // @[Modules.scala 166:64:@47815.4]
  wire [13:0] _T_99772; // @[Modules.scala 166:64:@47816.4]
  wire [13:0] buffer_14_464; // @[Modules.scala 166:64:@47817.4]
  wire [14:0] _T_99774; // @[Modules.scala 166:64:@47819.4]
  wire [13:0] _T_99775; // @[Modules.scala 166:64:@47820.4]
  wire [13:0] buffer_14_465; // @[Modules.scala 166:64:@47821.4]
  wire [14:0] _T_99777; // @[Modules.scala 166:64:@47823.4]
  wire [13:0] _T_99778; // @[Modules.scala 166:64:@47824.4]
  wire [13:0] buffer_14_466; // @[Modules.scala 166:64:@47825.4]
  wire [14:0] _T_99780; // @[Modules.scala 166:64:@47827.4]
  wire [13:0] _T_99781; // @[Modules.scala 166:64:@47828.4]
  wire [13:0] buffer_14_467; // @[Modules.scala 166:64:@47829.4]
  wire [14:0] _T_99783; // @[Modules.scala 166:64:@47831.4]
  wire [13:0] _T_99784; // @[Modules.scala 166:64:@47832.4]
  wire [13:0] buffer_14_468; // @[Modules.scala 166:64:@47833.4]
  wire [14:0] _T_99786; // @[Modules.scala 166:64:@47835.4]
  wire [13:0] _T_99787; // @[Modules.scala 166:64:@47836.4]
  wire [13:0] buffer_14_469; // @[Modules.scala 166:64:@47837.4]
  wire [14:0] _T_99789; // @[Modules.scala 166:64:@47839.4]
  wire [13:0] _T_99790; // @[Modules.scala 166:64:@47840.4]
  wire [13:0] buffer_14_470; // @[Modules.scala 166:64:@47841.4]
  wire [14:0] _T_99792; // @[Modules.scala 166:64:@47843.4]
  wire [13:0] _T_99793; // @[Modules.scala 166:64:@47844.4]
  wire [13:0] buffer_14_471; // @[Modules.scala 166:64:@47845.4]
  wire [14:0] _T_99795; // @[Modules.scala 166:64:@47847.4]
  wire [13:0] _T_99796; // @[Modules.scala 166:64:@47848.4]
  wire [13:0] buffer_14_472; // @[Modules.scala 166:64:@47849.4]
  wire [14:0] _T_99798; // @[Modules.scala 166:64:@47851.4]
  wire [13:0] _T_99799; // @[Modules.scala 166:64:@47852.4]
  wire [13:0] buffer_14_473; // @[Modules.scala 166:64:@47853.4]
  wire [14:0] _T_99801; // @[Modules.scala 166:64:@47855.4]
  wire [13:0] _T_99802; // @[Modules.scala 166:64:@47856.4]
  wire [13:0] buffer_14_474; // @[Modules.scala 166:64:@47857.4]
  wire [14:0] _T_99804; // @[Modules.scala 166:64:@47859.4]
  wire [13:0] _T_99805; // @[Modules.scala 166:64:@47860.4]
  wire [13:0] buffer_14_475; // @[Modules.scala 166:64:@47861.4]
  wire [14:0] _T_99807; // @[Modules.scala 166:64:@47863.4]
  wire [13:0] _T_99808; // @[Modules.scala 166:64:@47864.4]
  wire [13:0] buffer_14_476; // @[Modules.scala 166:64:@47865.4]
  wire [14:0] _T_99810; // @[Modules.scala 166:64:@47867.4]
  wire [13:0] _T_99811; // @[Modules.scala 166:64:@47868.4]
  wire [13:0] buffer_14_477; // @[Modules.scala 166:64:@47869.4]
  wire [14:0] _T_99813; // @[Modules.scala 166:64:@47871.4]
  wire [13:0] _T_99814; // @[Modules.scala 166:64:@47872.4]
  wire [13:0] buffer_14_478; // @[Modules.scala 166:64:@47873.4]
  wire [14:0] _T_99816; // @[Modules.scala 166:64:@47875.4]
  wire [13:0] _T_99817; // @[Modules.scala 166:64:@47876.4]
  wire [13:0] buffer_14_479; // @[Modules.scala 166:64:@47877.4]
  wire [14:0] _T_99819; // @[Modules.scala 166:64:@47879.4]
  wire [13:0] _T_99820; // @[Modules.scala 166:64:@47880.4]
  wire [13:0] buffer_14_480; // @[Modules.scala 166:64:@47881.4]
  wire [14:0] _T_99822; // @[Modules.scala 166:64:@47883.4]
  wire [13:0] _T_99823; // @[Modules.scala 166:64:@47884.4]
  wire [13:0] buffer_14_481; // @[Modules.scala 166:64:@47885.4]
  wire [14:0] _T_99825; // @[Modules.scala 166:64:@47887.4]
  wire [13:0] _T_99826; // @[Modules.scala 166:64:@47888.4]
  wire [13:0] buffer_14_482; // @[Modules.scala 166:64:@47889.4]
  wire [14:0] _T_99828; // @[Modules.scala 166:64:@47891.4]
  wire [13:0] _T_99829; // @[Modules.scala 166:64:@47892.4]
  wire [13:0] buffer_14_483; // @[Modules.scala 166:64:@47893.4]
  wire [14:0] _T_99831; // @[Modules.scala 166:64:@47895.4]
  wire [13:0] _T_99832; // @[Modules.scala 166:64:@47896.4]
  wire [13:0] buffer_14_484; // @[Modules.scala 166:64:@47897.4]
  wire [14:0] _T_99834; // @[Modules.scala 166:64:@47899.4]
  wire [13:0] _T_99835; // @[Modules.scala 166:64:@47900.4]
  wire [13:0] buffer_14_485; // @[Modules.scala 166:64:@47901.4]
  wire [14:0] _T_99837; // @[Modules.scala 166:64:@47903.4]
  wire [13:0] _T_99838; // @[Modules.scala 166:64:@47904.4]
  wire [13:0] buffer_14_486; // @[Modules.scala 166:64:@47905.4]
  wire [14:0] _T_99840; // @[Modules.scala 166:64:@47907.4]
  wire [13:0] _T_99841; // @[Modules.scala 166:64:@47908.4]
  wire [13:0] buffer_14_487; // @[Modules.scala 166:64:@47909.4]
  wire [14:0] _T_99843; // @[Modules.scala 166:64:@47911.4]
  wire [13:0] _T_99844; // @[Modules.scala 166:64:@47912.4]
  wire [13:0] buffer_14_488; // @[Modules.scala 166:64:@47913.4]
  wire [14:0] _T_99846; // @[Modules.scala 166:64:@47915.4]
  wire [13:0] _T_99847; // @[Modules.scala 166:64:@47916.4]
  wire [13:0] buffer_14_489; // @[Modules.scala 166:64:@47917.4]
  wire [14:0] _T_99849; // @[Modules.scala 166:64:@47919.4]
  wire [13:0] _T_99850; // @[Modules.scala 166:64:@47920.4]
  wire [13:0] buffer_14_490; // @[Modules.scala 166:64:@47921.4]
  wire [14:0] _T_99852; // @[Modules.scala 166:64:@47923.4]
  wire [13:0] _T_99853; // @[Modules.scala 166:64:@47924.4]
  wire [13:0] buffer_14_491; // @[Modules.scala 166:64:@47925.4]
  wire [14:0] _T_99855; // @[Modules.scala 166:64:@47927.4]
  wire [13:0] _T_99856; // @[Modules.scala 166:64:@47928.4]
  wire [13:0] buffer_14_492; // @[Modules.scala 166:64:@47929.4]
  wire [14:0] _T_99858; // @[Modules.scala 166:64:@47931.4]
  wire [13:0] _T_99859; // @[Modules.scala 166:64:@47932.4]
  wire [13:0] buffer_14_493; // @[Modules.scala 166:64:@47933.4]
  wire [14:0] _T_99861; // @[Modules.scala 166:64:@47935.4]
  wire [13:0] _T_99862; // @[Modules.scala 166:64:@47936.4]
  wire [13:0] buffer_14_494; // @[Modules.scala 166:64:@47937.4]
  wire [14:0] _T_99864; // @[Modules.scala 166:64:@47939.4]
  wire [13:0] _T_99865; // @[Modules.scala 166:64:@47940.4]
  wire [13:0] buffer_14_495; // @[Modules.scala 166:64:@47941.4]
  wire [14:0] _T_99867; // @[Modules.scala 166:64:@47943.4]
  wire [13:0] _T_99868; // @[Modules.scala 166:64:@47944.4]
  wire [13:0] buffer_14_496; // @[Modules.scala 166:64:@47945.4]
  wire [14:0] _T_99870; // @[Modules.scala 166:64:@47947.4]
  wire [13:0] _T_99871; // @[Modules.scala 166:64:@47948.4]
  wire [13:0] buffer_14_497; // @[Modules.scala 166:64:@47949.4]
  wire [14:0] _T_99873; // @[Modules.scala 166:64:@47951.4]
  wire [13:0] _T_99874; // @[Modules.scala 166:64:@47952.4]
  wire [13:0] buffer_14_498; // @[Modules.scala 166:64:@47953.4]
  wire [14:0] _T_99876; // @[Modules.scala 166:64:@47955.4]
  wire [13:0] _T_99877; // @[Modules.scala 166:64:@47956.4]
  wire [13:0] buffer_14_499; // @[Modules.scala 166:64:@47957.4]
  wire [14:0] _T_99879; // @[Modules.scala 166:64:@47959.4]
  wire [13:0] _T_99880; // @[Modules.scala 166:64:@47960.4]
  wire [13:0] buffer_14_500; // @[Modules.scala 166:64:@47961.4]
  wire [14:0] _T_99882; // @[Modules.scala 166:64:@47963.4]
  wire [13:0] _T_99883; // @[Modules.scala 166:64:@47964.4]
  wire [13:0] buffer_14_501; // @[Modules.scala 166:64:@47965.4]
  wire [14:0] _T_99885; // @[Modules.scala 166:64:@47967.4]
  wire [13:0] _T_99886; // @[Modules.scala 166:64:@47968.4]
  wire [13:0] buffer_14_502; // @[Modules.scala 166:64:@47969.4]
  wire [14:0] _T_99888; // @[Modules.scala 166:64:@47971.4]
  wire [13:0] _T_99889; // @[Modules.scala 166:64:@47972.4]
  wire [13:0] buffer_14_503; // @[Modules.scala 166:64:@47973.4]
  wire [14:0] _T_99891; // @[Modules.scala 166:64:@47975.4]
  wire [13:0] _T_99892; // @[Modules.scala 166:64:@47976.4]
  wire [13:0] buffer_14_504; // @[Modules.scala 166:64:@47977.4]
  wire [14:0] _T_99894; // @[Modules.scala 166:64:@47979.4]
  wire [13:0] _T_99895; // @[Modules.scala 166:64:@47980.4]
  wire [13:0] buffer_14_505; // @[Modules.scala 166:64:@47981.4]
  wire [14:0] _T_99897; // @[Modules.scala 166:64:@47983.4]
  wire [13:0] _T_99898; // @[Modules.scala 166:64:@47984.4]
  wire [13:0] buffer_14_506; // @[Modules.scala 166:64:@47985.4]
  wire [14:0] _T_99900; // @[Modules.scala 166:64:@47987.4]
  wire [13:0] _T_99901; // @[Modules.scala 166:64:@47988.4]
  wire [13:0] buffer_14_507; // @[Modules.scala 166:64:@47989.4]
  wire [14:0] _T_99903; // @[Modules.scala 166:64:@47991.4]
  wire [13:0] _T_99904; // @[Modules.scala 166:64:@47992.4]
  wire [13:0] buffer_14_508; // @[Modules.scala 166:64:@47993.4]
  wire [14:0] _T_99906; // @[Modules.scala 166:64:@47995.4]
  wire [13:0] _T_99907; // @[Modules.scala 166:64:@47996.4]
  wire [13:0] buffer_14_509; // @[Modules.scala 166:64:@47997.4]
  wire [14:0] _T_99909; // @[Modules.scala 166:64:@47999.4]
  wire [13:0] _T_99910; // @[Modules.scala 166:64:@48000.4]
  wire [13:0] buffer_14_510; // @[Modules.scala 166:64:@48001.4]
  wire [14:0] _T_99912; // @[Modules.scala 166:64:@48003.4]
  wire [13:0] _T_99913; // @[Modules.scala 166:64:@48004.4]
  wire [13:0] buffer_14_511; // @[Modules.scala 166:64:@48005.4]
  wire [14:0] _T_99915; // @[Modules.scala 166:64:@48007.4]
  wire [13:0] _T_99916; // @[Modules.scala 166:64:@48008.4]
  wire [13:0] buffer_14_512; // @[Modules.scala 166:64:@48009.4]
  wire [14:0] _T_99918; // @[Modules.scala 166:64:@48011.4]
  wire [13:0] _T_99919; // @[Modules.scala 166:64:@48012.4]
  wire [13:0] buffer_14_513; // @[Modules.scala 166:64:@48013.4]
  wire [14:0] _T_99921; // @[Modules.scala 166:64:@48015.4]
  wire [13:0] _T_99922; // @[Modules.scala 166:64:@48016.4]
  wire [13:0] buffer_14_514; // @[Modules.scala 166:64:@48017.4]
  wire [14:0] _T_99924; // @[Modules.scala 166:64:@48019.4]
  wire [13:0] _T_99925; // @[Modules.scala 166:64:@48020.4]
  wire [13:0] buffer_14_515; // @[Modules.scala 166:64:@48021.4]
  wire [14:0] _T_99927; // @[Modules.scala 166:64:@48023.4]
  wire [13:0] _T_99928; // @[Modules.scala 166:64:@48024.4]
  wire [13:0] buffer_14_516; // @[Modules.scala 166:64:@48025.4]
  wire [14:0] _T_99930; // @[Modules.scala 166:64:@48027.4]
  wire [13:0] _T_99931; // @[Modules.scala 166:64:@48028.4]
  wire [13:0] buffer_14_517; // @[Modules.scala 166:64:@48029.4]
  wire [14:0] _T_99933; // @[Modules.scala 166:64:@48031.4]
  wire [13:0] _T_99934; // @[Modules.scala 166:64:@48032.4]
  wire [13:0] buffer_14_518; // @[Modules.scala 166:64:@48033.4]
  wire [14:0] _T_99936; // @[Modules.scala 166:64:@48035.4]
  wire [13:0] _T_99937; // @[Modules.scala 166:64:@48036.4]
  wire [13:0] buffer_14_519; // @[Modules.scala 166:64:@48037.4]
  wire [14:0] _T_99939; // @[Modules.scala 166:64:@48039.4]
  wire [13:0] _T_99940; // @[Modules.scala 166:64:@48040.4]
  wire [13:0] buffer_14_520; // @[Modules.scala 166:64:@48041.4]
  wire [14:0] _T_99942; // @[Modules.scala 166:64:@48043.4]
  wire [13:0] _T_99943; // @[Modules.scala 166:64:@48044.4]
  wire [13:0] buffer_14_521; // @[Modules.scala 166:64:@48045.4]
  wire [14:0] _T_99945; // @[Modules.scala 166:64:@48047.4]
  wire [13:0] _T_99946; // @[Modules.scala 166:64:@48048.4]
  wire [13:0] buffer_14_522; // @[Modules.scala 166:64:@48049.4]
  wire [14:0] _T_99948; // @[Modules.scala 166:64:@48051.4]
  wire [13:0] _T_99949; // @[Modules.scala 166:64:@48052.4]
  wire [13:0] buffer_14_523; // @[Modules.scala 166:64:@48053.4]
  wire [14:0] _T_99954; // @[Modules.scala 166:64:@48059.4]
  wire [13:0] _T_99955; // @[Modules.scala 166:64:@48060.4]
  wire [13:0] buffer_14_525; // @[Modules.scala 166:64:@48061.4]
  wire [14:0] _T_99957; // @[Modules.scala 166:64:@48063.4]
  wire [13:0] _T_99958; // @[Modules.scala 166:64:@48064.4]
  wire [13:0] buffer_14_526; // @[Modules.scala 166:64:@48065.4]
  wire [14:0] _T_99960; // @[Modules.scala 166:64:@48067.4]
  wire [13:0] _T_99961; // @[Modules.scala 166:64:@48068.4]
  wire [13:0] buffer_14_527; // @[Modules.scala 166:64:@48069.4]
  wire [14:0] _T_99963; // @[Modules.scala 166:64:@48071.4]
  wire [13:0] _T_99964; // @[Modules.scala 166:64:@48072.4]
  wire [13:0] buffer_14_528; // @[Modules.scala 166:64:@48073.4]
  wire [14:0] _T_99966; // @[Modules.scala 166:64:@48075.4]
  wire [13:0] _T_99967; // @[Modules.scala 166:64:@48076.4]
  wire [13:0] buffer_14_529; // @[Modules.scala 166:64:@48077.4]
  wire [14:0] _T_99969; // @[Modules.scala 166:64:@48079.4]
  wire [13:0] _T_99970; // @[Modules.scala 166:64:@48080.4]
  wire [13:0] buffer_14_530; // @[Modules.scala 166:64:@48081.4]
  wire [14:0] _T_99972; // @[Modules.scala 166:64:@48083.4]
  wire [13:0] _T_99973; // @[Modules.scala 166:64:@48084.4]
  wire [13:0] buffer_14_531; // @[Modules.scala 166:64:@48085.4]
  wire [14:0] _T_99975; // @[Modules.scala 166:64:@48087.4]
  wire [13:0] _T_99976; // @[Modules.scala 166:64:@48088.4]
  wire [13:0] buffer_14_532; // @[Modules.scala 166:64:@48089.4]
  wire [14:0] _T_99978; // @[Modules.scala 166:64:@48091.4]
  wire [13:0] _T_99979; // @[Modules.scala 166:64:@48092.4]
  wire [13:0] buffer_14_533; // @[Modules.scala 166:64:@48093.4]
  wire [14:0] _T_99981; // @[Modules.scala 166:64:@48095.4]
  wire [13:0] _T_99982; // @[Modules.scala 166:64:@48096.4]
  wire [13:0] buffer_14_534; // @[Modules.scala 166:64:@48097.4]
  wire [14:0] _T_99984; // @[Modules.scala 166:64:@48099.4]
  wire [13:0] _T_99985; // @[Modules.scala 166:64:@48100.4]
  wire [13:0] buffer_14_535; // @[Modules.scala 166:64:@48101.4]
  wire [14:0] _T_99987; // @[Modules.scala 166:64:@48103.4]
  wire [13:0] _T_99988; // @[Modules.scala 166:64:@48104.4]
  wire [13:0] buffer_14_536; // @[Modules.scala 166:64:@48105.4]
  wire [14:0] _T_99990; // @[Modules.scala 166:64:@48107.4]
  wire [13:0] _T_99991; // @[Modules.scala 166:64:@48108.4]
  wire [13:0] buffer_14_537; // @[Modules.scala 166:64:@48109.4]
  wire [14:0] _T_99993; // @[Modules.scala 166:64:@48111.4]
  wire [13:0] _T_99994; // @[Modules.scala 166:64:@48112.4]
  wire [13:0] buffer_14_538; // @[Modules.scala 166:64:@48113.4]
  wire [14:0] _T_99996; // @[Modules.scala 166:64:@48115.4]
  wire [13:0] _T_99997; // @[Modules.scala 166:64:@48116.4]
  wire [13:0] buffer_14_539; // @[Modules.scala 166:64:@48117.4]
  wire [14:0] _T_99999; // @[Modules.scala 166:64:@48119.4]
  wire [13:0] _T_100000; // @[Modules.scala 166:64:@48120.4]
  wire [13:0] buffer_14_540; // @[Modules.scala 166:64:@48121.4]
  wire [14:0] _T_100002; // @[Modules.scala 166:64:@48123.4]
  wire [13:0] _T_100003; // @[Modules.scala 166:64:@48124.4]
  wire [13:0] buffer_14_541; // @[Modules.scala 166:64:@48125.4]
  wire [14:0] _T_100005; // @[Modules.scala 166:64:@48127.4]
  wire [13:0] _T_100006; // @[Modules.scala 166:64:@48128.4]
  wire [13:0] buffer_14_542; // @[Modules.scala 166:64:@48129.4]
  wire [14:0] _T_100008; // @[Modules.scala 166:64:@48131.4]
  wire [13:0] _T_100009; // @[Modules.scala 166:64:@48132.4]
  wire [13:0] buffer_14_543; // @[Modules.scala 166:64:@48133.4]
  wire [14:0] _T_100011; // @[Modules.scala 166:64:@48135.4]
  wire [13:0] _T_100012; // @[Modules.scala 166:64:@48136.4]
  wire [13:0] buffer_14_544; // @[Modules.scala 166:64:@48137.4]
  wire [14:0] _T_100014; // @[Modules.scala 166:64:@48139.4]
  wire [13:0] _T_100015; // @[Modules.scala 166:64:@48140.4]
  wire [13:0] buffer_14_545; // @[Modules.scala 166:64:@48141.4]
  wire [14:0] _T_100017; // @[Modules.scala 166:64:@48143.4]
  wire [13:0] _T_100018; // @[Modules.scala 166:64:@48144.4]
  wire [13:0] buffer_14_546; // @[Modules.scala 166:64:@48145.4]
  wire [14:0] _T_100020; // @[Modules.scala 166:64:@48147.4]
  wire [13:0] _T_100021; // @[Modules.scala 166:64:@48148.4]
  wire [13:0] buffer_14_547; // @[Modules.scala 166:64:@48149.4]
  wire [14:0] _T_100023; // @[Modules.scala 166:64:@48151.4]
  wire [13:0] _T_100024; // @[Modules.scala 166:64:@48152.4]
  wire [13:0] buffer_14_548; // @[Modules.scala 166:64:@48153.4]
  wire [14:0] _T_100026; // @[Modules.scala 166:64:@48155.4]
  wire [13:0] _T_100027; // @[Modules.scala 166:64:@48156.4]
  wire [13:0] buffer_14_549; // @[Modules.scala 166:64:@48157.4]
  wire [14:0] _T_100029; // @[Modules.scala 166:64:@48159.4]
  wire [13:0] _T_100030; // @[Modules.scala 166:64:@48160.4]
  wire [13:0] buffer_14_550; // @[Modules.scala 166:64:@48161.4]
  wire [14:0] _T_100032; // @[Modules.scala 166:64:@48163.4]
  wire [13:0] _T_100033; // @[Modules.scala 166:64:@48164.4]
  wire [13:0] buffer_14_551; // @[Modules.scala 166:64:@48165.4]
  wire [14:0] _T_100035; // @[Modules.scala 166:64:@48167.4]
  wire [13:0] _T_100036; // @[Modules.scala 166:64:@48168.4]
  wire [13:0] buffer_14_552; // @[Modules.scala 166:64:@48169.4]
  wire [14:0] _T_100038; // @[Modules.scala 166:64:@48171.4]
  wire [13:0] _T_100039; // @[Modules.scala 166:64:@48172.4]
  wire [13:0] buffer_14_553; // @[Modules.scala 166:64:@48173.4]
  wire [14:0] _T_100041; // @[Modules.scala 166:64:@48175.4]
  wire [13:0] _T_100042; // @[Modules.scala 166:64:@48176.4]
  wire [13:0] buffer_14_554; // @[Modules.scala 166:64:@48177.4]
  wire [14:0] _T_100044; // @[Modules.scala 166:64:@48179.4]
  wire [13:0] _T_100045; // @[Modules.scala 166:64:@48180.4]
  wire [13:0] buffer_14_555; // @[Modules.scala 166:64:@48181.4]
  wire [14:0] _T_100047; // @[Modules.scala 166:64:@48183.4]
  wire [13:0] _T_100048; // @[Modules.scala 166:64:@48184.4]
  wire [13:0] buffer_14_556; // @[Modules.scala 166:64:@48185.4]
  wire [14:0] _T_100050; // @[Modules.scala 166:64:@48187.4]
  wire [13:0] _T_100051; // @[Modules.scala 166:64:@48188.4]
  wire [13:0] buffer_14_557; // @[Modules.scala 166:64:@48189.4]
  wire [14:0] _T_100053; // @[Modules.scala 166:64:@48191.4]
  wire [13:0] _T_100054; // @[Modules.scala 166:64:@48192.4]
  wire [13:0] buffer_14_558; // @[Modules.scala 166:64:@48193.4]
  wire [14:0] _T_100056; // @[Modules.scala 166:64:@48195.4]
  wire [13:0] _T_100057; // @[Modules.scala 166:64:@48196.4]
  wire [13:0] buffer_14_559; // @[Modules.scala 166:64:@48197.4]
  wire [14:0] _T_100059; // @[Modules.scala 166:64:@48199.4]
  wire [13:0] _T_100060; // @[Modules.scala 166:64:@48200.4]
  wire [13:0] buffer_14_560; // @[Modules.scala 166:64:@48201.4]
  wire [14:0] _T_100062; // @[Modules.scala 166:64:@48203.4]
  wire [13:0] _T_100063; // @[Modules.scala 166:64:@48204.4]
  wire [13:0] buffer_14_561; // @[Modules.scala 166:64:@48205.4]
  wire [14:0] _T_100065; // @[Modules.scala 166:64:@48207.4]
  wire [13:0] _T_100066; // @[Modules.scala 166:64:@48208.4]
  wire [13:0] buffer_14_562; // @[Modules.scala 166:64:@48209.4]
  wire [14:0] _T_100068; // @[Modules.scala 166:64:@48211.4]
  wire [13:0] _T_100069; // @[Modules.scala 166:64:@48212.4]
  wire [13:0] buffer_14_563; // @[Modules.scala 166:64:@48213.4]
  wire [14:0] _T_100071; // @[Modules.scala 166:64:@48215.4]
  wire [13:0] _T_100072; // @[Modules.scala 166:64:@48216.4]
  wire [13:0] buffer_14_564; // @[Modules.scala 166:64:@48217.4]
  wire [14:0] _T_100074; // @[Modules.scala 172:66:@48219.4]
  wire [13:0] _T_100075; // @[Modules.scala 172:66:@48220.4]
  wire [13:0] buffer_14_565; // @[Modules.scala 172:66:@48221.4]
  wire [14:0] _T_100077; // @[Modules.scala 160:64:@48223.4]
  wire [13:0] _T_100078; // @[Modules.scala 160:64:@48224.4]
  wire [13:0] buffer_14_566; // @[Modules.scala 160:64:@48225.4]
  wire [14:0] _T_100080; // @[Modules.scala 160:64:@48227.4]
  wire [13:0] _T_100081; // @[Modules.scala 160:64:@48228.4]
  wire [13:0] buffer_14_567; // @[Modules.scala 160:64:@48229.4]
  wire [14:0] _T_100083; // @[Modules.scala 160:64:@48231.4]
  wire [13:0] _T_100084; // @[Modules.scala 160:64:@48232.4]
  wire [13:0] buffer_14_568; // @[Modules.scala 160:64:@48233.4]
  wire [14:0] _T_100086; // @[Modules.scala 160:64:@48235.4]
  wire [13:0] _T_100087; // @[Modules.scala 160:64:@48236.4]
  wire [13:0] buffer_14_569; // @[Modules.scala 160:64:@48237.4]
  wire [14:0] _T_100089; // @[Modules.scala 160:64:@48239.4]
  wire [13:0] _T_100090; // @[Modules.scala 160:64:@48240.4]
  wire [13:0] buffer_14_570; // @[Modules.scala 160:64:@48241.4]
  wire [14:0] _T_100092; // @[Modules.scala 160:64:@48243.4]
  wire [13:0] _T_100093; // @[Modules.scala 160:64:@48244.4]
  wire [13:0] buffer_14_571; // @[Modules.scala 160:64:@48245.4]
  wire [14:0] _T_100095; // @[Modules.scala 160:64:@48247.4]
  wire [13:0] _T_100096; // @[Modules.scala 160:64:@48248.4]
  wire [13:0] buffer_14_572; // @[Modules.scala 160:64:@48249.4]
  wire [14:0] _T_100098; // @[Modules.scala 160:64:@48251.4]
  wire [13:0] _T_100099; // @[Modules.scala 160:64:@48252.4]
  wire [13:0] buffer_14_573; // @[Modules.scala 160:64:@48253.4]
  wire [14:0] _T_100101; // @[Modules.scala 160:64:@48255.4]
  wire [13:0] _T_100102; // @[Modules.scala 160:64:@48256.4]
  wire [13:0] buffer_14_574; // @[Modules.scala 160:64:@48257.4]
  wire [14:0] _T_100104; // @[Modules.scala 160:64:@48259.4]
  wire [13:0] _T_100105; // @[Modules.scala 160:64:@48260.4]
  wire [13:0] buffer_14_575; // @[Modules.scala 160:64:@48261.4]
  wire [14:0] _T_100107; // @[Modules.scala 160:64:@48263.4]
  wire [13:0] _T_100108; // @[Modules.scala 160:64:@48264.4]
  wire [13:0] buffer_14_576; // @[Modules.scala 160:64:@48265.4]
  wire [14:0] _T_100110; // @[Modules.scala 160:64:@48267.4]
  wire [13:0] _T_100111; // @[Modules.scala 160:64:@48268.4]
  wire [13:0] buffer_14_577; // @[Modules.scala 160:64:@48269.4]
  wire [14:0] _T_100113; // @[Modules.scala 160:64:@48271.4]
  wire [13:0] _T_100114; // @[Modules.scala 160:64:@48272.4]
  wire [13:0] buffer_14_578; // @[Modules.scala 160:64:@48273.4]
  wire [14:0] _T_100116; // @[Modules.scala 160:64:@48275.4]
  wire [13:0] _T_100117; // @[Modules.scala 160:64:@48276.4]
  wire [13:0] buffer_14_579; // @[Modules.scala 160:64:@48277.4]
  wire [14:0] _T_100119; // @[Modules.scala 160:64:@48279.4]
  wire [13:0] _T_100120; // @[Modules.scala 160:64:@48280.4]
  wire [13:0] buffer_14_580; // @[Modules.scala 160:64:@48281.4]
  wire [14:0] _T_100122; // @[Modules.scala 160:64:@48283.4]
  wire [13:0] _T_100123; // @[Modules.scala 160:64:@48284.4]
  wire [13:0] buffer_14_581; // @[Modules.scala 160:64:@48285.4]
  wire [14:0] _T_100125; // @[Modules.scala 160:64:@48287.4]
  wire [13:0] _T_100126; // @[Modules.scala 160:64:@48288.4]
  wire [13:0] buffer_14_582; // @[Modules.scala 160:64:@48289.4]
  wire [14:0] _T_100128; // @[Modules.scala 160:64:@48291.4]
  wire [13:0] _T_100129; // @[Modules.scala 160:64:@48292.4]
  wire [13:0] buffer_14_583; // @[Modules.scala 160:64:@48293.4]
  wire [14:0] _T_100131; // @[Modules.scala 160:64:@48295.4]
  wire [13:0] _T_100132; // @[Modules.scala 160:64:@48296.4]
  wire [13:0] buffer_14_584; // @[Modules.scala 160:64:@48297.4]
  wire [14:0] _T_100134; // @[Modules.scala 166:64:@48299.4]
  wire [13:0] _T_100135; // @[Modules.scala 166:64:@48300.4]
  wire [13:0] buffer_14_585; // @[Modules.scala 166:64:@48301.4]
  wire [14:0] _T_100137; // @[Modules.scala 166:64:@48303.4]
  wire [13:0] _T_100138; // @[Modules.scala 166:64:@48304.4]
  wire [13:0] buffer_14_586; // @[Modules.scala 166:64:@48305.4]
  wire [14:0] _T_100140; // @[Modules.scala 166:64:@48307.4]
  wire [13:0] _T_100141; // @[Modules.scala 166:64:@48308.4]
  wire [13:0] buffer_14_587; // @[Modules.scala 166:64:@48309.4]
  wire [14:0] _T_100143; // @[Modules.scala 166:64:@48311.4]
  wire [13:0] _T_100144; // @[Modules.scala 166:64:@48312.4]
  wire [13:0] buffer_14_588; // @[Modules.scala 166:64:@48313.4]
  wire [14:0] _T_100146; // @[Modules.scala 166:64:@48315.4]
  wire [13:0] _T_100147; // @[Modules.scala 166:64:@48316.4]
  wire [13:0] buffer_14_589; // @[Modules.scala 166:64:@48317.4]
  wire [14:0] _T_100149; // @[Modules.scala 166:64:@48319.4]
  wire [13:0] _T_100150; // @[Modules.scala 166:64:@48320.4]
  wire [13:0] buffer_14_590; // @[Modules.scala 166:64:@48321.4]
  wire [14:0] _T_100152; // @[Modules.scala 166:64:@48323.4]
  wire [13:0] _T_100153; // @[Modules.scala 166:64:@48324.4]
  wire [13:0] buffer_14_591; // @[Modules.scala 166:64:@48325.4]
  wire [14:0] _T_100155; // @[Modules.scala 166:64:@48327.4]
  wire [13:0] _T_100156; // @[Modules.scala 166:64:@48328.4]
  wire [13:0] buffer_14_592; // @[Modules.scala 166:64:@48329.4]
  wire [14:0] _T_100158; // @[Modules.scala 166:64:@48331.4]
  wire [13:0] _T_100159; // @[Modules.scala 166:64:@48332.4]
  wire [13:0] buffer_14_593; // @[Modules.scala 166:64:@48333.4]
  wire [14:0] _T_100161; // @[Modules.scala 166:64:@48335.4]
  wire [13:0] _T_100162; // @[Modules.scala 166:64:@48336.4]
  wire [13:0] buffer_14_594; // @[Modules.scala 166:64:@48337.4]
  wire [14:0] _T_100164; // @[Modules.scala 166:64:@48339.4]
  wire [13:0] _T_100165; // @[Modules.scala 166:64:@48340.4]
  wire [13:0] buffer_14_595; // @[Modules.scala 166:64:@48341.4]
  wire [14:0] _T_100167; // @[Modules.scala 166:64:@48343.4]
  wire [13:0] _T_100168; // @[Modules.scala 166:64:@48344.4]
  wire [13:0] buffer_14_596; // @[Modules.scala 166:64:@48345.4]
  wire [14:0] _T_100170; // @[Modules.scala 166:64:@48347.4]
  wire [13:0] _T_100171; // @[Modules.scala 166:64:@48348.4]
  wire [13:0] buffer_14_597; // @[Modules.scala 166:64:@48349.4]
  wire [14:0] _T_100173; // @[Modules.scala 172:66:@48351.4]
  wire [13:0] _T_100174; // @[Modules.scala 172:66:@48352.4]
  wire [13:0] buffer_14_598; // @[Modules.scala 172:66:@48353.4]
  wire [14:0] _T_100176; // @[Modules.scala 166:64:@48355.4]
  wire [13:0] _T_100177; // @[Modules.scala 166:64:@48356.4]
  wire [13:0] buffer_14_599; // @[Modules.scala 166:64:@48357.4]
  wire [14:0] _T_100179; // @[Modules.scala 166:64:@48359.4]
  wire [13:0] _T_100180; // @[Modules.scala 166:64:@48360.4]
  wire [13:0] buffer_14_600; // @[Modules.scala 166:64:@48361.4]
  wire [14:0] _T_100182; // @[Modules.scala 160:64:@48363.4]
  wire [13:0] _T_100183; // @[Modules.scala 160:64:@48364.4]
  wire [13:0] buffer_14_601; // @[Modules.scala 160:64:@48365.4]
  wire [14:0] _T_100185; // @[Modules.scala 172:66:@48367.4]
  wire [13:0] _T_100186; // @[Modules.scala 172:66:@48368.4]
  wire [13:0] buffer_14_602; // @[Modules.scala 172:66:@48369.4]
  wire [6:0] _T_100206; // @[Modules.scala 143:103:@48566.4]
  wire [5:0] _T_100207; // @[Modules.scala 143:103:@48567.4]
  wire [5:0] _T_100208; // @[Modules.scala 143:103:@48568.4]
  wire [5:0] _GEN_1060; // @[Modules.scala 143:103:@48632.4]
  wire [6:0] _T_100283; // @[Modules.scala 143:103:@48632.4]
  wire [5:0] _T_100284; // @[Modules.scala 143:103:@48633.4]
  wire [5:0] _T_100285; // @[Modules.scala 143:103:@48634.4]
  wire [6:0] _T_100416; // @[Modules.scala 143:103:@48746.4]
  wire [5:0] _T_100417; // @[Modules.scala 143:103:@48747.4]
  wire [5:0] _T_100418; // @[Modules.scala 143:103:@48748.4]
  wire [6:0] _T_100437; // @[Modules.scala 143:103:@48764.4]
  wire [5:0] _T_100438; // @[Modules.scala 143:103:@48765.4]
  wire [5:0] _T_100439; // @[Modules.scala 143:103:@48766.4]
  wire [5:0] _GEN_1068; // @[Modules.scala 143:103:@48830.4]
  wire [6:0] _T_100514; // @[Modules.scala 143:103:@48830.4]
  wire [5:0] _T_100515; // @[Modules.scala 143:103:@48831.4]
  wire [5:0] _T_100516; // @[Modules.scala 143:103:@48832.4]
  wire [5:0] _T_100528; // @[Modules.scala 143:103:@48842.4]
  wire [4:0] _T_100529; // @[Modules.scala 143:103:@48843.4]
  wire [4:0] _T_100530; // @[Modules.scala 143:103:@48844.4]
  wire [6:0] _T_100563; // @[Modules.scala 143:103:@48872.4]
  wire [5:0] _T_100564; // @[Modules.scala 143:103:@48873.4]
  wire [5:0] _T_100565; // @[Modules.scala 143:103:@48874.4]
  wire [5:0] _GEN_1069; // @[Modules.scala 143:103:@48878.4]
  wire [6:0] _T_100570; // @[Modules.scala 143:103:@48878.4]
  wire [5:0] _T_100571; // @[Modules.scala 143:103:@48879.4]
  wire [5:0] _T_100572; // @[Modules.scala 143:103:@48880.4]
  wire [5:0] _GEN_1073; // @[Modules.scala 143:103:@48902.4]
  wire [6:0] _T_100598; // @[Modules.scala 143:103:@48902.4]
  wire [5:0] _T_100599; // @[Modules.scala 143:103:@48903.4]
  wire [5:0] _T_100600; // @[Modules.scala 143:103:@48904.4]
  wire [6:0] _T_100605; // @[Modules.scala 143:103:@48908.4]
  wire [5:0] _T_100606; // @[Modules.scala 143:103:@48909.4]
  wire [5:0] _T_100607; // @[Modules.scala 143:103:@48910.4]
  wire [6:0] _T_100633; // @[Modules.scala 143:103:@48932.4]
  wire [5:0] _T_100634; // @[Modules.scala 143:103:@48933.4]
  wire [5:0] _T_100635; // @[Modules.scala 143:103:@48934.4]
  wire [6:0] _T_100682; // @[Modules.scala 143:103:@48974.4]
  wire [5:0] _T_100683; // @[Modules.scala 143:103:@48975.4]
  wire [5:0] _T_100684; // @[Modules.scala 143:103:@48976.4]
  wire [5:0] _T_100689; // @[Modules.scala 143:103:@48980.4]
  wire [4:0] _T_100690; // @[Modules.scala 143:103:@48981.4]
  wire [4:0] _T_100691; // @[Modules.scala 143:103:@48982.4]
  wire [6:0] _T_100696; // @[Modules.scala 143:103:@48986.4]
  wire [5:0] _T_100697; // @[Modules.scala 143:103:@48987.4]
  wire [5:0] _T_100698; // @[Modules.scala 143:103:@48988.4]
  wire [5:0] _T_100731; // @[Modules.scala 143:103:@49016.4]
  wire [4:0] _T_100732; // @[Modules.scala 143:103:@49017.4]
  wire [4:0] _T_100733; // @[Modules.scala 143:103:@49018.4]
  wire [5:0] _T_100745; // @[Modules.scala 143:103:@49028.4]
  wire [4:0] _T_100746; // @[Modules.scala 143:103:@49029.4]
  wire [4:0] _T_100747; // @[Modules.scala 143:103:@49030.4]
  wire [6:0] _T_100752; // @[Modules.scala 143:103:@49034.4]
  wire [5:0] _T_100753; // @[Modules.scala 143:103:@49035.4]
  wire [5:0] _T_100754; // @[Modules.scala 143:103:@49036.4]
  wire [6:0] _T_100759; // @[Modules.scala 143:103:@49040.4]
  wire [5:0] _T_100760; // @[Modules.scala 143:103:@49041.4]
  wire [5:0] _T_100761; // @[Modules.scala 143:103:@49042.4]
  wire [5:0] _T_100801; // @[Modules.scala 143:103:@49076.4]
  wire [4:0] _T_100802; // @[Modules.scala 143:103:@49077.4]
  wire [4:0] _T_100803; // @[Modules.scala 143:103:@49078.4]
  wire [6:0] _T_100808; // @[Modules.scala 143:103:@49082.4]
  wire [5:0] _T_100809; // @[Modules.scala 143:103:@49083.4]
  wire [5:0] _T_100810; // @[Modules.scala 143:103:@49084.4]
  wire [5:0] _T_100815; // @[Modules.scala 143:103:@49088.4]
  wire [4:0] _T_100816; // @[Modules.scala 143:103:@49089.4]
  wire [4:0] _T_100817; // @[Modules.scala 143:103:@49090.4]
  wire [6:0] _T_100829; // @[Modules.scala 143:103:@49100.4]
  wire [5:0] _T_100830; // @[Modules.scala 143:103:@49101.4]
  wire [5:0] _T_100831; // @[Modules.scala 143:103:@49102.4]
  wire [5:0] _T_100857; // @[Modules.scala 143:103:@49124.4]
  wire [4:0] _T_100858; // @[Modules.scala 143:103:@49125.4]
  wire [4:0] _T_100859; // @[Modules.scala 143:103:@49126.4]
  wire [5:0] _GEN_1083; // @[Modules.scala 143:103:@49136.4]
  wire [6:0] _T_100871; // @[Modules.scala 143:103:@49136.4]
  wire [5:0] _T_100872; // @[Modules.scala 143:103:@49137.4]
  wire [5:0] _T_100873; // @[Modules.scala 143:103:@49138.4]
  wire [5:0] _GEN_1084; // @[Modules.scala 143:103:@49148.4]
  wire [6:0] _T_100885; // @[Modules.scala 143:103:@49148.4]
  wire [5:0] _T_100886; // @[Modules.scala 143:103:@49149.4]
  wire [5:0] _T_100887; // @[Modules.scala 143:103:@49150.4]
  wire [5:0] _T_100934; // @[Modules.scala 143:103:@49190.4]
  wire [4:0] _T_100935; // @[Modules.scala 143:103:@49191.4]
  wire [4:0] _T_100936; // @[Modules.scala 143:103:@49192.4]
  wire [6:0] _T_101018; // @[Modules.scala 143:103:@49262.4]
  wire [5:0] _T_101019; // @[Modules.scala 143:103:@49263.4]
  wire [5:0] _T_101020; // @[Modules.scala 143:103:@49264.4]
  wire [6:0] _T_101046; // @[Modules.scala 143:103:@49286.4]
  wire [5:0] _T_101047; // @[Modules.scala 143:103:@49287.4]
  wire [5:0] _T_101048; // @[Modules.scala 143:103:@49288.4]
  wire [5:0] _GEN_1091; // @[Modules.scala 143:103:@49292.4]
  wire [6:0] _T_101053; // @[Modules.scala 143:103:@49292.4]
  wire [5:0] _T_101054; // @[Modules.scala 143:103:@49293.4]
  wire [5:0] _T_101055; // @[Modules.scala 143:103:@49294.4]
  wire [5:0] _T_101067; // @[Modules.scala 143:103:@49304.4]
  wire [4:0] _T_101068; // @[Modules.scala 143:103:@49305.4]
  wire [4:0] _T_101069; // @[Modules.scala 143:103:@49306.4]
  wire [5:0] _GEN_1092; // @[Modules.scala 143:103:@49310.4]
  wire [6:0] _T_101074; // @[Modules.scala 143:103:@49310.4]
  wire [5:0] _T_101075; // @[Modules.scala 143:103:@49311.4]
  wire [5:0] _T_101076; // @[Modules.scala 143:103:@49312.4]
  wire [5:0] _T_101116; // @[Modules.scala 143:103:@49346.4]
  wire [4:0] _T_101117; // @[Modules.scala 143:103:@49347.4]
  wire [4:0] _T_101118; // @[Modules.scala 143:103:@49348.4]
  wire [6:0] _T_101137; // @[Modules.scala 143:103:@49364.4]
  wire [5:0] _T_101138; // @[Modules.scala 143:103:@49365.4]
  wire [5:0] _T_101139; // @[Modules.scala 143:103:@49366.4]
  wire [6:0] _T_101158; // @[Modules.scala 143:103:@49382.4]
  wire [5:0] _T_101159; // @[Modules.scala 143:103:@49383.4]
  wire [5:0] _T_101160; // @[Modules.scala 143:103:@49384.4]
  wire [6:0] _T_101165; // @[Modules.scala 143:103:@49388.4]
  wire [5:0] _T_101166; // @[Modules.scala 143:103:@49389.4]
  wire [5:0] _T_101167; // @[Modules.scala 143:103:@49390.4]
  wire [6:0] _T_101200; // @[Modules.scala 143:103:@49418.4]
  wire [5:0] _T_101201; // @[Modules.scala 143:103:@49419.4]
  wire [5:0] _T_101202; // @[Modules.scala 143:103:@49420.4]
  wire [6:0] _T_101242; // @[Modules.scala 143:103:@49454.4]
  wire [5:0] _T_101243; // @[Modules.scala 143:103:@49455.4]
  wire [5:0] _T_101244; // @[Modules.scala 143:103:@49456.4]
  wire [6:0] _T_101368; // @[Modules.scala 143:103:@49562.4]
  wire [5:0] _T_101369; // @[Modules.scala 143:103:@49563.4]
  wire [5:0] _T_101370; // @[Modules.scala 143:103:@49564.4]
  wire [6:0] _T_101382; // @[Modules.scala 143:103:@49574.4]
  wire [5:0] _T_101383; // @[Modules.scala 143:103:@49575.4]
  wire [5:0] _T_101384; // @[Modules.scala 143:103:@49576.4]
  wire [6:0] _T_101417; // @[Modules.scala 143:103:@49604.4]
  wire [5:0] _T_101418; // @[Modules.scala 143:103:@49605.4]
  wire [5:0] _T_101419; // @[Modules.scala 143:103:@49606.4]
  wire [6:0] _T_101459; // @[Modules.scala 143:103:@49640.4]
  wire [5:0] _T_101460; // @[Modules.scala 143:103:@49641.4]
  wire [5:0] _T_101461; // @[Modules.scala 143:103:@49642.4]
  wire [5:0] _GEN_1110; // @[Modules.scala 143:103:@49646.4]
  wire [6:0] _T_101466; // @[Modules.scala 143:103:@49646.4]
  wire [5:0] _T_101467; // @[Modules.scala 143:103:@49647.4]
  wire [5:0] _T_101468; // @[Modules.scala 143:103:@49648.4]
  wire [5:0] _T_101473; // @[Modules.scala 143:103:@49652.4]
  wire [4:0] _T_101474; // @[Modules.scala 143:103:@49653.4]
  wire [4:0] _T_101475; // @[Modules.scala 143:103:@49654.4]
  wire [6:0] _T_101480; // @[Modules.scala 143:103:@49658.4]
  wire [5:0] _T_101481; // @[Modules.scala 143:103:@49659.4]
  wire [5:0] _T_101482; // @[Modules.scala 143:103:@49660.4]
  wire [6:0] _T_101536; // @[Modules.scala 143:103:@49706.4]
  wire [5:0] _T_101537; // @[Modules.scala 143:103:@49707.4]
  wire [5:0] _T_101538; // @[Modules.scala 143:103:@49708.4]
  wire [5:0] _T_101564; // @[Modules.scala 143:103:@49730.4]
  wire [4:0] _T_101565; // @[Modules.scala 143:103:@49731.4]
  wire [4:0] _T_101566; // @[Modules.scala 143:103:@49732.4]
  wire [6:0] _T_101627; // @[Modules.scala 143:103:@49784.4]
  wire [5:0] _T_101628; // @[Modules.scala 143:103:@49785.4]
  wire [5:0] _T_101629; // @[Modules.scala 143:103:@49786.4]
  wire [6:0] _T_101697; // @[Modules.scala 143:103:@49844.4]
  wire [5:0] _T_101698; // @[Modules.scala 143:103:@49845.4]
  wire [5:0] _T_101699; // @[Modules.scala 143:103:@49846.4]
  wire [5:0] _T_101704; // @[Modules.scala 143:103:@49850.4]
  wire [4:0] _T_101705; // @[Modules.scala 143:103:@49851.4]
  wire [4:0] _T_101706; // @[Modules.scala 143:103:@49852.4]
  wire [6:0] _T_101753; // @[Modules.scala 143:103:@49892.4]
  wire [5:0] _T_101754; // @[Modules.scala 143:103:@49893.4]
  wire [5:0] _T_101755; // @[Modules.scala 143:103:@49894.4]
  wire [6:0] _T_101760; // @[Modules.scala 143:103:@49898.4]
  wire [5:0] _T_101761; // @[Modules.scala 143:103:@49899.4]
  wire [5:0] _T_101762; // @[Modules.scala 143:103:@49900.4]
  wire [5:0] _GEN_1118; // @[Modules.scala 143:103:@49940.4]
  wire [6:0] _T_101809; // @[Modules.scala 143:103:@49940.4]
  wire [5:0] _T_101810; // @[Modules.scala 143:103:@49941.4]
  wire [5:0] _T_101811; // @[Modules.scala 143:103:@49942.4]
  wire [6:0] _T_101851; // @[Modules.scala 143:103:@49976.4]
  wire [5:0] _T_101852; // @[Modules.scala 143:103:@49977.4]
  wire [5:0] _T_101853; // @[Modules.scala 143:103:@49978.4]
  wire [6:0] _T_101879; // @[Modules.scala 143:103:@50000.4]
  wire [5:0] _T_101880; // @[Modules.scala 143:103:@50001.4]
  wire [5:0] _T_101881; // @[Modules.scala 143:103:@50002.4]
  wire [4:0] _T_101890; // @[Modules.scala 143:74:@50010.4]
  wire [5:0] _T_101893; // @[Modules.scala 143:103:@50012.4]
  wire [4:0] _T_101894; // @[Modules.scala 143:103:@50013.4]
  wire [4:0] _T_101895; // @[Modules.scala 143:103:@50014.4]
  wire [6:0] _T_101928; // @[Modules.scala 143:103:@50042.4]
  wire [5:0] _T_101929; // @[Modules.scala 143:103:@50043.4]
  wire [5:0] _T_101930; // @[Modules.scala 143:103:@50044.4]
  wire [6:0] _T_101935; // @[Modules.scala 143:103:@50048.4]
  wire [5:0] _T_101936; // @[Modules.scala 143:103:@50049.4]
  wire [5:0] _T_101937; // @[Modules.scala 143:103:@50050.4]
  wire [6:0] _T_101963; // @[Modules.scala 143:103:@50072.4]
  wire [5:0] _T_101964; // @[Modules.scala 143:103:@50073.4]
  wire [5:0] _T_101965; // @[Modules.scala 143:103:@50074.4]
  wire [5:0] _GEN_1125; // @[Modules.scala 143:103:@50090.4]
  wire [6:0] _T_101984; // @[Modules.scala 143:103:@50090.4]
  wire [5:0] _T_101985; // @[Modules.scala 143:103:@50091.4]
  wire [5:0] _T_101986; // @[Modules.scala 143:103:@50092.4]
  wire [6:0] _T_102012; // @[Modules.scala 143:103:@50114.4]
  wire [5:0] _T_102013; // @[Modules.scala 143:103:@50115.4]
  wire [5:0] _T_102014; // @[Modules.scala 143:103:@50116.4]
  wire [6:0] _T_102152; // @[Modules.scala 143:103:@50234.4]
  wire [5:0] _T_102153; // @[Modules.scala 143:103:@50235.4]
  wire [5:0] _T_102154; // @[Modules.scala 143:103:@50236.4]
  wire [5:0] _T_102208; // @[Modules.scala 143:103:@50282.4]
  wire [4:0] _T_102209; // @[Modules.scala 143:103:@50283.4]
  wire [4:0] _T_102210; // @[Modules.scala 143:103:@50284.4]
  wire [6:0] _T_102313; // @[Modules.scala 143:103:@50372.4]
  wire [5:0] _T_102314; // @[Modules.scala 143:103:@50373.4]
  wire [5:0] _T_102315; // @[Modules.scala 143:103:@50374.4]
  wire [6:0] _T_102341; // @[Modules.scala 143:103:@50396.4]
  wire [5:0] _T_102342; // @[Modules.scala 143:103:@50397.4]
  wire [5:0] _T_102343; // @[Modules.scala 143:103:@50398.4]
  wire [14:0] _T_102344; // @[Modules.scala 160:64:@50400.4]
  wire [13:0] _T_102345; // @[Modules.scala 160:64:@50401.4]
  wire [13:0] buffer_15_308; // @[Modules.scala 160:64:@50402.4]
  wire [13:0] buffer_15_2; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102347; // @[Modules.scala 160:64:@50404.4]
  wire [13:0] _T_102348; // @[Modules.scala 160:64:@50405.4]
  wire [13:0] buffer_15_309; // @[Modules.scala 160:64:@50406.4]
  wire [13:0] buffer_15_13; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102362; // @[Modules.scala 160:64:@50424.4]
  wire [13:0] _T_102363; // @[Modules.scala 160:64:@50425.4]
  wire [13:0] buffer_15_314; // @[Modules.scala 160:64:@50426.4]
  wire [14:0] _T_102380; // @[Modules.scala 160:64:@50448.4]
  wire [13:0] _T_102381; // @[Modules.scala 160:64:@50449.4]
  wire [13:0] buffer_15_320; // @[Modules.scala 160:64:@50450.4]
  wire [13:0] buffer_15_32; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102392; // @[Modules.scala 160:64:@50464.4]
  wire [13:0] _T_102393; // @[Modules.scala 160:64:@50465.4]
  wire [13:0] buffer_15_324; // @[Modules.scala 160:64:@50466.4]
  wire [13:0] buffer_15_35; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102395; // @[Modules.scala 160:64:@50468.4]
  wire [13:0] _T_102396; // @[Modules.scala 160:64:@50469.4]
  wire [13:0] buffer_15_325; // @[Modules.scala 160:64:@50470.4]
  wire [14:0] _T_102410; // @[Modules.scala 160:64:@50488.4]
  wire [13:0] _T_102411; // @[Modules.scala 160:64:@50489.4]
  wire [13:0] buffer_15_330; // @[Modules.scala 160:64:@50490.4]
  wire [13:0] buffer_15_46; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102413; // @[Modules.scala 160:64:@50492.4]
  wire [13:0] _T_102414; // @[Modules.scala 160:64:@50493.4]
  wire [13:0] buffer_15_331; // @[Modules.scala 160:64:@50494.4]
  wire [13:0] buffer_15_48; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102416; // @[Modules.scala 160:64:@50496.4]
  wire [13:0] _T_102417; // @[Modules.scala 160:64:@50497.4]
  wire [13:0] buffer_15_332; // @[Modules.scala 160:64:@50498.4]
  wire [13:0] buffer_15_53; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102422; // @[Modules.scala 160:64:@50504.4]
  wire [13:0] _T_102423; // @[Modules.scala 160:64:@50505.4]
  wire [13:0] buffer_15_334; // @[Modules.scala 160:64:@50506.4]
  wire [13:0] buffer_15_54; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102425; // @[Modules.scala 160:64:@50508.4]
  wire [13:0] _T_102426; // @[Modules.scala 160:64:@50509.4]
  wire [13:0] buffer_15_335; // @[Modules.scala 160:64:@50510.4]
  wire [14:0] _T_102428; // @[Modules.scala 160:64:@50512.4]
  wire [13:0] _T_102429; // @[Modules.scala 160:64:@50513.4]
  wire [13:0] buffer_15_336; // @[Modules.scala 160:64:@50514.4]
  wire [13:0] buffer_15_58; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_59; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102431; // @[Modules.scala 160:64:@50516.4]
  wire [13:0] _T_102432; // @[Modules.scala 160:64:@50517.4]
  wire [13:0] buffer_15_337; // @[Modules.scala 160:64:@50518.4]
  wire [13:0] buffer_15_63; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102437; // @[Modules.scala 160:64:@50524.4]
  wire [13:0] _T_102438; // @[Modules.scala 160:64:@50525.4]
  wire [13:0] buffer_15_339; // @[Modules.scala 160:64:@50526.4]
  wire [14:0] _T_102440; // @[Modules.scala 160:64:@50528.4]
  wire [13:0] _T_102441; // @[Modules.scala 160:64:@50529.4]
  wire [13:0] buffer_15_340; // @[Modules.scala 160:64:@50530.4]
  wire [14:0] _T_102443; // @[Modules.scala 160:64:@50532.4]
  wire [13:0] _T_102444; // @[Modules.scala 160:64:@50533.4]
  wire [13:0] buffer_15_341; // @[Modules.scala 160:64:@50534.4]
  wire [14:0] _T_102446; // @[Modules.scala 160:64:@50536.4]
  wire [13:0] _T_102447; // @[Modules.scala 160:64:@50537.4]
  wire [13:0] buffer_15_342; // @[Modules.scala 160:64:@50538.4]
  wire [13:0] buffer_15_70; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_71; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102449; // @[Modules.scala 160:64:@50540.4]
  wire [13:0] _T_102450; // @[Modules.scala 160:64:@50541.4]
  wire [13:0] buffer_15_343; // @[Modules.scala 160:64:@50542.4]
  wire [13:0] buffer_15_72; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102452; // @[Modules.scala 160:64:@50544.4]
  wire [13:0] _T_102453; // @[Modules.scala 160:64:@50545.4]
  wire [13:0] buffer_15_344; // @[Modules.scala 160:64:@50546.4]
  wire [14:0] _T_102455; // @[Modules.scala 160:64:@50548.4]
  wire [13:0] _T_102456; // @[Modules.scala 160:64:@50549.4]
  wire [13:0] buffer_15_345; // @[Modules.scala 160:64:@50550.4]
  wire [13:0] buffer_15_77; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102458; // @[Modules.scala 160:64:@50552.4]
  wire [13:0] _T_102459; // @[Modules.scala 160:64:@50553.4]
  wire [13:0] buffer_15_346; // @[Modules.scala 160:64:@50554.4]
  wire [13:0] buffer_15_79; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102461; // @[Modules.scala 160:64:@50556.4]
  wire [13:0] _T_102462; // @[Modules.scala 160:64:@50557.4]
  wire [13:0] buffer_15_347; // @[Modules.scala 160:64:@50558.4]
  wire [13:0] buffer_15_80; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_81; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102464; // @[Modules.scala 160:64:@50560.4]
  wire [13:0] _T_102465; // @[Modules.scala 160:64:@50561.4]
  wire [13:0] buffer_15_348; // @[Modules.scala 160:64:@50562.4]
  wire [14:0] _T_102470; // @[Modules.scala 160:64:@50568.4]
  wire [13:0] _T_102471; // @[Modules.scala 160:64:@50569.4]
  wire [13:0] buffer_15_350; // @[Modules.scala 160:64:@50570.4]
  wire [13:0] buffer_15_87; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102473; // @[Modules.scala 160:64:@50572.4]
  wire [13:0] _T_102474; // @[Modules.scala 160:64:@50573.4]
  wire [13:0] buffer_15_351; // @[Modules.scala 160:64:@50574.4]
  wire [13:0] buffer_15_88; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_89; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102476; // @[Modules.scala 160:64:@50576.4]
  wire [13:0] _T_102477; // @[Modules.scala 160:64:@50577.4]
  wire [13:0] buffer_15_352; // @[Modules.scala 160:64:@50578.4]
  wire [13:0] buffer_15_91; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102479; // @[Modules.scala 160:64:@50580.4]
  wire [13:0] _T_102480; // @[Modules.scala 160:64:@50581.4]
  wire [13:0] buffer_15_353; // @[Modules.scala 160:64:@50582.4]
  wire [13:0] buffer_15_95; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102485; // @[Modules.scala 160:64:@50588.4]
  wire [13:0] _T_102486; // @[Modules.scala 160:64:@50589.4]
  wire [13:0] buffer_15_355; // @[Modules.scala 160:64:@50590.4]
  wire [13:0] buffer_15_97; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102488; // @[Modules.scala 160:64:@50592.4]
  wire [13:0] _T_102489; // @[Modules.scala 160:64:@50593.4]
  wire [13:0] buffer_15_356; // @[Modules.scala 160:64:@50594.4]
  wire [13:0] buffer_15_99; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102491; // @[Modules.scala 160:64:@50596.4]
  wire [13:0] _T_102492; // @[Modules.scala 160:64:@50597.4]
  wire [13:0] buffer_15_357; // @[Modules.scala 160:64:@50598.4]
  wire [14:0] _T_102494; // @[Modules.scala 160:64:@50600.4]
  wire [13:0] _T_102495; // @[Modules.scala 160:64:@50601.4]
  wire [13:0] buffer_15_358; // @[Modules.scala 160:64:@50602.4]
  wire [14:0] _T_102497; // @[Modules.scala 160:64:@50604.4]
  wire [13:0] _T_102498; // @[Modules.scala 160:64:@50605.4]
  wire [13:0] buffer_15_359; // @[Modules.scala 160:64:@50606.4]
  wire [14:0] _T_102500; // @[Modules.scala 160:64:@50608.4]
  wire [13:0] _T_102501; // @[Modules.scala 160:64:@50609.4]
  wire [13:0] buffer_15_360; // @[Modules.scala 160:64:@50610.4]
  wire [13:0] buffer_15_106; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102503; // @[Modules.scala 160:64:@50612.4]
  wire [13:0] _T_102504; // @[Modules.scala 160:64:@50613.4]
  wire [13:0] buffer_15_361; // @[Modules.scala 160:64:@50614.4]
  wire [14:0] _T_102506; // @[Modules.scala 160:64:@50616.4]
  wire [13:0] _T_102507; // @[Modules.scala 160:64:@50617.4]
  wire [13:0] buffer_15_362; // @[Modules.scala 160:64:@50618.4]
  wire [14:0] _T_102509; // @[Modules.scala 160:64:@50620.4]
  wire [13:0] _T_102510; // @[Modules.scala 160:64:@50621.4]
  wire [13:0] buffer_15_363; // @[Modules.scala 160:64:@50622.4]
  wire [14:0] _T_102515; // @[Modules.scala 160:64:@50628.4]
  wire [13:0] _T_102516; // @[Modules.scala 160:64:@50629.4]
  wire [13:0] buffer_15_365; // @[Modules.scala 160:64:@50630.4]
  wire [14:0] _T_102518; // @[Modules.scala 160:64:@50632.4]
  wire [13:0] _T_102519; // @[Modules.scala 160:64:@50633.4]
  wire [13:0] buffer_15_366; // @[Modules.scala 160:64:@50634.4]
  wire [13:0] buffer_15_118; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102521; // @[Modules.scala 160:64:@50636.4]
  wire [13:0] _T_102522; // @[Modules.scala 160:64:@50637.4]
  wire [13:0] buffer_15_367; // @[Modules.scala 160:64:@50638.4]
  wire [14:0] _T_102524; // @[Modules.scala 160:64:@50640.4]
  wire [13:0] _T_102525; // @[Modules.scala 160:64:@50641.4]
  wire [13:0] buffer_15_368; // @[Modules.scala 160:64:@50642.4]
  wire [13:0] buffer_15_122; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_123; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102527; // @[Modules.scala 160:64:@50644.4]
  wire [13:0] _T_102528; // @[Modules.scala 160:64:@50645.4]
  wire [13:0] buffer_15_369; // @[Modules.scala 160:64:@50646.4]
  wire [13:0] buffer_15_125; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102530; // @[Modules.scala 160:64:@50648.4]
  wire [13:0] _T_102531; // @[Modules.scala 160:64:@50649.4]
  wire [13:0] buffer_15_370; // @[Modules.scala 160:64:@50650.4]
  wire [13:0] buffer_15_126; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102533; // @[Modules.scala 160:64:@50652.4]
  wire [13:0] _T_102534; // @[Modules.scala 160:64:@50653.4]
  wire [13:0] buffer_15_371; // @[Modules.scala 160:64:@50654.4]
  wire [13:0] buffer_15_132; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102542; // @[Modules.scala 160:64:@50664.4]
  wire [13:0] _T_102543; // @[Modules.scala 160:64:@50665.4]
  wire [13:0] buffer_15_374; // @[Modules.scala 160:64:@50666.4]
  wire [13:0] buffer_15_135; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102545; // @[Modules.scala 160:64:@50668.4]
  wire [13:0] _T_102546; // @[Modules.scala 160:64:@50669.4]
  wire [13:0] buffer_15_375; // @[Modules.scala 160:64:@50670.4]
  wire [14:0] _T_102548; // @[Modules.scala 160:64:@50672.4]
  wire [13:0] _T_102549; // @[Modules.scala 160:64:@50673.4]
  wire [13:0] buffer_15_376; // @[Modules.scala 160:64:@50674.4]
  wire [13:0] buffer_15_138; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_139; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102551; // @[Modules.scala 160:64:@50676.4]
  wire [13:0] _T_102552; // @[Modules.scala 160:64:@50677.4]
  wire [13:0] buffer_15_377; // @[Modules.scala 160:64:@50678.4]
  wire [14:0] _T_102554; // @[Modules.scala 160:64:@50680.4]
  wire [13:0] _T_102555; // @[Modules.scala 160:64:@50681.4]
  wire [13:0] buffer_15_378; // @[Modules.scala 160:64:@50682.4]
  wire [13:0] buffer_15_144; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102560; // @[Modules.scala 160:64:@50688.4]
  wire [13:0] _T_102561; // @[Modules.scala 160:64:@50689.4]
  wire [13:0] buffer_15_380; // @[Modules.scala 160:64:@50690.4]
  wire [14:0] _T_102563; // @[Modules.scala 160:64:@50692.4]
  wire [13:0] _T_102564; // @[Modules.scala 160:64:@50693.4]
  wire [13:0] buffer_15_381; // @[Modules.scala 160:64:@50694.4]
  wire [14:0] _T_102566; // @[Modules.scala 160:64:@50696.4]
  wire [13:0] _T_102567; // @[Modules.scala 160:64:@50697.4]
  wire [13:0] buffer_15_382; // @[Modules.scala 160:64:@50698.4]
  wire [13:0] buffer_15_150; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102569; // @[Modules.scala 160:64:@50700.4]
  wire [13:0] _T_102570; // @[Modules.scala 160:64:@50701.4]
  wire [13:0] buffer_15_383; // @[Modules.scala 160:64:@50702.4]
  wire [14:0] _T_102572; // @[Modules.scala 160:64:@50704.4]
  wire [13:0] _T_102573; // @[Modules.scala 160:64:@50705.4]
  wire [13:0] buffer_15_384; // @[Modules.scala 160:64:@50706.4]
  wire [14:0] _T_102578; // @[Modules.scala 160:64:@50712.4]
  wire [13:0] _T_102579; // @[Modules.scala 160:64:@50713.4]
  wire [13:0] buffer_15_386; // @[Modules.scala 160:64:@50714.4]
  wire [14:0] _T_102587; // @[Modules.scala 160:64:@50724.4]
  wire [13:0] _T_102588; // @[Modules.scala 160:64:@50725.4]
  wire [13:0] buffer_15_389; // @[Modules.scala 160:64:@50726.4]
  wire [14:0] _T_102590; // @[Modules.scala 160:64:@50728.4]
  wire [13:0] _T_102591; // @[Modules.scala 160:64:@50729.4]
  wire [13:0] buffer_15_390; // @[Modules.scala 160:64:@50730.4]
  wire [14:0] _T_102593; // @[Modules.scala 160:64:@50732.4]
  wire [13:0] _T_102594; // @[Modules.scala 160:64:@50733.4]
  wire [13:0] buffer_15_391; // @[Modules.scala 160:64:@50734.4]
  wire [13:0] buffer_15_168; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102596; // @[Modules.scala 160:64:@50736.4]
  wire [13:0] _T_102597; // @[Modules.scala 160:64:@50737.4]
  wire [13:0] buffer_15_392; // @[Modules.scala 160:64:@50738.4]
  wire [13:0] buffer_15_170; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102599; // @[Modules.scala 160:64:@50740.4]
  wire [13:0] _T_102600; // @[Modules.scala 160:64:@50741.4]
  wire [13:0] buffer_15_393; // @[Modules.scala 160:64:@50742.4]
  wire [14:0] _T_102602; // @[Modules.scala 160:64:@50744.4]
  wire [13:0] _T_102603; // @[Modules.scala 160:64:@50745.4]
  wire [13:0] buffer_15_394; // @[Modules.scala 160:64:@50746.4]
  wire [13:0] buffer_15_175; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102605; // @[Modules.scala 160:64:@50748.4]
  wire [13:0] _T_102606; // @[Modules.scala 160:64:@50749.4]
  wire [13:0] buffer_15_395; // @[Modules.scala 160:64:@50750.4]
  wire [14:0] _T_102611; // @[Modules.scala 160:64:@50756.4]
  wire [13:0] _T_102612; // @[Modules.scala 160:64:@50757.4]
  wire [13:0] buffer_15_397; // @[Modules.scala 160:64:@50758.4]
  wire [13:0] buffer_15_181; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102614; // @[Modules.scala 160:64:@50760.4]
  wire [13:0] _T_102615; // @[Modules.scala 160:64:@50761.4]
  wire [13:0] buffer_15_398; // @[Modules.scala 160:64:@50762.4]
  wire [13:0] buffer_15_182; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_183; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102617; // @[Modules.scala 160:64:@50764.4]
  wire [13:0] _T_102618; // @[Modules.scala 160:64:@50765.4]
  wire [13:0] buffer_15_399; // @[Modules.scala 160:64:@50766.4]
  wire [13:0] buffer_15_184; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102620; // @[Modules.scala 160:64:@50768.4]
  wire [13:0] _T_102621; // @[Modules.scala 160:64:@50769.4]
  wire [13:0] buffer_15_400; // @[Modules.scala 160:64:@50770.4]
  wire [14:0] _T_102626; // @[Modules.scala 160:64:@50776.4]
  wire [13:0] _T_102627; // @[Modules.scala 160:64:@50777.4]
  wire [13:0] buffer_15_402; // @[Modules.scala 160:64:@50778.4]
  wire [14:0] _T_102629; // @[Modules.scala 160:64:@50780.4]
  wire [13:0] _T_102630; // @[Modules.scala 160:64:@50781.4]
  wire [13:0] buffer_15_403; // @[Modules.scala 160:64:@50782.4]
  wire [13:0] buffer_15_192; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102632; // @[Modules.scala 160:64:@50784.4]
  wire [13:0] _T_102633; // @[Modules.scala 160:64:@50785.4]
  wire [13:0] buffer_15_404; // @[Modules.scala 160:64:@50786.4]
  wire [13:0] buffer_15_196; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102638; // @[Modules.scala 160:64:@50792.4]
  wire [13:0] _T_102639; // @[Modules.scala 160:64:@50793.4]
  wire [13:0] buffer_15_406; // @[Modules.scala 160:64:@50794.4]
  wire [13:0] buffer_15_205; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102650; // @[Modules.scala 160:64:@50808.4]
  wire [13:0] _T_102651; // @[Modules.scala 160:64:@50809.4]
  wire [13:0] buffer_15_410; // @[Modules.scala 160:64:@50810.4]
  wire [14:0] _T_102659; // @[Modules.scala 160:64:@50820.4]
  wire [13:0] _T_102660; // @[Modules.scala 160:64:@50821.4]
  wire [13:0] buffer_15_413; // @[Modules.scala 160:64:@50822.4]
  wire [14:0] _T_102662; // @[Modules.scala 160:64:@50824.4]
  wire [13:0] _T_102663; // @[Modules.scala 160:64:@50825.4]
  wire [13:0] buffer_15_414; // @[Modules.scala 160:64:@50826.4]
  wire [13:0] buffer_15_215; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102665; // @[Modules.scala 160:64:@50828.4]
  wire [13:0] _T_102666; // @[Modules.scala 160:64:@50829.4]
  wire [13:0] buffer_15_415; // @[Modules.scala 160:64:@50830.4]
  wire [13:0] buffer_15_216; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102668; // @[Modules.scala 160:64:@50832.4]
  wire [13:0] _T_102669; // @[Modules.scala 160:64:@50833.4]
  wire [13:0] buffer_15_416; // @[Modules.scala 160:64:@50834.4]
  wire [14:0] _T_102671; // @[Modules.scala 160:64:@50836.4]
  wire [13:0] _T_102672; // @[Modules.scala 160:64:@50837.4]
  wire [13:0] buffer_15_417; // @[Modules.scala 160:64:@50838.4]
  wire [14:0] _T_102674; // @[Modules.scala 160:64:@50840.4]
  wire [13:0] _T_102675; // @[Modules.scala 160:64:@50841.4]
  wire [13:0] buffer_15_418; // @[Modules.scala 160:64:@50842.4]
  wire [13:0] buffer_15_223; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102677; // @[Modules.scala 160:64:@50844.4]
  wire [13:0] _T_102678; // @[Modules.scala 160:64:@50845.4]
  wire [13:0] buffer_15_419; // @[Modules.scala 160:64:@50846.4]
  wire [13:0] buffer_15_224; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102680; // @[Modules.scala 160:64:@50848.4]
  wire [13:0] _T_102681; // @[Modules.scala 160:64:@50849.4]
  wire [13:0] buffer_15_420; // @[Modules.scala 160:64:@50850.4]
  wire [14:0] _T_102683; // @[Modules.scala 160:64:@50852.4]
  wire [13:0] _T_102684; // @[Modules.scala 160:64:@50853.4]
  wire [13:0] buffer_15_421; // @[Modules.scala 160:64:@50854.4]
  wire [14:0] _T_102686; // @[Modules.scala 160:64:@50856.4]
  wire [13:0] _T_102687; // @[Modules.scala 160:64:@50857.4]
  wire [13:0] buffer_15_422; // @[Modules.scala 160:64:@50858.4]
  wire [13:0] buffer_15_231; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102689; // @[Modules.scala 160:64:@50860.4]
  wire [13:0] _T_102690; // @[Modules.scala 160:64:@50861.4]
  wire [13:0] buffer_15_423; // @[Modules.scala 160:64:@50862.4]
  wire [13:0] buffer_15_237; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102698; // @[Modules.scala 160:64:@50872.4]
  wire [13:0] _T_102699; // @[Modules.scala 160:64:@50873.4]
  wire [13:0] buffer_15_426; // @[Modules.scala 160:64:@50874.4]
  wire [14:0] _T_102701; // @[Modules.scala 160:64:@50876.4]
  wire [13:0] _T_102702; // @[Modules.scala 160:64:@50877.4]
  wire [13:0] buffer_15_427; // @[Modules.scala 160:64:@50878.4]
  wire [13:0] buffer_15_241; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102704; // @[Modules.scala 160:64:@50880.4]
  wire [13:0] _T_102705; // @[Modules.scala 160:64:@50881.4]
  wire [13:0] buffer_15_428; // @[Modules.scala 160:64:@50882.4]
  wire [13:0] buffer_15_243; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102707; // @[Modules.scala 160:64:@50884.4]
  wire [13:0] _T_102708; // @[Modules.scala 160:64:@50885.4]
  wire [13:0] buffer_15_429; // @[Modules.scala 160:64:@50886.4]
  wire [13:0] buffer_15_248; // @[Modules.scala 112:22:@8.4]
  wire [13:0] buffer_15_249; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102716; // @[Modules.scala 160:64:@50896.4]
  wire [13:0] _T_102717; // @[Modules.scala 160:64:@50897.4]
  wire [13:0] buffer_15_432; // @[Modules.scala 160:64:@50898.4]
  wire [14:0] _T_102719; // @[Modules.scala 160:64:@50900.4]
  wire [13:0] _T_102720; // @[Modules.scala 160:64:@50901.4]
  wire [13:0] buffer_15_433; // @[Modules.scala 160:64:@50902.4]
  wire [13:0] buffer_15_253; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102722; // @[Modules.scala 160:64:@50904.4]
  wire [13:0] _T_102723; // @[Modules.scala 160:64:@50905.4]
  wire [13:0] buffer_15_434; // @[Modules.scala 160:64:@50906.4]
  wire [13:0] buffer_15_256; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102728; // @[Modules.scala 160:64:@50912.4]
  wire [13:0] _T_102729; // @[Modules.scala 160:64:@50913.4]
  wire [13:0] buffer_15_436; // @[Modules.scala 160:64:@50914.4]
  wire [14:0] _T_102731; // @[Modules.scala 160:64:@50916.4]
  wire [13:0] _T_102732; // @[Modules.scala 160:64:@50917.4]
  wire [13:0] buffer_15_437; // @[Modules.scala 160:64:@50918.4]
  wire [13:0] buffer_15_260; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102734; // @[Modules.scala 160:64:@50920.4]
  wire [13:0] _T_102735; // @[Modules.scala 160:64:@50921.4]
  wire [13:0] buffer_15_438; // @[Modules.scala 160:64:@50922.4]
  wire [14:0] _T_102737; // @[Modules.scala 160:64:@50924.4]
  wire [13:0] _T_102738; // @[Modules.scala 160:64:@50925.4]
  wire [13:0] buffer_15_439; // @[Modules.scala 160:64:@50926.4]
  wire [14:0] _T_102743; // @[Modules.scala 160:64:@50932.4]
  wire [13:0] _T_102744; // @[Modules.scala 160:64:@50933.4]
  wire [13:0] buffer_15_441; // @[Modules.scala 160:64:@50934.4]
  wire [14:0] _T_102752; // @[Modules.scala 160:64:@50944.4]
  wire [13:0] _T_102753; // @[Modules.scala 160:64:@50945.4]
  wire [13:0] buffer_15_444; // @[Modules.scala 160:64:@50946.4]
  wire [14:0] _T_102755; // @[Modules.scala 160:64:@50948.4]
  wire [13:0] _T_102756; // @[Modules.scala 160:64:@50949.4]
  wire [13:0] buffer_15_445; // @[Modules.scala 160:64:@50950.4]
  wire [14:0] _T_102758; // @[Modules.scala 160:64:@50952.4]
  wire [13:0] _T_102759; // @[Modules.scala 160:64:@50953.4]
  wire [13:0] buffer_15_446; // @[Modules.scala 160:64:@50954.4]
  wire [13:0] buffer_15_280; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102764; // @[Modules.scala 160:64:@50960.4]
  wire [13:0] _T_102765; // @[Modules.scala 160:64:@50961.4]
  wire [13:0] buffer_15_448; // @[Modules.scala 160:64:@50962.4]
  wire [13:0] buffer_15_288; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102776; // @[Modules.scala 160:64:@50976.4]
  wire [13:0] _T_102777; // @[Modules.scala 160:64:@50977.4]
  wire [13:0] buffer_15_452; // @[Modules.scala 160:64:@50978.4]
  wire [13:0] buffer_15_303; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102797; // @[Modules.scala 160:64:@51004.4]
  wire [13:0] _T_102798; // @[Modules.scala 160:64:@51005.4]
  wire [13:0] buffer_15_459; // @[Modules.scala 160:64:@51006.4]
  wire [13:0] buffer_15_307; // @[Modules.scala 112:22:@8.4]
  wire [14:0] _T_102803; // @[Modules.scala 160:64:@51012.4]
  wire [13:0] _T_102804; // @[Modules.scala 160:64:@51013.4]
  wire [13:0] buffer_15_461; // @[Modules.scala 160:64:@51014.4]
  wire [14:0] _T_102806; // @[Modules.scala 160:64:@51016.4]
  wire [13:0] _T_102807; // @[Modules.scala 160:64:@51017.4]
  wire [13:0] buffer_15_462; // @[Modules.scala 160:64:@51018.4]
  wire [14:0] _T_102815; // @[Modules.scala 160:64:@51028.4]
  wire [13:0] _T_102816; // @[Modules.scala 160:64:@51029.4]
  wire [13:0] buffer_15_465; // @[Modules.scala 160:64:@51030.4]
  wire [14:0] _T_102824; // @[Modules.scala 160:64:@51040.4]
  wire [13:0] _T_102825; // @[Modules.scala 160:64:@51041.4]
  wire [13:0] buffer_15_468; // @[Modules.scala 160:64:@51042.4]
  wire [14:0] _T_102830; // @[Modules.scala 160:64:@51048.4]
  wire [13:0] _T_102831; // @[Modules.scala 160:64:@51049.4]
  wire [13:0] buffer_15_470; // @[Modules.scala 160:64:@51050.4]
  wire [14:0] _T_102836; // @[Modules.scala 160:64:@51056.4]
  wire [13:0] _T_102837; // @[Modules.scala 160:64:@51057.4]
  wire [13:0] buffer_15_472; // @[Modules.scala 160:64:@51058.4]
  wire [14:0] _T_102839; // @[Modules.scala 160:64:@51060.4]
  wire [13:0] _T_102840; // @[Modules.scala 160:64:@51061.4]
  wire [13:0] buffer_15_473; // @[Modules.scala 160:64:@51062.4]
  wire [14:0] _T_102842; // @[Modules.scala 160:64:@51064.4]
  wire [13:0] _T_102843; // @[Modules.scala 160:64:@51065.4]
  wire [13:0] buffer_15_474; // @[Modules.scala 160:64:@51066.4]
  wire [14:0] _T_102845; // @[Modules.scala 160:64:@51068.4]
  wire [13:0] _T_102846; // @[Modules.scala 160:64:@51069.4]
  wire [13:0] buffer_15_475; // @[Modules.scala 160:64:@51070.4]
  wire [14:0] _T_102848; // @[Modules.scala 160:64:@51072.4]
  wire [13:0] _T_102849; // @[Modules.scala 160:64:@51073.4]
  wire [13:0] buffer_15_476; // @[Modules.scala 160:64:@51074.4]
  wire [14:0] _T_102851; // @[Modules.scala 160:64:@51076.4]
  wire [13:0] _T_102852; // @[Modules.scala 160:64:@51077.4]
  wire [13:0] buffer_15_477; // @[Modules.scala 160:64:@51078.4]
  wire [14:0] _T_102854; // @[Modules.scala 160:64:@51080.4]
  wire [13:0] _T_102855; // @[Modules.scala 160:64:@51081.4]
  wire [13:0] buffer_15_478; // @[Modules.scala 160:64:@51082.4]
  wire [14:0] _T_102857; // @[Modules.scala 160:64:@51084.4]
  wire [13:0] _T_102858; // @[Modules.scala 160:64:@51085.4]
  wire [13:0] buffer_15_479; // @[Modules.scala 160:64:@51086.4]
  wire [14:0] _T_102860; // @[Modules.scala 160:64:@51088.4]
  wire [13:0] _T_102861; // @[Modules.scala 160:64:@51089.4]
  wire [13:0] buffer_15_480; // @[Modules.scala 160:64:@51090.4]
  wire [14:0] _T_102863; // @[Modules.scala 160:64:@51092.4]
  wire [13:0] _T_102864; // @[Modules.scala 160:64:@51093.4]
  wire [13:0] buffer_15_481; // @[Modules.scala 160:64:@51094.4]
  wire [14:0] _T_102866; // @[Modules.scala 160:64:@51096.4]
  wire [13:0] _T_102867; // @[Modules.scala 160:64:@51097.4]
  wire [13:0] buffer_15_482; // @[Modules.scala 160:64:@51098.4]
  wire [14:0] _T_102869; // @[Modules.scala 160:64:@51100.4]
  wire [13:0] _T_102870; // @[Modules.scala 160:64:@51101.4]
  wire [13:0] buffer_15_483; // @[Modules.scala 160:64:@51102.4]
  wire [14:0] _T_102872; // @[Modules.scala 160:64:@51104.4]
  wire [13:0] _T_102873; // @[Modules.scala 160:64:@51105.4]
  wire [13:0] buffer_15_484; // @[Modules.scala 160:64:@51106.4]
  wire [14:0] _T_102875; // @[Modules.scala 160:64:@51108.4]
  wire [13:0] _T_102876; // @[Modules.scala 160:64:@51109.4]
  wire [13:0] buffer_15_485; // @[Modules.scala 160:64:@51110.4]
  wire [14:0] _T_102878; // @[Modules.scala 160:64:@51112.4]
  wire [13:0] _T_102879; // @[Modules.scala 160:64:@51113.4]
  wire [13:0] buffer_15_486; // @[Modules.scala 160:64:@51114.4]
  wire [14:0] _T_102881; // @[Modules.scala 160:64:@51116.4]
  wire [13:0] _T_102882; // @[Modules.scala 160:64:@51117.4]
  wire [13:0] buffer_15_487; // @[Modules.scala 160:64:@51118.4]
  wire [14:0] _T_102884; // @[Modules.scala 160:64:@51120.4]
  wire [13:0] _T_102885; // @[Modules.scala 160:64:@51121.4]
  wire [13:0] buffer_15_488; // @[Modules.scala 160:64:@51122.4]
  wire [14:0] _T_102887; // @[Modules.scala 160:64:@51124.4]
  wire [13:0] _T_102888; // @[Modules.scala 160:64:@51125.4]
  wire [13:0] buffer_15_489; // @[Modules.scala 160:64:@51126.4]
  wire [14:0] _T_102890; // @[Modules.scala 160:64:@51128.4]
  wire [13:0] _T_102891; // @[Modules.scala 160:64:@51129.4]
  wire [13:0] buffer_15_490; // @[Modules.scala 160:64:@51130.4]
  wire [14:0] _T_102893; // @[Modules.scala 160:64:@51132.4]
  wire [13:0] _T_102894; // @[Modules.scala 160:64:@51133.4]
  wire [13:0] buffer_15_491; // @[Modules.scala 160:64:@51134.4]
  wire [14:0] _T_102896; // @[Modules.scala 160:64:@51136.4]
  wire [13:0] _T_102897; // @[Modules.scala 160:64:@51137.4]
  wire [13:0] buffer_15_492; // @[Modules.scala 160:64:@51138.4]
  wire [14:0] _T_102899; // @[Modules.scala 160:64:@51140.4]
  wire [13:0] _T_102900; // @[Modules.scala 160:64:@51141.4]
  wire [13:0] buffer_15_493; // @[Modules.scala 160:64:@51142.4]
  wire [14:0] _T_102902; // @[Modules.scala 160:64:@51144.4]
  wire [13:0] _T_102903; // @[Modules.scala 160:64:@51145.4]
  wire [13:0] buffer_15_494; // @[Modules.scala 160:64:@51146.4]
  wire [14:0] _T_102905; // @[Modules.scala 160:64:@51148.4]
  wire [13:0] _T_102906; // @[Modules.scala 160:64:@51149.4]
  wire [13:0] buffer_15_495; // @[Modules.scala 160:64:@51150.4]
  wire [14:0] _T_102908; // @[Modules.scala 160:64:@51152.4]
  wire [13:0] _T_102909; // @[Modules.scala 160:64:@51153.4]
  wire [13:0] buffer_15_496; // @[Modules.scala 160:64:@51154.4]
  wire [14:0] _T_102911; // @[Modules.scala 160:64:@51156.4]
  wire [13:0] _T_102912; // @[Modules.scala 160:64:@51157.4]
  wire [13:0] buffer_15_497; // @[Modules.scala 160:64:@51158.4]
  wire [14:0] _T_102914; // @[Modules.scala 160:64:@51160.4]
  wire [13:0] _T_102915; // @[Modules.scala 160:64:@51161.4]
  wire [13:0] buffer_15_498; // @[Modules.scala 160:64:@51162.4]
  wire [14:0] _T_102917; // @[Modules.scala 160:64:@51164.4]
  wire [13:0] _T_102918; // @[Modules.scala 160:64:@51165.4]
  wire [13:0] buffer_15_499; // @[Modules.scala 160:64:@51166.4]
  wire [14:0] _T_102920; // @[Modules.scala 160:64:@51168.4]
  wire [13:0] _T_102921; // @[Modules.scala 160:64:@51169.4]
  wire [13:0] buffer_15_500; // @[Modules.scala 160:64:@51170.4]
  wire [14:0] _T_102923; // @[Modules.scala 160:64:@51172.4]
  wire [13:0] _T_102924; // @[Modules.scala 160:64:@51173.4]
  wire [13:0] buffer_15_501; // @[Modules.scala 160:64:@51174.4]
  wire [14:0] _T_102926; // @[Modules.scala 160:64:@51176.4]
  wire [13:0] _T_102927; // @[Modules.scala 160:64:@51177.4]
  wire [13:0] buffer_15_502; // @[Modules.scala 160:64:@51178.4]
  wire [14:0] _T_102929; // @[Modules.scala 160:64:@51180.4]
  wire [13:0] _T_102930; // @[Modules.scala 160:64:@51181.4]
  wire [13:0] buffer_15_503; // @[Modules.scala 160:64:@51182.4]
  wire [14:0] _T_102932; // @[Modules.scala 160:64:@51184.4]
  wire [13:0] _T_102933; // @[Modules.scala 160:64:@51185.4]
  wire [13:0] buffer_15_504; // @[Modules.scala 160:64:@51186.4]
  wire [14:0] _T_102935; // @[Modules.scala 160:64:@51188.4]
  wire [13:0] _T_102936; // @[Modules.scala 160:64:@51189.4]
  wire [13:0] buffer_15_505; // @[Modules.scala 160:64:@51190.4]
  wire [14:0] _T_102938; // @[Modules.scala 160:64:@51192.4]
  wire [13:0] _T_102939; // @[Modules.scala 160:64:@51193.4]
  wire [13:0] buffer_15_506; // @[Modules.scala 160:64:@51194.4]
  wire [14:0] _T_102941; // @[Modules.scala 160:64:@51196.4]
  wire [13:0] _T_102942; // @[Modules.scala 160:64:@51197.4]
  wire [13:0] buffer_15_507; // @[Modules.scala 160:64:@51198.4]
  wire [14:0] _T_102944; // @[Modules.scala 160:64:@51200.4]
  wire [13:0] _T_102945; // @[Modules.scala 160:64:@51201.4]
  wire [13:0] buffer_15_508; // @[Modules.scala 160:64:@51202.4]
  wire [14:0] _T_102947; // @[Modules.scala 160:64:@51204.4]
  wire [13:0] _T_102948; // @[Modules.scala 160:64:@51205.4]
  wire [13:0] buffer_15_509; // @[Modules.scala 160:64:@51206.4]
  wire [14:0] _T_102950; // @[Modules.scala 160:64:@51208.4]
  wire [13:0] _T_102951; // @[Modules.scala 160:64:@51209.4]
  wire [13:0] buffer_15_510; // @[Modules.scala 160:64:@51210.4]
  wire [14:0] _T_102953; // @[Modules.scala 160:64:@51212.4]
  wire [13:0] _T_102954; // @[Modules.scala 160:64:@51213.4]
  wire [13:0] buffer_15_511; // @[Modules.scala 160:64:@51214.4]
  wire [14:0] _T_102956; // @[Modules.scala 160:64:@51216.4]
  wire [13:0] _T_102957; // @[Modules.scala 160:64:@51217.4]
  wire [13:0] buffer_15_512; // @[Modules.scala 160:64:@51218.4]
  wire [14:0] _T_102959; // @[Modules.scala 160:64:@51220.4]
  wire [13:0] _T_102960; // @[Modules.scala 160:64:@51221.4]
  wire [13:0] buffer_15_513; // @[Modules.scala 160:64:@51222.4]
  wire [14:0] _T_102962; // @[Modules.scala 160:64:@51224.4]
  wire [13:0] _T_102963; // @[Modules.scala 160:64:@51225.4]
  wire [13:0] buffer_15_514; // @[Modules.scala 160:64:@51226.4]
  wire [14:0] _T_102965; // @[Modules.scala 160:64:@51228.4]
  wire [13:0] _T_102966; // @[Modules.scala 160:64:@51229.4]
  wire [13:0] buffer_15_515; // @[Modules.scala 160:64:@51230.4]
  wire [14:0] _T_102968; // @[Modules.scala 160:64:@51232.4]
  wire [13:0] _T_102969; // @[Modules.scala 160:64:@51233.4]
  wire [13:0] buffer_15_516; // @[Modules.scala 160:64:@51234.4]
  wire [14:0] _T_102971; // @[Modules.scala 160:64:@51236.4]
  wire [13:0] _T_102972; // @[Modules.scala 160:64:@51237.4]
  wire [13:0] buffer_15_517; // @[Modules.scala 160:64:@51238.4]
  wire [14:0] _T_102974; // @[Modules.scala 160:64:@51240.4]
  wire [13:0] _T_102975; // @[Modules.scala 160:64:@51241.4]
  wire [13:0] buffer_15_518; // @[Modules.scala 160:64:@51242.4]
  wire [14:0] _T_102977; // @[Modules.scala 160:64:@51244.4]
  wire [13:0] _T_102978; // @[Modules.scala 160:64:@51245.4]
  wire [13:0] buffer_15_519; // @[Modules.scala 160:64:@51246.4]
  wire [14:0] _T_102980; // @[Modules.scala 160:64:@51248.4]
  wire [13:0] _T_102981; // @[Modules.scala 160:64:@51249.4]
  wire [13:0] buffer_15_520; // @[Modules.scala 160:64:@51250.4]
  wire [14:0] _T_102983; // @[Modules.scala 160:64:@51252.4]
  wire [13:0] _T_102984; // @[Modules.scala 160:64:@51253.4]
  wire [13:0] buffer_15_521; // @[Modules.scala 160:64:@51254.4]
  wire [14:0] _T_102986; // @[Modules.scala 160:64:@51256.4]
  wire [13:0] _T_102987; // @[Modules.scala 160:64:@51257.4]
  wire [13:0] buffer_15_522; // @[Modules.scala 160:64:@51258.4]
  wire [14:0] _T_102989; // @[Modules.scala 160:64:@51260.4]
  wire [13:0] _T_102990; // @[Modules.scala 160:64:@51261.4]
  wire [13:0] buffer_15_523; // @[Modules.scala 160:64:@51262.4]
  wire [14:0] _T_102992; // @[Modules.scala 160:64:@51264.4]
  wire [13:0] _T_102993; // @[Modules.scala 160:64:@51265.4]
  wire [13:0] buffer_15_524; // @[Modules.scala 160:64:@51266.4]
  wire [14:0] _T_102995; // @[Modules.scala 160:64:@51268.4]
  wire [13:0] _T_102996; // @[Modules.scala 160:64:@51269.4]
  wire [13:0] buffer_15_525; // @[Modules.scala 160:64:@51270.4]
  wire [14:0] _T_102998; // @[Modules.scala 160:64:@51272.4]
  wire [13:0] _T_102999; // @[Modules.scala 160:64:@51273.4]
  wire [13:0] buffer_15_526; // @[Modules.scala 160:64:@51274.4]
  wire [14:0] _T_103001; // @[Modules.scala 160:64:@51276.4]
  wire [13:0] _T_103002; // @[Modules.scala 160:64:@51277.4]
  wire [13:0] buffer_15_527; // @[Modules.scala 160:64:@51278.4]
  wire [14:0] _T_103004; // @[Modules.scala 160:64:@51280.4]
  wire [13:0] _T_103005; // @[Modules.scala 160:64:@51281.4]
  wire [13:0] buffer_15_528; // @[Modules.scala 160:64:@51282.4]
  wire [14:0] _T_103007; // @[Modules.scala 160:64:@51284.4]
  wire [13:0] _T_103008; // @[Modules.scala 160:64:@51285.4]
  wire [13:0] buffer_15_529; // @[Modules.scala 160:64:@51286.4]
  wire [14:0] _T_103010; // @[Modules.scala 160:64:@51288.4]
  wire [13:0] _T_103011; // @[Modules.scala 160:64:@51289.4]
  wire [13:0] buffer_15_530; // @[Modules.scala 160:64:@51290.4]
  wire [14:0] _T_103013; // @[Modules.scala 160:64:@51292.4]
  wire [13:0] _T_103014; // @[Modules.scala 160:64:@51293.4]
  wire [13:0] buffer_15_531; // @[Modules.scala 160:64:@51294.4]
  wire [14:0] _T_103016; // @[Modules.scala 160:64:@51296.4]
  wire [13:0] _T_103017; // @[Modules.scala 160:64:@51297.4]
  wire [13:0] buffer_15_532; // @[Modules.scala 160:64:@51298.4]
  wire [14:0] _T_103022; // @[Modules.scala 160:64:@51304.4]
  wire [13:0] _T_103023; // @[Modules.scala 160:64:@51305.4]
  wire [13:0] buffer_15_534; // @[Modules.scala 160:64:@51306.4]
  wire [14:0] _T_103025; // @[Modules.scala 160:64:@51308.4]
  wire [13:0] _T_103026; // @[Modules.scala 160:64:@51309.4]
  wire [13:0] buffer_15_535; // @[Modules.scala 160:64:@51310.4]
  wire [14:0] _T_103031; // @[Modules.scala 160:64:@51316.4]
  wire [13:0] _T_103032; // @[Modules.scala 160:64:@51317.4]
  wire [13:0] buffer_15_537; // @[Modules.scala 160:64:@51318.4]
  wire [14:0] _T_103034; // @[Modules.scala 160:64:@51320.4]
  wire [13:0] _T_103035; // @[Modules.scala 160:64:@51321.4]
  wire [13:0] buffer_15_538; // @[Modules.scala 160:64:@51322.4]
  wire [14:0] _T_103037; // @[Modules.scala 166:64:@51324.4]
  wire [13:0] _T_103038; // @[Modules.scala 166:64:@51325.4]
  wire [13:0] buffer_15_539; // @[Modules.scala 166:64:@51326.4]
  wire [14:0] _T_103040; // @[Modules.scala 166:64:@51328.4]
  wire [13:0] _T_103041; // @[Modules.scala 166:64:@51329.4]
  wire [13:0] buffer_15_540; // @[Modules.scala 166:64:@51330.4]
  wire [14:0] _T_103046; // @[Modules.scala 166:64:@51336.4]
  wire [13:0] _T_103047; // @[Modules.scala 166:64:@51337.4]
  wire [13:0] buffer_15_542; // @[Modules.scala 166:64:@51338.4]
  wire [14:0] _T_103049; // @[Modules.scala 166:64:@51340.4]
  wire [13:0] _T_103050; // @[Modules.scala 166:64:@51341.4]
  wire [13:0] buffer_15_543; // @[Modules.scala 166:64:@51342.4]
  wire [14:0] _T_103052; // @[Modules.scala 166:64:@51344.4]
  wire [13:0] _T_103053; // @[Modules.scala 166:64:@51345.4]
  wire [13:0] buffer_15_544; // @[Modules.scala 166:64:@51346.4]
  wire [14:0] _T_103055; // @[Modules.scala 166:64:@51348.4]
  wire [13:0] _T_103056; // @[Modules.scala 166:64:@51349.4]
  wire [13:0] buffer_15_545; // @[Modules.scala 166:64:@51350.4]
  wire [14:0] _T_103058; // @[Modules.scala 166:64:@51352.4]
  wire [13:0] _T_103059; // @[Modules.scala 166:64:@51353.4]
  wire [13:0] buffer_15_546; // @[Modules.scala 166:64:@51354.4]
  wire [14:0] _T_103061; // @[Modules.scala 166:64:@51356.4]
  wire [13:0] _T_103062; // @[Modules.scala 166:64:@51357.4]
  wire [13:0] buffer_15_547; // @[Modules.scala 166:64:@51358.4]
  wire [14:0] _T_103064; // @[Modules.scala 166:64:@51360.4]
  wire [13:0] _T_103065; // @[Modules.scala 166:64:@51361.4]
  wire [13:0] buffer_15_548; // @[Modules.scala 166:64:@51362.4]
  wire [14:0] _T_103067; // @[Modules.scala 166:64:@51364.4]
  wire [13:0] _T_103068; // @[Modules.scala 166:64:@51365.4]
  wire [13:0] buffer_15_549; // @[Modules.scala 166:64:@51366.4]
  wire [14:0] _T_103070; // @[Modules.scala 166:64:@51368.4]
  wire [13:0] _T_103071; // @[Modules.scala 166:64:@51369.4]
  wire [13:0] buffer_15_550; // @[Modules.scala 166:64:@51370.4]
  wire [14:0] _T_103073; // @[Modules.scala 166:64:@51372.4]
  wire [13:0] _T_103074; // @[Modules.scala 166:64:@51373.4]
  wire [13:0] buffer_15_551; // @[Modules.scala 166:64:@51374.4]
  wire [14:0] _T_103076; // @[Modules.scala 166:64:@51376.4]
  wire [13:0] _T_103077; // @[Modules.scala 166:64:@51377.4]
  wire [13:0] buffer_15_552; // @[Modules.scala 166:64:@51378.4]
  wire [14:0] _T_103079; // @[Modules.scala 166:64:@51380.4]
  wire [13:0] _T_103080; // @[Modules.scala 166:64:@51381.4]
  wire [13:0] buffer_15_553; // @[Modules.scala 166:64:@51382.4]
  wire [14:0] _T_103082; // @[Modules.scala 166:64:@51384.4]
  wire [13:0] _T_103083; // @[Modules.scala 166:64:@51385.4]
  wire [13:0] buffer_15_554; // @[Modules.scala 166:64:@51386.4]
  wire [14:0] _T_103085; // @[Modules.scala 166:64:@51388.4]
  wire [13:0] _T_103086; // @[Modules.scala 166:64:@51389.4]
  wire [13:0] buffer_15_555; // @[Modules.scala 166:64:@51390.4]
  wire [14:0] _T_103088; // @[Modules.scala 166:64:@51392.4]
  wire [13:0] _T_103089; // @[Modules.scala 166:64:@51393.4]
  wire [13:0] buffer_15_556; // @[Modules.scala 166:64:@51394.4]
  wire [14:0] _T_103091; // @[Modules.scala 166:64:@51396.4]
  wire [13:0] _T_103092; // @[Modules.scala 166:64:@51397.4]
  wire [13:0] buffer_15_557; // @[Modules.scala 166:64:@51398.4]
  wire [14:0] _T_103094; // @[Modules.scala 166:64:@51400.4]
  wire [13:0] _T_103095; // @[Modules.scala 166:64:@51401.4]
  wire [13:0] buffer_15_558; // @[Modules.scala 166:64:@51402.4]
  wire [14:0] _T_103097; // @[Modules.scala 166:64:@51404.4]
  wire [13:0] _T_103098; // @[Modules.scala 166:64:@51405.4]
  wire [13:0] buffer_15_559; // @[Modules.scala 166:64:@51406.4]
  wire [14:0] _T_103100; // @[Modules.scala 166:64:@51408.4]
  wire [13:0] _T_103101; // @[Modules.scala 166:64:@51409.4]
  wire [13:0] buffer_15_560; // @[Modules.scala 166:64:@51410.4]
  wire [14:0] _T_103103; // @[Modules.scala 166:64:@51412.4]
  wire [13:0] _T_103104; // @[Modules.scala 166:64:@51413.4]
  wire [13:0] buffer_15_561; // @[Modules.scala 166:64:@51414.4]
  wire [14:0] _T_103106; // @[Modules.scala 166:64:@51416.4]
  wire [13:0] _T_103107; // @[Modules.scala 166:64:@51417.4]
  wire [13:0] buffer_15_562; // @[Modules.scala 166:64:@51418.4]
  wire [14:0] _T_103109; // @[Modules.scala 166:64:@51420.4]
  wire [13:0] _T_103110; // @[Modules.scala 166:64:@51421.4]
  wire [13:0] buffer_15_563; // @[Modules.scala 166:64:@51422.4]
  wire [14:0] _T_103112; // @[Modules.scala 166:64:@51424.4]
  wire [13:0] _T_103113; // @[Modules.scala 166:64:@51425.4]
  wire [13:0] buffer_15_564; // @[Modules.scala 166:64:@51426.4]
  wire [14:0] _T_103115; // @[Modules.scala 166:64:@51428.4]
  wire [13:0] _T_103116; // @[Modules.scala 166:64:@51429.4]
  wire [13:0] buffer_15_565; // @[Modules.scala 166:64:@51430.4]
  wire [14:0] _T_103118; // @[Modules.scala 166:64:@51432.4]
  wire [13:0] _T_103119; // @[Modules.scala 166:64:@51433.4]
  wire [13:0] buffer_15_566; // @[Modules.scala 166:64:@51434.4]
  wire [14:0] _T_103121; // @[Modules.scala 166:64:@51436.4]
  wire [13:0] _T_103122; // @[Modules.scala 166:64:@51437.4]
  wire [13:0] buffer_15_567; // @[Modules.scala 166:64:@51438.4]
  wire [14:0] _T_103124; // @[Modules.scala 166:64:@51440.4]
  wire [13:0] _T_103125; // @[Modules.scala 166:64:@51441.4]
  wire [13:0] buffer_15_568; // @[Modules.scala 166:64:@51442.4]
  wire [14:0] _T_103127; // @[Modules.scala 166:64:@51444.4]
  wire [13:0] _T_103128; // @[Modules.scala 166:64:@51445.4]
  wire [13:0] buffer_15_569; // @[Modules.scala 166:64:@51446.4]
  wire [14:0] _T_103130; // @[Modules.scala 166:64:@51448.4]
  wire [13:0] _T_103131; // @[Modules.scala 166:64:@51449.4]
  wire [13:0] buffer_15_570; // @[Modules.scala 166:64:@51450.4]
  wire [14:0] _T_103133; // @[Modules.scala 166:64:@51452.4]
  wire [13:0] _T_103134; // @[Modules.scala 166:64:@51453.4]
  wire [13:0] buffer_15_571; // @[Modules.scala 166:64:@51454.4]
  wire [14:0] _T_103136; // @[Modules.scala 166:64:@51456.4]
  wire [13:0] _T_103137; // @[Modules.scala 166:64:@51457.4]
  wire [13:0] buffer_15_572; // @[Modules.scala 166:64:@51458.4]
  wire [14:0] _T_103139; // @[Modules.scala 166:64:@51460.4]
  wire [13:0] _T_103140; // @[Modules.scala 166:64:@51461.4]
  wire [13:0] buffer_15_573; // @[Modules.scala 166:64:@51462.4]
  wire [14:0] _T_103142; // @[Modules.scala 166:64:@51464.4]
  wire [13:0] _T_103143; // @[Modules.scala 166:64:@51465.4]
  wire [13:0] buffer_15_574; // @[Modules.scala 166:64:@51466.4]
  wire [14:0] _T_103145; // @[Modules.scala 166:64:@51468.4]
  wire [13:0] _T_103146; // @[Modules.scala 166:64:@51469.4]
  wire [13:0] buffer_15_575; // @[Modules.scala 166:64:@51470.4]
  wire [14:0] _T_103148; // @[Modules.scala 166:64:@51472.4]
  wire [13:0] _T_103149; // @[Modules.scala 166:64:@51473.4]
  wire [13:0] buffer_15_576; // @[Modules.scala 166:64:@51474.4]
  wire [14:0] _T_103151; // @[Modules.scala 160:64:@51476.4]
  wire [13:0] _T_103152; // @[Modules.scala 160:64:@51477.4]
  wire [13:0] buffer_15_577; // @[Modules.scala 160:64:@51478.4]
  wire [14:0] _T_103154; // @[Modules.scala 160:64:@51480.4]
  wire [13:0] _T_103155; // @[Modules.scala 160:64:@51481.4]
  wire [13:0] buffer_15_578; // @[Modules.scala 160:64:@51482.4]
  wire [14:0] _T_103157; // @[Modules.scala 160:64:@51484.4]
  wire [13:0] _T_103158; // @[Modules.scala 160:64:@51485.4]
  wire [13:0] buffer_15_579; // @[Modules.scala 160:64:@51486.4]
  wire [14:0] _T_103160; // @[Modules.scala 160:64:@51488.4]
  wire [13:0] _T_103161; // @[Modules.scala 160:64:@51489.4]
  wire [13:0] buffer_15_580; // @[Modules.scala 160:64:@51490.4]
  wire [14:0] _T_103163; // @[Modules.scala 160:64:@51492.4]
  wire [13:0] _T_103164; // @[Modules.scala 160:64:@51493.4]
  wire [13:0] buffer_15_581; // @[Modules.scala 160:64:@51494.4]
  wire [14:0] _T_103166; // @[Modules.scala 160:64:@51496.4]
  wire [13:0] _T_103167; // @[Modules.scala 160:64:@51497.4]
  wire [13:0] buffer_15_582; // @[Modules.scala 160:64:@51498.4]
  wire [14:0] _T_103169; // @[Modules.scala 160:64:@51500.4]
  wire [13:0] _T_103170; // @[Modules.scala 160:64:@51501.4]
  wire [13:0] buffer_15_583; // @[Modules.scala 160:64:@51502.4]
  wire [14:0] _T_103172; // @[Modules.scala 160:64:@51504.4]
  wire [13:0] _T_103173; // @[Modules.scala 160:64:@51505.4]
  wire [13:0] buffer_15_584; // @[Modules.scala 160:64:@51506.4]
  wire [14:0] _T_103175; // @[Modules.scala 160:64:@51508.4]
  wire [13:0] _T_103176; // @[Modules.scala 160:64:@51509.4]
  wire [13:0] buffer_15_585; // @[Modules.scala 160:64:@51510.4]
  wire [14:0] _T_103178; // @[Modules.scala 160:64:@51512.4]
  wire [13:0] _T_103179; // @[Modules.scala 160:64:@51513.4]
  wire [13:0] buffer_15_586; // @[Modules.scala 160:64:@51514.4]
  wire [14:0] _T_103181; // @[Modules.scala 160:64:@51516.4]
  wire [13:0] _T_103182; // @[Modules.scala 160:64:@51517.4]
  wire [13:0] buffer_15_587; // @[Modules.scala 160:64:@51518.4]
  wire [14:0] _T_103184; // @[Modules.scala 160:64:@51520.4]
  wire [13:0] _T_103185; // @[Modules.scala 160:64:@51521.4]
  wire [13:0] buffer_15_588; // @[Modules.scala 160:64:@51522.4]
  wire [14:0] _T_103187; // @[Modules.scala 160:64:@51524.4]
  wire [13:0] _T_103188; // @[Modules.scala 160:64:@51525.4]
  wire [13:0] buffer_15_589; // @[Modules.scala 160:64:@51526.4]
  wire [14:0] _T_103190; // @[Modules.scala 160:64:@51528.4]
  wire [13:0] _T_103191; // @[Modules.scala 160:64:@51529.4]
  wire [13:0] buffer_15_590; // @[Modules.scala 160:64:@51530.4]
  wire [14:0] _T_103193; // @[Modules.scala 160:64:@51532.4]
  wire [13:0] _T_103194; // @[Modules.scala 160:64:@51533.4]
  wire [13:0] buffer_15_591; // @[Modules.scala 160:64:@51534.4]
  wire [14:0] _T_103196; // @[Modules.scala 160:64:@51536.4]
  wire [13:0] _T_103197; // @[Modules.scala 160:64:@51537.4]
  wire [13:0] buffer_15_592; // @[Modules.scala 160:64:@51538.4]
  wire [14:0] _T_103199; // @[Modules.scala 160:64:@51540.4]
  wire [13:0] _T_103200; // @[Modules.scala 160:64:@51541.4]
  wire [13:0] buffer_15_593; // @[Modules.scala 160:64:@51542.4]
  wire [14:0] _T_103202; // @[Modules.scala 160:64:@51544.4]
  wire [13:0] _T_103203; // @[Modules.scala 160:64:@51545.4]
  wire [13:0] buffer_15_594; // @[Modules.scala 160:64:@51546.4]
  wire [14:0] _T_103205; // @[Modules.scala 160:64:@51548.4]
  wire [13:0] _T_103206; // @[Modules.scala 160:64:@51549.4]
  wire [13:0] buffer_15_595; // @[Modules.scala 160:64:@51550.4]
  wire [14:0] _T_103208; // @[Modules.scala 166:64:@51552.4]
  wire [13:0] _T_103209; // @[Modules.scala 166:64:@51553.4]
  wire [13:0] buffer_15_596; // @[Modules.scala 166:64:@51554.4]
  wire [14:0] _T_103211; // @[Modules.scala 166:64:@51556.4]
  wire [13:0] _T_103212; // @[Modules.scala 166:64:@51557.4]
  wire [13:0] buffer_15_597; // @[Modules.scala 166:64:@51558.4]
  wire [14:0] _T_103214; // @[Modules.scala 166:64:@51560.4]
  wire [13:0] _T_103215; // @[Modules.scala 166:64:@51561.4]
  wire [13:0] buffer_15_598; // @[Modules.scala 166:64:@51562.4]
  wire [14:0] _T_103217; // @[Modules.scala 166:64:@51564.4]
  wire [13:0] _T_103218; // @[Modules.scala 166:64:@51565.4]
  wire [13:0] buffer_15_599; // @[Modules.scala 166:64:@51566.4]
  wire [14:0] _T_103220; // @[Modules.scala 166:64:@51568.4]
  wire [13:0] _T_103221; // @[Modules.scala 166:64:@51569.4]
  wire [13:0] buffer_15_600; // @[Modules.scala 166:64:@51570.4]
  wire [14:0] _T_103223; // @[Modules.scala 166:64:@51572.4]
  wire [13:0] _T_103224; // @[Modules.scala 166:64:@51573.4]
  wire [13:0] buffer_15_601; // @[Modules.scala 166:64:@51574.4]
  wire [14:0] _T_103226; // @[Modules.scala 166:64:@51576.4]
  wire [13:0] _T_103227; // @[Modules.scala 166:64:@51577.4]
  wire [13:0] buffer_15_602; // @[Modules.scala 166:64:@51578.4]
  wire [14:0] _T_103229; // @[Modules.scala 166:64:@51580.4]
  wire [13:0] _T_103230; // @[Modules.scala 166:64:@51581.4]
  wire [13:0] buffer_15_603; // @[Modules.scala 166:64:@51582.4]
  wire [14:0] _T_103232; // @[Modules.scala 166:64:@51584.4]
  wire [13:0] _T_103233; // @[Modules.scala 166:64:@51585.4]
  wire [13:0] buffer_15_604; // @[Modules.scala 166:64:@51586.4]
  wire [14:0] _T_103235; // @[Modules.scala 172:66:@51588.4]
  wire [13:0] _T_103236; // @[Modules.scala 172:66:@51589.4]
  wire [13:0] buffer_15_605; // @[Modules.scala 172:66:@51590.4]
  wire [14:0] _T_103238; // @[Modules.scala 160:64:@51592.4]
  wire [13:0] _T_103239; // @[Modules.scala 160:64:@51593.4]
  wire [13:0] buffer_15_606; // @[Modules.scala 160:64:@51594.4]
  wire [14:0] _T_103241; // @[Modules.scala 160:64:@51596.4]
  wire [13:0] _T_103242; // @[Modules.scala 160:64:@51597.4]
  wire [13:0] buffer_15_607; // @[Modules.scala 160:64:@51598.4]
  wire [14:0] _T_103244; // @[Modules.scala 160:64:@51600.4]
  wire [13:0] _T_103245; // @[Modules.scala 160:64:@51601.4]
  wire [13:0] buffer_15_608; // @[Modules.scala 160:64:@51602.4]
  wire [14:0] _T_103247; // @[Modules.scala 160:64:@51604.4]
  wire [13:0] _T_103248; // @[Modules.scala 160:64:@51605.4]
  wire [13:0] buffer_15_609; // @[Modules.scala 160:64:@51606.4]
  wire [14:0] _T_103250; // @[Modules.scala 160:64:@51608.4]
  wire [13:0] _T_103251; // @[Modules.scala 160:64:@51609.4]
  wire [13:0] buffer_15_610; // @[Modules.scala 160:64:@51610.4]
  wire [14:0] _T_103253; // @[Modules.scala 166:64:@51612.4]
  wire [13:0] _T_103254; // @[Modules.scala 166:64:@51613.4]
  wire [13:0] buffer_15_611; // @[Modules.scala 166:64:@51614.4]
  wire [14:0] _T_103256; // @[Modules.scala 166:64:@51616.4]
  wire [13:0] _T_103257; // @[Modules.scala 166:64:@51617.4]
  wire [13:0] buffer_15_612; // @[Modules.scala 166:64:@51618.4]
  wire [14:0] _T_103259; // @[Modules.scala 160:64:@51620.4]
  wire [13:0] _T_103260; // @[Modules.scala 160:64:@51621.4]
  wire [13:0] buffer_15_613; // @[Modules.scala 160:64:@51622.4]
  wire [14:0] _T_103262; // @[Modules.scala 172:66:@51624.4]
  wire [13:0] _T_103263; // @[Modules.scala 172:66:@51625.4]
  wire [13:0] buffer_15_614; // @[Modules.scala 172:66:@51626.4]
  assign _T_54199 = $signed(4'sh1) * $signed(io_in_12); // @[Modules.scala 150:74:@9.4]
  assign _T_54201 = $signed(4'sh1) * $signed(io_in_13); // @[Modules.scala 151:80:@10.4]
  assign _T_54202 = $signed(_T_54199) + $signed(_T_54201); // @[Modules.scala 150:103:@11.4]
  assign _T_54203 = _T_54202[5:0]; // @[Modules.scala 150:103:@12.4]
  assign _T_54204 = $signed(_T_54203); // @[Modules.scala 150:103:@13.4]
  assign _T_54206 = $signed(4'sh1) * $signed(io_in_14); // @[Modules.scala 150:74:@15.4]
  assign _T_54208 = $signed(4'sh1) * $signed(io_in_15); // @[Modules.scala 151:80:@16.4]
  assign _T_54209 = $signed(_T_54206) + $signed(_T_54208); // @[Modules.scala 150:103:@17.4]
  assign _T_54210 = _T_54209[5:0]; // @[Modules.scala 150:103:@18.4]
  assign _T_54211 = $signed(_T_54210); // @[Modules.scala 150:103:@19.4]
  assign _T_54213 = $signed(-4'sh1) * $signed(io_in_28); // @[Modules.scala 150:74:@21.4]
  assign _T_54215 = $signed(4'sh1) * $signed(io_in_32); // @[Modules.scala 151:80:@22.4]
  assign _GEN_0 = {{1{_T_54213[4]}},_T_54213}; // @[Modules.scala 150:103:@23.4]
  assign _T_54216 = $signed(_GEN_0) + $signed(_T_54215); // @[Modules.scala 150:103:@23.4]
  assign _T_54217 = _T_54216[5:0]; // @[Modules.scala 150:103:@24.4]
  assign _T_54218 = $signed(_T_54217); // @[Modules.scala 150:103:@25.4]
  assign _T_54220 = $signed(4'sh1) * $signed(io_in_33); // @[Modules.scala 150:74:@27.4]
  assign _T_54222 = $signed(4'sh1) * $signed(io_in_36); // @[Modules.scala 151:80:@28.4]
  assign _T_54223 = $signed(_T_54220) + $signed(_T_54222); // @[Modules.scala 150:103:@29.4]
  assign _T_54224 = _T_54223[5:0]; // @[Modules.scala 150:103:@30.4]
  assign _T_54225 = $signed(_T_54224); // @[Modules.scala 150:103:@31.4]
  assign _T_54227 = $signed(4'sh1) * $signed(io_in_37); // @[Modules.scala 150:74:@33.4]
  assign _T_54229 = $signed(4'sh1) * $signed(io_in_38); // @[Modules.scala 151:80:@34.4]
  assign _T_54230 = $signed(_T_54227) + $signed(_T_54229); // @[Modules.scala 150:103:@35.4]
  assign _T_54231 = _T_54230[5:0]; // @[Modules.scala 150:103:@36.4]
  assign _T_54232 = $signed(_T_54231); // @[Modules.scala 150:103:@37.4]
  assign _T_54234 = $signed(4'sh1) * $signed(io_in_39); // @[Modules.scala 150:74:@39.4]
  assign _T_54236 = $signed(4'sh1) * $signed(io_in_40); // @[Modules.scala 151:80:@40.4]
  assign _T_54237 = $signed(_T_54234) + $signed(_T_54236); // @[Modules.scala 150:103:@41.4]
  assign _T_54238 = _T_54237[5:0]; // @[Modules.scala 150:103:@42.4]
  assign _T_54239 = $signed(_T_54238); // @[Modules.scala 150:103:@43.4]
  assign _T_54241 = $signed(4'sh1) * $signed(io_in_41); // @[Modules.scala 150:74:@45.4]
  assign _T_54243 = $signed(4'sh1) * $signed(io_in_42); // @[Modules.scala 151:80:@46.4]
  assign _T_54244 = $signed(_T_54241) + $signed(_T_54243); // @[Modules.scala 150:103:@47.4]
  assign _T_54245 = _T_54244[5:0]; // @[Modules.scala 150:103:@48.4]
  assign _T_54246 = $signed(_T_54245); // @[Modules.scala 150:103:@49.4]
  assign _T_54248 = $signed(4'sh1) * $signed(io_in_43); // @[Modules.scala 150:74:@51.4]
  assign _T_54250 = $signed(4'sh1) * $signed(io_in_44); // @[Modules.scala 151:80:@52.4]
  assign _T_54251 = $signed(_T_54248) + $signed(_T_54250); // @[Modules.scala 150:103:@53.4]
  assign _T_54252 = _T_54251[5:0]; // @[Modules.scala 150:103:@54.4]
  assign _T_54253 = $signed(_T_54252); // @[Modules.scala 150:103:@55.4]
  assign _T_54255 = $signed(4'sh1) * $signed(io_in_45); // @[Modules.scala 150:74:@57.4]
  assign _T_54257 = $signed(4'sh1) * $signed(io_in_46); // @[Modules.scala 151:80:@58.4]
  assign _T_54258 = $signed(_T_54255) + $signed(_T_54257); // @[Modules.scala 150:103:@59.4]
  assign _T_54259 = _T_54258[5:0]; // @[Modules.scala 150:103:@60.4]
  assign _T_54260 = $signed(_T_54259); // @[Modules.scala 150:103:@61.4]
  assign _T_54262 = $signed(4'sh1) * $signed(io_in_47); // @[Modules.scala 150:74:@63.4]
  assign _T_54264 = $signed(4'sh1) * $signed(io_in_48); // @[Modules.scala 151:80:@64.4]
  assign _T_54265 = $signed(_T_54262) + $signed(_T_54264); // @[Modules.scala 150:103:@65.4]
  assign _T_54266 = _T_54265[5:0]; // @[Modules.scala 150:103:@66.4]
  assign _T_54267 = $signed(_T_54266); // @[Modules.scala 150:103:@67.4]
  assign _T_54269 = $signed(4'sh1) * $signed(io_in_49); // @[Modules.scala 150:74:@69.4]
  assign _T_54271 = $signed(4'sh1) * $signed(io_in_50); // @[Modules.scala 151:80:@70.4]
  assign _T_54272 = $signed(_T_54269) + $signed(_T_54271); // @[Modules.scala 150:103:@71.4]
  assign _T_54273 = _T_54272[5:0]; // @[Modules.scala 150:103:@72.4]
  assign _T_54274 = $signed(_T_54273); // @[Modules.scala 150:103:@73.4]
  assign _T_54276 = $signed(4'sh1) * $signed(io_in_51); // @[Modules.scala 150:74:@75.4]
  assign _T_54278 = $signed(4'sh1) * $signed(io_in_59); // @[Modules.scala 151:80:@76.4]
  assign _T_54279 = $signed(_T_54276) + $signed(_T_54278); // @[Modules.scala 150:103:@77.4]
  assign _T_54280 = _T_54279[5:0]; // @[Modules.scala 150:103:@78.4]
  assign _T_54281 = $signed(_T_54280); // @[Modules.scala 150:103:@79.4]
  assign _T_54283 = $signed(4'sh1) * $signed(io_in_61); // @[Modules.scala 150:74:@81.4]
  assign _T_54285 = $signed(4'sh1) * $signed(io_in_62); // @[Modules.scala 151:80:@82.4]
  assign _T_54286 = $signed(_T_54283) + $signed(_T_54285); // @[Modules.scala 150:103:@83.4]
  assign _T_54287 = _T_54286[5:0]; // @[Modules.scala 150:103:@84.4]
  assign _T_54288 = $signed(_T_54287); // @[Modules.scala 150:103:@85.4]
  assign _T_54290 = $signed(4'sh1) * $signed(io_in_63); // @[Modules.scala 150:74:@87.4]
  assign _T_54292 = $signed(4'sh1) * $signed(io_in_64); // @[Modules.scala 151:80:@88.4]
  assign _T_54293 = $signed(_T_54290) + $signed(_T_54292); // @[Modules.scala 150:103:@89.4]
  assign _T_54294 = _T_54293[5:0]; // @[Modules.scala 150:103:@90.4]
  assign _T_54295 = $signed(_T_54294); // @[Modules.scala 150:103:@91.4]
  assign _T_54297 = $signed(4'sh1) * $signed(io_in_65); // @[Modules.scala 150:74:@93.4]
  assign _T_54299 = $signed(4'sh1) * $signed(io_in_66); // @[Modules.scala 151:80:@94.4]
  assign _T_54300 = $signed(_T_54297) + $signed(_T_54299); // @[Modules.scala 150:103:@95.4]
  assign _T_54301 = _T_54300[5:0]; // @[Modules.scala 150:103:@96.4]
  assign _T_54302 = $signed(_T_54301); // @[Modules.scala 150:103:@97.4]
  assign _T_54304 = $signed(4'sh1) * $signed(io_in_67); // @[Modules.scala 150:74:@99.4]
  assign _T_54306 = $signed(4'sh1) * $signed(io_in_68); // @[Modules.scala 151:80:@100.4]
  assign _T_54307 = $signed(_T_54304) + $signed(_T_54306); // @[Modules.scala 150:103:@101.4]
  assign _T_54308 = _T_54307[5:0]; // @[Modules.scala 150:103:@102.4]
  assign _T_54309 = $signed(_T_54308); // @[Modules.scala 150:103:@103.4]
  assign _T_54311 = $signed(4'sh1) * $signed(io_in_69); // @[Modules.scala 150:74:@105.4]
  assign _T_54313 = $signed(4'sh1) * $signed(io_in_70); // @[Modules.scala 151:80:@106.4]
  assign _T_54314 = $signed(_T_54311) + $signed(_T_54313); // @[Modules.scala 150:103:@107.4]
  assign _T_54315 = _T_54314[5:0]; // @[Modules.scala 150:103:@108.4]
  assign _T_54316 = $signed(_T_54315); // @[Modules.scala 150:103:@109.4]
  assign _T_54318 = $signed(4'sh1) * $signed(io_in_71); // @[Modules.scala 150:74:@111.4]
  assign _T_54320 = $signed(4'sh1) * $signed(io_in_72); // @[Modules.scala 151:80:@112.4]
  assign _T_54321 = $signed(_T_54318) + $signed(_T_54320); // @[Modules.scala 150:103:@113.4]
  assign _T_54322 = _T_54321[5:0]; // @[Modules.scala 150:103:@114.4]
  assign _T_54323 = $signed(_T_54322); // @[Modules.scala 150:103:@115.4]
  assign _T_54325 = $signed(4'sh1) * $signed(io_in_73); // @[Modules.scala 150:74:@117.4]
  assign _T_54327 = $signed(4'sh1) * $signed(io_in_74); // @[Modules.scala 151:80:@118.4]
  assign _T_54328 = $signed(_T_54325) + $signed(_T_54327); // @[Modules.scala 150:103:@119.4]
  assign _T_54329 = _T_54328[5:0]; // @[Modules.scala 150:103:@120.4]
  assign _T_54330 = $signed(_T_54329); // @[Modules.scala 150:103:@121.4]
  assign _T_54332 = $signed(4'sh1) * $signed(io_in_75); // @[Modules.scala 150:74:@123.4]
  assign _T_54334 = $signed(4'sh1) * $signed(io_in_76); // @[Modules.scala 151:80:@124.4]
  assign _T_54335 = $signed(_T_54332) + $signed(_T_54334); // @[Modules.scala 150:103:@125.4]
  assign _T_54336 = _T_54335[5:0]; // @[Modules.scala 150:103:@126.4]
  assign _T_54337 = $signed(_T_54336); // @[Modules.scala 150:103:@127.4]
  assign _T_54339 = $signed(4'sh1) * $signed(io_in_77); // @[Modules.scala 150:74:@129.4]
  assign _T_54341 = $signed(4'sh1) * $signed(io_in_78); // @[Modules.scala 151:80:@130.4]
  assign _T_54342 = $signed(_T_54339) + $signed(_T_54341); // @[Modules.scala 150:103:@131.4]
  assign _T_54343 = _T_54342[5:0]; // @[Modules.scala 150:103:@132.4]
  assign _T_54344 = $signed(_T_54343); // @[Modules.scala 150:103:@133.4]
  assign _T_54346 = $signed(4'sh1) * $signed(io_in_79); // @[Modules.scala 150:74:@135.4]
  assign _T_54348 = $signed(4'sh1) * $signed(io_in_80); // @[Modules.scala 151:80:@136.4]
  assign _T_54349 = $signed(_T_54346) + $signed(_T_54348); // @[Modules.scala 150:103:@137.4]
  assign _T_54350 = _T_54349[5:0]; // @[Modules.scala 150:103:@138.4]
  assign _T_54351 = $signed(_T_54350); // @[Modules.scala 150:103:@139.4]
  assign _T_54353 = $signed(4'sh1) * $signed(io_in_81); // @[Modules.scala 150:74:@141.4]
  assign _T_54355 = $signed(-4'sh1) * $signed(io_in_86); // @[Modules.scala 151:80:@142.4]
  assign _GEN_1 = {{1{_T_54355[4]}},_T_54355}; // @[Modules.scala 150:103:@143.4]
  assign _T_54356 = $signed(_T_54353) + $signed(_GEN_1); // @[Modules.scala 150:103:@143.4]
  assign _T_54357 = _T_54356[5:0]; // @[Modules.scala 150:103:@144.4]
  assign _T_54358 = $signed(_T_54357); // @[Modules.scala 150:103:@145.4]
  assign _T_54360 = $signed(4'sh1) * $signed(io_in_87); // @[Modules.scala 150:74:@147.4]
  assign _T_54362 = $signed(4'sh1) * $signed(io_in_88); // @[Modules.scala 151:80:@148.4]
  assign _T_54363 = $signed(_T_54360) + $signed(_T_54362); // @[Modules.scala 150:103:@149.4]
  assign _T_54364 = _T_54363[5:0]; // @[Modules.scala 150:103:@150.4]
  assign _T_54365 = $signed(_T_54364); // @[Modules.scala 150:103:@151.4]
  assign _T_54367 = $signed(4'sh1) * $signed(io_in_89); // @[Modules.scala 150:74:@153.4]
  assign _T_54369 = $signed(4'sh1) * $signed(io_in_90); // @[Modules.scala 151:80:@154.4]
  assign _T_54370 = $signed(_T_54367) + $signed(_T_54369); // @[Modules.scala 150:103:@155.4]
  assign _T_54371 = _T_54370[5:0]; // @[Modules.scala 150:103:@156.4]
  assign _T_54372 = $signed(_T_54371); // @[Modules.scala 150:103:@157.4]
  assign _T_54374 = $signed(4'sh1) * $signed(io_in_91); // @[Modules.scala 150:74:@159.4]
  assign _T_54376 = $signed(4'sh1) * $signed(io_in_92); // @[Modules.scala 151:80:@160.4]
  assign _T_54377 = $signed(_T_54374) + $signed(_T_54376); // @[Modules.scala 150:103:@161.4]
  assign _T_54378 = _T_54377[5:0]; // @[Modules.scala 150:103:@162.4]
  assign _T_54379 = $signed(_T_54378); // @[Modules.scala 150:103:@163.4]
  assign _T_54381 = $signed(4'sh1) * $signed(io_in_93); // @[Modules.scala 150:74:@165.4]
  assign _T_54383 = $signed(4'sh1) * $signed(io_in_94); // @[Modules.scala 151:80:@166.4]
  assign _T_54384 = $signed(_T_54381) + $signed(_T_54383); // @[Modules.scala 150:103:@167.4]
  assign _T_54385 = _T_54384[5:0]; // @[Modules.scala 150:103:@168.4]
  assign _T_54386 = $signed(_T_54385); // @[Modules.scala 150:103:@169.4]
  assign _T_54388 = $signed(4'sh1) * $signed(io_in_95); // @[Modules.scala 150:74:@171.4]
  assign _T_54390 = $signed(4'sh1) * $signed(io_in_96); // @[Modules.scala 151:80:@172.4]
  assign _T_54391 = $signed(_T_54388) + $signed(_T_54390); // @[Modules.scala 150:103:@173.4]
  assign _T_54392 = _T_54391[5:0]; // @[Modules.scala 150:103:@174.4]
  assign _T_54393 = $signed(_T_54392); // @[Modules.scala 150:103:@175.4]
  assign _T_54395 = $signed(4'sh1) * $signed(io_in_97); // @[Modules.scala 150:74:@177.4]
  assign _T_54397 = $signed(4'sh1) * $signed(io_in_98); // @[Modules.scala 151:80:@178.4]
  assign _T_54398 = $signed(_T_54395) + $signed(_T_54397); // @[Modules.scala 150:103:@179.4]
  assign _T_54399 = _T_54398[5:0]; // @[Modules.scala 150:103:@180.4]
  assign _T_54400 = $signed(_T_54399); // @[Modules.scala 150:103:@181.4]
  assign _T_54402 = $signed(4'sh1) * $signed(io_in_99); // @[Modules.scala 150:74:@183.4]
  assign _T_54404 = $signed(4'sh1) * $signed(io_in_100); // @[Modules.scala 151:80:@184.4]
  assign _T_54405 = $signed(_T_54402) + $signed(_T_54404); // @[Modules.scala 150:103:@185.4]
  assign _T_54406 = _T_54405[5:0]; // @[Modules.scala 150:103:@186.4]
  assign _T_54407 = $signed(_T_54406); // @[Modules.scala 150:103:@187.4]
  assign _T_54409 = $signed(4'sh1) * $signed(io_in_101); // @[Modules.scala 150:74:@189.4]
  assign _T_54411 = $signed(4'sh1) * $signed(io_in_102); // @[Modules.scala 151:80:@190.4]
  assign _T_54412 = $signed(_T_54409) + $signed(_T_54411); // @[Modules.scala 150:103:@191.4]
  assign _T_54413 = _T_54412[5:0]; // @[Modules.scala 150:103:@192.4]
  assign _T_54414 = $signed(_T_54413); // @[Modules.scala 150:103:@193.4]
  assign _T_54416 = $signed(4'sh1) * $signed(io_in_103); // @[Modules.scala 150:74:@195.4]
  assign _T_54418 = $signed(4'sh1) * $signed(io_in_104); // @[Modules.scala 151:80:@196.4]
  assign _T_54419 = $signed(_T_54416) + $signed(_T_54418); // @[Modules.scala 150:103:@197.4]
  assign _T_54420 = _T_54419[5:0]; // @[Modules.scala 150:103:@198.4]
  assign _T_54421 = $signed(_T_54420); // @[Modules.scala 150:103:@199.4]
  assign _T_54423 = $signed(4'sh1) * $signed(io_in_105); // @[Modules.scala 150:74:@201.4]
  assign _T_54425 = $signed(4'sh1) * $signed(io_in_106); // @[Modules.scala 151:80:@202.4]
  assign _T_54426 = $signed(_T_54423) + $signed(_T_54425); // @[Modules.scala 150:103:@203.4]
  assign _T_54427 = _T_54426[5:0]; // @[Modules.scala 150:103:@204.4]
  assign _T_54428 = $signed(_T_54427); // @[Modules.scala 150:103:@205.4]
  assign _T_54430 = $signed(4'sh1) * $signed(io_in_107); // @[Modules.scala 150:74:@207.4]
  assign _T_54432 = $signed(4'sh1) * $signed(io_in_108); // @[Modules.scala 151:80:@208.4]
  assign _T_54433 = $signed(_T_54430) + $signed(_T_54432); // @[Modules.scala 150:103:@209.4]
  assign _T_54434 = _T_54433[5:0]; // @[Modules.scala 150:103:@210.4]
  assign _T_54435 = $signed(_T_54434); // @[Modules.scala 150:103:@211.4]
  assign _T_54437 = $signed(4'sh1) * $signed(io_in_109); // @[Modules.scala 150:74:@213.4]
  assign _T_54439 = $signed(-4'sh1) * $signed(io_in_110); // @[Modules.scala 151:80:@214.4]
  assign _GEN_2 = {{1{_T_54439[4]}},_T_54439}; // @[Modules.scala 150:103:@215.4]
  assign _T_54440 = $signed(_T_54437) + $signed(_GEN_2); // @[Modules.scala 150:103:@215.4]
  assign _T_54441 = _T_54440[5:0]; // @[Modules.scala 150:103:@216.4]
  assign _T_54442 = $signed(_T_54441); // @[Modules.scala 150:103:@217.4]
  assign _T_54444 = $signed(4'sh1) * $signed(io_in_113); // @[Modules.scala 150:74:@219.4]
  assign _T_54446 = $signed(-4'sh1) * $signed(io_in_114); // @[Modules.scala 151:80:@220.4]
  assign _GEN_3 = {{1{_T_54446[4]}},_T_54446}; // @[Modules.scala 150:103:@221.4]
  assign _T_54447 = $signed(_T_54444) + $signed(_GEN_3); // @[Modules.scala 150:103:@221.4]
  assign _T_54448 = _T_54447[5:0]; // @[Modules.scala 150:103:@222.4]
  assign _T_54449 = $signed(_T_54448); // @[Modules.scala 150:103:@223.4]
  assign _T_54451 = $signed(4'sh1) * $signed(io_in_116); // @[Modules.scala 150:74:@225.4]
  assign _T_54453 = $signed(-4'sh1) * $signed(io_in_117); // @[Modules.scala 151:80:@226.4]
  assign _GEN_4 = {{1{_T_54453[4]}},_T_54453}; // @[Modules.scala 150:103:@227.4]
  assign _T_54454 = $signed(_T_54451) + $signed(_GEN_4); // @[Modules.scala 150:103:@227.4]
  assign _T_54455 = _T_54454[5:0]; // @[Modules.scala 150:103:@228.4]
  assign _T_54456 = $signed(_T_54455); // @[Modules.scala 150:103:@229.4]
  assign _T_54458 = $signed(-4'sh1) * $signed(io_in_118); // @[Modules.scala 150:74:@231.4]
  assign _T_54460 = $signed(4'sh1) * $signed(io_in_120); // @[Modules.scala 151:80:@232.4]
  assign _GEN_5 = {{1{_T_54458[4]}},_T_54458}; // @[Modules.scala 150:103:@233.4]
  assign _T_54461 = $signed(_GEN_5) + $signed(_T_54460); // @[Modules.scala 150:103:@233.4]
  assign _T_54462 = _T_54461[5:0]; // @[Modules.scala 150:103:@234.4]
  assign _T_54463 = $signed(_T_54462); // @[Modules.scala 150:103:@235.4]
  assign _T_54465 = $signed(4'sh1) * $signed(io_in_121); // @[Modules.scala 150:74:@237.4]
  assign _T_54467 = $signed(4'sh1) * $signed(io_in_122); // @[Modules.scala 151:80:@238.4]
  assign _T_54468 = $signed(_T_54465) + $signed(_T_54467); // @[Modules.scala 150:103:@239.4]
  assign _T_54469 = _T_54468[5:0]; // @[Modules.scala 150:103:@240.4]
  assign _T_54470 = $signed(_T_54469); // @[Modules.scala 150:103:@241.4]
  assign _T_54472 = $signed(4'sh1) * $signed(io_in_123); // @[Modules.scala 150:74:@243.4]
  assign _T_54474 = $signed(4'sh1) * $signed(io_in_124); // @[Modules.scala 151:80:@244.4]
  assign _T_54475 = $signed(_T_54472) + $signed(_T_54474); // @[Modules.scala 150:103:@245.4]
  assign _T_54476 = _T_54475[5:0]; // @[Modules.scala 150:103:@246.4]
  assign _T_54477 = $signed(_T_54476); // @[Modules.scala 150:103:@247.4]
  assign _T_54479 = $signed(4'sh1) * $signed(io_in_125); // @[Modules.scala 150:74:@249.4]
  assign _T_54481 = $signed(4'sh1) * $signed(io_in_126); // @[Modules.scala 151:80:@250.4]
  assign _T_54482 = $signed(_T_54479) + $signed(_T_54481); // @[Modules.scala 150:103:@251.4]
  assign _T_54483 = _T_54482[5:0]; // @[Modules.scala 150:103:@252.4]
  assign _T_54484 = $signed(_T_54483); // @[Modules.scala 150:103:@253.4]
  assign _T_54486 = $signed(4'sh1) * $signed(io_in_128); // @[Modules.scala 150:74:@255.4]
  assign _T_54488 = $signed(4'sh1) * $signed(io_in_129); // @[Modules.scala 151:80:@256.4]
  assign _T_54489 = $signed(_T_54486) + $signed(_T_54488); // @[Modules.scala 150:103:@257.4]
  assign _T_54490 = _T_54489[5:0]; // @[Modules.scala 150:103:@258.4]
  assign _T_54491 = $signed(_T_54490); // @[Modules.scala 150:103:@259.4]
  assign _T_54493 = $signed(4'sh1) * $signed(io_in_130); // @[Modules.scala 150:74:@261.4]
  assign _T_54495 = $signed(4'sh1) * $signed(io_in_131); // @[Modules.scala 151:80:@262.4]
  assign _T_54496 = $signed(_T_54493) + $signed(_T_54495); // @[Modules.scala 150:103:@263.4]
  assign _T_54497 = _T_54496[5:0]; // @[Modules.scala 150:103:@264.4]
  assign _T_54498 = $signed(_T_54497); // @[Modules.scala 150:103:@265.4]
  assign _T_54500 = $signed(4'sh1) * $signed(io_in_133); // @[Modules.scala 150:74:@267.4]
  assign _T_54502 = $signed(4'sh1) * $signed(io_in_134); // @[Modules.scala 151:80:@268.4]
  assign _T_54503 = $signed(_T_54500) + $signed(_T_54502); // @[Modules.scala 150:103:@269.4]
  assign _T_54504 = _T_54503[5:0]; // @[Modules.scala 150:103:@270.4]
  assign _T_54505 = $signed(_T_54504); // @[Modules.scala 150:103:@271.4]
  assign _T_54507 = $signed(-4'sh1) * $signed(io_in_135); // @[Modules.scala 150:74:@273.4]
  assign _T_54509 = $signed(-4'sh1) * $signed(io_in_136); // @[Modules.scala 151:80:@274.4]
  assign _T_54510 = $signed(_T_54507) + $signed(_T_54509); // @[Modules.scala 150:103:@275.4]
  assign _T_54511 = _T_54510[4:0]; // @[Modules.scala 150:103:@276.4]
  assign _T_54512 = $signed(_T_54511); // @[Modules.scala 150:103:@277.4]
  assign _T_54514 = $signed(-4'sh1) * $signed(io_in_137); // @[Modules.scala 150:74:@279.4]
  assign _T_54516 = $signed(4'sh1) * $signed(io_in_138); // @[Modules.scala 151:80:@280.4]
  assign _GEN_6 = {{1{_T_54514[4]}},_T_54514}; // @[Modules.scala 150:103:@281.4]
  assign _T_54517 = $signed(_GEN_6) + $signed(_T_54516); // @[Modules.scala 150:103:@281.4]
  assign _T_54518 = _T_54517[5:0]; // @[Modules.scala 150:103:@282.4]
  assign _T_54519 = $signed(_T_54518); // @[Modules.scala 150:103:@283.4]
  assign _T_54521 = $signed(4'sh1) * $signed(io_in_143); // @[Modules.scala 150:74:@285.4]
  assign _T_54523 = $signed(-4'sh1) * $signed(io_in_146); // @[Modules.scala 151:80:@286.4]
  assign _GEN_7 = {{1{_T_54523[4]}},_T_54523}; // @[Modules.scala 150:103:@287.4]
  assign _T_54524 = $signed(_T_54521) + $signed(_GEN_7); // @[Modules.scala 150:103:@287.4]
  assign _T_54525 = _T_54524[5:0]; // @[Modules.scala 150:103:@288.4]
  assign _T_54526 = $signed(_T_54525); // @[Modules.scala 150:103:@289.4]
  assign _T_54528 = $signed(-4'sh1) * $signed(io_in_147); // @[Modules.scala 150:74:@291.4]
  assign _T_54530 = $signed(4'sh1) * $signed(io_in_148); // @[Modules.scala 151:80:@292.4]
  assign _GEN_8 = {{1{_T_54528[4]}},_T_54528}; // @[Modules.scala 150:103:@293.4]
  assign _T_54531 = $signed(_GEN_8) + $signed(_T_54530); // @[Modules.scala 150:103:@293.4]
  assign _T_54532 = _T_54531[5:0]; // @[Modules.scala 150:103:@294.4]
  assign _T_54533 = $signed(_T_54532); // @[Modules.scala 150:103:@295.4]
  assign _T_54535 = $signed(4'sh1) * $signed(io_in_149); // @[Modules.scala 150:74:@297.4]
  assign _T_54537 = $signed(4'sh1) * $signed(io_in_150); // @[Modules.scala 151:80:@298.4]
  assign _T_54538 = $signed(_T_54535) + $signed(_T_54537); // @[Modules.scala 150:103:@299.4]
  assign _T_54539 = _T_54538[5:0]; // @[Modules.scala 150:103:@300.4]
  assign _T_54540 = $signed(_T_54539); // @[Modules.scala 150:103:@301.4]
  assign _T_54542 = $signed(4'sh1) * $signed(io_in_151); // @[Modules.scala 150:74:@303.4]
  assign _T_54544 = $signed(-4'sh1) * $signed(io_in_156); // @[Modules.scala 151:80:@304.4]
  assign _GEN_9 = {{1{_T_54544[4]}},_T_54544}; // @[Modules.scala 150:103:@305.4]
  assign _T_54545 = $signed(_T_54542) + $signed(_GEN_9); // @[Modules.scala 150:103:@305.4]
  assign _T_54546 = _T_54545[5:0]; // @[Modules.scala 150:103:@306.4]
  assign _T_54547 = $signed(_T_54546); // @[Modules.scala 150:103:@307.4]
  assign _T_54549 = $signed(-4'sh1) * $signed(io_in_157); // @[Modules.scala 150:74:@309.4]
  assign _T_54551 = $signed(-4'sh1) * $signed(io_in_160); // @[Modules.scala 151:80:@310.4]
  assign _T_54552 = $signed(_T_54549) + $signed(_T_54551); // @[Modules.scala 150:103:@311.4]
  assign _T_54553 = _T_54552[4:0]; // @[Modules.scala 150:103:@312.4]
  assign _T_54554 = $signed(_T_54553); // @[Modules.scala 150:103:@313.4]
  assign _T_54556 = $signed(4'sh1) * $signed(io_in_161); // @[Modules.scala 150:74:@315.4]
  assign _T_54558 = $signed(-4'sh1) * $signed(io_in_162); // @[Modules.scala 151:80:@316.4]
  assign _GEN_10 = {{1{_T_54558[4]}},_T_54558}; // @[Modules.scala 150:103:@317.4]
  assign _T_54559 = $signed(_T_54556) + $signed(_GEN_10); // @[Modules.scala 150:103:@317.4]
  assign _T_54560 = _T_54559[5:0]; // @[Modules.scala 150:103:@318.4]
  assign _T_54561 = $signed(_T_54560); // @[Modules.scala 150:103:@319.4]
  assign _T_54563 = $signed(-4'sh1) * $signed(io_in_163); // @[Modules.scala 150:74:@321.4]
  assign _T_54565 = $signed(-4'sh1) * $signed(io_in_164); // @[Modules.scala 151:80:@322.4]
  assign _T_54566 = $signed(_T_54563) + $signed(_T_54565); // @[Modules.scala 150:103:@323.4]
  assign _T_54567 = _T_54566[4:0]; // @[Modules.scala 150:103:@324.4]
  assign _T_54568 = $signed(_T_54567); // @[Modules.scala 150:103:@325.4]
  assign _T_54570 = $signed(-4'sh1) * $signed(io_in_165); // @[Modules.scala 150:74:@327.4]
  assign _T_54572 = $signed(4'sh1) * $signed(io_in_166); // @[Modules.scala 151:80:@328.4]
  assign _GEN_11 = {{1{_T_54570[4]}},_T_54570}; // @[Modules.scala 150:103:@329.4]
  assign _T_54573 = $signed(_GEN_11) + $signed(_T_54572); // @[Modules.scala 150:103:@329.4]
  assign _T_54574 = _T_54573[5:0]; // @[Modules.scala 150:103:@330.4]
  assign _T_54575 = $signed(_T_54574); // @[Modules.scala 150:103:@331.4]
  assign _T_54577 = $signed(4'sh1) * $signed(io_in_167); // @[Modules.scala 150:74:@333.4]
  assign _T_54579 = $signed(-4'sh1) * $signed(io_in_169); // @[Modules.scala 151:80:@334.4]
  assign _GEN_12 = {{1{_T_54579[4]}},_T_54579}; // @[Modules.scala 150:103:@335.4]
  assign _T_54580 = $signed(_T_54577) + $signed(_GEN_12); // @[Modules.scala 150:103:@335.4]
  assign _T_54581 = _T_54580[5:0]; // @[Modules.scala 150:103:@336.4]
  assign _T_54582 = $signed(_T_54581); // @[Modules.scala 150:103:@337.4]
  assign _T_54584 = $signed(-4'sh1) * $signed(io_in_170); // @[Modules.scala 150:74:@339.4]
  assign _T_54586 = $signed(4'sh1) * $signed(io_in_171); // @[Modules.scala 151:80:@340.4]
  assign _GEN_13 = {{1{_T_54584[4]}},_T_54584}; // @[Modules.scala 150:103:@341.4]
  assign _T_54587 = $signed(_GEN_13) + $signed(_T_54586); // @[Modules.scala 150:103:@341.4]
  assign _T_54588 = _T_54587[5:0]; // @[Modules.scala 150:103:@342.4]
  assign _T_54589 = $signed(_T_54588); // @[Modules.scala 150:103:@343.4]
  assign _T_54591 = $signed(4'sh1) * $signed(io_in_172); // @[Modules.scala 150:74:@345.4]
  assign _T_54593 = $signed(4'sh1) * $signed(io_in_173); // @[Modules.scala 151:80:@346.4]
  assign _T_54594 = $signed(_T_54591) + $signed(_T_54593); // @[Modules.scala 150:103:@347.4]
  assign _T_54595 = _T_54594[5:0]; // @[Modules.scala 150:103:@348.4]
  assign _T_54596 = $signed(_T_54595); // @[Modules.scala 150:103:@349.4]
  assign _T_54598 = $signed(4'sh1) * $signed(io_in_174); // @[Modules.scala 150:74:@351.4]
  assign _T_54600 = $signed(4'sh1) * $signed(io_in_175); // @[Modules.scala 151:80:@352.4]
  assign _T_54601 = $signed(_T_54598) + $signed(_T_54600); // @[Modules.scala 150:103:@353.4]
  assign _T_54602 = _T_54601[5:0]; // @[Modules.scala 150:103:@354.4]
  assign _T_54603 = $signed(_T_54602); // @[Modules.scala 150:103:@355.4]
  assign _T_54605 = $signed(4'sh1) * $signed(io_in_176); // @[Modules.scala 150:74:@357.4]
  assign _T_54607 = $signed(-4'sh1) * $signed(io_in_178); // @[Modules.scala 151:80:@358.4]
  assign _GEN_14 = {{1{_T_54607[4]}},_T_54607}; // @[Modules.scala 150:103:@359.4]
  assign _T_54608 = $signed(_T_54605) + $signed(_GEN_14); // @[Modules.scala 150:103:@359.4]
  assign _T_54609 = _T_54608[5:0]; // @[Modules.scala 150:103:@360.4]
  assign _T_54610 = $signed(_T_54609); // @[Modules.scala 150:103:@361.4]
  assign _T_54612 = $signed(-4'sh1) * $signed(io_in_180); // @[Modules.scala 150:74:@363.4]
  assign _T_54614 = $signed(-4'sh1) * $signed(io_in_181); // @[Modules.scala 151:80:@364.4]
  assign _T_54615 = $signed(_T_54612) + $signed(_T_54614); // @[Modules.scala 150:103:@365.4]
  assign _T_54616 = _T_54615[4:0]; // @[Modules.scala 150:103:@366.4]
  assign _T_54617 = $signed(_T_54616); // @[Modules.scala 150:103:@367.4]
  assign _T_54619 = $signed(-4'sh1) * $signed(io_in_183); // @[Modules.scala 150:74:@369.4]
  assign _T_54621 = $signed(-4'sh1) * $signed(io_in_184); // @[Modules.scala 151:80:@370.4]
  assign _T_54622 = $signed(_T_54619) + $signed(_T_54621); // @[Modules.scala 150:103:@371.4]
  assign _T_54623 = _T_54622[4:0]; // @[Modules.scala 150:103:@372.4]
  assign _T_54624 = $signed(_T_54623); // @[Modules.scala 150:103:@373.4]
  assign _T_54626 = $signed(-4'sh1) * $signed(io_in_185); // @[Modules.scala 150:74:@375.4]
  assign _T_54628 = $signed(-4'sh1) * $signed(io_in_186); // @[Modules.scala 151:80:@376.4]
  assign _T_54629 = $signed(_T_54626) + $signed(_T_54628); // @[Modules.scala 150:103:@377.4]
  assign _T_54630 = _T_54629[4:0]; // @[Modules.scala 150:103:@378.4]
  assign _T_54631 = $signed(_T_54630); // @[Modules.scala 150:103:@379.4]
  assign _T_54633 = $signed(-4'sh1) * $signed(io_in_187); // @[Modules.scala 150:74:@381.4]
  assign _T_54635 = $signed(-4'sh1) * $signed(io_in_190); // @[Modules.scala 151:80:@382.4]
  assign _T_54636 = $signed(_T_54633) + $signed(_T_54635); // @[Modules.scala 150:103:@383.4]
  assign _T_54637 = _T_54636[4:0]; // @[Modules.scala 150:103:@384.4]
  assign _T_54638 = $signed(_T_54637); // @[Modules.scala 150:103:@385.4]
  assign _T_54640 = $signed(-4'sh1) * $signed(io_in_191); // @[Modules.scala 150:74:@387.4]
  assign _T_54642 = $signed(-4'sh1) * $signed(io_in_192); // @[Modules.scala 151:80:@388.4]
  assign _T_54643 = $signed(_T_54640) + $signed(_T_54642); // @[Modules.scala 150:103:@389.4]
  assign _T_54644 = _T_54643[4:0]; // @[Modules.scala 150:103:@390.4]
  assign _T_54645 = $signed(_T_54644); // @[Modules.scala 150:103:@391.4]
  assign _T_54647 = $signed(-4'sh1) * $signed(io_in_193); // @[Modules.scala 150:74:@393.4]
  assign _T_54649 = $signed(-4'sh1) * $signed(io_in_194); // @[Modules.scala 151:80:@394.4]
  assign _T_54650 = $signed(_T_54647) + $signed(_T_54649); // @[Modules.scala 150:103:@395.4]
  assign _T_54651 = _T_54650[4:0]; // @[Modules.scala 150:103:@396.4]
  assign _T_54652 = $signed(_T_54651); // @[Modules.scala 150:103:@397.4]
  assign _T_54654 = $signed(4'sh1) * $signed(io_in_195); // @[Modules.scala 150:74:@399.4]
  assign _T_54656 = $signed(-4'sh1) * $signed(io_in_196); // @[Modules.scala 151:80:@400.4]
  assign _GEN_15 = {{1{_T_54656[4]}},_T_54656}; // @[Modules.scala 150:103:@401.4]
  assign _T_54657 = $signed(_T_54654) + $signed(_GEN_15); // @[Modules.scala 150:103:@401.4]
  assign _T_54658 = _T_54657[5:0]; // @[Modules.scala 150:103:@402.4]
  assign _T_54659 = $signed(_T_54658); // @[Modules.scala 150:103:@403.4]
  assign _T_54661 = $signed(4'sh1) * $signed(io_in_197); // @[Modules.scala 150:74:@405.4]
  assign _T_54663 = $signed(4'sh1) * $signed(io_in_198); // @[Modules.scala 151:80:@406.4]
  assign _T_54664 = $signed(_T_54661) + $signed(_T_54663); // @[Modules.scala 150:103:@407.4]
  assign _T_54665 = _T_54664[5:0]; // @[Modules.scala 150:103:@408.4]
  assign _T_54666 = $signed(_T_54665); // @[Modules.scala 150:103:@409.4]
  assign _T_54668 = $signed(4'sh1) * $signed(io_in_199); // @[Modules.scala 150:74:@411.4]
  assign _T_54670 = $signed(4'sh1) * $signed(io_in_200); // @[Modules.scala 151:80:@412.4]
  assign _T_54671 = $signed(_T_54668) + $signed(_T_54670); // @[Modules.scala 150:103:@413.4]
  assign _T_54672 = _T_54671[5:0]; // @[Modules.scala 150:103:@414.4]
  assign _T_54673 = $signed(_T_54672); // @[Modules.scala 150:103:@415.4]
  assign _T_54675 = $signed(4'sh1) * $signed(io_in_201); // @[Modules.scala 150:74:@417.4]
  assign _T_54677 = $signed(4'sh1) * $signed(io_in_202); // @[Modules.scala 151:80:@418.4]
  assign _T_54678 = $signed(_T_54675) + $signed(_T_54677); // @[Modules.scala 150:103:@419.4]
  assign _T_54679 = _T_54678[5:0]; // @[Modules.scala 150:103:@420.4]
  assign _T_54680 = $signed(_T_54679); // @[Modules.scala 150:103:@421.4]
  assign _T_54682 = $signed(4'sh1) * $signed(io_in_203); // @[Modules.scala 150:74:@423.4]
  assign _T_54684 = $signed(-4'sh1) * $signed(io_in_205); // @[Modules.scala 151:80:@424.4]
  assign _GEN_16 = {{1{_T_54684[4]}},_T_54684}; // @[Modules.scala 150:103:@425.4]
  assign _T_54685 = $signed(_T_54682) + $signed(_GEN_16); // @[Modules.scala 150:103:@425.4]
  assign _T_54686 = _T_54685[5:0]; // @[Modules.scala 150:103:@426.4]
  assign _T_54687 = $signed(_T_54686); // @[Modules.scala 150:103:@427.4]
  assign _T_54689 = $signed(4'sh1) * $signed(io_in_206); // @[Modules.scala 150:74:@429.4]
  assign _T_54691 = $signed(-4'sh1) * $signed(io_in_212); // @[Modules.scala 151:80:@430.4]
  assign _GEN_17 = {{1{_T_54691[4]}},_T_54691}; // @[Modules.scala 150:103:@431.4]
  assign _T_54692 = $signed(_T_54689) + $signed(_GEN_17); // @[Modules.scala 150:103:@431.4]
  assign _T_54693 = _T_54692[5:0]; // @[Modules.scala 150:103:@432.4]
  assign _T_54694 = $signed(_T_54693); // @[Modules.scala 150:103:@433.4]
  assign _T_54696 = $signed(-4'sh1) * $signed(io_in_213); // @[Modules.scala 150:74:@435.4]
  assign _T_54698 = $signed(-4'sh1) * $signed(io_in_214); // @[Modules.scala 151:80:@436.4]
  assign _T_54699 = $signed(_T_54696) + $signed(_T_54698); // @[Modules.scala 150:103:@437.4]
  assign _T_54700 = _T_54699[4:0]; // @[Modules.scala 150:103:@438.4]
  assign _T_54701 = $signed(_T_54700); // @[Modules.scala 150:103:@439.4]
  assign _T_54703 = $signed(-4'sh1) * $signed(io_in_216); // @[Modules.scala 150:74:@441.4]
  assign _T_54705 = $signed(-4'sh1) * $signed(io_in_217); // @[Modules.scala 151:80:@442.4]
  assign _T_54706 = $signed(_T_54703) + $signed(_T_54705); // @[Modules.scala 150:103:@443.4]
  assign _T_54707 = _T_54706[4:0]; // @[Modules.scala 150:103:@444.4]
  assign _T_54708 = $signed(_T_54707); // @[Modules.scala 150:103:@445.4]
  assign _T_54710 = $signed(-4'sh1) * $signed(io_in_218); // @[Modules.scala 150:74:@447.4]
  assign _T_54712 = $signed(-4'sh1) * $signed(io_in_219); // @[Modules.scala 151:80:@448.4]
  assign _T_54713 = $signed(_T_54710) + $signed(_T_54712); // @[Modules.scala 150:103:@449.4]
  assign _T_54714 = _T_54713[4:0]; // @[Modules.scala 150:103:@450.4]
  assign _T_54715 = $signed(_T_54714); // @[Modules.scala 150:103:@451.4]
  assign _T_54717 = $signed(-4'sh1) * $signed(io_in_220); // @[Modules.scala 150:74:@453.4]
  assign _T_54719 = $signed(-4'sh1) * $signed(io_in_221); // @[Modules.scala 151:80:@454.4]
  assign _T_54720 = $signed(_T_54717) + $signed(_T_54719); // @[Modules.scala 150:103:@455.4]
  assign _T_54721 = _T_54720[4:0]; // @[Modules.scala 150:103:@456.4]
  assign _T_54722 = $signed(_T_54721); // @[Modules.scala 150:103:@457.4]
  assign _T_54724 = $signed(4'sh1) * $signed(io_in_223); // @[Modules.scala 150:74:@459.4]
  assign _T_54726 = $signed(-4'sh1) * $signed(io_in_224); // @[Modules.scala 151:80:@460.4]
  assign _GEN_18 = {{1{_T_54726[4]}},_T_54726}; // @[Modules.scala 150:103:@461.4]
  assign _T_54727 = $signed(_T_54724) + $signed(_GEN_18); // @[Modules.scala 150:103:@461.4]
  assign _T_54728 = _T_54727[5:0]; // @[Modules.scala 150:103:@462.4]
  assign _T_54729 = $signed(_T_54728); // @[Modules.scala 150:103:@463.4]
  assign _T_54731 = $signed(4'sh1) * $signed(io_in_225); // @[Modules.scala 150:74:@465.4]
  assign _T_54733 = $signed(4'sh1) * $signed(io_in_226); // @[Modules.scala 151:80:@466.4]
  assign _T_54734 = $signed(_T_54731) + $signed(_T_54733); // @[Modules.scala 150:103:@467.4]
  assign _T_54735 = _T_54734[5:0]; // @[Modules.scala 150:103:@468.4]
  assign _T_54736 = $signed(_T_54735); // @[Modules.scala 150:103:@469.4]
  assign _T_54738 = $signed(4'sh1) * $signed(io_in_227); // @[Modules.scala 150:74:@471.4]
  assign _T_54740 = $signed(4'sh1) * $signed(io_in_228); // @[Modules.scala 151:80:@472.4]
  assign _T_54741 = $signed(_T_54738) + $signed(_T_54740); // @[Modules.scala 150:103:@473.4]
  assign _T_54742 = _T_54741[5:0]; // @[Modules.scala 150:103:@474.4]
  assign _T_54743 = $signed(_T_54742); // @[Modules.scala 150:103:@475.4]
  assign _T_54745 = $signed(4'sh1) * $signed(io_in_229); // @[Modules.scala 150:74:@477.4]
  assign _T_54747 = $signed(4'sh1) * $signed(io_in_230); // @[Modules.scala 151:80:@478.4]
  assign _T_54748 = $signed(_T_54745) + $signed(_T_54747); // @[Modules.scala 150:103:@479.4]
  assign _T_54749 = _T_54748[5:0]; // @[Modules.scala 150:103:@480.4]
  assign _T_54750 = $signed(_T_54749); // @[Modules.scala 150:103:@481.4]
  assign _T_54752 = $signed(4'sh1) * $signed(io_in_231); // @[Modules.scala 150:74:@483.4]
  assign _T_54754 = $signed(4'sh1) * $signed(io_in_232); // @[Modules.scala 151:80:@484.4]
  assign _T_54755 = $signed(_T_54752) + $signed(_T_54754); // @[Modules.scala 150:103:@485.4]
  assign _T_54756 = _T_54755[5:0]; // @[Modules.scala 150:103:@486.4]
  assign _T_54757 = $signed(_T_54756); // @[Modules.scala 150:103:@487.4]
  assign _T_54759 = $signed(-4'sh1) * $signed(io_in_233); // @[Modules.scala 150:74:@489.4]
  assign _T_54761 = $signed(4'sh1) * $signed(io_in_235); // @[Modules.scala 151:80:@490.4]
  assign _GEN_19 = {{1{_T_54759[4]}},_T_54759}; // @[Modules.scala 150:103:@491.4]
  assign _T_54762 = $signed(_GEN_19) + $signed(_T_54761); // @[Modules.scala 150:103:@491.4]
  assign _T_54763 = _T_54762[5:0]; // @[Modules.scala 150:103:@492.4]
  assign _T_54764 = $signed(_T_54763); // @[Modules.scala 150:103:@493.4]
  assign _T_54766 = $signed(4'sh1) * $signed(io_in_238); // @[Modules.scala 150:74:@495.4]
  assign _T_54768 = $signed(-4'sh1) * $signed(io_in_240); // @[Modules.scala 151:80:@496.4]
  assign _GEN_20 = {{1{_T_54768[4]}},_T_54768}; // @[Modules.scala 150:103:@497.4]
  assign _T_54769 = $signed(_T_54766) + $signed(_GEN_20); // @[Modules.scala 150:103:@497.4]
  assign _T_54770 = _T_54769[5:0]; // @[Modules.scala 150:103:@498.4]
  assign _T_54771 = $signed(_T_54770); // @[Modules.scala 150:103:@499.4]
  assign _T_54773 = $signed(-4'sh1) * $signed(io_in_241); // @[Modules.scala 150:74:@501.4]
  assign _T_54775 = $signed(-4'sh1) * $signed(io_in_242); // @[Modules.scala 151:80:@502.4]
  assign _T_54776 = $signed(_T_54773) + $signed(_T_54775); // @[Modules.scala 150:103:@503.4]
  assign _T_54777 = _T_54776[4:0]; // @[Modules.scala 150:103:@504.4]
  assign _T_54778 = $signed(_T_54777); // @[Modules.scala 150:103:@505.4]
  assign _T_54780 = $signed(-4'sh1) * $signed(io_in_243); // @[Modules.scala 150:74:@507.4]
  assign _T_54782 = $signed(-4'sh1) * $signed(io_in_244); // @[Modules.scala 151:80:@508.4]
  assign _T_54783 = $signed(_T_54780) + $signed(_T_54782); // @[Modules.scala 150:103:@509.4]
  assign _T_54784 = _T_54783[4:0]; // @[Modules.scala 150:103:@510.4]
  assign _T_54785 = $signed(_T_54784); // @[Modules.scala 150:103:@511.4]
  assign _T_54787 = $signed(-4'sh1) * $signed(io_in_245); // @[Modules.scala 150:74:@513.4]
  assign _T_54789 = $signed(-4'sh1) * $signed(io_in_246); // @[Modules.scala 151:80:@514.4]
  assign _T_54790 = $signed(_T_54787) + $signed(_T_54789); // @[Modules.scala 150:103:@515.4]
  assign _T_54791 = _T_54790[4:0]; // @[Modules.scala 150:103:@516.4]
  assign _T_54792 = $signed(_T_54791); // @[Modules.scala 150:103:@517.4]
  assign _T_54794 = $signed(-4'sh1) * $signed(io_in_247); // @[Modules.scala 150:74:@519.4]
  assign _T_54796 = $signed(-4'sh1) * $signed(io_in_248); // @[Modules.scala 151:80:@520.4]
  assign _T_54797 = $signed(_T_54794) + $signed(_T_54796); // @[Modules.scala 150:103:@521.4]
  assign _T_54798 = _T_54797[4:0]; // @[Modules.scala 150:103:@522.4]
  assign _T_54799 = $signed(_T_54798); // @[Modules.scala 150:103:@523.4]
  assign _T_54801 = $signed(-4'sh1) * $signed(io_in_249); // @[Modules.scala 150:74:@525.4]
  assign _T_54803 = $signed(-4'sh1) * $signed(io_in_250); // @[Modules.scala 151:80:@526.4]
  assign _T_54804 = $signed(_T_54801) + $signed(_T_54803); // @[Modules.scala 150:103:@527.4]
  assign _T_54805 = _T_54804[4:0]; // @[Modules.scala 150:103:@528.4]
  assign _T_54806 = $signed(_T_54805); // @[Modules.scala 150:103:@529.4]
  assign _T_54808 = $signed(4'sh1) * $signed(io_in_251); // @[Modules.scala 150:74:@531.4]
  assign _T_54810 = $signed(-4'sh1) * $signed(io_in_252); // @[Modules.scala 151:80:@532.4]
  assign _GEN_21 = {{1{_T_54810[4]}},_T_54810}; // @[Modules.scala 150:103:@533.4]
  assign _T_54811 = $signed(_T_54808) + $signed(_GEN_21); // @[Modules.scala 150:103:@533.4]
  assign _T_54812 = _T_54811[5:0]; // @[Modules.scala 150:103:@534.4]
  assign _T_54813 = $signed(_T_54812); // @[Modules.scala 150:103:@535.4]
  assign _T_54815 = $signed(4'sh1) * $signed(io_in_253); // @[Modules.scala 150:74:@537.4]
  assign _T_54817 = $signed(4'sh1) * $signed(io_in_254); // @[Modules.scala 151:80:@538.4]
  assign _T_54818 = $signed(_T_54815) + $signed(_T_54817); // @[Modules.scala 150:103:@539.4]
  assign _T_54819 = _T_54818[5:0]; // @[Modules.scala 150:103:@540.4]
  assign _T_54820 = $signed(_T_54819); // @[Modules.scala 150:103:@541.4]
  assign _T_54822 = $signed(4'sh1) * $signed(io_in_256); // @[Modules.scala 150:74:@543.4]
  assign _T_54824 = $signed(4'sh1) * $signed(io_in_260); // @[Modules.scala 151:80:@544.4]
  assign _T_54825 = $signed(_T_54822) + $signed(_T_54824); // @[Modules.scala 150:103:@545.4]
  assign _T_54826 = _T_54825[5:0]; // @[Modules.scala 150:103:@546.4]
  assign _T_54827 = $signed(_T_54826); // @[Modules.scala 150:103:@547.4]
  assign _T_54829 = $signed(-4'sh1) * $signed(io_in_261); // @[Modules.scala 150:74:@549.4]
  assign _T_54831 = $signed(-4'sh1) * $signed(io_in_262); // @[Modules.scala 151:80:@550.4]
  assign _T_54832 = $signed(_T_54829) + $signed(_T_54831); // @[Modules.scala 150:103:@551.4]
  assign _T_54833 = _T_54832[4:0]; // @[Modules.scala 150:103:@552.4]
  assign _T_54834 = $signed(_T_54833); // @[Modules.scala 150:103:@553.4]
  assign _T_54836 = $signed(-4'sh1) * $signed(io_in_263); // @[Modules.scala 150:74:@555.4]
  assign _T_54838 = $signed(-4'sh1) * $signed(io_in_264); // @[Modules.scala 151:80:@556.4]
  assign _T_54839 = $signed(_T_54836) + $signed(_T_54838); // @[Modules.scala 150:103:@557.4]
  assign _T_54840 = _T_54839[4:0]; // @[Modules.scala 150:103:@558.4]
  assign _T_54841 = $signed(_T_54840); // @[Modules.scala 150:103:@559.4]
  assign _T_54843 = $signed(-4'sh1) * $signed(io_in_265); // @[Modules.scala 150:74:@561.4]
  assign _T_54845 = $signed(4'sh1) * $signed(io_in_266); // @[Modules.scala 151:80:@562.4]
  assign _GEN_22 = {{1{_T_54843[4]}},_T_54843}; // @[Modules.scala 150:103:@563.4]
  assign _T_54846 = $signed(_GEN_22) + $signed(_T_54845); // @[Modules.scala 150:103:@563.4]
  assign _T_54847 = _T_54846[5:0]; // @[Modules.scala 150:103:@564.4]
  assign _T_54848 = $signed(_T_54847); // @[Modules.scala 150:103:@565.4]
  assign _T_54850 = $signed(4'sh1) * $signed(io_in_267); // @[Modules.scala 150:74:@567.4]
  assign _T_54852 = $signed(-4'sh1) * $signed(io_in_268); // @[Modules.scala 151:80:@568.4]
  assign _GEN_23 = {{1{_T_54852[4]}},_T_54852}; // @[Modules.scala 150:103:@569.4]
  assign _T_54853 = $signed(_T_54850) + $signed(_GEN_23); // @[Modules.scala 150:103:@569.4]
  assign _T_54854 = _T_54853[5:0]; // @[Modules.scala 150:103:@570.4]
  assign _T_54855 = $signed(_T_54854); // @[Modules.scala 150:103:@571.4]
  assign _T_54857 = $signed(-4'sh1) * $signed(io_in_269); // @[Modules.scala 150:74:@573.4]
  assign _T_54859 = $signed(-4'sh1) * $signed(io_in_270); // @[Modules.scala 151:80:@574.4]
  assign _T_54860 = $signed(_T_54857) + $signed(_T_54859); // @[Modules.scala 150:103:@575.4]
  assign _T_54861 = _T_54860[4:0]; // @[Modules.scala 150:103:@576.4]
  assign _T_54862 = $signed(_T_54861); // @[Modules.scala 150:103:@577.4]
  assign _T_54864 = $signed(-4'sh1) * $signed(io_in_271); // @[Modules.scala 150:74:@579.4]
  assign _T_54866 = $signed(-4'sh1) * $signed(io_in_272); // @[Modules.scala 151:80:@580.4]
  assign _T_54867 = $signed(_T_54864) + $signed(_T_54866); // @[Modules.scala 150:103:@581.4]
  assign _T_54868 = _T_54867[4:0]; // @[Modules.scala 150:103:@582.4]
  assign _T_54869 = $signed(_T_54868); // @[Modules.scala 150:103:@583.4]
  assign _T_54871 = $signed(-4'sh1) * $signed(io_in_273); // @[Modules.scala 150:74:@585.4]
  assign _T_54873 = $signed(-4'sh1) * $signed(io_in_274); // @[Modules.scala 151:80:@586.4]
  assign _T_54874 = $signed(_T_54871) + $signed(_T_54873); // @[Modules.scala 150:103:@587.4]
  assign _T_54875 = _T_54874[4:0]; // @[Modules.scala 150:103:@588.4]
  assign _T_54876 = $signed(_T_54875); // @[Modules.scala 150:103:@589.4]
  assign _T_54878 = $signed(-4'sh1) * $signed(io_in_275); // @[Modules.scala 150:74:@591.4]
  assign _T_54880 = $signed(-4'sh1) * $signed(io_in_276); // @[Modules.scala 151:80:@592.4]
  assign _T_54881 = $signed(_T_54878) + $signed(_T_54880); // @[Modules.scala 150:103:@593.4]
  assign _T_54882 = _T_54881[4:0]; // @[Modules.scala 150:103:@594.4]
  assign _T_54883 = $signed(_T_54882); // @[Modules.scala 150:103:@595.4]
  assign _T_54885 = $signed(-4'sh1) * $signed(io_in_277); // @[Modules.scala 150:74:@597.4]
  assign _T_54887 = $signed(-4'sh1) * $signed(io_in_278); // @[Modules.scala 151:80:@598.4]
  assign _T_54888 = $signed(_T_54885) + $signed(_T_54887); // @[Modules.scala 150:103:@599.4]
  assign _T_54889 = _T_54888[4:0]; // @[Modules.scala 150:103:@600.4]
  assign _T_54890 = $signed(_T_54889); // @[Modules.scala 150:103:@601.4]
  assign _T_54892 = $signed(-4'sh1) * $signed(io_in_279); // @[Modules.scala 150:74:@603.4]
  assign _T_54894 = $signed(-4'sh1) * $signed(io_in_280); // @[Modules.scala 151:80:@604.4]
  assign _T_54895 = $signed(_T_54892) + $signed(_T_54894); // @[Modules.scala 150:103:@605.4]
  assign _T_54896 = _T_54895[4:0]; // @[Modules.scala 150:103:@606.4]
  assign _T_54897 = $signed(_T_54896); // @[Modules.scala 150:103:@607.4]
  assign _T_54899 = $signed(4'sh1) * $signed(io_in_281); // @[Modules.scala 150:74:@609.4]
  assign _T_54901 = $signed(4'sh1) * $signed(io_in_282); // @[Modules.scala 151:80:@610.4]
  assign _T_54902 = $signed(_T_54899) + $signed(_T_54901); // @[Modules.scala 150:103:@611.4]
  assign _T_54903 = _T_54902[5:0]; // @[Modules.scala 150:103:@612.4]
  assign _T_54904 = $signed(_T_54903); // @[Modules.scala 150:103:@613.4]
  assign _T_54906 = $signed(4'sh1) * $signed(io_in_283); // @[Modules.scala 150:74:@615.4]
  assign _T_54908 = $signed(-4'sh1) * $signed(io_in_284); // @[Modules.scala 151:80:@616.4]
  assign _GEN_24 = {{1{_T_54908[4]}},_T_54908}; // @[Modules.scala 150:103:@617.4]
  assign _T_54909 = $signed(_T_54906) + $signed(_GEN_24); // @[Modules.scala 150:103:@617.4]
  assign _T_54910 = _T_54909[5:0]; // @[Modules.scala 150:103:@618.4]
  assign _T_54911 = $signed(_T_54910); // @[Modules.scala 150:103:@619.4]
  assign _T_54913 = $signed(-4'sh1) * $signed(io_in_285); // @[Modules.scala 150:74:@621.4]
  assign _T_54915 = $signed(-4'sh1) * $signed(io_in_286); // @[Modules.scala 151:80:@622.4]
  assign _T_54916 = $signed(_T_54913) + $signed(_T_54915); // @[Modules.scala 150:103:@623.4]
  assign _T_54917 = _T_54916[4:0]; // @[Modules.scala 150:103:@624.4]
  assign _T_54918 = $signed(_T_54917); // @[Modules.scala 150:103:@625.4]
  assign _T_54920 = $signed(-4'sh1) * $signed(io_in_287); // @[Modules.scala 150:74:@627.4]
  assign _T_54922 = $signed(-4'sh1) * $signed(io_in_288); // @[Modules.scala 151:80:@628.4]
  assign _T_54923 = $signed(_T_54920) + $signed(_T_54922); // @[Modules.scala 150:103:@629.4]
  assign _T_54924 = _T_54923[4:0]; // @[Modules.scala 150:103:@630.4]
  assign _T_54925 = $signed(_T_54924); // @[Modules.scala 150:103:@631.4]
  assign _T_54927 = $signed(-4'sh1) * $signed(io_in_289); // @[Modules.scala 150:74:@633.4]
  assign _T_54929 = $signed(-4'sh1) * $signed(io_in_290); // @[Modules.scala 151:80:@634.4]
  assign _T_54930 = $signed(_T_54927) + $signed(_T_54929); // @[Modules.scala 150:103:@635.4]
  assign _T_54931 = _T_54930[4:0]; // @[Modules.scala 150:103:@636.4]
  assign _T_54932 = $signed(_T_54931); // @[Modules.scala 150:103:@637.4]
  assign _T_54934 = $signed(-4'sh1) * $signed(io_in_291); // @[Modules.scala 150:74:@639.4]
  assign _T_54936 = $signed(-4'sh1) * $signed(io_in_292); // @[Modules.scala 151:80:@640.4]
  assign _T_54937 = $signed(_T_54934) + $signed(_T_54936); // @[Modules.scala 150:103:@641.4]
  assign _T_54938 = _T_54937[4:0]; // @[Modules.scala 150:103:@642.4]
  assign _T_54939 = $signed(_T_54938); // @[Modules.scala 150:103:@643.4]
  assign _T_54941 = $signed(-4'sh1) * $signed(io_in_293); // @[Modules.scala 150:74:@645.4]
  assign _T_54943 = $signed(4'sh1) * $signed(io_in_294); // @[Modules.scala 151:80:@646.4]
  assign _GEN_25 = {{1{_T_54941[4]}},_T_54941}; // @[Modules.scala 150:103:@647.4]
  assign _T_54944 = $signed(_GEN_25) + $signed(_T_54943); // @[Modules.scala 150:103:@647.4]
  assign _T_54945 = _T_54944[5:0]; // @[Modules.scala 150:103:@648.4]
  assign _T_54946 = $signed(_T_54945); // @[Modules.scala 150:103:@649.4]
  assign _T_54948 = $signed(4'sh1) * $signed(io_in_295); // @[Modules.scala 150:74:@651.4]
  assign _T_54950 = $signed(4'sh1) * $signed(io_in_296); // @[Modules.scala 151:80:@652.4]
  assign _T_54951 = $signed(_T_54948) + $signed(_T_54950); // @[Modules.scala 150:103:@653.4]
  assign _T_54952 = _T_54951[5:0]; // @[Modules.scala 150:103:@654.4]
  assign _T_54953 = $signed(_T_54952); // @[Modules.scala 150:103:@655.4]
  assign _T_54955 = $signed(-4'sh1) * $signed(io_in_298); // @[Modules.scala 150:74:@657.4]
  assign _T_54957 = $signed(-4'sh1) * $signed(io_in_299); // @[Modules.scala 151:80:@658.4]
  assign _T_54958 = $signed(_T_54955) + $signed(_T_54957); // @[Modules.scala 150:103:@659.4]
  assign _T_54959 = _T_54958[4:0]; // @[Modules.scala 150:103:@660.4]
  assign _T_54960 = $signed(_T_54959); // @[Modules.scala 150:103:@661.4]
  assign _T_54962 = $signed(-4'sh1) * $signed(io_in_300); // @[Modules.scala 150:74:@663.4]
  assign _T_54964 = $signed(-4'sh1) * $signed(io_in_301); // @[Modules.scala 151:80:@664.4]
  assign _T_54965 = $signed(_T_54962) + $signed(_T_54964); // @[Modules.scala 150:103:@665.4]
  assign _T_54966 = _T_54965[4:0]; // @[Modules.scala 150:103:@666.4]
  assign _T_54967 = $signed(_T_54966); // @[Modules.scala 150:103:@667.4]
  assign _T_54969 = $signed(-4'sh1) * $signed(io_in_302); // @[Modules.scala 150:74:@669.4]
  assign _T_54971 = $signed(-4'sh1) * $signed(io_in_303); // @[Modules.scala 151:80:@670.4]
  assign _T_54972 = $signed(_T_54969) + $signed(_T_54971); // @[Modules.scala 150:103:@671.4]
  assign _T_54973 = _T_54972[4:0]; // @[Modules.scala 150:103:@672.4]
  assign _T_54974 = $signed(_T_54973); // @[Modules.scala 150:103:@673.4]
  assign _T_54976 = $signed(-4'sh1) * $signed(io_in_304); // @[Modules.scala 150:74:@675.4]
  assign _T_54978 = $signed(-4'sh1) * $signed(io_in_305); // @[Modules.scala 151:80:@676.4]
  assign _T_54979 = $signed(_T_54976) + $signed(_T_54978); // @[Modules.scala 150:103:@677.4]
  assign _T_54980 = _T_54979[4:0]; // @[Modules.scala 150:103:@678.4]
  assign _T_54981 = $signed(_T_54980); // @[Modules.scala 150:103:@679.4]
  assign _T_54983 = $signed(-4'sh1) * $signed(io_in_306); // @[Modules.scala 150:74:@681.4]
  assign _T_54985 = $signed(-4'sh1) * $signed(io_in_308); // @[Modules.scala 151:80:@682.4]
  assign _T_54986 = $signed(_T_54983) + $signed(_T_54985); // @[Modules.scala 150:103:@683.4]
  assign _T_54987 = _T_54986[4:0]; // @[Modules.scala 150:103:@684.4]
  assign _T_54988 = $signed(_T_54987); // @[Modules.scala 150:103:@685.4]
  assign _T_54990 = $signed(4'sh1) * $signed(io_in_309); // @[Modules.scala 150:74:@687.4]
  assign _T_54992 = $signed(-4'sh1) * $signed(io_in_310); // @[Modules.scala 151:80:@688.4]
  assign _GEN_26 = {{1{_T_54992[4]}},_T_54992}; // @[Modules.scala 150:103:@689.4]
  assign _T_54993 = $signed(_T_54990) + $signed(_GEN_26); // @[Modules.scala 150:103:@689.4]
  assign _T_54994 = _T_54993[5:0]; // @[Modules.scala 150:103:@690.4]
  assign _T_54995 = $signed(_T_54994); // @[Modules.scala 150:103:@691.4]
  assign _T_54997 = $signed(4'sh1) * $signed(io_in_311); // @[Modules.scala 150:74:@693.4]
  assign _T_54999 = $signed(-4'sh1) * $signed(io_in_312); // @[Modules.scala 151:80:@694.4]
  assign _GEN_27 = {{1{_T_54999[4]}},_T_54999}; // @[Modules.scala 150:103:@695.4]
  assign _T_55000 = $signed(_T_54997) + $signed(_GEN_27); // @[Modules.scala 150:103:@695.4]
  assign _T_55001 = _T_55000[5:0]; // @[Modules.scala 150:103:@696.4]
  assign _T_55002 = $signed(_T_55001); // @[Modules.scala 150:103:@697.4]
  assign _T_55004 = $signed(-4'sh1) * $signed(io_in_313); // @[Modules.scala 150:74:@699.4]
  assign _T_55006 = $signed(-4'sh1) * $signed(io_in_314); // @[Modules.scala 151:80:@700.4]
  assign _T_55007 = $signed(_T_55004) + $signed(_T_55006); // @[Modules.scala 150:103:@701.4]
  assign _T_55008 = _T_55007[4:0]; // @[Modules.scala 150:103:@702.4]
  assign _T_55009 = $signed(_T_55008); // @[Modules.scala 150:103:@703.4]
  assign _T_55011 = $signed(-4'sh1) * $signed(io_in_315); // @[Modules.scala 150:74:@705.4]
  assign _T_55013 = $signed(-4'sh1) * $signed(io_in_316); // @[Modules.scala 151:80:@706.4]
  assign _T_55014 = $signed(_T_55011) + $signed(_T_55013); // @[Modules.scala 150:103:@707.4]
  assign _T_55015 = _T_55014[4:0]; // @[Modules.scala 150:103:@708.4]
  assign _T_55016 = $signed(_T_55015); // @[Modules.scala 150:103:@709.4]
  assign _T_55018 = $signed(-4'sh1) * $signed(io_in_317); // @[Modules.scala 150:74:@711.4]
  assign _T_55020 = $signed(-4'sh1) * $signed(io_in_318); // @[Modules.scala 151:80:@712.4]
  assign _T_55021 = $signed(_T_55018) + $signed(_T_55020); // @[Modules.scala 150:103:@713.4]
  assign _T_55022 = _T_55021[4:0]; // @[Modules.scala 150:103:@714.4]
  assign _T_55023 = $signed(_T_55022); // @[Modules.scala 150:103:@715.4]
  assign _T_55025 = $signed(-4'sh1) * $signed(io_in_319); // @[Modules.scala 150:74:@717.4]
  assign _T_55027 = $signed(-4'sh1) * $signed(io_in_320); // @[Modules.scala 151:80:@718.4]
  assign _T_55028 = $signed(_T_55025) + $signed(_T_55027); // @[Modules.scala 150:103:@719.4]
  assign _T_55029 = _T_55028[4:0]; // @[Modules.scala 150:103:@720.4]
  assign _T_55030 = $signed(_T_55029); // @[Modules.scala 150:103:@721.4]
  assign _T_55032 = $signed(-4'sh1) * $signed(io_in_321); // @[Modules.scala 150:74:@723.4]
  assign _T_55034 = $signed(4'sh1) * $signed(io_in_323); // @[Modules.scala 151:80:@724.4]
  assign _GEN_28 = {{1{_T_55032[4]}},_T_55032}; // @[Modules.scala 150:103:@725.4]
  assign _T_55035 = $signed(_GEN_28) + $signed(_T_55034); // @[Modules.scala 150:103:@725.4]
  assign _T_55036 = _T_55035[5:0]; // @[Modules.scala 150:103:@726.4]
  assign _T_55037 = $signed(_T_55036); // @[Modules.scala 150:103:@727.4]
  assign _T_55039 = $signed(-4'sh1) * $signed(io_in_324); // @[Modules.scala 150:74:@729.4]
  assign _T_55041 = $signed(-4'sh1) * $signed(io_in_325); // @[Modules.scala 151:80:@730.4]
  assign _T_55042 = $signed(_T_55039) + $signed(_T_55041); // @[Modules.scala 150:103:@731.4]
  assign _T_55043 = _T_55042[4:0]; // @[Modules.scala 150:103:@732.4]
  assign _T_55044 = $signed(_T_55043); // @[Modules.scala 150:103:@733.4]
  assign _T_55046 = $signed(-4'sh1) * $signed(io_in_326); // @[Modules.scala 150:74:@735.4]
  assign _T_55048 = $signed(-4'sh1) * $signed(io_in_327); // @[Modules.scala 151:80:@736.4]
  assign _T_55049 = $signed(_T_55046) + $signed(_T_55048); // @[Modules.scala 150:103:@737.4]
  assign _T_55050 = _T_55049[4:0]; // @[Modules.scala 150:103:@738.4]
  assign _T_55051 = $signed(_T_55050); // @[Modules.scala 150:103:@739.4]
  assign _T_55053 = $signed(-4'sh1) * $signed(io_in_328); // @[Modules.scala 150:74:@741.4]
  assign _T_55055 = $signed(-4'sh1) * $signed(io_in_329); // @[Modules.scala 151:80:@742.4]
  assign _T_55056 = $signed(_T_55053) + $signed(_T_55055); // @[Modules.scala 150:103:@743.4]
  assign _T_55057 = _T_55056[4:0]; // @[Modules.scala 150:103:@744.4]
  assign _T_55058 = $signed(_T_55057); // @[Modules.scala 150:103:@745.4]
  assign _T_55060 = $signed(-4'sh1) * $signed(io_in_330); // @[Modules.scala 150:74:@747.4]
  assign _T_55062 = $signed(-4'sh1) * $signed(io_in_331); // @[Modules.scala 151:80:@748.4]
  assign _T_55063 = $signed(_T_55060) + $signed(_T_55062); // @[Modules.scala 150:103:@749.4]
  assign _T_55064 = _T_55063[4:0]; // @[Modules.scala 150:103:@750.4]
  assign _T_55065 = $signed(_T_55064); // @[Modules.scala 150:103:@751.4]
  assign _T_55067 = $signed(-4'sh1) * $signed(io_in_332); // @[Modules.scala 150:74:@753.4]
  assign _T_55069 = $signed(-4'sh1) * $signed(io_in_333); // @[Modules.scala 151:80:@754.4]
  assign _T_55070 = $signed(_T_55067) + $signed(_T_55069); // @[Modules.scala 150:103:@755.4]
  assign _T_55071 = _T_55070[4:0]; // @[Modules.scala 150:103:@756.4]
  assign _T_55072 = $signed(_T_55071); // @[Modules.scala 150:103:@757.4]
  assign _T_55074 = $signed(-4'sh1) * $signed(io_in_336); // @[Modules.scala 150:74:@759.4]
  assign _T_55076 = $signed(4'sh1) * $signed(io_in_337); // @[Modules.scala 151:80:@760.4]
  assign _GEN_29 = {{1{_T_55074[4]}},_T_55074}; // @[Modules.scala 150:103:@761.4]
  assign _T_55077 = $signed(_GEN_29) + $signed(_T_55076); // @[Modules.scala 150:103:@761.4]
  assign _T_55078 = _T_55077[5:0]; // @[Modules.scala 150:103:@762.4]
  assign _T_55079 = $signed(_T_55078); // @[Modules.scala 150:103:@763.4]
  assign _T_55081 = $signed(4'sh1) * $signed(io_in_338); // @[Modules.scala 150:74:@765.4]
  assign _T_55083 = $signed(4'sh1) * $signed(io_in_339); // @[Modules.scala 151:80:@766.4]
  assign _T_55084 = $signed(_T_55081) + $signed(_T_55083); // @[Modules.scala 150:103:@767.4]
  assign _T_55085 = _T_55084[5:0]; // @[Modules.scala 150:103:@768.4]
  assign _T_55086 = $signed(_T_55085); // @[Modules.scala 150:103:@769.4]
  assign _T_55088 = $signed(-4'sh1) * $signed(io_in_340); // @[Modules.scala 150:74:@771.4]
  assign _T_55090 = $signed(-4'sh1) * $signed(io_in_341); // @[Modules.scala 151:80:@772.4]
  assign _T_55091 = $signed(_T_55088) + $signed(_T_55090); // @[Modules.scala 150:103:@773.4]
  assign _T_55092 = _T_55091[4:0]; // @[Modules.scala 150:103:@774.4]
  assign _T_55093 = $signed(_T_55092); // @[Modules.scala 150:103:@775.4]
  assign _T_55095 = $signed(-4'sh1) * $signed(io_in_342); // @[Modules.scala 150:74:@777.4]
  assign _T_55097 = $signed(-4'sh1) * $signed(io_in_343); // @[Modules.scala 151:80:@778.4]
  assign _T_55098 = $signed(_T_55095) + $signed(_T_55097); // @[Modules.scala 150:103:@779.4]
  assign _T_55099 = _T_55098[4:0]; // @[Modules.scala 150:103:@780.4]
  assign _T_55100 = $signed(_T_55099); // @[Modules.scala 150:103:@781.4]
  assign _T_55102 = $signed(-4'sh1) * $signed(io_in_344); // @[Modules.scala 150:74:@783.4]
  assign _T_55104 = $signed(-4'sh1) * $signed(io_in_345); // @[Modules.scala 151:80:@784.4]
  assign _T_55105 = $signed(_T_55102) + $signed(_T_55104); // @[Modules.scala 150:103:@785.4]
  assign _T_55106 = _T_55105[4:0]; // @[Modules.scala 150:103:@786.4]
  assign _T_55107 = $signed(_T_55106); // @[Modules.scala 150:103:@787.4]
  assign _T_55109 = $signed(-4'sh1) * $signed(io_in_346); // @[Modules.scala 150:74:@789.4]
  assign _T_55111 = $signed(-4'sh1) * $signed(io_in_347); // @[Modules.scala 151:80:@790.4]
  assign _T_55112 = $signed(_T_55109) + $signed(_T_55111); // @[Modules.scala 150:103:@791.4]
  assign _T_55113 = _T_55112[4:0]; // @[Modules.scala 150:103:@792.4]
  assign _T_55114 = $signed(_T_55113); // @[Modules.scala 150:103:@793.4]
  assign _T_55116 = $signed(-4'sh1) * $signed(io_in_348); // @[Modules.scala 150:74:@795.4]
  assign _T_55118 = $signed(-4'sh1) * $signed(io_in_349); // @[Modules.scala 151:80:@796.4]
  assign _T_55119 = $signed(_T_55116) + $signed(_T_55118); // @[Modules.scala 150:103:@797.4]
  assign _T_55120 = _T_55119[4:0]; // @[Modules.scala 150:103:@798.4]
  assign _T_55121 = $signed(_T_55120); // @[Modules.scala 150:103:@799.4]
  assign _T_55123 = $signed(4'sh1) * $signed(io_in_350); // @[Modules.scala 150:74:@801.4]
  assign _T_55125 = $signed(4'sh1) * $signed(io_in_351); // @[Modules.scala 151:80:@802.4]
  assign _T_55126 = $signed(_T_55123) + $signed(_T_55125); // @[Modules.scala 150:103:@803.4]
  assign _T_55127 = _T_55126[5:0]; // @[Modules.scala 150:103:@804.4]
  assign _T_55128 = $signed(_T_55127); // @[Modules.scala 150:103:@805.4]
  assign _T_55130 = $signed(-4'sh1) * $signed(io_in_352); // @[Modules.scala 150:74:@807.4]
  assign _T_55132 = $signed(-4'sh1) * $signed(io_in_353); // @[Modules.scala 151:80:@808.4]
  assign _T_55133 = $signed(_T_55130) + $signed(_T_55132); // @[Modules.scala 150:103:@809.4]
  assign _T_55134 = _T_55133[4:0]; // @[Modules.scala 150:103:@810.4]
  assign _T_55135 = $signed(_T_55134); // @[Modules.scala 150:103:@811.4]
  assign _T_55137 = $signed(4'sh1) * $signed(io_in_356); // @[Modules.scala 150:74:@813.4]
  assign _T_55139 = $signed(-4'sh1) * $signed(io_in_357); // @[Modules.scala 151:80:@814.4]
  assign _GEN_30 = {{1{_T_55139[4]}},_T_55139}; // @[Modules.scala 150:103:@815.4]
  assign _T_55140 = $signed(_T_55137) + $signed(_GEN_30); // @[Modules.scala 150:103:@815.4]
  assign _T_55141 = _T_55140[5:0]; // @[Modules.scala 150:103:@816.4]
  assign _T_55142 = $signed(_T_55141); // @[Modules.scala 150:103:@817.4]
  assign _T_55144 = $signed(-4'sh1) * $signed(io_in_358); // @[Modules.scala 150:74:@819.4]
  assign _T_55146 = $signed(-4'sh1) * $signed(io_in_359); // @[Modules.scala 151:80:@820.4]
  assign _T_55147 = $signed(_T_55144) + $signed(_T_55146); // @[Modules.scala 150:103:@821.4]
  assign _T_55148 = _T_55147[4:0]; // @[Modules.scala 150:103:@822.4]
  assign _T_55149 = $signed(_T_55148); // @[Modules.scala 150:103:@823.4]
  assign _T_55151 = $signed(4'sh1) * $signed(io_in_360); // @[Modules.scala 150:74:@825.4]
  assign _T_55153 = $signed(-4'sh1) * $signed(io_in_361); // @[Modules.scala 151:80:@826.4]
  assign _GEN_31 = {{1{_T_55153[4]}},_T_55153}; // @[Modules.scala 150:103:@827.4]
  assign _T_55154 = $signed(_T_55151) + $signed(_GEN_31); // @[Modules.scala 150:103:@827.4]
  assign _T_55155 = _T_55154[5:0]; // @[Modules.scala 150:103:@828.4]
  assign _T_55156 = $signed(_T_55155); // @[Modules.scala 150:103:@829.4]
  assign _T_55158 = $signed(-4'sh1) * $signed(io_in_362); // @[Modules.scala 150:74:@831.4]
  assign _T_55160 = $signed(4'sh1) * $signed(io_in_363); // @[Modules.scala 151:80:@832.4]
  assign _GEN_32 = {{1{_T_55158[4]}},_T_55158}; // @[Modules.scala 150:103:@833.4]
  assign _T_55161 = $signed(_GEN_32) + $signed(_T_55160); // @[Modules.scala 150:103:@833.4]
  assign _T_55162 = _T_55161[5:0]; // @[Modules.scala 150:103:@834.4]
  assign _T_55163 = $signed(_T_55162); // @[Modules.scala 150:103:@835.4]
  assign _T_55165 = $signed(4'sh1) * $signed(io_in_364); // @[Modules.scala 150:74:@837.4]
  assign _T_55167 = $signed(4'sh1) * $signed(io_in_365); // @[Modules.scala 151:80:@838.4]
  assign _T_55168 = $signed(_T_55165) + $signed(_T_55167); // @[Modules.scala 150:103:@839.4]
  assign _T_55169 = _T_55168[5:0]; // @[Modules.scala 150:103:@840.4]
  assign _T_55170 = $signed(_T_55169); // @[Modules.scala 150:103:@841.4]
  assign _T_55172 = $signed(4'sh1) * $signed(io_in_366); // @[Modules.scala 150:74:@843.4]
  assign _T_55174 = $signed(4'sh1) * $signed(io_in_367); // @[Modules.scala 151:80:@844.4]
  assign _T_55175 = $signed(_T_55172) + $signed(_T_55174); // @[Modules.scala 150:103:@845.4]
  assign _T_55176 = _T_55175[5:0]; // @[Modules.scala 150:103:@846.4]
  assign _T_55177 = $signed(_T_55176); // @[Modules.scala 150:103:@847.4]
  assign _T_55179 = $signed(-4'sh1) * $signed(io_in_368); // @[Modules.scala 150:74:@849.4]
  assign _T_55181 = $signed(-4'sh1) * $signed(io_in_369); // @[Modules.scala 151:80:@850.4]
  assign _T_55182 = $signed(_T_55179) + $signed(_T_55181); // @[Modules.scala 150:103:@851.4]
  assign _T_55183 = _T_55182[4:0]; // @[Modules.scala 150:103:@852.4]
  assign _T_55184 = $signed(_T_55183); // @[Modules.scala 150:103:@853.4]
  assign _T_55186 = $signed(-4'sh1) * $signed(io_in_370); // @[Modules.scala 150:74:@855.4]
  assign _T_55188 = $signed(-4'sh1) * $signed(io_in_371); // @[Modules.scala 151:80:@856.4]
  assign _T_55189 = $signed(_T_55186) + $signed(_T_55188); // @[Modules.scala 150:103:@857.4]
  assign _T_55190 = _T_55189[4:0]; // @[Modules.scala 150:103:@858.4]
  assign _T_55191 = $signed(_T_55190); // @[Modules.scala 150:103:@859.4]
  assign _T_55193 = $signed(-4'sh1) * $signed(io_in_372); // @[Modules.scala 150:74:@861.4]
  assign _T_55195 = $signed(-4'sh1) * $signed(io_in_373); // @[Modules.scala 151:80:@862.4]
  assign _T_55196 = $signed(_T_55193) + $signed(_T_55195); // @[Modules.scala 150:103:@863.4]
  assign _T_55197 = _T_55196[4:0]; // @[Modules.scala 150:103:@864.4]
  assign _T_55198 = $signed(_T_55197); // @[Modules.scala 150:103:@865.4]
  assign _T_55200 = $signed(-4'sh1) * $signed(io_in_374); // @[Modules.scala 150:74:@867.4]
  assign _T_55202 = $signed(-4'sh1) * $signed(io_in_375); // @[Modules.scala 151:80:@868.4]
  assign _T_55203 = $signed(_T_55200) + $signed(_T_55202); // @[Modules.scala 150:103:@869.4]
  assign _T_55204 = _T_55203[4:0]; // @[Modules.scala 150:103:@870.4]
  assign _T_55205 = $signed(_T_55204); // @[Modules.scala 150:103:@871.4]
  assign _T_55207 = $signed(-4'sh1) * $signed(io_in_376); // @[Modules.scala 150:74:@873.4]
  assign _T_55209 = $signed(-4'sh1) * $signed(io_in_377); // @[Modules.scala 151:80:@874.4]
  assign _T_55210 = $signed(_T_55207) + $signed(_T_55209); // @[Modules.scala 150:103:@875.4]
  assign _T_55211 = _T_55210[4:0]; // @[Modules.scala 150:103:@876.4]
  assign _T_55212 = $signed(_T_55211); // @[Modules.scala 150:103:@877.4]
  assign _T_55214 = $signed(4'sh1) * $signed(io_in_378); // @[Modules.scala 150:74:@879.4]
  assign _T_55216 = $signed(-4'sh1) * $signed(io_in_381); // @[Modules.scala 151:80:@880.4]
  assign _GEN_33 = {{1{_T_55216[4]}},_T_55216}; // @[Modules.scala 150:103:@881.4]
  assign _T_55217 = $signed(_T_55214) + $signed(_GEN_33); // @[Modules.scala 150:103:@881.4]
  assign _T_55218 = _T_55217[5:0]; // @[Modules.scala 150:103:@882.4]
  assign _T_55219 = $signed(_T_55218); // @[Modules.scala 150:103:@883.4]
  assign _T_55221 = $signed(4'sh1) * $signed(io_in_382); // @[Modules.scala 150:74:@885.4]
  assign _T_55223 = $signed(-4'sh1) * $signed(io_in_384); // @[Modules.scala 151:80:@886.4]
  assign _GEN_34 = {{1{_T_55223[4]}},_T_55223}; // @[Modules.scala 150:103:@887.4]
  assign _T_55224 = $signed(_T_55221) + $signed(_GEN_34); // @[Modules.scala 150:103:@887.4]
  assign _T_55225 = _T_55224[5:0]; // @[Modules.scala 150:103:@888.4]
  assign _T_55226 = $signed(_T_55225); // @[Modules.scala 150:103:@889.4]
  assign _T_55228 = $signed(-4'sh1) * $signed(io_in_386); // @[Modules.scala 150:74:@891.4]
  assign _T_55230 = $signed(4'sh1) * $signed(io_in_387); // @[Modules.scala 151:80:@892.4]
  assign _GEN_35 = {{1{_T_55228[4]}},_T_55228}; // @[Modules.scala 150:103:@893.4]
  assign _T_55231 = $signed(_GEN_35) + $signed(_T_55230); // @[Modules.scala 150:103:@893.4]
  assign _T_55232 = _T_55231[5:0]; // @[Modules.scala 150:103:@894.4]
  assign _T_55233 = $signed(_T_55232); // @[Modules.scala 150:103:@895.4]
  assign _T_55235 = $signed(4'sh1) * $signed(io_in_388); // @[Modules.scala 150:74:@897.4]
  assign _T_55237 = $signed(-4'sh1) * $signed(io_in_389); // @[Modules.scala 151:80:@898.4]
  assign _GEN_36 = {{1{_T_55237[4]}},_T_55237}; // @[Modules.scala 150:103:@899.4]
  assign _T_55238 = $signed(_T_55235) + $signed(_GEN_36); // @[Modules.scala 150:103:@899.4]
  assign _T_55239 = _T_55238[5:0]; // @[Modules.scala 150:103:@900.4]
  assign _T_55240 = $signed(_T_55239); // @[Modules.scala 150:103:@901.4]
  assign _T_55242 = $signed(-4'sh1) * $signed(io_in_390); // @[Modules.scala 150:74:@903.4]
  assign _T_55244 = $signed(4'sh1) * $signed(io_in_391); // @[Modules.scala 151:80:@904.4]
  assign _GEN_37 = {{1{_T_55242[4]}},_T_55242}; // @[Modules.scala 150:103:@905.4]
  assign _T_55245 = $signed(_GEN_37) + $signed(_T_55244); // @[Modules.scala 150:103:@905.4]
  assign _T_55246 = _T_55245[5:0]; // @[Modules.scala 150:103:@906.4]
  assign _T_55247 = $signed(_T_55246); // @[Modules.scala 150:103:@907.4]
  assign _T_55249 = $signed(4'sh1) * $signed(io_in_392); // @[Modules.scala 150:74:@909.4]
  assign _T_55251 = $signed(-4'sh1) * $signed(io_in_393); // @[Modules.scala 151:80:@910.4]
  assign _GEN_38 = {{1{_T_55251[4]}},_T_55251}; // @[Modules.scala 150:103:@911.4]
  assign _T_55252 = $signed(_T_55249) + $signed(_GEN_38); // @[Modules.scala 150:103:@911.4]
  assign _T_55253 = _T_55252[5:0]; // @[Modules.scala 150:103:@912.4]
  assign _T_55254 = $signed(_T_55253); // @[Modules.scala 150:103:@913.4]
  assign _T_55256 = $signed(4'sh1) * $signed(io_in_394); // @[Modules.scala 150:74:@915.4]
  assign _T_55258 = $signed(4'sh1) * $signed(io_in_395); // @[Modules.scala 151:80:@916.4]
  assign _T_55259 = $signed(_T_55256) + $signed(_T_55258); // @[Modules.scala 150:103:@917.4]
  assign _T_55260 = _T_55259[5:0]; // @[Modules.scala 150:103:@918.4]
  assign _T_55261 = $signed(_T_55260); // @[Modules.scala 150:103:@919.4]
  assign _T_55263 = $signed(-4'sh1) * $signed(io_in_396); // @[Modules.scala 150:74:@921.4]
  assign _T_55265 = $signed(-4'sh1) * $signed(io_in_397); // @[Modules.scala 151:80:@922.4]
  assign _T_55266 = $signed(_T_55263) + $signed(_T_55265); // @[Modules.scala 150:103:@923.4]
  assign _T_55267 = _T_55266[4:0]; // @[Modules.scala 150:103:@924.4]
  assign _T_55268 = $signed(_T_55267); // @[Modules.scala 150:103:@925.4]
  assign _T_55270 = $signed(-4'sh1) * $signed(io_in_398); // @[Modules.scala 150:74:@927.4]
  assign _T_55272 = $signed(-4'sh1) * $signed(io_in_399); // @[Modules.scala 151:80:@928.4]
  assign _T_55273 = $signed(_T_55270) + $signed(_T_55272); // @[Modules.scala 150:103:@929.4]
  assign _T_55274 = _T_55273[4:0]; // @[Modules.scala 150:103:@930.4]
  assign _T_55275 = $signed(_T_55274); // @[Modules.scala 150:103:@931.4]
  assign _T_55277 = $signed(-4'sh1) * $signed(io_in_400); // @[Modules.scala 150:74:@933.4]
  assign _T_55279 = $signed(-4'sh1) * $signed(io_in_401); // @[Modules.scala 151:80:@934.4]
  assign _T_55280 = $signed(_T_55277) + $signed(_T_55279); // @[Modules.scala 150:103:@935.4]
  assign _T_55281 = _T_55280[4:0]; // @[Modules.scala 150:103:@936.4]
  assign _T_55282 = $signed(_T_55281); // @[Modules.scala 150:103:@937.4]
  assign _T_55284 = $signed(-4'sh1) * $signed(io_in_402); // @[Modules.scala 150:74:@939.4]
  assign _T_55286 = $signed(-4'sh1) * $signed(io_in_403); // @[Modules.scala 151:80:@940.4]
  assign _T_55287 = $signed(_T_55284) + $signed(_T_55286); // @[Modules.scala 150:103:@941.4]
  assign _T_55288 = _T_55287[4:0]; // @[Modules.scala 150:103:@942.4]
  assign _T_55289 = $signed(_T_55288); // @[Modules.scala 150:103:@943.4]
  assign _T_55291 = $signed(-4'sh1) * $signed(io_in_404); // @[Modules.scala 150:74:@945.4]
  assign _T_55293 = $signed(4'sh1) * $signed(io_in_406); // @[Modules.scala 151:80:@946.4]
  assign _GEN_39 = {{1{_T_55291[4]}},_T_55291}; // @[Modules.scala 150:103:@947.4]
  assign _T_55294 = $signed(_GEN_39) + $signed(_T_55293); // @[Modules.scala 150:103:@947.4]
  assign _T_55295 = _T_55294[5:0]; // @[Modules.scala 150:103:@948.4]
  assign _T_55296 = $signed(_T_55295); // @[Modules.scala 150:103:@949.4]
  assign _T_55298 = $signed(4'sh1) * $signed(io_in_407); // @[Modules.scala 150:74:@951.4]
  assign _T_55300 = $signed(-4'sh1) * $signed(io_in_408); // @[Modules.scala 151:80:@952.4]
  assign _GEN_40 = {{1{_T_55300[4]}},_T_55300}; // @[Modules.scala 150:103:@953.4]
  assign _T_55301 = $signed(_T_55298) + $signed(_GEN_40); // @[Modules.scala 150:103:@953.4]
  assign _T_55302 = _T_55301[5:0]; // @[Modules.scala 150:103:@954.4]
  assign _T_55303 = $signed(_T_55302); // @[Modules.scala 150:103:@955.4]
  assign _T_55305 = $signed(-4'sh1) * $signed(io_in_409); // @[Modules.scala 150:74:@957.4]
  assign _T_55307 = $signed(4'sh1) * $signed(io_in_410); // @[Modules.scala 151:80:@958.4]
  assign _GEN_41 = {{1{_T_55305[4]}},_T_55305}; // @[Modules.scala 150:103:@959.4]
  assign _T_55308 = $signed(_GEN_41) + $signed(_T_55307); // @[Modules.scala 150:103:@959.4]
  assign _T_55309 = _T_55308[5:0]; // @[Modules.scala 150:103:@960.4]
  assign _T_55310 = $signed(_T_55309); // @[Modules.scala 150:103:@961.4]
  assign _T_55312 = $signed(4'sh1) * $signed(io_in_411); // @[Modules.scala 150:74:@963.4]
  assign _T_55314 = $signed(4'sh1) * $signed(io_in_413); // @[Modules.scala 151:80:@964.4]
  assign _T_55315 = $signed(_T_55312) + $signed(_T_55314); // @[Modules.scala 150:103:@965.4]
  assign _T_55316 = _T_55315[5:0]; // @[Modules.scala 150:103:@966.4]
  assign _T_55317 = $signed(_T_55316); // @[Modules.scala 150:103:@967.4]
  assign _T_55319 = $signed(4'sh1) * $signed(io_in_416); // @[Modules.scala 150:74:@969.4]
  assign _T_55321 = $signed(-4'sh1) * $signed(io_in_417); // @[Modules.scala 151:80:@970.4]
  assign _GEN_42 = {{1{_T_55321[4]}},_T_55321}; // @[Modules.scala 150:103:@971.4]
  assign _T_55322 = $signed(_T_55319) + $signed(_GEN_42); // @[Modules.scala 150:103:@971.4]
  assign _T_55323 = _T_55322[5:0]; // @[Modules.scala 150:103:@972.4]
  assign _T_55324 = $signed(_T_55323); // @[Modules.scala 150:103:@973.4]
  assign _T_55326 = $signed(4'sh1) * $signed(io_in_418); // @[Modules.scala 150:74:@975.4]
  assign _T_55328 = $signed(4'sh1) * $signed(io_in_420); // @[Modules.scala 151:80:@976.4]
  assign _T_55329 = $signed(_T_55326) + $signed(_T_55328); // @[Modules.scala 150:103:@977.4]
  assign _T_55330 = _T_55329[5:0]; // @[Modules.scala 150:103:@978.4]
  assign _T_55331 = $signed(_T_55330); // @[Modules.scala 150:103:@979.4]
  assign _T_55333 = $signed(-4'sh1) * $signed(io_in_421); // @[Modules.scala 150:74:@981.4]
  assign _T_55335 = $signed(4'sh1) * $signed(io_in_422); // @[Modules.scala 151:80:@982.4]
  assign _GEN_43 = {{1{_T_55333[4]}},_T_55333}; // @[Modules.scala 150:103:@983.4]
  assign _T_55336 = $signed(_GEN_43) + $signed(_T_55335); // @[Modules.scala 150:103:@983.4]
  assign _T_55337 = _T_55336[5:0]; // @[Modules.scala 150:103:@984.4]
  assign _T_55338 = $signed(_T_55337); // @[Modules.scala 150:103:@985.4]
  assign _T_55340 = $signed(4'sh1) * $signed(io_in_423); // @[Modules.scala 150:74:@987.4]
  assign _T_55342 = $signed(-4'sh1) * $signed(io_in_424); // @[Modules.scala 151:80:@988.4]
  assign _GEN_44 = {{1{_T_55342[4]}},_T_55342}; // @[Modules.scala 150:103:@989.4]
  assign _T_55343 = $signed(_T_55340) + $signed(_GEN_44); // @[Modules.scala 150:103:@989.4]
  assign _T_55344 = _T_55343[5:0]; // @[Modules.scala 150:103:@990.4]
  assign _T_55345 = $signed(_T_55344); // @[Modules.scala 150:103:@991.4]
  assign _T_55347 = $signed(-4'sh1) * $signed(io_in_425); // @[Modules.scala 150:74:@993.4]
  assign _T_55349 = $signed(-4'sh1) * $signed(io_in_426); // @[Modules.scala 151:80:@994.4]
  assign _T_55350 = $signed(_T_55347) + $signed(_T_55349); // @[Modules.scala 150:103:@995.4]
  assign _T_55351 = _T_55350[4:0]; // @[Modules.scala 150:103:@996.4]
  assign _T_55352 = $signed(_T_55351); // @[Modules.scala 150:103:@997.4]
  assign _T_55354 = $signed(-4'sh1) * $signed(io_in_427); // @[Modules.scala 150:74:@999.4]
  assign _T_55356 = $signed(-4'sh1) * $signed(io_in_429); // @[Modules.scala 151:80:@1000.4]
  assign _T_55357 = $signed(_T_55354) + $signed(_T_55356); // @[Modules.scala 150:103:@1001.4]
  assign _T_55358 = _T_55357[4:0]; // @[Modules.scala 150:103:@1002.4]
  assign _T_55359 = $signed(_T_55358); // @[Modules.scala 150:103:@1003.4]
  assign _T_55361 = $signed(-4'sh1) * $signed(io_in_430); // @[Modules.scala 150:74:@1005.4]
  assign _T_55363 = $signed(4'sh1) * $signed(io_in_432); // @[Modules.scala 151:80:@1006.4]
  assign _GEN_45 = {{1{_T_55361[4]}},_T_55361}; // @[Modules.scala 150:103:@1007.4]
  assign _T_55364 = $signed(_GEN_45) + $signed(_T_55363); // @[Modules.scala 150:103:@1007.4]
  assign _T_55365 = _T_55364[5:0]; // @[Modules.scala 150:103:@1008.4]
  assign _T_55366 = $signed(_T_55365); // @[Modules.scala 150:103:@1009.4]
  assign _T_55368 = $signed(4'sh1) * $signed(io_in_433); // @[Modules.scala 150:74:@1011.4]
  assign _T_55370 = $signed(4'sh1) * $signed(io_in_434); // @[Modules.scala 151:80:@1012.4]
  assign _T_55371 = $signed(_T_55368) + $signed(_T_55370); // @[Modules.scala 150:103:@1013.4]
  assign _T_55372 = _T_55371[5:0]; // @[Modules.scala 150:103:@1014.4]
  assign _T_55373 = $signed(_T_55372); // @[Modules.scala 150:103:@1015.4]
  assign _T_55375 = $signed(4'sh1) * $signed(io_in_435); // @[Modules.scala 150:74:@1017.4]
  assign _T_55377 = $signed(-4'sh1) * $signed(io_in_436); // @[Modules.scala 151:80:@1018.4]
  assign _GEN_46 = {{1{_T_55377[4]}},_T_55377}; // @[Modules.scala 150:103:@1019.4]
  assign _T_55378 = $signed(_T_55375) + $signed(_GEN_46); // @[Modules.scala 150:103:@1019.4]
  assign _T_55379 = _T_55378[5:0]; // @[Modules.scala 150:103:@1020.4]
  assign _T_55380 = $signed(_T_55379); // @[Modules.scala 150:103:@1021.4]
  assign _T_55382 = $signed(-4'sh1) * $signed(io_in_437); // @[Modules.scala 150:74:@1023.4]
  assign _T_55384 = $signed(4'sh1) * $signed(io_in_438); // @[Modules.scala 151:80:@1024.4]
  assign _GEN_47 = {{1{_T_55382[4]}},_T_55382}; // @[Modules.scala 150:103:@1025.4]
  assign _T_55385 = $signed(_GEN_47) + $signed(_T_55384); // @[Modules.scala 150:103:@1025.4]
  assign _T_55386 = _T_55385[5:0]; // @[Modules.scala 150:103:@1026.4]
  assign _T_55387 = $signed(_T_55386); // @[Modules.scala 150:103:@1027.4]
  assign _T_55389 = $signed(4'sh1) * $signed(io_in_439); // @[Modules.scala 150:74:@1029.4]
  assign _T_55391 = $signed(4'sh1) * $signed(io_in_440); // @[Modules.scala 151:80:@1030.4]
  assign _T_55392 = $signed(_T_55389) + $signed(_T_55391); // @[Modules.scala 150:103:@1031.4]
  assign _T_55393 = _T_55392[5:0]; // @[Modules.scala 150:103:@1032.4]
  assign _T_55394 = $signed(_T_55393); // @[Modules.scala 150:103:@1033.4]
  assign _T_55396 = $signed(4'sh1) * $signed(io_in_441); // @[Modules.scala 150:74:@1035.4]
  assign _T_55398 = $signed(-4'sh1) * $signed(io_in_442); // @[Modules.scala 151:80:@1036.4]
  assign _GEN_48 = {{1{_T_55398[4]}},_T_55398}; // @[Modules.scala 150:103:@1037.4]
  assign _T_55399 = $signed(_T_55396) + $signed(_GEN_48); // @[Modules.scala 150:103:@1037.4]
  assign _T_55400 = _T_55399[5:0]; // @[Modules.scala 150:103:@1038.4]
  assign _T_55401 = $signed(_T_55400); // @[Modules.scala 150:103:@1039.4]
  assign _T_55403 = $signed(-4'sh1) * $signed(io_in_443); // @[Modules.scala 150:74:@1041.4]
  assign _T_55405 = $signed(4'sh1) * $signed(io_in_445); // @[Modules.scala 151:80:@1042.4]
  assign _GEN_49 = {{1{_T_55403[4]}},_T_55403}; // @[Modules.scala 150:103:@1043.4]
  assign _T_55406 = $signed(_GEN_49) + $signed(_T_55405); // @[Modules.scala 150:103:@1043.4]
  assign _T_55407 = _T_55406[5:0]; // @[Modules.scala 150:103:@1044.4]
  assign _T_55408 = $signed(_T_55407); // @[Modules.scala 150:103:@1045.4]
  assign _T_55410 = $signed(4'sh1) * $signed(io_in_446); // @[Modules.scala 150:74:@1047.4]
  assign _T_55412 = $signed(4'sh1) * $signed(io_in_447); // @[Modules.scala 151:80:@1048.4]
  assign _T_55413 = $signed(_T_55410) + $signed(_T_55412); // @[Modules.scala 150:103:@1049.4]
  assign _T_55414 = _T_55413[5:0]; // @[Modules.scala 150:103:@1050.4]
  assign _T_55415 = $signed(_T_55414); // @[Modules.scala 150:103:@1051.4]
  assign _T_55417 = $signed(-4'sh1) * $signed(io_in_448); // @[Modules.scala 150:74:@1053.4]
  assign _T_55419 = $signed(-4'sh1) * $signed(io_in_449); // @[Modules.scala 151:80:@1054.4]
  assign _T_55420 = $signed(_T_55417) + $signed(_T_55419); // @[Modules.scala 150:103:@1055.4]
  assign _T_55421 = _T_55420[4:0]; // @[Modules.scala 150:103:@1056.4]
  assign _T_55422 = $signed(_T_55421); // @[Modules.scala 150:103:@1057.4]
  assign _T_55424 = $signed(4'sh1) * $signed(io_in_450); // @[Modules.scala 150:74:@1059.4]
  assign _T_55426 = $signed(4'sh1) * $signed(io_in_451); // @[Modules.scala 151:80:@1060.4]
  assign _T_55427 = $signed(_T_55424) + $signed(_T_55426); // @[Modules.scala 150:103:@1061.4]
  assign _T_55428 = _T_55427[5:0]; // @[Modules.scala 150:103:@1062.4]
  assign _T_55429 = $signed(_T_55428); // @[Modules.scala 150:103:@1063.4]
  assign _T_55431 = $signed(-4'sh1) * $signed(io_in_452); // @[Modules.scala 150:74:@1065.4]
  assign _T_55433 = $signed(-4'sh1) * $signed(io_in_453); // @[Modules.scala 151:80:@1066.4]
  assign _T_55434 = $signed(_T_55431) + $signed(_T_55433); // @[Modules.scala 150:103:@1067.4]
  assign _T_55435 = _T_55434[4:0]; // @[Modules.scala 150:103:@1068.4]
  assign _T_55436 = $signed(_T_55435); // @[Modules.scala 150:103:@1069.4]
  assign _T_55438 = $signed(4'sh1) * $signed(io_in_455); // @[Modules.scala 150:74:@1071.4]
  assign _T_55440 = $signed(4'sh1) * $signed(io_in_457); // @[Modules.scala 151:80:@1072.4]
  assign _T_55441 = $signed(_T_55438) + $signed(_T_55440); // @[Modules.scala 150:103:@1073.4]
  assign _T_55442 = _T_55441[5:0]; // @[Modules.scala 150:103:@1074.4]
  assign _T_55443 = $signed(_T_55442); // @[Modules.scala 150:103:@1075.4]
  assign _T_55445 = $signed(4'sh1) * $signed(io_in_458); // @[Modules.scala 150:74:@1077.4]
  assign _T_55447 = $signed(4'sh1) * $signed(io_in_459); // @[Modules.scala 151:80:@1078.4]
  assign _T_55448 = $signed(_T_55445) + $signed(_T_55447); // @[Modules.scala 150:103:@1079.4]
  assign _T_55449 = _T_55448[5:0]; // @[Modules.scala 150:103:@1080.4]
  assign _T_55450 = $signed(_T_55449); // @[Modules.scala 150:103:@1081.4]
  assign _T_55452 = $signed(4'sh1) * $signed(io_in_461); // @[Modules.scala 150:74:@1083.4]
  assign _T_55454 = $signed(4'sh1) * $signed(io_in_462); // @[Modules.scala 151:80:@1084.4]
  assign _T_55455 = $signed(_T_55452) + $signed(_T_55454); // @[Modules.scala 150:103:@1085.4]
  assign _T_55456 = _T_55455[5:0]; // @[Modules.scala 150:103:@1086.4]
  assign _T_55457 = $signed(_T_55456); // @[Modules.scala 150:103:@1087.4]
  assign _T_55459 = $signed(4'sh1) * $signed(io_in_463); // @[Modules.scala 150:74:@1089.4]
  assign _T_55461 = $signed(-4'sh1) * $signed(io_in_465); // @[Modules.scala 151:80:@1090.4]
  assign _GEN_50 = {{1{_T_55461[4]}},_T_55461}; // @[Modules.scala 150:103:@1091.4]
  assign _T_55462 = $signed(_T_55459) + $signed(_GEN_50); // @[Modules.scala 150:103:@1091.4]
  assign _T_55463 = _T_55462[5:0]; // @[Modules.scala 150:103:@1092.4]
  assign _T_55464 = $signed(_T_55463); // @[Modules.scala 150:103:@1093.4]
  assign _T_55466 = $signed(-4'sh1) * $signed(io_in_466); // @[Modules.scala 150:74:@1095.4]
  assign _T_55468 = $signed(4'sh1) * $signed(io_in_467); // @[Modules.scala 151:80:@1096.4]
  assign _GEN_51 = {{1{_T_55466[4]}},_T_55466}; // @[Modules.scala 150:103:@1097.4]
  assign _T_55469 = $signed(_GEN_51) + $signed(_T_55468); // @[Modules.scala 150:103:@1097.4]
  assign _T_55470 = _T_55469[5:0]; // @[Modules.scala 150:103:@1098.4]
  assign _T_55471 = $signed(_T_55470); // @[Modules.scala 150:103:@1099.4]
  assign _T_55473 = $signed(4'sh1) * $signed(io_in_469); // @[Modules.scala 150:74:@1101.4]
  assign _T_55475 = $signed(-4'sh1) * $signed(io_in_471); // @[Modules.scala 151:80:@1102.4]
  assign _GEN_52 = {{1{_T_55475[4]}},_T_55475}; // @[Modules.scala 150:103:@1103.4]
  assign _T_55476 = $signed(_T_55473) + $signed(_GEN_52); // @[Modules.scala 150:103:@1103.4]
  assign _T_55477 = _T_55476[5:0]; // @[Modules.scala 150:103:@1104.4]
  assign _T_55478 = $signed(_T_55477); // @[Modules.scala 150:103:@1105.4]
  assign _T_55480 = $signed(4'sh1) * $signed(io_in_473); // @[Modules.scala 150:74:@1107.4]
  assign _T_55482 = $signed(4'sh1) * $signed(io_in_474); // @[Modules.scala 151:80:@1108.4]
  assign _T_55483 = $signed(_T_55480) + $signed(_T_55482); // @[Modules.scala 150:103:@1109.4]
  assign _T_55484 = _T_55483[5:0]; // @[Modules.scala 150:103:@1110.4]
  assign _T_55485 = $signed(_T_55484); // @[Modules.scala 150:103:@1111.4]
  assign _T_55487 = $signed(-4'sh1) * $signed(io_in_477); // @[Modules.scala 150:74:@1113.4]
  assign _T_55489 = $signed(4'sh1) * $signed(io_in_478); // @[Modules.scala 151:80:@1114.4]
  assign _GEN_53 = {{1{_T_55487[4]}},_T_55487}; // @[Modules.scala 150:103:@1115.4]
  assign _T_55490 = $signed(_GEN_53) + $signed(_T_55489); // @[Modules.scala 150:103:@1115.4]
  assign _T_55491 = _T_55490[5:0]; // @[Modules.scala 150:103:@1116.4]
  assign _T_55492 = $signed(_T_55491); // @[Modules.scala 150:103:@1117.4]
  assign _T_55494 = $signed(4'sh1) * $signed(io_in_479); // @[Modules.scala 150:74:@1119.4]
  assign _T_55496 = $signed(4'sh1) * $signed(io_in_480); // @[Modules.scala 151:80:@1120.4]
  assign _T_55497 = $signed(_T_55494) + $signed(_T_55496); // @[Modules.scala 150:103:@1121.4]
  assign _T_55498 = _T_55497[5:0]; // @[Modules.scala 150:103:@1122.4]
  assign _T_55499 = $signed(_T_55498); // @[Modules.scala 150:103:@1123.4]
  assign _T_55501 = $signed(4'sh1) * $signed(io_in_482); // @[Modules.scala 150:74:@1125.4]
  assign _T_55503 = $signed(-4'sh1) * $signed(io_in_485); // @[Modules.scala 151:80:@1126.4]
  assign _GEN_54 = {{1{_T_55503[4]}},_T_55503}; // @[Modules.scala 150:103:@1127.4]
  assign _T_55504 = $signed(_T_55501) + $signed(_GEN_54); // @[Modules.scala 150:103:@1127.4]
  assign _T_55505 = _T_55504[5:0]; // @[Modules.scala 150:103:@1128.4]
  assign _T_55506 = $signed(_T_55505); // @[Modules.scala 150:103:@1129.4]
  assign _T_55508 = $signed(4'sh1) * $signed(io_in_486); // @[Modules.scala 150:74:@1131.4]
  assign _T_55510 = $signed(4'sh1) * $signed(io_in_487); // @[Modules.scala 151:80:@1132.4]
  assign _T_55511 = $signed(_T_55508) + $signed(_T_55510); // @[Modules.scala 150:103:@1133.4]
  assign _T_55512 = _T_55511[5:0]; // @[Modules.scala 150:103:@1134.4]
  assign _T_55513 = $signed(_T_55512); // @[Modules.scala 150:103:@1135.4]
  assign _T_55515 = $signed(4'sh1) * $signed(io_in_488); // @[Modules.scala 150:74:@1137.4]
  assign _T_55517 = $signed(4'sh1) * $signed(io_in_489); // @[Modules.scala 151:80:@1138.4]
  assign _T_55518 = $signed(_T_55515) + $signed(_T_55517); // @[Modules.scala 150:103:@1139.4]
  assign _T_55519 = _T_55518[5:0]; // @[Modules.scala 150:103:@1140.4]
  assign _T_55520 = $signed(_T_55519); // @[Modules.scala 150:103:@1141.4]
  assign _T_55522 = $signed(4'sh1) * $signed(io_in_490); // @[Modules.scala 150:74:@1143.4]
  assign _T_55524 = $signed(4'sh1) * $signed(io_in_491); // @[Modules.scala 151:80:@1144.4]
  assign _T_55525 = $signed(_T_55522) + $signed(_T_55524); // @[Modules.scala 150:103:@1145.4]
  assign _T_55526 = _T_55525[5:0]; // @[Modules.scala 150:103:@1146.4]
  assign _T_55527 = $signed(_T_55526); // @[Modules.scala 150:103:@1147.4]
  assign _T_55529 = $signed(-4'sh1) * $signed(io_in_492); // @[Modules.scala 150:74:@1149.4]
  assign _T_55531 = $signed(-4'sh1) * $signed(io_in_493); // @[Modules.scala 151:80:@1150.4]
  assign _T_55532 = $signed(_T_55529) + $signed(_T_55531); // @[Modules.scala 150:103:@1151.4]
  assign _T_55533 = _T_55532[4:0]; // @[Modules.scala 150:103:@1152.4]
  assign _T_55534 = $signed(_T_55533); // @[Modules.scala 150:103:@1153.4]
  assign _T_55536 = $signed(-4'sh1) * $signed(io_in_494); // @[Modules.scala 150:74:@1155.4]
  assign _T_55538 = $signed(4'sh1) * $signed(io_in_497); // @[Modules.scala 151:80:@1156.4]
  assign _GEN_55 = {{1{_T_55536[4]}},_T_55536}; // @[Modules.scala 150:103:@1157.4]
  assign _T_55539 = $signed(_GEN_55) + $signed(_T_55538); // @[Modules.scala 150:103:@1157.4]
  assign _T_55540 = _T_55539[5:0]; // @[Modules.scala 150:103:@1158.4]
  assign _T_55541 = $signed(_T_55540); // @[Modules.scala 150:103:@1159.4]
  assign _T_55543 = $signed(4'sh1) * $signed(io_in_499); // @[Modules.scala 150:74:@1161.4]
  assign _T_55545 = $signed(4'sh1) * $signed(io_in_500); // @[Modules.scala 151:80:@1162.4]
  assign _T_55546 = $signed(_T_55543) + $signed(_T_55545); // @[Modules.scala 150:103:@1163.4]
  assign _T_55547 = _T_55546[5:0]; // @[Modules.scala 150:103:@1164.4]
  assign _T_55548 = $signed(_T_55547); // @[Modules.scala 150:103:@1165.4]
  assign _T_55550 = $signed(4'sh1) * $signed(io_in_501); // @[Modules.scala 150:74:@1167.4]
  assign _T_55552 = $signed(4'sh1) * $signed(io_in_502); // @[Modules.scala 151:80:@1168.4]
  assign _T_55553 = $signed(_T_55550) + $signed(_T_55552); // @[Modules.scala 150:103:@1169.4]
  assign _T_55554 = _T_55553[5:0]; // @[Modules.scala 150:103:@1170.4]
  assign _T_55555 = $signed(_T_55554); // @[Modules.scala 150:103:@1171.4]
  assign _T_55557 = $signed(4'sh1) * $signed(io_in_503); // @[Modules.scala 150:74:@1173.4]
  assign _T_55559 = $signed(-4'sh1) * $signed(io_in_504); // @[Modules.scala 151:80:@1174.4]
  assign _GEN_56 = {{1{_T_55559[4]}},_T_55559}; // @[Modules.scala 150:103:@1175.4]
  assign _T_55560 = $signed(_T_55557) + $signed(_GEN_56); // @[Modules.scala 150:103:@1175.4]
  assign _T_55561 = _T_55560[5:0]; // @[Modules.scala 150:103:@1176.4]
  assign _T_55562 = $signed(_T_55561); // @[Modules.scala 150:103:@1177.4]
  assign _T_55564 = $signed(4'sh1) * $signed(io_in_505); // @[Modules.scala 150:74:@1179.4]
  assign _T_55566 = $signed(4'sh1) * $signed(io_in_506); // @[Modules.scala 151:80:@1180.4]
  assign _T_55567 = $signed(_T_55564) + $signed(_T_55566); // @[Modules.scala 150:103:@1181.4]
  assign _T_55568 = _T_55567[5:0]; // @[Modules.scala 150:103:@1182.4]
  assign _T_55569 = $signed(_T_55568); // @[Modules.scala 150:103:@1183.4]
  assign _T_55571 = $signed(4'sh1) * $signed(io_in_507); // @[Modules.scala 150:74:@1185.4]
  assign _T_55573 = $signed(4'sh1) * $signed(io_in_508); // @[Modules.scala 151:80:@1186.4]
  assign _T_55574 = $signed(_T_55571) + $signed(_T_55573); // @[Modules.scala 150:103:@1187.4]
  assign _T_55575 = _T_55574[5:0]; // @[Modules.scala 150:103:@1188.4]
  assign _T_55576 = $signed(_T_55575); // @[Modules.scala 150:103:@1189.4]
  assign _T_55578 = $signed(4'sh1) * $signed(io_in_509); // @[Modules.scala 150:74:@1191.4]
  assign _T_55580 = $signed(-4'sh1) * $signed(io_in_510); // @[Modules.scala 151:80:@1192.4]
  assign _GEN_57 = {{1{_T_55580[4]}},_T_55580}; // @[Modules.scala 150:103:@1193.4]
  assign _T_55581 = $signed(_T_55578) + $signed(_GEN_57); // @[Modules.scala 150:103:@1193.4]
  assign _T_55582 = _T_55581[5:0]; // @[Modules.scala 150:103:@1194.4]
  assign _T_55583 = $signed(_T_55582); // @[Modules.scala 150:103:@1195.4]
  assign _T_55585 = $signed(-4'sh1) * $signed(io_in_512); // @[Modules.scala 150:74:@1197.4]
  assign _T_55587 = $signed(4'sh1) * $signed(io_in_513); // @[Modules.scala 151:80:@1198.4]
  assign _GEN_58 = {{1{_T_55585[4]}},_T_55585}; // @[Modules.scala 150:103:@1199.4]
  assign _T_55588 = $signed(_GEN_58) + $signed(_T_55587); // @[Modules.scala 150:103:@1199.4]
  assign _T_55589 = _T_55588[5:0]; // @[Modules.scala 150:103:@1200.4]
  assign _T_55590 = $signed(_T_55589); // @[Modules.scala 150:103:@1201.4]
  assign _T_55592 = $signed(4'sh1) * $signed(io_in_514); // @[Modules.scala 150:74:@1203.4]
  assign _T_55594 = $signed(4'sh1) * $signed(io_in_515); // @[Modules.scala 151:80:@1204.4]
  assign _T_55595 = $signed(_T_55592) + $signed(_T_55594); // @[Modules.scala 150:103:@1205.4]
  assign _T_55596 = _T_55595[5:0]; // @[Modules.scala 150:103:@1206.4]
  assign _T_55597 = $signed(_T_55596); // @[Modules.scala 150:103:@1207.4]
  assign _T_55599 = $signed(4'sh1) * $signed(io_in_516); // @[Modules.scala 150:74:@1209.4]
  assign _T_55601 = $signed(4'sh1) * $signed(io_in_517); // @[Modules.scala 151:80:@1210.4]
  assign _T_55602 = $signed(_T_55599) + $signed(_T_55601); // @[Modules.scala 150:103:@1211.4]
  assign _T_55603 = _T_55602[5:0]; // @[Modules.scala 150:103:@1212.4]
  assign _T_55604 = $signed(_T_55603); // @[Modules.scala 150:103:@1213.4]
  assign _T_55606 = $signed(4'sh1) * $signed(io_in_518); // @[Modules.scala 150:74:@1215.4]
  assign _T_55608 = $signed(-4'sh1) * $signed(io_in_519); // @[Modules.scala 151:80:@1216.4]
  assign _GEN_59 = {{1{_T_55608[4]}},_T_55608}; // @[Modules.scala 150:103:@1217.4]
  assign _T_55609 = $signed(_T_55606) + $signed(_GEN_59); // @[Modules.scala 150:103:@1217.4]
  assign _T_55610 = _T_55609[5:0]; // @[Modules.scala 150:103:@1218.4]
  assign _T_55611 = $signed(_T_55610); // @[Modules.scala 150:103:@1219.4]
  assign _T_55613 = $signed(-4'sh1) * $signed(io_in_520); // @[Modules.scala 150:74:@1221.4]
  assign _T_55615 = $signed(4'sh1) * $signed(io_in_521); // @[Modules.scala 151:80:@1222.4]
  assign _GEN_60 = {{1{_T_55613[4]}},_T_55613}; // @[Modules.scala 150:103:@1223.4]
  assign _T_55616 = $signed(_GEN_60) + $signed(_T_55615); // @[Modules.scala 150:103:@1223.4]
  assign _T_55617 = _T_55616[5:0]; // @[Modules.scala 150:103:@1224.4]
  assign _T_55618 = $signed(_T_55617); // @[Modules.scala 150:103:@1225.4]
  assign _T_55620 = $signed(4'sh1) * $signed(io_in_523); // @[Modules.scala 150:74:@1227.4]
  assign _T_55622 = $signed(4'sh1) * $signed(io_in_524); // @[Modules.scala 151:80:@1228.4]
  assign _T_55623 = $signed(_T_55620) + $signed(_T_55622); // @[Modules.scala 150:103:@1229.4]
  assign _T_55624 = _T_55623[5:0]; // @[Modules.scala 150:103:@1230.4]
  assign _T_55625 = $signed(_T_55624); // @[Modules.scala 150:103:@1231.4]
  assign _T_55627 = $signed(4'sh1) * $signed(io_in_526); // @[Modules.scala 150:74:@1233.4]
  assign _T_55629 = $signed(4'sh1) * $signed(io_in_527); // @[Modules.scala 151:80:@1234.4]
  assign _T_55630 = $signed(_T_55627) + $signed(_T_55629); // @[Modules.scala 150:103:@1235.4]
  assign _T_55631 = _T_55630[5:0]; // @[Modules.scala 150:103:@1236.4]
  assign _T_55632 = $signed(_T_55631); // @[Modules.scala 150:103:@1237.4]
  assign _T_55634 = $signed(4'sh1) * $signed(io_in_528); // @[Modules.scala 150:74:@1239.4]
  assign _T_55636 = $signed(4'sh1) * $signed(io_in_529); // @[Modules.scala 151:80:@1240.4]
  assign _T_55637 = $signed(_T_55634) + $signed(_T_55636); // @[Modules.scala 150:103:@1241.4]
  assign _T_55638 = _T_55637[5:0]; // @[Modules.scala 150:103:@1242.4]
  assign _T_55639 = $signed(_T_55638); // @[Modules.scala 150:103:@1243.4]
  assign _T_55641 = $signed(4'sh1) * $signed(io_in_530); // @[Modules.scala 150:74:@1245.4]
  assign _T_55643 = $signed(4'sh1) * $signed(io_in_531); // @[Modules.scala 151:80:@1246.4]
  assign _T_55644 = $signed(_T_55641) + $signed(_T_55643); // @[Modules.scala 150:103:@1247.4]
  assign _T_55645 = _T_55644[5:0]; // @[Modules.scala 150:103:@1248.4]
  assign _T_55646 = $signed(_T_55645); // @[Modules.scala 150:103:@1249.4]
  assign _T_55648 = $signed(-4'sh1) * $signed(io_in_532); // @[Modules.scala 150:74:@1251.4]
  assign _T_55650 = $signed(4'sh1) * $signed(io_in_533); // @[Modules.scala 151:80:@1252.4]
  assign _GEN_61 = {{1{_T_55648[4]}},_T_55648}; // @[Modules.scala 150:103:@1253.4]
  assign _T_55651 = $signed(_GEN_61) + $signed(_T_55650); // @[Modules.scala 150:103:@1253.4]
  assign _T_55652 = _T_55651[5:0]; // @[Modules.scala 150:103:@1254.4]
  assign _T_55653 = $signed(_T_55652); // @[Modules.scala 150:103:@1255.4]
  assign _T_55655 = $signed(4'sh1) * $signed(io_in_534); // @[Modules.scala 150:74:@1257.4]
  assign _T_55657 = $signed(4'sh1) * $signed(io_in_535); // @[Modules.scala 151:80:@1258.4]
  assign _T_55658 = $signed(_T_55655) + $signed(_T_55657); // @[Modules.scala 150:103:@1259.4]
  assign _T_55659 = _T_55658[5:0]; // @[Modules.scala 150:103:@1260.4]
  assign _T_55660 = $signed(_T_55659); // @[Modules.scala 150:103:@1261.4]
  assign _T_55662 = $signed(4'sh1) * $signed(io_in_536); // @[Modules.scala 150:74:@1263.4]
  assign _T_55664 = $signed(4'sh1) * $signed(io_in_537); // @[Modules.scala 151:80:@1264.4]
  assign _T_55665 = $signed(_T_55662) + $signed(_T_55664); // @[Modules.scala 150:103:@1265.4]
  assign _T_55666 = _T_55665[5:0]; // @[Modules.scala 150:103:@1266.4]
  assign _T_55667 = $signed(_T_55666); // @[Modules.scala 150:103:@1267.4]
  assign _T_55669 = $signed(4'sh1) * $signed(io_in_539); // @[Modules.scala 150:74:@1269.4]
  assign _T_55671 = $signed(4'sh1) * $signed(io_in_540); // @[Modules.scala 151:80:@1270.4]
  assign _T_55672 = $signed(_T_55669) + $signed(_T_55671); // @[Modules.scala 150:103:@1271.4]
  assign _T_55673 = _T_55672[5:0]; // @[Modules.scala 150:103:@1272.4]
  assign _T_55674 = $signed(_T_55673); // @[Modules.scala 150:103:@1273.4]
  assign _T_55676 = $signed(4'sh1) * $signed(io_in_541); // @[Modules.scala 150:74:@1275.4]
  assign _T_55678 = $signed(4'sh1) * $signed(io_in_542); // @[Modules.scala 151:80:@1276.4]
  assign _T_55679 = $signed(_T_55676) + $signed(_T_55678); // @[Modules.scala 150:103:@1277.4]
  assign _T_55680 = _T_55679[5:0]; // @[Modules.scala 150:103:@1278.4]
  assign _T_55681 = $signed(_T_55680); // @[Modules.scala 150:103:@1279.4]
  assign _T_55683 = $signed(4'sh1) * $signed(io_in_543); // @[Modules.scala 150:74:@1281.4]
  assign _T_55685 = $signed(4'sh1) * $signed(io_in_544); // @[Modules.scala 151:80:@1282.4]
  assign _T_55686 = $signed(_T_55683) + $signed(_T_55685); // @[Modules.scala 150:103:@1283.4]
  assign _T_55687 = _T_55686[5:0]; // @[Modules.scala 150:103:@1284.4]
  assign _T_55688 = $signed(_T_55687); // @[Modules.scala 150:103:@1285.4]
  assign _T_55690 = $signed(4'sh1) * $signed(io_in_545); // @[Modules.scala 150:74:@1287.4]
  assign _T_55692 = $signed(4'sh1) * $signed(io_in_546); // @[Modules.scala 151:80:@1288.4]
  assign _T_55693 = $signed(_T_55690) + $signed(_T_55692); // @[Modules.scala 150:103:@1289.4]
  assign _T_55694 = _T_55693[5:0]; // @[Modules.scala 150:103:@1290.4]
  assign _T_55695 = $signed(_T_55694); // @[Modules.scala 150:103:@1291.4]
  assign _T_55697 = $signed(4'sh1) * $signed(io_in_547); // @[Modules.scala 150:74:@1293.4]
  assign _T_55699 = $signed(4'sh1) * $signed(io_in_548); // @[Modules.scala 151:80:@1294.4]
  assign _T_55700 = $signed(_T_55697) + $signed(_T_55699); // @[Modules.scala 150:103:@1295.4]
  assign _T_55701 = _T_55700[5:0]; // @[Modules.scala 150:103:@1296.4]
  assign _T_55702 = $signed(_T_55701); // @[Modules.scala 150:103:@1297.4]
  assign _T_55704 = $signed(4'sh1) * $signed(io_in_549); // @[Modules.scala 150:74:@1299.4]
  assign _T_55706 = $signed(4'sh1) * $signed(io_in_551); // @[Modules.scala 151:80:@1300.4]
  assign _T_55707 = $signed(_T_55704) + $signed(_T_55706); // @[Modules.scala 150:103:@1301.4]
  assign _T_55708 = _T_55707[5:0]; // @[Modules.scala 150:103:@1302.4]
  assign _T_55709 = $signed(_T_55708); // @[Modules.scala 150:103:@1303.4]
  assign _T_55711 = $signed(4'sh1) * $signed(io_in_552); // @[Modules.scala 150:74:@1305.4]
  assign _T_55713 = $signed(4'sh1) * $signed(io_in_556); // @[Modules.scala 151:80:@1306.4]
  assign _T_55714 = $signed(_T_55711) + $signed(_T_55713); // @[Modules.scala 150:103:@1307.4]
  assign _T_55715 = _T_55714[5:0]; // @[Modules.scala 150:103:@1308.4]
  assign _T_55716 = $signed(_T_55715); // @[Modules.scala 150:103:@1309.4]
  assign _T_55718 = $signed(4'sh1) * $signed(io_in_557); // @[Modules.scala 150:74:@1311.4]
  assign _T_55720 = $signed(4'sh1) * $signed(io_in_558); // @[Modules.scala 151:80:@1312.4]
  assign _T_55721 = $signed(_T_55718) + $signed(_T_55720); // @[Modules.scala 150:103:@1313.4]
  assign _T_55722 = _T_55721[5:0]; // @[Modules.scala 150:103:@1314.4]
  assign _T_55723 = $signed(_T_55722); // @[Modules.scala 150:103:@1315.4]
  assign _T_55725 = $signed(-4'sh1) * $signed(io_in_559); // @[Modules.scala 150:74:@1317.4]
  assign _T_55727 = $signed(4'sh1) * $signed(io_in_562); // @[Modules.scala 151:80:@1318.4]
  assign _GEN_62 = {{1{_T_55725[4]}},_T_55725}; // @[Modules.scala 150:103:@1319.4]
  assign _T_55728 = $signed(_GEN_62) + $signed(_T_55727); // @[Modules.scala 150:103:@1319.4]
  assign _T_55729 = _T_55728[5:0]; // @[Modules.scala 150:103:@1320.4]
  assign _T_55730 = $signed(_T_55729); // @[Modules.scala 150:103:@1321.4]
  assign _T_55732 = $signed(4'sh1) * $signed(io_in_563); // @[Modules.scala 150:74:@1323.4]
  assign _T_55734 = $signed(4'sh1) * $signed(io_in_564); // @[Modules.scala 151:80:@1324.4]
  assign _T_55735 = $signed(_T_55732) + $signed(_T_55734); // @[Modules.scala 150:103:@1325.4]
  assign _T_55736 = _T_55735[5:0]; // @[Modules.scala 150:103:@1326.4]
  assign _T_55737 = $signed(_T_55736); // @[Modules.scala 150:103:@1327.4]
  assign _T_55739 = $signed(4'sh1) * $signed(io_in_565); // @[Modules.scala 150:74:@1329.4]
  assign _T_55741 = $signed(4'sh1) * $signed(io_in_566); // @[Modules.scala 151:80:@1330.4]
  assign _T_55742 = $signed(_T_55739) + $signed(_T_55741); // @[Modules.scala 150:103:@1331.4]
  assign _T_55743 = _T_55742[5:0]; // @[Modules.scala 150:103:@1332.4]
  assign _T_55744 = $signed(_T_55743); // @[Modules.scala 150:103:@1333.4]
  assign _T_55746 = $signed(4'sh1) * $signed(io_in_567); // @[Modules.scala 150:74:@1335.4]
  assign _T_55748 = $signed(4'sh1) * $signed(io_in_570); // @[Modules.scala 151:80:@1336.4]
  assign _T_55749 = $signed(_T_55746) + $signed(_T_55748); // @[Modules.scala 150:103:@1337.4]
  assign _T_55750 = _T_55749[5:0]; // @[Modules.scala 150:103:@1338.4]
  assign _T_55751 = $signed(_T_55750); // @[Modules.scala 150:103:@1339.4]
  assign _T_55753 = $signed(4'sh1) * $signed(io_in_571); // @[Modules.scala 150:74:@1341.4]
  assign _T_55755 = $signed(4'sh1) * $signed(io_in_572); // @[Modules.scala 151:80:@1342.4]
  assign _T_55756 = $signed(_T_55753) + $signed(_T_55755); // @[Modules.scala 150:103:@1343.4]
  assign _T_55757 = _T_55756[5:0]; // @[Modules.scala 150:103:@1344.4]
  assign _T_55758 = $signed(_T_55757); // @[Modules.scala 150:103:@1345.4]
  assign _T_55760 = $signed(4'sh1) * $signed(io_in_573); // @[Modules.scala 150:74:@1347.4]
  assign _T_55762 = $signed(4'sh1) * $signed(io_in_574); // @[Modules.scala 151:80:@1348.4]
  assign _T_55763 = $signed(_T_55760) + $signed(_T_55762); // @[Modules.scala 150:103:@1349.4]
  assign _T_55764 = _T_55763[5:0]; // @[Modules.scala 150:103:@1350.4]
  assign _T_55765 = $signed(_T_55764); // @[Modules.scala 150:103:@1351.4]
  assign _T_55767 = $signed(4'sh1) * $signed(io_in_578); // @[Modules.scala 150:74:@1353.4]
  assign _T_55769 = $signed(-4'sh1) * $signed(io_in_580); // @[Modules.scala 151:80:@1354.4]
  assign _GEN_63 = {{1{_T_55769[4]}},_T_55769}; // @[Modules.scala 150:103:@1355.4]
  assign _T_55770 = $signed(_T_55767) + $signed(_GEN_63); // @[Modules.scala 150:103:@1355.4]
  assign _T_55771 = _T_55770[5:0]; // @[Modules.scala 150:103:@1356.4]
  assign _T_55772 = $signed(_T_55771); // @[Modules.scala 150:103:@1357.4]
  assign _T_55774 = $signed(-4'sh1) * $signed(io_in_582); // @[Modules.scala 150:74:@1359.4]
  assign _T_55776 = $signed(4'sh1) * $signed(io_in_583); // @[Modules.scala 151:80:@1360.4]
  assign _GEN_64 = {{1{_T_55774[4]}},_T_55774}; // @[Modules.scala 150:103:@1361.4]
  assign _T_55777 = $signed(_GEN_64) + $signed(_T_55776); // @[Modules.scala 150:103:@1361.4]
  assign _T_55778 = _T_55777[5:0]; // @[Modules.scala 150:103:@1362.4]
  assign _T_55779 = $signed(_T_55778); // @[Modules.scala 150:103:@1363.4]
  assign _T_55781 = $signed(4'sh1) * $signed(io_in_584); // @[Modules.scala 150:74:@1365.4]
  assign _T_55783 = $signed(4'sh1) * $signed(io_in_585); // @[Modules.scala 151:80:@1366.4]
  assign _T_55784 = $signed(_T_55781) + $signed(_T_55783); // @[Modules.scala 150:103:@1367.4]
  assign _T_55785 = _T_55784[5:0]; // @[Modules.scala 150:103:@1368.4]
  assign _T_55786 = $signed(_T_55785); // @[Modules.scala 150:103:@1369.4]
  assign _T_55788 = $signed(4'sh1) * $signed(io_in_587); // @[Modules.scala 150:74:@1371.4]
  assign _T_55790 = $signed(4'sh1) * $signed(io_in_588); // @[Modules.scala 151:80:@1372.4]
  assign _T_55791 = $signed(_T_55788) + $signed(_T_55790); // @[Modules.scala 150:103:@1373.4]
  assign _T_55792 = _T_55791[5:0]; // @[Modules.scala 150:103:@1374.4]
  assign _T_55793 = $signed(_T_55792); // @[Modules.scala 150:103:@1375.4]
  assign _T_55795 = $signed(4'sh1) * $signed(io_in_589); // @[Modules.scala 150:74:@1377.4]
  assign _T_55797 = $signed(4'sh1) * $signed(io_in_590); // @[Modules.scala 151:80:@1378.4]
  assign _T_55798 = $signed(_T_55795) + $signed(_T_55797); // @[Modules.scala 150:103:@1379.4]
  assign _T_55799 = _T_55798[5:0]; // @[Modules.scala 150:103:@1380.4]
  assign _T_55800 = $signed(_T_55799); // @[Modules.scala 150:103:@1381.4]
  assign _T_55802 = $signed(4'sh1) * $signed(io_in_591); // @[Modules.scala 150:74:@1383.4]
  assign _T_55804 = $signed(4'sh1) * $signed(io_in_592); // @[Modules.scala 151:80:@1384.4]
  assign _T_55805 = $signed(_T_55802) + $signed(_T_55804); // @[Modules.scala 150:103:@1385.4]
  assign _T_55806 = _T_55805[5:0]; // @[Modules.scala 150:103:@1386.4]
  assign _T_55807 = $signed(_T_55806); // @[Modules.scala 150:103:@1387.4]
  assign _T_55809 = $signed(4'sh1) * $signed(io_in_593); // @[Modules.scala 150:74:@1389.4]
  assign _T_55811 = $signed(4'sh1) * $signed(io_in_594); // @[Modules.scala 151:80:@1390.4]
  assign _T_55812 = $signed(_T_55809) + $signed(_T_55811); // @[Modules.scala 150:103:@1391.4]
  assign _T_55813 = _T_55812[5:0]; // @[Modules.scala 150:103:@1392.4]
  assign _T_55814 = $signed(_T_55813); // @[Modules.scala 150:103:@1393.4]
  assign _T_55816 = $signed(4'sh1) * $signed(io_in_596); // @[Modules.scala 150:74:@1395.4]
  assign _T_55818 = $signed(4'sh1) * $signed(io_in_598); // @[Modules.scala 151:80:@1396.4]
  assign _T_55819 = $signed(_T_55816) + $signed(_T_55818); // @[Modules.scala 150:103:@1397.4]
  assign _T_55820 = _T_55819[5:0]; // @[Modules.scala 150:103:@1398.4]
  assign _T_55821 = $signed(_T_55820); // @[Modules.scala 150:103:@1399.4]
  assign _T_55823 = $signed(4'sh1) * $signed(io_in_599); // @[Modules.scala 150:74:@1401.4]
  assign _T_55825 = $signed(4'sh1) * $signed(io_in_601); // @[Modules.scala 151:80:@1402.4]
  assign _T_55826 = $signed(_T_55823) + $signed(_T_55825); // @[Modules.scala 150:103:@1403.4]
  assign _T_55827 = _T_55826[5:0]; // @[Modules.scala 150:103:@1404.4]
  assign _T_55828 = $signed(_T_55827); // @[Modules.scala 150:103:@1405.4]
  assign _T_55830 = $signed(4'sh1) * $signed(io_in_602); // @[Modules.scala 150:74:@1407.4]
  assign _T_55832 = $signed(4'sh1) * $signed(io_in_603); // @[Modules.scala 151:80:@1408.4]
  assign _T_55833 = $signed(_T_55830) + $signed(_T_55832); // @[Modules.scala 150:103:@1409.4]
  assign _T_55834 = _T_55833[5:0]; // @[Modules.scala 150:103:@1410.4]
  assign _T_55835 = $signed(_T_55834); // @[Modules.scala 150:103:@1411.4]
  assign _T_55837 = $signed(-4'sh1) * $signed(io_in_608); // @[Modules.scala 150:74:@1413.4]
  assign _T_55839 = $signed(4'sh1) * $signed(io_in_609); // @[Modules.scala 151:80:@1414.4]
  assign _GEN_65 = {{1{_T_55837[4]}},_T_55837}; // @[Modules.scala 150:103:@1415.4]
  assign _T_55840 = $signed(_GEN_65) + $signed(_T_55839); // @[Modules.scala 150:103:@1415.4]
  assign _T_55841 = _T_55840[5:0]; // @[Modules.scala 150:103:@1416.4]
  assign _T_55842 = $signed(_T_55841); // @[Modules.scala 150:103:@1417.4]
  assign _T_55844 = $signed(4'sh1) * $signed(io_in_610); // @[Modules.scala 150:74:@1419.4]
  assign _T_55846 = $signed(4'sh1) * $signed(io_in_611); // @[Modules.scala 151:80:@1420.4]
  assign _T_55847 = $signed(_T_55844) + $signed(_T_55846); // @[Modules.scala 150:103:@1421.4]
  assign _T_55848 = _T_55847[5:0]; // @[Modules.scala 150:103:@1422.4]
  assign _T_55849 = $signed(_T_55848); // @[Modules.scala 150:103:@1423.4]
  assign _T_55851 = $signed(4'sh1) * $signed(io_in_612); // @[Modules.scala 150:74:@1425.4]
  assign _T_55853 = $signed(4'sh1) * $signed(io_in_613); // @[Modules.scala 151:80:@1426.4]
  assign _T_55854 = $signed(_T_55851) + $signed(_T_55853); // @[Modules.scala 150:103:@1427.4]
  assign _T_55855 = _T_55854[5:0]; // @[Modules.scala 150:103:@1428.4]
  assign _T_55856 = $signed(_T_55855); // @[Modules.scala 150:103:@1429.4]
  assign _T_55858 = $signed(4'sh1) * $signed(io_in_614); // @[Modules.scala 150:74:@1431.4]
  assign _T_55860 = $signed(4'sh1) * $signed(io_in_616); // @[Modules.scala 151:80:@1432.4]
  assign _T_55861 = $signed(_T_55858) + $signed(_T_55860); // @[Modules.scala 150:103:@1433.4]
  assign _T_55862 = _T_55861[5:0]; // @[Modules.scala 150:103:@1434.4]
  assign _T_55863 = $signed(_T_55862); // @[Modules.scala 150:103:@1435.4]
  assign _T_55865 = $signed(4'sh1) * $signed(io_in_617); // @[Modules.scala 150:74:@1437.4]
  assign _T_55867 = $signed(4'sh1) * $signed(io_in_618); // @[Modules.scala 151:80:@1438.4]
  assign _T_55868 = $signed(_T_55865) + $signed(_T_55867); // @[Modules.scala 150:103:@1439.4]
  assign _T_55869 = _T_55868[5:0]; // @[Modules.scala 150:103:@1440.4]
  assign _T_55870 = $signed(_T_55869); // @[Modules.scala 150:103:@1441.4]
  assign _T_55872 = $signed(4'sh1) * $signed(io_in_619); // @[Modules.scala 150:74:@1443.4]
  assign _T_55874 = $signed(4'sh1) * $signed(io_in_620); // @[Modules.scala 151:80:@1444.4]
  assign _T_55875 = $signed(_T_55872) + $signed(_T_55874); // @[Modules.scala 150:103:@1445.4]
  assign _T_55876 = _T_55875[5:0]; // @[Modules.scala 150:103:@1446.4]
  assign _T_55877 = $signed(_T_55876); // @[Modules.scala 150:103:@1447.4]
  assign _T_55879 = $signed(4'sh1) * $signed(io_in_621); // @[Modules.scala 150:74:@1449.4]
  assign _T_55881 = $signed(4'sh1) * $signed(io_in_622); // @[Modules.scala 151:80:@1450.4]
  assign _T_55882 = $signed(_T_55879) + $signed(_T_55881); // @[Modules.scala 150:103:@1451.4]
  assign _T_55883 = _T_55882[5:0]; // @[Modules.scala 150:103:@1452.4]
  assign _T_55884 = $signed(_T_55883); // @[Modules.scala 150:103:@1453.4]
  assign _T_55886 = $signed(-4'sh1) * $signed(io_in_623); // @[Modules.scala 150:74:@1455.4]
  assign _T_55888 = $signed(4'sh1) * $signed(io_in_625); // @[Modules.scala 151:80:@1456.4]
  assign _GEN_66 = {{1{_T_55886[4]}},_T_55886}; // @[Modules.scala 150:103:@1457.4]
  assign _T_55889 = $signed(_GEN_66) + $signed(_T_55888); // @[Modules.scala 150:103:@1457.4]
  assign _T_55890 = _T_55889[5:0]; // @[Modules.scala 150:103:@1458.4]
  assign _T_55891 = $signed(_T_55890); // @[Modules.scala 150:103:@1459.4]
  assign _T_55893 = $signed(-4'sh1) * $signed(io_in_627); // @[Modules.scala 150:74:@1461.4]
  assign _T_55895 = $signed(-4'sh1) * $signed(io_in_628); // @[Modules.scala 151:80:@1462.4]
  assign _T_55896 = $signed(_T_55893) + $signed(_T_55895); // @[Modules.scala 150:103:@1463.4]
  assign _T_55897 = _T_55896[4:0]; // @[Modules.scala 150:103:@1464.4]
  assign _T_55898 = $signed(_T_55897); // @[Modules.scala 150:103:@1465.4]
  assign _T_55900 = $signed(-4'sh1) * $signed(io_in_629); // @[Modules.scala 150:74:@1467.4]
  assign _T_55902 = $signed(-4'sh1) * $signed(io_in_630); // @[Modules.scala 151:80:@1468.4]
  assign _T_55903 = $signed(_T_55900) + $signed(_T_55902); // @[Modules.scala 150:103:@1469.4]
  assign _T_55904 = _T_55903[4:0]; // @[Modules.scala 150:103:@1470.4]
  assign _T_55905 = $signed(_T_55904); // @[Modules.scala 150:103:@1471.4]
  assign _T_55907 = $signed(-4'sh1) * $signed(io_in_631); // @[Modules.scala 150:74:@1473.4]
  assign _T_55909 = $signed(-4'sh1) * $signed(io_in_632); // @[Modules.scala 151:80:@1474.4]
  assign _T_55910 = $signed(_T_55907) + $signed(_T_55909); // @[Modules.scala 150:103:@1475.4]
  assign _T_55911 = _T_55910[4:0]; // @[Modules.scala 150:103:@1476.4]
  assign _T_55912 = $signed(_T_55911); // @[Modules.scala 150:103:@1477.4]
  assign _T_55914 = $signed(-4'sh1) * $signed(io_in_633); // @[Modules.scala 150:74:@1479.4]
  assign _T_55916 = $signed(-4'sh1) * $signed(io_in_634); // @[Modules.scala 151:80:@1480.4]
  assign _T_55917 = $signed(_T_55914) + $signed(_T_55916); // @[Modules.scala 150:103:@1481.4]
  assign _T_55918 = _T_55917[4:0]; // @[Modules.scala 150:103:@1482.4]
  assign _T_55919 = $signed(_T_55918); // @[Modules.scala 150:103:@1483.4]
  assign _T_55921 = $signed(4'sh1) * $signed(io_in_635); // @[Modules.scala 150:74:@1485.4]
  assign _T_55923 = $signed(4'sh1) * $signed(io_in_636); // @[Modules.scala 151:80:@1486.4]
  assign _T_55924 = $signed(_T_55921) + $signed(_T_55923); // @[Modules.scala 150:103:@1487.4]
  assign _T_55925 = _T_55924[5:0]; // @[Modules.scala 150:103:@1488.4]
  assign _T_55926 = $signed(_T_55925); // @[Modules.scala 150:103:@1489.4]
  assign _T_55928 = $signed(4'sh1) * $signed(io_in_637); // @[Modules.scala 150:74:@1491.4]
  assign _T_55930 = $signed(4'sh1) * $signed(io_in_638); // @[Modules.scala 151:80:@1492.4]
  assign _T_55931 = $signed(_T_55928) + $signed(_T_55930); // @[Modules.scala 150:103:@1493.4]
  assign _T_55932 = _T_55931[5:0]; // @[Modules.scala 150:103:@1494.4]
  assign _T_55933 = $signed(_T_55932); // @[Modules.scala 150:103:@1495.4]
  assign _T_55935 = $signed(4'sh1) * $signed(io_in_639); // @[Modules.scala 150:74:@1497.4]
  assign _T_55937 = $signed(4'sh1) * $signed(io_in_640); // @[Modules.scala 151:80:@1498.4]
  assign _T_55938 = $signed(_T_55935) + $signed(_T_55937); // @[Modules.scala 150:103:@1499.4]
  assign _T_55939 = _T_55938[5:0]; // @[Modules.scala 150:103:@1500.4]
  assign _T_55940 = $signed(_T_55939); // @[Modules.scala 150:103:@1501.4]
  assign _T_55942 = $signed(4'sh1) * $signed(io_in_641); // @[Modules.scala 150:74:@1503.4]
  assign _T_55944 = $signed(4'sh1) * $signed(io_in_642); // @[Modules.scala 151:80:@1504.4]
  assign _T_55945 = $signed(_T_55942) + $signed(_T_55944); // @[Modules.scala 150:103:@1505.4]
  assign _T_55946 = _T_55945[5:0]; // @[Modules.scala 150:103:@1506.4]
  assign _T_55947 = $signed(_T_55946); // @[Modules.scala 150:103:@1507.4]
  assign _T_55949 = $signed(4'sh1) * $signed(io_in_646); // @[Modules.scala 150:74:@1509.4]
  assign _T_55951 = $signed(4'sh1) * $signed(io_in_647); // @[Modules.scala 151:80:@1510.4]
  assign _T_55952 = $signed(_T_55949) + $signed(_T_55951); // @[Modules.scala 150:103:@1511.4]
  assign _T_55953 = _T_55952[5:0]; // @[Modules.scala 150:103:@1512.4]
  assign _T_55954 = $signed(_T_55953); // @[Modules.scala 150:103:@1513.4]
  assign _T_55956 = $signed(4'sh1) * $signed(io_in_648); // @[Modules.scala 150:74:@1515.4]
  assign _T_55958 = $signed(4'sh1) * $signed(io_in_649); // @[Modules.scala 151:80:@1516.4]
  assign _T_55959 = $signed(_T_55956) + $signed(_T_55958); // @[Modules.scala 150:103:@1517.4]
  assign _T_55960 = _T_55959[5:0]; // @[Modules.scala 150:103:@1518.4]
  assign _T_55961 = $signed(_T_55960); // @[Modules.scala 150:103:@1519.4]
  assign _T_55963 = $signed(4'sh1) * $signed(io_in_650); // @[Modules.scala 150:74:@1521.4]
  assign _T_55965 = $signed(4'sh1) * $signed(io_in_651); // @[Modules.scala 151:80:@1522.4]
  assign _T_55966 = $signed(_T_55963) + $signed(_T_55965); // @[Modules.scala 150:103:@1523.4]
  assign _T_55967 = _T_55966[5:0]; // @[Modules.scala 150:103:@1524.4]
  assign _T_55968 = $signed(_T_55967); // @[Modules.scala 150:103:@1525.4]
  assign _T_55970 = $signed(-4'sh1) * $signed(io_in_652); // @[Modules.scala 150:74:@1527.4]
  assign _T_55972 = $signed(-4'sh1) * $signed(io_in_653); // @[Modules.scala 151:80:@1528.4]
  assign _T_55973 = $signed(_T_55970) + $signed(_T_55972); // @[Modules.scala 150:103:@1529.4]
  assign _T_55974 = _T_55973[4:0]; // @[Modules.scala 150:103:@1530.4]
  assign _T_55975 = $signed(_T_55974); // @[Modules.scala 150:103:@1531.4]
  assign _T_55977 = $signed(-4'sh1) * $signed(io_in_654); // @[Modules.scala 150:74:@1533.4]
  assign _T_55979 = $signed(-4'sh1) * $signed(io_in_655); // @[Modules.scala 151:80:@1534.4]
  assign _T_55980 = $signed(_T_55977) + $signed(_T_55979); // @[Modules.scala 150:103:@1535.4]
  assign _T_55981 = _T_55980[4:0]; // @[Modules.scala 150:103:@1536.4]
  assign _T_55982 = $signed(_T_55981); // @[Modules.scala 150:103:@1537.4]
  assign _T_55984 = $signed(-4'sh1) * $signed(io_in_656); // @[Modules.scala 150:74:@1539.4]
  assign _T_55986 = $signed(-4'sh1) * $signed(io_in_657); // @[Modules.scala 151:80:@1540.4]
  assign _T_55987 = $signed(_T_55984) + $signed(_T_55986); // @[Modules.scala 150:103:@1541.4]
  assign _T_55988 = _T_55987[4:0]; // @[Modules.scala 150:103:@1542.4]
  assign _T_55989 = $signed(_T_55988); // @[Modules.scala 150:103:@1543.4]
  assign _T_55991 = $signed(-4'sh1) * $signed(io_in_658); // @[Modules.scala 150:74:@1545.4]
  assign _T_55993 = $signed(-4'sh1) * $signed(io_in_659); // @[Modules.scala 151:80:@1546.4]
  assign _T_55994 = $signed(_T_55991) + $signed(_T_55993); // @[Modules.scala 150:103:@1547.4]
  assign _T_55995 = _T_55994[4:0]; // @[Modules.scala 150:103:@1548.4]
  assign _T_55996 = $signed(_T_55995); // @[Modules.scala 150:103:@1549.4]
  assign _T_55998 = $signed(-4'sh1) * $signed(io_in_660); // @[Modules.scala 150:74:@1551.4]
  assign _T_56000 = $signed(-4'sh1) * $signed(io_in_661); // @[Modules.scala 151:80:@1552.4]
  assign _T_56001 = $signed(_T_55998) + $signed(_T_56000); // @[Modules.scala 150:103:@1553.4]
  assign _T_56002 = _T_56001[4:0]; // @[Modules.scala 150:103:@1554.4]
  assign _T_56003 = $signed(_T_56002); // @[Modules.scala 150:103:@1555.4]
  assign _T_56005 = $signed(-4'sh1) * $signed(io_in_662); // @[Modules.scala 150:74:@1557.4]
  assign _T_56007 = $signed(-4'sh1) * $signed(io_in_663); // @[Modules.scala 151:80:@1558.4]
  assign _T_56008 = $signed(_T_56005) + $signed(_T_56007); // @[Modules.scala 150:103:@1559.4]
  assign _T_56009 = _T_56008[4:0]; // @[Modules.scala 150:103:@1560.4]
  assign _T_56010 = $signed(_T_56009); // @[Modules.scala 150:103:@1561.4]
  assign _T_56012 = $signed(-4'sh1) * $signed(io_in_664); // @[Modules.scala 150:74:@1563.4]
  assign _T_56014 = $signed(-4'sh1) * $signed(io_in_665); // @[Modules.scala 151:80:@1564.4]
  assign _T_56015 = $signed(_T_56012) + $signed(_T_56014); // @[Modules.scala 150:103:@1565.4]
  assign _T_56016 = _T_56015[4:0]; // @[Modules.scala 150:103:@1566.4]
  assign _T_56017 = $signed(_T_56016); // @[Modules.scala 150:103:@1567.4]
  assign _T_56019 = $signed(4'sh1) * $signed(io_in_667); // @[Modules.scala 150:74:@1569.4]
  assign _T_56021 = $signed(4'sh1) * $signed(io_in_669); // @[Modules.scala 151:80:@1570.4]
  assign _T_56022 = $signed(_T_56019) + $signed(_T_56021); // @[Modules.scala 150:103:@1571.4]
  assign _T_56023 = _T_56022[5:0]; // @[Modules.scala 150:103:@1572.4]
  assign _T_56024 = $signed(_T_56023); // @[Modules.scala 150:103:@1573.4]
  assign _T_56026 = $signed(4'sh1) * $signed(io_in_670); // @[Modules.scala 150:74:@1575.4]
  assign _T_56028 = $signed(-4'sh1) * $signed(io_in_674); // @[Modules.scala 151:80:@1576.4]
  assign _GEN_67 = {{1{_T_56028[4]}},_T_56028}; // @[Modules.scala 150:103:@1577.4]
  assign _T_56029 = $signed(_T_56026) + $signed(_GEN_67); // @[Modules.scala 150:103:@1577.4]
  assign _T_56030 = _T_56029[5:0]; // @[Modules.scala 150:103:@1578.4]
  assign _T_56031 = $signed(_T_56030); // @[Modules.scala 150:103:@1579.4]
  assign _T_56033 = $signed(4'sh1) * $signed(io_in_675); // @[Modules.scala 150:74:@1581.4]
  assign _T_56035 = $signed(4'sh1) * $signed(io_in_676); // @[Modules.scala 151:80:@1582.4]
  assign _T_56036 = $signed(_T_56033) + $signed(_T_56035); // @[Modules.scala 150:103:@1583.4]
  assign _T_56037 = _T_56036[5:0]; // @[Modules.scala 150:103:@1584.4]
  assign _T_56038 = $signed(_T_56037); // @[Modules.scala 150:103:@1585.4]
  assign _T_56040 = $signed(4'sh1) * $signed(io_in_677); // @[Modules.scala 150:74:@1587.4]
  assign _T_56042 = $signed(4'sh1) * $signed(io_in_678); // @[Modules.scala 151:80:@1588.4]
  assign _T_56043 = $signed(_T_56040) + $signed(_T_56042); // @[Modules.scala 150:103:@1589.4]
  assign _T_56044 = _T_56043[5:0]; // @[Modules.scala 150:103:@1590.4]
  assign _T_56045 = $signed(_T_56044); // @[Modules.scala 150:103:@1591.4]
  assign _T_56047 = $signed(4'sh1) * $signed(io_in_679); // @[Modules.scala 150:74:@1593.4]
  assign _T_56049 = $signed(-4'sh1) * $signed(io_in_680); // @[Modules.scala 151:80:@1594.4]
  assign _GEN_68 = {{1{_T_56049[4]}},_T_56049}; // @[Modules.scala 150:103:@1595.4]
  assign _T_56050 = $signed(_T_56047) + $signed(_GEN_68); // @[Modules.scala 150:103:@1595.4]
  assign _T_56051 = _T_56050[5:0]; // @[Modules.scala 150:103:@1596.4]
  assign _T_56052 = $signed(_T_56051); // @[Modules.scala 150:103:@1597.4]
  assign _T_56054 = $signed(-4'sh1) * $signed(io_in_681); // @[Modules.scala 150:74:@1599.4]
  assign _T_56056 = $signed(-4'sh1) * $signed(io_in_682); // @[Modules.scala 151:80:@1600.4]
  assign _T_56057 = $signed(_T_56054) + $signed(_T_56056); // @[Modules.scala 150:103:@1601.4]
  assign _T_56058 = _T_56057[4:0]; // @[Modules.scala 150:103:@1602.4]
  assign _T_56059 = $signed(_T_56058); // @[Modules.scala 150:103:@1603.4]
  assign _T_56061 = $signed(-4'sh1) * $signed(io_in_685); // @[Modules.scala 150:74:@1605.4]
  assign _T_56063 = $signed(-4'sh1) * $signed(io_in_686); // @[Modules.scala 151:80:@1606.4]
  assign _T_56064 = $signed(_T_56061) + $signed(_T_56063); // @[Modules.scala 150:103:@1607.4]
  assign _T_56065 = _T_56064[4:0]; // @[Modules.scala 150:103:@1608.4]
  assign _T_56066 = $signed(_T_56065); // @[Modules.scala 150:103:@1609.4]
  assign _T_56068 = $signed(-4'sh1) * $signed(io_in_687); // @[Modules.scala 150:74:@1611.4]
  assign _T_56070 = $signed(-4'sh1) * $signed(io_in_688); // @[Modules.scala 151:80:@1612.4]
  assign _T_56071 = $signed(_T_56068) + $signed(_T_56070); // @[Modules.scala 150:103:@1613.4]
  assign _T_56072 = _T_56071[4:0]; // @[Modules.scala 150:103:@1614.4]
  assign _T_56073 = $signed(_T_56072); // @[Modules.scala 150:103:@1615.4]
  assign _T_56075 = $signed(-4'sh1) * $signed(io_in_689); // @[Modules.scala 150:74:@1617.4]
  assign _T_56077 = $signed(-4'sh1) * $signed(io_in_690); // @[Modules.scala 151:80:@1618.4]
  assign _T_56078 = $signed(_T_56075) + $signed(_T_56077); // @[Modules.scala 150:103:@1619.4]
  assign _T_56079 = _T_56078[4:0]; // @[Modules.scala 150:103:@1620.4]
  assign _T_56080 = $signed(_T_56079); // @[Modules.scala 150:103:@1621.4]
  assign _T_56082 = $signed(-4'sh1) * $signed(io_in_691); // @[Modules.scala 150:74:@1623.4]
  assign _T_56084 = $signed(-4'sh1) * $signed(io_in_692); // @[Modules.scala 151:80:@1624.4]
  assign _T_56085 = $signed(_T_56082) + $signed(_T_56084); // @[Modules.scala 150:103:@1625.4]
  assign _T_56086 = _T_56085[4:0]; // @[Modules.scala 150:103:@1626.4]
  assign _T_56087 = $signed(_T_56086); // @[Modules.scala 150:103:@1627.4]
  assign _T_56089 = $signed(-4'sh1) * $signed(io_in_693); // @[Modules.scala 150:74:@1629.4]
  assign _T_56091 = $signed(-4'sh1) * $signed(io_in_694); // @[Modules.scala 151:80:@1630.4]
  assign _T_56092 = $signed(_T_56089) + $signed(_T_56091); // @[Modules.scala 150:103:@1631.4]
  assign _T_56093 = _T_56092[4:0]; // @[Modules.scala 150:103:@1632.4]
  assign _T_56094 = $signed(_T_56093); // @[Modules.scala 150:103:@1633.4]
  assign _T_56096 = $signed(-4'sh1) * $signed(io_in_695); // @[Modules.scala 150:74:@1635.4]
  assign _T_56098 = $signed(4'sh1) * $signed(io_in_696); // @[Modules.scala 151:80:@1636.4]
  assign _GEN_69 = {{1{_T_56096[4]}},_T_56096}; // @[Modules.scala 150:103:@1637.4]
  assign _T_56099 = $signed(_GEN_69) + $signed(_T_56098); // @[Modules.scala 150:103:@1637.4]
  assign _T_56100 = _T_56099[5:0]; // @[Modules.scala 150:103:@1638.4]
  assign _T_56101 = $signed(_T_56100); // @[Modules.scala 150:103:@1639.4]
  assign _T_56103 = $signed(4'sh1) * $signed(io_in_697); // @[Modules.scala 150:74:@1641.4]
  assign _T_56105 = $signed(4'sh1) * $signed(io_in_698); // @[Modules.scala 151:80:@1642.4]
  assign _T_56106 = $signed(_T_56103) + $signed(_T_56105); // @[Modules.scala 150:103:@1643.4]
  assign _T_56107 = _T_56106[5:0]; // @[Modules.scala 150:103:@1644.4]
  assign _T_56108 = $signed(_T_56107); // @[Modules.scala 150:103:@1645.4]
  assign _T_56110 = $signed(4'sh1) * $signed(io_in_702); // @[Modules.scala 150:74:@1647.4]
  assign _T_56112 = $signed(4'sh1) * $signed(io_in_703); // @[Modules.scala 151:80:@1648.4]
  assign _T_56113 = $signed(_T_56110) + $signed(_T_56112); // @[Modules.scala 150:103:@1649.4]
  assign _T_56114 = _T_56113[5:0]; // @[Modules.scala 150:103:@1650.4]
  assign _T_56115 = $signed(_T_56114); // @[Modules.scala 150:103:@1651.4]
  assign _T_56117 = $signed(4'sh1) * $signed(io_in_704); // @[Modules.scala 150:74:@1653.4]
  assign _T_56119 = $signed(-4'sh1) * $signed(io_in_706); // @[Modules.scala 151:80:@1654.4]
  assign _GEN_70 = {{1{_T_56119[4]}},_T_56119}; // @[Modules.scala 150:103:@1655.4]
  assign _T_56120 = $signed(_T_56117) + $signed(_GEN_70); // @[Modules.scala 150:103:@1655.4]
  assign _T_56121 = _T_56120[5:0]; // @[Modules.scala 150:103:@1656.4]
  assign _T_56122 = $signed(_T_56121); // @[Modules.scala 150:103:@1657.4]
  assign _T_56124 = $signed(-4'sh1) * $signed(io_in_707); // @[Modules.scala 150:74:@1659.4]
  assign _T_56126 = $signed(4'sh1) * $signed(io_in_708); // @[Modules.scala 151:80:@1660.4]
  assign _GEN_71 = {{1{_T_56124[4]}},_T_56124}; // @[Modules.scala 150:103:@1661.4]
  assign _T_56127 = $signed(_GEN_71) + $signed(_T_56126); // @[Modules.scala 150:103:@1661.4]
  assign _T_56128 = _T_56127[5:0]; // @[Modules.scala 150:103:@1662.4]
  assign _T_56129 = $signed(_T_56128); // @[Modules.scala 150:103:@1663.4]
  assign _T_56131 = $signed(4'sh1) * $signed(io_in_709); // @[Modules.scala 150:74:@1665.4]
  assign _T_56133 = $signed(4'sh1) * $signed(io_in_710); // @[Modules.scala 151:80:@1666.4]
  assign _T_56134 = $signed(_T_56131) + $signed(_T_56133); // @[Modules.scala 150:103:@1667.4]
  assign _T_56135 = _T_56134[5:0]; // @[Modules.scala 150:103:@1668.4]
  assign _T_56136 = $signed(_T_56135); // @[Modules.scala 150:103:@1669.4]
  assign _T_56138 = $signed(4'sh1) * $signed(io_in_711); // @[Modules.scala 150:74:@1671.4]
  assign _T_56140 = $signed(4'sh1) * $signed(io_in_712); // @[Modules.scala 151:80:@1672.4]
  assign _T_56141 = $signed(_T_56138) + $signed(_T_56140); // @[Modules.scala 150:103:@1673.4]
  assign _T_56142 = _T_56141[5:0]; // @[Modules.scala 150:103:@1674.4]
  assign _T_56143 = $signed(_T_56142); // @[Modules.scala 150:103:@1675.4]
  assign _T_56145 = $signed(-4'sh1) * $signed(io_in_713); // @[Modules.scala 150:74:@1677.4]
  assign _T_56147 = $signed(-4'sh1) * $signed(io_in_714); // @[Modules.scala 151:80:@1678.4]
  assign _T_56148 = $signed(_T_56145) + $signed(_T_56147); // @[Modules.scala 150:103:@1679.4]
  assign _T_56149 = _T_56148[4:0]; // @[Modules.scala 150:103:@1680.4]
  assign _T_56150 = $signed(_T_56149); // @[Modules.scala 150:103:@1681.4]
  assign _T_56152 = $signed(-4'sh1) * $signed(io_in_715); // @[Modules.scala 150:74:@1683.4]
  assign _T_56154 = $signed(-4'sh1) * $signed(io_in_716); // @[Modules.scala 151:80:@1684.4]
  assign _T_56155 = $signed(_T_56152) + $signed(_T_56154); // @[Modules.scala 150:103:@1685.4]
  assign _T_56156 = _T_56155[4:0]; // @[Modules.scala 150:103:@1686.4]
  assign _T_56157 = $signed(_T_56156); // @[Modules.scala 150:103:@1687.4]
  assign _T_56159 = $signed(-4'sh1) * $signed(io_in_717); // @[Modules.scala 150:74:@1689.4]
  assign _T_56161 = $signed(-4'sh1) * $signed(io_in_718); // @[Modules.scala 151:80:@1690.4]
  assign _T_56162 = $signed(_T_56159) + $signed(_T_56161); // @[Modules.scala 150:103:@1691.4]
  assign _T_56163 = _T_56162[4:0]; // @[Modules.scala 150:103:@1692.4]
  assign _T_56164 = $signed(_T_56163); // @[Modules.scala 150:103:@1693.4]
  assign _T_56166 = $signed(-4'sh1) * $signed(io_in_719); // @[Modules.scala 150:74:@1695.4]
  assign _T_56168 = $signed(-4'sh1) * $signed(io_in_720); // @[Modules.scala 151:80:@1696.4]
  assign _T_56169 = $signed(_T_56166) + $signed(_T_56168); // @[Modules.scala 150:103:@1697.4]
  assign _T_56170 = _T_56169[4:0]; // @[Modules.scala 150:103:@1698.4]
  assign _T_56171 = $signed(_T_56170); // @[Modules.scala 150:103:@1699.4]
  assign _T_56173 = $signed(-4'sh1) * $signed(io_in_721); // @[Modules.scala 150:74:@1701.4]
  assign _T_56175 = $signed(-4'sh1) * $signed(io_in_722); // @[Modules.scala 151:80:@1702.4]
  assign _T_56176 = $signed(_T_56173) + $signed(_T_56175); // @[Modules.scala 150:103:@1703.4]
  assign _T_56177 = _T_56176[4:0]; // @[Modules.scala 150:103:@1704.4]
  assign _T_56178 = $signed(_T_56177); // @[Modules.scala 150:103:@1705.4]
  assign _T_56180 = $signed(-4'sh1) * $signed(io_in_723); // @[Modules.scala 150:74:@1707.4]
  assign _T_56182 = $signed(-4'sh1) * $signed(io_in_724); // @[Modules.scala 151:80:@1708.4]
  assign _T_56183 = $signed(_T_56180) + $signed(_T_56182); // @[Modules.scala 150:103:@1709.4]
  assign _T_56184 = _T_56183[4:0]; // @[Modules.scala 150:103:@1710.4]
  assign _T_56185 = $signed(_T_56184); // @[Modules.scala 150:103:@1711.4]
  assign _T_56187 = $signed(-4'sh1) * $signed(io_in_725); // @[Modules.scala 150:74:@1713.4]
  assign _T_56189 = $signed(-4'sh1) * $signed(io_in_726); // @[Modules.scala 151:80:@1714.4]
  assign _T_56190 = $signed(_T_56187) + $signed(_T_56189); // @[Modules.scala 150:103:@1715.4]
  assign _T_56191 = _T_56190[4:0]; // @[Modules.scala 150:103:@1716.4]
  assign _T_56192 = $signed(_T_56191); // @[Modules.scala 150:103:@1717.4]
  assign _T_56194 = $signed(-4'sh1) * $signed(io_in_731); // @[Modules.scala 150:74:@1719.4]
  assign _T_56196 = $signed(4'sh1) * $signed(io_in_736); // @[Modules.scala 151:80:@1720.4]
  assign _GEN_72 = {{1{_T_56194[4]}},_T_56194}; // @[Modules.scala 150:103:@1721.4]
  assign _T_56197 = $signed(_GEN_72) + $signed(_T_56196); // @[Modules.scala 150:103:@1721.4]
  assign _T_56198 = _T_56197[5:0]; // @[Modules.scala 150:103:@1722.4]
  assign _T_56199 = $signed(_T_56198); // @[Modules.scala 150:103:@1723.4]
  assign _T_56201 = $signed(4'sh1) * $signed(io_in_737); // @[Modules.scala 150:74:@1725.4]
  assign _T_56203 = $signed(4'sh1) * $signed(io_in_738); // @[Modules.scala 151:80:@1726.4]
  assign _T_56204 = $signed(_T_56201) + $signed(_T_56203); // @[Modules.scala 150:103:@1727.4]
  assign _T_56205 = _T_56204[5:0]; // @[Modules.scala 150:103:@1728.4]
  assign _T_56206 = $signed(_T_56205); // @[Modules.scala 150:103:@1729.4]
  assign _T_56208 = $signed(4'sh1) * $signed(io_in_739); // @[Modules.scala 150:74:@1731.4]
  assign _T_56210 = $signed(4'sh1) * $signed(io_in_740); // @[Modules.scala 151:80:@1732.4]
  assign _T_56211 = $signed(_T_56208) + $signed(_T_56210); // @[Modules.scala 150:103:@1733.4]
  assign _T_56212 = _T_56211[5:0]; // @[Modules.scala 150:103:@1734.4]
  assign _T_56213 = $signed(_T_56212); // @[Modules.scala 150:103:@1735.4]
  assign _T_56215 = $signed(-4'sh1) * $signed(io_in_742); // @[Modules.scala 150:74:@1737.4]
  assign _T_56217 = $signed(4'sh1) * $signed(io_in_744); // @[Modules.scala 151:80:@1738.4]
  assign _GEN_73 = {{1{_T_56215[4]}},_T_56215}; // @[Modules.scala 150:103:@1739.4]
  assign _T_56218 = $signed(_GEN_73) + $signed(_T_56217); // @[Modules.scala 150:103:@1739.4]
  assign _T_56219 = _T_56218[5:0]; // @[Modules.scala 150:103:@1740.4]
  assign _T_56220 = $signed(_T_56219); // @[Modules.scala 150:103:@1741.4]
  assign _T_56222 = $signed(4'sh1) * $signed(io_in_745); // @[Modules.scala 150:74:@1743.4]
  assign _T_56224 = $signed(-4'sh1) * $signed(io_in_746); // @[Modules.scala 151:80:@1744.4]
  assign _GEN_74 = {{1{_T_56224[4]}},_T_56224}; // @[Modules.scala 150:103:@1745.4]
  assign _T_56225 = $signed(_T_56222) + $signed(_GEN_74); // @[Modules.scala 150:103:@1745.4]
  assign _T_56226 = _T_56225[5:0]; // @[Modules.scala 150:103:@1746.4]
  assign _T_56227 = $signed(_T_56226); // @[Modules.scala 150:103:@1747.4]
  assign _T_56229 = $signed(-4'sh1) * $signed(io_in_747); // @[Modules.scala 150:74:@1749.4]
  assign _T_56231 = $signed(-4'sh1) * $signed(io_in_748); // @[Modules.scala 151:80:@1750.4]
  assign _T_56232 = $signed(_T_56229) + $signed(_T_56231); // @[Modules.scala 150:103:@1751.4]
  assign _T_56233 = _T_56232[4:0]; // @[Modules.scala 150:103:@1752.4]
  assign _T_56234 = $signed(_T_56233); // @[Modules.scala 150:103:@1753.4]
  assign _T_56236 = $signed(-4'sh1) * $signed(io_in_749); // @[Modules.scala 150:74:@1755.4]
  assign _T_56238 = $signed(-4'sh1) * $signed(io_in_750); // @[Modules.scala 151:80:@1756.4]
  assign _T_56239 = $signed(_T_56236) + $signed(_T_56238); // @[Modules.scala 150:103:@1757.4]
  assign _T_56240 = _T_56239[4:0]; // @[Modules.scala 150:103:@1758.4]
  assign _T_56241 = $signed(_T_56240); // @[Modules.scala 150:103:@1759.4]
  assign _T_56243 = $signed(-4'sh1) * $signed(io_in_751); // @[Modules.scala 150:74:@1761.4]
  assign _T_56245 = $signed(4'sh1) * $signed(io_in_752); // @[Modules.scala 151:80:@1762.4]
  assign _GEN_75 = {{1{_T_56243[4]}},_T_56243}; // @[Modules.scala 150:103:@1763.4]
  assign _T_56246 = $signed(_GEN_75) + $signed(_T_56245); // @[Modules.scala 150:103:@1763.4]
  assign _T_56247 = _T_56246[5:0]; // @[Modules.scala 150:103:@1764.4]
  assign _T_56248 = $signed(_T_56247); // @[Modules.scala 150:103:@1765.4]
  assign _T_56250 = $signed(4'sh1) * $signed(io_in_760); // @[Modules.scala 150:74:@1767.4]
  assign _T_56252 = $signed(4'sh1) * $signed(io_in_761); // @[Modules.scala 151:80:@1768.4]
  assign _T_56253 = $signed(_T_56250) + $signed(_T_56252); // @[Modules.scala 150:103:@1769.4]
  assign _T_56254 = _T_56253[5:0]; // @[Modules.scala 150:103:@1770.4]
  assign _T_56255 = $signed(_T_56254); // @[Modules.scala 150:103:@1771.4]
  assign _T_56257 = $signed(-4'sh1) * $signed(io_in_763); // @[Modules.scala 150:74:@1773.4]
  assign _T_56259 = $signed(-4'sh1) * $signed(io_in_764); // @[Modules.scala 151:80:@1774.4]
  assign _T_56260 = $signed(_T_56257) + $signed(_T_56259); // @[Modules.scala 150:103:@1775.4]
  assign _T_56261 = _T_56260[4:0]; // @[Modules.scala 150:103:@1776.4]
  assign _T_56262 = $signed(_T_56261); // @[Modules.scala 150:103:@1777.4]
  assign _T_56264 = $signed(4'sh1) * $signed(io_in_765); // @[Modules.scala 150:74:@1779.4]
  assign _T_56266 = $signed(4'sh1) * $signed(io_in_766); // @[Modules.scala 151:80:@1780.4]
  assign _T_56267 = $signed(_T_56264) + $signed(_T_56266); // @[Modules.scala 150:103:@1781.4]
  assign _T_56268 = _T_56267[5:0]; // @[Modules.scala 150:103:@1782.4]
  assign _T_56269 = $signed(_T_56268); // @[Modules.scala 150:103:@1783.4]
  assign _T_56271 = $signed(4'sh1) * $signed(io_in_767); // @[Modules.scala 150:74:@1785.4]
  assign _T_56273 = $signed(4'sh1) * $signed(io_in_769); // @[Modules.scala 151:80:@1786.4]
  assign _T_56274 = $signed(_T_56271) + $signed(_T_56273); // @[Modules.scala 150:103:@1787.4]
  assign _T_56275 = _T_56274[5:0]; // @[Modules.scala 150:103:@1788.4]
  assign _T_56276 = $signed(_T_56275); // @[Modules.scala 150:103:@1789.4]
  assign _T_56278 = $signed(4'sh1) * $signed(io_in_770); // @[Modules.scala 150:74:@1791.4]
  assign _T_56280 = $signed(4'sh1) * $signed(io_in_771); // @[Modules.scala 151:80:@1792.4]
  assign _T_56281 = $signed(_T_56278) + $signed(_T_56280); // @[Modules.scala 150:103:@1793.4]
  assign _T_56282 = _T_56281[5:0]; // @[Modules.scala 150:103:@1794.4]
  assign _T_56283 = $signed(_T_56282); // @[Modules.scala 150:103:@1795.4]
  assign _T_56285 = $signed(4'sh1) * $signed(io_in_772); // @[Modules.scala 150:74:@1797.4]
  assign _T_56287 = $signed(4'sh1) * $signed(io_in_773); // @[Modules.scala 151:80:@1798.4]
  assign _T_56288 = $signed(_T_56285) + $signed(_T_56287); // @[Modules.scala 150:103:@1799.4]
  assign _T_56289 = _T_56288[5:0]; // @[Modules.scala 150:103:@1800.4]
  assign _T_56290 = $signed(_T_56289); // @[Modules.scala 150:103:@1801.4]
  assign _T_56292 = $signed(-4'sh1) * $signed(io_in_775); // @[Modules.scala 150:74:@1803.4]
  assign _T_56294 = $signed(-4'sh1) * $signed(io_in_776); // @[Modules.scala 151:80:@1804.4]
  assign _T_56295 = $signed(_T_56292) + $signed(_T_56294); // @[Modules.scala 150:103:@1805.4]
  assign _T_56296 = _T_56295[4:0]; // @[Modules.scala 150:103:@1806.4]
  assign _T_56297 = $signed(_T_56296); // @[Modules.scala 150:103:@1807.4]
  assign _T_56299 = $signed(4'sh1) * $signed(io_in_777); // @[Modules.scala 150:74:@1809.4]
  assign _T_56301 = $signed(4'sh1) * $signed(io_in_778); // @[Modules.scala 151:80:@1810.4]
  assign _T_56302 = $signed(_T_56299) + $signed(_T_56301); // @[Modules.scala 150:103:@1811.4]
  assign _T_56303 = _T_56302[5:0]; // @[Modules.scala 150:103:@1812.4]
  assign _T_56304 = $signed(_T_56303); // @[Modules.scala 150:103:@1813.4]
  assign _T_56306 = $signed(4'sh1) * $signed(io_in_779); // @[Modules.scala 153:80:@1815.4]
  assign buffer_0_0 = {{8{_T_54204[5]}},_T_54204}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_1 = {{8{_T_54211[5]}},_T_54211}; // @[Modules.scala 112:22:@8.4]
  assign _T_56307 = $signed(buffer_0_0) + $signed(buffer_0_1); // @[Modules.scala 160:64:@1817.4]
  assign _T_56308 = _T_56307[13:0]; // @[Modules.scala 160:64:@1818.4]
  assign buffer_0_302 = $signed(_T_56308); // @[Modules.scala 160:64:@1819.4]
  assign buffer_0_2 = {{8{_T_54218[5]}},_T_54218}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_3 = {{8{_T_54225[5]}},_T_54225}; // @[Modules.scala 112:22:@8.4]
  assign _T_56310 = $signed(buffer_0_2) + $signed(buffer_0_3); // @[Modules.scala 160:64:@1821.4]
  assign _T_56311 = _T_56310[13:0]; // @[Modules.scala 160:64:@1822.4]
  assign buffer_0_303 = $signed(_T_56311); // @[Modules.scala 160:64:@1823.4]
  assign buffer_0_4 = {{8{_T_54232[5]}},_T_54232}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_5 = {{8{_T_54239[5]}},_T_54239}; // @[Modules.scala 112:22:@8.4]
  assign _T_56313 = $signed(buffer_0_4) + $signed(buffer_0_5); // @[Modules.scala 160:64:@1825.4]
  assign _T_56314 = _T_56313[13:0]; // @[Modules.scala 160:64:@1826.4]
  assign buffer_0_304 = $signed(_T_56314); // @[Modules.scala 160:64:@1827.4]
  assign buffer_0_6 = {{8{_T_54246[5]}},_T_54246}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_7 = {{8{_T_54253[5]}},_T_54253}; // @[Modules.scala 112:22:@8.4]
  assign _T_56316 = $signed(buffer_0_6) + $signed(buffer_0_7); // @[Modules.scala 160:64:@1829.4]
  assign _T_56317 = _T_56316[13:0]; // @[Modules.scala 160:64:@1830.4]
  assign buffer_0_305 = $signed(_T_56317); // @[Modules.scala 160:64:@1831.4]
  assign buffer_0_8 = {{8{_T_54260[5]}},_T_54260}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_9 = {{8{_T_54267[5]}},_T_54267}; // @[Modules.scala 112:22:@8.4]
  assign _T_56319 = $signed(buffer_0_8) + $signed(buffer_0_9); // @[Modules.scala 160:64:@1833.4]
  assign _T_56320 = _T_56319[13:0]; // @[Modules.scala 160:64:@1834.4]
  assign buffer_0_306 = $signed(_T_56320); // @[Modules.scala 160:64:@1835.4]
  assign buffer_0_10 = {{8{_T_54274[5]}},_T_54274}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_11 = {{8{_T_54281[5]}},_T_54281}; // @[Modules.scala 112:22:@8.4]
  assign _T_56322 = $signed(buffer_0_10) + $signed(buffer_0_11); // @[Modules.scala 160:64:@1837.4]
  assign _T_56323 = _T_56322[13:0]; // @[Modules.scala 160:64:@1838.4]
  assign buffer_0_307 = $signed(_T_56323); // @[Modules.scala 160:64:@1839.4]
  assign buffer_0_12 = {{8{_T_54288[5]}},_T_54288}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_13 = {{8{_T_54295[5]}},_T_54295}; // @[Modules.scala 112:22:@8.4]
  assign _T_56325 = $signed(buffer_0_12) + $signed(buffer_0_13); // @[Modules.scala 160:64:@1841.4]
  assign _T_56326 = _T_56325[13:0]; // @[Modules.scala 160:64:@1842.4]
  assign buffer_0_308 = $signed(_T_56326); // @[Modules.scala 160:64:@1843.4]
  assign buffer_0_14 = {{8{_T_54302[5]}},_T_54302}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_15 = {{8{_T_54309[5]}},_T_54309}; // @[Modules.scala 112:22:@8.4]
  assign _T_56328 = $signed(buffer_0_14) + $signed(buffer_0_15); // @[Modules.scala 160:64:@1845.4]
  assign _T_56329 = _T_56328[13:0]; // @[Modules.scala 160:64:@1846.4]
  assign buffer_0_309 = $signed(_T_56329); // @[Modules.scala 160:64:@1847.4]
  assign buffer_0_16 = {{8{_T_54316[5]}},_T_54316}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_17 = {{8{_T_54323[5]}},_T_54323}; // @[Modules.scala 112:22:@8.4]
  assign _T_56331 = $signed(buffer_0_16) + $signed(buffer_0_17); // @[Modules.scala 160:64:@1849.4]
  assign _T_56332 = _T_56331[13:0]; // @[Modules.scala 160:64:@1850.4]
  assign buffer_0_310 = $signed(_T_56332); // @[Modules.scala 160:64:@1851.4]
  assign buffer_0_18 = {{8{_T_54330[5]}},_T_54330}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_19 = {{8{_T_54337[5]}},_T_54337}; // @[Modules.scala 112:22:@8.4]
  assign _T_56334 = $signed(buffer_0_18) + $signed(buffer_0_19); // @[Modules.scala 160:64:@1853.4]
  assign _T_56335 = _T_56334[13:0]; // @[Modules.scala 160:64:@1854.4]
  assign buffer_0_311 = $signed(_T_56335); // @[Modules.scala 160:64:@1855.4]
  assign buffer_0_20 = {{8{_T_54344[5]}},_T_54344}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_21 = {{8{_T_54351[5]}},_T_54351}; // @[Modules.scala 112:22:@8.4]
  assign _T_56337 = $signed(buffer_0_20) + $signed(buffer_0_21); // @[Modules.scala 160:64:@1857.4]
  assign _T_56338 = _T_56337[13:0]; // @[Modules.scala 160:64:@1858.4]
  assign buffer_0_312 = $signed(_T_56338); // @[Modules.scala 160:64:@1859.4]
  assign buffer_0_22 = {{8{_T_54358[5]}},_T_54358}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_23 = {{8{_T_54365[5]}},_T_54365}; // @[Modules.scala 112:22:@8.4]
  assign _T_56340 = $signed(buffer_0_22) + $signed(buffer_0_23); // @[Modules.scala 160:64:@1861.4]
  assign _T_56341 = _T_56340[13:0]; // @[Modules.scala 160:64:@1862.4]
  assign buffer_0_313 = $signed(_T_56341); // @[Modules.scala 160:64:@1863.4]
  assign buffer_0_24 = {{8{_T_54372[5]}},_T_54372}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_25 = {{8{_T_54379[5]}},_T_54379}; // @[Modules.scala 112:22:@8.4]
  assign _T_56343 = $signed(buffer_0_24) + $signed(buffer_0_25); // @[Modules.scala 160:64:@1865.4]
  assign _T_56344 = _T_56343[13:0]; // @[Modules.scala 160:64:@1866.4]
  assign buffer_0_314 = $signed(_T_56344); // @[Modules.scala 160:64:@1867.4]
  assign buffer_0_26 = {{8{_T_54386[5]}},_T_54386}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_27 = {{8{_T_54393[5]}},_T_54393}; // @[Modules.scala 112:22:@8.4]
  assign _T_56346 = $signed(buffer_0_26) + $signed(buffer_0_27); // @[Modules.scala 160:64:@1869.4]
  assign _T_56347 = _T_56346[13:0]; // @[Modules.scala 160:64:@1870.4]
  assign buffer_0_315 = $signed(_T_56347); // @[Modules.scala 160:64:@1871.4]
  assign buffer_0_28 = {{8{_T_54400[5]}},_T_54400}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_29 = {{8{_T_54407[5]}},_T_54407}; // @[Modules.scala 112:22:@8.4]
  assign _T_56349 = $signed(buffer_0_28) + $signed(buffer_0_29); // @[Modules.scala 160:64:@1873.4]
  assign _T_56350 = _T_56349[13:0]; // @[Modules.scala 160:64:@1874.4]
  assign buffer_0_316 = $signed(_T_56350); // @[Modules.scala 160:64:@1875.4]
  assign buffer_0_30 = {{8{_T_54414[5]}},_T_54414}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_31 = {{8{_T_54421[5]}},_T_54421}; // @[Modules.scala 112:22:@8.4]
  assign _T_56352 = $signed(buffer_0_30) + $signed(buffer_0_31); // @[Modules.scala 160:64:@1877.4]
  assign _T_56353 = _T_56352[13:0]; // @[Modules.scala 160:64:@1878.4]
  assign buffer_0_317 = $signed(_T_56353); // @[Modules.scala 160:64:@1879.4]
  assign buffer_0_32 = {{8{_T_54428[5]}},_T_54428}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_33 = {{8{_T_54435[5]}},_T_54435}; // @[Modules.scala 112:22:@8.4]
  assign _T_56355 = $signed(buffer_0_32) + $signed(buffer_0_33); // @[Modules.scala 160:64:@1881.4]
  assign _T_56356 = _T_56355[13:0]; // @[Modules.scala 160:64:@1882.4]
  assign buffer_0_318 = $signed(_T_56356); // @[Modules.scala 160:64:@1883.4]
  assign buffer_0_34 = {{8{_T_54442[5]}},_T_54442}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_35 = {{8{_T_54449[5]}},_T_54449}; // @[Modules.scala 112:22:@8.4]
  assign _T_56358 = $signed(buffer_0_34) + $signed(buffer_0_35); // @[Modules.scala 160:64:@1885.4]
  assign _T_56359 = _T_56358[13:0]; // @[Modules.scala 160:64:@1886.4]
  assign buffer_0_319 = $signed(_T_56359); // @[Modules.scala 160:64:@1887.4]
  assign buffer_0_36 = {{8{_T_54456[5]}},_T_54456}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_37 = {{8{_T_54463[5]}},_T_54463}; // @[Modules.scala 112:22:@8.4]
  assign _T_56361 = $signed(buffer_0_36) + $signed(buffer_0_37); // @[Modules.scala 160:64:@1889.4]
  assign _T_56362 = _T_56361[13:0]; // @[Modules.scala 160:64:@1890.4]
  assign buffer_0_320 = $signed(_T_56362); // @[Modules.scala 160:64:@1891.4]
  assign buffer_0_38 = {{8{_T_54470[5]}},_T_54470}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_39 = {{8{_T_54477[5]}},_T_54477}; // @[Modules.scala 112:22:@8.4]
  assign _T_56364 = $signed(buffer_0_38) + $signed(buffer_0_39); // @[Modules.scala 160:64:@1893.4]
  assign _T_56365 = _T_56364[13:0]; // @[Modules.scala 160:64:@1894.4]
  assign buffer_0_321 = $signed(_T_56365); // @[Modules.scala 160:64:@1895.4]
  assign buffer_0_40 = {{8{_T_54484[5]}},_T_54484}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_41 = {{8{_T_54491[5]}},_T_54491}; // @[Modules.scala 112:22:@8.4]
  assign _T_56367 = $signed(buffer_0_40) + $signed(buffer_0_41); // @[Modules.scala 160:64:@1897.4]
  assign _T_56368 = _T_56367[13:0]; // @[Modules.scala 160:64:@1898.4]
  assign buffer_0_322 = $signed(_T_56368); // @[Modules.scala 160:64:@1899.4]
  assign buffer_0_42 = {{8{_T_54498[5]}},_T_54498}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_43 = {{8{_T_54505[5]}},_T_54505}; // @[Modules.scala 112:22:@8.4]
  assign _T_56370 = $signed(buffer_0_42) + $signed(buffer_0_43); // @[Modules.scala 160:64:@1901.4]
  assign _T_56371 = _T_56370[13:0]; // @[Modules.scala 160:64:@1902.4]
  assign buffer_0_323 = $signed(_T_56371); // @[Modules.scala 160:64:@1903.4]
  assign buffer_0_44 = {{9{_T_54512[4]}},_T_54512}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_45 = {{8{_T_54519[5]}},_T_54519}; // @[Modules.scala 112:22:@8.4]
  assign _T_56373 = $signed(buffer_0_44) + $signed(buffer_0_45); // @[Modules.scala 160:64:@1905.4]
  assign _T_56374 = _T_56373[13:0]; // @[Modules.scala 160:64:@1906.4]
  assign buffer_0_324 = $signed(_T_56374); // @[Modules.scala 160:64:@1907.4]
  assign buffer_0_46 = {{8{_T_54526[5]}},_T_54526}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_47 = {{8{_T_54533[5]}},_T_54533}; // @[Modules.scala 112:22:@8.4]
  assign _T_56376 = $signed(buffer_0_46) + $signed(buffer_0_47); // @[Modules.scala 160:64:@1909.4]
  assign _T_56377 = _T_56376[13:0]; // @[Modules.scala 160:64:@1910.4]
  assign buffer_0_325 = $signed(_T_56377); // @[Modules.scala 160:64:@1911.4]
  assign buffer_0_48 = {{8{_T_54540[5]}},_T_54540}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_49 = {{8{_T_54547[5]}},_T_54547}; // @[Modules.scala 112:22:@8.4]
  assign _T_56379 = $signed(buffer_0_48) + $signed(buffer_0_49); // @[Modules.scala 160:64:@1913.4]
  assign _T_56380 = _T_56379[13:0]; // @[Modules.scala 160:64:@1914.4]
  assign buffer_0_326 = $signed(_T_56380); // @[Modules.scala 160:64:@1915.4]
  assign buffer_0_50 = {{9{_T_54554[4]}},_T_54554}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_51 = {{8{_T_54561[5]}},_T_54561}; // @[Modules.scala 112:22:@8.4]
  assign _T_56382 = $signed(buffer_0_50) + $signed(buffer_0_51); // @[Modules.scala 160:64:@1917.4]
  assign _T_56383 = _T_56382[13:0]; // @[Modules.scala 160:64:@1918.4]
  assign buffer_0_327 = $signed(_T_56383); // @[Modules.scala 160:64:@1919.4]
  assign buffer_0_52 = {{9{_T_54568[4]}},_T_54568}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_53 = {{8{_T_54575[5]}},_T_54575}; // @[Modules.scala 112:22:@8.4]
  assign _T_56385 = $signed(buffer_0_52) + $signed(buffer_0_53); // @[Modules.scala 160:64:@1921.4]
  assign _T_56386 = _T_56385[13:0]; // @[Modules.scala 160:64:@1922.4]
  assign buffer_0_328 = $signed(_T_56386); // @[Modules.scala 160:64:@1923.4]
  assign buffer_0_54 = {{8{_T_54582[5]}},_T_54582}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_55 = {{8{_T_54589[5]}},_T_54589}; // @[Modules.scala 112:22:@8.4]
  assign _T_56388 = $signed(buffer_0_54) + $signed(buffer_0_55); // @[Modules.scala 160:64:@1925.4]
  assign _T_56389 = _T_56388[13:0]; // @[Modules.scala 160:64:@1926.4]
  assign buffer_0_329 = $signed(_T_56389); // @[Modules.scala 160:64:@1927.4]
  assign buffer_0_56 = {{8{_T_54596[5]}},_T_54596}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_57 = {{8{_T_54603[5]}},_T_54603}; // @[Modules.scala 112:22:@8.4]
  assign _T_56391 = $signed(buffer_0_56) + $signed(buffer_0_57); // @[Modules.scala 160:64:@1929.4]
  assign _T_56392 = _T_56391[13:0]; // @[Modules.scala 160:64:@1930.4]
  assign buffer_0_330 = $signed(_T_56392); // @[Modules.scala 160:64:@1931.4]
  assign buffer_0_58 = {{8{_T_54610[5]}},_T_54610}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_59 = {{9{_T_54617[4]}},_T_54617}; // @[Modules.scala 112:22:@8.4]
  assign _T_56394 = $signed(buffer_0_58) + $signed(buffer_0_59); // @[Modules.scala 160:64:@1933.4]
  assign _T_56395 = _T_56394[13:0]; // @[Modules.scala 160:64:@1934.4]
  assign buffer_0_331 = $signed(_T_56395); // @[Modules.scala 160:64:@1935.4]
  assign buffer_0_60 = {{9{_T_54624[4]}},_T_54624}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_61 = {{9{_T_54631[4]}},_T_54631}; // @[Modules.scala 112:22:@8.4]
  assign _T_56397 = $signed(buffer_0_60) + $signed(buffer_0_61); // @[Modules.scala 160:64:@1937.4]
  assign _T_56398 = _T_56397[13:0]; // @[Modules.scala 160:64:@1938.4]
  assign buffer_0_332 = $signed(_T_56398); // @[Modules.scala 160:64:@1939.4]
  assign buffer_0_62 = {{9{_T_54638[4]}},_T_54638}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_63 = {{9{_T_54645[4]}},_T_54645}; // @[Modules.scala 112:22:@8.4]
  assign _T_56400 = $signed(buffer_0_62) + $signed(buffer_0_63); // @[Modules.scala 160:64:@1941.4]
  assign _T_56401 = _T_56400[13:0]; // @[Modules.scala 160:64:@1942.4]
  assign buffer_0_333 = $signed(_T_56401); // @[Modules.scala 160:64:@1943.4]
  assign buffer_0_64 = {{9{_T_54652[4]}},_T_54652}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_65 = {{8{_T_54659[5]}},_T_54659}; // @[Modules.scala 112:22:@8.4]
  assign _T_56403 = $signed(buffer_0_64) + $signed(buffer_0_65); // @[Modules.scala 160:64:@1945.4]
  assign _T_56404 = _T_56403[13:0]; // @[Modules.scala 160:64:@1946.4]
  assign buffer_0_334 = $signed(_T_56404); // @[Modules.scala 160:64:@1947.4]
  assign buffer_0_66 = {{8{_T_54666[5]}},_T_54666}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_67 = {{8{_T_54673[5]}},_T_54673}; // @[Modules.scala 112:22:@8.4]
  assign _T_56406 = $signed(buffer_0_66) + $signed(buffer_0_67); // @[Modules.scala 160:64:@1949.4]
  assign _T_56407 = _T_56406[13:0]; // @[Modules.scala 160:64:@1950.4]
  assign buffer_0_335 = $signed(_T_56407); // @[Modules.scala 160:64:@1951.4]
  assign buffer_0_68 = {{8{_T_54680[5]}},_T_54680}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_69 = {{8{_T_54687[5]}},_T_54687}; // @[Modules.scala 112:22:@8.4]
  assign _T_56409 = $signed(buffer_0_68) + $signed(buffer_0_69); // @[Modules.scala 160:64:@1953.4]
  assign _T_56410 = _T_56409[13:0]; // @[Modules.scala 160:64:@1954.4]
  assign buffer_0_336 = $signed(_T_56410); // @[Modules.scala 160:64:@1955.4]
  assign buffer_0_70 = {{8{_T_54694[5]}},_T_54694}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_71 = {{9{_T_54701[4]}},_T_54701}; // @[Modules.scala 112:22:@8.4]
  assign _T_56412 = $signed(buffer_0_70) + $signed(buffer_0_71); // @[Modules.scala 160:64:@1957.4]
  assign _T_56413 = _T_56412[13:0]; // @[Modules.scala 160:64:@1958.4]
  assign buffer_0_337 = $signed(_T_56413); // @[Modules.scala 160:64:@1959.4]
  assign buffer_0_72 = {{9{_T_54708[4]}},_T_54708}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_73 = {{9{_T_54715[4]}},_T_54715}; // @[Modules.scala 112:22:@8.4]
  assign _T_56415 = $signed(buffer_0_72) + $signed(buffer_0_73); // @[Modules.scala 160:64:@1961.4]
  assign _T_56416 = _T_56415[13:0]; // @[Modules.scala 160:64:@1962.4]
  assign buffer_0_338 = $signed(_T_56416); // @[Modules.scala 160:64:@1963.4]
  assign buffer_0_74 = {{9{_T_54722[4]}},_T_54722}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_75 = {{8{_T_54729[5]}},_T_54729}; // @[Modules.scala 112:22:@8.4]
  assign _T_56418 = $signed(buffer_0_74) + $signed(buffer_0_75); // @[Modules.scala 160:64:@1965.4]
  assign _T_56419 = _T_56418[13:0]; // @[Modules.scala 160:64:@1966.4]
  assign buffer_0_339 = $signed(_T_56419); // @[Modules.scala 160:64:@1967.4]
  assign buffer_0_76 = {{8{_T_54736[5]}},_T_54736}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_77 = {{8{_T_54743[5]}},_T_54743}; // @[Modules.scala 112:22:@8.4]
  assign _T_56421 = $signed(buffer_0_76) + $signed(buffer_0_77); // @[Modules.scala 160:64:@1969.4]
  assign _T_56422 = _T_56421[13:0]; // @[Modules.scala 160:64:@1970.4]
  assign buffer_0_340 = $signed(_T_56422); // @[Modules.scala 160:64:@1971.4]
  assign buffer_0_78 = {{8{_T_54750[5]}},_T_54750}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_79 = {{8{_T_54757[5]}},_T_54757}; // @[Modules.scala 112:22:@8.4]
  assign _T_56424 = $signed(buffer_0_78) + $signed(buffer_0_79); // @[Modules.scala 160:64:@1973.4]
  assign _T_56425 = _T_56424[13:0]; // @[Modules.scala 160:64:@1974.4]
  assign buffer_0_341 = $signed(_T_56425); // @[Modules.scala 160:64:@1975.4]
  assign buffer_0_80 = {{8{_T_54764[5]}},_T_54764}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_81 = {{8{_T_54771[5]}},_T_54771}; // @[Modules.scala 112:22:@8.4]
  assign _T_56427 = $signed(buffer_0_80) + $signed(buffer_0_81); // @[Modules.scala 160:64:@1977.4]
  assign _T_56428 = _T_56427[13:0]; // @[Modules.scala 160:64:@1978.4]
  assign buffer_0_342 = $signed(_T_56428); // @[Modules.scala 160:64:@1979.4]
  assign buffer_0_82 = {{9{_T_54778[4]}},_T_54778}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_83 = {{9{_T_54785[4]}},_T_54785}; // @[Modules.scala 112:22:@8.4]
  assign _T_56430 = $signed(buffer_0_82) + $signed(buffer_0_83); // @[Modules.scala 160:64:@1981.4]
  assign _T_56431 = _T_56430[13:0]; // @[Modules.scala 160:64:@1982.4]
  assign buffer_0_343 = $signed(_T_56431); // @[Modules.scala 160:64:@1983.4]
  assign buffer_0_84 = {{9{_T_54792[4]}},_T_54792}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_85 = {{9{_T_54799[4]}},_T_54799}; // @[Modules.scala 112:22:@8.4]
  assign _T_56433 = $signed(buffer_0_84) + $signed(buffer_0_85); // @[Modules.scala 160:64:@1985.4]
  assign _T_56434 = _T_56433[13:0]; // @[Modules.scala 160:64:@1986.4]
  assign buffer_0_344 = $signed(_T_56434); // @[Modules.scala 160:64:@1987.4]
  assign buffer_0_86 = {{9{_T_54806[4]}},_T_54806}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_87 = {{8{_T_54813[5]}},_T_54813}; // @[Modules.scala 112:22:@8.4]
  assign _T_56436 = $signed(buffer_0_86) + $signed(buffer_0_87); // @[Modules.scala 160:64:@1989.4]
  assign _T_56437 = _T_56436[13:0]; // @[Modules.scala 160:64:@1990.4]
  assign buffer_0_345 = $signed(_T_56437); // @[Modules.scala 160:64:@1991.4]
  assign buffer_0_88 = {{8{_T_54820[5]}},_T_54820}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_89 = {{8{_T_54827[5]}},_T_54827}; // @[Modules.scala 112:22:@8.4]
  assign _T_56439 = $signed(buffer_0_88) + $signed(buffer_0_89); // @[Modules.scala 160:64:@1993.4]
  assign _T_56440 = _T_56439[13:0]; // @[Modules.scala 160:64:@1994.4]
  assign buffer_0_346 = $signed(_T_56440); // @[Modules.scala 160:64:@1995.4]
  assign buffer_0_90 = {{9{_T_54834[4]}},_T_54834}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_91 = {{9{_T_54841[4]}},_T_54841}; // @[Modules.scala 112:22:@8.4]
  assign _T_56442 = $signed(buffer_0_90) + $signed(buffer_0_91); // @[Modules.scala 160:64:@1997.4]
  assign _T_56443 = _T_56442[13:0]; // @[Modules.scala 160:64:@1998.4]
  assign buffer_0_347 = $signed(_T_56443); // @[Modules.scala 160:64:@1999.4]
  assign buffer_0_92 = {{8{_T_54848[5]}},_T_54848}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_93 = {{8{_T_54855[5]}},_T_54855}; // @[Modules.scala 112:22:@8.4]
  assign _T_56445 = $signed(buffer_0_92) + $signed(buffer_0_93); // @[Modules.scala 160:64:@2001.4]
  assign _T_56446 = _T_56445[13:0]; // @[Modules.scala 160:64:@2002.4]
  assign buffer_0_348 = $signed(_T_56446); // @[Modules.scala 160:64:@2003.4]
  assign buffer_0_94 = {{9{_T_54862[4]}},_T_54862}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_95 = {{9{_T_54869[4]}},_T_54869}; // @[Modules.scala 112:22:@8.4]
  assign _T_56448 = $signed(buffer_0_94) + $signed(buffer_0_95); // @[Modules.scala 160:64:@2005.4]
  assign _T_56449 = _T_56448[13:0]; // @[Modules.scala 160:64:@2006.4]
  assign buffer_0_349 = $signed(_T_56449); // @[Modules.scala 160:64:@2007.4]
  assign buffer_0_96 = {{9{_T_54876[4]}},_T_54876}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_97 = {{9{_T_54883[4]}},_T_54883}; // @[Modules.scala 112:22:@8.4]
  assign _T_56451 = $signed(buffer_0_96) + $signed(buffer_0_97); // @[Modules.scala 160:64:@2009.4]
  assign _T_56452 = _T_56451[13:0]; // @[Modules.scala 160:64:@2010.4]
  assign buffer_0_350 = $signed(_T_56452); // @[Modules.scala 160:64:@2011.4]
  assign buffer_0_98 = {{9{_T_54890[4]}},_T_54890}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_99 = {{9{_T_54897[4]}},_T_54897}; // @[Modules.scala 112:22:@8.4]
  assign _T_56454 = $signed(buffer_0_98) + $signed(buffer_0_99); // @[Modules.scala 160:64:@2013.4]
  assign _T_56455 = _T_56454[13:0]; // @[Modules.scala 160:64:@2014.4]
  assign buffer_0_351 = $signed(_T_56455); // @[Modules.scala 160:64:@2015.4]
  assign buffer_0_100 = {{8{_T_54904[5]}},_T_54904}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_101 = {{8{_T_54911[5]}},_T_54911}; // @[Modules.scala 112:22:@8.4]
  assign _T_56457 = $signed(buffer_0_100) + $signed(buffer_0_101); // @[Modules.scala 160:64:@2017.4]
  assign _T_56458 = _T_56457[13:0]; // @[Modules.scala 160:64:@2018.4]
  assign buffer_0_352 = $signed(_T_56458); // @[Modules.scala 160:64:@2019.4]
  assign buffer_0_102 = {{9{_T_54918[4]}},_T_54918}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_103 = {{9{_T_54925[4]}},_T_54925}; // @[Modules.scala 112:22:@8.4]
  assign _T_56460 = $signed(buffer_0_102) + $signed(buffer_0_103); // @[Modules.scala 160:64:@2021.4]
  assign _T_56461 = _T_56460[13:0]; // @[Modules.scala 160:64:@2022.4]
  assign buffer_0_353 = $signed(_T_56461); // @[Modules.scala 160:64:@2023.4]
  assign buffer_0_104 = {{9{_T_54932[4]}},_T_54932}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_105 = {{9{_T_54939[4]}},_T_54939}; // @[Modules.scala 112:22:@8.4]
  assign _T_56463 = $signed(buffer_0_104) + $signed(buffer_0_105); // @[Modules.scala 160:64:@2025.4]
  assign _T_56464 = _T_56463[13:0]; // @[Modules.scala 160:64:@2026.4]
  assign buffer_0_354 = $signed(_T_56464); // @[Modules.scala 160:64:@2027.4]
  assign buffer_0_106 = {{8{_T_54946[5]}},_T_54946}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_107 = {{8{_T_54953[5]}},_T_54953}; // @[Modules.scala 112:22:@8.4]
  assign _T_56466 = $signed(buffer_0_106) + $signed(buffer_0_107); // @[Modules.scala 160:64:@2029.4]
  assign _T_56467 = _T_56466[13:0]; // @[Modules.scala 160:64:@2030.4]
  assign buffer_0_355 = $signed(_T_56467); // @[Modules.scala 160:64:@2031.4]
  assign buffer_0_108 = {{9{_T_54960[4]}},_T_54960}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_109 = {{9{_T_54967[4]}},_T_54967}; // @[Modules.scala 112:22:@8.4]
  assign _T_56469 = $signed(buffer_0_108) + $signed(buffer_0_109); // @[Modules.scala 160:64:@2033.4]
  assign _T_56470 = _T_56469[13:0]; // @[Modules.scala 160:64:@2034.4]
  assign buffer_0_356 = $signed(_T_56470); // @[Modules.scala 160:64:@2035.4]
  assign buffer_0_110 = {{9{_T_54974[4]}},_T_54974}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_111 = {{9{_T_54981[4]}},_T_54981}; // @[Modules.scala 112:22:@8.4]
  assign _T_56472 = $signed(buffer_0_110) + $signed(buffer_0_111); // @[Modules.scala 160:64:@2037.4]
  assign _T_56473 = _T_56472[13:0]; // @[Modules.scala 160:64:@2038.4]
  assign buffer_0_357 = $signed(_T_56473); // @[Modules.scala 160:64:@2039.4]
  assign buffer_0_112 = {{9{_T_54988[4]}},_T_54988}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_113 = {{8{_T_54995[5]}},_T_54995}; // @[Modules.scala 112:22:@8.4]
  assign _T_56475 = $signed(buffer_0_112) + $signed(buffer_0_113); // @[Modules.scala 160:64:@2041.4]
  assign _T_56476 = _T_56475[13:0]; // @[Modules.scala 160:64:@2042.4]
  assign buffer_0_358 = $signed(_T_56476); // @[Modules.scala 160:64:@2043.4]
  assign buffer_0_114 = {{8{_T_55002[5]}},_T_55002}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_115 = {{9{_T_55009[4]}},_T_55009}; // @[Modules.scala 112:22:@8.4]
  assign _T_56478 = $signed(buffer_0_114) + $signed(buffer_0_115); // @[Modules.scala 160:64:@2045.4]
  assign _T_56479 = _T_56478[13:0]; // @[Modules.scala 160:64:@2046.4]
  assign buffer_0_359 = $signed(_T_56479); // @[Modules.scala 160:64:@2047.4]
  assign buffer_0_116 = {{9{_T_55016[4]}},_T_55016}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_117 = {{9{_T_55023[4]}},_T_55023}; // @[Modules.scala 112:22:@8.4]
  assign _T_56481 = $signed(buffer_0_116) + $signed(buffer_0_117); // @[Modules.scala 160:64:@2049.4]
  assign _T_56482 = _T_56481[13:0]; // @[Modules.scala 160:64:@2050.4]
  assign buffer_0_360 = $signed(_T_56482); // @[Modules.scala 160:64:@2051.4]
  assign buffer_0_118 = {{9{_T_55030[4]}},_T_55030}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_119 = {{8{_T_55037[5]}},_T_55037}; // @[Modules.scala 112:22:@8.4]
  assign _T_56484 = $signed(buffer_0_118) + $signed(buffer_0_119); // @[Modules.scala 160:64:@2053.4]
  assign _T_56485 = _T_56484[13:0]; // @[Modules.scala 160:64:@2054.4]
  assign buffer_0_361 = $signed(_T_56485); // @[Modules.scala 160:64:@2055.4]
  assign buffer_0_120 = {{9{_T_55044[4]}},_T_55044}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_121 = {{9{_T_55051[4]}},_T_55051}; // @[Modules.scala 112:22:@8.4]
  assign _T_56487 = $signed(buffer_0_120) + $signed(buffer_0_121); // @[Modules.scala 160:64:@2057.4]
  assign _T_56488 = _T_56487[13:0]; // @[Modules.scala 160:64:@2058.4]
  assign buffer_0_362 = $signed(_T_56488); // @[Modules.scala 160:64:@2059.4]
  assign buffer_0_122 = {{9{_T_55058[4]}},_T_55058}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_123 = {{9{_T_55065[4]}},_T_55065}; // @[Modules.scala 112:22:@8.4]
  assign _T_56490 = $signed(buffer_0_122) + $signed(buffer_0_123); // @[Modules.scala 160:64:@2061.4]
  assign _T_56491 = _T_56490[13:0]; // @[Modules.scala 160:64:@2062.4]
  assign buffer_0_363 = $signed(_T_56491); // @[Modules.scala 160:64:@2063.4]
  assign buffer_0_124 = {{9{_T_55072[4]}},_T_55072}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_125 = {{8{_T_55079[5]}},_T_55079}; // @[Modules.scala 112:22:@8.4]
  assign _T_56493 = $signed(buffer_0_124) + $signed(buffer_0_125); // @[Modules.scala 160:64:@2065.4]
  assign _T_56494 = _T_56493[13:0]; // @[Modules.scala 160:64:@2066.4]
  assign buffer_0_364 = $signed(_T_56494); // @[Modules.scala 160:64:@2067.4]
  assign buffer_0_126 = {{8{_T_55086[5]}},_T_55086}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_127 = {{9{_T_55093[4]}},_T_55093}; // @[Modules.scala 112:22:@8.4]
  assign _T_56496 = $signed(buffer_0_126) + $signed(buffer_0_127); // @[Modules.scala 160:64:@2069.4]
  assign _T_56497 = _T_56496[13:0]; // @[Modules.scala 160:64:@2070.4]
  assign buffer_0_365 = $signed(_T_56497); // @[Modules.scala 160:64:@2071.4]
  assign buffer_0_128 = {{9{_T_55100[4]}},_T_55100}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_129 = {{9{_T_55107[4]}},_T_55107}; // @[Modules.scala 112:22:@8.4]
  assign _T_56499 = $signed(buffer_0_128) + $signed(buffer_0_129); // @[Modules.scala 160:64:@2073.4]
  assign _T_56500 = _T_56499[13:0]; // @[Modules.scala 160:64:@2074.4]
  assign buffer_0_366 = $signed(_T_56500); // @[Modules.scala 160:64:@2075.4]
  assign buffer_0_130 = {{9{_T_55114[4]}},_T_55114}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_131 = {{9{_T_55121[4]}},_T_55121}; // @[Modules.scala 112:22:@8.4]
  assign _T_56502 = $signed(buffer_0_130) + $signed(buffer_0_131); // @[Modules.scala 160:64:@2077.4]
  assign _T_56503 = _T_56502[13:0]; // @[Modules.scala 160:64:@2078.4]
  assign buffer_0_367 = $signed(_T_56503); // @[Modules.scala 160:64:@2079.4]
  assign buffer_0_132 = {{8{_T_55128[5]}},_T_55128}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_133 = {{9{_T_55135[4]}},_T_55135}; // @[Modules.scala 112:22:@8.4]
  assign _T_56505 = $signed(buffer_0_132) + $signed(buffer_0_133); // @[Modules.scala 160:64:@2081.4]
  assign _T_56506 = _T_56505[13:0]; // @[Modules.scala 160:64:@2082.4]
  assign buffer_0_368 = $signed(_T_56506); // @[Modules.scala 160:64:@2083.4]
  assign buffer_0_134 = {{8{_T_55142[5]}},_T_55142}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_135 = {{9{_T_55149[4]}},_T_55149}; // @[Modules.scala 112:22:@8.4]
  assign _T_56508 = $signed(buffer_0_134) + $signed(buffer_0_135); // @[Modules.scala 160:64:@2085.4]
  assign _T_56509 = _T_56508[13:0]; // @[Modules.scala 160:64:@2086.4]
  assign buffer_0_369 = $signed(_T_56509); // @[Modules.scala 160:64:@2087.4]
  assign buffer_0_136 = {{8{_T_55156[5]}},_T_55156}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_137 = {{8{_T_55163[5]}},_T_55163}; // @[Modules.scala 112:22:@8.4]
  assign _T_56511 = $signed(buffer_0_136) + $signed(buffer_0_137); // @[Modules.scala 160:64:@2089.4]
  assign _T_56512 = _T_56511[13:0]; // @[Modules.scala 160:64:@2090.4]
  assign buffer_0_370 = $signed(_T_56512); // @[Modules.scala 160:64:@2091.4]
  assign buffer_0_138 = {{8{_T_55170[5]}},_T_55170}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_139 = {{8{_T_55177[5]}},_T_55177}; // @[Modules.scala 112:22:@8.4]
  assign _T_56514 = $signed(buffer_0_138) + $signed(buffer_0_139); // @[Modules.scala 160:64:@2093.4]
  assign _T_56515 = _T_56514[13:0]; // @[Modules.scala 160:64:@2094.4]
  assign buffer_0_371 = $signed(_T_56515); // @[Modules.scala 160:64:@2095.4]
  assign buffer_0_140 = {{9{_T_55184[4]}},_T_55184}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_141 = {{9{_T_55191[4]}},_T_55191}; // @[Modules.scala 112:22:@8.4]
  assign _T_56517 = $signed(buffer_0_140) + $signed(buffer_0_141); // @[Modules.scala 160:64:@2097.4]
  assign _T_56518 = _T_56517[13:0]; // @[Modules.scala 160:64:@2098.4]
  assign buffer_0_372 = $signed(_T_56518); // @[Modules.scala 160:64:@2099.4]
  assign buffer_0_142 = {{9{_T_55198[4]}},_T_55198}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_143 = {{9{_T_55205[4]}},_T_55205}; // @[Modules.scala 112:22:@8.4]
  assign _T_56520 = $signed(buffer_0_142) + $signed(buffer_0_143); // @[Modules.scala 160:64:@2101.4]
  assign _T_56521 = _T_56520[13:0]; // @[Modules.scala 160:64:@2102.4]
  assign buffer_0_373 = $signed(_T_56521); // @[Modules.scala 160:64:@2103.4]
  assign buffer_0_144 = {{9{_T_55212[4]}},_T_55212}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_145 = {{8{_T_55219[5]}},_T_55219}; // @[Modules.scala 112:22:@8.4]
  assign _T_56523 = $signed(buffer_0_144) + $signed(buffer_0_145); // @[Modules.scala 160:64:@2105.4]
  assign _T_56524 = _T_56523[13:0]; // @[Modules.scala 160:64:@2106.4]
  assign buffer_0_374 = $signed(_T_56524); // @[Modules.scala 160:64:@2107.4]
  assign buffer_0_146 = {{8{_T_55226[5]}},_T_55226}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_147 = {{8{_T_55233[5]}},_T_55233}; // @[Modules.scala 112:22:@8.4]
  assign _T_56526 = $signed(buffer_0_146) + $signed(buffer_0_147); // @[Modules.scala 160:64:@2109.4]
  assign _T_56527 = _T_56526[13:0]; // @[Modules.scala 160:64:@2110.4]
  assign buffer_0_375 = $signed(_T_56527); // @[Modules.scala 160:64:@2111.4]
  assign buffer_0_148 = {{8{_T_55240[5]}},_T_55240}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_149 = {{8{_T_55247[5]}},_T_55247}; // @[Modules.scala 112:22:@8.4]
  assign _T_56529 = $signed(buffer_0_148) + $signed(buffer_0_149); // @[Modules.scala 160:64:@2113.4]
  assign _T_56530 = _T_56529[13:0]; // @[Modules.scala 160:64:@2114.4]
  assign buffer_0_376 = $signed(_T_56530); // @[Modules.scala 160:64:@2115.4]
  assign buffer_0_150 = {{8{_T_55254[5]}},_T_55254}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_151 = {{8{_T_55261[5]}},_T_55261}; // @[Modules.scala 112:22:@8.4]
  assign _T_56532 = $signed(buffer_0_150) + $signed(buffer_0_151); // @[Modules.scala 160:64:@2117.4]
  assign _T_56533 = _T_56532[13:0]; // @[Modules.scala 160:64:@2118.4]
  assign buffer_0_377 = $signed(_T_56533); // @[Modules.scala 160:64:@2119.4]
  assign buffer_0_152 = {{9{_T_55268[4]}},_T_55268}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_153 = {{9{_T_55275[4]}},_T_55275}; // @[Modules.scala 112:22:@8.4]
  assign _T_56535 = $signed(buffer_0_152) + $signed(buffer_0_153); // @[Modules.scala 160:64:@2121.4]
  assign _T_56536 = _T_56535[13:0]; // @[Modules.scala 160:64:@2122.4]
  assign buffer_0_378 = $signed(_T_56536); // @[Modules.scala 160:64:@2123.4]
  assign buffer_0_154 = {{9{_T_55282[4]}},_T_55282}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_155 = {{9{_T_55289[4]}},_T_55289}; // @[Modules.scala 112:22:@8.4]
  assign _T_56538 = $signed(buffer_0_154) + $signed(buffer_0_155); // @[Modules.scala 160:64:@2125.4]
  assign _T_56539 = _T_56538[13:0]; // @[Modules.scala 160:64:@2126.4]
  assign buffer_0_379 = $signed(_T_56539); // @[Modules.scala 160:64:@2127.4]
  assign buffer_0_156 = {{8{_T_55296[5]}},_T_55296}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_157 = {{8{_T_55303[5]}},_T_55303}; // @[Modules.scala 112:22:@8.4]
  assign _T_56541 = $signed(buffer_0_156) + $signed(buffer_0_157); // @[Modules.scala 160:64:@2129.4]
  assign _T_56542 = _T_56541[13:0]; // @[Modules.scala 160:64:@2130.4]
  assign buffer_0_380 = $signed(_T_56542); // @[Modules.scala 160:64:@2131.4]
  assign buffer_0_158 = {{8{_T_55310[5]}},_T_55310}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_159 = {{8{_T_55317[5]}},_T_55317}; // @[Modules.scala 112:22:@8.4]
  assign _T_56544 = $signed(buffer_0_158) + $signed(buffer_0_159); // @[Modules.scala 160:64:@2133.4]
  assign _T_56545 = _T_56544[13:0]; // @[Modules.scala 160:64:@2134.4]
  assign buffer_0_381 = $signed(_T_56545); // @[Modules.scala 160:64:@2135.4]
  assign buffer_0_160 = {{8{_T_55324[5]}},_T_55324}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_161 = {{8{_T_55331[5]}},_T_55331}; // @[Modules.scala 112:22:@8.4]
  assign _T_56547 = $signed(buffer_0_160) + $signed(buffer_0_161); // @[Modules.scala 160:64:@2137.4]
  assign _T_56548 = _T_56547[13:0]; // @[Modules.scala 160:64:@2138.4]
  assign buffer_0_382 = $signed(_T_56548); // @[Modules.scala 160:64:@2139.4]
  assign buffer_0_162 = {{8{_T_55338[5]}},_T_55338}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_163 = {{8{_T_55345[5]}},_T_55345}; // @[Modules.scala 112:22:@8.4]
  assign _T_56550 = $signed(buffer_0_162) + $signed(buffer_0_163); // @[Modules.scala 160:64:@2141.4]
  assign _T_56551 = _T_56550[13:0]; // @[Modules.scala 160:64:@2142.4]
  assign buffer_0_383 = $signed(_T_56551); // @[Modules.scala 160:64:@2143.4]
  assign buffer_0_164 = {{9{_T_55352[4]}},_T_55352}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_165 = {{9{_T_55359[4]}},_T_55359}; // @[Modules.scala 112:22:@8.4]
  assign _T_56553 = $signed(buffer_0_164) + $signed(buffer_0_165); // @[Modules.scala 160:64:@2145.4]
  assign _T_56554 = _T_56553[13:0]; // @[Modules.scala 160:64:@2146.4]
  assign buffer_0_384 = $signed(_T_56554); // @[Modules.scala 160:64:@2147.4]
  assign buffer_0_166 = {{8{_T_55366[5]}},_T_55366}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_167 = {{8{_T_55373[5]}},_T_55373}; // @[Modules.scala 112:22:@8.4]
  assign _T_56556 = $signed(buffer_0_166) + $signed(buffer_0_167); // @[Modules.scala 160:64:@2149.4]
  assign _T_56557 = _T_56556[13:0]; // @[Modules.scala 160:64:@2150.4]
  assign buffer_0_385 = $signed(_T_56557); // @[Modules.scala 160:64:@2151.4]
  assign buffer_0_168 = {{8{_T_55380[5]}},_T_55380}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_169 = {{8{_T_55387[5]}},_T_55387}; // @[Modules.scala 112:22:@8.4]
  assign _T_56559 = $signed(buffer_0_168) + $signed(buffer_0_169); // @[Modules.scala 160:64:@2153.4]
  assign _T_56560 = _T_56559[13:0]; // @[Modules.scala 160:64:@2154.4]
  assign buffer_0_386 = $signed(_T_56560); // @[Modules.scala 160:64:@2155.4]
  assign buffer_0_170 = {{8{_T_55394[5]}},_T_55394}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_171 = {{8{_T_55401[5]}},_T_55401}; // @[Modules.scala 112:22:@8.4]
  assign _T_56562 = $signed(buffer_0_170) + $signed(buffer_0_171); // @[Modules.scala 160:64:@2157.4]
  assign _T_56563 = _T_56562[13:0]; // @[Modules.scala 160:64:@2158.4]
  assign buffer_0_387 = $signed(_T_56563); // @[Modules.scala 160:64:@2159.4]
  assign buffer_0_172 = {{8{_T_55408[5]}},_T_55408}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_173 = {{8{_T_55415[5]}},_T_55415}; // @[Modules.scala 112:22:@8.4]
  assign _T_56565 = $signed(buffer_0_172) + $signed(buffer_0_173); // @[Modules.scala 160:64:@2161.4]
  assign _T_56566 = _T_56565[13:0]; // @[Modules.scala 160:64:@2162.4]
  assign buffer_0_388 = $signed(_T_56566); // @[Modules.scala 160:64:@2163.4]
  assign buffer_0_174 = {{9{_T_55422[4]}},_T_55422}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_175 = {{8{_T_55429[5]}},_T_55429}; // @[Modules.scala 112:22:@8.4]
  assign _T_56568 = $signed(buffer_0_174) + $signed(buffer_0_175); // @[Modules.scala 160:64:@2165.4]
  assign _T_56569 = _T_56568[13:0]; // @[Modules.scala 160:64:@2166.4]
  assign buffer_0_389 = $signed(_T_56569); // @[Modules.scala 160:64:@2167.4]
  assign buffer_0_176 = {{9{_T_55436[4]}},_T_55436}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_177 = {{8{_T_55443[5]}},_T_55443}; // @[Modules.scala 112:22:@8.4]
  assign _T_56571 = $signed(buffer_0_176) + $signed(buffer_0_177); // @[Modules.scala 160:64:@2169.4]
  assign _T_56572 = _T_56571[13:0]; // @[Modules.scala 160:64:@2170.4]
  assign buffer_0_390 = $signed(_T_56572); // @[Modules.scala 160:64:@2171.4]
  assign buffer_0_178 = {{8{_T_55450[5]}},_T_55450}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_179 = {{8{_T_55457[5]}},_T_55457}; // @[Modules.scala 112:22:@8.4]
  assign _T_56574 = $signed(buffer_0_178) + $signed(buffer_0_179); // @[Modules.scala 160:64:@2173.4]
  assign _T_56575 = _T_56574[13:0]; // @[Modules.scala 160:64:@2174.4]
  assign buffer_0_391 = $signed(_T_56575); // @[Modules.scala 160:64:@2175.4]
  assign buffer_0_180 = {{8{_T_55464[5]}},_T_55464}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_181 = {{8{_T_55471[5]}},_T_55471}; // @[Modules.scala 112:22:@8.4]
  assign _T_56577 = $signed(buffer_0_180) + $signed(buffer_0_181); // @[Modules.scala 160:64:@2177.4]
  assign _T_56578 = _T_56577[13:0]; // @[Modules.scala 160:64:@2178.4]
  assign buffer_0_392 = $signed(_T_56578); // @[Modules.scala 160:64:@2179.4]
  assign buffer_0_182 = {{8{_T_55478[5]}},_T_55478}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_183 = {{8{_T_55485[5]}},_T_55485}; // @[Modules.scala 112:22:@8.4]
  assign _T_56580 = $signed(buffer_0_182) + $signed(buffer_0_183); // @[Modules.scala 160:64:@2181.4]
  assign _T_56581 = _T_56580[13:0]; // @[Modules.scala 160:64:@2182.4]
  assign buffer_0_393 = $signed(_T_56581); // @[Modules.scala 160:64:@2183.4]
  assign buffer_0_184 = {{8{_T_55492[5]}},_T_55492}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_185 = {{8{_T_55499[5]}},_T_55499}; // @[Modules.scala 112:22:@8.4]
  assign _T_56583 = $signed(buffer_0_184) + $signed(buffer_0_185); // @[Modules.scala 160:64:@2185.4]
  assign _T_56584 = _T_56583[13:0]; // @[Modules.scala 160:64:@2186.4]
  assign buffer_0_394 = $signed(_T_56584); // @[Modules.scala 160:64:@2187.4]
  assign buffer_0_186 = {{8{_T_55506[5]}},_T_55506}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_187 = {{8{_T_55513[5]}},_T_55513}; // @[Modules.scala 112:22:@8.4]
  assign _T_56586 = $signed(buffer_0_186) + $signed(buffer_0_187); // @[Modules.scala 160:64:@2189.4]
  assign _T_56587 = _T_56586[13:0]; // @[Modules.scala 160:64:@2190.4]
  assign buffer_0_395 = $signed(_T_56587); // @[Modules.scala 160:64:@2191.4]
  assign buffer_0_188 = {{8{_T_55520[5]}},_T_55520}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_189 = {{8{_T_55527[5]}},_T_55527}; // @[Modules.scala 112:22:@8.4]
  assign _T_56589 = $signed(buffer_0_188) + $signed(buffer_0_189); // @[Modules.scala 160:64:@2193.4]
  assign _T_56590 = _T_56589[13:0]; // @[Modules.scala 160:64:@2194.4]
  assign buffer_0_396 = $signed(_T_56590); // @[Modules.scala 160:64:@2195.4]
  assign buffer_0_190 = {{9{_T_55534[4]}},_T_55534}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_191 = {{8{_T_55541[5]}},_T_55541}; // @[Modules.scala 112:22:@8.4]
  assign _T_56592 = $signed(buffer_0_190) + $signed(buffer_0_191); // @[Modules.scala 160:64:@2197.4]
  assign _T_56593 = _T_56592[13:0]; // @[Modules.scala 160:64:@2198.4]
  assign buffer_0_397 = $signed(_T_56593); // @[Modules.scala 160:64:@2199.4]
  assign buffer_0_192 = {{8{_T_55548[5]}},_T_55548}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_193 = {{8{_T_55555[5]}},_T_55555}; // @[Modules.scala 112:22:@8.4]
  assign _T_56595 = $signed(buffer_0_192) + $signed(buffer_0_193); // @[Modules.scala 160:64:@2201.4]
  assign _T_56596 = _T_56595[13:0]; // @[Modules.scala 160:64:@2202.4]
  assign buffer_0_398 = $signed(_T_56596); // @[Modules.scala 160:64:@2203.4]
  assign buffer_0_194 = {{8{_T_55562[5]}},_T_55562}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_195 = {{8{_T_55569[5]}},_T_55569}; // @[Modules.scala 112:22:@8.4]
  assign _T_56598 = $signed(buffer_0_194) + $signed(buffer_0_195); // @[Modules.scala 160:64:@2205.4]
  assign _T_56599 = _T_56598[13:0]; // @[Modules.scala 160:64:@2206.4]
  assign buffer_0_399 = $signed(_T_56599); // @[Modules.scala 160:64:@2207.4]
  assign buffer_0_196 = {{8{_T_55576[5]}},_T_55576}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_197 = {{8{_T_55583[5]}},_T_55583}; // @[Modules.scala 112:22:@8.4]
  assign _T_56601 = $signed(buffer_0_196) + $signed(buffer_0_197); // @[Modules.scala 160:64:@2209.4]
  assign _T_56602 = _T_56601[13:0]; // @[Modules.scala 160:64:@2210.4]
  assign buffer_0_400 = $signed(_T_56602); // @[Modules.scala 160:64:@2211.4]
  assign buffer_0_198 = {{8{_T_55590[5]}},_T_55590}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_199 = {{8{_T_55597[5]}},_T_55597}; // @[Modules.scala 112:22:@8.4]
  assign _T_56604 = $signed(buffer_0_198) + $signed(buffer_0_199); // @[Modules.scala 160:64:@2213.4]
  assign _T_56605 = _T_56604[13:0]; // @[Modules.scala 160:64:@2214.4]
  assign buffer_0_401 = $signed(_T_56605); // @[Modules.scala 160:64:@2215.4]
  assign buffer_0_200 = {{8{_T_55604[5]}},_T_55604}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_201 = {{8{_T_55611[5]}},_T_55611}; // @[Modules.scala 112:22:@8.4]
  assign _T_56607 = $signed(buffer_0_200) + $signed(buffer_0_201); // @[Modules.scala 160:64:@2217.4]
  assign _T_56608 = _T_56607[13:0]; // @[Modules.scala 160:64:@2218.4]
  assign buffer_0_402 = $signed(_T_56608); // @[Modules.scala 160:64:@2219.4]
  assign buffer_0_202 = {{8{_T_55618[5]}},_T_55618}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_203 = {{8{_T_55625[5]}},_T_55625}; // @[Modules.scala 112:22:@8.4]
  assign _T_56610 = $signed(buffer_0_202) + $signed(buffer_0_203); // @[Modules.scala 160:64:@2221.4]
  assign _T_56611 = _T_56610[13:0]; // @[Modules.scala 160:64:@2222.4]
  assign buffer_0_403 = $signed(_T_56611); // @[Modules.scala 160:64:@2223.4]
  assign buffer_0_204 = {{8{_T_55632[5]}},_T_55632}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_205 = {{8{_T_55639[5]}},_T_55639}; // @[Modules.scala 112:22:@8.4]
  assign _T_56613 = $signed(buffer_0_204) + $signed(buffer_0_205); // @[Modules.scala 160:64:@2225.4]
  assign _T_56614 = _T_56613[13:0]; // @[Modules.scala 160:64:@2226.4]
  assign buffer_0_404 = $signed(_T_56614); // @[Modules.scala 160:64:@2227.4]
  assign buffer_0_206 = {{8{_T_55646[5]}},_T_55646}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_207 = {{8{_T_55653[5]}},_T_55653}; // @[Modules.scala 112:22:@8.4]
  assign _T_56616 = $signed(buffer_0_206) + $signed(buffer_0_207); // @[Modules.scala 160:64:@2229.4]
  assign _T_56617 = _T_56616[13:0]; // @[Modules.scala 160:64:@2230.4]
  assign buffer_0_405 = $signed(_T_56617); // @[Modules.scala 160:64:@2231.4]
  assign buffer_0_208 = {{8{_T_55660[5]}},_T_55660}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_209 = {{8{_T_55667[5]}},_T_55667}; // @[Modules.scala 112:22:@8.4]
  assign _T_56619 = $signed(buffer_0_208) + $signed(buffer_0_209); // @[Modules.scala 160:64:@2233.4]
  assign _T_56620 = _T_56619[13:0]; // @[Modules.scala 160:64:@2234.4]
  assign buffer_0_406 = $signed(_T_56620); // @[Modules.scala 160:64:@2235.4]
  assign buffer_0_210 = {{8{_T_55674[5]}},_T_55674}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_211 = {{8{_T_55681[5]}},_T_55681}; // @[Modules.scala 112:22:@8.4]
  assign _T_56622 = $signed(buffer_0_210) + $signed(buffer_0_211); // @[Modules.scala 160:64:@2237.4]
  assign _T_56623 = _T_56622[13:0]; // @[Modules.scala 160:64:@2238.4]
  assign buffer_0_407 = $signed(_T_56623); // @[Modules.scala 160:64:@2239.4]
  assign buffer_0_212 = {{8{_T_55688[5]}},_T_55688}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_213 = {{8{_T_55695[5]}},_T_55695}; // @[Modules.scala 112:22:@8.4]
  assign _T_56625 = $signed(buffer_0_212) + $signed(buffer_0_213); // @[Modules.scala 160:64:@2241.4]
  assign _T_56626 = _T_56625[13:0]; // @[Modules.scala 160:64:@2242.4]
  assign buffer_0_408 = $signed(_T_56626); // @[Modules.scala 160:64:@2243.4]
  assign buffer_0_214 = {{8{_T_55702[5]}},_T_55702}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_215 = {{8{_T_55709[5]}},_T_55709}; // @[Modules.scala 112:22:@8.4]
  assign _T_56628 = $signed(buffer_0_214) + $signed(buffer_0_215); // @[Modules.scala 160:64:@2245.4]
  assign _T_56629 = _T_56628[13:0]; // @[Modules.scala 160:64:@2246.4]
  assign buffer_0_409 = $signed(_T_56629); // @[Modules.scala 160:64:@2247.4]
  assign buffer_0_216 = {{8{_T_55716[5]}},_T_55716}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_217 = {{8{_T_55723[5]}},_T_55723}; // @[Modules.scala 112:22:@8.4]
  assign _T_56631 = $signed(buffer_0_216) + $signed(buffer_0_217); // @[Modules.scala 160:64:@2249.4]
  assign _T_56632 = _T_56631[13:0]; // @[Modules.scala 160:64:@2250.4]
  assign buffer_0_410 = $signed(_T_56632); // @[Modules.scala 160:64:@2251.4]
  assign buffer_0_218 = {{8{_T_55730[5]}},_T_55730}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_219 = {{8{_T_55737[5]}},_T_55737}; // @[Modules.scala 112:22:@8.4]
  assign _T_56634 = $signed(buffer_0_218) + $signed(buffer_0_219); // @[Modules.scala 160:64:@2253.4]
  assign _T_56635 = _T_56634[13:0]; // @[Modules.scala 160:64:@2254.4]
  assign buffer_0_411 = $signed(_T_56635); // @[Modules.scala 160:64:@2255.4]
  assign buffer_0_220 = {{8{_T_55744[5]}},_T_55744}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_221 = {{8{_T_55751[5]}},_T_55751}; // @[Modules.scala 112:22:@8.4]
  assign _T_56637 = $signed(buffer_0_220) + $signed(buffer_0_221); // @[Modules.scala 160:64:@2257.4]
  assign _T_56638 = _T_56637[13:0]; // @[Modules.scala 160:64:@2258.4]
  assign buffer_0_412 = $signed(_T_56638); // @[Modules.scala 160:64:@2259.4]
  assign buffer_0_222 = {{8{_T_55758[5]}},_T_55758}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_223 = {{8{_T_55765[5]}},_T_55765}; // @[Modules.scala 112:22:@8.4]
  assign _T_56640 = $signed(buffer_0_222) + $signed(buffer_0_223); // @[Modules.scala 160:64:@2261.4]
  assign _T_56641 = _T_56640[13:0]; // @[Modules.scala 160:64:@2262.4]
  assign buffer_0_413 = $signed(_T_56641); // @[Modules.scala 160:64:@2263.4]
  assign buffer_0_224 = {{8{_T_55772[5]}},_T_55772}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_225 = {{8{_T_55779[5]}},_T_55779}; // @[Modules.scala 112:22:@8.4]
  assign _T_56643 = $signed(buffer_0_224) + $signed(buffer_0_225); // @[Modules.scala 160:64:@2265.4]
  assign _T_56644 = _T_56643[13:0]; // @[Modules.scala 160:64:@2266.4]
  assign buffer_0_414 = $signed(_T_56644); // @[Modules.scala 160:64:@2267.4]
  assign buffer_0_226 = {{8{_T_55786[5]}},_T_55786}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_227 = {{8{_T_55793[5]}},_T_55793}; // @[Modules.scala 112:22:@8.4]
  assign _T_56646 = $signed(buffer_0_226) + $signed(buffer_0_227); // @[Modules.scala 160:64:@2269.4]
  assign _T_56647 = _T_56646[13:0]; // @[Modules.scala 160:64:@2270.4]
  assign buffer_0_415 = $signed(_T_56647); // @[Modules.scala 160:64:@2271.4]
  assign buffer_0_228 = {{8{_T_55800[5]}},_T_55800}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_229 = {{8{_T_55807[5]}},_T_55807}; // @[Modules.scala 112:22:@8.4]
  assign _T_56649 = $signed(buffer_0_228) + $signed(buffer_0_229); // @[Modules.scala 160:64:@2273.4]
  assign _T_56650 = _T_56649[13:0]; // @[Modules.scala 160:64:@2274.4]
  assign buffer_0_416 = $signed(_T_56650); // @[Modules.scala 160:64:@2275.4]
  assign buffer_0_230 = {{8{_T_55814[5]}},_T_55814}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_231 = {{8{_T_55821[5]}},_T_55821}; // @[Modules.scala 112:22:@8.4]
  assign _T_56652 = $signed(buffer_0_230) + $signed(buffer_0_231); // @[Modules.scala 160:64:@2277.4]
  assign _T_56653 = _T_56652[13:0]; // @[Modules.scala 160:64:@2278.4]
  assign buffer_0_417 = $signed(_T_56653); // @[Modules.scala 160:64:@2279.4]
  assign buffer_0_232 = {{8{_T_55828[5]}},_T_55828}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_233 = {{8{_T_55835[5]}},_T_55835}; // @[Modules.scala 112:22:@8.4]
  assign _T_56655 = $signed(buffer_0_232) + $signed(buffer_0_233); // @[Modules.scala 160:64:@2281.4]
  assign _T_56656 = _T_56655[13:0]; // @[Modules.scala 160:64:@2282.4]
  assign buffer_0_418 = $signed(_T_56656); // @[Modules.scala 160:64:@2283.4]
  assign buffer_0_234 = {{8{_T_55842[5]}},_T_55842}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_235 = {{8{_T_55849[5]}},_T_55849}; // @[Modules.scala 112:22:@8.4]
  assign _T_56658 = $signed(buffer_0_234) + $signed(buffer_0_235); // @[Modules.scala 160:64:@2285.4]
  assign _T_56659 = _T_56658[13:0]; // @[Modules.scala 160:64:@2286.4]
  assign buffer_0_419 = $signed(_T_56659); // @[Modules.scala 160:64:@2287.4]
  assign buffer_0_236 = {{8{_T_55856[5]}},_T_55856}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_237 = {{8{_T_55863[5]}},_T_55863}; // @[Modules.scala 112:22:@8.4]
  assign _T_56661 = $signed(buffer_0_236) + $signed(buffer_0_237); // @[Modules.scala 160:64:@2289.4]
  assign _T_56662 = _T_56661[13:0]; // @[Modules.scala 160:64:@2290.4]
  assign buffer_0_420 = $signed(_T_56662); // @[Modules.scala 160:64:@2291.4]
  assign buffer_0_238 = {{8{_T_55870[5]}},_T_55870}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_239 = {{8{_T_55877[5]}},_T_55877}; // @[Modules.scala 112:22:@8.4]
  assign _T_56664 = $signed(buffer_0_238) + $signed(buffer_0_239); // @[Modules.scala 160:64:@2293.4]
  assign _T_56665 = _T_56664[13:0]; // @[Modules.scala 160:64:@2294.4]
  assign buffer_0_421 = $signed(_T_56665); // @[Modules.scala 160:64:@2295.4]
  assign buffer_0_240 = {{8{_T_55884[5]}},_T_55884}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_241 = {{8{_T_55891[5]}},_T_55891}; // @[Modules.scala 112:22:@8.4]
  assign _T_56667 = $signed(buffer_0_240) + $signed(buffer_0_241); // @[Modules.scala 160:64:@2297.4]
  assign _T_56668 = _T_56667[13:0]; // @[Modules.scala 160:64:@2298.4]
  assign buffer_0_422 = $signed(_T_56668); // @[Modules.scala 160:64:@2299.4]
  assign buffer_0_242 = {{9{_T_55898[4]}},_T_55898}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_243 = {{9{_T_55905[4]}},_T_55905}; // @[Modules.scala 112:22:@8.4]
  assign _T_56670 = $signed(buffer_0_242) + $signed(buffer_0_243); // @[Modules.scala 160:64:@2301.4]
  assign _T_56671 = _T_56670[13:0]; // @[Modules.scala 160:64:@2302.4]
  assign buffer_0_423 = $signed(_T_56671); // @[Modules.scala 160:64:@2303.4]
  assign buffer_0_244 = {{9{_T_55912[4]}},_T_55912}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_245 = {{9{_T_55919[4]}},_T_55919}; // @[Modules.scala 112:22:@8.4]
  assign _T_56673 = $signed(buffer_0_244) + $signed(buffer_0_245); // @[Modules.scala 160:64:@2305.4]
  assign _T_56674 = _T_56673[13:0]; // @[Modules.scala 160:64:@2306.4]
  assign buffer_0_424 = $signed(_T_56674); // @[Modules.scala 160:64:@2307.4]
  assign buffer_0_246 = {{8{_T_55926[5]}},_T_55926}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_247 = {{8{_T_55933[5]}},_T_55933}; // @[Modules.scala 112:22:@8.4]
  assign _T_56676 = $signed(buffer_0_246) + $signed(buffer_0_247); // @[Modules.scala 160:64:@2309.4]
  assign _T_56677 = _T_56676[13:0]; // @[Modules.scala 160:64:@2310.4]
  assign buffer_0_425 = $signed(_T_56677); // @[Modules.scala 160:64:@2311.4]
  assign buffer_0_248 = {{8{_T_55940[5]}},_T_55940}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_249 = {{8{_T_55947[5]}},_T_55947}; // @[Modules.scala 112:22:@8.4]
  assign _T_56679 = $signed(buffer_0_248) + $signed(buffer_0_249); // @[Modules.scala 160:64:@2313.4]
  assign _T_56680 = _T_56679[13:0]; // @[Modules.scala 160:64:@2314.4]
  assign buffer_0_426 = $signed(_T_56680); // @[Modules.scala 160:64:@2315.4]
  assign buffer_0_250 = {{8{_T_55954[5]}},_T_55954}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_251 = {{8{_T_55961[5]}},_T_55961}; // @[Modules.scala 112:22:@8.4]
  assign _T_56682 = $signed(buffer_0_250) + $signed(buffer_0_251); // @[Modules.scala 160:64:@2317.4]
  assign _T_56683 = _T_56682[13:0]; // @[Modules.scala 160:64:@2318.4]
  assign buffer_0_427 = $signed(_T_56683); // @[Modules.scala 160:64:@2319.4]
  assign buffer_0_252 = {{8{_T_55968[5]}},_T_55968}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_253 = {{9{_T_55975[4]}},_T_55975}; // @[Modules.scala 112:22:@8.4]
  assign _T_56685 = $signed(buffer_0_252) + $signed(buffer_0_253); // @[Modules.scala 160:64:@2321.4]
  assign _T_56686 = _T_56685[13:0]; // @[Modules.scala 160:64:@2322.4]
  assign buffer_0_428 = $signed(_T_56686); // @[Modules.scala 160:64:@2323.4]
  assign buffer_0_254 = {{9{_T_55982[4]}},_T_55982}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_255 = {{9{_T_55989[4]}},_T_55989}; // @[Modules.scala 112:22:@8.4]
  assign _T_56688 = $signed(buffer_0_254) + $signed(buffer_0_255); // @[Modules.scala 160:64:@2325.4]
  assign _T_56689 = _T_56688[13:0]; // @[Modules.scala 160:64:@2326.4]
  assign buffer_0_429 = $signed(_T_56689); // @[Modules.scala 160:64:@2327.4]
  assign buffer_0_256 = {{9{_T_55996[4]}},_T_55996}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_257 = {{9{_T_56003[4]}},_T_56003}; // @[Modules.scala 112:22:@8.4]
  assign _T_56691 = $signed(buffer_0_256) + $signed(buffer_0_257); // @[Modules.scala 160:64:@2329.4]
  assign _T_56692 = _T_56691[13:0]; // @[Modules.scala 160:64:@2330.4]
  assign buffer_0_430 = $signed(_T_56692); // @[Modules.scala 160:64:@2331.4]
  assign buffer_0_258 = {{9{_T_56010[4]}},_T_56010}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_259 = {{9{_T_56017[4]}},_T_56017}; // @[Modules.scala 112:22:@8.4]
  assign _T_56694 = $signed(buffer_0_258) + $signed(buffer_0_259); // @[Modules.scala 160:64:@2333.4]
  assign _T_56695 = _T_56694[13:0]; // @[Modules.scala 160:64:@2334.4]
  assign buffer_0_431 = $signed(_T_56695); // @[Modules.scala 160:64:@2335.4]
  assign buffer_0_260 = {{8{_T_56024[5]}},_T_56024}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_261 = {{8{_T_56031[5]}},_T_56031}; // @[Modules.scala 112:22:@8.4]
  assign _T_56697 = $signed(buffer_0_260) + $signed(buffer_0_261); // @[Modules.scala 160:64:@2337.4]
  assign _T_56698 = _T_56697[13:0]; // @[Modules.scala 160:64:@2338.4]
  assign buffer_0_432 = $signed(_T_56698); // @[Modules.scala 160:64:@2339.4]
  assign buffer_0_262 = {{8{_T_56038[5]}},_T_56038}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_263 = {{8{_T_56045[5]}},_T_56045}; // @[Modules.scala 112:22:@8.4]
  assign _T_56700 = $signed(buffer_0_262) + $signed(buffer_0_263); // @[Modules.scala 160:64:@2341.4]
  assign _T_56701 = _T_56700[13:0]; // @[Modules.scala 160:64:@2342.4]
  assign buffer_0_433 = $signed(_T_56701); // @[Modules.scala 160:64:@2343.4]
  assign buffer_0_264 = {{8{_T_56052[5]}},_T_56052}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_265 = {{9{_T_56059[4]}},_T_56059}; // @[Modules.scala 112:22:@8.4]
  assign _T_56703 = $signed(buffer_0_264) + $signed(buffer_0_265); // @[Modules.scala 160:64:@2345.4]
  assign _T_56704 = _T_56703[13:0]; // @[Modules.scala 160:64:@2346.4]
  assign buffer_0_434 = $signed(_T_56704); // @[Modules.scala 160:64:@2347.4]
  assign buffer_0_266 = {{9{_T_56066[4]}},_T_56066}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_267 = {{9{_T_56073[4]}},_T_56073}; // @[Modules.scala 112:22:@8.4]
  assign _T_56706 = $signed(buffer_0_266) + $signed(buffer_0_267); // @[Modules.scala 160:64:@2349.4]
  assign _T_56707 = _T_56706[13:0]; // @[Modules.scala 160:64:@2350.4]
  assign buffer_0_435 = $signed(_T_56707); // @[Modules.scala 160:64:@2351.4]
  assign buffer_0_268 = {{9{_T_56080[4]}},_T_56080}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_269 = {{9{_T_56087[4]}},_T_56087}; // @[Modules.scala 112:22:@8.4]
  assign _T_56709 = $signed(buffer_0_268) + $signed(buffer_0_269); // @[Modules.scala 160:64:@2353.4]
  assign _T_56710 = _T_56709[13:0]; // @[Modules.scala 160:64:@2354.4]
  assign buffer_0_436 = $signed(_T_56710); // @[Modules.scala 160:64:@2355.4]
  assign buffer_0_270 = {{9{_T_56094[4]}},_T_56094}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_271 = {{8{_T_56101[5]}},_T_56101}; // @[Modules.scala 112:22:@8.4]
  assign _T_56712 = $signed(buffer_0_270) + $signed(buffer_0_271); // @[Modules.scala 160:64:@2357.4]
  assign _T_56713 = _T_56712[13:0]; // @[Modules.scala 160:64:@2358.4]
  assign buffer_0_437 = $signed(_T_56713); // @[Modules.scala 160:64:@2359.4]
  assign buffer_0_272 = {{8{_T_56108[5]}},_T_56108}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_273 = {{8{_T_56115[5]}},_T_56115}; // @[Modules.scala 112:22:@8.4]
  assign _T_56715 = $signed(buffer_0_272) + $signed(buffer_0_273); // @[Modules.scala 160:64:@2361.4]
  assign _T_56716 = _T_56715[13:0]; // @[Modules.scala 160:64:@2362.4]
  assign buffer_0_438 = $signed(_T_56716); // @[Modules.scala 160:64:@2363.4]
  assign buffer_0_274 = {{8{_T_56122[5]}},_T_56122}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_275 = {{8{_T_56129[5]}},_T_56129}; // @[Modules.scala 112:22:@8.4]
  assign _T_56718 = $signed(buffer_0_274) + $signed(buffer_0_275); // @[Modules.scala 160:64:@2365.4]
  assign _T_56719 = _T_56718[13:0]; // @[Modules.scala 160:64:@2366.4]
  assign buffer_0_439 = $signed(_T_56719); // @[Modules.scala 160:64:@2367.4]
  assign buffer_0_276 = {{8{_T_56136[5]}},_T_56136}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_277 = {{8{_T_56143[5]}},_T_56143}; // @[Modules.scala 112:22:@8.4]
  assign _T_56721 = $signed(buffer_0_276) + $signed(buffer_0_277); // @[Modules.scala 160:64:@2369.4]
  assign _T_56722 = _T_56721[13:0]; // @[Modules.scala 160:64:@2370.4]
  assign buffer_0_440 = $signed(_T_56722); // @[Modules.scala 160:64:@2371.4]
  assign buffer_0_278 = {{9{_T_56150[4]}},_T_56150}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_279 = {{9{_T_56157[4]}},_T_56157}; // @[Modules.scala 112:22:@8.4]
  assign _T_56724 = $signed(buffer_0_278) + $signed(buffer_0_279); // @[Modules.scala 160:64:@2373.4]
  assign _T_56725 = _T_56724[13:0]; // @[Modules.scala 160:64:@2374.4]
  assign buffer_0_441 = $signed(_T_56725); // @[Modules.scala 160:64:@2375.4]
  assign buffer_0_280 = {{9{_T_56164[4]}},_T_56164}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_281 = {{9{_T_56171[4]}},_T_56171}; // @[Modules.scala 112:22:@8.4]
  assign _T_56727 = $signed(buffer_0_280) + $signed(buffer_0_281); // @[Modules.scala 160:64:@2377.4]
  assign _T_56728 = _T_56727[13:0]; // @[Modules.scala 160:64:@2378.4]
  assign buffer_0_442 = $signed(_T_56728); // @[Modules.scala 160:64:@2379.4]
  assign buffer_0_282 = {{9{_T_56178[4]}},_T_56178}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_283 = {{9{_T_56185[4]}},_T_56185}; // @[Modules.scala 112:22:@8.4]
  assign _T_56730 = $signed(buffer_0_282) + $signed(buffer_0_283); // @[Modules.scala 160:64:@2381.4]
  assign _T_56731 = _T_56730[13:0]; // @[Modules.scala 160:64:@2382.4]
  assign buffer_0_443 = $signed(_T_56731); // @[Modules.scala 160:64:@2383.4]
  assign buffer_0_284 = {{9{_T_56192[4]}},_T_56192}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_285 = {{8{_T_56199[5]}},_T_56199}; // @[Modules.scala 112:22:@8.4]
  assign _T_56733 = $signed(buffer_0_284) + $signed(buffer_0_285); // @[Modules.scala 160:64:@2385.4]
  assign _T_56734 = _T_56733[13:0]; // @[Modules.scala 160:64:@2386.4]
  assign buffer_0_444 = $signed(_T_56734); // @[Modules.scala 160:64:@2387.4]
  assign buffer_0_286 = {{8{_T_56206[5]}},_T_56206}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_287 = {{8{_T_56213[5]}},_T_56213}; // @[Modules.scala 112:22:@8.4]
  assign _T_56736 = $signed(buffer_0_286) + $signed(buffer_0_287); // @[Modules.scala 160:64:@2389.4]
  assign _T_56737 = _T_56736[13:0]; // @[Modules.scala 160:64:@2390.4]
  assign buffer_0_445 = $signed(_T_56737); // @[Modules.scala 160:64:@2391.4]
  assign buffer_0_288 = {{8{_T_56220[5]}},_T_56220}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_289 = {{8{_T_56227[5]}},_T_56227}; // @[Modules.scala 112:22:@8.4]
  assign _T_56739 = $signed(buffer_0_288) + $signed(buffer_0_289); // @[Modules.scala 160:64:@2393.4]
  assign _T_56740 = _T_56739[13:0]; // @[Modules.scala 160:64:@2394.4]
  assign buffer_0_446 = $signed(_T_56740); // @[Modules.scala 160:64:@2395.4]
  assign buffer_0_290 = {{9{_T_56234[4]}},_T_56234}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_291 = {{9{_T_56241[4]}},_T_56241}; // @[Modules.scala 112:22:@8.4]
  assign _T_56742 = $signed(buffer_0_290) + $signed(buffer_0_291); // @[Modules.scala 160:64:@2397.4]
  assign _T_56743 = _T_56742[13:0]; // @[Modules.scala 160:64:@2398.4]
  assign buffer_0_447 = $signed(_T_56743); // @[Modules.scala 160:64:@2399.4]
  assign buffer_0_292 = {{8{_T_56248[5]}},_T_56248}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_293 = {{8{_T_56255[5]}},_T_56255}; // @[Modules.scala 112:22:@8.4]
  assign _T_56745 = $signed(buffer_0_292) + $signed(buffer_0_293); // @[Modules.scala 160:64:@2401.4]
  assign _T_56746 = _T_56745[13:0]; // @[Modules.scala 160:64:@2402.4]
  assign buffer_0_448 = $signed(_T_56746); // @[Modules.scala 160:64:@2403.4]
  assign buffer_0_294 = {{9{_T_56262[4]}},_T_56262}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_295 = {{8{_T_56269[5]}},_T_56269}; // @[Modules.scala 112:22:@8.4]
  assign _T_56748 = $signed(buffer_0_294) + $signed(buffer_0_295); // @[Modules.scala 160:64:@2405.4]
  assign _T_56749 = _T_56748[13:0]; // @[Modules.scala 160:64:@2406.4]
  assign buffer_0_449 = $signed(_T_56749); // @[Modules.scala 160:64:@2407.4]
  assign buffer_0_296 = {{8{_T_56276[5]}},_T_56276}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_297 = {{8{_T_56283[5]}},_T_56283}; // @[Modules.scala 112:22:@8.4]
  assign _T_56751 = $signed(buffer_0_296) + $signed(buffer_0_297); // @[Modules.scala 160:64:@2409.4]
  assign _T_56752 = _T_56751[13:0]; // @[Modules.scala 160:64:@2410.4]
  assign buffer_0_450 = $signed(_T_56752); // @[Modules.scala 160:64:@2411.4]
  assign buffer_0_298 = {{8{_T_56290[5]}},_T_56290}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_299 = {{9{_T_56297[4]}},_T_56297}; // @[Modules.scala 112:22:@8.4]
  assign _T_56754 = $signed(buffer_0_298) + $signed(buffer_0_299); // @[Modules.scala 160:64:@2413.4]
  assign _T_56755 = _T_56754[13:0]; // @[Modules.scala 160:64:@2414.4]
  assign buffer_0_451 = $signed(_T_56755); // @[Modules.scala 160:64:@2415.4]
  assign buffer_0_300 = {{8{_T_56304[5]}},_T_56304}; // @[Modules.scala 112:22:@8.4]
  assign buffer_0_301 = {{8{_T_56306[5]}},_T_56306}; // @[Modules.scala 112:22:@8.4]
  assign _T_56757 = $signed(buffer_0_300) + $signed(buffer_0_301); // @[Modules.scala 160:64:@2417.4]
  assign _T_56758 = _T_56757[13:0]; // @[Modules.scala 160:64:@2418.4]
  assign buffer_0_452 = $signed(_T_56758); // @[Modules.scala 160:64:@2419.4]
  assign _T_56760 = $signed(buffer_0_302) + $signed(buffer_0_303); // @[Modules.scala 166:64:@2421.4]
  assign _T_56761 = _T_56760[13:0]; // @[Modules.scala 166:64:@2422.4]
  assign buffer_0_453 = $signed(_T_56761); // @[Modules.scala 166:64:@2423.4]
  assign _T_56763 = $signed(buffer_0_304) + $signed(buffer_0_305); // @[Modules.scala 166:64:@2425.4]
  assign _T_56764 = _T_56763[13:0]; // @[Modules.scala 166:64:@2426.4]
  assign buffer_0_454 = $signed(_T_56764); // @[Modules.scala 166:64:@2427.4]
  assign _T_56766 = $signed(buffer_0_306) + $signed(buffer_0_307); // @[Modules.scala 166:64:@2429.4]
  assign _T_56767 = _T_56766[13:0]; // @[Modules.scala 166:64:@2430.4]
  assign buffer_0_455 = $signed(_T_56767); // @[Modules.scala 166:64:@2431.4]
  assign _T_56769 = $signed(buffer_0_308) + $signed(buffer_0_309); // @[Modules.scala 166:64:@2433.4]
  assign _T_56770 = _T_56769[13:0]; // @[Modules.scala 166:64:@2434.4]
  assign buffer_0_456 = $signed(_T_56770); // @[Modules.scala 166:64:@2435.4]
  assign _T_56772 = $signed(buffer_0_310) + $signed(buffer_0_311); // @[Modules.scala 166:64:@2437.4]
  assign _T_56773 = _T_56772[13:0]; // @[Modules.scala 166:64:@2438.4]
  assign buffer_0_457 = $signed(_T_56773); // @[Modules.scala 166:64:@2439.4]
  assign _T_56775 = $signed(buffer_0_312) + $signed(buffer_0_313); // @[Modules.scala 166:64:@2441.4]
  assign _T_56776 = _T_56775[13:0]; // @[Modules.scala 166:64:@2442.4]
  assign buffer_0_458 = $signed(_T_56776); // @[Modules.scala 166:64:@2443.4]
  assign _T_56778 = $signed(buffer_0_314) + $signed(buffer_0_315); // @[Modules.scala 166:64:@2445.4]
  assign _T_56779 = _T_56778[13:0]; // @[Modules.scala 166:64:@2446.4]
  assign buffer_0_459 = $signed(_T_56779); // @[Modules.scala 166:64:@2447.4]
  assign _T_56781 = $signed(buffer_0_316) + $signed(buffer_0_317); // @[Modules.scala 166:64:@2449.4]
  assign _T_56782 = _T_56781[13:0]; // @[Modules.scala 166:64:@2450.4]
  assign buffer_0_460 = $signed(_T_56782); // @[Modules.scala 166:64:@2451.4]
  assign _T_56784 = $signed(buffer_0_318) + $signed(buffer_0_319); // @[Modules.scala 166:64:@2453.4]
  assign _T_56785 = _T_56784[13:0]; // @[Modules.scala 166:64:@2454.4]
  assign buffer_0_461 = $signed(_T_56785); // @[Modules.scala 166:64:@2455.4]
  assign _T_56787 = $signed(buffer_0_320) + $signed(buffer_0_321); // @[Modules.scala 166:64:@2457.4]
  assign _T_56788 = _T_56787[13:0]; // @[Modules.scala 166:64:@2458.4]
  assign buffer_0_462 = $signed(_T_56788); // @[Modules.scala 166:64:@2459.4]
  assign _T_56790 = $signed(buffer_0_322) + $signed(buffer_0_323); // @[Modules.scala 166:64:@2461.4]
  assign _T_56791 = _T_56790[13:0]; // @[Modules.scala 166:64:@2462.4]
  assign buffer_0_463 = $signed(_T_56791); // @[Modules.scala 166:64:@2463.4]
  assign _T_56793 = $signed(buffer_0_324) + $signed(buffer_0_325); // @[Modules.scala 166:64:@2465.4]
  assign _T_56794 = _T_56793[13:0]; // @[Modules.scala 166:64:@2466.4]
  assign buffer_0_464 = $signed(_T_56794); // @[Modules.scala 166:64:@2467.4]
  assign _T_56796 = $signed(buffer_0_326) + $signed(buffer_0_327); // @[Modules.scala 166:64:@2469.4]
  assign _T_56797 = _T_56796[13:0]; // @[Modules.scala 166:64:@2470.4]
  assign buffer_0_465 = $signed(_T_56797); // @[Modules.scala 166:64:@2471.4]
  assign _T_56799 = $signed(buffer_0_328) + $signed(buffer_0_329); // @[Modules.scala 166:64:@2473.4]
  assign _T_56800 = _T_56799[13:0]; // @[Modules.scala 166:64:@2474.4]
  assign buffer_0_466 = $signed(_T_56800); // @[Modules.scala 166:64:@2475.4]
  assign _T_56802 = $signed(buffer_0_330) + $signed(buffer_0_331); // @[Modules.scala 166:64:@2477.4]
  assign _T_56803 = _T_56802[13:0]; // @[Modules.scala 166:64:@2478.4]
  assign buffer_0_467 = $signed(_T_56803); // @[Modules.scala 166:64:@2479.4]
  assign _T_56805 = $signed(buffer_0_332) + $signed(buffer_0_333); // @[Modules.scala 166:64:@2481.4]
  assign _T_56806 = _T_56805[13:0]; // @[Modules.scala 166:64:@2482.4]
  assign buffer_0_468 = $signed(_T_56806); // @[Modules.scala 166:64:@2483.4]
  assign _T_56808 = $signed(buffer_0_334) + $signed(buffer_0_335); // @[Modules.scala 166:64:@2485.4]
  assign _T_56809 = _T_56808[13:0]; // @[Modules.scala 166:64:@2486.4]
  assign buffer_0_469 = $signed(_T_56809); // @[Modules.scala 166:64:@2487.4]
  assign _T_56811 = $signed(buffer_0_336) + $signed(buffer_0_337); // @[Modules.scala 166:64:@2489.4]
  assign _T_56812 = _T_56811[13:0]; // @[Modules.scala 166:64:@2490.4]
  assign buffer_0_470 = $signed(_T_56812); // @[Modules.scala 166:64:@2491.4]
  assign _T_56814 = $signed(buffer_0_338) + $signed(buffer_0_339); // @[Modules.scala 166:64:@2493.4]
  assign _T_56815 = _T_56814[13:0]; // @[Modules.scala 166:64:@2494.4]
  assign buffer_0_471 = $signed(_T_56815); // @[Modules.scala 166:64:@2495.4]
  assign _T_56817 = $signed(buffer_0_340) + $signed(buffer_0_341); // @[Modules.scala 166:64:@2497.4]
  assign _T_56818 = _T_56817[13:0]; // @[Modules.scala 166:64:@2498.4]
  assign buffer_0_472 = $signed(_T_56818); // @[Modules.scala 166:64:@2499.4]
  assign _T_56820 = $signed(buffer_0_342) + $signed(buffer_0_343); // @[Modules.scala 166:64:@2501.4]
  assign _T_56821 = _T_56820[13:0]; // @[Modules.scala 166:64:@2502.4]
  assign buffer_0_473 = $signed(_T_56821); // @[Modules.scala 166:64:@2503.4]
  assign _T_56823 = $signed(buffer_0_344) + $signed(buffer_0_345); // @[Modules.scala 166:64:@2505.4]
  assign _T_56824 = _T_56823[13:0]; // @[Modules.scala 166:64:@2506.4]
  assign buffer_0_474 = $signed(_T_56824); // @[Modules.scala 166:64:@2507.4]
  assign _T_56826 = $signed(buffer_0_346) + $signed(buffer_0_347); // @[Modules.scala 166:64:@2509.4]
  assign _T_56827 = _T_56826[13:0]; // @[Modules.scala 166:64:@2510.4]
  assign buffer_0_475 = $signed(_T_56827); // @[Modules.scala 166:64:@2511.4]
  assign _T_56829 = $signed(buffer_0_348) + $signed(buffer_0_349); // @[Modules.scala 166:64:@2513.4]
  assign _T_56830 = _T_56829[13:0]; // @[Modules.scala 166:64:@2514.4]
  assign buffer_0_476 = $signed(_T_56830); // @[Modules.scala 166:64:@2515.4]
  assign _T_56832 = $signed(buffer_0_350) + $signed(buffer_0_351); // @[Modules.scala 166:64:@2517.4]
  assign _T_56833 = _T_56832[13:0]; // @[Modules.scala 166:64:@2518.4]
  assign buffer_0_477 = $signed(_T_56833); // @[Modules.scala 166:64:@2519.4]
  assign _T_56835 = $signed(buffer_0_352) + $signed(buffer_0_353); // @[Modules.scala 166:64:@2521.4]
  assign _T_56836 = _T_56835[13:0]; // @[Modules.scala 166:64:@2522.4]
  assign buffer_0_478 = $signed(_T_56836); // @[Modules.scala 166:64:@2523.4]
  assign _T_56838 = $signed(buffer_0_354) + $signed(buffer_0_355); // @[Modules.scala 166:64:@2525.4]
  assign _T_56839 = _T_56838[13:0]; // @[Modules.scala 166:64:@2526.4]
  assign buffer_0_479 = $signed(_T_56839); // @[Modules.scala 166:64:@2527.4]
  assign _T_56841 = $signed(buffer_0_356) + $signed(buffer_0_357); // @[Modules.scala 166:64:@2529.4]
  assign _T_56842 = _T_56841[13:0]; // @[Modules.scala 166:64:@2530.4]
  assign buffer_0_480 = $signed(_T_56842); // @[Modules.scala 166:64:@2531.4]
  assign _T_56844 = $signed(buffer_0_358) + $signed(buffer_0_359); // @[Modules.scala 166:64:@2533.4]
  assign _T_56845 = _T_56844[13:0]; // @[Modules.scala 166:64:@2534.4]
  assign buffer_0_481 = $signed(_T_56845); // @[Modules.scala 166:64:@2535.4]
  assign _T_56847 = $signed(buffer_0_360) + $signed(buffer_0_361); // @[Modules.scala 166:64:@2537.4]
  assign _T_56848 = _T_56847[13:0]; // @[Modules.scala 166:64:@2538.4]
  assign buffer_0_482 = $signed(_T_56848); // @[Modules.scala 166:64:@2539.4]
  assign _T_56850 = $signed(buffer_0_362) + $signed(buffer_0_363); // @[Modules.scala 166:64:@2541.4]
  assign _T_56851 = _T_56850[13:0]; // @[Modules.scala 166:64:@2542.4]
  assign buffer_0_483 = $signed(_T_56851); // @[Modules.scala 166:64:@2543.4]
  assign _T_56853 = $signed(buffer_0_364) + $signed(buffer_0_365); // @[Modules.scala 166:64:@2545.4]
  assign _T_56854 = _T_56853[13:0]; // @[Modules.scala 166:64:@2546.4]
  assign buffer_0_484 = $signed(_T_56854); // @[Modules.scala 166:64:@2547.4]
  assign _T_56856 = $signed(buffer_0_366) + $signed(buffer_0_367); // @[Modules.scala 166:64:@2549.4]
  assign _T_56857 = _T_56856[13:0]; // @[Modules.scala 166:64:@2550.4]
  assign buffer_0_485 = $signed(_T_56857); // @[Modules.scala 166:64:@2551.4]
  assign _T_56859 = $signed(buffer_0_368) + $signed(buffer_0_369); // @[Modules.scala 166:64:@2553.4]
  assign _T_56860 = _T_56859[13:0]; // @[Modules.scala 166:64:@2554.4]
  assign buffer_0_486 = $signed(_T_56860); // @[Modules.scala 166:64:@2555.4]
  assign _T_56862 = $signed(buffer_0_370) + $signed(buffer_0_371); // @[Modules.scala 166:64:@2557.4]
  assign _T_56863 = _T_56862[13:0]; // @[Modules.scala 166:64:@2558.4]
  assign buffer_0_487 = $signed(_T_56863); // @[Modules.scala 166:64:@2559.4]
  assign _T_56865 = $signed(buffer_0_372) + $signed(buffer_0_373); // @[Modules.scala 166:64:@2561.4]
  assign _T_56866 = _T_56865[13:0]; // @[Modules.scala 166:64:@2562.4]
  assign buffer_0_488 = $signed(_T_56866); // @[Modules.scala 166:64:@2563.4]
  assign _T_56868 = $signed(buffer_0_374) + $signed(buffer_0_375); // @[Modules.scala 166:64:@2565.4]
  assign _T_56869 = _T_56868[13:0]; // @[Modules.scala 166:64:@2566.4]
  assign buffer_0_489 = $signed(_T_56869); // @[Modules.scala 166:64:@2567.4]
  assign _T_56871 = $signed(buffer_0_376) + $signed(buffer_0_377); // @[Modules.scala 166:64:@2569.4]
  assign _T_56872 = _T_56871[13:0]; // @[Modules.scala 166:64:@2570.4]
  assign buffer_0_490 = $signed(_T_56872); // @[Modules.scala 166:64:@2571.4]
  assign _T_56874 = $signed(buffer_0_378) + $signed(buffer_0_379); // @[Modules.scala 166:64:@2573.4]
  assign _T_56875 = _T_56874[13:0]; // @[Modules.scala 166:64:@2574.4]
  assign buffer_0_491 = $signed(_T_56875); // @[Modules.scala 166:64:@2575.4]
  assign _T_56877 = $signed(buffer_0_380) + $signed(buffer_0_381); // @[Modules.scala 166:64:@2577.4]
  assign _T_56878 = _T_56877[13:0]; // @[Modules.scala 166:64:@2578.4]
  assign buffer_0_492 = $signed(_T_56878); // @[Modules.scala 166:64:@2579.4]
  assign _T_56880 = $signed(buffer_0_382) + $signed(buffer_0_383); // @[Modules.scala 166:64:@2581.4]
  assign _T_56881 = _T_56880[13:0]; // @[Modules.scala 166:64:@2582.4]
  assign buffer_0_493 = $signed(_T_56881); // @[Modules.scala 166:64:@2583.4]
  assign _T_56883 = $signed(buffer_0_384) + $signed(buffer_0_385); // @[Modules.scala 166:64:@2585.4]
  assign _T_56884 = _T_56883[13:0]; // @[Modules.scala 166:64:@2586.4]
  assign buffer_0_494 = $signed(_T_56884); // @[Modules.scala 166:64:@2587.4]
  assign _T_56886 = $signed(buffer_0_386) + $signed(buffer_0_387); // @[Modules.scala 166:64:@2589.4]
  assign _T_56887 = _T_56886[13:0]; // @[Modules.scala 166:64:@2590.4]
  assign buffer_0_495 = $signed(_T_56887); // @[Modules.scala 166:64:@2591.4]
  assign _T_56889 = $signed(buffer_0_388) + $signed(buffer_0_389); // @[Modules.scala 166:64:@2593.4]
  assign _T_56890 = _T_56889[13:0]; // @[Modules.scala 166:64:@2594.4]
  assign buffer_0_496 = $signed(_T_56890); // @[Modules.scala 166:64:@2595.4]
  assign _T_56892 = $signed(buffer_0_390) + $signed(buffer_0_391); // @[Modules.scala 166:64:@2597.4]
  assign _T_56893 = _T_56892[13:0]; // @[Modules.scala 166:64:@2598.4]
  assign buffer_0_497 = $signed(_T_56893); // @[Modules.scala 166:64:@2599.4]
  assign _T_56895 = $signed(buffer_0_392) + $signed(buffer_0_393); // @[Modules.scala 166:64:@2601.4]
  assign _T_56896 = _T_56895[13:0]; // @[Modules.scala 166:64:@2602.4]
  assign buffer_0_498 = $signed(_T_56896); // @[Modules.scala 166:64:@2603.4]
  assign _T_56898 = $signed(buffer_0_394) + $signed(buffer_0_395); // @[Modules.scala 166:64:@2605.4]
  assign _T_56899 = _T_56898[13:0]; // @[Modules.scala 166:64:@2606.4]
  assign buffer_0_499 = $signed(_T_56899); // @[Modules.scala 166:64:@2607.4]
  assign _T_56901 = $signed(buffer_0_396) + $signed(buffer_0_397); // @[Modules.scala 166:64:@2609.4]
  assign _T_56902 = _T_56901[13:0]; // @[Modules.scala 166:64:@2610.4]
  assign buffer_0_500 = $signed(_T_56902); // @[Modules.scala 166:64:@2611.4]
  assign _T_56904 = $signed(buffer_0_398) + $signed(buffer_0_399); // @[Modules.scala 166:64:@2613.4]
  assign _T_56905 = _T_56904[13:0]; // @[Modules.scala 166:64:@2614.4]
  assign buffer_0_501 = $signed(_T_56905); // @[Modules.scala 166:64:@2615.4]
  assign _T_56907 = $signed(buffer_0_400) + $signed(buffer_0_401); // @[Modules.scala 166:64:@2617.4]
  assign _T_56908 = _T_56907[13:0]; // @[Modules.scala 166:64:@2618.4]
  assign buffer_0_502 = $signed(_T_56908); // @[Modules.scala 166:64:@2619.4]
  assign _T_56910 = $signed(buffer_0_402) + $signed(buffer_0_403); // @[Modules.scala 166:64:@2621.4]
  assign _T_56911 = _T_56910[13:0]; // @[Modules.scala 166:64:@2622.4]
  assign buffer_0_503 = $signed(_T_56911); // @[Modules.scala 166:64:@2623.4]
  assign _T_56913 = $signed(buffer_0_404) + $signed(buffer_0_405); // @[Modules.scala 166:64:@2625.4]
  assign _T_56914 = _T_56913[13:0]; // @[Modules.scala 166:64:@2626.4]
  assign buffer_0_504 = $signed(_T_56914); // @[Modules.scala 166:64:@2627.4]
  assign _T_56916 = $signed(buffer_0_406) + $signed(buffer_0_407); // @[Modules.scala 166:64:@2629.4]
  assign _T_56917 = _T_56916[13:0]; // @[Modules.scala 166:64:@2630.4]
  assign buffer_0_505 = $signed(_T_56917); // @[Modules.scala 166:64:@2631.4]
  assign _T_56919 = $signed(buffer_0_408) + $signed(buffer_0_409); // @[Modules.scala 166:64:@2633.4]
  assign _T_56920 = _T_56919[13:0]; // @[Modules.scala 166:64:@2634.4]
  assign buffer_0_506 = $signed(_T_56920); // @[Modules.scala 166:64:@2635.4]
  assign _T_56922 = $signed(buffer_0_410) + $signed(buffer_0_411); // @[Modules.scala 166:64:@2637.4]
  assign _T_56923 = _T_56922[13:0]; // @[Modules.scala 166:64:@2638.4]
  assign buffer_0_507 = $signed(_T_56923); // @[Modules.scala 166:64:@2639.4]
  assign _T_56925 = $signed(buffer_0_412) + $signed(buffer_0_413); // @[Modules.scala 166:64:@2641.4]
  assign _T_56926 = _T_56925[13:0]; // @[Modules.scala 166:64:@2642.4]
  assign buffer_0_508 = $signed(_T_56926); // @[Modules.scala 166:64:@2643.4]
  assign _T_56928 = $signed(buffer_0_414) + $signed(buffer_0_415); // @[Modules.scala 166:64:@2645.4]
  assign _T_56929 = _T_56928[13:0]; // @[Modules.scala 166:64:@2646.4]
  assign buffer_0_509 = $signed(_T_56929); // @[Modules.scala 166:64:@2647.4]
  assign _T_56931 = $signed(buffer_0_416) + $signed(buffer_0_417); // @[Modules.scala 166:64:@2649.4]
  assign _T_56932 = _T_56931[13:0]; // @[Modules.scala 166:64:@2650.4]
  assign buffer_0_510 = $signed(_T_56932); // @[Modules.scala 166:64:@2651.4]
  assign _T_56934 = $signed(buffer_0_418) + $signed(buffer_0_419); // @[Modules.scala 166:64:@2653.4]
  assign _T_56935 = _T_56934[13:0]; // @[Modules.scala 166:64:@2654.4]
  assign buffer_0_511 = $signed(_T_56935); // @[Modules.scala 166:64:@2655.4]
  assign _T_56937 = $signed(buffer_0_420) + $signed(buffer_0_421); // @[Modules.scala 166:64:@2657.4]
  assign _T_56938 = _T_56937[13:0]; // @[Modules.scala 166:64:@2658.4]
  assign buffer_0_512 = $signed(_T_56938); // @[Modules.scala 166:64:@2659.4]
  assign _T_56940 = $signed(buffer_0_422) + $signed(buffer_0_423); // @[Modules.scala 166:64:@2661.4]
  assign _T_56941 = _T_56940[13:0]; // @[Modules.scala 166:64:@2662.4]
  assign buffer_0_513 = $signed(_T_56941); // @[Modules.scala 166:64:@2663.4]
  assign _T_56943 = $signed(buffer_0_424) + $signed(buffer_0_425); // @[Modules.scala 166:64:@2665.4]
  assign _T_56944 = _T_56943[13:0]; // @[Modules.scala 166:64:@2666.4]
  assign buffer_0_514 = $signed(_T_56944); // @[Modules.scala 166:64:@2667.4]
  assign _T_56946 = $signed(buffer_0_426) + $signed(buffer_0_427); // @[Modules.scala 166:64:@2669.4]
  assign _T_56947 = _T_56946[13:0]; // @[Modules.scala 166:64:@2670.4]
  assign buffer_0_515 = $signed(_T_56947); // @[Modules.scala 166:64:@2671.4]
  assign _T_56949 = $signed(buffer_0_428) + $signed(buffer_0_429); // @[Modules.scala 166:64:@2673.4]
  assign _T_56950 = _T_56949[13:0]; // @[Modules.scala 166:64:@2674.4]
  assign buffer_0_516 = $signed(_T_56950); // @[Modules.scala 166:64:@2675.4]
  assign _T_56952 = $signed(buffer_0_430) + $signed(buffer_0_431); // @[Modules.scala 166:64:@2677.4]
  assign _T_56953 = _T_56952[13:0]; // @[Modules.scala 166:64:@2678.4]
  assign buffer_0_517 = $signed(_T_56953); // @[Modules.scala 166:64:@2679.4]
  assign _T_56955 = $signed(buffer_0_432) + $signed(buffer_0_433); // @[Modules.scala 166:64:@2681.4]
  assign _T_56956 = _T_56955[13:0]; // @[Modules.scala 166:64:@2682.4]
  assign buffer_0_518 = $signed(_T_56956); // @[Modules.scala 166:64:@2683.4]
  assign _T_56958 = $signed(buffer_0_434) + $signed(buffer_0_435); // @[Modules.scala 166:64:@2685.4]
  assign _T_56959 = _T_56958[13:0]; // @[Modules.scala 166:64:@2686.4]
  assign buffer_0_519 = $signed(_T_56959); // @[Modules.scala 166:64:@2687.4]
  assign _T_56961 = $signed(buffer_0_436) + $signed(buffer_0_437); // @[Modules.scala 166:64:@2689.4]
  assign _T_56962 = _T_56961[13:0]; // @[Modules.scala 166:64:@2690.4]
  assign buffer_0_520 = $signed(_T_56962); // @[Modules.scala 166:64:@2691.4]
  assign _T_56964 = $signed(buffer_0_438) + $signed(buffer_0_439); // @[Modules.scala 166:64:@2693.4]
  assign _T_56965 = _T_56964[13:0]; // @[Modules.scala 166:64:@2694.4]
  assign buffer_0_521 = $signed(_T_56965); // @[Modules.scala 166:64:@2695.4]
  assign _T_56967 = $signed(buffer_0_440) + $signed(buffer_0_441); // @[Modules.scala 166:64:@2697.4]
  assign _T_56968 = _T_56967[13:0]; // @[Modules.scala 166:64:@2698.4]
  assign buffer_0_522 = $signed(_T_56968); // @[Modules.scala 166:64:@2699.4]
  assign _T_56970 = $signed(buffer_0_442) + $signed(buffer_0_443); // @[Modules.scala 166:64:@2701.4]
  assign _T_56971 = _T_56970[13:0]; // @[Modules.scala 166:64:@2702.4]
  assign buffer_0_523 = $signed(_T_56971); // @[Modules.scala 166:64:@2703.4]
  assign _T_56973 = $signed(buffer_0_444) + $signed(buffer_0_445); // @[Modules.scala 166:64:@2705.4]
  assign _T_56974 = _T_56973[13:0]; // @[Modules.scala 166:64:@2706.4]
  assign buffer_0_524 = $signed(_T_56974); // @[Modules.scala 166:64:@2707.4]
  assign _T_56976 = $signed(buffer_0_446) + $signed(buffer_0_447); // @[Modules.scala 166:64:@2709.4]
  assign _T_56977 = _T_56976[13:0]; // @[Modules.scala 166:64:@2710.4]
  assign buffer_0_525 = $signed(_T_56977); // @[Modules.scala 166:64:@2711.4]
  assign _T_56979 = $signed(buffer_0_448) + $signed(buffer_0_449); // @[Modules.scala 166:64:@2713.4]
  assign _T_56980 = _T_56979[13:0]; // @[Modules.scala 166:64:@2714.4]
  assign buffer_0_526 = $signed(_T_56980); // @[Modules.scala 166:64:@2715.4]
  assign _T_56982 = $signed(buffer_0_450) + $signed(buffer_0_451); // @[Modules.scala 166:64:@2717.4]
  assign _T_56983 = _T_56982[13:0]; // @[Modules.scala 166:64:@2718.4]
  assign buffer_0_527 = $signed(_T_56983); // @[Modules.scala 166:64:@2719.4]
  assign _T_56985 = $signed(buffer_0_453) + $signed(buffer_0_454); // @[Modules.scala 166:64:@2721.4]
  assign _T_56986 = _T_56985[13:0]; // @[Modules.scala 166:64:@2722.4]
  assign buffer_0_528 = $signed(_T_56986); // @[Modules.scala 166:64:@2723.4]
  assign _T_56988 = $signed(buffer_0_455) + $signed(buffer_0_456); // @[Modules.scala 166:64:@2725.4]
  assign _T_56989 = _T_56988[13:0]; // @[Modules.scala 166:64:@2726.4]
  assign buffer_0_529 = $signed(_T_56989); // @[Modules.scala 166:64:@2727.4]
  assign _T_56991 = $signed(buffer_0_457) + $signed(buffer_0_458); // @[Modules.scala 166:64:@2729.4]
  assign _T_56992 = _T_56991[13:0]; // @[Modules.scala 166:64:@2730.4]
  assign buffer_0_530 = $signed(_T_56992); // @[Modules.scala 166:64:@2731.4]
  assign _T_56994 = $signed(buffer_0_459) + $signed(buffer_0_460); // @[Modules.scala 166:64:@2733.4]
  assign _T_56995 = _T_56994[13:0]; // @[Modules.scala 166:64:@2734.4]
  assign buffer_0_531 = $signed(_T_56995); // @[Modules.scala 166:64:@2735.4]
  assign _T_56997 = $signed(buffer_0_461) + $signed(buffer_0_462); // @[Modules.scala 166:64:@2737.4]
  assign _T_56998 = _T_56997[13:0]; // @[Modules.scala 166:64:@2738.4]
  assign buffer_0_532 = $signed(_T_56998); // @[Modules.scala 166:64:@2739.4]
  assign _T_57000 = $signed(buffer_0_463) + $signed(buffer_0_464); // @[Modules.scala 166:64:@2741.4]
  assign _T_57001 = _T_57000[13:0]; // @[Modules.scala 166:64:@2742.4]
  assign buffer_0_533 = $signed(_T_57001); // @[Modules.scala 166:64:@2743.4]
  assign _T_57003 = $signed(buffer_0_465) + $signed(buffer_0_466); // @[Modules.scala 166:64:@2745.4]
  assign _T_57004 = _T_57003[13:0]; // @[Modules.scala 166:64:@2746.4]
  assign buffer_0_534 = $signed(_T_57004); // @[Modules.scala 166:64:@2747.4]
  assign _T_57006 = $signed(buffer_0_467) + $signed(buffer_0_468); // @[Modules.scala 166:64:@2749.4]
  assign _T_57007 = _T_57006[13:0]; // @[Modules.scala 166:64:@2750.4]
  assign buffer_0_535 = $signed(_T_57007); // @[Modules.scala 166:64:@2751.4]
  assign _T_57009 = $signed(buffer_0_469) + $signed(buffer_0_470); // @[Modules.scala 166:64:@2753.4]
  assign _T_57010 = _T_57009[13:0]; // @[Modules.scala 166:64:@2754.4]
  assign buffer_0_536 = $signed(_T_57010); // @[Modules.scala 166:64:@2755.4]
  assign _T_57012 = $signed(buffer_0_471) + $signed(buffer_0_472); // @[Modules.scala 166:64:@2757.4]
  assign _T_57013 = _T_57012[13:0]; // @[Modules.scala 166:64:@2758.4]
  assign buffer_0_537 = $signed(_T_57013); // @[Modules.scala 166:64:@2759.4]
  assign _T_57015 = $signed(buffer_0_473) + $signed(buffer_0_474); // @[Modules.scala 166:64:@2761.4]
  assign _T_57016 = _T_57015[13:0]; // @[Modules.scala 166:64:@2762.4]
  assign buffer_0_538 = $signed(_T_57016); // @[Modules.scala 166:64:@2763.4]
  assign _T_57018 = $signed(buffer_0_475) + $signed(buffer_0_476); // @[Modules.scala 166:64:@2765.4]
  assign _T_57019 = _T_57018[13:0]; // @[Modules.scala 166:64:@2766.4]
  assign buffer_0_539 = $signed(_T_57019); // @[Modules.scala 166:64:@2767.4]
  assign _T_57021 = $signed(buffer_0_477) + $signed(buffer_0_478); // @[Modules.scala 166:64:@2769.4]
  assign _T_57022 = _T_57021[13:0]; // @[Modules.scala 166:64:@2770.4]
  assign buffer_0_540 = $signed(_T_57022); // @[Modules.scala 166:64:@2771.4]
  assign _T_57024 = $signed(buffer_0_479) + $signed(buffer_0_480); // @[Modules.scala 166:64:@2773.4]
  assign _T_57025 = _T_57024[13:0]; // @[Modules.scala 166:64:@2774.4]
  assign buffer_0_541 = $signed(_T_57025); // @[Modules.scala 166:64:@2775.4]
  assign _T_57027 = $signed(buffer_0_481) + $signed(buffer_0_482); // @[Modules.scala 166:64:@2777.4]
  assign _T_57028 = _T_57027[13:0]; // @[Modules.scala 166:64:@2778.4]
  assign buffer_0_542 = $signed(_T_57028); // @[Modules.scala 166:64:@2779.4]
  assign _T_57030 = $signed(buffer_0_483) + $signed(buffer_0_484); // @[Modules.scala 166:64:@2781.4]
  assign _T_57031 = _T_57030[13:0]; // @[Modules.scala 166:64:@2782.4]
  assign buffer_0_543 = $signed(_T_57031); // @[Modules.scala 166:64:@2783.4]
  assign _T_57033 = $signed(buffer_0_485) + $signed(buffer_0_486); // @[Modules.scala 166:64:@2785.4]
  assign _T_57034 = _T_57033[13:0]; // @[Modules.scala 166:64:@2786.4]
  assign buffer_0_544 = $signed(_T_57034); // @[Modules.scala 166:64:@2787.4]
  assign _T_57036 = $signed(buffer_0_487) + $signed(buffer_0_488); // @[Modules.scala 166:64:@2789.4]
  assign _T_57037 = _T_57036[13:0]; // @[Modules.scala 166:64:@2790.4]
  assign buffer_0_545 = $signed(_T_57037); // @[Modules.scala 166:64:@2791.4]
  assign _T_57039 = $signed(buffer_0_489) + $signed(buffer_0_490); // @[Modules.scala 166:64:@2793.4]
  assign _T_57040 = _T_57039[13:0]; // @[Modules.scala 166:64:@2794.4]
  assign buffer_0_546 = $signed(_T_57040); // @[Modules.scala 166:64:@2795.4]
  assign _T_57042 = $signed(buffer_0_491) + $signed(buffer_0_492); // @[Modules.scala 166:64:@2797.4]
  assign _T_57043 = _T_57042[13:0]; // @[Modules.scala 166:64:@2798.4]
  assign buffer_0_547 = $signed(_T_57043); // @[Modules.scala 166:64:@2799.4]
  assign _T_57045 = $signed(buffer_0_493) + $signed(buffer_0_494); // @[Modules.scala 166:64:@2801.4]
  assign _T_57046 = _T_57045[13:0]; // @[Modules.scala 166:64:@2802.4]
  assign buffer_0_548 = $signed(_T_57046); // @[Modules.scala 166:64:@2803.4]
  assign _T_57048 = $signed(buffer_0_495) + $signed(buffer_0_496); // @[Modules.scala 166:64:@2805.4]
  assign _T_57049 = _T_57048[13:0]; // @[Modules.scala 166:64:@2806.4]
  assign buffer_0_549 = $signed(_T_57049); // @[Modules.scala 166:64:@2807.4]
  assign _T_57051 = $signed(buffer_0_497) + $signed(buffer_0_498); // @[Modules.scala 166:64:@2809.4]
  assign _T_57052 = _T_57051[13:0]; // @[Modules.scala 166:64:@2810.4]
  assign buffer_0_550 = $signed(_T_57052); // @[Modules.scala 166:64:@2811.4]
  assign _T_57054 = $signed(buffer_0_499) + $signed(buffer_0_500); // @[Modules.scala 166:64:@2813.4]
  assign _T_57055 = _T_57054[13:0]; // @[Modules.scala 166:64:@2814.4]
  assign buffer_0_551 = $signed(_T_57055); // @[Modules.scala 166:64:@2815.4]
  assign _T_57057 = $signed(buffer_0_501) + $signed(buffer_0_502); // @[Modules.scala 166:64:@2817.4]
  assign _T_57058 = _T_57057[13:0]; // @[Modules.scala 166:64:@2818.4]
  assign buffer_0_552 = $signed(_T_57058); // @[Modules.scala 166:64:@2819.4]
  assign _T_57060 = $signed(buffer_0_503) + $signed(buffer_0_504); // @[Modules.scala 166:64:@2821.4]
  assign _T_57061 = _T_57060[13:0]; // @[Modules.scala 166:64:@2822.4]
  assign buffer_0_553 = $signed(_T_57061); // @[Modules.scala 166:64:@2823.4]
  assign _T_57063 = $signed(buffer_0_505) + $signed(buffer_0_506); // @[Modules.scala 166:64:@2825.4]
  assign _T_57064 = _T_57063[13:0]; // @[Modules.scala 166:64:@2826.4]
  assign buffer_0_554 = $signed(_T_57064); // @[Modules.scala 166:64:@2827.4]
  assign _T_57066 = $signed(buffer_0_507) + $signed(buffer_0_508); // @[Modules.scala 166:64:@2829.4]
  assign _T_57067 = _T_57066[13:0]; // @[Modules.scala 166:64:@2830.4]
  assign buffer_0_555 = $signed(_T_57067); // @[Modules.scala 166:64:@2831.4]
  assign _T_57069 = $signed(buffer_0_509) + $signed(buffer_0_510); // @[Modules.scala 166:64:@2833.4]
  assign _T_57070 = _T_57069[13:0]; // @[Modules.scala 166:64:@2834.4]
  assign buffer_0_556 = $signed(_T_57070); // @[Modules.scala 166:64:@2835.4]
  assign _T_57072 = $signed(buffer_0_511) + $signed(buffer_0_512); // @[Modules.scala 166:64:@2837.4]
  assign _T_57073 = _T_57072[13:0]; // @[Modules.scala 166:64:@2838.4]
  assign buffer_0_557 = $signed(_T_57073); // @[Modules.scala 166:64:@2839.4]
  assign _T_57075 = $signed(buffer_0_513) + $signed(buffer_0_514); // @[Modules.scala 166:64:@2841.4]
  assign _T_57076 = _T_57075[13:0]; // @[Modules.scala 166:64:@2842.4]
  assign buffer_0_558 = $signed(_T_57076); // @[Modules.scala 166:64:@2843.4]
  assign _T_57078 = $signed(buffer_0_515) + $signed(buffer_0_516); // @[Modules.scala 166:64:@2845.4]
  assign _T_57079 = _T_57078[13:0]; // @[Modules.scala 166:64:@2846.4]
  assign buffer_0_559 = $signed(_T_57079); // @[Modules.scala 166:64:@2847.4]
  assign _T_57081 = $signed(buffer_0_517) + $signed(buffer_0_518); // @[Modules.scala 166:64:@2849.4]
  assign _T_57082 = _T_57081[13:0]; // @[Modules.scala 166:64:@2850.4]
  assign buffer_0_560 = $signed(_T_57082); // @[Modules.scala 166:64:@2851.4]
  assign _T_57084 = $signed(buffer_0_519) + $signed(buffer_0_520); // @[Modules.scala 166:64:@2853.4]
  assign _T_57085 = _T_57084[13:0]; // @[Modules.scala 166:64:@2854.4]
  assign buffer_0_561 = $signed(_T_57085); // @[Modules.scala 166:64:@2855.4]
  assign _T_57087 = $signed(buffer_0_521) + $signed(buffer_0_522); // @[Modules.scala 166:64:@2857.4]
  assign _T_57088 = _T_57087[13:0]; // @[Modules.scala 166:64:@2858.4]
  assign buffer_0_562 = $signed(_T_57088); // @[Modules.scala 166:64:@2859.4]
  assign _T_57090 = $signed(buffer_0_523) + $signed(buffer_0_524); // @[Modules.scala 166:64:@2861.4]
  assign _T_57091 = _T_57090[13:0]; // @[Modules.scala 166:64:@2862.4]
  assign buffer_0_563 = $signed(_T_57091); // @[Modules.scala 166:64:@2863.4]
  assign _T_57093 = $signed(buffer_0_525) + $signed(buffer_0_526); // @[Modules.scala 166:64:@2865.4]
  assign _T_57094 = _T_57093[13:0]; // @[Modules.scala 166:64:@2866.4]
  assign buffer_0_564 = $signed(_T_57094); // @[Modules.scala 166:64:@2867.4]
  assign _T_57096 = $signed(buffer_0_527) + $signed(buffer_0_452); // @[Modules.scala 172:66:@2869.4]
  assign _T_57097 = _T_57096[13:0]; // @[Modules.scala 172:66:@2870.4]
  assign buffer_0_565 = $signed(_T_57097); // @[Modules.scala 172:66:@2871.4]
  assign _T_57099 = $signed(buffer_0_528) + $signed(buffer_0_529); // @[Modules.scala 160:64:@2873.4]
  assign _T_57100 = _T_57099[13:0]; // @[Modules.scala 160:64:@2874.4]
  assign buffer_0_566 = $signed(_T_57100); // @[Modules.scala 160:64:@2875.4]
  assign _T_57102 = $signed(buffer_0_530) + $signed(buffer_0_531); // @[Modules.scala 160:64:@2877.4]
  assign _T_57103 = _T_57102[13:0]; // @[Modules.scala 160:64:@2878.4]
  assign buffer_0_567 = $signed(_T_57103); // @[Modules.scala 160:64:@2879.4]
  assign _T_57105 = $signed(buffer_0_532) + $signed(buffer_0_533); // @[Modules.scala 160:64:@2881.4]
  assign _T_57106 = _T_57105[13:0]; // @[Modules.scala 160:64:@2882.4]
  assign buffer_0_568 = $signed(_T_57106); // @[Modules.scala 160:64:@2883.4]
  assign _T_57108 = $signed(buffer_0_534) + $signed(buffer_0_535); // @[Modules.scala 160:64:@2885.4]
  assign _T_57109 = _T_57108[13:0]; // @[Modules.scala 160:64:@2886.4]
  assign buffer_0_569 = $signed(_T_57109); // @[Modules.scala 160:64:@2887.4]
  assign _T_57111 = $signed(buffer_0_536) + $signed(buffer_0_537); // @[Modules.scala 160:64:@2889.4]
  assign _T_57112 = _T_57111[13:0]; // @[Modules.scala 160:64:@2890.4]
  assign buffer_0_570 = $signed(_T_57112); // @[Modules.scala 160:64:@2891.4]
  assign _T_57114 = $signed(buffer_0_538) + $signed(buffer_0_539); // @[Modules.scala 160:64:@2893.4]
  assign _T_57115 = _T_57114[13:0]; // @[Modules.scala 160:64:@2894.4]
  assign buffer_0_571 = $signed(_T_57115); // @[Modules.scala 160:64:@2895.4]
  assign _T_57117 = $signed(buffer_0_540) + $signed(buffer_0_541); // @[Modules.scala 160:64:@2897.4]
  assign _T_57118 = _T_57117[13:0]; // @[Modules.scala 160:64:@2898.4]
  assign buffer_0_572 = $signed(_T_57118); // @[Modules.scala 160:64:@2899.4]
  assign _T_57120 = $signed(buffer_0_542) + $signed(buffer_0_543); // @[Modules.scala 160:64:@2901.4]
  assign _T_57121 = _T_57120[13:0]; // @[Modules.scala 160:64:@2902.4]
  assign buffer_0_573 = $signed(_T_57121); // @[Modules.scala 160:64:@2903.4]
  assign _T_57123 = $signed(buffer_0_544) + $signed(buffer_0_545); // @[Modules.scala 160:64:@2905.4]
  assign _T_57124 = _T_57123[13:0]; // @[Modules.scala 160:64:@2906.4]
  assign buffer_0_574 = $signed(_T_57124); // @[Modules.scala 160:64:@2907.4]
  assign _T_57126 = $signed(buffer_0_546) + $signed(buffer_0_547); // @[Modules.scala 160:64:@2909.4]
  assign _T_57127 = _T_57126[13:0]; // @[Modules.scala 160:64:@2910.4]
  assign buffer_0_575 = $signed(_T_57127); // @[Modules.scala 160:64:@2911.4]
  assign _T_57129 = $signed(buffer_0_548) + $signed(buffer_0_549); // @[Modules.scala 160:64:@2913.4]
  assign _T_57130 = _T_57129[13:0]; // @[Modules.scala 160:64:@2914.4]
  assign buffer_0_576 = $signed(_T_57130); // @[Modules.scala 160:64:@2915.4]
  assign _T_57132 = $signed(buffer_0_550) + $signed(buffer_0_551); // @[Modules.scala 160:64:@2917.4]
  assign _T_57133 = _T_57132[13:0]; // @[Modules.scala 160:64:@2918.4]
  assign buffer_0_577 = $signed(_T_57133); // @[Modules.scala 160:64:@2919.4]
  assign _T_57135 = $signed(buffer_0_552) + $signed(buffer_0_553); // @[Modules.scala 160:64:@2921.4]
  assign _T_57136 = _T_57135[13:0]; // @[Modules.scala 160:64:@2922.4]
  assign buffer_0_578 = $signed(_T_57136); // @[Modules.scala 160:64:@2923.4]
  assign _T_57138 = $signed(buffer_0_554) + $signed(buffer_0_555); // @[Modules.scala 160:64:@2925.4]
  assign _T_57139 = _T_57138[13:0]; // @[Modules.scala 160:64:@2926.4]
  assign buffer_0_579 = $signed(_T_57139); // @[Modules.scala 160:64:@2927.4]
  assign _T_57141 = $signed(buffer_0_556) + $signed(buffer_0_557); // @[Modules.scala 160:64:@2929.4]
  assign _T_57142 = _T_57141[13:0]; // @[Modules.scala 160:64:@2930.4]
  assign buffer_0_580 = $signed(_T_57142); // @[Modules.scala 160:64:@2931.4]
  assign _T_57144 = $signed(buffer_0_558) + $signed(buffer_0_559); // @[Modules.scala 160:64:@2933.4]
  assign _T_57145 = _T_57144[13:0]; // @[Modules.scala 160:64:@2934.4]
  assign buffer_0_581 = $signed(_T_57145); // @[Modules.scala 160:64:@2935.4]
  assign _T_57147 = $signed(buffer_0_560) + $signed(buffer_0_561); // @[Modules.scala 160:64:@2937.4]
  assign _T_57148 = _T_57147[13:0]; // @[Modules.scala 160:64:@2938.4]
  assign buffer_0_582 = $signed(_T_57148); // @[Modules.scala 160:64:@2939.4]
  assign _T_57150 = $signed(buffer_0_562) + $signed(buffer_0_563); // @[Modules.scala 160:64:@2941.4]
  assign _T_57151 = _T_57150[13:0]; // @[Modules.scala 160:64:@2942.4]
  assign buffer_0_583 = $signed(_T_57151); // @[Modules.scala 160:64:@2943.4]
  assign _T_57153 = $signed(buffer_0_564) + $signed(buffer_0_565); // @[Modules.scala 160:64:@2945.4]
  assign _T_57154 = _T_57153[13:0]; // @[Modules.scala 160:64:@2946.4]
  assign buffer_0_584 = $signed(_T_57154); // @[Modules.scala 160:64:@2947.4]
  assign _T_57156 = $signed(buffer_0_566) + $signed(buffer_0_567); // @[Modules.scala 166:64:@2949.4]
  assign _T_57157 = _T_57156[13:0]; // @[Modules.scala 166:64:@2950.4]
  assign buffer_0_585 = $signed(_T_57157); // @[Modules.scala 166:64:@2951.4]
  assign _T_57159 = $signed(buffer_0_568) + $signed(buffer_0_569); // @[Modules.scala 166:64:@2953.4]
  assign _T_57160 = _T_57159[13:0]; // @[Modules.scala 166:64:@2954.4]
  assign buffer_0_586 = $signed(_T_57160); // @[Modules.scala 166:64:@2955.4]
  assign _T_57162 = $signed(buffer_0_570) + $signed(buffer_0_571); // @[Modules.scala 166:64:@2957.4]
  assign _T_57163 = _T_57162[13:0]; // @[Modules.scala 166:64:@2958.4]
  assign buffer_0_587 = $signed(_T_57163); // @[Modules.scala 166:64:@2959.4]
  assign _T_57165 = $signed(buffer_0_572) + $signed(buffer_0_573); // @[Modules.scala 166:64:@2961.4]
  assign _T_57166 = _T_57165[13:0]; // @[Modules.scala 166:64:@2962.4]
  assign buffer_0_588 = $signed(_T_57166); // @[Modules.scala 166:64:@2963.4]
  assign _T_57168 = $signed(buffer_0_574) + $signed(buffer_0_575); // @[Modules.scala 166:64:@2965.4]
  assign _T_57169 = _T_57168[13:0]; // @[Modules.scala 166:64:@2966.4]
  assign buffer_0_589 = $signed(_T_57169); // @[Modules.scala 166:64:@2967.4]
  assign _T_57171 = $signed(buffer_0_576) + $signed(buffer_0_577); // @[Modules.scala 166:64:@2969.4]
  assign _T_57172 = _T_57171[13:0]; // @[Modules.scala 166:64:@2970.4]
  assign buffer_0_590 = $signed(_T_57172); // @[Modules.scala 166:64:@2971.4]
  assign _T_57174 = $signed(buffer_0_578) + $signed(buffer_0_579); // @[Modules.scala 166:64:@2973.4]
  assign _T_57175 = _T_57174[13:0]; // @[Modules.scala 166:64:@2974.4]
  assign buffer_0_591 = $signed(_T_57175); // @[Modules.scala 166:64:@2975.4]
  assign _T_57177 = $signed(buffer_0_580) + $signed(buffer_0_581); // @[Modules.scala 166:64:@2977.4]
  assign _T_57178 = _T_57177[13:0]; // @[Modules.scala 166:64:@2978.4]
  assign buffer_0_592 = $signed(_T_57178); // @[Modules.scala 166:64:@2979.4]
  assign _T_57180 = $signed(buffer_0_582) + $signed(buffer_0_583); // @[Modules.scala 166:64:@2981.4]
  assign _T_57181 = _T_57180[13:0]; // @[Modules.scala 166:64:@2982.4]
  assign buffer_0_593 = $signed(_T_57181); // @[Modules.scala 166:64:@2983.4]
  assign _T_57183 = $signed(buffer_0_585) + $signed(buffer_0_586); // @[Modules.scala 166:64:@2985.4]
  assign _T_57184 = _T_57183[13:0]; // @[Modules.scala 166:64:@2986.4]
  assign buffer_0_594 = $signed(_T_57184); // @[Modules.scala 166:64:@2987.4]
  assign _T_57186 = $signed(buffer_0_587) + $signed(buffer_0_588); // @[Modules.scala 166:64:@2989.4]
  assign _T_57187 = _T_57186[13:0]; // @[Modules.scala 166:64:@2990.4]
  assign buffer_0_595 = $signed(_T_57187); // @[Modules.scala 166:64:@2991.4]
  assign _T_57189 = $signed(buffer_0_589) + $signed(buffer_0_590); // @[Modules.scala 166:64:@2993.4]
  assign _T_57190 = _T_57189[13:0]; // @[Modules.scala 166:64:@2994.4]
  assign buffer_0_596 = $signed(_T_57190); // @[Modules.scala 166:64:@2995.4]
  assign _T_57192 = $signed(buffer_0_591) + $signed(buffer_0_592); // @[Modules.scala 166:64:@2997.4]
  assign _T_57193 = _T_57192[13:0]; // @[Modules.scala 166:64:@2998.4]
  assign buffer_0_597 = $signed(_T_57193); // @[Modules.scala 166:64:@2999.4]
  assign _T_57195 = $signed(buffer_0_593) + $signed(buffer_0_584); // @[Modules.scala 172:66:@3001.4]
  assign _T_57196 = _T_57195[13:0]; // @[Modules.scala 172:66:@3002.4]
  assign buffer_0_598 = $signed(_T_57196); // @[Modules.scala 172:66:@3003.4]
  assign _T_57198 = $signed(buffer_0_594) + $signed(buffer_0_595); // @[Modules.scala 166:64:@3005.4]
  assign _T_57199 = _T_57198[13:0]; // @[Modules.scala 166:64:@3006.4]
  assign buffer_0_599 = $signed(_T_57199); // @[Modules.scala 166:64:@3007.4]
  assign _T_57201 = $signed(buffer_0_596) + $signed(buffer_0_597); // @[Modules.scala 166:64:@3009.4]
  assign _T_57202 = _T_57201[13:0]; // @[Modules.scala 166:64:@3010.4]
  assign buffer_0_600 = $signed(_T_57202); // @[Modules.scala 166:64:@3011.4]
  assign _T_57204 = $signed(buffer_0_599) + $signed(buffer_0_600); // @[Modules.scala 160:64:@3013.4]
  assign _T_57205 = _T_57204[13:0]; // @[Modules.scala 160:64:@3014.4]
  assign buffer_0_601 = $signed(_T_57205); // @[Modules.scala 160:64:@3015.4]
  assign _T_57207 = $signed(buffer_0_601) + $signed(buffer_0_598); // @[Modules.scala 172:66:@3017.4]
  assign _T_57208 = _T_57207[13:0]; // @[Modules.scala 172:66:@3018.4]
  assign buffer_0_602 = $signed(_T_57208); // @[Modules.scala 172:66:@3019.4]
  assign _T_57225 = $signed(4'sh1) * $signed(io_in_19); // @[Modules.scala 143:74:@3214.4]
  assign _T_57227 = $signed(-4'sh1) * $signed(io_in_32); // @[Modules.scala 144:80:@3215.4]
  assign _GEN_76 = {{1{_T_57227[4]}},_T_57227}; // @[Modules.scala 143:103:@3216.4]
  assign _T_57228 = $signed(_T_57225) + $signed(_GEN_76); // @[Modules.scala 143:103:@3216.4]
  assign _T_57229 = _T_57228[5:0]; // @[Modules.scala 143:103:@3217.4]
  assign _T_57230 = $signed(_T_57229); // @[Modules.scala 143:103:@3218.4]
  assign _T_57232 = $signed(4'sh1) * $signed(io_in_34); // @[Modules.scala 143:74:@3220.4]
  assign _T_57234 = $signed(4'sh1) * $signed(io_in_35); // @[Modules.scala 144:80:@3221.4]
  assign _T_57235 = $signed(_T_57232) + $signed(_T_57234); // @[Modules.scala 143:103:@3222.4]
  assign _T_57236 = _T_57235[5:0]; // @[Modules.scala 143:103:@3223.4]
  assign _T_57237 = $signed(_T_57236); // @[Modules.scala 143:103:@3224.4]
  assign _T_57239 = $signed(-4'sh1) * $signed(io_in_36); // @[Modules.scala 143:74:@3226.4]
  assign _T_57241 = $signed(-4'sh1) * $signed(io_in_37); // @[Modules.scala 144:80:@3227.4]
  assign _T_57242 = $signed(_T_57239) + $signed(_T_57241); // @[Modules.scala 143:103:@3228.4]
  assign _T_57243 = _T_57242[4:0]; // @[Modules.scala 143:103:@3229.4]
  assign _T_57244 = $signed(_T_57243); // @[Modules.scala 143:103:@3230.4]
  assign _T_57248 = $signed(-4'sh1) * $signed(io_in_40); // @[Modules.scala 144:80:@3233.4]
  assign _GEN_77 = {{1{_T_57248[4]}},_T_57248}; // @[Modules.scala 143:103:@3234.4]
  assign _T_57249 = $signed(_T_54229) + $signed(_GEN_77); // @[Modules.scala 143:103:@3234.4]
  assign _T_57250 = _T_57249[5:0]; // @[Modules.scala 143:103:@3235.4]
  assign _T_57251 = $signed(_T_57250); // @[Modules.scala 143:103:@3236.4]
  assign _T_57253 = $signed(-4'sh1) * $signed(io_in_41); // @[Modules.scala 143:74:@3238.4]
  assign _T_57255 = $signed(-4'sh1) * $signed(io_in_42); // @[Modules.scala 144:80:@3239.4]
  assign _T_57256 = $signed(_T_57253) + $signed(_T_57255); // @[Modules.scala 143:103:@3240.4]
  assign _T_57257 = _T_57256[4:0]; // @[Modules.scala 143:103:@3241.4]
  assign _T_57258 = $signed(_T_57257); // @[Modules.scala 143:103:@3242.4]
  assign _T_57260 = $signed(-4'sh1) * $signed(io_in_43); // @[Modules.scala 143:74:@3244.4]
  assign _T_57262 = $signed(-4'sh1) * $signed(io_in_45); // @[Modules.scala 144:80:@3245.4]
  assign _T_57263 = $signed(_T_57260) + $signed(_T_57262); // @[Modules.scala 143:103:@3246.4]
  assign _T_57264 = _T_57263[4:0]; // @[Modules.scala 143:103:@3247.4]
  assign _T_57265 = $signed(_T_57264); // @[Modules.scala 143:103:@3248.4]
  assign _T_57267 = $signed(-4'sh1) * $signed(io_in_46); // @[Modules.scala 143:74:@3250.4]
  assign _GEN_78 = {{1{_T_57267[4]}},_T_57267}; // @[Modules.scala 143:103:@3252.4]
  assign _T_57270 = $signed(_GEN_78) + $signed(_T_54264); // @[Modules.scala 143:103:@3252.4]
  assign _T_57271 = _T_57270[5:0]; // @[Modules.scala 143:103:@3253.4]
  assign _T_57272 = $signed(_T_57271); // @[Modules.scala 143:103:@3254.4]
  assign _T_57274 = $signed(-4'sh1) * $signed(io_in_49); // @[Modules.scala 143:74:@3256.4]
  assign _T_57276 = $signed(-4'sh1) * $signed(io_in_50); // @[Modules.scala 144:80:@3257.4]
  assign _T_57277 = $signed(_T_57274) + $signed(_T_57276); // @[Modules.scala 143:103:@3258.4]
  assign _T_57278 = _T_57277[4:0]; // @[Modules.scala 143:103:@3259.4]
  assign _T_57279 = $signed(_T_57278); // @[Modules.scala 143:103:@3260.4]
  assign _T_57281 = $signed(-4'sh1) * $signed(io_in_51); // @[Modules.scala 143:74:@3262.4]
  assign _GEN_79 = {{1{_T_57281[4]}},_T_57281}; // @[Modules.scala 143:103:@3264.4]
  assign _T_57284 = $signed(_GEN_79) + $signed(_T_54278); // @[Modules.scala 143:103:@3264.4]
  assign _T_57285 = _T_57284[5:0]; // @[Modules.scala 143:103:@3265.4]
  assign _T_57286 = $signed(_T_57285); // @[Modules.scala 143:103:@3266.4]
  assign _T_57288 = $signed(-4'sh1) * $signed(io_in_60); // @[Modules.scala 143:74:@3268.4]
  assign _GEN_80 = {{1{_T_57288[4]}},_T_57288}; // @[Modules.scala 143:103:@3270.4]
  assign _T_57291 = $signed(_GEN_80) + $signed(_T_54283); // @[Modules.scala 143:103:@3270.4]
  assign _T_57292 = _T_57291[5:0]; // @[Modules.scala 143:103:@3271.4]
  assign _T_57293 = $signed(_T_57292); // @[Modules.scala 143:103:@3272.4]
  assign _T_57297 = $signed(-4'sh1) * $signed(io_in_63); // @[Modules.scala 144:80:@3275.4]
  assign _GEN_81 = {{1{_T_57297[4]}},_T_57297}; // @[Modules.scala 143:103:@3276.4]
  assign _T_57298 = $signed(_T_54285) + $signed(_GEN_81); // @[Modules.scala 143:103:@3276.4]
  assign _T_57299 = _T_57298[5:0]; // @[Modules.scala 143:103:@3277.4]
  assign _T_57300 = $signed(_T_57299); // @[Modules.scala 143:103:@3278.4]
  assign _T_57302 = $signed(-4'sh1) * $signed(io_in_64); // @[Modules.scala 143:74:@3280.4]
  assign _T_57304 = $signed(-4'sh1) * $signed(io_in_65); // @[Modules.scala 144:80:@3281.4]
  assign _T_57305 = $signed(_T_57302) + $signed(_T_57304); // @[Modules.scala 143:103:@3282.4]
  assign _T_57306 = _T_57305[4:0]; // @[Modules.scala 143:103:@3283.4]
  assign _T_57307 = $signed(_T_57306); // @[Modules.scala 143:103:@3284.4]
  assign _T_57309 = $signed(-4'sh1) * $signed(io_in_66); // @[Modules.scala 143:74:@3286.4]
  assign _T_57311 = $signed(-4'sh1) * $signed(io_in_67); // @[Modules.scala 144:80:@3287.4]
  assign _T_57312 = $signed(_T_57309) + $signed(_T_57311); // @[Modules.scala 143:103:@3288.4]
  assign _T_57313 = _T_57312[4:0]; // @[Modules.scala 143:103:@3289.4]
  assign _T_57314 = $signed(_T_57313); // @[Modules.scala 143:103:@3290.4]
  assign _T_57316 = $signed(-4'sh1) * $signed(io_in_68); // @[Modules.scala 143:74:@3292.4]
  assign _T_57318 = $signed(-4'sh1) * $signed(io_in_69); // @[Modules.scala 144:80:@3293.4]
  assign _T_57319 = $signed(_T_57316) + $signed(_T_57318); // @[Modules.scala 143:103:@3294.4]
  assign _T_57320 = _T_57319[4:0]; // @[Modules.scala 143:103:@3295.4]
  assign _T_57321 = $signed(_T_57320); // @[Modules.scala 143:103:@3296.4]
  assign _T_57323 = $signed(-4'sh1) * $signed(io_in_70); // @[Modules.scala 143:74:@3298.4]
  assign _T_57325 = $signed(-4'sh1) * $signed(io_in_71); // @[Modules.scala 144:80:@3299.4]
  assign _T_57326 = $signed(_T_57323) + $signed(_T_57325); // @[Modules.scala 143:103:@3300.4]
  assign _T_57327 = _T_57326[4:0]; // @[Modules.scala 143:103:@3301.4]
  assign _T_57328 = $signed(_T_57327); // @[Modules.scala 143:103:@3302.4]
  assign _T_57330 = $signed(-4'sh1) * $signed(io_in_72); // @[Modules.scala 143:74:@3304.4]
  assign _T_57332 = $signed(-4'sh1) * $signed(io_in_73); // @[Modules.scala 144:80:@3305.4]
  assign _T_57333 = $signed(_T_57330) + $signed(_T_57332); // @[Modules.scala 143:103:@3306.4]
  assign _T_57334 = _T_57333[4:0]; // @[Modules.scala 143:103:@3307.4]
  assign _T_57335 = $signed(_T_57334); // @[Modules.scala 143:103:@3308.4]
  assign _T_57337 = $signed(-4'sh1) * $signed(io_in_74); // @[Modules.scala 143:74:@3310.4]
  assign _T_57339 = $signed(-4'sh1) * $signed(io_in_75); // @[Modules.scala 144:80:@3311.4]
  assign _T_57340 = $signed(_T_57337) + $signed(_T_57339); // @[Modules.scala 143:103:@3312.4]
  assign _T_57341 = _T_57340[4:0]; // @[Modules.scala 143:103:@3313.4]
  assign _T_57342 = $signed(_T_57341); // @[Modules.scala 143:103:@3314.4]
  assign _T_57347 = $signed(_T_54334) + $signed(_T_54339); // @[Modules.scala 143:103:@3318.4]
  assign _T_57348 = _T_57347[5:0]; // @[Modules.scala 143:103:@3319.4]
  assign _T_57349 = $signed(_T_57348); // @[Modules.scala 143:103:@3320.4]
  assign _T_57354 = $signed(_T_54341) + $signed(_T_54346); // @[Modules.scala 143:103:@3324.4]
  assign _T_57355 = _T_57354[5:0]; // @[Modules.scala 143:103:@3325.4]
  assign _T_57356 = $signed(_T_57355); // @[Modules.scala 143:103:@3326.4]
  assign _T_57361 = $signed(_T_54348) + $signed(_T_54353); // @[Modules.scala 143:103:@3330.4]
  assign _T_57362 = _T_57361[5:0]; // @[Modules.scala 143:103:@3331.4]
  assign _T_57363 = $signed(_T_57362); // @[Modules.scala 143:103:@3332.4]
  assign _T_57368 = $signed(_GEN_1) + $signed(_T_54360); // @[Modules.scala 143:103:@3336.4]
  assign _T_57369 = _T_57368[5:0]; // @[Modules.scala 143:103:@3337.4]
  assign _T_57370 = $signed(_T_57369); // @[Modules.scala 143:103:@3338.4]
  assign _T_57375 = $signed(_T_54362) + $signed(_T_54367); // @[Modules.scala 143:103:@3342.4]
  assign _T_57376 = _T_57375[5:0]; // @[Modules.scala 143:103:@3343.4]
  assign _T_57377 = $signed(_T_57376); // @[Modules.scala 143:103:@3344.4]
  assign _T_57379 = $signed(-4'sh1) * $signed(io_in_90); // @[Modules.scala 143:74:@3346.4]
  assign _T_57381 = $signed(-4'sh1) * $signed(io_in_91); // @[Modules.scala 144:80:@3347.4]
  assign _T_57382 = $signed(_T_57379) + $signed(_T_57381); // @[Modules.scala 143:103:@3348.4]
  assign _T_57383 = _T_57382[4:0]; // @[Modules.scala 143:103:@3349.4]
  assign _T_57384 = $signed(_T_57383); // @[Modules.scala 143:103:@3350.4]
  assign _T_57386 = $signed(-4'sh1) * $signed(io_in_92); // @[Modules.scala 143:74:@3352.4]
  assign _T_57388 = $signed(-4'sh1) * $signed(io_in_93); // @[Modules.scala 144:80:@3353.4]
  assign _T_57389 = $signed(_T_57386) + $signed(_T_57388); // @[Modules.scala 143:103:@3354.4]
  assign _T_57390 = _T_57389[4:0]; // @[Modules.scala 143:103:@3355.4]
  assign _T_57391 = $signed(_T_57390); // @[Modules.scala 143:103:@3356.4]
  assign _T_57393 = $signed(-4'sh1) * $signed(io_in_94); // @[Modules.scala 143:74:@3358.4]
  assign _T_57395 = $signed(-4'sh1) * $signed(io_in_95); // @[Modules.scala 144:80:@3359.4]
  assign _T_57396 = $signed(_T_57393) + $signed(_T_57395); // @[Modules.scala 143:103:@3360.4]
  assign _T_57397 = _T_57396[4:0]; // @[Modules.scala 143:103:@3361.4]
  assign _T_57398 = $signed(_T_57397); // @[Modules.scala 143:103:@3362.4]
  assign _T_57400 = $signed(-4'sh1) * $signed(io_in_96); // @[Modules.scala 143:74:@3364.4]
  assign _T_57402 = $signed(-4'sh1) * $signed(io_in_97); // @[Modules.scala 144:80:@3365.4]
  assign _T_57403 = $signed(_T_57400) + $signed(_T_57402); // @[Modules.scala 143:103:@3366.4]
  assign _T_57404 = _T_57403[4:0]; // @[Modules.scala 143:103:@3367.4]
  assign _T_57405 = $signed(_T_57404); // @[Modules.scala 143:103:@3368.4]
  assign _T_57409 = $signed(-4'sh1) * $signed(io_in_101); // @[Modules.scala 144:80:@3371.4]
  assign _GEN_83 = {{1{_T_57409[4]}},_T_57409}; // @[Modules.scala 143:103:@3372.4]
  assign _T_57410 = $signed(_T_54402) + $signed(_GEN_83); // @[Modules.scala 143:103:@3372.4]
  assign _T_57411 = _T_57410[5:0]; // @[Modules.scala 143:103:@3373.4]
  assign _T_57412 = $signed(_T_57411); // @[Modules.scala 143:103:@3374.4]
  assign _T_57414 = $signed(-4'sh1) * $signed(io_in_102); // @[Modules.scala 143:74:@3376.4]
  assign _T_57416 = $signed(-4'sh1) * $signed(io_in_103); // @[Modules.scala 144:80:@3377.4]
  assign _T_57417 = $signed(_T_57414) + $signed(_T_57416); // @[Modules.scala 143:103:@3378.4]
  assign _T_57418 = _T_57417[4:0]; // @[Modules.scala 143:103:@3379.4]
  assign _T_57419 = $signed(_T_57418); // @[Modules.scala 143:103:@3380.4]
  assign _T_57421 = $signed(-4'sh1) * $signed(io_in_104); // @[Modules.scala 143:74:@3382.4]
  assign _T_57423 = $signed(-4'sh1) * $signed(io_in_105); // @[Modules.scala 144:80:@3383.4]
  assign _T_57424 = $signed(_T_57421) + $signed(_T_57423); // @[Modules.scala 143:103:@3384.4]
  assign _T_57425 = _T_57424[4:0]; // @[Modules.scala 143:103:@3385.4]
  assign _T_57426 = $signed(_T_57425); // @[Modules.scala 143:103:@3386.4]
  assign _T_57428 = $signed(-4'sh1) * $signed(io_in_106); // @[Modules.scala 143:74:@3388.4]
  assign _T_57430 = $signed(-4'sh1) * $signed(io_in_107); // @[Modules.scala 144:80:@3389.4]
  assign _T_57431 = $signed(_T_57428) + $signed(_T_57430); // @[Modules.scala 143:103:@3390.4]
  assign _T_57432 = _T_57431[4:0]; // @[Modules.scala 143:103:@3391.4]
  assign _T_57433 = $signed(_T_57432); // @[Modules.scala 143:103:@3392.4]
  assign _T_57435 = $signed(-4'sh1) * $signed(io_in_108); // @[Modules.scala 143:74:@3394.4]
  assign _GEN_84 = {{1{_T_57435[4]}},_T_57435}; // @[Modules.scala 143:103:@3396.4]
  assign _T_57438 = $signed(_GEN_84) + $signed(_T_54437); // @[Modules.scala 143:103:@3396.4]
  assign _T_57439 = _T_57438[5:0]; // @[Modules.scala 143:103:@3397.4]
  assign _T_57440 = $signed(_T_57439); // @[Modules.scala 143:103:@3398.4]
  assign _T_57442 = $signed(4'sh1) * $signed(io_in_110); // @[Modules.scala 143:74:@3400.4]
  assign _T_57445 = $signed(_T_57442) + $signed(_T_54444); // @[Modules.scala 143:103:@3402.4]
  assign _T_57446 = _T_57445[5:0]; // @[Modules.scala 143:103:@3403.4]
  assign _T_57447 = $signed(_T_57446); // @[Modules.scala 143:103:@3404.4]
  assign _T_57449 = $signed(4'sh1) * $signed(io_in_114); // @[Modules.scala 143:74:@3406.4]
  assign _T_57451 = $signed(4'sh1) * $signed(io_in_115); // @[Modules.scala 144:80:@3407.4]
  assign _T_57452 = $signed(_T_57449) + $signed(_T_57451); // @[Modules.scala 143:103:@3408.4]
  assign _T_57453 = _T_57452[5:0]; // @[Modules.scala 143:103:@3409.4]
  assign _T_57454 = $signed(_T_57453); // @[Modules.scala 143:103:@3410.4]
  assign _T_57456 = $signed(4'sh1) * $signed(io_in_117); // @[Modules.scala 143:74:@3412.4]
  assign _T_57458 = $signed(4'sh1) * $signed(io_in_118); // @[Modules.scala 144:80:@3413.4]
  assign _T_57459 = $signed(_T_57456) + $signed(_T_57458); // @[Modules.scala 143:103:@3414.4]
  assign _T_57460 = _T_57459[5:0]; // @[Modules.scala 143:103:@3415.4]
  assign _T_57461 = $signed(_T_57460); // @[Modules.scala 143:103:@3416.4]
  assign _T_57466 = $signed(_T_54460) + $signed(_T_54465); // @[Modules.scala 143:103:@3420.4]
  assign _T_57467 = _T_57466[5:0]; // @[Modules.scala 143:103:@3421.4]
  assign _T_57468 = $signed(_T_57467); // @[Modules.scala 143:103:@3422.4]
  assign _T_57473 = $signed(_T_54467) + $signed(_T_54472); // @[Modules.scala 143:103:@3426.4]
  assign _T_57474 = _T_57473[5:0]; // @[Modules.scala 143:103:@3427.4]
  assign _T_57475 = $signed(_T_57474); // @[Modules.scala 143:103:@3428.4]
  assign _T_57480 = $signed(_T_54474) + $signed(_T_54479); // @[Modules.scala 143:103:@3432.4]
  assign _T_57481 = _T_57480[5:0]; // @[Modules.scala 143:103:@3433.4]
  assign _T_57482 = $signed(_T_57481); // @[Modules.scala 143:103:@3434.4]
  assign _T_57486 = $signed(-4'sh1) * $signed(io_in_128); // @[Modules.scala 144:80:@3437.4]
  assign _GEN_85 = {{1{_T_57486[4]}},_T_57486}; // @[Modules.scala 143:103:@3438.4]
  assign _T_57487 = $signed(_T_54481) + $signed(_GEN_85); // @[Modules.scala 143:103:@3438.4]
  assign _T_57488 = _T_57487[5:0]; // @[Modules.scala 143:103:@3439.4]
  assign _T_57489 = $signed(_T_57488); // @[Modules.scala 143:103:@3440.4]
  assign _T_57498 = $signed(4'sh1) * $signed(io_in_132); // @[Modules.scala 143:74:@3448.4]
  assign _T_57501 = $signed(_T_57498) + $signed(_T_54500); // @[Modules.scala 143:103:@3450.4]
  assign _T_57502 = _T_57501[5:0]; // @[Modules.scala 143:103:@3451.4]
  assign _T_57503 = $signed(_T_57502); // @[Modules.scala 143:103:@3452.4]
  assign _T_57507 = $signed(4'sh1) * $signed(io_in_135); // @[Modules.scala 144:80:@3455.4]
  assign _T_57508 = $signed(_T_54502) + $signed(_T_57507); // @[Modules.scala 143:103:@3456.4]
  assign _T_57509 = _T_57508[5:0]; // @[Modules.scala 143:103:@3457.4]
  assign _T_57510 = $signed(_T_57509); // @[Modules.scala 143:103:@3458.4]
  assign _T_57512 = $signed(4'sh1) * $signed(io_in_136); // @[Modules.scala 143:74:@3460.4]
  assign _T_57514 = $signed(4'sh1) * $signed(io_in_137); // @[Modules.scala 144:80:@3461.4]
  assign _T_57515 = $signed(_T_57512) + $signed(_T_57514); // @[Modules.scala 143:103:@3462.4]
  assign _T_57516 = _T_57515[5:0]; // @[Modules.scala 143:103:@3463.4]
  assign _T_57517 = $signed(_T_57516); // @[Modules.scala 143:103:@3464.4]
  assign _T_57521 = $signed(-4'sh1) * $signed(io_in_139); // @[Modules.scala 144:80:@3467.4]
  assign _GEN_86 = {{1{_T_57521[4]}},_T_57521}; // @[Modules.scala 143:103:@3468.4]
  assign _T_57522 = $signed(_T_54516) + $signed(_GEN_86); // @[Modules.scala 143:103:@3468.4]
  assign _T_57523 = _T_57522[5:0]; // @[Modules.scala 143:103:@3469.4]
  assign _T_57524 = $signed(_T_57523); // @[Modules.scala 143:103:@3470.4]
  assign _T_57526 = $signed(4'sh1) * $signed(io_in_142); // @[Modules.scala 143:74:@3472.4]
  assign _T_57529 = $signed(_T_57526) + $signed(_T_54521); // @[Modules.scala 143:103:@3474.4]
  assign _T_57530 = _T_57529[5:0]; // @[Modules.scala 143:103:@3475.4]
  assign _T_57531 = $signed(_T_57530); // @[Modules.scala 143:103:@3476.4]
  assign _T_57533 = $signed(4'sh1) * $signed(io_in_144); // @[Modules.scala 143:74:@3478.4]
  assign _T_57535 = $signed(4'sh1) * $signed(io_in_145); // @[Modules.scala 144:80:@3479.4]
  assign _T_57536 = $signed(_T_57533) + $signed(_T_57535); // @[Modules.scala 143:103:@3480.4]
  assign _T_57537 = _T_57536[5:0]; // @[Modules.scala 143:103:@3481.4]
  assign _T_57538 = $signed(_T_57537); // @[Modules.scala 143:103:@3482.4]
  assign _T_57540 = $signed(4'sh1) * $signed(io_in_146); // @[Modules.scala 143:74:@3484.4]
  assign _T_57542 = $signed(4'sh1) * $signed(io_in_147); // @[Modules.scala 144:80:@3485.4]
  assign _T_57543 = $signed(_T_57540) + $signed(_T_57542); // @[Modules.scala 143:103:@3486.4]
  assign _T_57544 = _T_57543[5:0]; // @[Modules.scala 143:103:@3487.4]
  assign _T_57545 = $signed(_T_57544); // @[Modules.scala 143:103:@3488.4]
  assign _T_57556 = $signed(4'sh1) * $signed(io_in_152); // @[Modules.scala 144:80:@3497.4]
  assign _T_57557 = $signed(_T_54542) + $signed(_T_57556); // @[Modules.scala 143:103:@3498.4]
  assign _T_57558 = _T_57557[5:0]; // @[Modules.scala 143:103:@3499.4]
  assign _T_57559 = $signed(_T_57558); // @[Modules.scala 143:103:@3500.4]
  assign _T_57561 = $signed(-4'sh1) * $signed(io_in_154); // @[Modules.scala 143:74:@3502.4]
  assign _T_57563 = $signed(-4'sh1) * $signed(io_in_155); // @[Modules.scala 144:80:@3503.4]
  assign _T_57564 = $signed(_T_57561) + $signed(_T_57563); // @[Modules.scala 143:103:@3504.4]
  assign _T_57565 = _T_57564[4:0]; // @[Modules.scala 143:103:@3505.4]
  assign _T_57566 = $signed(_T_57565); // @[Modules.scala 143:103:@3506.4]
  assign _T_57571 = $signed(_T_54544) + $signed(_T_54549); // @[Modules.scala 143:103:@3510.4]
  assign _T_57572 = _T_57571[4:0]; // @[Modules.scala 143:103:@3511.4]
  assign _T_57573 = $signed(_T_57572); // @[Modules.scala 143:103:@3512.4]
  assign _T_57575 = $signed(-4'sh1) * $signed(io_in_158); // @[Modules.scala 143:74:@3514.4]
  assign _GEN_87 = {{1{_T_57575[4]}},_T_57575}; // @[Modules.scala 143:103:@3516.4]
  assign _T_57578 = $signed(_GEN_87) + $signed(_T_54556); // @[Modules.scala 143:103:@3516.4]
  assign _T_57579 = _T_57578[5:0]; // @[Modules.scala 143:103:@3517.4]
  assign _T_57580 = $signed(_T_57579); // @[Modules.scala 143:103:@3518.4]
  assign _T_57585 = $signed(_T_54558) + $signed(_T_54563); // @[Modules.scala 143:103:@3522.4]
  assign _T_57586 = _T_57585[4:0]; // @[Modules.scala 143:103:@3523.4]
  assign _T_57587 = $signed(_T_57586); // @[Modules.scala 143:103:@3524.4]
  assign _T_57592 = $signed(_T_54565) + $signed(_T_54570); // @[Modules.scala 143:103:@3528.4]
  assign _T_57593 = _T_57592[4:0]; // @[Modules.scala 143:103:@3529.4]
  assign _T_57594 = $signed(_T_57593); // @[Modules.scala 143:103:@3530.4]
  assign _T_57596 = $signed(-4'sh1) * $signed(io_in_166); // @[Modules.scala 143:74:@3532.4]
  assign _GEN_88 = {{1{_T_57596[4]}},_T_57596}; // @[Modules.scala 143:103:@3534.4]
  assign _T_57599 = $signed(_GEN_88) + $signed(_T_54577); // @[Modules.scala 143:103:@3534.4]
  assign _T_57600 = _T_57599[5:0]; // @[Modules.scala 143:103:@3535.4]
  assign _T_57601 = $signed(_T_57600); // @[Modules.scala 143:103:@3536.4]
  assign _T_57619 = $signed(-4'sh1) * $signed(io_in_177); // @[Modules.scala 144:80:@3551.4]
  assign _GEN_90 = {{1{_T_57619[4]}},_T_57619}; // @[Modules.scala 143:103:@3552.4]
  assign _T_57620 = $signed(_T_54598) + $signed(_GEN_90); // @[Modules.scala 143:103:@3552.4]
  assign _T_57621 = _T_57620[5:0]; // @[Modules.scala 143:103:@3553.4]
  assign _T_57622 = $signed(_T_57621); // @[Modules.scala 143:103:@3554.4]
  assign _T_57626 = $signed(4'sh1) * $signed(io_in_179); // @[Modules.scala 144:80:@3557.4]
  assign _T_57627 = $signed(_GEN_14) + $signed(_T_57626); // @[Modules.scala 143:103:@3558.4]
  assign _T_57628 = _T_57627[5:0]; // @[Modules.scala 143:103:@3559.4]
  assign _T_57629 = $signed(_T_57628); // @[Modules.scala 143:103:@3560.4]
  assign _T_57631 = $signed(4'sh1) * $signed(io_in_180); // @[Modules.scala 143:74:@3562.4]
  assign _T_57633 = $signed(4'sh1) * $signed(io_in_181); // @[Modules.scala 144:80:@3563.4]
  assign _T_57634 = $signed(_T_57631) + $signed(_T_57633); // @[Modules.scala 143:103:@3564.4]
  assign _T_57635 = _T_57634[5:0]; // @[Modules.scala 143:103:@3565.4]
  assign _T_57636 = $signed(_T_57635); // @[Modules.scala 143:103:@3566.4]
  assign _T_57638 = $signed(4'sh1) * $signed(io_in_182); // @[Modules.scala 143:74:@3568.4]
  assign _T_57640 = $signed(4'sh1) * $signed(io_in_183); // @[Modules.scala 144:80:@3569.4]
  assign _T_57641 = $signed(_T_57638) + $signed(_T_57640); // @[Modules.scala 143:103:@3570.4]
  assign _T_57642 = _T_57641[5:0]; // @[Modules.scala 143:103:@3571.4]
  assign _T_57643 = $signed(_T_57642); // @[Modules.scala 143:103:@3572.4]
  assign _T_57645 = $signed(4'sh1) * $signed(io_in_184); // @[Modules.scala 143:74:@3574.4]
  assign _GEN_92 = {{1{_T_54626[4]}},_T_54626}; // @[Modules.scala 143:103:@3576.4]
  assign _T_57648 = $signed(_T_57645) + $signed(_GEN_92); // @[Modules.scala 143:103:@3576.4]
  assign _T_57649 = _T_57648[5:0]; // @[Modules.scala 143:103:@3577.4]
  assign _T_57650 = $signed(_T_57649); // @[Modules.scala 143:103:@3578.4]
  assign _T_57655 = $signed(_T_54628) + $signed(_T_54633); // @[Modules.scala 143:103:@3582.4]
  assign _T_57656 = _T_57655[4:0]; // @[Modules.scala 143:103:@3583.4]
  assign _T_57657 = $signed(_T_57656); // @[Modules.scala 143:103:@3584.4]
  assign _T_57662 = $signed(_T_54635) + $signed(_T_54640); // @[Modules.scala 143:103:@3588.4]
  assign _T_57663 = _T_57662[4:0]; // @[Modules.scala 143:103:@3589.4]
  assign _T_57664 = $signed(_T_57663); // @[Modules.scala 143:103:@3590.4]
  assign _T_57669 = $signed(_T_54642) + $signed(_T_54647); // @[Modules.scala 143:103:@3594.4]
  assign _T_57670 = _T_57669[4:0]; // @[Modules.scala 143:103:@3595.4]
  assign _T_57671 = $signed(_T_57670); // @[Modules.scala 143:103:@3596.4]
  assign _T_57675 = $signed(4'sh1) * $signed(io_in_196); // @[Modules.scala 144:80:@3599.4]
  assign _GEN_93 = {{1{_T_54649[4]}},_T_54649}; // @[Modules.scala 143:103:@3600.4]
  assign _T_57676 = $signed(_GEN_93) + $signed(_T_57675); // @[Modules.scala 143:103:@3600.4]
  assign _T_57677 = _T_57676[5:0]; // @[Modules.scala 143:103:@3601.4]
  assign _T_57678 = $signed(_T_57677); // @[Modules.scala 143:103:@3602.4]
  assign _T_57701 = $signed(-4'sh1) * $signed(io_in_203); // @[Modules.scala 143:74:@3622.4]
  assign _T_57704 = $signed(_T_57701) + $signed(_T_54684); // @[Modules.scala 143:103:@3624.4]
  assign _T_57705 = _T_57704[4:0]; // @[Modules.scala 143:103:@3625.4]
  assign _T_57706 = $signed(_T_57705); // @[Modules.scala 143:103:@3626.4]
  assign _T_57708 = $signed(4'sh1) * $signed(io_in_207); // @[Modules.scala 143:74:@3628.4]
  assign _T_57710 = $signed(4'sh1) * $signed(io_in_208); // @[Modules.scala 144:80:@3629.4]
  assign _T_57711 = $signed(_T_57708) + $signed(_T_57710); // @[Modules.scala 143:103:@3630.4]
  assign _T_57712 = _T_57711[5:0]; // @[Modules.scala 143:103:@3631.4]
  assign _T_57713 = $signed(_T_57712); // @[Modules.scala 143:103:@3632.4]
  assign _T_57715 = $signed(4'sh1) * $signed(io_in_209); // @[Modules.scala 143:74:@3634.4]
  assign _T_57717 = $signed(4'sh1) * $signed(io_in_210); // @[Modules.scala 144:80:@3635.4]
  assign _T_57718 = $signed(_T_57715) + $signed(_T_57717); // @[Modules.scala 143:103:@3636.4]
  assign _T_57719 = _T_57718[5:0]; // @[Modules.scala 143:103:@3637.4]
  assign _T_57720 = $signed(_T_57719); // @[Modules.scala 143:103:@3638.4]
  assign _T_57722 = $signed(4'sh1) * $signed(io_in_211); // @[Modules.scala 143:74:@3640.4]
  assign _T_57724 = $signed(4'sh1) * $signed(io_in_212); // @[Modules.scala 144:80:@3641.4]
  assign _T_57725 = $signed(_T_57722) + $signed(_T_57724); // @[Modules.scala 143:103:@3642.4]
  assign _T_57726 = _T_57725[5:0]; // @[Modules.scala 143:103:@3643.4]
  assign _T_57727 = $signed(_T_57726); // @[Modules.scala 143:103:@3644.4]
  assign _T_57729 = $signed(4'sh1) * $signed(io_in_213); // @[Modules.scala 143:74:@3646.4]
  assign _GEN_94 = {{1{_T_54698[4]}},_T_54698}; // @[Modules.scala 143:103:@3648.4]
  assign _T_57732 = $signed(_T_57729) + $signed(_GEN_94); // @[Modules.scala 143:103:@3648.4]
  assign _T_57733 = _T_57732[5:0]; // @[Modules.scala 143:103:@3649.4]
  assign _T_57734 = $signed(_T_57733); // @[Modules.scala 143:103:@3650.4]
  assign _T_57736 = $signed(4'sh1) * $signed(io_in_215); // @[Modules.scala 143:74:@3652.4]
  assign _T_57738 = $signed(4'sh1) * $signed(io_in_216); // @[Modules.scala 144:80:@3653.4]
  assign _T_57739 = $signed(_T_57736) + $signed(_T_57738); // @[Modules.scala 143:103:@3654.4]
  assign _T_57740 = _T_57739[5:0]; // @[Modules.scala 143:103:@3655.4]
  assign _T_57741 = $signed(_T_57740); // @[Modules.scala 143:103:@3656.4]
  assign _T_57757 = $signed(-4'sh1) * $signed(io_in_222); // @[Modules.scala 143:74:@3670.4]
  assign _T_57759 = $signed(-4'sh1) * $signed(io_in_223); // @[Modules.scala 144:80:@3671.4]
  assign _T_57760 = $signed(_T_57757) + $signed(_T_57759); // @[Modules.scala 143:103:@3672.4]
  assign _T_57761 = _T_57760[4:0]; // @[Modules.scala 143:103:@3673.4]
  assign _T_57762 = $signed(_T_57761); // @[Modules.scala 143:103:@3674.4]
  assign _T_57764 = $signed(4'sh1) * $signed(io_in_224); // @[Modules.scala 143:74:@3676.4]
  assign _T_57767 = $signed(_T_57764) + $signed(_T_54731); // @[Modules.scala 143:103:@3678.4]
  assign _T_57768 = _T_57767[5:0]; // @[Modules.scala 143:103:@3679.4]
  assign _T_57769 = $signed(_T_57768); // @[Modules.scala 143:103:@3680.4]
  assign _T_57774 = $signed(_T_54733) + $signed(_T_54738); // @[Modules.scala 143:103:@3684.4]
  assign _T_57775 = _T_57774[5:0]; // @[Modules.scala 143:103:@3685.4]
  assign _T_57776 = $signed(_T_57775); // @[Modules.scala 143:103:@3686.4]
  assign _T_57781 = $signed(_T_54740) + $signed(_T_54745); // @[Modules.scala 143:103:@3690.4]
  assign _T_57782 = _T_57781[5:0]; // @[Modules.scala 143:103:@3691.4]
  assign _T_57783 = $signed(_T_57782); // @[Modules.scala 143:103:@3692.4]
  assign _T_57787 = $signed(-4'sh1) * $signed(io_in_231); // @[Modules.scala 144:80:@3695.4]
  assign _GEN_95 = {{1{_T_57787[4]}},_T_57787}; // @[Modules.scala 143:103:@3696.4]
  assign _T_57788 = $signed(_T_54747) + $signed(_GEN_95); // @[Modules.scala 143:103:@3696.4]
  assign _T_57789 = _T_57788[5:0]; // @[Modules.scala 143:103:@3697.4]
  assign _T_57790 = $signed(_T_57789); // @[Modules.scala 143:103:@3698.4]
  assign _T_57794 = $signed(-4'sh1) * $signed(io_in_235); // @[Modules.scala 144:80:@3701.4]
  assign _T_57795 = $signed(_T_54759) + $signed(_T_57794); // @[Modules.scala 143:103:@3702.4]
  assign _T_57796 = _T_57795[4:0]; // @[Modules.scala 143:103:@3703.4]
  assign _T_57797 = $signed(_T_57796); // @[Modules.scala 143:103:@3704.4]
  assign _T_57799 = $signed(4'sh1) * $signed(io_in_237); // @[Modules.scala 143:74:@3706.4]
  assign _T_57802 = $signed(_T_57799) + $signed(_T_54766); // @[Modules.scala 143:103:@3708.4]
  assign _T_57803 = _T_57802[5:0]; // @[Modules.scala 143:103:@3709.4]
  assign _T_57804 = $signed(_T_57803); // @[Modules.scala 143:103:@3710.4]
  assign _T_57806 = $signed(4'sh1) * $signed(io_in_239); // @[Modules.scala 143:74:@3712.4]
  assign _T_57808 = $signed(4'sh1) * $signed(io_in_240); // @[Modules.scala 144:80:@3713.4]
  assign _T_57809 = $signed(_T_57806) + $signed(_T_57808); // @[Modules.scala 143:103:@3714.4]
  assign _T_57810 = _T_57809[5:0]; // @[Modules.scala 143:103:@3715.4]
  assign _T_57811 = $signed(_T_57810); // @[Modules.scala 143:103:@3716.4]
  assign _T_57813 = $signed(4'sh1) * $signed(io_in_241); // @[Modules.scala 143:74:@3718.4]
  assign _T_57815 = $signed(4'sh1) * $signed(io_in_242); // @[Modules.scala 144:80:@3719.4]
  assign _T_57816 = $signed(_T_57813) + $signed(_T_57815); // @[Modules.scala 143:103:@3720.4]
  assign _T_57817 = _T_57816[5:0]; // @[Modules.scala 143:103:@3721.4]
  assign _T_57818 = $signed(_T_57817); // @[Modules.scala 143:103:@3722.4]
  assign _T_57848 = $signed(-4'sh1) * $signed(io_in_251); // @[Modules.scala 143:74:@3748.4]
  assign _T_57850 = $signed(4'sh1) * $signed(io_in_252); // @[Modules.scala 144:80:@3749.4]
  assign _GEN_96 = {{1{_T_57848[4]}},_T_57848}; // @[Modules.scala 143:103:@3750.4]
  assign _T_57851 = $signed(_GEN_96) + $signed(_T_57850); // @[Modules.scala 143:103:@3750.4]
  assign _T_57852 = _T_57851[5:0]; // @[Modules.scala 143:103:@3751.4]
  assign _T_57853 = $signed(_T_57852); // @[Modules.scala 143:103:@3752.4]
  assign _T_57857 = $signed(4'sh1) * $signed(io_in_255); // @[Modules.scala 144:80:@3755.4]
  assign _T_57858 = $signed(_T_54817) + $signed(_T_57857); // @[Modules.scala 143:103:@3756.4]
  assign _T_57859 = _T_57858[5:0]; // @[Modules.scala 143:103:@3757.4]
  assign _T_57860 = $signed(_T_57859); // @[Modules.scala 143:103:@3758.4]
  assign _T_57864 = $signed(4'sh1) * $signed(io_in_257); // @[Modules.scala 144:80:@3761.4]
  assign _T_57865 = $signed(_T_54822) + $signed(_T_57864); // @[Modules.scala 143:103:@3762.4]
  assign _T_57866 = _T_57865[5:0]; // @[Modules.scala 143:103:@3763.4]
  assign _T_57867 = $signed(_T_57866); // @[Modules.scala 143:103:@3764.4]
  assign _T_57869 = $signed(-4'sh1) * $signed(io_in_259); // @[Modules.scala 143:74:@3766.4]
  assign _T_57872 = $signed(_T_57869) + $signed(_T_54831); // @[Modules.scala 143:103:@3768.4]
  assign _T_57873 = _T_57872[4:0]; // @[Modules.scala 143:103:@3769.4]
  assign _T_57874 = $signed(_T_57873); // @[Modules.scala 143:103:@3770.4]
  assign _T_57886 = $signed(_T_54845) + $signed(_T_54850); // @[Modules.scala 143:103:@3780.4]
  assign _T_57887 = _T_57886[5:0]; // @[Modules.scala 143:103:@3781.4]
  assign _T_57888 = $signed(_T_57887); // @[Modules.scala 143:103:@3782.4]
  assign _T_57890 = $signed(4'sh1) * $signed(io_in_268); // @[Modules.scala 143:74:@3784.4]
  assign _T_57892 = $signed(4'sh1) * $signed(io_in_269); // @[Modules.scala 144:80:@3785.4]
  assign _T_57893 = $signed(_T_57890) + $signed(_T_57892); // @[Modules.scala 143:103:@3786.4]
  assign _T_57894 = _T_57893[5:0]; // @[Modules.scala 143:103:@3787.4]
  assign _T_57895 = $signed(_T_57894); // @[Modules.scala 143:103:@3788.4]
  assign _T_57897 = $signed(4'sh1) * $signed(io_in_270); // @[Modules.scala 143:74:@3790.4]
  assign _T_57899 = $signed(4'sh1) * $signed(io_in_271); // @[Modules.scala 144:80:@3791.4]
  assign _T_57900 = $signed(_T_57897) + $signed(_T_57899); // @[Modules.scala 143:103:@3792.4]
  assign _T_57901 = _T_57900[5:0]; // @[Modules.scala 143:103:@3793.4]
  assign _T_57902 = $signed(_T_57901); // @[Modules.scala 143:103:@3794.4]
  assign _T_57904 = $signed(4'sh1) * $signed(io_in_272); // @[Modules.scala 143:74:@3796.4]
  assign _GEN_97 = {{1{_T_54873[4]}},_T_54873}; // @[Modules.scala 143:103:@3798.4]
  assign _T_57907 = $signed(_T_57904) + $signed(_GEN_97); // @[Modules.scala 143:103:@3798.4]
  assign _T_57908 = _T_57907[5:0]; // @[Modules.scala 143:103:@3799.4]
  assign _T_57909 = $signed(_T_57908); // @[Modules.scala 143:103:@3800.4]
  assign _T_57927 = $signed(4'sh1) * $signed(io_in_280); // @[Modules.scala 144:80:@3815.4]
  assign _GEN_98 = {{1{_T_54892[4]}},_T_54892}; // @[Modules.scala 143:103:@3816.4]
  assign _T_57928 = $signed(_GEN_98) + $signed(_T_57927); // @[Modules.scala 143:103:@3816.4]
  assign _T_57929 = _T_57928[5:0]; // @[Modules.scala 143:103:@3817.4]
  assign _T_57930 = $signed(_T_57929); // @[Modules.scala 143:103:@3818.4]
  assign _T_57941 = $signed(4'sh1) * $signed(io_in_284); // @[Modules.scala 144:80:@3827.4]
  assign _T_57942 = $signed(_T_54906) + $signed(_T_57941); // @[Modules.scala 143:103:@3828.4]
  assign _T_57943 = _T_57942[5:0]; // @[Modules.scala 143:103:@3829.4]
  assign _T_57944 = $signed(_T_57943); // @[Modules.scala 143:103:@3830.4]
  assign _T_57949 = $signed(_T_54922) + $signed(_T_54927); // @[Modules.scala 143:103:@3834.4]
  assign _T_57950 = _T_57949[4:0]; // @[Modules.scala 143:103:@3835.4]
  assign _T_57951 = $signed(_T_57950); // @[Modules.scala 143:103:@3836.4]
  assign _T_57956 = $signed(_T_54929) + $signed(_T_54934); // @[Modules.scala 143:103:@3840.4]
  assign _T_57957 = _T_57956[4:0]; // @[Modules.scala 143:103:@3841.4]
  assign _T_57958 = $signed(_T_57957); // @[Modules.scala 143:103:@3842.4]
  assign _T_57962 = $signed(4'sh1) * $signed(io_in_293); // @[Modules.scala 144:80:@3845.4]
  assign _GEN_99 = {{1{_T_54936[4]}},_T_54936}; // @[Modules.scala 143:103:@3846.4]
  assign _T_57963 = $signed(_GEN_99) + $signed(_T_57962); // @[Modules.scala 143:103:@3846.4]
  assign _T_57964 = _T_57963[5:0]; // @[Modules.scala 143:103:@3847.4]
  assign _T_57965 = $signed(_T_57964); // @[Modules.scala 143:103:@3848.4]
  assign _T_57970 = $signed(_T_54943) + $signed(_T_54948); // @[Modules.scala 143:103:@3852.4]
  assign _T_57971 = _T_57970[5:0]; // @[Modules.scala 143:103:@3853.4]
  assign _T_57972 = $signed(_T_57971); // @[Modules.scala 143:103:@3854.4]
  assign _T_57976 = $signed(4'sh1) * $signed(io_in_297); // @[Modules.scala 144:80:@3857.4]
  assign _T_57977 = $signed(_T_54950) + $signed(_T_57976); // @[Modules.scala 143:103:@3858.4]
  assign _T_57978 = _T_57977[5:0]; // @[Modules.scala 143:103:@3859.4]
  assign _T_57979 = $signed(_T_57978); // @[Modules.scala 143:103:@3860.4]
  assign _T_57981 = $signed(4'sh1) * $signed(io_in_298); // @[Modules.scala 143:74:@3862.4]
  assign _T_57983 = $signed(4'sh1) * $signed(io_in_299); // @[Modules.scala 144:80:@3863.4]
  assign _T_57984 = $signed(_T_57981) + $signed(_T_57983); // @[Modules.scala 143:103:@3864.4]
  assign _T_57985 = _T_57984[5:0]; // @[Modules.scala 143:103:@3865.4]
  assign _T_57986 = $signed(_T_57985); // @[Modules.scala 143:103:@3866.4]
  assign _T_57988 = $signed(4'sh1) * $signed(io_in_300); // @[Modules.scala 143:74:@3868.4]
  assign _T_57990 = $signed(4'sh1) * $signed(io_in_301); // @[Modules.scala 144:80:@3869.4]
  assign _T_57991 = $signed(_T_57988) + $signed(_T_57990); // @[Modules.scala 143:103:@3870.4]
  assign _T_57992 = _T_57991[5:0]; // @[Modules.scala 143:103:@3871.4]
  assign _T_57993 = $signed(_T_57992); // @[Modules.scala 143:103:@3872.4]
  assign _T_57998 = $signed(_T_54971) + $signed(_T_54976); // @[Modules.scala 143:103:@3876.4]
  assign _T_57999 = _T_57998[4:0]; // @[Modules.scala 143:103:@3877.4]
  assign _T_58000 = $signed(_T_57999); // @[Modules.scala 143:103:@3878.4]
  assign _T_58005 = $signed(_T_54978) + $signed(_T_54983); // @[Modules.scala 143:103:@3882.4]
  assign _T_58006 = _T_58005[4:0]; // @[Modules.scala 143:103:@3883.4]
  assign _T_58007 = $signed(_T_58006); // @[Modules.scala 143:103:@3884.4]
  assign _T_58009 = $signed(4'sh1) * $signed(io_in_307); // @[Modules.scala 143:74:@3886.4]
  assign _T_58011 = $signed(4'sh1) * $signed(io_in_308); // @[Modules.scala 144:80:@3887.4]
  assign _T_58012 = $signed(_T_58009) + $signed(_T_58011); // @[Modules.scala 143:103:@3888.4]
  assign _T_58013 = _T_58012[5:0]; // @[Modules.scala 143:103:@3889.4]
  assign _T_58014 = $signed(_T_58013); // @[Modules.scala 143:103:@3890.4]
  assign _T_58018 = $signed(4'sh1) * $signed(io_in_310); // @[Modules.scala 144:80:@3893.4]
  assign _T_58019 = $signed(_T_54990) + $signed(_T_58018); // @[Modules.scala 143:103:@3894.4]
  assign _T_58020 = _T_58019[5:0]; // @[Modules.scala 143:103:@3895.4]
  assign _T_58021 = $signed(_T_58020); // @[Modules.scala 143:103:@3896.4]
  assign _T_58025 = $signed(4'sh1) * $signed(io_in_312); // @[Modules.scala 144:80:@3899.4]
  assign _T_58026 = $signed(_T_54997) + $signed(_T_58025); // @[Modules.scala 143:103:@3900.4]
  assign _T_58027 = _T_58026[5:0]; // @[Modules.scala 143:103:@3901.4]
  assign _T_58028 = $signed(_T_58027); // @[Modules.scala 143:103:@3902.4]
  assign _T_58032 = $signed(4'sh1) * $signed(io_in_314); // @[Modules.scala 144:80:@3905.4]
  assign _GEN_100 = {{1{_T_55004[4]}},_T_55004}; // @[Modules.scala 143:103:@3906.4]
  assign _T_58033 = $signed(_GEN_100) + $signed(_T_58032); // @[Modules.scala 143:103:@3906.4]
  assign _T_58034 = _T_58033[5:0]; // @[Modules.scala 143:103:@3907.4]
  assign _T_58035 = $signed(_T_58034); // @[Modules.scala 143:103:@3908.4]
  assign _T_58040 = $signed(_T_55013) + $signed(_T_55018); // @[Modules.scala 143:103:@3912.4]
  assign _T_58041 = _T_58040[4:0]; // @[Modules.scala 143:103:@3913.4]
  assign _T_58042 = $signed(_T_58041); // @[Modules.scala 143:103:@3914.4]
  assign _T_58047 = $signed(_T_55020) + $signed(_T_55025); // @[Modules.scala 143:103:@3918.4]
  assign _T_58048 = _T_58047[4:0]; // @[Modules.scala 143:103:@3919.4]
  assign _T_58049 = $signed(_T_58048); // @[Modules.scala 143:103:@3920.4]
  assign _T_58053 = $signed(4'sh1) * $signed(io_in_321); // @[Modules.scala 144:80:@3923.4]
  assign _GEN_101 = {{1{_T_55027[4]}},_T_55027}; // @[Modules.scala 143:103:@3924.4]
  assign _T_58054 = $signed(_GEN_101) + $signed(_T_58053); // @[Modules.scala 143:103:@3924.4]
  assign _T_58055 = _T_58054[5:0]; // @[Modules.scala 143:103:@3925.4]
  assign _T_58056 = $signed(_T_58055); // @[Modules.scala 143:103:@3926.4]
  assign _T_58058 = $signed(4'sh1) * $signed(io_in_322); // @[Modules.scala 143:74:@3928.4]
  assign _T_58061 = $signed(_T_58058) + $signed(_T_55034); // @[Modules.scala 143:103:@3930.4]
  assign _T_58062 = _T_58061[5:0]; // @[Modules.scala 143:103:@3931.4]
  assign _T_58063 = $signed(_T_58062); // @[Modules.scala 143:103:@3932.4]
  assign _T_58065 = $signed(4'sh1) * $signed(io_in_324); // @[Modules.scala 143:74:@3934.4]
  assign _T_58067 = $signed(4'sh1) * $signed(io_in_325); // @[Modules.scala 144:80:@3935.4]
  assign _T_58068 = $signed(_T_58065) + $signed(_T_58067); // @[Modules.scala 143:103:@3936.4]
  assign _T_58069 = _T_58068[5:0]; // @[Modules.scala 143:103:@3937.4]
  assign _T_58070 = $signed(_T_58069); // @[Modules.scala 143:103:@3938.4]
  assign _T_58072 = $signed(4'sh1) * $signed(io_in_326); // @[Modules.scala 143:74:@3940.4]
  assign _T_58074 = $signed(4'sh1) * $signed(io_in_327); // @[Modules.scala 144:80:@3941.4]
  assign _T_58075 = $signed(_T_58072) + $signed(_T_58074); // @[Modules.scala 143:103:@3942.4]
  assign _T_58076 = _T_58075[5:0]; // @[Modules.scala 143:103:@3943.4]
  assign _T_58077 = $signed(_T_58076); // @[Modules.scala 143:103:@3944.4]
  assign _T_58079 = $signed(4'sh1) * $signed(io_in_328); // @[Modules.scala 143:74:@3946.4]
  assign _T_58081 = $signed(4'sh1) * $signed(io_in_329); // @[Modules.scala 144:80:@3947.4]
  assign _T_58082 = $signed(_T_58079) + $signed(_T_58081); // @[Modules.scala 143:103:@3948.4]
  assign _T_58083 = _T_58082[5:0]; // @[Modules.scala 143:103:@3949.4]
  assign _T_58084 = $signed(_T_58083); // @[Modules.scala 143:103:@3950.4]
  assign _T_58089 = $signed(_T_55062) + $signed(_T_55067); // @[Modules.scala 143:103:@3954.4]
  assign _T_58090 = _T_58089[4:0]; // @[Modules.scala 143:103:@3955.4]
  assign _T_58091 = $signed(_T_58090); // @[Modules.scala 143:103:@3956.4]
  assign _T_58095 = $signed(-4'sh1) * $signed(io_in_334); // @[Modules.scala 144:80:@3959.4]
  assign _T_58096 = $signed(_T_55069) + $signed(_T_58095); // @[Modules.scala 143:103:@3960.4]
  assign _T_58097 = _T_58096[4:0]; // @[Modules.scala 143:103:@3961.4]
  assign _T_58098 = $signed(_T_58097); // @[Modules.scala 143:103:@3962.4]
  assign _T_58100 = $signed(4'sh1) * $signed(io_in_335); // @[Modules.scala 143:74:@3964.4]
  assign _T_58102 = $signed(4'sh1) * $signed(io_in_336); // @[Modules.scala 144:80:@3965.4]
  assign _T_58103 = $signed(_T_58100) + $signed(_T_58102); // @[Modules.scala 143:103:@3966.4]
  assign _T_58104 = _T_58103[5:0]; // @[Modules.scala 143:103:@3967.4]
  assign _T_58105 = $signed(_T_58104); // @[Modules.scala 143:103:@3968.4]
  assign _T_58107 = $signed(-4'sh1) * $signed(io_in_337); // @[Modules.scala 143:74:@3970.4]
  assign _T_58109 = $signed(-4'sh1) * $signed(io_in_338); // @[Modules.scala 144:80:@3971.4]
  assign _T_58110 = $signed(_T_58107) + $signed(_T_58109); // @[Modules.scala 143:103:@3972.4]
  assign _T_58111 = _T_58110[4:0]; // @[Modules.scala 143:103:@3973.4]
  assign _T_58112 = $signed(_T_58111); // @[Modules.scala 143:103:@3974.4]
  assign _T_58116 = $signed(4'sh1) * $signed(io_in_340); // @[Modules.scala 144:80:@3977.4]
  assign _T_58117 = $signed(_T_55083) + $signed(_T_58116); // @[Modules.scala 143:103:@3978.4]
  assign _T_58118 = _T_58117[5:0]; // @[Modules.scala 143:103:@3979.4]
  assign _T_58119 = $signed(_T_58118); // @[Modules.scala 143:103:@3980.4]
  assign _T_58121 = $signed(4'sh1) * $signed(io_in_341); // @[Modules.scala 143:74:@3982.4]
  assign _GEN_102 = {{1{_T_55102[4]}},_T_55102}; // @[Modules.scala 143:103:@3984.4]
  assign _T_58124 = $signed(_T_58121) + $signed(_GEN_102); // @[Modules.scala 143:103:@3984.4]
  assign _T_58125 = _T_58124[5:0]; // @[Modules.scala 143:103:@3985.4]
  assign _T_58126 = $signed(_T_58125); // @[Modules.scala 143:103:@3986.4]
  assign _T_58131 = $signed(_T_55104) + $signed(_T_55109); // @[Modules.scala 143:103:@3990.4]
  assign _T_58132 = _T_58131[4:0]; // @[Modules.scala 143:103:@3991.4]
  assign _T_58133 = $signed(_T_58132); // @[Modules.scala 143:103:@3992.4]
  assign _T_58138 = $signed(_T_55111) + $signed(_T_55116); // @[Modules.scala 143:103:@3996.4]
  assign _T_58139 = _T_58138[4:0]; // @[Modules.scala 143:103:@3997.4]
  assign _T_58140 = $signed(_T_58139); // @[Modules.scala 143:103:@3998.4]
  assign _T_58142 = $signed(4'sh1) * $signed(io_in_349); // @[Modules.scala 143:74:@4000.4]
  assign _T_58145 = $signed(_T_58142) + $signed(_T_55123); // @[Modules.scala 143:103:@4002.4]
  assign _T_58146 = _T_58145[5:0]; // @[Modules.scala 143:103:@4003.4]
  assign _T_58147 = $signed(_T_58146); // @[Modules.scala 143:103:@4004.4]
  assign _T_58151 = $signed(4'sh1) * $signed(io_in_352); // @[Modules.scala 144:80:@4007.4]
  assign _T_58152 = $signed(_T_55125) + $signed(_T_58151); // @[Modules.scala 143:103:@4008.4]
  assign _T_58153 = _T_58152[5:0]; // @[Modules.scala 143:103:@4009.4]
  assign _T_58154 = $signed(_T_58153); // @[Modules.scala 143:103:@4010.4]
  assign _T_58156 = $signed(4'sh1) * $signed(io_in_353); // @[Modules.scala 143:74:@4012.4]
  assign _T_58158 = $signed(4'sh1) * $signed(io_in_354); // @[Modules.scala 144:80:@4013.4]
  assign _T_58159 = $signed(_T_58156) + $signed(_T_58158); // @[Modules.scala 143:103:@4014.4]
  assign _T_58160 = _T_58159[5:0]; // @[Modules.scala 143:103:@4015.4]
  assign _T_58161 = $signed(_T_58160); // @[Modules.scala 143:103:@4016.4]
  assign _T_58163 = $signed(4'sh1) * $signed(io_in_355); // @[Modules.scala 143:74:@4018.4]
  assign _T_58166 = $signed(_T_58163) + $signed(_T_55137); // @[Modules.scala 143:103:@4020.4]
  assign _T_58167 = _T_58166[5:0]; // @[Modules.scala 143:103:@4021.4]
  assign _T_58168 = $signed(_T_58167); // @[Modules.scala 143:103:@4022.4]
  assign _T_58170 = $signed(4'sh1) * $signed(io_in_357); // @[Modules.scala 143:74:@4024.4]
  assign _T_58172 = $signed(-4'sh1) * $signed(io_in_360); // @[Modules.scala 144:80:@4025.4]
  assign _GEN_103 = {{1{_T_58172[4]}},_T_58172}; // @[Modules.scala 143:103:@4026.4]
  assign _T_58173 = $signed(_T_58170) + $signed(_GEN_103); // @[Modules.scala 143:103:@4026.4]
  assign _T_58174 = _T_58173[5:0]; // @[Modules.scala 143:103:@4027.4]
  assign _T_58175 = $signed(_T_58174); // @[Modules.scala 143:103:@4028.4]
  assign _T_58177 = $signed(4'sh1) * $signed(io_in_361); // @[Modules.scala 143:74:@4030.4]
  assign _T_58180 = $signed(_T_58177) + $signed(_GEN_32); // @[Modules.scala 143:103:@4032.4]
  assign _T_58181 = _T_58180[5:0]; // @[Modules.scala 143:103:@4033.4]
  assign _T_58182 = $signed(_T_58181); // @[Modules.scala 143:103:@4034.4]
  assign _T_58187 = $signed(_T_55160) + $signed(_T_55165); // @[Modules.scala 143:103:@4038.4]
  assign _T_58188 = _T_58187[5:0]; // @[Modules.scala 143:103:@4039.4]
  assign _T_58189 = $signed(_T_58188); // @[Modules.scala 143:103:@4040.4]
  assign _T_58191 = $signed(-4'sh1) * $signed(io_in_365); // @[Modules.scala 143:74:@4042.4]
  assign _T_58193 = $signed(-4'sh1) * $signed(io_in_366); // @[Modules.scala 144:80:@4043.4]
  assign _T_58194 = $signed(_T_58191) + $signed(_T_58193); // @[Modules.scala 143:103:@4044.4]
  assign _T_58195 = _T_58194[4:0]; // @[Modules.scala 143:103:@4045.4]
  assign _T_58196 = $signed(_T_58195); // @[Modules.scala 143:103:@4046.4]
  assign _T_58200 = $signed(4'sh1) * $signed(io_in_368); // @[Modules.scala 144:80:@4049.4]
  assign _T_58201 = $signed(_T_55174) + $signed(_T_58200); // @[Modules.scala 143:103:@4050.4]
  assign _T_58202 = _T_58201[5:0]; // @[Modules.scala 143:103:@4051.4]
  assign _T_58203 = $signed(_T_58202); // @[Modules.scala 143:103:@4052.4]
  assign _T_58205 = $signed(4'sh1) * $signed(io_in_369); // @[Modules.scala 143:74:@4054.4]
  assign _T_58207 = $signed(4'sh1) * $signed(io_in_370); // @[Modules.scala 144:80:@4055.4]
  assign _T_58208 = $signed(_T_58205) + $signed(_T_58207); // @[Modules.scala 143:103:@4056.4]
  assign _T_58209 = _T_58208[5:0]; // @[Modules.scala 143:103:@4057.4]
  assign _T_58210 = $signed(_T_58209); // @[Modules.scala 143:103:@4058.4]
  assign _T_58212 = $signed(4'sh1) * $signed(io_in_372); // @[Modules.scala 143:74:@4060.4]
  assign _GEN_105 = {{1{_T_55200[4]}},_T_55200}; // @[Modules.scala 143:103:@4062.4]
  assign _T_58215 = $signed(_T_58212) + $signed(_GEN_105); // @[Modules.scala 143:103:@4062.4]
  assign _T_58216 = _T_58215[5:0]; // @[Modules.scala 143:103:@4063.4]
  assign _T_58217 = $signed(_T_58216); // @[Modules.scala 143:103:@4064.4]
  assign _T_58222 = $signed(_T_55202) + $signed(_T_55207); // @[Modules.scala 143:103:@4068.4]
  assign _T_58223 = _T_58222[4:0]; // @[Modules.scala 143:103:@4069.4]
  assign _T_58224 = $signed(_T_58223); // @[Modules.scala 143:103:@4070.4]
  assign _T_58226 = $signed(4'sh1) * $signed(io_in_377); // @[Modules.scala 143:74:@4072.4]
  assign _T_58229 = $signed(_T_58226) + $signed(_T_55214); // @[Modules.scala 143:103:@4074.4]
  assign _T_58230 = _T_58229[5:0]; // @[Modules.scala 143:103:@4075.4]
  assign _T_58231 = $signed(_T_58230); // @[Modules.scala 143:103:@4076.4]
  assign _T_58233 = $signed(4'sh1) * $signed(io_in_379); // @[Modules.scala 143:74:@4078.4]
  assign _T_58235 = $signed(4'sh1) * $signed(io_in_380); // @[Modules.scala 144:80:@4079.4]
  assign _T_58236 = $signed(_T_58233) + $signed(_T_58235); // @[Modules.scala 143:103:@4080.4]
  assign _T_58237 = _T_58236[5:0]; // @[Modules.scala 143:103:@4081.4]
  assign _T_58238 = $signed(_T_58237); // @[Modules.scala 143:103:@4082.4]
  assign _T_58240 = $signed(4'sh1) * $signed(io_in_381); // @[Modules.scala 143:74:@4084.4]
  assign _T_58243 = $signed(_T_58240) + $signed(_T_55221); // @[Modules.scala 143:103:@4086.4]
  assign _T_58244 = _T_58243[5:0]; // @[Modules.scala 143:103:@4087.4]
  assign _T_58245 = $signed(_T_58244); // @[Modules.scala 143:103:@4088.4]
  assign _T_58247 = $signed(4'sh1) * $signed(io_in_383); // @[Modules.scala 143:74:@4090.4]
  assign _T_58249 = $signed(4'sh1) * $signed(io_in_384); // @[Modules.scala 144:80:@4091.4]
  assign _T_58250 = $signed(_T_58247) + $signed(_T_58249); // @[Modules.scala 143:103:@4092.4]
  assign _T_58251 = _T_58250[5:0]; // @[Modules.scala 143:103:@4093.4]
  assign _T_58252 = $signed(_T_58251); // @[Modules.scala 143:103:@4094.4]
  assign _T_58254 = $signed(-4'sh1) * $signed(io_in_385); // @[Modules.scala 143:74:@4096.4]
  assign _T_58257 = $signed(_T_58254) + $signed(_T_55228); // @[Modules.scala 143:103:@4098.4]
  assign _T_58258 = _T_58257[4:0]; // @[Modules.scala 143:103:@4099.4]
  assign _T_58259 = $signed(_T_58258); // @[Modules.scala 143:103:@4100.4]
  assign _T_58261 = $signed(-4'sh1) * $signed(io_in_387); // @[Modules.scala 143:74:@4102.4]
  assign _T_58263 = $signed(-4'sh1) * $signed(io_in_388); // @[Modules.scala 144:80:@4103.4]
  assign _T_58264 = $signed(_T_58261) + $signed(_T_58263); // @[Modules.scala 143:103:@4104.4]
  assign _T_58265 = _T_58264[4:0]; // @[Modules.scala 143:103:@4105.4]
  assign _T_58266 = $signed(_T_58265); // @[Modules.scala 143:103:@4106.4]
  assign _T_58268 = $signed(4'sh1) * $signed(io_in_389); // @[Modules.scala 143:74:@4108.4]
  assign _T_58270 = $signed(4'sh1) * $signed(io_in_390); // @[Modules.scala 144:80:@4109.4]
  assign _T_58271 = $signed(_T_58268) + $signed(_T_58270); // @[Modules.scala 143:103:@4110.4]
  assign _T_58272 = _T_58271[5:0]; // @[Modules.scala 143:103:@4111.4]
  assign _T_58273 = $signed(_T_58272); // @[Modules.scala 143:103:@4112.4]
  assign _T_58277 = $signed(-4'sh1) * $signed(io_in_392); // @[Modules.scala 144:80:@4115.4]
  assign _GEN_106 = {{1{_T_58277[4]}},_T_58277}; // @[Modules.scala 143:103:@4116.4]
  assign _T_58278 = $signed(_T_55244) + $signed(_GEN_106); // @[Modules.scala 143:103:@4116.4]
  assign _T_58279 = _T_58278[5:0]; // @[Modules.scala 143:103:@4117.4]
  assign _T_58280 = $signed(_T_58279); // @[Modules.scala 143:103:@4118.4]
  assign _T_58282 = $signed(4'sh1) * $signed(io_in_393); // @[Modules.scala 143:74:@4120.4]
  assign _T_58285 = $signed(_T_58282) + $signed(_T_55258); // @[Modules.scala 143:103:@4122.4]
  assign _T_58286 = _T_58285[5:0]; // @[Modules.scala 143:103:@4123.4]
  assign _T_58287 = $signed(_T_58286); // @[Modules.scala 143:103:@4124.4]
  assign _T_58289 = $signed(4'sh1) * $signed(io_in_396); // @[Modules.scala 143:74:@4126.4]
  assign _T_58291 = $signed(4'sh1) * $signed(io_in_397); // @[Modules.scala 144:80:@4127.4]
  assign _T_58292 = $signed(_T_58289) + $signed(_T_58291); // @[Modules.scala 143:103:@4128.4]
  assign _T_58293 = _T_58292[5:0]; // @[Modules.scala 143:103:@4129.4]
  assign _T_58294 = $signed(_T_58293); // @[Modules.scala 143:103:@4130.4]
  assign _T_58296 = $signed(4'sh1) * $signed(io_in_400); // @[Modules.scala 143:74:@4132.4]
  assign _GEN_107 = {{1{_T_55284[4]}},_T_55284}; // @[Modules.scala 143:103:@4134.4]
  assign _T_58299 = $signed(_T_58296) + $signed(_GEN_107); // @[Modules.scala 143:103:@4134.4]
  assign _T_58300 = _T_58299[5:0]; // @[Modules.scala 143:103:@4135.4]
  assign _T_58301 = $signed(_T_58300); // @[Modules.scala 143:103:@4136.4]
  assign _T_58306 = $signed(_T_55286) + $signed(_T_55291); // @[Modules.scala 143:103:@4140.4]
  assign _T_58307 = _T_58306[4:0]; // @[Modules.scala 143:103:@4141.4]
  assign _T_58308 = $signed(_T_58307); // @[Modules.scala 143:103:@4142.4]
  assign _T_58310 = $signed(4'sh1) * $signed(io_in_405); // @[Modules.scala 143:74:@4144.4]
  assign _T_58313 = $signed(_T_58310) + $signed(_T_55293); // @[Modules.scala 143:103:@4146.4]
  assign _T_58314 = _T_58313[5:0]; // @[Modules.scala 143:103:@4147.4]
  assign _T_58315 = $signed(_T_58314); // @[Modules.scala 143:103:@4148.4]
  assign _T_58326 = $signed(-4'sh1) * $signed(io_in_412); // @[Modules.scala 144:80:@4157.4]
  assign _T_58327 = $signed(_T_55305) + $signed(_T_58326); // @[Modules.scala 143:103:@4158.4]
  assign _T_58328 = _T_58327[4:0]; // @[Modules.scala 143:103:@4159.4]
  assign _T_58329 = $signed(_T_58328); // @[Modules.scala 143:103:@4160.4]
  assign _T_58331 = $signed(-4'sh1) * $signed(io_in_413); // @[Modules.scala 143:74:@4162.4]
  assign _T_58333 = $signed(-4'sh1) * $signed(io_in_414); // @[Modules.scala 144:80:@4163.4]
  assign _T_58334 = $signed(_T_58331) + $signed(_T_58333); // @[Modules.scala 143:103:@4164.4]
  assign _T_58335 = _T_58334[4:0]; // @[Modules.scala 143:103:@4165.4]
  assign _T_58336 = $signed(_T_58335); // @[Modules.scala 143:103:@4166.4]
  assign _T_58338 = $signed(-4'sh1) * $signed(io_in_415); // @[Modules.scala 143:74:@4168.4]
  assign _T_58340 = $signed(-4'sh1) * $signed(io_in_416); // @[Modules.scala 144:80:@4169.4]
  assign _T_58341 = $signed(_T_58338) + $signed(_T_58340); // @[Modules.scala 143:103:@4170.4]
  assign _T_58342 = _T_58341[4:0]; // @[Modules.scala 143:103:@4171.4]
  assign _T_58343 = $signed(_T_58342); // @[Modules.scala 143:103:@4172.4]
  assign _T_58347 = $signed(-4'sh1) * $signed(io_in_418); // @[Modules.scala 144:80:@4175.4]
  assign _T_58348 = $signed(_T_55321) + $signed(_T_58347); // @[Modules.scala 143:103:@4176.4]
  assign _T_58349 = _T_58348[4:0]; // @[Modules.scala 143:103:@4177.4]
  assign _T_58350 = $signed(_T_58349); // @[Modules.scala 143:103:@4178.4]
  assign _T_58352 = $signed(-4'sh1) * $signed(io_in_420); // @[Modules.scala 143:74:@4180.4]
  assign _T_58355 = $signed(_T_58352) + $signed(_T_55333); // @[Modules.scala 143:103:@4182.4]
  assign _T_58356 = _T_58355[4:0]; // @[Modules.scala 143:103:@4183.4]
  assign _T_58357 = $signed(_T_58356); // @[Modules.scala 143:103:@4184.4]
  assign _T_58361 = $signed(4'sh1) * $signed(io_in_424); // @[Modules.scala 144:80:@4187.4]
  assign _T_58362 = $signed(_T_55340) + $signed(_T_58361); // @[Modules.scala 143:103:@4188.4]
  assign _T_58363 = _T_58362[5:0]; // @[Modules.scala 143:103:@4189.4]
  assign _T_58364 = $signed(_T_58363); // @[Modules.scala 143:103:@4190.4]
  assign _T_58375 = $signed(-4'sh1) * $signed(io_in_428); // @[Modules.scala 144:80:@4199.4]
  assign _T_58376 = $signed(_T_55354) + $signed(_T_58375); // @[Modules.scala 143:103:@4200.4]
  assign _T_58377 = _T_58376[4:0]; // @[Modules.scala 143:103:@4201.4]
  assign _T_58378 = $signed(_T_58377); // @[Modules.scala 143:103:@4202.4]
  assign _T_58382 = $signed(-4'sh1) * $signed(io_in_431); // @[Modules.scala 144:80:@4205.4]
  assign _T_58383 = $signed(_T_55361) + $signed(_T_58382); // @[Modules.scala 143:103:@4206.4]
  assign _T_58384 = _T_58383[4:0]; // @[Modules.scala 143:103:@4207.4]
  assign _T_58385 = $signed(_T_58384); // @[Modules.scala 143:103:@4208.4]
  assign _T_58387 = $signed(-4'sh1) * $signed(io_in_432); // @[Modules.scala 143:74:@4210.4]
  assign _GEN_109 = {{1{_T_58387[4]}},_T_58387}; // @[Modules.scala 143:103:@4212.4]
  assign _T_58390 = $signed(_GEN_109) + $signed(_T_55368); // @[Modules.scala 143:103:@4212.4]
  assign _T_58391 = _T_58390[5:0]; // @[Modules.scala 143:103:@4213.4]
  assign _T_58392 = $signed(_T_58391); // @[Modules.scala 143:103:@4214.4]
  assign _T_58397 = $signed(_T_55370) + $signed(_GEN_47); // @[Modules.scala 143:103:@4218.4]
  assign _T_58398 = _T_58397[5:0]; // @[Modules.scala 143:103:@4219.4]
  assign _T_58399 = $signed(_T_58398); // @[Modules.scala 143:103:@4220.4]
  assign _T_58401 = $signed(-4'sh1) * $signed(io_in_441); // @[Modules.scala 143:74:@4222.4]
  assign _T_58403 = $signed(4'sh1) * $signed(io_in_442); // @[Modules.scala 144:80:@4223.4]
  assign _GEN_111 = {{1{_T_58401[4]}},_T_58401}; // @[Modules.scala 143:103:@4224.4]
  assign _T_58404 = $signed(_GEN_111) + $signed(_T_58403); // @[Modules.scala 143:103:@4224.4]
  assign _T_58405 = _T_58404[5:0]; // @[Modules.scala 143:103:@4225.4]
  assign _T_58406 = $signed(_T_58405); // @[Modules.scala 143:103:@4226.4]
  assign _T_58410 = $signed(-4'sh1) * $signed(io_in_444); // @[Modules.scala 144:80:@4229.4]
  assign _T_58411 = $signed(_T_55403) + $signed(_T_58410); // @[Modules.scala 143:103:@4230.4]
  assign _T_58412 = _T_58411[4:0]; // @[Modules.scala 143:103:@4231.4]
  assign _T_58413 = $signed(_T_58412); // @[Modules.scala 143:103:@4232.4]
  assign _T_58415 = $signed(-4'sh1) * $signed(io_in_445); // @[Modules.scala 143:74:@4234.4]
  assign _T_58417 = $signed(-4'sh1) * $signed(io_in_446); // @[Modules.scala 144:80:@4235.4]
  assign _T_58418 = $signed(_T_58415) + $signed(_T_58417); // @[Modules.scala 143:103:@4236.4]
  assign _T_58419 = _T_58418[4:0]; // @[Modules.scala 143:103:@4237.4]
  assign _T_58420 = $signed(_T_58419); // @[Modules.scala 143:103:@4238.4]
  assign _T_58424 = $signed(4'sh1) * $signed(io_in_448); // @[Modules.scala 144:80:@4241.4]
  assign _T_58425 = $signed(_T_55412) + $signed(_T_58424); // @[Modules.scala 143:103:@4242.4]
  assign _T_58426 = _T_58425[5:0]; // @[Modules.scala 143:103:@4243.4]
  assign _T_58427 = $signed(_T_58426); // @[Modules.scala 143:103:@4244.4]
  assign _GEN_112 = {{1{_T_55419[4]}},_T_55419}; // @[Modules.scala 143:103:@4248.4]
  assign _T_58432 = $signed(_GEN_112) + $signed(_T_55424); // @[Modules.scala 143:103:@4248.4]
  assign _T_58433 = _T_58432[5:0]; // @[Modules.scala 143:103:@4249.4]
  assign _T_58434 = $signed(_T_58433); // @[Modules.scala 143:103:@4250.4]
  assign _T_58438 = $signed(4'sh1) * $signed(io_in_452); // @[Modules.scala 144:80:@4253.4]
  assign _T_58439 = $signed(_T_55426) + $signed(_T_58438); // @[Modules.scala 143:103:@4254.4]
  assign _T_58440 = _T_58439[5:0]; // @[Modules.scala 143:103:@4255.4]
  assign _T_58441 = $signed(_T_58440); // @[Modules.scala 143:103:@4256.4]
  assign _T_58445 = $signed(-4'sh1) * $signed(io_in_454); // @[Modules.scala 144:80:@4259.4]
  assign _T_58446 = $signed(_T_55433) + $signed(_T_58445); // @[Modules.scala 143:103:@4260.4]
  assign _T_58447 = _T_58446[4:0]; // @[Modules.scala 143:103:@4261.4]
  assign _T_58448 = $signed(_T_58447); // @[Modules.scala 143:103:@4262.4]
  assign _T_58450 = $signed(-4'sh1) * $signed(io_in_455); // @[Modules.scala 143:74:@4264.4]
  assign _T_58452 = $signed(-4'sh1) * $signed(io_in_456); // @[Modules.scala 144:80:@4265.4]
  assign _T_58453 = $signed(_T_58450) + $signed(_T_58452); // @[Modules.scala 143:103:@4266.4]
  assign _T_58454 = _T_58453[4:0]; // @[Modules.scala 143:103:@4267.4]
  assign _T_58455 = $signed(_T_58454); // @[Modules.scala 143:103:@4268.4]
  assign _T_58457 = $signed(-4'sh1) * $signed(io_in_457); // @[Modules.scala 143:74:@4270.4]
  assign _T_58459 = $signed(-4'sh1) * $signed(io_in_458); // @[Modules.scala 144:80:@4271.4]
  assign _T_58460 = $signed(_T_58457) + $signed(_T_58459); // @[Modules.scala 143:103:@4272.4]
  assign _T_58461 = _T_58460[4:0]; // @[Modules.scala 143:103:@4273.4]
  assign _T_58462 = $signed(_T_58461); // @[Modules.scala 143:103:@4274.4]
  assign _T_58464 = $signed(-4'sh1) * $signed(io_in_459); // @[Modules.scala 143:74:@4276.4]
  assign _T_58466 = $signed(-4'sh1) * $signed(io_in_460); // @[Modules.scala 144:80:@4277.4]
  assign _T_58467 = $signed(_T_58464) + $signed(_T_58466); // @[Modules.scala 143:103:@4278.4]
  assign _T_58468 = _T_58467[4:0]; // @[Modules.scala 143:103:@4279.4]
  assign _T_58469 = $signed(_T_58468); // @[Modules.scala 143:103:@4280.4]
  assign _T_58471 = $signed(-4'sh1) * $signed(io_in_463); // @[Modules.scala 143:74:@4282.4]
  assign _T_58473 = $signed(-4'sh1) * $signed(io_in_464); // @[Modules.scala 144:80:@4283.4]
  assign _T_58474 = $signed(_T_58471) + $signed(_T_58473); // @[Modules.scala 143:103:@4284.4]
  assign _T_58475 = _T_58474[4:0]; // @[Modules.scala 143:103:@4285.4]
  assign _T_58476 = $signed(_T_58475); // @[Modules.scala 143:103:@4286.4]
  assign _T_58478 = $signed(4'sh1) * $signed(io_in_465); // @[Modules.scala 143:74:@4288.4]
  assign _T_58480 = $signed(4'sh1) * $signed(io_in_466); // @[Modules.scala 144:80:@4289.4]
  assign _T_58481 = $signed(_T_58478) + $signed(_T_58480); // @[Modules.scala 143:103:@4290.4]
  assign _T_58482 = _T_58481[5:0]; // @[Modules.scala 143:103:@4291.4]
  assign _T_58483 = $signed(_T_58482); // @[Modules.scala 143:103:@4292.4]
  assign _T_58485 = $signed(4'sh1) * $signed(io_in_470); // @[Modules.scala 143:74:@4294.4]
  assign _T_58488 = $signed(_T_58485) + $signed(_GEN_52); // @[Modules.scala 143:103:@4296.4]
  assign _T_58489 = _T_58488[5:0]; // @[Modules.scala 143:103:@4297.4]
  assign _T_58490 = $signed(_T_58489); // @[Modules.scala 143:103:@4298.4]
  assign _T_58492 = $signed(-4'sh1) * $signed(io_in_472); // @[Modules.scala 143:74:@4300.4]
  assign _T_58494 = $signed(-4'sh1) * $signed(io_in_473); // @[Modules.scala 144:80:@4301.4]
  assign _T_58495 = $signed(_T_58492) + $signed(_T_58494); // @[Modules.scala 143:103:@4302.4]
  assign _T_58496 = _T_58495[4:0]; // @[Modules.scala 143:103:@4303.4]
  assign _T_58497 = $signed(_T_58496); // @[Modules.scala 143:103:@4304.4]
  assign _T_58501 = $signed(4'sh1) * $signed(io_in_475); // @[Modules.scala 144:80:@4307.4]
  assign _T_58502 = $signed(_T_55482) + $signed(_T_58501); // @[Modules.scala 143:103:@4308.4]
  assign _T_58503 = _T_58502[5:0]; // @[Modules.scala 143:103:@4309.4]
  assign _T_58504 = $signed(_T_58503); // @[Modules.scala 143:103:@4310.4]
  assign _T_58520 = $signed(-4'sh1) * $signed(io_in_481); // @[Modules.scala 143:74:@4324.4]
  assign _T_58522 = $signed(-4'sh1) * $signed(io_in_482); // @[Modules.scala 144:80:@4325.4]
  assign _T_58523 = $signed(_T_58520) + $signed(_T_58522); // @[Modules.scala 143:103:@4326.4]
  assign _T_58524 = _T_58523[4:0]; // @[Modules.scala 143:103:@4327.4]
  assign _T_58525 = $signed(_T_58524); // @[Modules.scala 143:103:@4328.4]
  assign _T_58527 = $signed(-4'sh1) * $signed(io_in_483); // @[Modules.scala 143:74:@4330.4]
  assign _T_58529 = $signed(-4'sh1) * $signed(io_in_484); // @[Modules.scala 144:80:@4331.4]
  assign _T_58530 = $signed(_T_58527) + $signed(_T_58529); // @[Modules.scala 143:103:@4332.4]
  assign _T_58531 = _T_58530[4:0]; // @[Modules.scala 143:103:@4333.4]
  assign _T_58532 = $signed(_T_58531); // @[Modules.scala 143:103:@4334.4]
  assign _T_58536 = $signed(-4'sh1) * $signed(io_in_486); // @[Modules.scala 144:80:@4337.4]
  assign _T_58537 = $signed(_T_55503) + $signed(_T_58536); // @[Modules.scala 143:103:@4338.4]
  assign _T_58538 = _T_58537[4:0]; // @[Modules.scala 143:103:@4339.4]
  assign _T_58539 = $signed(_T_58538); // @[Modules.scala 143:103:@4340.4]
  assign _T_58541 = $signed(-4'sh1) * $signed(io_in_487); // @[Modules.scala 143:74:@4342.4]
  assign _T_58543 = $signed(-4'sh1) * $signed(io_in_488); // @[Modules.scala 144:80:@4343.4]
  assign _T_58544 = $signed(_T_58541) + $signed(_T_58543); // @[Modules.scala 143:103:@4344.4]
  assign _T_58545 = _T_58544[4:0]; // @[Modules.scala 143:103:@4345.4]
  assign _T_58546 = $signed(_T_58545); // @[Modules.scala 143:103:@4346.4]
  assign _T_58548 = $signed(-4'sh1) * $signed(io_in_490); // @[Modules.scala 143:74:@4348.4]
  assign _T_58550 = $signed(-4'sh1) * $signed(io_in_491); // @[Modules.scala 144:80:@4349.4]
  assign _T_58551 = $signed(_T_58548) + $signed(_T_58550); // @[Modules.scala 143:103:@4350.4]
  assign _T_58552 = _T_58551[4:0]; // @[Modules.scala 143:103:@4351.4]
  assign _T_58553 = $signed(_T_58552); // @[Modules.scala 143:103:@4352.4]
  assign _T_58557 = $signed(4'sh1) * $signed(io_in_494); // @[Modules.scala 144:80:@4355.4]
  assign _GEN_115 = {{1{_T_55529[4]}},_T_55529}; // @[Modules.scala 143:103:@4356.4]
  assign _T_58558 = $signed(_GEN_115) + $signed(_T_58557); // @[Modules.scala 143:103:@4356.4]
  assign _T_58559 = _T_58558[5:0]; // @[Modules.scala 143:103:@4357.4]
  assign _T_58560 = $signed(_T_58559); // @[Modules.scala 143:103:@4358.4]
  assign _T_58562 = $signed(-4'sh1) * $signed(io_in_495); // @[Modules.scala 143:74:@4360.4]
  assign _T_58564 = $signed(-4'sh1) * $signed(io_in_496); // @[Modules.scala 144:80:@4361.4]
  assign _T_58565 = $signed(_T_58562) + $signed(_T_58564); // @[Modules.scala 143:103:@4362.4]
  assign _T_58566 = _T_58565[4:0]; // @[Modules.scala 143:103:@4363.4]
  assign _T_58567 = $signed(_T_58566); // @[Modules.scala 143:103:@4364.4]
  assign _T_58569 = $signed(4'sh1) * $signed(io_in_498); // @[Modules.scala 143:74:@4366.4]
  assign _T_58571 = $signed(-4'sh1) * $signed(io_in_499); // @[Modules.scala 144:80:@4367.4]
  assign _GEN_116 = {{1{_T_58571[4]}},_T_58571}; // @[Modules.scala 143:103:@4368.4]
  assign _T_58572 = $signed(_T_58569) + $signed(_GEN_116); // @[Modules.scala 143:103:@4368.4]
  assign _T_58573 = _T_58572[5:0]; // @[Modules.scala 143:103:@4369.4]
  assign _T_58574 = $signed(_T_58573); // @[Modules.scala 143:103:@4370.4]
  assign _T_58576 = $signed(-4'sh1) * $signed(io_in_500); // @[Modules.scala 143:74:@4372.4]
  assign _T_58578 = $signed(-4'sh1) * $signed(io_in_501); // @[Modules.scala 144:80:@4373.4]
  assign _T_58579 = $signed(_T_58576) + $signed(_T_58578); // @[Modules.scala 143:103:@4374.4]
  assign _T_58580 = _T_58579[4:0]; // @[Modules.scala 143:103:@4375.4]
  assign _T_58581 = $signed(_T_58580); // @[Modules.scala 143:103:@4376.4]
  assign _T_58586 = $signed(_T_55552) + $signed(_T_55557); // @[Modules.scala 143:103:@4380.4]
  assign _T_58587 = _T_58586[5:0]; // @[Modules.scala 143:103:@4381.4]
  assign _T_58588 = $signed(_T_58587); // @[Modules.scala 143:103:@4382.4]
  assign _T_58590 = $signed(4'sh1) * $signed(io_in_504); // @[Modules.scala 143:74:@4384.4]
  assign _T_58593 = $signed(_T_58590) + $signed(_T_55566); // @[Modules.scala 143:103:@4386.4]
  assign _T_58594 = _T_58593[5:0]; // @[Modules.scala 143:103:@4387.4]
  assign _T_58595 = $signed(_T_58594); // @[Modules.scala 143:103:@4388.4]
  assign _T_58599 = $signed(-4'sh1) * $signed(io_in_509); // @[Modules.scala 144:80:@4391.4]
  assign _GEN_117 = {{1{_T_58599[4]}},_T_58599}; // @[Modules.scala 143:103:@4392.4]
  assign _T_58600 = $signed(_T_55571) + $signed(_GEN_117); // @[Modules.scala 143:103:@4392.4]
  assign _T_58601 = _T_58600[5:0]; // @[Modules.scala 143:103:@4393.4]
  assign _T_58602 = $signed(_T_58601); // @[Modules.scala 143:103:@4394.4]
  assign _T_58606 = $signed(-4'sh1) * $signed(io_in_511); // @[Modules.scala 144:80:@4397.4]
  assign _T_58607 = $signed(_T_55580) + $signed(_T_58606); // @[Modules.scala 143:103:@4398.4]
  assign _T_58608 = _T_58607[4:0]; // @[Modules.scala 143:103:@4399.4]
  assign _T_58609 = $signed(_T_58608); // @[Modules.scala 143:103:@4400.4]
  assign _T_58613 = $signed(-4'sh1) * $signed(io_in_513); // @[Modules.scala 144:80:@4403.4]
  assign _T_58614 = $signed(_T_55585) + $signed(_T_58613); // @[Modules.scala 143:103:@4404.4]
  assign _T_58615 = _T_58614[4:0]; // @[Modules.scala 143:103:@4405.4]
  assign _T_58616 = $signed(_T_58615); // @[Modules.scala 143:103:@4406.4]
  assign _T_58618 = $signed(-4'sh1) * $signed(io_in_514); // @[Modules.scala 143:74:@4408.4]
  assign _T_58620 = $signed(-4'sh1) * $signed(io_in_515); // @[Modules.scala 144:80:@4409.4]
  assign _T_58621 = $signed(_T_58618) + $signed(_T_58620); // @[Modules.scala 143:103:@4410.4]
  assign _T_58622 = _T_58621[4:0]; // @[Modules.scala 143:103:@4411.4]
  assign _T_58623 = $signed(_T_58622); // @[Modules.scala 143:103:@4412.4]
  assign _T_58625 = $signed(-4'sh1) * $signed(io_in_516); // @[Modules.scala 143:74:@4414.4]
  assign _T_58627 = $signed(-4'sh1) * $signed(io_in_517); // @[Modules.scala 144:80:@4415.4]
  assign _T_58628 = $signed(_T_58625) + $signed(_T_58627); // @[Modules.scala 143:103:@4416.4]
  assign _T_58629 = _T_58628[4:0]; // @[Modules.scala 143:103:@4417.4]
  assign _T_58630 = $signed(_T_58629); // @[Modules.scala 143:103:@4418.4]
  assign _T_58632 = $signed(4'sh1) * $signed(io_in_519); // @[Modules.scala 143:74:@4420.4]
  assign _T_58635 = $signed(_T_58632) + $signed(_GEN_60); // @[Modules.scala 143:103:@4422.4]
  assign _T_58636 = _T_58635[5:0]; // @[Modules.scala 143:103:@4423.4]
  assign _T_58637 = $signed(_T_58636); // @[Modules.scala 143:103:@4424.4]
  assign _T_58639 = $signed(-4'sh1) * $signed(io_in_527); // @[Modules.scala 143:74:@4426.4]
  assign _T_58641 = $signed(-4'sh1) * $signed(io_in_528); // @[Modules.scala 144:80:@4427.4]
  assign _T_58642 = $signed(_T_58639) + $signed(_T_58641); // @[Modules.scala 143:103:@4428.4]
  assign _T_58643 = _T_58642[4:0]; // @[Modules.scala 143:103:@4429.4]
  assign _T_58644 = $signed(_T_58643); // @[Modules.scala 143:103:@4430.4]
  assign _T_58646 = $signed(-4'sh1) * $signed(io_in_529); // @[Modules.scala 143:74:@4432.4]
  assign _T_58648 = $signed(-4'sh1) * $signed(io_in_530); // @[Modules.scala 144:80:@4433.4]
  assign _T_58649 = $signed(_T_58646) + $signed(_T_58648); // @[Modules.scala 143:103:@4434.4]
  assign _T_58650 = _T_58649[4:0]; // @[Modules.scala 143:103:@4435.4]
  assign _T_58651 = $signed(_T_58650); // @[Modules.scala 143:103:@4436.4]
  assign _T_58655 = $signed(4'sh1) * $signed(io_in_532); // @[Modules.scala 144:80:@4439.4]
  assign _T_58656 = $signed(_T_55643) + $signed(_T_58655); // @[Modules.scala 143:103:@4440.4]
  assign _T_58657 = _T_58656[5:0]; // @[Modules.scala 143:103:@4441.4]
  assign _T_58658 = $signed(_T_58657); // @[Modules.scala 143:103:@4442.4]
  assign _T_58660 = $signed(-4'sh1) * $signed(io_in_533); // @[Modules.scala 143:74:@4444.4]
  assign _GEN_119 = {{1{_T_58660[4]}},_T_58660}; // @[Modules.scala 143:103:@4446.4]
  assign _T_58663 = $signed(_GEN_119) + $signed(_T_55655); // @[Modules.scala 143:103:@4446.4]
  assign _T_58664 = _T_58663[5:0]; // @[Modules.scala 143:103:@4447.4]
  assign _T_58665 = $signed(_T_58664); // @[Modules.scala 143:103:@4448.4]
  assign _T_58670 = $signed(_T_55657) + $signed(_T_55662); // @[Modules.scala 143:103:@4452.4]
  assign _T_58671 = _T_58670[5:0]; // @[Modules.scala 143:103:@4453.4]
  assign _T_58672 = $signed(_T_58671); // @[Modules.scala 143:103:@4454.4]
  assign _T_58674 = $signed(-4'sh1) * $signed(io_in_537); // @[Modules.scala 143:74:@4456.4]
  assign _T_58676 = $signed(-4'sh1) * $signed(io_in_538); // @[Modules.scala 144:80:@4457.4]
  assign _T_58677 = $signed(_T_58674) + $signed(_T_58676); // @[Modules.scala 143:103:@4458.4]
  assign _T_58678 = _T_58677[4:0]; // @[Modules.scala 143:103:@4459.4]
  assign _T_58679 = $signed(_T_58678); // @[Modules.scala 143:103:@4460.4]
  assign _T_58681 = $signed(-4'sh1) * $signed(io_in_540); // @[Modules.scala 143:74:@4462.4]
  assign _T_58683 = $signed(-4'sh1) * $signed(io_in_541); // @[Modules.scala 144:80:@4463.4]
  assign _T_58684 = $signed(_T_58681) + $signed(_T_58683); // @[Modules.scala 143:103:@4464.4]
  assign _T_58685 = _T_58684[4:0]; // @[Modules.scala 143:103:@4465.4]
  assign _T_58686 = $signed(_T_58685); // @[Modules.scala 143:103:@4466.4]
  assign _T_58688 = $signed(-4'sh1) * $signed(io_in_542); // @[Modules.scala 143:74:@4468.4]
  assign _T_58690 = $signed(-4'sh1) * $signed(io_in_543); // @[Modules.scala 144:80:@4469.4]
  assign _T_58691 = $signed(_T_58688) + $signed(_T_58690); // @[Modules.scala 143:103:@4470.4]
  assign _T_58692 = _T_58691[4:0]; // @[Modules.scala 143:103:@4471.4]
  assign _T_58693 = $signed(_T_58692); // @[Modules.scala 143:103:@4472.4]
  assign _T_58695 = $signed(-4'sh1) * $signed(io_in_544); // @[Modules.scala 143:74:@4474.4]
  assign _T_58697 = $signed(-4'sh1) * $signed(io_in_545); // @[Modules.scala 144:80:@4475.4]
  assign _T_58698 = $signed(_T_58695) + $signed(_T_58697); // @[Modules.scala 143:103:@4476.4]
  assign _T_58699 = _T_58698[4:0]; // @[Modules.scala 143:103:@4477.4]
  assign _T_58700 = $signed(_T_58699); // @[Modules.scala 143:103:@4478.4]
  assign _T_58704 = $signed(-4'sh1) * $signed(io_in_548); // @[Modules.scala 144:80:@4481.4]
  assign _GEN_120 = {{1{_T_58704[4]}},_T_58704}; // @[Modules.scala 143:103:@4482.4]
  assign _T_58705 = $signed(_T_55692) + $signed(_GEN_120); // @[Modules.scala 143:103:@4482.4]
  assign _T_58706 = _T_58705[5:0]; // @[Modules.scala 143:103:@4483.4]
  assign _T_58707 = $signed(_T_58706); // @[Modules.scala 143:103:@4484.4]
  assign _T_58709 = $signed(-4'sh1) * $signed(io_in_549); // @[Modules.scala 143:74:@4486.4]
  assign _T_58711 = $signed(-4'sh1) * $signed(io_in_550); // @[Modules.scala 144:80:@4487.4]
  assign _T_58712 = $signed(_T_58709) + $signed(_T_58711); // @[Modules.scala 143:103:@4488.4]
  assign _T_58713 = _T_58712[4:0]; // @[Modules.scala 143:103:@4489.4]
  assign _T_58714 = $signed(_T_58713); // @[Modules.scala 143:103:@4490.4]
  assign _T_58718 = $signed(-4'sh1) * $signed(io_in_553); // @[Modules.scala 144:80:@4493.4]
  assign _GEN_121 = {{1{_T_58718[4]}},_T_58718}; // @[Modules.scala 143:103:@4494.4]
  assign _T_58719 = $signed(_T_55706) + $signed(_GEN_121); // @[Modules.scala 143:103:@4494.4]
  assign _T_58720 = _T_58719[5:0]; // @[Modules.scala 143:103:@4495.4]
  assign _T_58721 = $signed(_T_58720); // @[Modules.scala 143:103:@4496.4]
  assign _T_58723 = $signed(-4'sh1) * $signed(io_in_554); // @[Modules.scala 143:74:@4498.4]
  assign _T_58725 = $signed(-4'sh1) * $signed(io_in_555); // @[Modules.scala 144:80:@4499.4]
  assign _T_58726 = $signed(_T_58723) + $signed(_T_58725); // @[Modules.scala 143:103:@4500.4]
  assign _T_58727 = _T_58726[4:0]; // @[Modules.scala 143:103:@4501.4]
  assign _T_58728 = $signed(_T_58727); // @[Modules.scala 143:103:@4502.4]
  assign _T_58730 = $signed(-4'sh1) * $signed(io_in_556); // @[Modules.scala 143:74:@4504.4]
  assign _T_58732 = $signed(-4'sh1) * $signed(io_in_557); // @[Modules.scala 144:80:@4505.4]
  assign _T_58733 = $signed(_T_58730) + $signed(_T_58732); // @[Modules.scala 143:103:@4506.4]
  assign _T_58734 = _T_58733[4:0]; // @[Modules.scala 143:103:@4507.4]
  assign _T_58735 = $signed(_T_58734); // @[Modules.scala 143:103:@4508.4]
  assign _T_58737 = $signed(-4'sh1) * $signed(io_in_558); // @[Modules.scala 143:74:@4510.4]
  assign _T_58740 = $signed(_T_58737) + $signed(_T_55725); // @[Modules.scala 143:103:@4512.4]
  assign _T_58741 = _T_58740[4:0]; // @[Modules.scala 143:103:@4513.4]
  assign _T_58742 = $signed(_T_58741); // @[Modules.scala 143:103:@4514.4]
  assign _T_58747 = $signed(_T_55727) + $signed(_T_55732); // @[Modules.scala 143:103:@4518.4]
  assign _T_58748 = _T_58747[5:0]; // @[Modules.scala 143:103:@4519.4]
  assign _T_58749 = $signed(_T_58748); // @[Modules.scala 143:103:@4520.4]
  assign _T_58753 = $signed(-4'sh1) * $signed(io_in_565); // @[Modules.scala 144:80:@4523.4]
  assign _GEN_122 = {{1{_T_58753[4]}},_T_58753}; // @[Modules.scala 143:103:@4524.4]
  assign _T_58754 = $signed(_T_55734) + $signed(_GEN_122); // @[Modules.scala 143:103:@4524.4]
  assign _T_58755 = _T_58754[5:0]; // @[Modules.scala 143:103:@4525.4]
  assign _T_58756 = $signed(_T_58755); // @[Modules.scala 143:103:@4526.4]
  assign _T_58758 = $signed(-4'sh1) * $signed(io_in_566); // @[Modules.scala 143:74:@4528.4]
  assign _T_58760 = $signed(-4'sh1) * $signed(io_in_571); // @[Modules.scala 144:80:@4529.4]
  assign _T_58761 = $signed(_T_58758) + $signed(_T_58760); // @[Modules.scala 143:103:@4530.4]
  assign _T_58762 = _T_58761[4:0]; // @[Modules.scala 143:103:@4531.4]
  assign _T_58763 = $signed(_T_58762); // @[Modules.scala 143:103:@4532.4]
  assign _T_58765 = $signed(-4'sh1) * $signed(io_in_572); // @[Modules.scala 143:74:@4534.4]
  assign _T_58767 = $signed(-4'sh1) * $signed(io_in_573); // @[Modules.scala 144:80:@4535.4]
  assign _T_58768 = $signed(_T_58765) + $signed(_T_58767); // @[Modules.scala 143:103:@4536.4]
  assign _T_58769 = _T_58768[4:0]; // @[Modules.scala 143:103:@4537.4]
  assign _T_58770 = $signed(_T_58769); // @[Modules.scala 143:103:@4538.4]
  assign _T_58774 = $signed(-4'sh1) * $signed(io_in_576); // @[Modules.scala 144:80:@4541.4]
  assign _GEN_123 = {{1{_T_58774[4]}},_T_58774}; // @[Modules.scala 143:103:@4542.4]
  assign _T_58775 = $signed(_T_55762) + $signed(_GEN_123); // @[Modules.scala 143:103:@4542.4]
  assign _T_58776 = _T_58775[5:0]; // @[Modules.scala 143:103:@4543.4]
  assign _T_58777 = $signed(_T_58776); // @[Modules.scala 143:103:@4544.4]
  assign _T_58779 = $signed(-4'sh1) * $signed(io_in_577); // @[Modules.scala 143:74:@4546.4]
  assign _T_58781 = $signed(-4'sh1) * $signed(io_in_578); // @[Modules.scala 144:80:@4547.4]
  assign _T_58782 = $signed(_T_58779) + $signed(_T_58781); // @[Modules.scala 143:103:@4548.4]
  assign _T_58783 = _T_58782[4:0]; // @[Modules.scala 143:103:@4549.4]
  assign _T_58784 = $signed(_T_58783); // @[Modules.scala 143:103:@4550.4]
  assign _T_58786 = $signed(4'sh1) * $signed(io_in_579); // @[Modules.scala 143:74:@4552.4]
  assign _T_58788 = $signed(4'sh1) * $signed(io_in_580); // @[Modules.scala 144:80:@4553.4]
  assign _T_58789 = $signed(_T_58786) + $signed(_T_58788); // @[Modules.scala 143:103:@4554.4]
  assign _T_58790 = _T_58789[5:0]; // @[Modules.scala 143:103:@4555.4]
  assign _T_58791 = $signed(_T_58790); // @[Modules.scala 143:103:@4556.4]
  assign _T_58793 = $signed(-4'sh1) * $signed(io_in_581); // @[Modules.scala 143:74:@4558.4]
  assign _T_58796 = $signed(_T_58793) + $signed(_T_55774); // @[Modules.scala 143:103:@4560.4]
  assign _T_58797 = _T_58796[4:0]; // @[Modules.scala 143:103:@4561.4]
  assign _T_58798 = $signed(_T_58797); // @[Modules.scala 143:103:@4562.4]
  assign _T_58800 = $signed(-4'sh1) * $signed(io_in_583); // @[Modules.scala 143:74:@4564.4]
  assign _T_58802 = $signed(-4'sh1) * $signed(io_in_584); // @[Modules.scala 144:80:@4565.4]
  assign _T_58803 = $signed(_T_58800) + $signed(_T_58802); // @[Modules.scala 143:103:@4566.4]
  assign _T_58804 = _T_58803[4:0]; // @[Modules.scala 143:103:@4567.4]
  assign _T_58805 = $signed(_T_58804); // @[Modules.scala 143:103:@4568.4]
  assign _T_58807 = $signed(-4'sh1) * $signed(io_in_585); // @[Modules.scala 143:74:@4570.4]
  assign _T_58809 = $signed(4'sh1) * $signed(io_in_586); // @[Modules.scala 144:80:@4571.4]
  assign _GEN_124 = {{1{_T_58807[4]}},_T_58807}; // @[Modules.scala 143:103:@4572.4]
  assign _T_58810 = $signed(_GEN_124) + $signed(_T_58809); // @[Modules.scala 143:103:@4572.4]
  assign _T_58811 = _T_58810[5:0]; // @[Modules.scala 143:103:@4573.4]
  assign _T_58812 = $signed(_T_58811); // @[Modules.scala 143:103:@4574.4]
  assign _T_58814 = $signed(-4'sh1) * $signed(io_in_587); // @[Modules.scala 143:74:@4576.4]
  assign _T_58816 = $signed(-4'sh1) * $signed(io_in_588); // @[Modules.scala 144:80:@4577.4]
  assign _T_58817 = $signed(_T_58814) + $signed(_T_58816); // @[Modules.scala 143:103:@4578.4]
  assign _T_58818 = _T_58817[4:0]; // @[Modules.scala 143:103:@4579.4]
  assign _T_58819 = $signed(_T_58818); // @[Modules.scala 143:103:@4580.4]
  assign _T_58837 = $signed(-4'sh1) * $signed(io_in_595); // @[Modules.scala 144:80:@4595.4]
  assign _GEN_125 = {{1{_T_58837[4]}},_T_58837}; // @[Modules.scala 143:103:@4596.4]
  assign _T_58838 = $signed(_T_55809) + $signed(_GEN_125); // @[Modules.scala 143:103:@4596.4]
  assign _T_58839 = _T_58838[5:0]; // @[Modules.scala 143:103:@4597.4]
  assign _T_58840 = $signed(_T_58839); // @[Modules.scala 143:103:@4598.4]
  assign _T_58844 = $signed(-4'sh1) * $signed(io_in_600); // @[Modules.scala 144:80:@4601.4]
  assign _GEN_126 = {{1{_T_58844[4]}},_T_58844}; // @[Modules.scala 143:103:@4602.4]
  assign _T_58845 = $signed(_T_55816) + $signed(_GEN_126); // @[Modules.scala 143:103:@4602.4]
  assign _T_58846 = _T_58845[5:0]; // @[Modules.scala 143:103:@4603.4]
  assign _T_58847 = $signed(_T_58846); // @[Modules.scala 143:103:@4604.4]
  assign _T_58849 = $signed(-4'sh1) * $signed(io_in_601); // @[Modules.scala 143:74:@4606.4]
  assign _T_58851 = $signed(-4'sh1) * $signed(io_in_605); // @[Modules.scala 144:80:@4607.4]
  assign _T_58852 = $signed(_T_58849) + $signed(_T_58851); // @[Modules.scala 143:103:@4608.4]
  assign _T_58853 = _T_58852[4:0]; // @[Modules.scala 143:103:@4609.4]
  assign _T_58854 = $signed(_T_58853); // @[Modules.scala 143:103:@4610.4]
  assign _T_58856 = $signed(-4'sh1) * $signed(io_in_606); // @[Modules.scala 143:74:@4612.4]
  assign _T_58858 = $signed(4'sh1) * $signed(io_in_607); // @[Modules.scala 144:80:@4613.4]
  assign _GEN_127 = {{1{_T_58856[4]}},_T_58856}; // @[Modules.scala 143:103:@4614.4]
  assign _T_58859 = $signed(_GEN_127) + $signed(_T_58858); // @[Modules.scala 143:103:@4614.4]
  assign _T_58860 = _T_58859[5:0]; // @[Modules.scala 143:103:@4615.4]
  assign _T_58861 = $signed(_T_58860); // @[Modules.scala 143:103:@4616.4]
  assign _T_58865 = $signed(-4'sh1) * $signed(io_in_609); // @[Modules.scala 144:80:@4619.4]
  assign _T_58866 = $signed(_T_55837) + $signed(_T_58865); // @[Modules.scala 143:103:@4620.4]
  assign _T_58867 = _T_58866[4:0]; // @[Modules.scala 143:103:@4621.4]
  assign _T_58868 = $signed(_T_58867); // @[Modules.scala 143:103:@4622.4]
  assign _T_58870 = $signed(-4'sh1) * $signed(io_in_610); // @[Modules.scala 143:74:@4624.4]
  assign _T_58872 = $signed(-4'sh1) * $signed(io_in_611); // @[Modules.scala 144:80:@4625.4]
  assign _T_58873 = $signed(_T_58870) + $signed(_T_58872); // @[Modules.scala 143:103:@4626.4]
  assign _T_58874 = _T_58873[4:0]; // @[Modules.scala 143:103:@4627.4]
  assign _T_58875 = $signed(_T_58874); // @[Modules.scala 143:103:@4628.4]
  assign _T_58877 = $signed(-4'sh1) * $signed(io_in_612); // @[Modules.scala 143:74:@4630.4]
  assign _T_58879 = $signed(-4'sh1) * $signed(io_in_613); // @[Modules.scala 144:80:@4631.4]
  assign _T_58880 = $signed(_T_58877) + $signed(_T_58879); // @[Modules.scala 143:103:@4632.4]
  assign _T_58881 = _T_58880[4:0]; // @[Modules.scala 143:103:@4633.4]
  assign _T_58882 = $signed(_T_58881); // @[Modules.scala 143:103:@4634.4]
  assign _T_58886 = $signed(-4'sh1) * $signed(io_in_616); // @[Modules.scala 144:80:@4637.4]
  assign _GEN_128 = {{1{_T_58886[4]}},_T_58886}; // @[Modules.scala 143:103:@4638.4]
  assign _T_58887 = $signed(_T_55858) + $signed(_GEN_128); // @[Modules.scala 143:103:@4638.4]
  assign _T_58888 = _T_58887[5:0]; // @[Modules.scala 143:103:@4639.4]
  assign _T_58889 = $signed(_T_58888); // @[Modules.scala 143:103:@4640.4]
  assign _T_58891 = $signed(-4'sh1) * $signed(io_in_617); // @[Modules.scala 143:74:@4642.4]
  assign _GEN_129 = {{1{_T_58891[4]}},_T_58891}; // @[Modules.scala 143:103:@4644.4]
  assign _T_58894 = $signed(_GEN_129) + $signed(_T_55867); // @[Modules.scala 143:103:@4644.4]
  assign _T_58895 = _T_58894[5:0]; // @[Modules.scala 143:103:@4645.4]
  assign _T_58896 = $signed(_T_58895); // @[Modules.scala 143:103:@4646.4]
  assign _T_58912 = $signed(4'sh1) * $signed(io_in_624); // @[Modules.scala 143:74:@4660.4]
  assign _T_58915 = $signed(_T_58912) + $signed(_T_55888); // @[Modules.scala 143:103:@4662.4]
  assign _T_58916 = _T_58915[5:0]; // @[Modules.scala 143:103:@4663.4]
  assign _T_58917 = $signed(_T_58916); // @[Modules.scala 143:103:@4664.4]
  assign _T_58919 = $signed(4'sh1) * $signed(io_in_626); // @[Modules.scala 143:74:@4666.4]
  assign _GEN_130 = {{1{_T_55895[4]}},_T_55895}; // @[Modules.scala 143:103:@4668.4]
  assign _T_58922 = $signed(_T_58919) + $signed(_GEN_130); // @[Modules.scala 143:103:@4668.4]
  assign _T_58923 = _T_58922[5:0]; // @[Modules.scala 143:103:@4669.4]
  assign _T_58924 = $signed(_T_58923); // @[Modules.scala 143:103:@4670.4]
  assign _T_58929 = $signed(_T_55900) + $signed(_T_55907); // @[Modules.scala 143:103:@4674.4]
  assign _T_58930 = _T_58929[4:0]; // @[Modules.scala 143:103:@4675.4]
  assign _T_58931 = $signed(_T_58930); // @[Modules.scala 143:103:@4676.4]
  assign _T_58933 = $signed(4'sh1) * $signed(io_in_633); // @[Modules.scala 143:74:@4678.4]
  assign _GEN_131 = {{1{_T_55916[4]}},_T_55916}; // @[Modules.scala 143:103:@4680.4]
  assign _T_58936 = $signed(_T_58933) + $signed(_GEN_131); // @[Modules.scala 143:103:@4680.4]
  assign _T_58937 = _T_58936[5:0]; // @[Modules.scala 143:103:@4681.4]
  assign _T_58938 = $signed(_T_58937); // @[Modules.scala 143:103:@4682.4]
  assign _T_58940 = $signed(-4'sh1) * $signed(io_in_636); // @[Modules.scala 143:74:@4684.4]
  assign _T_58942 = $signed(-4'sh1) * $signed(io_in_637); // @[Modules.scala 144:80:@4685.4]
  assign _T_58943 = $signed(_T_58940) + $signed(_T_58942); // @[Modules.scala 143:103:@4686.4]
  assign _T_58944 = _T_58943[4:0]; // @[Modules.scala 143:103:@4687.4]
  assign _T_58945 = $signed(_T_58944); // @[Modules.scala 143:103:@4688.4]
  assign _T_58947 = $signed(-4'sh1) * $signed(io_in_638); // @[Modules.scala 143:74:@4690.4]
  assign _T_58949 = $signed(-4'sh1) * $signed(io_in_639); // @[Modules.scala 144:80:@4691.4]
  assign _T_58950 = $signed(_T_58947) + $signed(_T_58949); // @[Modules.scala 143:103:@4692.4]
  assign _T_58951 = _T_58950[4:0]; // @[Modules.scala 143:103:@4693.4]
  assign _T_58952 = $signed(_T_58951); // @[Modules.scala 143:103:@4694.4]
  assign _T_58954 = $signed(-4'sh1) * $signed(io_in_640); // @[Modules.scala 143:74:@4696.4]
  assign _GEN_132 = {{1{_T_58954[4]}},_T_58954}; // @[Modules.scala 143:103:@4698.4]
  assign _T_58957 = $signed(_GEN_132) + $signed(_T_55942); // @[Modules.scala 143:103:@4698.4]
  assign _T_58958 = _T_58957[5:0]; // @[Modules.scala 143:103:@4699.4]
  assign _T_58959 = $signed(_T_58958); // @[Modules.scala 143:103:@4700.4]
  assign _T_58964 = $signed(_T_55944) + $signed(_T_55949); // @[Modules.scala 143:103:@4704.4]
  assign _T_58965 = _T_58964[5:0]; // @[Modules.scala 143:103:@4705.4]
  assign _T_58966 = $signed(_T_58965); // @[Modules.scala 143:103:@4706.4]
  assign _T_58982 = $signed(4'sh1) * $signed(io_in_652); // @[Modules.scala 143:74:@4720.4]
  assign _T_58984 = $signed(4'sh1) * $signed(io_in_655); // @[Modules.scala 144:80:@4721.4]
  assign _T_58985 = $signed(_T_58982) + $signed(_T_58984); // @[Modules.scala 143:103:@4722.4]
  assign _T_58986 = _T_58985[5:0]; // @[Modules.scala 143:103:@4723.4]
  assign _T_58987 = $signed(_T_58986); // @[Modules.scala 143:103:@4724.4]
  assign _T_58992 = $signed(_T_55986) + $signed(_T_55991); // @[Modules.scala 143:103:@4728.4]
  assign _T_58993 = _T_58992[4:0]; // @[Modules.scala 143:103:@4729.4]
  assign _T_58994 = $signed(_T_58993); // @[Modules.scala 143:103:@4730.4]
  assign _T_58999 = $signed(_T_55993) + $signed(_T_55998); // @[Modules.scala 143:103:@4734.4]
  assign _T_59000 = _T_58999[4:0]; // @[Modules.scala 143:103:@4735.4]
  assign _T_59001 = $signed(_T_59000); // @[Modules.scala 143:103:@4736.4]
  assign _T_59003 = $signed(4'sh1) * $signed(io_in_661); // @[Modules.scala 143:74:@4738.4]
  assign _T_59005 = $signed(4'sh1) * $signed(io_in_663); // @[Modules.scala 144:80:@4739.4]
  assign _T_59006 = $signed(_T_59003) + $signed(_T_59005); // @[Modules.scala 143:103:@4740.4]
  assign _T_59007 = _T_59006[5:0]; // @[Modules.scala 143:103:@4741.4]
  assign _T_59008 = $signed(_T_59007); // @[Modules.scala 143:103:@4742.4]
  assign _T_59017 = $signed(-4'sh1) * $signed(io_in_666); // @[Modules.scala 143:74:@4750.4]
  assign _T_59019 = $signed(-4'sh1) * $signed(io_in_667); // @[Modules.scala 144:80:@4751.4]
  assign _T_59020 = $signed(_T_59017) + $signed(_T_59019); // @[Modules.scala 143:103:@4752.4]
  assign _T_59021 = _T_59020[4:0]; // @[Modules.scala 143:103:@4753.4]
  assign _T_59022 = $signed(_T_59021); // @[Modules.scala 143:103:@4754.4]
  assign _T_59024 = $signed(-4'sh1) * $signed(io_in_668); // @[Modules.scala 143:74:@4756.4]
  assign _GEN_133 = {{1{_T_59024[4]}},_T_59024}; // @[Modules.scala 143:103:@4758.4]
  assign _T_59027 = $signed(_GEN_133) + $signed(_T_56021); // @[Modules.scala 143:103:@4758.4]
  assign _T_59028 = _T_59027[5:0]; // @[Modules.scala 143:103:@4759.4]
  assign _T_59029 = $signed(_T_59028); // @[Modules.scala 143:103:@4760.4]
  assign _T_59033 = $signed(4'sh1) * $signed(io_in_674); // @[Modules.scala 144:80:@4763.4]
  assign _T_59034 = $signed(_T_56026) + $signed(_T_59033); // @[Modules.scala 143:103:@4764.4]
  assign _T_59035 = _T_59034[5:0]; // @[Modules.scala 143:103:@4765.4]
  assign _T_59036 = $signed(_T_59035); // @[Modules.scala 143:103:@4766.4]
  assign _T_59054 = $signed(4'sh1) * $signed(io_in_680); // @[Modules.scala 144:80:@4781.4]
  assign _T_59055 = $signed(_T_56047) + $signed(_T_59054); // @[Modules.scala 143:103:@4782.4]
  assign _T_59056 = _T_59055[5:0]; // @[Modules.scala 143:103:@4783.4]
  assign _T_59057 = $signed(_T_59056); // @[Modules.scala 143:103:@4784.4]
  assign _T_59059 = $signed(4'sh1) * $signed(io_in_681); // @[Modules.scala 143:74:@4786.4]
  assign _T_59061 = $signed(4'sh1) * $signed(io_in_683); // @[Modules.scala 144:80:@4787.4]
  assign _T_59062 = $signed(_T_59059) + $signed(_T_59061); // @[Modules.scala 143:103:@4788.4]
  assign _T_59063 = _T_59062[5:0]; // @[Modules.scala 143:103:@4789.4]
  assign _T_59064 = $signed(_T_59063); // @[Modules.scala 143:103:@4790.4]
  assign _T_59066 = $signed(-4'sh1) * $signed(io_in_684); // @[Modules.scala 143:74:@4792.4]
  assign _T_59069 = $signed(_T_59066) + $signed(_T_56061); // @[Modules.scala 143:103:@4794.4]
  assign _T_59070 = _T_59069[4:0]; // @[Modules.scala 143:103:@4795.4]
  assign _T_59071 = $signed(_T_59070); // @[Modules.scala 143:103:@4796.4]
  assign _T_59075 = $signed(4'sh1) * $signed(io_in_687); // @[Modules.scala 144:80:@4799.4]
  assign _GEN_134 = {{1{_T_56063[4]}},_T_56063}; // @[Modules.scala 143:103:@4800.4]
  assign _T_59076 = $signed(_GEN_134) + $signed(_T_59075); // @[Modules.scala 143:103:@4800.4]
  assign _T_59077 = _T_59076[5:0]; // @[Modules.scala 143:103:@4801.4]
  assign _T_59078 = $signed(_T_59077); // @[Modules.scala 143:103:@4802.4]
  assign _T_59080 = $signed(4'sh1) * $signed(io_in_688); // @[Modules.scala 143:74:@4804.4]
  assign _T_59082 = $signed(4'sh1) * $signed(io_in_689); // @[Modules.scala 144:80:@4805.4]
  assign _T_59083 = $signed(_T_59080) + $signed(_T_59082); // @[Modules.scala 143:103:@4806.4]
  assign _T_59084 = _T_59083[5:0]; // @[Modules.scala 143:103:@4807.4]
  assign _T_59085 = $signed(_T_59084); // @[Modules.scala 143:103:@4808.4]
  assign _T_59087 = $signed(4'sh1) * $signed(io_in_690); // @[Modules.scala 143:74:@4810.4]
  assign _T_59089 = $signed(4'sh1) * $signed(io_in_691); // @[Modules.scala 144:80:@4811.4]
  assign _T_59090 = $signed(_T_59087) + $signed(_T_59089); // @[Modules.scala 143:103:@4812.4]
  assign _T_59091 = _T_59090[5:0]; // @[Modules.scala 143:103:@4813.4]
  assign _T_59092 = $signed(_T_59091); // @[Modules.scala 143:103:@4814.4]
  assign _T_59094 = $signed(4'sh1) * $signed(io_in_692); // @[Modules.scala 143:74:@4816.4]
  assign _GEN_135 = {{1{_T_56089[4]}},_T_56089}; // @[Modules.scala 143:103:@4818.4]
  assign _T_59097 = $signed(_T_59094) + $signed(_GEN_135); // @[Modules.scala 143:103:@4818.4]
  assign _T_59098 = _T_59097[5:0]; // @[Modules.scala 143:103:@4819.4]
  assign _T_59099 = $signed(_T_59098); // @[Modules.scala 143:103:@4820.4]
  assign _T_59104 = $signed(_T_56091) + $signed(_T_56096); // @[Modules.scala 143:103:@4824.4]
  assign _T_59105 = _T_59104[4:0]; // @[Modules.scala 143:103:@4825.4]
  assign _T_59106 = $signed(_T_59105); // @[Modules.scala 143:103:@4826.4]
  assign _T_59108 = $signed(-4'sh1) * $signed(io_in_696); // @[Modules.scala 143:74:@4828.4]
  assign _GEN_136 = {{1{_T_59108[4]}},_T_59108}; // @[Modules.scala 143:103:@4830.4]
  assign _T_59111 = $signed(_GEN_136) + $signed(_T_56105); // @[Modules.scala 143:103:@4830.4]
  assign _T_59112 = _T_59111[5:0]; // @[Modules.scala 143:103:@4831.4]
  assign _T_59113 = $signed(_T_59112); // @[Modules.scala 143:103:@4832.4]
  assign _T_59115 = $signed(-4'sh1) * $signed(io_in_699); // @[Modules.scala 143:74:@4834.4]
  assign _GEN_137 = {{1{_T_59115[4]}},_T_59115}; // @[Modules.scala 143:103:@4836.4]
  assign _T_59118 = $signed(_GEN_137) + $signed(_T_56110); // @[Modules.scala 143:103:@4836.4]
  assign _T_59119 = _T_59118[5:0]; // @[Modules.scala 143:103:@4837.4]
  assign _T_59120 = $signed(_T_59119); // @[Modules.scala 143:103:@4838.4]
  assign _T_59122 = $signed(-4'sh1) * $signed(io_in_703); // @[Modules.scala 143:74:@4840.4]
  assign _T_59124 = $signed(4'sh1) * $signed(io_in_705); // @[Modules.scala 144:80:@4841.4]
  assign _GEN_138 = {{1{_T_59122[4]}},_T_59122}; // @[Modules.scala 143:103:@4842.4]
  assign _T_59125 = $signed(_GEN_138) + $signed(_T_59124); // @[Modules.scala 143:103:@4842.4]
  assign _T_59126 = _T_59125[5:0]; // @[Modules.scala 143:103:@4843.4]
  assign _T_59127 = $signed(_T_59126); // @[Modules.scala 143:103:@4844.4]
  assign _T_59129 = $signed(4'sh1) * $signed(io_in_706); // @[Modules.scala 143:74:@4846.4]
  assign _T_59131 = $signed(4'sh1) * $signed(io_in_707); // @[Modules.scala 144:80:@4847.4]
  assign _T_59132 = $signed(_T_59129) + $signed(_T_59131); // @[Modules.scala 143:103:@4848.4]
  assign _T_59133 = _T_59132[5:0]; // @[Modules.scala 143:103:@4849.4]
  assign _T_59134 = $signed(_T_59133); // @[Modules.scala 143:103:@4850.4]
  assign _T_59139 = $signed(_T_56126) + $signed(_T_56131); // @[Modules.scala 143:103:@4854.4]
  assign _T_59140 = _T_59139[5:0]; // @[Modules.scala 143:103:@4855.4]
  assign _T_59141 = $signed(_T_59140); // @[Modules.scala 143:103:@4856.4]
  assign _T_59146 = $signed(_T_56133) + $signed(_T_56138); // @[Modules.scala 143:103:@4860.4]
  assign _T_59147 = _T_59146[5:0]; // @[Modules.scala 143:103:@4861.4]
  assign _T_59148 = $signed(_T_59147); // @[Modules.scala 143:103:@4862.4]
  assign _T_59152 = $signed(4'sh1) * $signed(io_in_713); // @[Modules.scala 144:80:@4865.4]
  assign _T_59153 = $signed(_T_56140) + $signed(_T_59152); // @[Modules.scala 143:103:@4866.4]
  assign _T_59154 = _T_59153[5:0]; // @[Modules.scala 143:103:@4867.4]
  assign _T_59155 = $signed(_T_59154); // @[Modules.scala 143:103:@4868.4]
  assign _T_59157 = $signed(4'sh1) * $signed(io_in_714); // @[Modules.scala 143:74:@4870.4]
  assign _T_59159 = $signed(4'sh1) * $signed(io_in_715); // @[Modules.scala 144:80:@4871.4]
  assign _T_59160 = $signed(_T_59157) + $signed(_T_59159); // @[Modules.scala 143:103:@4872.4]
  assign _T_59161 = _T_59160[5:0]; // @[Modules.scala 143:103:@4873.4]
  assign _T_59162 = $signed(_T_59161); // @[Modules.scala 143:103:@4874.4]
  assign _T_59164 = $signed(4'sh1) * $signed(io_in_716); // @[Modules.scala 143:74:@4876.4]
  assign _T_59166 = $signed(4'sh1) * $signed(io_in_717); // @[Modules.scala 144:80:@4877.4]
  assign _T_59167 = $signed(_T_59164) + $signed(_T_59166); // @[Modules.scala 143:103:@4878.4]
  assign _T_59168 = _T_59167[5:0]; // @[Modules.scala 143:103:@4879.4]
  assign _T_59169 = $signed(_T_59168); // @[Modules.scala 143:103:@4880.4]
  assign _T_59171 = $signed(4'sh1) * $signed(io_in_718); // @[Modules.scala 143:74:@4882.4]
  assign _T_59173 = $signed(4'sh1) * $signed(io_in_719); // @[Modules.scala 144:80:@4883.4]
  assign _T_59174 = $signed(_T_59171) + $signed(_T_59173); // @[Modules.scala 143:103:@4884.4]
  assign _T_59175 = _T_59174[5:0]; // @[Modules.scala 143:103:@4885.4]
  assign _T_59176 = $signed(_T_59175); // @[Modules.scala 143:103:@4886.4]
  assign _T_59178 = $signed(4'sh1) * $signed(io_in_720); // @[Modules.scala 143:74:@4888.4]
  assign _T_59180 = $signed(4'sh1) * $signed(io_in_721); // @[Modules.scala 144:80:@4889.4]
  assign _T_59181 = $signed(_T_59178) + $signed(_T_59180); // @[Modules.scala 143:103:@4890.4]
  assign _T_59182 = _T_59181[5:0]; // @[Modules.scala 143:103:@4891.4]
  assign _T_59183 = $signed(_T_59182); // @[Modules.scala 143:103:@4892.4]
  assign _T_59185 = $signed(4'sh1) * $signed(io_in_725); // @[Modules.scala 143:74:@4894.4]
  assign _GEN_139 = {{1{_T_56189[4]}},_T_56189}; // @[Modules.scala 143:103:@4896.4]
  assign _T_59188 = $signed(_T_59185) + $signed(_GEN_139); // @[Modules.scala 143:103:@4896.4]
  assign _T_59189 = _T_59188[5:0]; // @[Modules.scala 143:103:@4897.4]
  assign _T_59190 = $signed(_T_59189); // @[Modules.scala 143:103:@4898.4]
  assign _T_59194 = $signed(-4'sh1) * $signed(io_in_732); // @[Modules.scala 144:80:@4901.4]
  assign _T_59195 = $signed(_T_56194) + $signed(_T_59194); // @[Modules.scala 143:103:@4902.4]
  assign _T_59196 = _T_59195[4:0]; // @[Modules.scala 143:103:@4903.4]
  assign _T_59197 = $signed(_T_59196); // @[Modules.scala 143:103:@4904.4]
  assign _T_59199 = $signed(-4'sh1) * $signed(io_in_733); // @[Modules.scala 143:74:@4906.4]
  assign _T_59201 = $signed(4'sh1) * $signed(io_in_734); // @[Modules.scala 144:80:@4907.4]
  assign _GEN_140 = {{1{_T_59199[4]}},_T_59199}; // @[Modules.scala 143:103:@4908.4]
  assign _T_59202 = $signed(_GEN_140) + $signed(_T_59201); // @[Modules.scala 143:103:@4908.4]
  assign _T_59203 = _T_59202[5:0]; // @[Modules.scala 143:103:@4909.4]
  assign _T_59204 = $signed(_T_59203); // @[Modules.scala 143:103:@4910.4]
  assign _T_59206 = $signed(4'sh1) * $signed(io_in_735); // @[Modules.scala 143:74:@4912.4]
  assign _T_59209 = $signed(_T_59206) + $signed(_T_56196); // @[Modules.scala 143:103:@4914.4]
  assign _T_59210 = _T_59209[5:0]; // @[Modules.scala 143:103:@4915.4]
  assign _T_59211 = $signed(_T_59210); // @[Modules.scala 143:103:@4916.4]
  assign _T_59227 = $signed(4'sh1) * $signed(io_in_741); // @[Modules.scala 143:74:@4930.4]
  assign _T_59229 = $signed(4'sh1) * $signed(io_in_742); // @[Modules.scala 144:80:@4931.4]
  assign _T_59230 = $signed(_T_59227) + $signed(_T_59229); // @[Modules.scala 143:103:@4932.4]
  assign _T_59231 = _T_59230[5:0]; // @[Modules.scala 143:103:@4933.4]
  assign _T_59232 = $signed(_T_59231); // @[Modules.scala 143:103:@4934.4]
  assign _T_59234 = $signed(4'sh1) * $signed(io_in_743); // @[Modules.scala 143:74:@4936.4]
  assign _T_59237 = $signed(_T_59234) + $signed(_T_56217); // @[Modules.scala 143:103:@4938.4]
  assign _T_59238 = _T_59237[5:0]; // @[Modules.scala 143:103:@4939.4]
  assign _T_59239 = $signed(_T_59238); // @[Modules.scala 143:103:@4940.4]
  assign _T_59243 = $signed(4'sh1) * $signed(io_in_746); // @[Modules.scala 144:80:@4943.4]
  assign _T_59244 = $signed(_T_56222) + $signed(_T_59243); // @[Modules.scala 143:103:@4944.4]
  assign _T_59245 = _T_59244[5:0]; // @[Modules.scala 143:103:@4945.4]
  assign _T_59246 = $signed(_T_59245); // @[Modules.scala 143:103:@4946.4]
  assign _T_59248 = $signed(4'sh1) * $signed(io_in_747); // @[Modules.scala 143:74:@4948.4]
  assign _T_59250 = $signed(4'sh1) * $signed(io_in_748); // @[Modules.scala 144:80:@4949.4]
  assign _T_59251 = $signed(_T_59248) + $signed(_T_59250); // @[Modules.scala 143:103:@4950.4]
  assign _T_59252 = _T_59251[5:0]; // @[Modules.scala 143:103:@4951.4]
  assign _T_59253 = $signed(_T_59252); // @[Modules.scala 143:103:@4952.4]
  assign _T_59255 = $signed(4'sh1) * $signed(io_in_749); // @[Modules.scala 143:74:@4954.4]
  assign _T_59258 = $signed(_T_59255) + $signed(_GEN_75); // @[Modules.scala 143:103:@4956.4]
  assign _T_59259 = _T_59258[5:0]; // @[Modules.scala 143:103:@4957.4]
  assign _T_59260 = $signed(_T_59259); // @[Modules.scala 143:103:@4958.4]
  assign _T_59264 = $signed(4'sh1) * $signed(io_in_753); // @[Modules.scala 144:80:@4961.4]
  assign _T_59265 = $signed(_T_56245) + $signed(_T_59264); // @[Modules.scala 143:103:@4962.4]
  assign _T_59266 = _T_59265[5:0]; // @[Modules.scala 143:103:@4963.4]
  assign _T_59267 = $signed(_T_59266); // @[Modules.scala 143:103:@4964.4]
  assign _T_59269 = $signed(-4'sh1) * $signed(io_in_760); // @[Modules.scala 143:74:@4966.4]
  assign _GEN_142 = {{1{_T_59269[4]}},_T_59269}; // @[Modules.scala 143:103:@4968.4]
  assign _T_59272 = $signed(_GEN_142) + $signed(_T_56252); // @[Modules.scala 143:103:@4968.4]
  assign _T_59273 = _T_59272[5:0]; // @[Modules.scala 143:103:@4969.4]
  assign _T_59274 = $signed(_T_59273); // @[Modules.scala 143:103:@4970.4]
  assign _T_59276 = $signed(4'sh1) * $signed(io_in_762); // @[Modules.scala 143:74:@4972.4]
  assign _T_59278 = $signed(4'sh1) * $signed(io_in_764); // @[Modules.scala 144:80:@4973.4]
  assign _T_59279 = $signed(_T_59276) + $signed(_T_59278); // @[Modules.scala 143:103:@4974.4]
  assign _T_59280 = _T_59279[5:0]; // @[Modules.scala 143:103:@4975.4]
  assign _T_59281 = $signed(_T_59280); // @[Modules.scala 143:103:@4976.4]
  assign _T_59290 = $signed(-4'sh1) * $signed(io_in_767); // @[Modules.scala 143:74:@4984.4]
  assign _T_59292 = $signed(-4'sh1) * $signed(io_in_768); // @[Modules.scala 144:80:@4985.4]
  assign _T_59293 = $signed(_T_59290) + $signed(_T_59292); // @[Modules.scala 143:103:@4986.4]
  assign _T_59294 = _T_59293[4:0]; // @[Modules.scala 143:103:@4987.4]
  assign _T_59295 = $signed(_T_59294); // @[Modules.scala 143:103:@4988.4]
  assign _T_59300 = $signed(_T_56273) + $signed(_T_56278); // @[Modules.scala 143:103:@4992.4]
  assign _T_59301 = _T_59300[5:0]; // @[Modules.scala 143:103:@4993.4]
  assign _T_59302 = $signed(_T_59301); // @[Modules.scala 143:103:@4994.4]
  assign _T_59307 = $signed(_T_56280) + $signed(_T_56285); // @[Modules.scala 143:103:@4998.4]
  assign _T_59308 = _T_59307[5:0]; // @[Modules.scala 143:103:@4999.4]
  assign _T_59309 = $signed(_T_59308); // @[Modules.scala 143:103:@5000.4]
  assign _T_59313 = $signed(4'sh1) * $signed(io_in_774); // @[Modules.scala 144:80:@5003.4]
  assign _T_59314 = $signed(_T_56287) + $signed(_T_59313); // @[Modules.scala 143:103:@5004.4]
  assign _T_59315 = _T_59314[5:0]; // @[Modules.scala 143:103:@5005.4]
  assign _T_59316 = $signed(_T_59315); // @[Modules.scala 143:103:@5006.4]
  assign _T_59318 = $signed(4'sh1) * $signed(io_in_775); // @[Modules.scala 143:74:@5008.4]
  assign _T_59320 = $signed(4'sh1) * $signed(io_in_776); // @[Modules.scala 144:80:@5009.4]
  assign _T_59321 = $signed(_T_59318) + $signed(_T_59320); // @[Modules.scala 143:103:@5010.4]
  assign _T_59322 = _T_59321[5:0]; // @[Modules.scala 143:103:@5011.4]
  assign _T_59323 = $signed(_T_59322); // @[Modules.scala 143:103:@5012.4]
  assign _T_59327 = $signed(-4'sh1) * $signed(io_in_778); // @[Modules.scala 144:80:@5015.4]
  assign _GEN_143 = {{1{_T_59327[4]}},_T_59327}; // @[Modules.scala 143:103:@5016.4]
  assign _T_59328 = $signed(_T_56299) + $signed(_GEN_143); // @[Modules.scala 143:103:@5016.4]
  assign _T_59329 = _T_59328[5:0]; // @[Modules.scala 143:103:@5017.4]
  assign _T_59330 = $signed(_T_59329); // @[Modules.scala 143:103:@5018.4]
  assign _T_59332 = $signed(-4'sh1) * $signed(io_in_779); // @[Modules.scala 143:74:@5020.4]
  assign _T_59334 = $signed(-4'sh1) * $signed(io_in_780); // @[Modules.scala 144:80:@5021.4]
  assign _T_59335 = $signed(_T_59332) + $signed(_T_59334); // @[Modules.scala 143:103:@5022.4]
  assign _T_59336 = _T_59335[4:0]; // @[Modules.scala 143:103:@5023.4]
  assign _T_59337 = $signed(_T_59336); // @[Modules.scala 143:103:@5024.4]
  assign buffer_1_2 = {{8{_T_57230[5]}},_T_57230}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_3 = {{8{_T_57237[5]}},_T_57237}; // @[Modules.scala 112:22:@8.4]
  assign _T_59341 = $signed(buffer_1_2) + $signed(buffer_1_3); // @[Modules.scala 160:64:@5030.4]
  assign _T_59342 = _T_59341[13:0]; // @[Modules.scala 160:64:@5031.4]
  assign buffer_1_305 = $signed(_T_59342); // @[Modules.scala 160:64:@5032.4]
  assign buffer_1_4 = {{9{_T_57244[4]}},_T_57244}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_5 = {{8{_T_57251[5]}},_T_57251}; // @[Modules.scala 112:22:@8.4]
  assign _T_59344 = $signed(buffer_1_4) + $signed(buffer_1_5); // @[Modules.scala 160:64:@5034.4]
  assign _T_59345 = _T_59344[13:0]; // @[Modules.scala 160:64:@5035.4]
  assign buffer_1_306 = $signed(_T_59345); // @[Modules.scala 160:64:@5036.4]
  assign buffer_1_6 = {{9{_T_57258[4]}},_T_57258}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_7 = {{9{_T_57265[4]}},_T_57265}; // @[Modules.scala 112:22:@8.4]
  assign _T_59347 = $signed(buffer_1_6) + $signed(buffer_1_7); // @[Modules.scala 160:64:@5038.4]
  assign _T_59348 = _T_59347[13:0]; // @[Modules.scala 160:64:@5039.4]
  assign buffer_1_307 = $signed(_T_59348); // @[Modules.scala 160:64:@5040.4]
  assign buffer_1_8 = {{8{_T_57272[5]}},_T_57272}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_9 = {{9{_T_57279[4]}},_T_57279}; // @[Modules.scala 112:22:@8.4]
  assign _T_59350 = $signed(buffer_1_8) + $signed(buffer_1_9); // @[Modules.scala 160:64:@5042.4]
  assign _T_59351 = _T_59350[13:0]; // @[Modules.scala 160:64:@5043.4]
  assign buffer_1_308 = $signed(_T_59351); // @[Modules.scala 160:64:@5044.4]
  assign buffer_1_10 = {{8{_T_57286[5]}},_T_57286}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_11 = {{8{_T_57293[5]}},_T_57293}; // @[Modules.scala 112:22:@8.4]
  assign _T_59353 = $signed(buffer_1_10) + $signed(buffer_1_11); // @[Modules.scala 160:64:@5046.4]
  assign _T_59354 = _T_59353[13:0]; // @[Modules.scala 160:64:@5047.4]
  assign buffer_1_309 = $signed(_T_59354); // @[Modules.scala 160:64:@5048.4]
  assign buffer_1_12 = {{8{_T_57300[5]}},_T_57300}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_13 = {{9{_T_57307[4]}},_T_57307}; // @[Modules.scala 112:22:@8.4]
  assign _T_59356 = $signed(buffer_1_12) + $signed(buffer_1_13); // @[Modules.scala 160:64:@5050.4]
  assign _T_59357 = _T_59356[13:0]; // @[Modules.scala 160:64:@5051.4]
  assign buffer_1_310 = $signed(_T_59357); // @[Modules.scala 160:64:@5052.4]
  assign buffer_1_14 = {{9{_T_57314[4]}},_T_57314}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_15 = {{9{_T_57321[4]}},_T_57321}; // @[Modules.scala 112:22:@8.4]
  assign _T_59359 = $signed(buffer_1_14) + $signed(buffer_1_15); // @[Modules.scala 160:64:@5054.4]
  assign _T_59360 = _T_59359[13:0]; // @[Modules.scala 160:64:@5055.4]
  assign buffer_1_311 = $signed(_T_59360); // @[Modules.scala 160:64:@5056.4]
  assign buffer_1_16 = {{9{_T_57328[4]}},_T_57328}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_17 = {{9{_T_57335[4]}},_T_57335}; // @[Modules.scala 112:22:@8.4]
  assign _T_59362 = $signed(buffer_1_16) + $signed(buffer_1_17); // @[Modules.scala 160:64:@5058.4]
  assign _T_59363 = _T_59362[13:0]; // @[Modules.scala 160:64:@5059.4]
  assign buffer_1_312 = $signed(_T_59363); // @[Modules.scala 160:64:@5060.4]
  assign buffer_1_18 = {{9{_T_57342[4]}},_T_57342}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_19 = {{8{_T_57349[5]}},_T_57349}; // @[Modules.scala 112:22:@8.4]
  assign _T_59365 = $signed(buffer_1_18) + $signed(buffer_1_19); // @[Modules.scala 160:64:@5062.4]
  assign _T_59366 = _T_59365[13:0]; // @[Modules.scala 160:64:@5063.4]
  assign buffer_1_313 = $signed(_T_59366); // @[Modules.scala 160:64:@5064.4]
  assign buffer_1_20 = {{8{_T_57356[5]}},_T_57356}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_21 = {{8{_T_57363[5]}},_T_57363}; // @[Modules.scala 112:22:@8.4]
  assign _T_59368 = $signed(buffer_1_20) + $signed(buffer_1_21); // @[Modules.scala 160:64:@5066.4]
  assign _T_59369 = _T_59368[13:0]; // @[Modules.scala 160:64:@5067.4]
  assign buffer_1_314 = $signed(_T_59369); // @[Modules.scala 160:64:@5068.4]
  assign buffer_1_22 = {{8{_T_57370[5]}},_T_57370}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_23 = {{8{_T_57377[5]}},_T_57377}; // @[Modules.scala 112:22:@8.4]
  assign _T_59371 = $signed(buffer_1_22) + $signed(buffer_1_23); // @[Modules.scala 160:64:@5070.4]
  assign _T_59372 = _T_59371[13:0]; // @[Modules.scala 160:64:@5071.4]
  assign buffer_1_315 = $signed(_T_59372); // @[Modules.scala 160:64:@5072.4]
  assign buffer_1_24 = {{9{_T_57384[4]}},_T_57384}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_25 = {{9{_T_57391[4]}},_T_57391}; // @[Modules.scala 112:22:@8.4]
  assign _T_59374 = $signed(buffer_1_24) + $signed(buffer_1_25); // @[Modules.scala 160:64:@5074.4]
  assign _T_59375 = _T_59374[13:0]; // @[Modules.scala 160:64:@5075.4]
  assign buffer_1_316 = $signed(_T_59375); // @[Modules.scala 160:64:@5076.4]
  assign buffer_1_26 = {{9{_T_57398[4]}},_T_57398}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_27 = {{9{_T_57405[4]}},_T_57405}; // @[Modules.scala 112:22:@8.4]
  assign _T_59377 = $signed(buffer_1_26) + $signed(buffer_1_27); // @[Modules.scala 160:64:@5078.4]
  assign _T_59378 = _T_59377[13:0]; // @[Modules.scala 160:64:@5079.4]
  assign buffer_1_317 = $signed(_T_59378); // @[Modules.scala 160:64:@5080.4]
  assign buffer_1_28 = {{8{_T_57412[5]}},_T_57412}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_29 = {{9{_T_57419[4]}},_T_57419}; // @[Modules.scala 112:22:@8.4]
  assign _T_59380 = $signed(buffer_1_28) + $signed(buffer_1_29); // @[Modules.scala 160:64:@5082.4]
  assign _T_59381 = _T_59380[13:0]; // @[Modules.scala 160:64:@5083.4]
  assign buffer_1_318 = $signed(_T_59381); // @[Modules.scala 160:64:@5084.4]
  assign buffer_1_30 = {{9{_T_57426[4]}},_T_57426}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_31 = {{9{_T_57433[4]}},_T_57433}; // @[Modules.scala 112:22:@8.4]
  assign _T_59383 = $signed(buffer_1_30) + $signed(buffer_1_31); // @[Modules.scala 160:64:@5086.4]
  assign _T_59384 = _T_59383[13:0]; // @[Modules.scala 160:64:@5087.4]
  assign buffer_1_319 = $signed(_T_59384); // @[Modules.scala 160:64:@5088.4]
  assign buffer_1_32 = {{8{_T_57440[5]}},_T_57440}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_33 = {{8{_T_57447[5]}},_T_57447}; // @[Modules.scala 112:22:@8.4]
  assign _T_59386 = $signed(buffer_1_32) + $signed(buffer_1_33); // @[Modules.scala 160:64:@5090.4]
  assign _T_59387 = _T_59386[13:0]; // @[Modules.scala 160:64:@5091.4]
  assign buffer_1_320 = $signed(_T_59387); // @[Modules.scala 160:64:@5092.4]
  assign buffer_1_34 = {{8{_T_57454[5]}},_T_57454}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_35 = {{8{_T_57461[5]}},_T_57461}; // @[Modules.scala 112:22:@8.4]
  assign _T_59389 = $signed(buffer_1_34) + $signed(buffer_1_35); // @[Modules.scala 160:64:@5094.4]
  assign _T_59390 = _T_59389[13:0]; // @[Modules.scala 160:64:@5095.4]
  assign buffer_1_321 = $signed(_T_59390); // @[Modules.scala 160:64:@5096.4]
  assign buffer_1_36 = {{8{_T_57468[5]}},_T_57468}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_37 = {{8{_T_57475[5]}},_T_57475}; // @[Modules.scala 112:22:@8.4]
  assign _T_59392 = $signed(buffer_1_36) + $signed(buffer_1_37); // @[Modules.scala 160:64:@5098.4]
  assign _T_59393 = _T_59392[13:0]; // @[Modules.scala 160:64:@5099.4]
  assign buffer_1_322 = $signed(_T_59393); // @[Modules.scala 160:64:@5100.4]
  assign buffer_1_38 = {{8{_T_57482[5]}},_T_57482}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_39 = {{8{_T_57489[5]}},_T_57489}; // @[Modules.scala 112:22:@8.4]
  assign _T_59395 = $signed(buffer_1_38) + $signed(buffer_1_39); // @[Modules.scala 160:64:@5102.4]
  assign _T_59396 = _T_59395[13:0]; // @[Modules.scala 160:64:@5103.4]
  assign buffer_1_323 = $signed(_T_59396); // @[Modules.scala 160:64:@5104.4]
  assign buffer_1_41 = {{8{_T_57503[5]}},_T_57503}; // @[Modules.scala 112:22:@8.4]
  assign _T_59398 = $signed(buffer_0_42) + $signed(buffer_1_41); // @[Modules.scala 160:64:@5106.4]
  assign _T_59399 = _T_59398[13:0]; // @[Modules.scala 160:64:@5107.4]
  assign buffer_1_324 = $signed(_T_59399); // @[Modules.scala 160:64:@5108.4]
  assign buffer_1_42 = {{8{_T_57510[5]}},_T_57510}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_43 = {{8{_T_57517[5]}},_T_57517}; // @[Modules.scala 112:22:@8.4]
  assign _T_59401 = $signed(buffer_1_42) + $signed(buffer_1_43); // @[Modules.scala 160:64:@5110.4]
  assign _T_59402 = _T_59401[13:0]; // @[Modules.scala 160:64:@5111.4]
  assign buffer_1_325 = $signed(_T_59402); // @[Modules.scala 160:64:@5112.4]
  assign buffer_1_44 = {{8{_T_57524[5]}},_T_57524}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_45 = {{8{_T_57531[5]}},_T_57531}; // @[Modules.scala 112:22:@8.4]
  assign _T_59404 = $signed(buffer_1_44) + $signed(buffer_1_45); // @[Modules.scala 160:64:@5114.4]
  assign _T_59405 = _T_59404[13:0]; // @[Modules.scala 160:64:@5115.4]
  assign buffer_1_326 = $signed(_T_59405); // @[Modules.scala 160:64:@5116.4]
  assign buffer_1_46 = {{8{_T_57538[5]}},_T_57538}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_47 = {{8{_T_57545[5]}},_T_57545}; // @[Modules.scala 112:22:@8.4]
  assign _T_59407 = $signed(buffer_1_46) + $signed(buffer_1_47); // @[Modules.scala 160:64:@5118.4]
  assign _T_59408 = _T_59407[13:0]; // @[Modules.scala 160:64:@5119.4]
  assign buffer_1_327 = $signed(_T_59408); // @[Modules.scala 160:64:@5120.4]
  assign buffer_1_49 = {{8{_T_57559[5]}},_T_57559}; // @[Modules.scala 112:22:@8.4]
  assign _T_59410 = $signed(buffer_0_48) + $signed(buffer_1_49); // @[Modules.scala 160:64:@5122.4]
  assign _T_59411 = _T_59410[13:0]; // @[Modules.scala 160:64:@5123.4]
  assign buffer_1_328 = $signed(_T_59411); // @[Modules.scala 160:64:@5124.4]
  assign buffer_1_50 = {{9{_T_57566[4]}},_T_57566}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_51 = {{9{_T_57573[4]}},_T_57573}; // @[Modules.scala 112:22:@8.4]
  assign _T_59413 = $signed(buffer_1_50) + $signed(buffer_1_51); // @[Modules.scala 160:64:@5126.4]
  assign _T_59414 = _T_59413[13:0]; // @[Modules.scala 160:64:@5127.4]
  assign buffer_1_329 = $signed(_T_59414); // @[Modules.scala 160:64:@5128.4]
  assign buffer_1_52 = {{8{_T_57580[5]}},_T_57580}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_53 = {{9{_T_57587[4]}},_T_57587}; // @[Modules.scala 112:22:@8.4]
  assign _T_59416 = $signed(buffer_1_52) + $signed(buffer_1_53); // @[Modules.scala 160:64:@5130.4]
  assign _T_59417 = _T_59416[13:0]; // @[Modules.scala 160:64:@5131.4]
  assign buffer_1_330 = $signed(_T_59417); // @[Modules.scala 160:64:@5132.4]
  assign buffer_1_54 = {{9{_T_57594[4]}},_T_57594}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_55 = {{8{_T_57601[5]}},_T_57601}; // @[Modules.scala 112:22:@8.4]
  assign _T_59419 = $signed(buffer_1_54) + $signed(buffer_1_55); // @[Modules.scala 160:64:@5134.4]
  assign _T_59420 = _T_59419[13:0]; // @[Modules.scala 160:64:@5135.4]
  assign buffer_1_331 = $signed(_T_59420); // @[Modules.scala 160:64:@5136.4]
  assign _T_59422 = $signed(buffer_0_55) + $signed(buffer_0_56); // @[Modules.scala 160:64:@5138.4]
  assign _T_59423 = _T_59422[13:0]; // @[Modules.scala 160:64:@5139.4]
  assign buffer_1_332 = $signed(_T_59423); // @[Modules.scala 160:64:@5140.4]
  assign buffer_1_58 = {{8{_T_57622[5]}},_T_57622}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_59 = {{8{_T_57629[5]}},_T_57629}; // @[Modules.scala 112:22:@8.4]
  assign _T_59425 = $signed(buffer_1_58) + $signed(buffer_1_59); // @[Modules.scala 160:64:@5142.4]
  assign _T_59426 = _T_59425[13:0]; // @[Modules.scala 160:64:@5143.4]
  assign buffer_1_333 = $signed(_T_59426); // @[Modules.scala 160:64:@5144.4]
  assign buffer_1_60 = {{8{_T_57636[5]}},_T_57636}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_61 = {{8{_T_57643[5]}},_T_57643}; // @[Modules.scala 112:22:@8.4]
  assign _T_59428 = $signed(buffer_1_60) + $signed(buffer_1_61); // @[Modules.scala 160:64:@5146.4]
  assign _T_59429 = _T_59428[13:0]; // @[Modules.scala 160:64:@5147.4]
  assign buffer_1_334 = $signed(_T_59429); // @[Modules.scala 160:64:@5148.4]
  assign buffer_1_62 = {{8{_T_57650[5]}},_T_57650}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_63 = {{9{_T_57657[4]}},_T_57657}; // @[Modules.scala 112:22:@8.4]
  assign _T_59431 = $signed(buffer_1_62) + $signed(buffer_1_63); // @[Modules.scala 160:64:@5150.4]
  assign _T_59432 = _T_59431[13:0]; // @[Modules.scala 160:64:@5151.4]
  assign buffer_1_335 = $signed(_T_59432); // @[Modules.scala 160:64:@5152.4]
  assign buffer_1_64 = {{9{_T_57664[4]}},_T_57664}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_65 = {{9{_T_57671[4]}},_T_57671}; // @[Modules.scala 112:22:@8.4]
  assign _T_59434 = $signed(buffer_1_64) + $signed(buffer_1_65); // @[Modules.scala 160:64:@5154.4]
  assign _T_59435 = _T_59434[13:0]; // @[Modules.scala 160:64:@5155.4]
  assign buffer_1_336 = $signed(_T_59435); // @[Modules.scala 160:64:@5156.4]
  assign buffer_1_66 = {{8{_T_57678[5]}},_T_57678}; // @[Modules.scala 112:22:@8.4]
  assign _T_59437 = $signed(buffer_1_66) + $signed(buffer_0_66); // @[Modules.scala 160:64:@5158.4]
  assign _T_59438 = _T_59437[13:0]; // @[Modules.scala 160:64:@5159.4]
  assign buffer_1_337 = $signed(_T_59438); // @[Modules.scala 160:64:@5160.4]
  assign _T_59440 = $signed(buffer_0_67) + $signed(buffer_0_68); // @[Modules.scala 160:64:@5162.4]
  assign _T_59441 = _T_59440[13:0]; // @[Modules.scala 160:64:@5163.4]
  assign buffer_1_338 = $signed(_T_59441); // @[Modules.scala 160:64:@5164.4]
  assign buffer_1_70 = {{9{_T_57706[4]}},_T_57706}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_71 = {{8{_T_57713[5]}},_T_57713}; // @[Modules.scala 112:22:@8.4]
  assign _T_59443 = $signed(buffer_1_70) + $signed(buffer_1_71); // @[Modules.scala 160:64:@5166.4]
  assign _T_59444 = _T_59443[13:0]; // @[Modules.scala 160:64:@5167.4]
  assign buffer_1_339 = $signed(_T_59444); // @[Modules.scala 160:64:@5168.4]
  assign buffer_1_72 = {{8{_T_57720[5]}},_T_57720}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_73 = {{8{_T_57727[5]}},_T_57727}; // @[Modules.scala 112:22:@8.4]
  assign _T_59446 = $signed(buffer_1_72) + $signed(buffer_1_73); // @[Modules.scala 160:64:@5170.4]
  assign _T_59447 = _T_59446[13:0]; // @[Modules.scala 160:64:@5171.4]
  assign buffer_1_340 = $signed(_T_59447); // @[Modules.scala 160:64:@5172.4]
  assign buffer_1_74 = {{8{_T_57734[5]}},_T_57734}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_75 = {{8{_T_57741[5]}},_T_57741}; // @[Modules.scala 112:22:@8.4]
  assign _T_59449 = $signed(buffer_1_74) + $signed(buffer_1_75); // @[Modules.scala 160:64:@5174.4]
  assign _T_59450 = _T_59449[13:0]; // @[Modules.scala 160:64:@5175.4]
  assign buffer_1_341 = $signed(_T_59450); // @[Modules.scala 160:64:@5176.4]
  assign _T_59452 = $signed(buffer_0_73) + $signed(buffer_0_74); // @[Modules.scala 160:64:@5178.4]
  assign _T_59453 = _T_59452[13:0]; // @[Modules.scala 160:64:@5179.4]
  assign buffer_1_342 = $signed(_T_59453); // @[Modules.scala 160:64:@5180.4]
  assign buffer_1_78 = {{9{_T_57762[4]}},_T_57762}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_79 = {{8{_T_57769[5]}},_T_57769}; // @[Modules.scala 112:22:@8.4]
  assign _T_59455 = $signed(buffer_1_78) + $signed(buffer_1_79); // @[Modules.scala 160:64:@5182.4]
  assign _T_59456 = _T_59455[13:0]; // @[Modules.scala 160:64:@5183.4]
  assign buffer_1_343 = $signed(_T_59456); // @[Modules.scala 160:64:@5184.4]
  assign buffer_1_80 = {{8{_T_57776[5]}},_T_57776}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_81 = {{8{_T_57783[5]}},_T_57783}; // @[Modules.scala 112:22:@8.4]
  assign _T_59458 = $signed(buffer_1_80) + $signed(buffer_1_81); // @[Modules.scala 160:64:@5186.4]
  assign _T_59459 = _T_59458[13:0]; // @[Modules.scala 160:64:@5187.4]
  assign buffer_1_344 = $signed(_T_59459); // @[Modules.scala 160:64:@5188.4]
  assign buffer_1_82 = {{8{_T_57790[5]}},_T_57790}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_83 = {{9{_T_57797[4]}},_T_57797}; // @[Modules.scala 112:22:@8.4]
  assign _T_59461 = $signed(buffer_1_82) + $signed(buffer_1_83); // @[Modules.scala 160:64:@5190.4]
  assign _T_59462 = _T_59461[13:0]; // @[Modules.scala 160:64:@5191.4]
  assign buffer_1_345 = $signed(_T_59462); // @[Modules.scala 160:64:@5192.4]
  assign buffer_1_84 = {{8{_T_57804[5]}},_T_57804}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_85 = {{8{_T_57811[5]}},_T_57811}; // @[Modules.scala 112:22:@8.4]
  assign _T_59464 = $signed(buffer_1_84) + $signed(buffer_1_85); // @[Modules.scala 160:64:@5194.4]
  assign _T_59465 = _T_59464[13:0]; // @[Modules.scala 160:64:@5195.4]
  assign buffer_1_346 = $signed(_T_59465); // @[Modules.scala 160:64:@5196.4]
  assign buffer_1_86 = {{8{_T_57818[5]}},_T_57818}; // @[Modules.scala 112:22:@8.4]
  assign _T_59467 = $signed(buffer_1_86) + $signed(buffer_0_83); // @[Modules.scala 160:64:@5198.4]
  assign _T_59468 = _T_59467[13:0]; // @[Modules.scala 160:64:@5199.4]
  assign buffer_1_347 = $signed(_T_59468); // @[Modules.scala 160:64:@5200.4]
  assign buffer_1_91 = {{8{_T_57853[5]}},_T_57853}; // @[Modules.scala 112:22:@8.4]
  assign _T_59473 = $signed(buffer_0_86) + $signed(buffer_1_91); // @[Modules.scala 160:64:@5206.4]
  assign _T_59474 = _T_59473[13:0]; // @[Modules.scala 160:64:@5207.4]
  assign buffer_1_349 = $signed(_T_59474); // @[Modules.scala 160:64:@5208.4]
  assign buffer_1_92 = {{8{_T_57860[5]}},_T_57860}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_93 = {{8{_T_57867[5]}},_T_57867}; // @[Modules.scala 112:22:@8.4]
  assign _T_59476 = $signed(buffer_1_92) + $signed(buffer_1_93); // @[Modules.scala 160:64:@5210.4]
  assign _T_59477 = _T_59476[13:0]; // @[Modules.scala 160:64:@5211.4]
  assign buffer_1_350 = $signed(_T_59477); // @[Modules.scala 160:64:@5212.4]
  assign buffer_1_94 = {{9{_T_57874[4]}},_T_57874}; // @[Modules.scala 112:22:@8.4]
  assign _T_59479 = $signed(buffer_1_94) + $signed(buffer_0_91); // @[Modules.scala 160:64:@5214.4]
  assign _T_59480 = _T_59479[13:0]; // @[Modules.scala 160:64:@5215.4]
  assign buffer_1_351 = $signed(_T_59480); // @[Modules.scala 160:64:@5216.4]
  assign buffer_1_96 = {{8{_T_57888[5]}},_T_57888}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_97 = {{8{_T_57895[5]}},_T_57895}; // @[Modules.scala 112:22:@8.4]
  assign _T_59482 = $signed(buffer_1_96) + $signed(buffer_1_97); // @[Modules.scala 160:64:@5218.4]
  assign _T_59483 = _T_59482[13:0]; // @[Modules.scala 160:64:@5219.4]
  assign buffer_1_352 = $signed(_T_59483); // @[Modules.scala 160:64:@5220.4]
  assign buffer_1_98 = {{8{_T_57902[5]}},_T_57902}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_99 = {{8{_T_57909[5]}},_T_57909}; // @[Modules.scala 112:22:@8.4]
  assign _T_59485 = $signed(buffer_1_98) + $signed(buffer_1_99); // @[Modules.scala 160:64:@5222.4]
  assign _T_59486 = _T_59485[13:0]; // @[Modules.scala 160:64:@5223.4]
  assign buffer_1_353 = $signed(_T_59486); // @[Modules.scala 160:64:@5224.4]
  assign _T_59488 = $signed(buffer_0_97) + $signed(buffer_0_98); // @[Modules.scala 160:64:@5226.4]
  assign _T_59489 = _T_59488[13:0]; // @[Modules.scala 160:64:@5227.4]
  assign buffer_1_354 = $signed(_T_59489); // @[Modules.scala 160:64:@5228.4]
  assign buffer_1_102 = {{8{_T_57930[5]}},_T_57930}; // @[Modules.scala 112:22:@8.4]
  assign _T_59491 = $signed(buffer_1_102) + $signed(buffer_0_100); // @[Modules.scala 160:64:@5230.4]
  assign _T_59492 = _T_59491[13:0]; // @[Modules.scala 160:64:@5231.4]
  assign buffer_1_355 = $signed(_T_59492); // @[Modules.scala 160:64:@5232.4]
  assign buffer_1_104 = {{8{_T_57944[5]}},_T_57944}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_105 = {{9{_T_57951[4]}},_T_57951}; // @[Modules.scala 112:22:@8.4]
  assign _T_59494 = $signed(buffer_1_104) + $signed(buffer_1_105); // @[Modules.scala 160:64:@5234.4]
  assign _T_59495 = _T_59494[13:0]; // @[Modules.scala 160:64:@5235.4]
  assign buffer_1_356 = $signed(_T_59495); // @[Modules.scala 160:64:@5236.4]
  assign buffer_1_106 = {{9{_T_57958[4]}},_T_57958}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_107 = {{8{_T_57965[5]}},_T_57965}; // @[Modules.scala 112:22:@8.4]
  assign _T_59497 = $signed(buffer_1_106) + $signed(buffer_1_107); // @[Modules.scala 160:64:@5238.4]
  assign _T_59498 = _T_59497[13:0]; // @[Modules.scala 160:64:@5239.4]
  assign buffer_1_357 = $signed(_T_59498); // @[Modules.scala 160:64:@5240.4]
  assign buffer_1_108 = {{8{_T_57972[5]}},_T_57972}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_109 = {{8{_T_57979[5]}},_T_57979}; // @[Modules.scala 112:22:@8.4]
  assign _T_59500 = $signed(buffer_1_108) + $signed(buffer_1_109); // @[Modules.scala 160:64:@5242.4]
  assign _T_59501 = _T_59500[13:0]; // @[Modules.scala 160:64:@5243.4]
  assign buffer_1_358 = $signed(_T_59501); // @[Modules.scala 160:64:@5244.4]
  assign buffer_1_110 = {{8{_T_57986[5]}},_T_57986}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_111 = {{8{_T_57993[5]}},_T_57993}; // @[Modules.scala 112:22:@8.4]
  assign _T_59503 = $signed(buffer_1_110) + $signed(buffer_1_111); // @[Modules.scala 160:64:@5246.4]
  assign _T_59504 = _T_59503[13:0]; // @[Modules.scala 160:64:@5247.4]
  assign buffer_1_359 = $signed(_T_59504); // @[Modules.scala 160:64:@5248.4]
  assign buffer_1_112 = {{9{_T_58000[4]}},_T_58000}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_113 = {{9{_T_58007[4]}},_T_58007}; // @[Modules.scala 112:22:@8.4]
  assign _T_59506 = $signed(buffer_1_112) + $signed(buffer_1_113); // @[Modules.scala 160:64:@5250.4]
  assign _T_59507 = _T_59506[13:0]; // @[Modules.scala 160:64:@5251.4]
  assign buffer_1_360 = $signed(_T_59507); // @[Modules.scala 160:64:@5252.4]
  assign buffer_1_114 = {{8{_T_58014[5]}},_T_58014}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_115 = {{8{_T_58021[5]}},_T_58021}; // @[Modules.scala 112:22:@8.4]
  assign _T_59509 = $signed(buffer_1_114) + $signed(buffer_1_115); // @[Modules.scala 160:64:@5254.4]
  assign _T_59510 = _T_59509[13:0]; // @[Modules.scala 160:64:@5255.4]
  assign buffer_1_361 = $signed(_T_59510); // @[Modules.scala 160:64:@5256.4]
  assign buffer_1_116 = {{8{_T_58028[5]}},_T_58028}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_117 = {{8{_T_58035[5]}},_T_58035}; // @[Modules.scala 112:22:@8.4]
  assign _T_59512 = $signed(buffer_1_116) + $signed(buffer_1_117); // @[Modules.scala 160:64:@5258.4]
  assign _T_59513 = _T_59512[13:0]; // @[Modules.scala 160:64:@5259.4]
  assign buffer_1_362 = $signed(_T_59513); // @[Modules.scala 160:64:@5260.4]
  assign buffer_1_118 = {{9{_T_58042[4]}},_T_58042}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_119 = {{9{_T_58049[4]}},_T_58049}; // @[Modules.scala 112:22:@8.4]
  assign _T_59515 = $signed(buffer_1_118) + $signed(buffer_1_119); // @[Modules.scala 160:64:@5262.4]
  assign _T_59516 = _T_59515[13:0]; // @[Modules.scala 160:64:@5263.4]
  assign buffer_1_363 = $signed(_T_59516); // @[Modules.scala 160:64:@5264.4]
  assign buffer_1_120 = {{8{_T_58056[5]}},_T_58056}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_121 = {{8{_T_58063[5]}},_T_58063}; // @[Modules.scala 112:22:@8.4]
  assign _T_59518 = $signed(buffer_1_120) + $signed(buffer_1_121); // @[Modules.scala 160:64:@5266.4]
  assign _T_59519 = _T_59518[13:0]; // @[Modules.scala 160:64:@5267.4]
  assign buffer_1_364 = $signed(_T_59519); // @[Modules.scala 160:64:@5268.4]
  assign buffer_1_122 = {{8{_T_58070[5]}},_T_58070}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_123 = {{8{_T_58077[5]}},_T_58077}; // @[Modules.scala 112:22:@8.4]
  assign _T_59521 = $signed(buffer_1_122) + $signed(buffer_1_123); // @[Modules.scala 160:64:@5270.4]
  assign _T_59522 = _T_59521[13:0]; // @[Modules.scala 160:64:@5271.4]
  assign buffer_1_365 = $signed(_T_59522); // @[Modules.scala 160:64:@5272.4]
  assign buffer_1_124 = {{8{_T_58084[5]}},_T_58084}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_125 = {{9{_T_58091[4]}},_T_58091}; // @[Modules.scala 112:22:@8.4]
  assign _T_59524 = $signed(buffer_1_124) + $signed(buffer_1_125); // @[Modules.scala 160:64:@5274.4]
  assign _T_59525 = _T_59524[13:0]; // @[Modules.scala 160:64:@5275.4]
  assign buffer_1_366 = $signed(_T_59525); // @[Modules.scala 160:64:@5276.4]
  assign buffer_1_126 = {{9{_T_58098[4]}},_T_58098}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_127 = {{8{_T_58105[5]}},_T_58105}; // @[Modules.scala 112:22:@8.4]
  assign _T_59527 = $signed(buffer_1_126) + $signed(buffer_1_127); // @[Modules.scala 160:64:@5278.4]
  assign _T_59528 = _T_59527[13:0]; // @[Modules.scala 160:64:@5279.4]
  assign buffer_1_367 = $signed(_T_59528); // @[Modules.scala 160:64:@5280.4]
  assign buffer_1_128 = {{9{_T_58112[4]}},_T_58112}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_129 = {{8{_T_58119[5]}},_T_58119}; // @[Modules.scala 112:22:@8.4]
  assign _T_59530 = $signed(buffer_1_128) + $signed(buffer_1_129); // @[Modules.scala 160:64:@5282.4]
  assign _T_59531 = _T_59530[13:0]; // @[Modules.scala 160:64:@5283.4]
  assign buffer_1_368 = $signed(_T_59531); // @[Modules.scala 160:64:@5284.4]
  assign buffer_1_130 = {{8{_T_58126[5]}},_T_58126}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_131 = {{9{_T_58133[4]}},_T_58133}; // @[Modules.scala 112:22:@8.4]
  assign _T_59533 = $signed(buffer_1_130) + $signed(buffer_1_131); // @[Modules.scala 160:64:@5286.4]
  assign _T_59534 = _T_59533[13:0]; // @[Modules.scala 160:64:@5287.4]
  assign buffer_1_369 = $signed(_T_59534); // @[Modules.scala 160:64:@5288.4]
  assign buffer_1_132 = {{9{_T_58140[4]}},_T_58140}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_133 = {{8{_T_58147[5]}},_T_58147}; // @[Modules.scala 112:22:@8.4]
  assign _T_59536 = $signed(buffer_1_132) + $signed(buffer_1_133); // @[Modules.scala 160:64:@5290.4]
  assign _T_59537 = _T_59536[13:0]; // @[Modules.scala 160:64:@5291.4]
  assign buffer_1_370 = $signed(_T_59537); // @[Modules.scala 160:64:@5292.4]
  assign buffer_1_134 = {{8{_T_58154[5]}},_T_58154}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_135 = {{8{_T_58161[5]}},_T_58161}; // @[Modules.scala 112:22:@8.4]
  assign _T_59539 = $signed(buffer_1_134) + $signed(buffer_1_135); // @[Modules.scala 160:64:@5294.4]
  assign _T_59540 = _T_59539[13:0]; // @[Modules.scala 160:64:@5295.4]
  assign buffer_1_371 = $signed(_T_59540); // @[Modules.scala 160:64:@5296.4]
  assign buffer_1_136 = {{8{_T_58168[5]}},_T_58168}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_137 = {{8{_T_58175[5]}},_T_58175}; // @[Modules.scala 112:22:@8.4]
  assign _T_59542 = $signed(buffer_1_136) + $signed(buffer_1_137); // @[Modules.scala 160:64:@5298.4]
  assign _T_59543 = _T_59542[13:0]; // @[Modules.scala 160:64:@5299.4]
  assign buffer_1_372 = $signed(_T_59543); // @[Modules.scala 160:64:@5300.4]
  assign buffer_1_138 = {{8{_T_58182[5]}},_T_58182}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_139 = {{8{_T_58189[5]}},_T_58189}; // @[Modules.scala 112:22:@8.4]
  assign _T_59545 = $signed(buffer_1_138) + $signed(buffer_1_139); // @[Modules.scala 160:64:@5302.4]
  assign _T_59546 = _T_59545[13:0]; // @[Modules.scala 160:64:@5303.4]
  assign buffer_1_373 = $signed(_T_59546); // @[Modules.scala 160:64:@5304.4]
  assign buffer_1_140 = {{9{_T_58196[4]}},_T_58196}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_141 = {{8{_T_58203[5]}},_T_58203}; // @[Modules.scala 112:22:@8.4]
  assign _T_59548 = $signed(buffer_1_140) + $signed(buffer_1_141); // @[Modules.scala 160:64:@5306.4]
  assign _T_59549 = _T_59548[13:0]; // @[Modules.scala 160:64:@5307.4]
  assign buffer_1_374 = $signed(_T_59549); // @[Modules.scala 160:64:@5308.4]
  assign buffer_1_142 = {{8{_T_58210[5]}},_T_58210}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_143 = {{8{_T_58217[5]}},_T_58217}; // @[Modules.scala 112:22:@8.4]
  assign _T_59551 = $signed(buffer_1_142) + $signed(buffer_1_143); // @[Modules.scala 160:64:@5310.4]
  assign _T_59552 = _T_59551[13:0]; // @[Modules.scala 160:64:@5311.4]
  assign buffer_1_375 = $signed(_T_59552); // @[Modules.scala 160:64:@5312.4]
  assign buffer_1_144 = {{9{_T_58224[4]}},_T_58224}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_145 = {{8{_T_58231[5]}},_T_58231}; // @[Modules.scala 112:22:@8.4]
  assign _T_59554 = $signed(buffer_1_144) + $signed(buffer_1_145); // @[Modules.scala 160:64:@5314.4]
  assign _T_59555 = _T_59554[13:0]; // @[Modules.scala 160:64:@5315.4]
  assign buffer_1_376 = $signed(_T_59555); // @[Modules.scala 160:64:@5316.4]
  assign buffer_1_146 = {{8{_T_58238[5]}},_T_58238}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_147 = {{8{_T_58245[5]}},_T_58245}; // @[Modules.scala 112:22:@8.4]
  assign _T_59557 = $signed(buffer_1_146) + $signed(buffer_1_147); // @[Modules.scala 160:64:@5318.4]
  assign _T_59558 = _T_59557[13:0]; // @[Modules.scala 160:64:@5319.4]
  assign buffer_1_377 = $signed(_T_59558); // @[Modules.scala 160:64:@5320.4]
  assign buffer_1_148 = {{8{_T_58252[5]}},_T_58252}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_149 = {{9{_T_58259[4]}},_T_58259}; // @[Modules.scala 112:22:@8.4]
  assign _T_59560 = $signed(buffer_1_148) + $signed(buffer_1_149); // @[Modules.scala 160:64:@5322.4]
  assign _T_59561 = _T_59560[13:0]; // @[Modules.scala 160:64:@5323.4]
  assign buffer_1_378 = $signed(_T_59561); // @[Modules.scala 160:64:@5324.4]
  assign buffer_1_150 = {{9{_T_58266[4]}},_T_58266}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_151 = {{8{_T_58273[5]}},_T_58273}; // @[Modules.scala 112:22:@8.4]
  assign _T_59563 = $signed(buffer_1_150) + $signed(buffer_1_151); // @[Modules.scala 160:64:@5326.4]
  assign _T_59564 = _T_59563[13:0]; // @[Modules.scala 160:64:@5327.4]
  assign buffer_1_379 = $signed(_T_59564); // @[Modules.scala 160:64:@5328.4]
  assign buffer_1_152 = {{8{_T_58280[5]}},_T_58280}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_153 = {{8{_T_58287[5]}},_T_58287}; // @[Modules.scala 112:22:@8.4]
  assign _T_59566 = $signed(buffer_1_152) + $signed(buffer_1_153); // @[Modules.scala 160:64:@5330.4]
  assign _T_59567 = _T_59566[13:0]; // @[Modules.scala 160:64:@5331.4]
  assign buffer_1_380 = $signed(_T_59567); // @[Modules.scala 160:64:@5332.4]
  assign buffer_1_154 = {{8{_T_58294[5]}},_T_58294}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_155 = {{8{_T_58301[5]}},_T_58301}; // @[Modules.scala 112:22:@8.4]
  assign _T_59569 = $signed(buffer_1_154) + $signed(buffer_1_155); // @[Modules.scala 160:64:@5334.4]
  assign _T_59570 = _T_59569[13:0]; // @[Modules.scala 160:64:@5335.4]
  assign buffer_1_381 = $signed(_T_59570); // @[Modules.scala 160:64:@5336.4]
  assign buffer_1_156 = {{9{_T_58308[4]}},_T_58308}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_157 = {{8{_T_58315[5]}},_T_58315}; // @[Modules.scala 112:22:@8.4]
  assign _T_59572 = $signed(buffer_1_156) + $signed(buffer_1_157); // @[Modules.scala 160:64:@5338.4]
  assign _T_59573 = _T_59572[13:0]; // @[Modules.scala 160:64:@5339.4]
  assign buffer_1_382 = $signed(_T_59573); // @[Modules.scala 160:64:@5340.4]
  assign buffer_1_159 = {{9{_T_58329[4]}},_T_58329}; // @[Modules.scala 112:22:@8.4]
  assign _T_59575 = $signed(buffer_0_157) + $signed(buffer_1_159); // @[Modules.scala 160:64:@5342.4]
  assign _T_59576 = _T_59575[13:0]; // @[Modules.scala 160:64:@5343.4]
  assign buffer_1_383 = $signed(_T_59576); // @[Modules.scala 160:64:@5344.4]
  assign buffer_1_160 = {{9{_T_58336[4]}},_T_58336}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_161 = {{9{_T_58343[4]}},_T_58343}; // @[Modules.scala 112:22:@8.4]
  assign _T_59578 = $signed(buffer_1_160) + $signed(buffer_1_161); // @[Modules.scala 160:64:@5346.4]
  assign _T_59579 = _T_59578[13:0]; // @[Modules.scala 160:64:@5347.4]
  assign buffer_1_384 = $signed(_T_59579); // @[Modules.scala 160:64:@5348.4]
  assign buffer_1_162 = {{9{_T_58350[4]}},_T_58350}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_163 = {{9{_T_58357[4]}},_T_58357}; // @[Modules.scala 112:22:@8.4]
  assign _T_59581 = $signed(buffer_1_162) + $signed(buffer_1_163); // @[Modules.scala 160:64:@5350.4]
  assign _T_59582 = _T_59581[13:0]; // @[Modules.scala 160:64:@5351.4]
  assign buffer_1_385 = $signed(_T_59582); // @[Modules.scala 160:64:@5352.4]
  assign buffer_1_164 = {{8{_T_58364[5]}},_T_58364}; // @[Modules.scala 112:22:@8.4]
  assign _T_59584 = $signed(buffer_1_164) + $signed(buffer_0_164); // @[Modules.scala 160:64:@5354.4]
  assign _T_59585 = _T_59584[13:0]; // @[Modules.scala 160:64:@5355.4]
  assign buffer_1_386 = $signed(_T_59585); // @[Modules.scala 160:64:@5356.4]
  assign buffer_1_166 = {{9{_T_58378[4]}},_T_58378}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_167 = {{9{_T_58385[4]}},_T_58385}; // @[Modules.scala 112:22:@8.4]
  assign _T_59587 = $signed(buffer_1_166) + $signed(buffer_1_167); // @[Modules.scala 160:64:@5358.4]
  assign _T_59588 = _T_59587[13:0]; // @[Modules.scala 160:64:@5359.4]
  assign buffer_1_387 = $signed(_T_59588); // @[Modules.scala 160:64:@5360.4]
  assign buffer_1_168 = {{8{_T_58392[5]}},_T_58392}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_169 = {{8{_T_58399[5]}},_T_58399}; // @[Modules.scala 112:22:@8.4]
  assign _T_59590 = $signed(buffer_1_168) + $signed(buffer_1_169); // @[Modules.scala 160:64:@5362.4]
  assign _T_59591 = _T_59590[13:0]; // @[Modules.scala 160:64:@5363.4]
  assign buffer_1_388 = $signed(_T_59591); // @[Modules.scala 160:64:@5364.4]
  assign buffer_1_170 = {{8{_T_58406[5]}},_T_58406}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_171 = {{9{_T_58413[4]}},_T_58413}; // @[Modules.scala 112:22:@8.4]
  assign _T_59593 = $signed(buffer_1_170) + $signed(buffer_1_171); // @[Modules.scala 160:64:@5366.4]
  assign _T_59594 = _T_59593[13:0]; // @[Modules.scala 160:64:@5367.4]
  assign buffer_1_389 = $signed(_T_59594); // @[Modules.scala 160:64:@5368.4]
  assign buffer_1_172 = {{9{_T_58420[4]}},_T_58420}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_173 = {{8{_T_58427[5]}},_T_58427}; // @[Modules.scala 112:22:@8.4]
  assign _T_59596 = $signed(buffer_1_172) + $signed(buffer_1_173); // @[Modules.scala 160:64:@5370.4]
  assign _T_59597 = _T_59596[13:0]; // @[Modules.scala 160:64:@5371.4]
  assign buffer_1_390 = $signed(_T_59597); // @[Modules.scala 160:64:@5372.4]
  assign buffer_1_174 = {{8{_T_58434[5]}},_T_58434}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_175 = {{8{_T_58441[5]}},_T_58441}; // @[Modules.scala 112:22:@8.4]
  assign _T_59599 = $signed(buffer_1_174) + $signed(buffer_1_175); // @[Modules.scala 160:64:@5374.4]
  assign _T_59600 = _T_59599[13:0]; // @[Modules.scala 160:64:@5375.4]
  assign buffer_1_391 = $signed(_T_59600); // @[Modules.scala 160:64:@5376.4]
  assign buffer_1_176 = {{9{_T_58448[4]}},_T_58448}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_177 = {{9{_T_58455[4]}},_T_58455}; // @[Modules.scala 112:22:@8.4]
  assign _T_59602 = $signed(buffer_1_176) + $signed(buffer_1_177); // @[Modules.scala 160:64:@5378.4]
  assign _T_59603 = _T_59602[13:0]; // @[Modules.scala 160:64:@5379.4]
  assign buffer_1_392 = $signed(_T_59603); // @[Modules.scala 160:64:@5380.4]
  assign buffer_1_178 = {{9{_T_58462[4]}},_T_58462}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_179 = {{9{_T_58469[4]}},_T_58469}; // @[Modules.scala 112:22:@8.4]
  assign _T_59605 = $signed(buffer_1_178) + $signed(buffer_1_179); // @[Modules.scala 160:64:@5382.4]
  assign _T_59606 = _T_59605[13:0]; // @[Modules.scala 160:64:@5383.4]
  assign buffer_1_393 = $signed(_T_59606); // @[Modules.scala 160:64:@5384.4]
  assign buffer_1_180 = {{9{_T_58476[4]}},_T_58476}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_181 = {{8{_T_58483[5]}},_T_58483}; // @[Modules.scala 112:22:@8.4]
  assign _T_59608 = $signed(buffer_1_180) + $signed(buffer_1_181); // @[Modules.scala 160:64:@5386.4]
  assign _T_59609 = _T_59608[13:0]; // @[Modules.scala 160:64:@5387.4]
  assign buffer_1_394 = $signed(_T_59609); // @[Modules.scala 160:64:@5388.4]
  assign buffer_1_182 = {{8{_T_58490[5]}},_T_58490}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_183 = {{9{_T_58497[4]}},_T_58497}; // @[Modules.scala 112:22:@8.4]
  assign _T_59611 = $signed(buffer_1_182) + $signed(buffer_1_183); // @[Modules.scala 160:64:@5390.4]
  assign _T_59612 = _T_59611[13:0]; // @[Modules.scala 160:64:@5391.4]
  assign buffer_1_395 = $signed(_T_59612); // @[Modules.scala 160:64:@5392.4]
  assign buffer_1_184 = {{8{_T_58504[5]}},_T_58504}; // @[Modules.scala 112:22:@8.4]
  assign _T_59614 = $signed(buffer_1_184) + $signed(buffer_0_184); // @[Modules.scala 160:64:@5394.4]
  assign _T_59615 = _T_59614[13:0]; // @[Modules.scala 160:64:@5395.4]
  assign buffer_1_396 = $signed(_T_59615); // @[Modules.scala 160:64:@5396.4]
  assign buffer_1_187 = {{9{_T_58525[4]}},_T_58525}; // @[Modules.scala 112:22:@8.4]
  assign _T_59617 = $signed(buffer_0_185) + $signed(buffer_1_187); // @[Modules.scala 160:64:@5398.4]
  assign _T_59618 = _T_59617[13:0]; // @[Modules.scala 160:64:@5399.4]
  assign buffer_1_397 = $signed(_T_59618); // @[Modules.scala 160:64:@5400.4]
  assign buffer_1_188 = {{9{_T_58532[4]}},_T_58532}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_189 = {{9{_T_58539[4]}},_T_58539}; // @[Modules.scala 112:22:@8.4]
  assign _T_59620 = $signed(buffer_1_188) + $signed(buffer_1_189); // @[Modules.scala 160:64:@5402.4]
  assign _T_59621 = _T_59620[13:0]; // @[Modules.scala 160:64:@5403.4]
  assign buffer_1_398 = $signed(_T_59621); // @[Modules.scala 160:64:@5404.4]
  assign buffer_1_190 = {{9{_T_58546[4]}},_T_58546}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_191 = {{9{_T_58553[4]}},_T_58553}; // @[Modules.scala 112:22:@8.4]
  assign _T_59623 = $signed(buffer_1_190) + $signed(buffer_1_191); // @[Modules.scala 160:64:@5406.4]
  assign _T_59624 = _T_59623[13:0]; // @[Modules.scala 160:64:@5407.4]
  assign buffer_1_399 = $signed(_T_59624); // @[Modules.scala 160:64:@5408.4]
  assign buffer_1_192 = {{8{_T_58560[5]}},_T_58560}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_193 = {{9{_T_58567[4]}},_T_58567}; // @[Modules.scala 112:22:@8.4]
  assign _T_59626 = $signed(buffer_1_192) + $signed(buffer_1_193); // @[Modules.scala 160:64:@5410.4]
  assign _T_59627 = _T_59626[13:0]; // @[Modules.scala 160:64:@5411.4]
  assign buffer_1_400 = $signed(_T_59627); // @[Modules.scala 160:64:@5412.4]
  assign buffer_1_194 = {{8{_T_58574[5]}},_T_58574}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_195 = {{9{_T_58581[4]}},_T_58581}; // @[Modules.scala 112:22:@8.4]
  assign _T_59629 = $signed(buffer_1_194) + $signed(buffer_1_195); // @[Modules.scala 160:64:@5414.4]
  assign _T_59630 = _T_59629[13:0]; // @[Modules.scala 160:64:@5415.4]
  assign buffer_1_401 = $signed(_T_59630); // @[Modules.scala 160:64:@5416.4]
  assign buffer_1_196 = {{8{_T_58588[5]}},_T_58588}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_197 = {{8{_T_58595[5]}},_T_58595}; // @[Modules.scala 112:22:@8.4]
  assign _T_59632 = $signed(buffer_1_196) + $signed(buffer_1_197); // @[Modules.scala 160:64:@5418.4]
  assign _T_59633 = _T_59632[13:0]; // @[Modules.scala 160:64:@5419.4]
  assign buffer_1_402 = $signed(_T_59633); // @[Modules.scala 160:64:@5420.4]
  assign buffer_1_198 = {{8{_T_58602[5]}},_T_58602}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_199 = {{9{_T_58609[4]}},_T_58609}; // @[Modules.scala 112:22:@8.4]
  assign _T_59635 = $signed(buffer_1_198) + $signed(buffer_1_199); // @[Modules.scala 160:64:@5422.4]
  assign _T_59636 = _T_59635[13:0]; // @[Modules.scala 160:64:@5423.4]
  assign buffer_1_403 = $signed(_T_59636); // @[Modules.scala 160:64:@5424.4]
  assign buffer_1_200 = {{9{_T_58616[4]}},_T_58616}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_201 = {{9{_T_58623[4]}},_T_58623}; // @[Modules.scala 112:22:@8.4]
  assign _T_59638 = $signed(buffer_1_200) + $signed(buffer_1_201); // @[Modules.scala 160:64:@5426.4]
  assign _T_59639 = _T_59638[13:0]; // @[Modules.scala 160:64:@5427.4]
  assign buffer_1_404 = $signed(_T_59639); // @[Modules.scala 160:64:@5428.4]
  assign buffer_1_202 = {{9{_T_58630[4]}},_T_58630}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_203 = {{8{_T_58637[5]}},_T_58637}; // @[Modules.scala 112:22:@8.4]
  assign _T_59641 = $signed(buffer_1_202) + $signed(buffer_1_203); // @[Modules.scala 160:64:@5430.4]
  assign _T_59642 = _T_59641[13:0]; // @[Modules.scala 160:64:@5431.4]
  assign buffer_1_405 = $signed(_T_59642); // @[Modules.scala 160:64:@5432.4]
  assign buffer_1_204 = {{9{_T_58644[4]}},_T_58644}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_205 = {{9{_T_58651[4]}},_T_58651}; // @[Modules.scala 112:22:@8.4]
  assign _T_59644 = $signed(buffer_1_204) + $signed(buffer_1_205); // @[Modules.scala 160:64:@5434.4]
  assign _T_59645 = _T_59644[13:0]; // @[Modules.scala 160:64:@5435.4]
  assign buffer_1_406 = $signed(_T_59645); // @[Modules.scala 160:64:@5436.4]
  assign buffer_1_206 = {{8{_T_58658[5]}},_T_58658}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_207 = {{8{_T_58665[5]}},_T_58665}; // @[Modules.scala 112:22:@8.4]
  assign _T_59647 = $signed(buffer_1_206) + $signed(buffer_1_207); // @[Modules.scala 160:64:@5438.4]
  assign _T_59648 = _T_59647[13:0]; // @[Modules.scala 160:64:@5439.4]
  assign buffer_1_407 = $signed(_T_59648); // @[Modules.scala 160:64:@5440.4]
  assign buffer_1_208 = {{8{_T_58672[5]}},_T_58672}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_209 = {{9{_T_58679[4]}},_T_58679}; // @[Modules.scala 112:22:@8.4]
  assign _T_59650 = $signed(buffer_1_208) + $signed(buffer_1_209); // @[Modules.scala 160:64:@5442.4]
  assign _T_59651 = _T_59650[13:0]; // @[Modules.scala 160:64:@5443.4]
  assign buffer_1_408 = $signed(_T_59651); // @[Modules.scala 160:64:@5444.4]
  assign buffer_1_210 = {{9{_T_58686[4]}},_T_58686}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_211 = {{9{_T_58693[4]}},_T_58693}; // @[Modules.scala 112:22:@8.4]
  assign _T_59653 = $signed(buffer_1_210) + $signed(buffer_1_211); // @[Modules.scala 160:64:@5446.4]
  assign _T_59654 = _T_59653[13:0]; // @[Modules.scala 160:64:@5447.4]
  assign buffer_1_409 = $signed(_T_59654); // @[Modules.scala 160:64:@5448.4]
  assign buffer_1_212 = {{9{_T_58700[4]}},_T_58700}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_213 = {{8{_T_58707[5]}},_T_58707}; // @[Modules.scala 112:22:@8.4]
  assign _T_59656 = $signed(buffer_1_212) + $signed(buffer_1_213); // @[Modules.scala 160:64:@5450.4]
  assign _T_59657 = _T_59656[13:0]; // @[Modules.scala 160:64:@5451.4]
  assign buffer_1_410 = $signed(_T_59657); // @[Modules.scala 160:64:@5452.4]
  assign buffer_1_214 = {{9{_T_58714[4]}},_T_58714}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_215 = {{8{_T_58721[5]}},_T_58721}; // @[Modules.scala 112:22:@8.4]
  assign _T_59659 = $signed(buffer_1_214) + $signed(buffer_1_215); // @[Modules.scala 160:64:@5454.4]
  assign _T_59660 = _T_59659[13:0]; // @[Modules.scala 160:64:@5455.4]
  assign buffer_1_411 = $signed(_T_59660); // @[Modules.scala 160:64:@5456.4]
  assign buffer_1_216 = {{9{_T_58728[4]}},_T_58728}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_217 = {{9{_T_58735[4]}},_T_58735}; // @[Modules.scala 112:22:@8.4]
  assign _T_59662 = $signed(buffer_1_216) + $signed(buffer_1_217); // @[Modules.scala 160:64:@5458.4]
  assign _T_59663 = _T_59662[13:0]; // @[Modules.scala 160:64:@5459.4]
  assign buffer_1_412 = $signed(_T_59663); // @[Modules.scala 160:64:@5460.4]
  assign buffer_1_218 = {{9{_T_58742[4]}},_T_58742}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_219 = {{8{_T_58749[5]}},_T_58749}; // @[Modules.scala 112:22:@8.4]
  assign _T_59665 = $signed(buffer_1_218) + $signed(buffer_1_219); // @[Modules.scala 160:64:@5462.4]
  assign _T_59666 = _T_59665[13:0]; // @[Modules.scala 160:64:@5463.4]
  assign buffer_1_413 = $signed(_T_59666); // @[Modules.scala 160:64:@5464.4]
  assign buffer_1_220 = {{8{_T_58756[5]}},_T_58756}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_221 = {{9{_T_58763[4]}},_T_58763}; // @[Modules.scala 112:22:@8.4]
  assign _T_59668 = $signed(buffer_1_220) + $signed(buffer_1_221); // @[Modules.scala 160:64:@5466.4]
  assign _T_59669 = _T_59668[13:0]; // @[Modules.scala 160:64:@5467.4]
  assign buffer_1_414 = $signed(_T_59669); // @[Modules.scala 160:64:@5468.4]
  assign buffer_1_222 = {{9{_T_58770[4]}},_T_58770}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_223 = {{8{_T_58777[5]}},_T_58777}; // @[Modules.scala 112:22:@8.4]
  assign _T_59671 = $signed(buffer_1_222) + $signed(buffer_1_223); // @[Modules.scala 160:64:@5470.4]
  assign _T_59672 = _T_59671[13:0]; // @[Modules.scala 160:64:@5471.4]
  assign buffer_1_415 = $signed(_T_59672); // @[Modules.scala 160:64:@5472.4]
  assign buffer_1_224 = {{9{_T_58784[4]}},_T_58784}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_225 = {{8{_T_58791[5]}},_T_58791}; // @[Modules.scala 112:22:@8.4]
  assign _T_59674 = $signed(buffer_1_224) + $signed(buffer_1_225); // @[Modules.scala 160:64:@5474.4]
  assign _T_59675 = _T_59674[13:0]; // @[Modules.scala 160:64:@5475.4]
  assign buffer_1_416 = $signed(_T_59675); // @[Modules.scala 160:64:@5476.4]
  assign buffer_1_226 = {{9{_T_58798[4]}},_T_58798}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_227 = {{9{_T_58805[4]}},_T_58805}; // @[Modules.scala 112:22:@8.4]
  assign _T_59677 = $signed(buffer_1_226) + $signed(buffer_1_227); // @[Modules.scala 160:64:@5478.4]
  assign _T_59678 = _T_59677[13:0]; // @[Modules.scala 160:64:@5479.4]
  assign buffer_1_417 = $signed(_T_59678); // @[Modules.scala 160:64:@5480.4]
  assign buffer_1_228 = {{8{_T_58812[5]}},_T_58812}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_229 = {{9{_T_58819[4]}},_T_58819}; // @[Modules.scala 112:22:@8.4]
  assign _T_59680 = $signed(buffer_1_228) + $signed(buffer_1_229); // @[Modules.scala 160:64:@5482.4]
  assign _T_59681 = _T_59680[13:0]; // @[Modules.scala 160:64:@5483.4]
  assign buffer_1_418 = $signed(_T_59681); // @[Modules.scala 160:64:@5484.4]
  assign buffer_1_232 = {{8{_T_58840[5]}},_T_58840}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_233 = {{8{_T_58847[5]}},_T_58847}; // @[Modules.scala 112:22:@8.4]
  assign _T_59686 = $signed(buffer_1_232) + $signed(buffer_1_233); // @[Modules.scala 160:64:@5490.4]
  assign _T_59687 = _T_59686[13:0]; // @[Modules.scala 160:64:@5491.4]
  assign buffer_1_420 = $signed(_T_59687); // @[Modules.scala 160:64:@5492.4]
  assign buffer_1_234 = {{9{_T_58854[4]}},_T_58854}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_235 = {{8{_T_58861[5]}},_T_58861}; // @[Modules.scala 112:22:@8.4]
  assign _T_59689 = $signed(buffer_1_234) + $signed(buffer_1_235); // @[Modules.scala 160:64:@5494.4]
  assign _T_59690 = _T_59689[13:0]; // @[Modules.scala 160:64:@5495.4]
  assign buffer_1_421 = $signed(_T_59690); // @[Modules.scala 160:64:@5496.4]
  assign buffer_1_236 = {{9{_T_58868[4]}},_T_58868}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_237 = {{9{_T_58875[4]}},_T_58875}; // @[Modules.scala 112:22:@8.4]
  assign _T_59692 = $signed(buffer_1_236) + $signed(buffer_1_237); // @[Modules.scala 160:64:@5498.4]
  assign _T_59693 = _T_59692[13:0]; // @[Modules.scala 160:64:@5499.4]
  assign buffer_1_422 = $signed(_T_59693); // @[Modules.scala 160:64:@5500.4]
  assign buffer_1_238 = {{9{_T_58882[4]}},_T_58882}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_239 = {{8{_T_58889[5]}},_T_58889}; // @[Modules.scala 112:22:@8.4]
  assign _T_59695 = $signed(buffer_1_238) + $signed(buffer_1_239); // @[Modules.scala 160:64:@5502.4]
  assign _T_59696 = _T_59695[13:0]; // @[Modules.scala 160:64:@5503.4]
  assign buffer_1_423 = $signed(_T_59696); // @[Modules.scala 160:64:@5504.4]
  assign buffer_1_240 = {{8{_T_58896[5]}},_T_58896}; // @[Modules.scala 112:22:@8.4]
  assign _T_59698 = $signed(buffer_1_240) + $signed(buffer_0_239); // @[Modules.scala 160:64:@5506.4]
  assign _T_59699 = _T_59698[13:0]; // @[Modules.scala 160:64:@5507.4]
  assign buffer_1_424 = $signed(_T_59699); // @[Modules.scala 160:64:@5508.4]
  assign buffer_1_243 = {{8{_T_58917[5]}},_T_58917}; // @[Modules.scala 112:22:@8.4]
  assign _T_59701 = $signed(buffer_0_240) + $signed(buffer_1_243); // @[Modules.scala 160:64:@5510.4]
  assign _T_59702 = _T_59701[13:0]; // @[Modules.scala 160:64:@5511.4]
  assign buffer_1_425 = $signed(_T_59702); // @[Modules.scala 160:64:@5512.4]
  assign buffer_1_244 = {{8{_T_58924[5]}},_T_58924}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_245 = {{9{_T_58931[4]}},_T_58931}; // @[Modules.scala 112:22:@8.4]
  assign _T_59704 = $signed(buffer_1_244) + $signed(buffer_1_245); // @[Modules.scala 160:64:@5514.4]
  assign _T_59705 = _T_59704[13:0]; // @[Modules.scala 160:64:@5515.4]
  assign buffer_1_426 = $signed(_T_59705); // @[Modules.scala 160:64:@5516.4]
  assign buffer_1_246 = {{8{_T_58938[5]}},_T_58938}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_247 = {{9{_T_58945[4]}},_T_58945}; // @[Modules.scala 112:22:@8.4]
  assign _T_59707 = $signed(buffer_1_246) + $signed(buffer_1_247); // @[Modules.scala 160:64:@5518.4]
  assign _T_59708 = _T_59707[13:0]; // @[Modules.scala 160:64:@5519.4]
  assign buffer_1_427 = $signed(_T_59708); // @[Modules.scala 160:64:@5520.4]
  assign buffer_1_248 = {{9{_T_58952[4]}},_T_58952}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_249 = {{8{_T_58959[5]}},_T_58959}; // @[Modules.scala 112:22:@8.4]
  assign _T_59710 = $signed(buffer_1_248) + $signed(buffer_1_249); // @[Modules.scala 160:64:@5522.4]
  assign _T_59711 = _T_59710[13:0]; // @[Modules.scala 160:64:@5523.4]
  assign buffer_1_428 = $signed(_T_59711); // @[Modules.scala 160:64:@5524.4]
  assign buffer_1_250 = {{8{_T_58966[5]}},_T_58966}; // @[Modules.scala 112:22:@8.4]
  assign _T_59713 = $signed(buffer_1_250) + $signed(buffer_0_251); // @[Modules.scala 160:64:@5526.4]
  assign _T_59714 = _T_59713[13:0]; // @[Modules.scala 160:64:@5527.4]
  assign buffer_1_429 = $signed(_T_59714); // @[Modules.scala 160:64:@5528.4]
  assign buffer_1_253 = {{8{_T_58987[5]}},_T_58987}; // @[Modules.scala 112:22:@8.4]
  assign _T_59716 = $signed(buffer_0_252) + $signed(buffer_1_253); // @[Modules.scala 160:64:@5530.4]
  assign _T_59717 = _T_59716[13:0]; // @[Modules.scala 160:64:@5531.4]
  assign buffer_1_430 = $signed(_T_59717); // @[Modules.scala 160:64:@5532.4]
  assign buffer_1_254 = {{9{_T_58994[4]}},_T_58994}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_255 = {{9{_T_59001[4]}},_T_59001}; // @[Modules.scala 112:22:@8.4]
  assign _T_59719 = $signed(buffer_1_254) + $signed(buffer_1_255); // @[Modules.scala 160:64:@5534.4]
  assign _T_59720 = _T_59719[13:0]; // @[Modules.scala 160:64:@5535.4]
  assign buffer_1_431 = $signed(_T_59720); // @[Modules.scala 160:64:@5536.4]
  assign buffer_1_256 = {{8{_T_59008[5]}},_T_59008}; // @[Modules.scala 112:22:@8.4]
  assign _T_59722 = $signed(buffer_1_256) + $signed(buffer_0_259); // @[Modules.scala 160:64:@5538.4]
  assign _T_59723 = _T_59722[13:0]; // @[Modules.scala 160:64:@5539.4]
  assign buffer_1_432 = $signed(_T_59723); // @[Modules.scala 160:64:@5540.4]
  assign buffer_1_258 = {{9{_T_59022[4]}},_T_59022}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_259 = {{8{_T_59029[5]}},_T_59029}; // @[Modules.scala 112:22:@8.4]
  assign _T_59725 = $signed(buffer_1_258) + $signed(buffer_1_259); // @[Modules.scala 160:64:@5542.4]
  assign _T_59726 = _T_59725[13:0]; // @[Modules.scala 160:64:@5543.4]
  assign buffer_1_433 = $signed(_T_59726); // @[Modules.scala 160:64:@5544.4]
  assign buffer_1_260 = {{8{_T_59036[5]}},_T_59036}; // @[Modules.scala 112:22:@8.4]
  assign _T_59728 = $signed(buffer_1_260) + $signed(buffer_0_262); // @[Modules.scala 160:64:@5546.4]
  assign _T_59729 = _T_59728[13:0]; // @[Modules.scala 160:64:@5547.4]
  assign buffer_1_434 = $signed(_T_59729); // @[Modules.scala 160:64:@5548.4]
  assign buffer_1_263 = {{8{_T_59057[5]}},_T_59057}; // @[Modules.scala 112:22:@8.4]
  assign _T_59731 = $signed(buffer_0_263) + $signed(buffer_1_263); // @[Modules.scala 160:64:@5550.4]
  assign _T_59732 = _T_59731[13:0]; // @[Modules.scala 160:64:@5551.4]
  assign buffer_1_435 = $signed(_T_59732); // @[Modules.scala 160:64:@5552.4]
  assign buffer_1_264 = {{8{_T_59064[5]}},_T_59064}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_265 = {{9{_T_59071[4]}},_T_59071}; // @[Modules.scala 112:22:@8.4]
  assign _T_59734 = $signed(buffer_1_264) + $signed(buffer_1_265); // @[Modules.scala 160:64:@5554.4]
  assign _T_59735 = _T_59734[13:0]; // @[Modules.scala 160:64:@5555.4]
  assign buffer_1_436 = $signed(_T_59735); // @[Modules.scala 160:64:@5556.4]
  assign buffer_1_266 = {{8{_T_59078[5]}},_T_59078}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_267 = {{8{_T_59085[5]}},_T_59085}; // @[Modules.scala 112:22:@8.4]
  assign _T_59737 = $signed(buffer_1_266) + $signed(buffer_1_267); // @[Modules.scala 160:64:@5558.4]
  assign _T_59738 = _T_59737[13:0]; // @[Modules.scala 160:64:@5559.4]
  assign buffer_1_437 = $signed(_T_59738); // @[Modules.scala 160:64:@5560.4]
  assign buffer_1_268 = {{8{_T_59092[5]}},_T_59092}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_269 = {{8{_T_59099[5]}},_T_59099}; // @[Modules.scala 112:22:@8.4]
  assign _T_59740 = $signed(buffer_1_268) + $signed(buffer_1_269); // @[Modules.scala 160:64:@5562.4]
  assign _T_59741 = _T_59740[13:0]; // @[Modules.scala 160:64:@5563.4]
  assign buffer_1_438 = $signed(_T_59741); // @[Modules.scala 160:64:@5564.4]
  assign buffer_1_270 = {{9{_T_59106[4]}},_T_59106}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_271 = {{8{_T_59113[5]}},_T_59113}; // @[Modules.scala 112:22:@8.4]
  assign _T_59743 = $signed(buffer_1_270) + $signed(buffer_1_271); // @[Modules.scala 160:64:@5566.4]
  assign _T_59744 = _T_59743[13:0]; // @[Modules.scala 160:64:@5567.4]
  assign buffer_1_439 = $signed(_T_59744); // @[Modules.scala 160:64:@5568.4]
  assign buffer_1_272 = {{8{_T_59120[5]}},_T_59120}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_273 = {{8{_T_59127[5]}},_T_59127}; // @[Modules.scala 112:22:@8.4]
  assign _T_59746 = $signed(buffer_1_272) + $signed(buffer_1_273); // @[Modules.scala 160:64:@5570.4]
  assign _T_59747 = _T_59746[13:0]; // @[Modules.scala 160:64:@5571.4]
  assign buffer_1_440 = $signed(_T_59747); // @[Modules.scala 160:64:@5572.4]
  assign buffer_1_274 = {{8{_T_59134[5]}},_T_59134}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_275 = {{8{_T_59141[5]}},_T_59141}; // @[Modules.scala 112:22:@8.4]
  assign _T_59749 = $signed(buffer_1_274) + $signed(buffer_1_275); // @[Modules.scala 160:64:@5574.4]
  assign _T_59750 = _T_59749[13:0]; // @[Modules.scala 160:64:@5575.4]
  assign buffer_1_441 = $signed(_T_59750); // @[Modules.scala 160:64:@5576.4]
  assign buffer_1_276 = {{8{_T_59148[5]}},_T_59148}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_277 = {{8{_T_59155[5]}},_T_59155}; // @[Modules.scala 112:22:@8.4]
  assign _T_59752 = $signed(buffer_1_276) + $signed(buffer_1_277); // @[Modules.scala 160:64:@5578.4]
  assign _T_59753 = _T_59752[13:0]; // @[Modules.scala 160:64:@5579.4]
  assign buffer_1_442 = $signed(_T_59753); // @[Modules.scala 160:64:@5580.4]
  assign buffer_1_278 = {{8{_T_59162[5]}},_T_59162}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_279 = {{8{_T_59169[5]}},_T_59169}; // @[Modules.scala 112:22:@8.4]
  assign _T_59755 = $signed(buffer_1_278) + $signed(buffer_1_279); // @[Modules.scala 160:64:@5582.4]
  assign _T_59756 = _T_59755[13:0]; // @[Modules.scala 160:64:@5583.4]
  assign buffer_1_443 = $signed(_T_59756); // @[Modules.scala 160:64:@5584.4]
  assign buffer_1_280 = {{8{_T_59176[5]}},_T_59176}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_281 = {{8{_T_59183[5]}},_T_59183}; // @[Modules.scala 112:22:@8.4]
  assign _T_59758 = $signed(buffer_1_280) + $signed(buffer_1_281); // @[Modules.scala 160:64:@5586.4]
  assign _T_59759 = _T_59758[13:0]; // @[Modules.scala 160:64:@5587.4]
  assign buffer_1_444 = $signed(_T_59759); // @[Modules.scala 160:64:@5588.4]
  assign buffer_1_282 = {{8{_T_59190[5]}},_T_59190}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_283 = {{9{_T_59197[4]}},_T_59197}; // @[Modules.scala 112:22:@8.4]
  assign _T_59761 = $signed(buffer_1_282) + $signed(buffer_1_283); // @[Modules.scala 160:64:@5590.4]
  assign _T_59762 = _T_59761[13:0]; // @[Modules.scala 160:64:@5591.4]
  assign buffer_1_445 = $signed(_T_59762); // @[Modules.scala 160:64:@5592.4]
  assign buffer_1_284 = {{8{_T_59204[5]}},_T_59204}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_285 = {{8{_T_59211[5]}},_T_59211}; // @[Modules.scala 112:22:@8.4]
  assign _T_59764 = $signed(buffer_1_284) + $signed(buffer_1_285); // @[Modules.scala 160:64:@5594.4]
  assign _T_59765 = _T_59764[13:0]; // @[Modules.scala 160:64:@5595.4]
  assign buffer_1_446 = $signed(_T_59765); // @[Modules.scala 160:64:@5596.4]
  assign buffer_1_288 = {{8{_T_59232[5]}},_T_59232}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_289 = {{8{_T_59239[5]}},_T_59239}; // @[Modules.scala 112:22:@8.4]
  assign _T_59770 = $signed(buffer_1_288) + $signed(buffer_1_289); // @[Modules.scala 160:64:@5602.4]
  assign _T_59771 = _T_59770[13:0]; // @[Modules.scala 160:64:@5603.4]
  assign buffer_1_448 = $signed(_T_59771); // @[Modules.scala 160:64:@5604.4]
  assign buffer_1_290 = {{8{_T_59246[5]}},_T_59246}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_291 = {{8{_T_59253[5]}},_T_59253}; // @[Modules.scala 112:22:@8.4]
  assign _T_59773 = $signed(buffer_1_290) + $signed(buffer_1_291); // @[Modules.scala 160:64:@5606.4]
  assign _T_59774 = _T_59773[13:0]; // @[Modules.scala 160:64:@5607.4]
  assign buffer_1_449 = $signed(_T_59774); // @[Modules.scala 160:64:@5608.4]
  assign buffer_1_292 = {{8{_T_59260[5]}},_T_59260}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_293 = {{8{_T_59267[5]}},_T_59267}; // @[Modules.scala 112:22:@8.4]
  assign _T_59776 = $signed(buffer_1_292) + $signed(buffer_1_293); // @[Modules.scala 160:64:@5610.4]
  assign _T_59777 = _T_59776[13:0]; // @[Modules.scala 160:64:@5611.4]
  assign buffer_1_450 = $signed(_T_59777); // @[Modules.scala 160:64:@5612.4]
  assign buffer_1_294 = {{8{_T_59274[5]}},_T_59274}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_295 = {{8{_T_59281[5]}},_T_59281}; // @[Modules.scala 112:22:@8.4]
  assign _T_59779 = $signed(buffer_1_294) + $signed(buffer_1_295); // @[Modules.scala 160:64:@5614.4]
  assign _T_59780 = _T_59779[13:0]; // @[Modules.scala 160:64:@5615.4]
  assign buffer_1_451 = $signed(_T_59780); // @[Modules.scala 160:64:@5616.4]
  assign buffer_1_297 = {{9{_T_59295[4]}},_T_59295}; // @[Modules.scala 112:22:@8.4]
  assign _T_59782 = $signed(buffer_0_295) + $signed(buffer_1_297); // @[Modules.scala 160:64:@5618.4]
  assign _T_59783 = _T_59782[13:0]; // @[Modules.scala 160:64:@5619.4]
  assign buffer_1_452 = $signed(_T_59783); // @[Modules.scala 160:64:@5620.4]
  assign buffer_1_298 = {{8{_T_59302[5]}},_T_59302}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_299 = {{8{_T_59309[5]}},_T_59309}; // @[Modules.scala 112:22:@8.4]
  assign _T_59785 = $signed(buffer_1_298) + $signed(buffer_1_299); // @[Modules.scala 160:64:@5622.4]
  assign _T_59786 = _T_59785[13:0]; // @[Modules.scala 160:64:@5623.4]
  assign buffer_1_453 = $signed(_T_59786); // @[Modules.scala 160:64:@5624.4]
  assign buffer_1_300 = {{8{_T_59316[5]}},_T_59316}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_301 = {{8{_T_59323[5]}},_T_59323}; // @[Modules.scala 112:22:@8.4]
  assign _T_59788 = $signed(buffer_1_300) + $signed(buffer_1_301); // @[Modules.scala 160:64:@5626.4]
  assign _T_59789 = _T_59788[13:0]; // @[Modules.scala 160:64:@5627.4]
  assign buffer_1_454 = $signed(_T_59789); // @[Modules.scala 160:64:@5628.4]
  assign buffer_1_302 = {{8{_T_59330[5]}},_T_59330}; // @[Modules.scala 112:22:@8.4]
  assign buffer_1_303 = {{9{_T_59337[4]}},_T_59337}; // @[Modules.scala 112:22:@8.4]
  assign _T_59791 = $signed(buffer_1_302) + $signed(buffer_1_303); // @[Modules.scala 160:64:@5630.4]
  assign _T_59792 = _T_59791[13:0]; // @[Modules.scala 160:64:@5631.4]
  assign buffer_1_455 = $signed(_T_59792); // @[Modules.scala 160:64:@5632.4]
  assign _T_59794 = $signed(buffer_0_302) + $signed(buffer_1_305); // @[Modules.scala 160:64:@5634.4]
  assign _T_59795 = _T_59794[13:0]; // @[Modules.scala 160:64:@5635.4]
  assign buffer_1_456 = $signed(_T_59795); // @[Modules.scala 160:64:@5636.4]
  assign _T_59797 = $signed(buffer_1_306) + $signed(buffer_1_307); // @[Modules.scala 160:64:@5638.4]
  assign _T_59798 = _T_59797[13:0]; // @[Modules.scala 160:64:@5639.4]
  assign buffer_1_457 = $signed(_T_59798); // @[Modules.scala 160:64:@5640.4]
  assign _T_59800 = $signed(buffer_1_308) + $signed(buffer_1_309); // @[Modules.scala 160:64:@5642.4]
  assign _T_59801 = _T_59800[13:0]; // @[Modules.scala 160:64:@5643.4]
  assign buffer_1_458 = $signed(_T_59801); // @[Modules.scala 160:64:@5644.4]
  assign _T_59803 = $signed(buffer_1_310) + $signed(buffer_1_311); // @[Modules.scala 160:64:@5646.4]
  assign _T_59804 = _T_59803[13:0]; // @[Modules.scala 160:64:@5647.4]
  assign buffer_1_459 = $signed(_T_59804); // @[Modules.scala 160:64:@5648.4]
  assign _T_59806 = $signed(buffer_1_312) + $signed(buffer_1_313); // @[Modules.scala 160:64:@5650.4]
  assign _T_59807 = _T_59806[13:0]; // @[Modules.scala 160:64:@5651.4]
  assign buffer_1_460 = $signed(_T_59807); // @[Modules.scala 160:64:@5652.4]
  assign _T_59809 = $signed(buffer_1_314) + $signed(buffer_1_315); // @[Modules.scala 160:64:@5654.4]
  assign _T_59810 = _T_59809[13:0]; // @[Modules.scala 160:64:@5655.4]
  assign buffer_1_461 = $signed(_T_59810); // @[Modules.scala 160:64:@5656.4]
  assign _T_59812 = $signed(buffer_1_316) + $signed(buffer_1_317); // @[Modules.scala 160:64:@5658.4]
  assign _T_59813 = _T_59812[13:0]; // @[Modules.scala 160:64:@5659.4]
  assign buffer_1_462 = $signed(_T_59813); // @[Modules.scala 160:64:@5660.4]
  assign _T_59815 = $signed(buffer_1_318) + $signed(buffer_1_319); // @[Modules.scala 160:64:@5662.4]
  assign _T_59816 = _T_59815[13:0]; // @[Modules.scala 160:64:@5663.4]
  assign buffer_1_463 = $signed(_T_59816); // @[Modules.scala 160:64:@5664.4]
  assign _T_59818 = $signed(buffer_1_320) + $signed(buffer_1_321); // @[Modules.scala 160:64:@5666.4]
  assign _T_59819 = _T_59818[13:0]; // @[Modules.scala 160:64:@5667.4]
  assign buffer_1_464 = $signed(_T_59819); // @[Modules.scala 160:64:@5668.4]
  assign _T_59821 = $signed(buffer_1_322) + $signed(buffer_1_323); // @[Modules.scala 160:64:@5670.4]
  assign _T_59822 = _T_59821[13:0]; // @[Modules.scala 160:64:@5671.4]
  assign buffer_1_465 = $signed(_T_59822); // @[Modules.scala 160:64:@5672.4]
  assign _T_59824 = $signed(buffer_1_324) + $signed(buffer_1_325); // @[Modules.scala 160:64:@5674.4]
  assign _T_59825 = _T_59824[13:0]; // @[Modules.scala 160:64:@5675.4]
  assign buffer_1_466 = $signed(_T_59825); // @[Modules.scala 160:64:@5676.4]
  assign _T_59827 = $signed(buffer_1_326) + $signed(buffer_1_327); // @[Modules.scala 160:64:@5678.4]
  assign _T_59828 = _T_59827[13:0]; // @[Modules.scala 160:64:@5679.4]
  assign buffer_1_467 = $signed(_T_59828); // @[Modules.scala 160:64:@5680.4]
  assign _T_59830 = $signed(buffer_1_328) + $signed(buffer_1_329); // @[Modules.scala 160:64:@5682.4]
  assign _T_59831 = _T_59830[13:0]; // @[Modules.scala 160:64:@5683.4]
  assign buffer_1_468 = $signed(_T_59831); // @[Modules.scala 160:64:@5684.4]
  assign _T_59833 = $signed(buffer_1_330) + $signed(buffer_1_331); // @[Modules.scala 160:64:@5686.4]
  assign _T_59834 = _T_59833[13:0]; // @[Modules.scala 160:64:@5687.4]
  assign buffer_1_469 = $signed(_T_59834); // @[Modules.scala 160:64:@5688.4]
  assign _T_59836 = $signed(buffer_1_332) + $signed(buffer_1_333); // @[Modules.scala 160:64:@5690.4]
  assign _T_59837 = _T_59836[13:0]; // @[Modules.scala 160:64:@5691.4]
  assign buffer_1_470 = $signed(_T_59837); // @[Modules.scala 160:64:@5692.4]
  assign _T_59839 = $signed(buffer_1_334) + $signed(buffer_1_335); // @[Modules.scala 160:64:@5694.4]
  assign _T_59840 = _T_59839[13:0]; // @[Modules.scala 160:64:@5695.4]
  assign buffer_1_471 = $signed(_T_59840); // @[Modules.scala 160:64:@5696.4]
  assign _T_59842 = $signed(buffer_1_336) + $signed(buffer_1_337); // @[Modules.scala 160:64:@5698.4]
  assign _T_59843 = _T_59842[13:0]; // @[Modules.scala 160:64:@5699.4]
  assign buffer_1_472 = $signed(_T_59843); // @[Modules.scala 160:64:@5700.4]
  assign _T_59845 = $signed(buffer_1_338) + $signed(buffer_1_339); // @[Modules.scala 160:64:@5702.4]
  assign _T_59846 = _T_59845[13:0]; // @[Modules.scala 160:64:@5703.4]
  assign buffer_1_473 = $signed(_T_59846); // @[Modules.scala 160:64:@5704.4]
  assign _T_59848 = $signed(buffer_1_340) + $signed(buffer_1_341); // @[Modules.scala 160:64:@5706.4]
  assign _T_59849 = _T_59848[13:0]; // @[Modules.scala 160:64:@5707.4]
  assign buffer_1_474 = $signed(_T_59849); // @[Modules.scala 160:64:@5708.4]
  assign _T_59851 = $signed(buffer_1_342) + $signed(buffer_1_343); // @[Modules.scala 160:64:@5710.4]
  assign _T_59852 = _T_59851[13:0]; // @[Modules.scala 160:64:@5711.4]
  assign buffer_1_475 = $signed(_T_59852); // @[Modules.scala 160:64:@5712.4]
  assign _T_59854 = $signed(buffer_1_344) + $signed(buffer_1_345); // @[Modules.scala 160:64:@5714.4]
  assign _T_59855 = _T_59854[13:0]; // @[Modules.scala 160:64:@5715.4]
  assign buffer_1_476 = $signed(_T_59855); // @[Modules.scala 160:64:@5716.4]
  assign _T_59857 = $signed(buffer_1_346) + $signed(buffer_1_347); // @[Modules.scala 160:64:@5718.4]
  assign _T_59858 = _T_59857[13:0]; // @[Modules.scala 160:64:@5719.4]
  assign buffer_1_477 = $signed(_T_59858); // @[Modules.scala 160:64:@5720.4]
  assign _T_59860 = $signed(buffer_0_344) + $signed(buffer_1_349); // @[Modules.scala 160:64:@5722.4]
  assign _T_59861 = _T_59860[13:0]; // @[Modules.scala 160:64:@5723.4]
  assign buffer_1_478 = $signed(_T_59861); // @[Modules.scala 160:64:@5724.4]
  assign _T_59863 = $signed(buffer_1_350) + $signed(buffer_1_351); // @[Modules.scala 160:64:@5726.4]
  assign _T_59864 = _T_59863[13:0]; // @[Modules.scala 160:64:@5727.4]
  assign buffer_1_479 = $signed(_T_59864); // @[Modules.scala 160:64:@5728.4]
  assign _T_59866 = $signed(buffer_1_352) + $signed(buffer_1_353); // @[Modules.scala 160:64:@5730.4]
  assign _T_59867 = _T_59866[13:0]; // @[Modules.scala 160:64:@5731.4]
  assign buffer_1_480 = $signed(_T_59867); // @[Modules.scala 160:64:@5732.4]
  assign _T_59869 = $signed(buffer_1_354) + $signed(buffer_1_355); // @[Modules.scala 160:64:@5734.4]
  assign _T_59870 = _T_59869[13:0]; // @[Modules.scala 160:64:@5735.4]
  assign buffer_1_481 = $signed(_T_59870); // @[Modules.scala 160:64:@5736.4]
  assign _T_59872 = $signed(buffer_1_356) + $signed(buffer_1_357); // @[Modules.scala 160:64:@5738.4]
  assign _T_59873 = _T_59872[13:0]; // @[Modules.scala 160:64:@5739.4]
  assign buffer_1_482 = $signed(_T_59873); // @[Modules.scala 160:64:@5740.4]
  assign _T_59875 = $signed(buffer_1_358) + $signed(buffer_1_359); // @[Modules.scala 160:64:@5742.4]
  assign _T_59876 = _T_59875[13:0]; // @[Modules.scala 160:64:@5743.4]
  assign buffer_1_483 = $signed(_T_59876); // @[Modules.scala 160:64:@5744.4]
  assign _T_59878 = $signed(buffer_1_360) + $signed(buffer_1_361); // @[Modules.scala 160:64:@5746.4]
  assign _T_59879 = _T_59878[13:0]; // @[Modules.scala 160:64:@5747.4]
  assign buffer_1_484 = $signed(_T_59879); // @[Modules.scala 160:64:@5748.4]
  assign _T_59881 = $signed(buffer_1_362) + $signed(buffer_1_363); // @[Modules.scala 160:64:@5750.4]
  assign _T_59882 = _T_59881[13:0]; // @[Modules.scala 160:64:@5751.4]
  assign buffer_1_485 = $signed(_T_59882); // @[Modules.scala 160:64:@5752.4]
  assign _T_59884 = $signed(buffer_1_364) + $signed(buffer_1_365); // @[Modules.scala 160:64:@5754.4]
  assign _T_59885 = _T_59884[13:0]; // @[Modules.scala 160:64:@5755.4]
  assign buffer_1_486 = $signed(_T_59885); // @[Modules.scala 160:64:@5756.4]
  assign _T_59887 = $signed(buffer_1_366) + $signed(buffer_1_367); // @[Modules.scala 160:64:@5758.4]
  assign _T_59888 = _T_59887[13:0]; // @[Modules.scala 160:64:@5759.4]
  assign buffer_1_487 = $signed(_T_59888); // @[Modules.scala 160:64:@5760.4]
  assign _T_59890 = $signed(buffer_1_368) + $signed(buffer_1_369); // @[Modules.scala 160:64:@5762.4]
  assign _T_59891 = _T_59890[13:0]; // @[Modules.scala 160:64:@5763.4]
  assign buffer_1_488 = $signed(_T_59891); // @[Modules.scala 160:64:@5764.4]
  assign _T_59893 = $signed(buffer_1_370) + $signed(buffer_1_371); // @[Modules.scala 160:64:@5766.4]
  assign _T_59894 = _T_59893[13:0]; // @[Modules.scala 160:64:@5767.4]
  assign buffer_1_489 = $signed(_T_59894); // @[Modules.scala 160:64:@5768.4]
  assign _T_59896 = $signed(buffer_1_372) + $signed(buffer_1_373); // @[Modules.scala 160:64:@5770.4]
  assign _T_59897 = _T_59896[13:0]; // @[Modules.scala 160:64:@5771.4]
  assign buffer_1_490 = $signed(_T_59897); // @[Modules.scala 160:64:@5772.4]
  assign _T_59899 = $signed(buffer_1_374) + $signed(buffer_1_375); // @[Modules.scala 160:64:@5774.4]
  assign _T_59900 = _T_59899[13:0]; // @[Modules.scala 160:64:@5775.4]
  assign buffer_1_491 = $signed(_T_59900); // @[Modules.scala 160:64:@5776.4]
  assign _T_59902 = $signed(buffer_1_376) + $signed(buffer_1_377); // @[Modules.scala 160:64:@5778.4]
  assign _T_59903 = _T_59902[13:0]; // @[Modules.scala 160:64:@5779.4]
  assign buffer_1_492 = $signed(_T_59903); // @[Modules.scala 160:64:@5780.4]
  assign _T_59905 = $signed(buffer_1_378) + $signed(buffer_1_379); // @[Modules.scala 160:64:@5782.4]
  assign _T_59906 = _T_59905[13:0]; // @[Modules.scala 160:64:@5783.4]
  assign buffer_1_493 = $signed(_T_59906); // @[Modules.scala 160:64:@5784.4]
  assign _T_59908 = $signed(buffer_1_380) + $signed(buffer_1_381); // @[Modules.scala 160:64:@5786.4]
  assign _T_59909 = _T_59908[13:0]; // @[Modules.scala 160:64:@5787.4]
  assign buffer_1_494 = $signed(_T_59909); // @[Modules.scala 160:64:@5788.4]
  assign _T_59911 = $signed(buffer_1_382) + $signed(buffer_1_383); // @[Modules.scala 160:64:@5790.4]
  assign _T_59912 = _T_59911[13:0]; // @[Modules.scala 160:64:@5791.4]
  assign buffer_1_495 = $signed(_T_59912); // @[Modules.scala 160:64:@5792.4]
  assign _T_59914 = $signed(buffer_1_384) + $signed(buffer_1_385); // @[Modules.scala 160:64:@5794.4]
  assign _T_59915 = _T_59914[13:0]; // @[Modules.scala 160:64:@5795.4]
  assign buffer_1_496 = $signed(_T_59915); // @[Modules.scala 160:64:@5796.4]
  assign _T_59917 = $signed(buffer_1_386) + $signed(buffer_1_387); // @[Modules.scala 160:64:@5798.4]
  assign _T_59918 = _T_59917[13:0]; // @[Modules.scala 160:64:@5799.4]
  assign buffer_1_497 = $signed(_T_59918); // @[Modules.scala 160:64:@5800.4]
  assign _T_59920 = $signed(buffer_1_388) + $signed(buffer_1_389); // @[Modules.scala 160:64:@5802.4]
  assign _T_59921 = _T_59920[13:0]; // @[Modules.scala 160:64:@5803.4]
  assign buffer_1_498 = $signed(_T_59921); // @[Modules.scala 160:64:@5804.4]
  assign _T_59923 = $signed(buffer_1_390) + $signed(buffer_1_391); // @[Modules.scala 160:64:@5806.4]
  assign _T_59924 = _T_59923[13:0]; // @[Modules.scala 160:64:@5807.4]
  assign buffer_1_499 = $signed(_T_59924); // @[Modules.scala 160:64:@5808.4]
  assign _T_59926 = $signed(buffer_1_392) + $signed(buffer_1_393); // @[Modules.scala 160:64:@5810.4]
  assign _T_59927 = _T_59926[13:0]; // @[Modules.scala 160:64:@5811.4]
  assign buffer_1_500 = $signed(_T_59927); // @[Modules.scala 160:64:@5812.4]
  assign _T_59929 = $signed(buffer_1_394) + $signed(buffer_1_395); // @[Modules.scala 160:64:@5814.4]
  assign _T_59930 = _T_59929[13:0]; // @[Modules.scala 160:64:@5815.4]
  assign buffer_1_501 = $signed(_T_59930); // @[Modules.scala 160:64:@5816.4]
  assign _T_59932 = $signed(buffer_1_396) + $signed(buffer_1_397); // @[Modules.scala 160:64:@5818.4]
  assign _T_59933 = _T_59932[13:0]; // @[Modules.scala 160:64:@5819.4]
  assign buffer_1_502 = $signed(_T_59933); // @[Modules.scala 160:64:@5820.4]
  assign _T_59935 = $signed(buffer_1_398) + $signed(buffer_1_399); // @[Modules.scala 160:64:@5822.4]
  assign _T_59936 = _T_59935[13:0]; // @[Modules.scala 160:64:@5823.4]
  assign buffer_1_503 = $signed(_T_59936); // @[Modules.scala 160:64:@5824.4]
  assign _T_59938 = $signed(buffer_1_400) + $signed(buffer_1_401); // @[Modules.scala 160:64:@5826.4]
  assign _T_59939 = _T_59938[13:0]; // @[Modules.scala 160:64:@5827.4]
  assign buffer_1_504 = $signed(_T_59939); // @[Modules.scala 160:64:@5828.4]
  assign _T_59941 = $signed(buffer_1_402) + $signed(buffer_1_403); // @[Modules.scala 160:64:@5830.4]
  assign _T_59942 = _T_59941[13:0]; // @[Modules.scala 160:64:@5831.4]
  assign buffer_1_505 = $signed(_T_59942); // @[Modules.scala 160:64:@5832.4]
  assign _T_59944 = $signed(buffer_1_404) + $signed(buffer_1_405); // @[Modules.scala 160:64:@5834.4]
  assign _T_59945 = _T_59944[13:0]; // @[Modules.scala 160:64:@5835.4]
  assign buffer_1_506 = $signed(_T_59945); // @[Modules.scala 160:64:@5836.4]
  assign _T_59947 = $signed(buffer_1_406) + $signed(buffer_1_407); // @[Modules.scala 160:64:@5838.4]
  assign _T_59948 = _T_59947[13:0]; // @[Modules.scala 160:64:@5839.4]
  assign buffer_1_507 = $signed(_T_59948); // @[Modules.scala 160:64:@5840.4]
  assign _T_59950 = $signed(buffer_1_408) + $signed(buffer_1_409); // @[Modules.scala 160:64:@5842.4]
  assign _T_59951 = _T_59950[13:0]; // @[Modules.scala 160:64:@5843.4]
  assign buffer_1_508 = $signed(_T_59951); // @[Modules.scala 160:64:@5844.4]
  assign _T_59953 = $signed(buffer_1_410) + $signed(buffer_1_411); // @[Modules.scala 160:64:@5846.4]
  assign _T_59954 = _T_59953[13:0]; // @[Modules.scala 160:64:@5847.4]
  assign buffer_1_509 = $signed(_T_59954); // @[Modules.scala 160:64:@5848.4]
  assign _T_59956 = $signed(buffer_1_412) + $signed(buffer_1_413); // @[Modules.scala 160:64:@5850.4]
  assign _T_59957 = _T_59956[13:0]; // @[Modules.scala 160:64:@5851.4]
  assign buffer_1_510 = $signed(_T_59957); // @[Modules.scala 160:64:@5852.4]
  assign _T_59959 = $signed(buffer_1_414) + $signed(buffer_1_415); // @[Modules.scala 160:64:@5854.4]
  assign _T_59960 = _T_59959[13:0]; // @[Modules.scala 160:64:@5855.4]
  assign buffer_1_511 = $signed(_T_59960); // @[Modules.scala 160:64:@5856.4]
  assign _T_59962 = $signed(buffer_1_416) + $signed(buffer_1_417); // @[Modules.scala 160:64:@5858.4]
  assign _T_59963 = _T_59962[13:0]; // @[Modules.scala 160:64:@5859.4]
  assign buffer_1_512 = $signed(_T_59963); // @[Modules.scala 160:64:@5860.4]
  assign _T_59965 = $signed(buffer_1_418) + $signed(buffer_0_416); // @[Modules.scala 160:64:@5862.4]
  assign _T_59966 = _T_59965[13:0]; // @[Modules.scala 160:64:@5863.4]
  assign buffer_1_513 = $signed(_T_59966); // @[Modules.scala 160:64:@5864.4]
  assign _T_59968 = $signed(buffer_1_420) + $signed(buffer_1_421); // @[Modules.scala 160:64:@5866.4]
  assign _T_59969 = _T_59968[13:0]; // @[Modules.scala 160:64:@5867.4]
  assign buffer_1_514 = $signed(_T_59969); // @[Modules.scala 160:64:@5868.4]
  assign _T_59971 = $signed(buffer_1_422) + $signed(buffer_1_423); // @[Modules.scala 160:64:@5870.4]
  assign _T_59972 = _T_59971[13:0]; // @[Modules.scala 160:64:@5871.4]
  assign buffer_1_515 = $signed(_T_59972); // @[Modules.scala 160:64:@5872.4]
  assign _T_59974 = $signed(buffer_1_424) + $signed(buffer_1_425); // @[Modules.scala 160:64:@5874.4]
  assign _T_59975 = _T_59974[13:0]; // @[Modules.scala 160:64:@5875.4]
  assign buffer_1_516 = $signed(_T_59975); // @[Modules.scala 160:64:@5876.4]
  assign _T_59977 = $signed(buffer_1_426) + $signed(buffer_1_427); // @[Modules.scala 160:64:@5878.4]
  assign _T_59978 = _T_59977[13:0]; // @[Modules.scala 160:64:@5879.4]
  assign buffer_1_517 = $signed(_T_59978); // @[Modules.scala 160:64:@5880.4]
  assign _T_59980 = $signed(buffer_1_428) + $signed(buffer_1_429); // @[Modules.scala 160:64:@5882.4]
  assign _T_59981 = _T_59980[13:0]; // @[Modules.scala 160:64:@5883.4]
  assign buffer_1_518 = $signed(_T_59981); // @[Modules.scala 160:64:@5884.4]
  assign _T_59983 = $signed(buffer_1_430) + $signed(buffer_1_431); // @[Modules.scala 160:64:@5886.4]
  assign _T_59984 = _T_59983[13:0]; // @[Modules.scala 160:64:@5887.4]
  assign buffer_1_519 = $signed(_T_59984); // @[Modules.scala 160:64:@5888.4]
  assign _T_59986 = $signed(buffer_1_432) + $signed(buffer_1_433); // @[Modules.scala 160:64:@5890.4]
  assign _T_59987 = _T_59986[13:0]; // @[Modules.scala 160:64:@5891.4]
  assign buffer_1_520 = $signed(_T_59987); // @[Modules.scala 160:64:@5892.4]
  assign _T_59989 = $signed(buffer_1_434) + $signed(buffer_1_435); // @[Modules.scala 160:64:@5894.4]
  assign _T_59990 = _T_59989[13:0]; // @[Modules.scala 160:64:@5895.4]
  assign buffer_1_521 = $signed(_T_59990); // @[Modules.scala 160:64:@5896.4]
  assign _T_59992 = $signed(buffer_1_436) + $signed(buffer_1_437); // @[Modules.scala 160:64:@5898.4]
  assign _T_59993 = _T_59992[13:0]; // @[Modules.scala 160:64:@5899.4]
  assign buffer_1_522 = $signed(_T_59993); // @[Modules.scala 160:64:@5900.4]
  assign _T_59995 = $signed(buffer_1_438) + $signed(buffer_1_439); // @[Modules.scala 160:64:@5902.4]
  assign _T_59996 = _T_59995[13:0]; // @[Modules.scala 160:64:@5903.4]
  assign buffer_1_523 = $signed(_T_59996); // @[Modules.scala 160:64:@5904.4]
  assign _T_59998 = $signed(buffer_1_440) + $signed(buffer_1_441); // @[Modules.scala 160:64:@5906.4]
  assign _T_59999 = _T_59998[13:0]; // @[Modules.scala 160:64:@5907.4]
  assign buffer_1_524 = $signed(_T_59999); // @[Modules.scala 160:64:@5908.4]
  assign _T_60001 = $signed(buffer_1_442) + $signed(buffer_1_443); // @[Modules.scala 160:64:@5910.4]
  assign _T_60002 = _T_60001[13:0]; // @[Modules.scala 160:64:@5911.4]
  assign buffer_1_525 = $signed(_T_60002); // @[Modules.scala 160:64:@5912.4]
  assign _T_60004 = $signed(buffer_1_444) + $signed(buffer_1_445); // @[Modules.scala 160:64:@5914.4]
  assign _T_60005 = _T_60004[13:0]; // @[Modules.scala 160:64:@5915.4]
  assign buffer_1_526 = $signed(_T_60005); // @[Modules.scala 160:64:@5916.4]
  assign _T_60007 = $signed(buffer_1_446) + $signed(buffer_0_445); // @[Modules.scala 160:64:@5918.4]
  assign _T_60008 = _T_60007[13:0]; // @[Modules.scala 160:64:@5919.4]
  assign buffer_1_527 = $signed(_T_60008); // @[Modules.scala 160:64:@5920.4]
  assign _T_60010 = $signed(buffer_1_448) + $signed(buffer_1_449); // @[Modules.scala 160:64:@5922.4]
  assign _T_60011 = _T_60010[13:0]; // @[Modules.scala 160:64:@5923.4]
  assign buffer_1_528 = $signed(_T_60011); // @[Modules.scala 160:64:@5924.4]
  assign _T_60013 = $signed(buffer_1_450) + $signed(buffer_1_451); // @[Modules.scala 160:64:@5926.4]
  assign _T_60014 = _T_60013[13:0]; // @[Modules.scala 160:64:@5927.4]
  assign buffer_1_529 = $signed(_T_60014); // @[Modules.scala 160:64:@5928.4]
  assign _T_60016 = $signed(buffer_1_452) + $signed(buffer_1_453); // @[Modules.scala 160:64:@5930.4]
  assign _T_60017 = _T_60016[13:0]; // @[Modules.scala 160:64:@5931.4]
  assign buffer_1_530 = $signed(_T_60017); // @[Modules.scala 160:64:@5932.4]
  assign _T_60019 = $signed(buffer_1_454) + $signed(buffer_1_455); // @[Modules.scala 160:64:@5934.4]
  assign _T_60020 = _T_60019[13:0]; // @[Modules.scala 160:64:@5935.4]
  assign buffer_1_531 = $signed(_T_60020); // @[Modules.scala 160:64:@5936.4]
  assign _T_60022 = $signed(buffer_1_456) + $signed(buffer_1_457); // @[Modules.scala 160:64:@5938.4]
  assign _T_60023 = _T_60022[13:0]; // @[Modules.scala 160:64:@5939.4]
  assign buffer_1_532 = $signed(_T_60023); // @[Modules.scala 160:64:@5940.4]
  assign _T_60025 = $signed(buffer_1_458) + $signed(buffer_1_459); // @[Modules.scala 160:64:@5942.4]
  assign _T_60026 = _T_60025[13:0]; // @[Modules.scala 160:64:@5943.4]
  assign buffer_1_533 = $signed(_T_60026); // @[Modules.scala 160:64:@5944.4]
  assign _T_60028 = $signed(buffer_1_460) + $signed(buffer_1_461); // @[Modules.scala 160:64:@5946.4]
  assign _T_60029 = _T_60028[13:0]; // @[Modules.scala 160:64:@5947.4]
  assign buffer_1_534 = $signed(_T_60029); // @[Modules.scala 160:64:@5948.4]
  assign _T_60031 = $signed(buffer_1_462) + $signed(buffer_1_463); // @[Modules.scala 160:64:@5950.4]
  assign _T_60032 = _T_60031[13:0]; // @[Modules.scala 160:64:@5951.4]
  assign buffer_1_535 = $signed(_T_60032); // @[Modules.scala 160:64:@5952.4]
  assign _T_60034 = $signed(buffer_1_464) + $signed(buffer_1_465); // @[Modules.scala 160:64:@5954.4]
  assign _T_60035 = _T_60034[13:0]; // @[Modules.scala 160:64:@5955.4]
  assign buffer_1_536 = $signed(_T_60035); // @[Modules.scala 160:64:@5956.4]
  assign _T_60037 = $signed(buffer_1_466) + $signed(buffer_1_467); // @[Modules.scala 160:64:@5958.4]
  assign _T_60038 = _T_60037[13:0]; // @[Modules.scala 160:64:@5959.4]
  assign buffer_1_537 = $signed(_T_60038); // @[Modules.scala 160:64:@5960.4]
  assign _T_60040 = $signed(buffer_1_468) + $signed(buffer_1_469); // @[Modules.scala 160:64:@5962.4]
  assign _T_60041 = _T_60040[13:0]; // @[Modules.scala 160:64:@5963.4]
  assign buffer_1_538 = $signed(_T_60041); // @[Modules.scala 160:64:@5964.4]
  assign _T_60043 = $signed(buffer_1_470) + $signed(buffer_1_471); // @[Modules.scala 160:64:@5966.4]
  assign _T_60044 = _T_60043[13:0]; // @[Modules.scala 160:64:@5967.4]
  assign buffer_1_539 = $signed(_T_60044); // @[Modules.scala 160:64:@5968.4]
  assign _T_60046 = $signed(buffer_1_472) + $signed(buffer_1_473); // @[Modules.scala 160:64:@5970.4]
  assign _T_60047 = _T_60046[13:0]; // @[Modules.scala 160:64:@5971.4]
  assign buffer_1_540 = $signed(_T_60047); // @[Modules.scala 160:64:@5972.4]
  assign _T_60049 = $signed(buffer_1_474) + $signed(buffer_1_475); // @[Modules.scala 160:64:@5974.4]
  assign _T_60050 = _T_60049[13:0]; // @[Modules.scala 160:64:@5975.4]
  assign buffer_1_541 = $signed(_T_60050); // @[Modules.scala 160:64:@5976.4]
  assign _T_60052 = $signed(buffer_1_476) + $signed(buffer_1_477); // @[Modules.scala 160:64:@5978.4]
  assign _T_60053 = _T_60052[13:0]; // @[Modules.scala 160:64:@5979.4]
  assign buffer_1_542 = $signed(_T_60053); // @[Modules.scala 160:64:@5980.4]
  assign _T_60055 = $signed(buffer_1_478) + $signed(buffer_1_479); // @[Modules.scala 160:64:@5982.4]
  assign _T_60056 = _T_60055[13:0]; // @[Modules.scala 160:64:@5983.4]
  assign buffer_1_543 = $signed(_T_60056); // @[Modules.scala 160:64:@5984.4]
  assign _T_60058 = $signed(buffer_1_480) + $signed(buffer_1_481); // @[Modules.scala 160:64:@5986.4]
  assign _T_60059 = _T_60058[13:0]; // @[Modules.scala 160:64:@5987.4]
  assign buffer_1_544 = $signed(_T_60059); // @[Modules.scala 160:64:@5988.4]
  assign _T_60061 = $signed(buffer_1_482) + $signed(buffer_1_483); // @[Modules.scala 160:64:@5990.4]
  assign _T_60062 = _T_60061[13:0]; // @[Modules.scala 160:64:@5991.4]
  assign buffer_1_545 = $signed(_T_60062); // @[Modules.scala 160:64:@5992.4]
  assign _T_60064 = $signed(buffer_1_484) + $signed(buffer_1_485); // @[Modules.scala 160:64:@5994.4]
  assign _T_60065 = _T_60064[13:0]; // @[Modules.scala 160:64:@5995.4]
  assign buffer_1_546 = $signed(_T_60065); // @[Modules.scala 160:64:@5996.4]
  assign _T_60067 = $signed(buffer_1_486) + $signed(buffer_1_487); // @[Modules.scala 160:64:@5998.4]
  assign _T_60068 = _T_60067[13:0]; // @[Modules.scala 160:64:@5999.4]
  assign buffer_1_547 = $signed(_T_60068); // @[Modules.scala 160:64:@6000.4]
  assign _T_60070 = $signed(buffer_1_488) + $signed(buffer_1_489); // @[Modules.scala 160:64:@6002.4]
  assign _T_60071 = _T_60070[13:0]; // @[Modules.scala 160:64:@6003.4]
  assign buffer_1_548 = $signed(_T_60071); // @[Modules.scala 160:64:@6004.4]
  assign _T_60073 = $signed(buffer_1_490) + $signed(buffer_1_491); // @[Modules.scala 160:64:@6006.4]
  assign _T_60074 = _T_60073[13:0]; // @[Modules.scala 160:64:@6007.4]
  assign buffer_1_549 = $signed(_T_60074); // @[Modules.scala 160:64:@6008.4]
  assign _T_60076 = $signed(buffer_1_492) + $signed(buffer_1_493); // @[Modules.scala 160:64:@6010.4]
  assign _T_60077 = _T_60076[13:0]; // @[Modules.scala 160:64:@6011.4]
  assign buffer_1_550 = $signed(_T_60077); // @[Modules.scala 160:64:@6012.4]
  assign _T_60079 = $signed(buffer_1_494) + $signed(buffer_1_495); // @[Modules.scala 160:64:@6014.4]
  assign _T_60080 = _T_60079[13:0]; // @[Modules.scala 160:64:@6015.4]
  assign buffer_1_551 = $signed(_T_60080); // @[Modules.scala 160:64:@6016.4]
  assign _T_60082 = $signed(buffer_1_496) + $signed(buffer_1_497); // @[Modules.scala 160:64:@6018.4]
  assign _T_60083 = _T_60082[13:0]; // @[Modules.scala 160:64:@6019.4]
  assign buffer_1_552 = $signed(_T_60083); // @[Modules.scala 160:64:@6020.4]
  assign _T_60085 = $signed(buffer_1_498) + $signed(buffer_1_499); // @[Modules.scala 160:64:@6022.4]
  assign _T_60086 = _T_60085[13:0]; // @[Modules.scala 160:64:@6023.4]
  assign buffer_1_553 = $signed(_T_60086); // @[Modules.scala 160:64:@6024.4]
  assign _T_60088 = $signed(buffer_1_500) + $signed(buffer_1_501); // @[Modules.scala 160:64:@6026.4]
  assign _T_60089 = _T_60088[13:0]; // @[Modules.scala 160:64:@6027.4]
  assign buffer_1_554 = $signed(_T_60089); // @[Modules.scala 160:64:@6028.4]
  assign _T_60091 = $signed(buffer_1_502) + $signed(buffer_1_503); // @[Modules.scala 160:64:@6030.4]
  assign _T_60092 = _T_60091[13:0]; // @[Modules.scala 160:64:@6031.4]
  assign buffer_1_555 = $signed(_T_60092); // @[Modules.scala 160:64:@6032.4]
  assign _T_60094 = $signed(buffer_1_504) + $signed(buffer_1_505); // @[Modules.scala 160:64:@6034.4]
  assign _T_60095 = _T_60094[13:0]; // @[Modules.scala 160:64:@6035.4]
  assign buffer_1_556 = $signed(_T_60095); // @[Modules.scala 160:64:@6036.4]
  assign _T_60097 = $signed(buffer_1_506) + $signed(buffer_1_507); // @[Modules.scala 160:64:@6038.4]
  assign _T_60098 = _T_60097[13:0]; // @[Modules.scala 160:64:@6039.4]
  assign buffer_1_557 = $signed(_T_60098); // @[Modules.scala 160:64:@6040.4]
  assign _T_60100 = $signed(buffer_1_508) + $signed(buffer_1_509); // @[Modules.scala 160:64:@6042.4]
  assign _T_60101 = _T_60100[13:0]; // @[Modules.scala 160:64:@6043.4]
  assign buffer_1_558 = $signed(_T_60101); // @[Modules.scala 160:64:@6044.4]
  assign _T_60103 = $signed(buffer_1_510) + $signed(buffer_1_511); // @[Modules.scala 160:64:@6046.4]
  assign _T_60104 = _T_60103[13:0]; // @[Modules.scala 160:64:@6047.4]
  assign buffer_1_559 = $signed(_T_60104); // @[Modules.scala 160:64:@6048.4]
  assign _T_60106 = $signed(buffer_1_512) + $signed(buffer_1_513); // @[Modules.scala 160:64:@6050.4]
  assign _T_60107 = _T_60106[13:0]; // @[Modules.scala 160:64:@6051.4]
  assign buffer_1_560 = $signed(_T_60107); // @[Modules.scala 160:64:@6052.4]
  assign _T_60109 = $signed(buffer_1_514) + $signed(buffer_1_515); // @[Modules.scala 160:64:@6054.4]
  assign _T_60110 = _T_60109[13:0]; // @[Modules.scala 160:64:@6055.4]
  assign buffer_1_561 = $signed(_T_60110); // @[Modules.scala 160:64:@6056.4]
  assign _T_60112 = $signed(buffer_1_516) + $signed(buffer_1_517); // @[Modules.scala 160:64:@6058.4]
  assign _T_60113 = _T_60112[13:0]; // @[Modules.scala 160:64:@6059.4]
  assign buffer_1_562 = $signed(_T_60113); // @[Modules.scala 160:64:@6060.4]
  assign _T_60115 = $signed(buffer_1_518) + $signed(buffer_1_519); // @[Modules.scala 160:64:@6062.4]
  assign _T_60116 = _T_60115[13:0]; // @[Modules.scala 160:64:@6063.4]
  assign buffer_1_563 = $signed(_T_60116); // @[Modules.scala 160:64:@6064.4]
  assign _T_60118 = $signed(buffer_1_520) + $signed(buffer_1_521); // @[Modules.scala 160:64:@6066.4]
  assign _T_60119 = _T_60118[13:0]; // @[Modules.scala 160:64:@6067.4]
  assign buffer_1_564 = $signed(_T_60119); // @[Modules.scala 160:64:@6068.4]
  assign _T_60121 = $signed(buffer_1_522) + $signed(buffer_1_523); // @[Modules.scala 160:64:@6070.4]
  assign _T_60122 = _T_60121[13:0]; // @[Modules.scala 160:64:@6071.4]
  assign buffer_1_565 = $signed(_T_60122); // @[Modules.scala 160:64:@6072.4]
  assign _T_60124 = $signed(buffer_1_524) + $signed(buffer_1_525); // @[Modules.scala 160:64:@6074.4]
  assign _T_60125 = _T_60124[13:0]; // @[Modules.scala 160:64:@6075.4]
  assign buffer_1_566 = $signed(_T_60125); // @[Modules.scala 160:64:@6076.4]
  assign _T_60127 = $signed(buffer_1_526) + $signed(buffer_1_527); // @[Modules.scala 160:64:@6078.4]
  assign _T_60128 = _T_60127[13:0]; // @[Modules.scala 160:64:@6079.4]
  assign buffer_1_567 = $signed(_T_60128); // @[Modules.scala 160:64:@6080.4]
  assign _T_60130 = $signed(buffer_1_528) + $signed(buffer_1_529); // @[Modules.scala 160:64:@6082.4]
  assign _T_60131 = _T_60130[13:0]; // @[Modules.scala 160:64:@6083.4]
  assign buffer_1_568 = $signed(_T_60131); // @[Modules.scala 160:64:@6084.4]
  assign _T_60133 = $signed(buffer_1_530) + $signed(buffer_1_531); // @[Modules.scala 160:64:@6086.4]
  assign _T_60134 = _T_60133[13:0]; // @[Modules.scala 160:64:@6087.4]
  assign buffer_1_569 = $signed(_T_60134); // @[Modules.scala 160:64:@6088.4]
  assign _T_60136 = $signed(buffer_1_532) + $signed(buffer_1_533); // @[Modules.scala 160:64:@6090.4]
  assign _T_60137 = _T_60136[13:0]; // @[Modules.scala 160:64:@6091.4]
  assign buffer_1_570 = $signed(_T_60137); // @[Modules.scala 160:64:@6092.4]
  assign _T_60139 = $signed(buffer_1_534) + $signed(buffer_1_535); // @[Modules.scala 160:64:@6094.4]
  assign _T_60140 = _T_60139[13:0]; // @[Modules.scala 160:64:@6095.4]
  assign buffer_1_571 = $signed(_T_60140); // @[Modules.scala 160:64:@6096.4]
  assign _T_60142 = $signed(buffer_1_536) + $signed(buffer_1_537); // @[Modules.scala 160:64:@6098.4]
  assign _T_60143 = _T_60142[13:0]; // @[Modules.scala 160:64:@6099.4]
  assign buffer_1_572 = $signed(_T_60143); // @[Modules.scala 160:64:@6100.4]
  assign _T_60145 = $signed(buffer_1_538) + $signed(buffer_1_539); // @[Modules.scala 160:64:@6102.4]
  assign _T_60146 = _T_60145[13:0]; // @[Modules.scala 160:64:@6103.4]
  assign buffer_1_573 = $signed(_T_60146); // @[Modules.scala 160:64:@6104.4]
  assign _T_60148 = $signed(buffer_1_540) + $signed(buffer_1_541); // @[Modules.scala 160:64:@6106.4]
  assign _T_60149 = _T_60148[13:0]; // @[Modules.scala 160:64:@6107.4]
  assign buffer_1_574 = $signed(_T_60149); // @[Modules.scala 160:64:@6108.4]
  assign _T_60151 = $signed(buffer_1_542) + $signed(buffer_1_543); // @[Modules.scala 160:64:@6110.4]
  assign _T_60152 = _T_60151[13:0]; // @[Modules.scala 160:64:@6111.4]
  assign buffer_1_575 = $signed(_T_60152); // @[Modules.scala 160:64:@6112.4]
  assign _T_60154 = $signed(buffer_1_544) + $signed(buffer_1_545); // @[Modules.scala 160:64:@6114.4]
  assign _T_60155 = _T_60154[13:0]; // @[Modules.scala 160:64:@6115.4]
  assign buffer_1_576 = $signed(_T_60155); // @[Modules.scala 160:64:@6116.4]
  assign _T_60157 = $signed(buffer_1_546) + $signed(buffer_1_547); // @[Modules.scala 160:64:@6118.4]
  assign _T_60158 = _T_60157[13:0]; // @[Modules.scala 160:64:@6119.4]
  assign buffer_1_577 = $signed(_T_60158); // @[Modules.scala 160:64:@6120.4]
  assign _T_60160 = $signed(buffer_1_548) + $signed(buffer_1_549); // @[Modules.scala 160:64:@6122.4]
  assign _T_60161 = _T_60160[13:0]; // @[Modules.scala 160:64:@6123.4]
  assign buffer_1_578 = $signed(_T_60161); // @[Modules.scala 160:64:@6124.4]
  assign _T_60163 = $signed(buffer_1_550) + $signed(buffer_1_551); // @[Modules.scala 160:64:@6126.4]
  assign _T_60164 = _T_60163[13:0]; // @[Modules.scala 160:64:@6127.4]
  assign buffer_1_579 = $signed(_T_60164); // @[Modules.scala 160:64:@6128.4]
  assign _T_60166 = $signed(buffer_1_552) + $signed(buffer_1_553); // @[Modules.scala 160:64:@6130.4]
  assign _T_60167 = _T_60166[13:0]; // @[Modules.scala 160:64:@6131.4]
  assign buffer_1_580 = $signed(_T_60167); // @[Modules.scala 160:64:@6132.4]
  assign _T_60169 = $signed(buffer_1_554) + $signed(buffer_1_555); // @[Modules.scala 160:64:@6134.4]
  assign _T_60170 = _T_60169[13:0]; // @[Modules.scala 160:64:@6135.4]
  assign buffer_1_581 = $signed(_T_60170); // @[Modules.scala 160:64:@6136.4]
  assign _T_60172 = $signed(buffer_1_556) + $signed(buffer_1_557); // @[Modules.scala 160:64:@6138.4]
  assign _T_60173 = _T_60172[13:0]; // @[Modules.scala 160:64:@6139.4]
  assign buffer_1_582 = $signed(_T_60173); // @[Modules.scala 160:64:@6140.4]
  assign _T_60175 = $signed(buffer_1_558) + $signed(buffer_1_559); // @[Modules.scala 160:64:@6142.4]
  assign _T_60176 = _T_60175[13:0]; // @[Modules.scala 160:64:@6143.4]
  assign buffer_1_583 = $signed(_T_60176); // @[Modules.scala 160:64:@6144.4]
  assign _T_60178 = $signed(buffer_1_560) + $signed(buffer_1_561); // @[Modules.scala 160:64:@6146.4]
  assign _T_60179 = _T_60178[13:0]; // @[Modules.scala 160:64:@6147.4]
  assign buffer_1_584 = $signed(_T_60179); // @[Modules.scala 160:64:@6148.4]
  assign _T_60181 = $signed(buffer_1_562) + $signed(buffer_1_563); // @[Modules.scala 160:64:@6150.4]
  assign _T_60182 = _T_60181[13:0]; // @[Modules.scala 160:64:@6151.4]
  assign buffer_1_585 = $signed(_T_60182); // @[Modules.scala 160:64:@6152.4]
  assign _T_60184 = $signed(buffer_1_564) + $signed(buffer_1_565); // @[Modules.scala 160:64:@6154.4]
  assign _T_60185 = _T_60184[13:0]; // @[Modules.scala 160:64:@6155.4]
  assign buffer_1_586 = $signed(_T_60185); // @[Modules.scala 160:64:@6156.4]
  assign _T_60187 = $signed(buffer_1_566) + $signed(buffer_1_567); // @[Modules.scala 160:64:@6158.4]
  assign _T_60188 = _T_60187[13:0]; // @[Modules.scala 160:64:@6159.4]
  assign buffer_1_587 = $signed(_T_60188); // @[Modules.scala 160:64:@6160.4]
  assign _T_60190 = $signed(buffer_1_568) + $signed(buffer_1_569); // @[Modules.scala 160:64:@6162.4]
  assign _T_60191 = _T_60190[13:0]; // @[Modules.scala 160:64:@6163.4]
  assign buffer_1_588 = $signed(_T_60191); // @[Modules.scala 160:64:@6164.4]
  assign _T_60193 = $signed(buffer_1_570) + $signed(buffer_1_571); // @[Modules.scala 166:64:@6166.4]
  assign _T_60194 = _T_60193[13:0]; // @[Modules.scala 166:64:@6167.4]
  assign buffer_1_589 = $signed(_T_60194); // @[Modules.scala 166:64:@6168.4]
  assign _T_60196 = $signed(buffer_1_572) + $signed(buffer_1_573); // @[Modules.scala 166:64:@6170.4]
  assign _T_60197 = _T_60196[13:0]; // @[Modules.scala 166:64:@6171.4]
  assign buffer_1_590 = $signed(_T_60197); // @[Modules.scala 166:64:@6172.4]
  assign _T_60199 = $signed(buffer_1_574) + $signed(buffer_1_575); // @[Modules.scala 166:64:@6174.4]
  assign _T_60200 = _T_60199[13:0]; // @[Modules.scala 166:64:@6175.4]
  assign buffer_1_591 = $signed(_T_60200); // @[Modules.scala 166:64:@6176.4]
  assign _T_60202 = $signed(buffer_1_576) + $signed(buffer_1_577); // @[Modules.scala 166:64:@6178.4]
  assign _T_60203 = _T_60202[13:0]; // @[Modules.scala 166:64:@6179.4]
  assign buffer_1_592 = $signed(_T_60203); // @[Modules.scala 166:64:@6180.4]
  assign _T_60205 = $signed(buffer_1_578) + $signed(buffer_1_579); // @[Modules.scala 166:64:@6182.4]
  assign _T_60206 = _T_60205[13:0]; // @[Modules.scala 166:64:@6183.4]
  assign buffer_1_593 = $signed(_T_60206); // @[Modules.scala 166:64:@6184.4]
  assign _T_60208 = $signed(buffer_1_580) + $signed(buffer_1_581); // @[Modules.scala 166:64:@6186.4]
  assign _T_60209 = _T_60208[13:0]; // @[Modules.scala 166:64:@6187.4]
  assign buffer_1_594 = $signed(_T_60209); // @[Modules.scala 166:64:@6188.4]
  assign _T_60211 = $signed(buffer_1_582) + $signed(buffer_1_583); // @[Modules.scala 166:64:@6190.4]
  assign _T_60212 = _T_60211[13:0]; // @[Modules.scala 166:64:@6191.4]
  assign buffer_1_595 = $signed(_T_60212); // @[Modules.scala 166:64:@6192.4]
  assign _T_60214 = $signed(buffer_1_584) + $signed(buffer_1_585); // @[Modules.scala 166:64:@6194.4]
  assign _T_60215 = _T_60214[13:0]; // @[Modules.scala 166:64:@6195.4]
  assign buffer_1_596 = $signed(_T_60215); // @[Modules.scala 166:64:@6196.4]
  assign _T_60217 = $signed(buffer_1_586) + $signed(buffer_1_587); // @[Modules.scala 166:64:@6198.4]
  assign _T_60218 = _T_60217[13:0]; // @[Modules.scala 166:64:@6199.4]
  assign buffer_1_597 = $signed(_T_60218); // @[Modules.scala 166:64:@6200.4]
  assign _T_60220 = $signed(buffer_1_589) + $signed(buffer_1_590); // @[Modules.scala 166:64:@6202.4]
  assign _T_60221 = _T_60220[13:0]; // @[Modules.scala 166:64:@6203.4]
  assign buffer_1_598 = $signed(_T_60221); // @[Modules.scala 166:64:@6204.4]
  assign _T_60223 = $signed(buffer_1_591) + $signed(buffer_1_592); // @[Modules.scala 166:64:@6206.4]
  assign _T_60224 = _T_60223[13:0]; // @[Modules.scala 166:64:@6207.4]
  assign buffer_1_599 = $signed(_T_60224); // @[Modules.scala 166:64:@6208.4]
  assign _T_60226 = $signed(buffer_1_593) + $signed(buffer_1_594); // @[Modules.scala 166:64:@6210.4]
  assign _T_60227 = _T_60226[13:0]; // @[Modules.scala 166:64:@6211.4]
  assign buffer_1_600 = $signed(_T_60227); // @[Modules.scala 166:64:@6212.4]
  assign _T_60229 = $signed(buffer_1_595) + $signed(buffer_1_596); // @[Modules.scala 166:64:@6214.4]
  assign _T_60230 = _T_60229[13:0]; // @[Modules.scala 166:64:@6215.4]
  assign buffer_1_601 = $signed(_T_60230); // @[Modules.scala 166:64:@6216.4]
  assign _T_60232 = $signed(buffer_1_597) + $signed(buffer_1_588); // @[Modules.scala 172:66:@6218.4]
  assign _T_60233 = _T_60232[13:0]; // @[Modules.scala 172:66:@6219.4]
  assign buffer_1_602 = $signed(_T_60233); // @[Modules.scala 172:66:@6220.4]
  assign _T_60235 = $signed(buffer_1_598) + $signed(buffer_1_599); // @[Modules.scala 166:64:@6222.4]
  assign _T_60236 = _T_60235[13:0]; // @[Modules.scala 166:64:@6223.4]
  assign buffer_1_603 = $signed(_T_60236); // @[Modules.scala 166:64:@6224.4]
  assign _T_60238 = $signed(buffer_1_600) + $signed(buffer_1_601); // @[Modules.scala 166:64:@6226.4]
  assign _T_60239 = _T_60238[13:0]; // @[Modules.scala 166:64:@6227.4]
  assign buffer_1_604 = $signed(_T_60239); // @[Modules.scala 166:64:@6228.4]
  assign _T_60241 = $signed(buffer_1_603) + $signed(buffer_1_604); // @[Modules.scala 160:64:@6230.4]
  assign _T_60242 = _T_60241[13:0]; // @[Modules.scala 160:64:@6231.4]
  assign buffer_1_605 = $signed(_T_60242); // @[Modules.scala 160:64:@6232.4]
  assign _T_60244 = $signed(buffer_1_605) + $signed(buffer_1_602); // @[Modules.scala 172:66:@6234.4]
  assign _T_60245 = _T_60244[13:0]; // @[Modules.scala 172:66:@6235.4]
  assign buffer_1_606 = $signed(_T_60245); // @[Modules.scala 172:66:@6236.4]
  assign _T_60248 = $signed(-4'sh1) * $signed(io_in_12); // @[Modules.scala 143:74:@6415.4]
  assign _T_60250 = $signed(-4'sh1) * $signed(io_in_13); // @[Modules.scala 144:80:@6416.4]
  assign _T_60251 = $signed(_T_60248) + $signed(_T_60250); // @[Modules.scala 143:103:@6417.4]
  assign _T_60252 = _T_60251[4:0]; // @[Modules.scala 143:103:@6418.4]
  assign _T_60253 = $signed(_T_60252); // @[Modules.scala 143:103:@6419.4]
  assign _T_60255 = $signed(-4'sh1) * $signed(io_in_14); // @[Modules.scala 143:74:@6421.4]
  assign _T_60257 = $signed(-4'sh1) * $signed(io_in_15); // @[Modules.scala 144:80:@6422.4]
  assign _T_60258 = $signed(_T_60255) + $signed(_T_60257); // @[Modules.scala 143:103:@6423.4]
  assign _T_60259 = _T_60258[4:0]; // @[Modules.scala 143:103:@6424.4]
  assign _T_60260 = $signed(_T_60259); // @[Modules.scala 143:103:@6425.4]
  assign _T_60264 = $signed(-4'sh1) * $signed(io_in_33); // @[Modules.scala 144:80:@6428.4]
  assign _T_60265 = $signed(_T_57227) + $signed(_T_60264); // @[Modules.scala 143:103:@6429.4]
  assign _T_60266 = _T_60265[4:0]; // @[Modules.scala 143:103:@6430.4]
  assign _T_60267 = $signed(_T_60266); // @[Modules.scala 143:103:@6431.4]
  assign _T_60269 = $signed(-4'sh1) * $signed(io_in_34); // @[Modules.scala 143:74:@6433.4]
  assign _T_60271 = $signed(-4'sh1) * $signed(io_in_35); // @[Modules.scala 144:80:@6434.4]
  assign _T_60272 = $signed(_T_60269) + $signed(_T_60271); // @[Modules.scala 143:103:@6435.4]
  assign _T_60273 = _T_60272[4:0]; // @[Modules.scala 143:103:@6436.4]
  assign _T_60274 = $signed(_T_60273); // @[Modules.scala 143:103:@6437.4]
  assign _T_60279 = $signed(_T_54222) + $signed(_T_54227); // @[Modules.scala 143:103:@6441.4]
  assign _T_60280 = _T_60279[5:0]; // @[Modules.scala 143:103:@6442.4]
  assign _T_60281 = $signed(_T_60280); // @[Modules.scala 143:103:@6443.4]
  assign _T_60286 = $signed(_T_54229) + $signed(_T_54234); // @[Modules.scala 143:103:@6447.4]
  assign _T_60287 = _T_60286[5:0]; // @[Modules.scala 143:103:@6448.4]
  assign _T_60288 = $signed(_T_60287); // @[Modules.scala 143:103:@6449.4]
  assign _T_60293 = $signed(_T_57248) + $signed(_T_57253); // @[Modules.scala 143:103:@6453.4]
  assign _T_60294 = _T_60293[4:0]; // @[Modules.scala 143:103:@6454.4]
  assign _T_60295 = $signed(_T_60294); // @[Modules.scala 143:103:@6455.4]
  assign _T_60299 = $signed(-4'sh1) * $signed(io_in_44); // @[Modules.scala 144:80:@6458.4]
  assign _GEN_144 = {{1{_T_60299[4]}},_T_60299}; // @[Modules.scala 143:103:@6459.4]
  assign _T_60300 = $signed(_T_54243) + $signed(_GEN_144); // @[Modules.scala 143:103:@6459.4]
  assign _T_60301 = _T_60300[5:0]; // @[Modules.scala 143:103:@6460.4]
  assign _T_60302 = $signed(_T_60301); // @[Modules.scala 143:103:@6461.4]
  assign _T_60307 = $signed(_T_57262) + $signed(_T_57267); // @[Modules.scala 143:103:@6465.4]
  assign _T_60308 = _T_60307[4:0]; // @[Modules.scala 143:103:@6466.4]
  assign _T_60309 = $signed(_T_60308); // @[Modules.scala 143:103:@6467.4]
  assign _T_60327 = $signed(-4'sh1) * $signed(io_in_59); // @[Modules.scala 144:80:@6482.4]
  assign _T_60328 = $signed(_T_57281) + $signed(_T_60327); // @[Modules.scala 143:103:@6483.4]
  assign _T_60329 = _T_60328[4:0]; // @[Modules.scala 143:103:@6484.4]
  assign _T_60330 = $signed(_T_60329); // @[Modules.scala 143:103:@6485.4]
  assign _T_60332 = $signed(-4'sh1) * $signed(io_in_61); // @[Modules.scala 143:74:@6487.4]
  assign _T_60334 = $signed(-4'sh1) * $signed(io_in_62); // @[Modules.scala 144:80:@6488.4]
  assign _T_60335 = $signed(_T_60332) + $signed(_T_60334); // @[Modules.scala 143:103:@6489.4]
  assign _T_60336 = _T_60335[4:0]; // @[Modules.scala 143:103:@6490.4]
  assign _T_60337 = $signed(_T_60336); // @[Modules.scala 143:103:@6491.4]
  assign _T_60342 = $signed(_T_57297) + $signed(_T_57309); // @[Modules.scala 143:103:@6495.4]
  assign _T_60343 = _T_60342[4:0]; // @[Modules.scala 143:103:@6496.4]
  assign _T_60344 = $signed(_T_60343); // @[Modules.scala 143:103:@6497.4]
  assign _T_60349 = $signed(_T_57311) + $signed(_T_57316); // @[Modules.scala 143:103:@6501.4]
  assign _T_60350 = _T_60349[4:0]; // @[Modules.scala 143:103:@6502.4]
  assign _T_60351 = $signed(_T_60350); // @[Modules.scala 143:103:@6503.4]
  assign _T_60356 = $signed(_T_57318) + $signed(_T_57323); // @[Modules.scala 143:103:@6507.4]
  assign _T_60357 = _T_60356[4:0]; // @[Modules.scala 143:103:@6508.4]
  assign _T_60358 = $signed(_T_60357); // @[Modules.scala 143:103:@6509.4]
  assign _T_60363 = $signed(_T_57325) + $signed(_T_57330); // @[Modules.scala 143:103:@6513.4]
  assign _T_60364 = _T_60363[4:0]; // @[Modules.scala 143:103:@6514.4]
  assign _T_60365 = $signed(_T_60364); // @[Modules.scala 143:103:@6515.4]
  assign _GEN_145 = {{1{_T_57332[4]}},_T_57332}; // @[Modules.scala 143:103:@6519.4]
  assign _T_60370 = $signed(_GEN_145) + $signed(_T_54332); // @[Modules.scala 143:103:@6519.4]
  assign _T_60371 = _T_60370[5:0]; // @[Modules.scala 143:103:@6520.4]
  assign _T_60372 = $signed(_T_60371); // @[Modules.scala 143:103:@6521.4]
  assign _T_60402 = $signed(-4'sh1) * $signed(io_in_88); // @[Modules.scala 143:74:@6547.4]
  assign _T_60404 = $signed(-4'sh1) * $signed(io_in_89); // @[Modules.scala 144:80:@6548.4]
  assign _T_60405 = $signed(_T_60402) + $signed(_T_60404); // @[Modules.scala 143:103:@6549.4]
  assign _T_60406 = _T_60405[4:0]; // @[Modules.scala 143:103:@6550.4]
  assign _T_60407 = $signed(_T_60406); // @[Modules.scala 143:103:@6551.4]
  assign _T_60412 = $signed(_T_54369) + $signed(_T_54374); // @[Modules.scala 143:103:@6555.4]
  assign _T_60413 = _T_60412[5:0]; // @[Modules.scala 143:103:@6556.4]
  assign _T_60414 = $signed(_T_60413); // @[Modules.scala 143:103:@6557.4]
  assign _GEN_147 = {{1{_T_57395[4]}},_T_57395}; // @[Modules.scala 143:103:@6561.4]
  assign _T_60419 = $signed(_T_54381) + $signed(_GEN_147); // @[Modules.scala 143:103:@6561.4]
  assign _T_60420 = _T_60419[5:0]; // @[Modules.scala 143:103:@6562.4]
  assign _T_60421 = $signed(_T_60420); // @[Modules.scala 143:103:@6563.4]
  assign _T_60430 = $signed(-4'sh1) * $signed(io_in_98); // @[Modules.scala 143:74:@6571.4]
  assign _GEN_148 = {{1{_T_60430[4]}},_T_60430}; // @[Modules.scala 143:103:@6573.4]
  assign _T_60433 = $signed(_GEN_148) + $signed(_T_54402); // @[Modules.scala 143:103:@6573.4]
  assign _T_60434 = _T_60433[5:0]; // @[Modules.scala 143:103:@6574.4]
  assign _T_60435 = $signed(_T_60434); // @[Modules.scala 143:103:@6575.4]
  assign _T_60440 = $signed(_T_54404) + $signed(_T_54409); // @[Modules.scala 143:103:@6579.4]
  assign _T_60441 = _T_60440[5:0]; // @[Modules.scala 143:103:@6580.4]
  assign _T_60442 = $signed(_T_60441); // @[Modules.scala 143:103:@6581.4]
  assign _T_60447 = $signed(_T_54411) + $signed(_T_54416); // @[Modules.scala 143:103:@6585.4]
  assign _T_60448 = _T_60447[5:0]; // @[Modules.scala 143:103:@6586.4]
  assign _T_60449 = $signed(_T_60448); // @[Modules.scala 143:103:@6587.4]
  assign _T_60454 = $signed(_T_54418) + $signed(_T_54423); // @[Modules.scala 143:103:@6591.4]
  assign _T_60455 = _T_60454[5:0]; // @[Modules.scala 143:103:@6592.4]
  assign _T_60456 = $signed(_T_60455); // @[Modules.scala 143:103:@6593.4]
  assign _T_60461 = $signed(_T_54425) + $signed(_T_54430); // @[Modules.scala 143:103:@6597.4]
  assign _T_60462 = _T_60461[5:0]; // @[Modules.scala 143:103:@6598.4]
  assign _T_60463 = $signed(_T_60462); // @[Modules.scala 143:103:@6599.4]
  assign _T_60468 = $signed(_T_54432) + $signed(_T_54437); // @[Modules.scala 143:103:@6603.4]
  assign _T_60469 = _T_60468[5:0]; // @[Modules.scala 143:103:@6604.4]
  assign _T_60470 = $signed(_T_60469); // @[Modules.scala 143:103:@6605.4]
  assign _T_60474 = $signed(-4'sh1) * $signed(io_in_113); // @[Modules.scala 144:80:@6608.4]
  assign _T_60475 = $signed(_T_54439) + $signed(_T_60474); // @[Modules.scala 143:103:@6609.4]
  assign _T_60476 = _T_60475[4:0]; // @[Modules.scala 143:103:@6610.4]
  assign _T_60477 = $signed(_T_60476); // @[Modules.scala 143:103:@6611.4]
  assign _T_60482 = $signed(_GEN_3) + $signed(_T_57456); // @[Modules.scala 143:103:@6615.4]
  assign _T_60483 = _T_60482[5:0]; // @[Modules.scala 143:103:@6616.4]
  assign _T_60484 = $signed(_T_60483); // @[Modules.scala 143:103:@6617.4]
  assign _T_60488 = $signed(4'sh1) * $signed(io_in_119); // @[Modules.scala 144:80:@6620.4]
  assign _T_60489 = $signed(_T_57458) + $signed(_T_60488); // @[Modules.scala 143:103:@6621.4]
  assign _T_60490 = _T_60489[5:0]; // @[Modules.scala 143:103:@6622.4]
  assign _T_60491 = $signed(_T_60490); // @[Modules.scala 143:103:@6623.4]
  assign _T_60495 = $signed(-4'sh1) * $signed(io_in_122); // @[Modules.scala 144:80:@6626.4]
  assign _GEN_150 = {{1{_T_60495[4]}},_T_60495}; // @[Modules.scala 143:103:@6627.4]
  assign _T_60496 = $signed(_T_54460) + $signed(_GEN_150); // @[Modules.scala 143:103:@6627.4]
  assign _T_60497 = _T_60496[5:0]; // @[Modules.scala 143:103:@6628.4]
  assign _T_60498 = $signed(_T_60497); // @[Modules.scala 143:103:@6629.4]
  assign _T_60500 = $signed(-4'sh1) * $signed(io_in_123); // @[Modules.scala 143:74:@6631.4]
  assign _T_60502 = $signed(-4'sh1) * $signed(io_in_124); // @[Modules.scala 144:80:@6632.4]
  assign _T_60503 = $signed(_T_60500) + $signed(_T_60502); // @[Modules.scala 143:103:@6633.4]
  assign _T_60504 = _T_60503[4:0]; // @[Modules.scala 143:103:@6634.4]
  assign _T_60505 = $signed(_T_60504); // @[Modules.scala 143:103:@6635.4]
  assign _T_60507 = $signed(-4'sh1) * $signed(io_in_125); // @[Modules.scala 143:74:@6637.4]
  assign _T_60509 = $signed(-4'sh1) * $signed(io_in_126); // @[Modules.scala 144:80:@6638.4]
  assign _T_60510 = $signed(_T_60507) + $signed(_T_60509); // @[Modules.scala 143:103:@6639.4]
  assign _T_60511 = _T_60510[4:0]; // @[Modules.scala 143:103:@6640.4]
  assign _T_60512 = $signed(_T_60511); // @[Modules.scala 143:103:@6641.4]
  assign _T_60514 = $signed(-4'sh1) * $signed(io_in_127); // @[Modules.scala 143:74:@6643.4]
  assign _GEN_151 = {{1{_T_60514[4]}},_T_60514}; // @[Modules.scala 143:103:@6645.4]
  assign _T_60517 = $signed(_GEN_151) + $signed(_T_54488); // @[Modules.scala 143:103:@6645.4]
  assign _T_60518 = _T_60517[5:0]; // @[Modules.scala 143:103:@6646.4]
  assign _T_60519 = $signed(_T_60518); // @[Modules.scala 143:103:@6647.4]
  assign _T_60544 = $signed(-4'sh1) * $signed(io_in_138); // @[Modules.scala 144:80:@6668.4]
  assign _GEN_152 = {{1{_T_60544[4]}},_T_60544}; // @[Modules.scala 143:103:@6669.4]
  assign _T_60545 = $signed(_T_57512) + $signed(_GEN_152); // @[Modules.scala 143:103:@6669.4]
  assign _T_60546 = _T_60545[5:0]; // @[Modules.scala 143:103:@6670.4]
  assign _T_60547 = $signed(_T_60546); // @[Modules.scala 143:103:@6671.4]
  assign _T_60549 = $signed(4'sh1) * $signed(io_in_139); // @[Modules.scala 143:74:@6673.4]
  assign _T_60551 = $signed(-4'sh1) * $signed(io_in_142); // @[Modules.scala 144:80:@6674.4]
  assign _GEN_153 = {{1{_T_60551[4]}},_T_60551}; // @[Modules.scala 143:103:@6675.4]
  assign _T_60552 = $signed(_T_60549) + $signed(_GEN_153); // @[Modules.scala 143:103:@6675.4]
  assign _T_60553 = _T_60552[5:0]; // @[Modules.scala 143:103:@6676.4]
  assign _T_60554 = $signed(_T_60553); // @[Modules.scala 143:103:@6677.4]
  assign _T_60556 = $signed(-4'sh1) * $signed(io_in_143); // @[Modules.scala 143:74:@6679.4]
  assign _GEN_154 = {{1{_T_60556[4]}},_T_60556}; // @[Modules.scala 143:103:@6681.4]
  assign _T_60559 = $signed(_GEN_154) + $signed(_T_57533); // @[Modules.scala 143:103:@6681.4]
  assign _T_60560 = _T_60559[5:0]; // @[Modules.scala 143:103:@6682.4]
  assign _T_60561 = $signed(_T_60560); // @[Modules.scala 143:103:@6683.4]
  assign _T_60563 = $signed(-4'sh1) * $signed(io_in_145); // @[Modules.scala 143:74:@6685.4]
  assign _T_60566 = $signed(_T_60563) + $signed(_T_54523); // @[Modules.scala 143:103:@6687.4]
  assign _T_60567 = _T_60566[4:0]; // @[Modules.scala 143:103:@6688.4]
  assign _T_60568 = $signed(_T_60567); // @[Modules.scala 143:103:@6689.4]
  assign _T_60573 = $signed(_T_57542) + $signed(_T_54530); // @[Modules.scala 143:103:@6693.4]
  assign _T_60574 = _T_60573[5:0]; // @[Modules.scala 143:103:@6694.4]
  assign _T_60575 = $signed(_T_60574); // @[Modules.scala 143:103:@6695.4]
  assign _T_60577 = $signed(-4'sh1) * $signed(io_in_150); // @[Modules.scala 143:74:@6697.4]
  assign _T_60579 = $signed(-4'sh1) * $signed(io_in_151); // @[Modules.scala 144:80:@6698.4]
  assign _T_60580 = $signed(_T_60577) + $signed(_T_60579); // @[Modules.scala 143:103:@6699.4]
  assign _T_60581 = _T_60580[4:0]; // @[Modules.scala 143:103:@6700.4]
  assign _T_60582 = $signed(_T_60581); // @[Modules.scala 143:103:@6701.4]
  assign _T_60584 = $signed(-4'sh1) * $signed(io_in_152); // @[Modules.scala 143:74:@6703.4]
  assign _T_60586 = $signed(-4'sh1) * $signed(io_in_153); // @[Modules.scala 144:80:@6704.4]
  assign _T_60587 = $signed(_T_60584) + $signed(_T_60586); // @[Modules.scala 143:103:@6705.4]
  assign _T_60588 = _T_60587[4:0]; // @[Modules.scala 143:103:@6706.4]
  assign _T_60589 = $signed(_T_60588); // @[Modules.scala 143:103:@6707.4]
  assign _T_60605 = $signed(4'sh1) * $signed(io_in_159); // @[Modules.scala 143:74:@6721.4]
  assign _T_60607 = $signed(-4'sh1) * $signed(io_in_161); // @[Modules.scala 144:80:@6722.4]
  assign _GEN_155 = {{1{_T_60607[4]}},_T_60607}; // @[Modules.scala 143:103:@6723.4]
  assign _T_60608 = $signed(_T_60605) + $signed(_GEN_155); // @[Modules.scala 143:103:@6723.4]
  assign _T_60609 = _T_60608[5:0]; // @[Modules.scala 143:103:@6724.4]
  assign _T_60610 = $signed(_T_60609); // @[Modules.scala 143:103:@6725.4]
  assign _T_60614 = $signed(4'sh1) * $signed(io_in_163); // @[Modules.scala 144:80:@6728.4]
  assign _T_60615 = $signed(_GEN_10) + $signed(_T_60614); // @[Modules.scala 143:103:@6729.4]
  assign _T_60616 = _T_60615[5:0]; // @[Modules.scala 143:103:@6730.4]
  assign _T_60617 = $signed(_T_60616); // @[Modules.scala 143:103:@6731.4]
  assign _T_60619 = $signed(4'sh1) * $signed(io_in_164); // @[Modules.scala 143:74:@6733.4]
  assign _T_60622 = $signed(_T_60619) + $signed(_GEN_11); // @[Modules.scala 143:103:@6735.4]
  assign _T_60623 = _T_60622[5:0]; // @[Modules.scala 143:103:@6736.4]
  assign _T_60624 = $signed(_T_60623); // @[Modules.scala 143:103:@6737.4]
  assign _T_60628 = $signed(4'sh1) * $signed(io_in_169); // @[Modules.scala 144:80:@6740.4]
  assign _T_60629 = $signed(_GEN_88) + $signed(_T_60628); // @[Modules.scala 143:103:@6741.4]
  assign _T_60630 = _T_60629[5:0]; // @[Modules.scala 143:103:@6742.4]
  assign _T_60631 = $signed(_T_60630); // @[Modules.scala 143:103:@6743.4]
  assign _T_60633 = $signed(4'sh1) * $signed(io_in_170); // @[Modules.scala 143:74:@6745.4]
  assign _T_60635 = $signed(-4'sh1) * $signed(io_in_171); // @[Modules.scala 144:80:@6746.4]
  assign _GEN_159 = {{1{_T_60635[4]}},_T_60635}; // @[Modules.scala 143:103:@6747.4]
  assign _T_60636 = $signed(_T_60633) + $signed(_GEN_159); // @[Modules.scala 143:103:@6747.4]
  assign _T_60637 = _T_60636[5:0]; // @[Modules.scala 143:103:@6748.4]
  assign _T_60638 = $signed(_T_60637); // @[Modules.scala 143:103:@6749.4]
  assign _T_60642 = $signed(-4'sh1) * $signed(io_in_173); // @[Modules.scala 144:80:@6752.4]
  assign _GEN_160 = {{1{_T_60642[4]}},_T_60642}; // @[Modules.scala 143:103:@6753.4]
  assign _T_60643 = $signed(_T_54591) + $signed(_GEN_160); // @[Modules.scala 143:103:@6753.4]
  assign _T_60644 = _T_60643[5:0]; // @[Modules.scala 143:103:@6754.4]
  assign _T_60645 = $signed(_T_60644); // @[Modules.scala 143:103:@6755.4]
  assign _T_60647 = $signed(-4'sh1) * $signed(io_in_174); // @[Modules.scala 143:74:@6757.4]
  assign _GEN_161 = {{1{_T_60647[4]}},_T_60647}; // @[Modules.scala 143:103:@6759.4]
  assign _T_60650 = $signed(_GEN_161) + $signed(_T_54600); // @[Modules.scala 143:103:@6759.4]
  assign _T_60651 = _T_60650[5:0]; // @[Modules.scala 143:103:@6760.4]
  assign _T_60652 = $signed(_T_60651); // @[Modules.scala 143:103:@6761.4]
  assign _T_60656 = $signed(-4'sh1) * $signed(io_in_179); // @[Modules.scala 144:80:@6764.4]
  assign _T_60657 = $signed(_T_54607) + $signed(_T_60656); // @[Modules.scala 143:103:@6765.4]
  assign _T_60658 = _T_60657[4:0]; // @[Modules.scala 143:103:@6766.4]
  assign _T_60659 = $signed(_T_60658); // @[Modules.scala 143:103:@6767.4]
  assign _T_60668 = $signed(-4'sh1) * $signed(io_in_182); // @[Modules.scala 143:74:@6775.4]
  assign _T_60671 = $signed(_T_60668) + $signed(_T_54619); // @[Modules.scala 143:103:@6777.4]
  assign _T_60672 = _T_60671[4:0]; // @[Modules.scala 143:103:@6778.4]
  assign _T_60673 = $signed(_T_60672); // @[Modules.scala 143:103:@6779.4]
  assign _T_60678 = $signed(_T_54621) + $signed(_T_54626); // @[Modules.scala 143:103:@6783.4]
  assign _T_60679 = _T_60678[4:0]; // @[Modules.scala 143:103:@6784.4]
  assign _T_60680 = $signed(_T_60679); // @[Modules.scala 143:103:@6785.4]
  assign _T_60689 = $signed(-4'sh1) * $signed(io_in_188); // @[Modules.scala 143:74:@6793.4]
  assign _T_60691 = $signed(-4'sh1) * $signed(io_in_189); // @[Modules.scala 144:80:@6794.4]
  assign _T_60692 = $signed(_T_60689) + $signed(_T_60691); // @[Modules.scala 143:103:@6795.4]
  assign _T_60693 = _T_60692[4:0]; // @[Modules.scala 143:103:@6796.4]
  assign _T_60694 = $signed(_T_60693); // @[Modules.scala 143:103:@6797.4]
  assign _T_60698 = $signed(4'sh1) * $signed(io_in_191); // @[Modules.scala 144:80:@6800.4]
  assign _GEN_162 = {{1{_T_54635[4]}},_T_54635}; // @[Modules.scala 143:103:@6801.4]
  assign _T_60699 = $signed(_GEN_162) + $signed(_T_60698); // @[Modules.scala 143:103:@6801.4]
  assign _T_60700 = _T_60699[5:0]; // @[Modules.scala 143:103:@6802.4]
  assign _T_60701 = $signed(_T_60700); // @[Modules.scala 143:103:@6803.4]
  assign _T_60717 = $signed(-4'sh1) * $signed(io_in_199); // @[Modules.scala 143:74:@6817.4]
  assign _T_60719 = $signed(-4'sh1) * $signed(io_in_200); // @[Modules.scala 144:80:@6818.4]
  assign _T_60720 = $signed(_T_60717) + $signed(_T_60719); // @[Modules.scala 143:103:@6819.4]
  assign _T_60721 = _T_60720[4:0]; // @[Modules.scala 143:103:@6820.4]
  assign _T_60722 = $signed(_T_60721); // @[Modules.scala 143:103:@6821.4]
  assign _T_60724 = $signed(-4'sh1) * $signed(io_in_201); // @[Modules.scala 143:74:@6823.4]
  assign _T_60726 = $signed(-4'sh1) * $signed(io_in_202); // @[Modules.scala 144:80:@6824.4]
  assign _T_60727 = $signed(_T_60724) + $signed(_T_60726); // @[Modules.scala 143:103:@6825.4]
  assign _T_60728 = _T_60727[4:0]; // @[Modules.scala 143:103:@6826.4]
  assign _T_60729 = $signed(_T_60728); // @[Modules.scala 143:103:@6827.4]
  assign _T_60733 = $signed(-4'sh1) * $signed(io_in_204); // @[Modules.scala 144:80:@6830.4]
  assign _GEN_164 = {{1{_T_60733[4]}},_T_60733}; // @[Modules.scala 143:103:@6831.4]
  assign _T_60734 = $signed(_T_54682) + $signed(_GEN_164); // @[Modules.scala 143:103:@6831.4]
  assign _T_60735 = _T_60734[5:0]; // @[Modules.scala 143:103:@6832.4]
  assign _T_60736 = $signed(_T_60735); // @[Modules.scala 143:103:@6833.4]
  assign _T_60740 = $signed(-4'sh1) * $signed(io_in_206); // @[Modules.scala 144:80:@6836.4]
  assign _T_60741 = $signed(_T_54684) + $signed(_T_60740); // @[Modules.scala 143:103:@6837.4]
  assign _T_60742 = _T_60741[4:0]; // @[Modules.scala 143:103:@6838.4]
  assign _T_60743 = $signed(_T_60742); // @[Modules.scala 143:103:@6839.4]
  assign _T_60745 = $signed(-4'sh1) * $signed(io_in_207); // @[Modules.scala 143:74:@6841.4]
  assign _T_60747 = $signed(-4'sh1) * $signed(io_in_208); // @[Modules.scala 144:80:@6842.4]
  assign _T_60748 = $signed(_T_60745) + $signed(_T_60747); // @[Modules.scala 143:103:@6843.4]
  assign _T_60749 = _T_60748[4:0]; // @[Modules.scala 143:103:@6844.4]
  assign _T_60750 = $signed(_T_60749); // @[Modules.scala 143:103:@6845.4]
  assign _T_60752 = $signed(-4'sh1) * $signed(io_in_209); // @[Modules.scala 143:74:@6847.4]
  assign _T_60754 = $signed(-4'sh1) * $signed(io_in_210); // @[Modules.scala 144:80:@6848.4]
  assign _T_60755 = $signed(_T_60752) + $signed(_T_60754); // @[Modules.scala 143:103:@6849.4]
  assign _T_60756 = _T_60755[4:0]; // @[Modules.scala 143:103:@6850.4]
  assign _T_60757 = $signed(_T_60756); // @[Modules.scala 143:103:@6851.4]
  assign _T_60759 = $signed(-4'sh1) * $signed(io_in_211); // @[Modules.scala 143:74:@6853.4]
  assign _T_60762 = $signed(_T_60759) + $signed(_T_54691); // @[Modules.scala 143:103:@6855.4]
  assign _T_60763 = _T_60762[4:0]; // @[Modules.scala 143:103:@6856.4]
  assign _T_60764 = $signed(_T_60763); // @[Modules.scala 143:103:@6857.4]
  assign _T_60773 = $signed(-4'sh1) * $signed(io_in_215); // @[Modules.scala 143:74:@6865.4]
  assign _T_60776 = $signed(_T_60773) + $signed(_T_54703); // @[Modules.scala 143:103:@6867.4]
  assign _T_60777 = _T_60776[4:0]; // @[Modules.scala 143:103:@6868.4]
  assign _T_60778 = $signed(_T_60777); // @[Modules.scala 143:103:@6869.4]
  assign _T_60783 = $signed(_T_54705) + $signed(_T_54710); // @[Modules.scala 143:103:@6873.4]
  assign _T_60784 = _T_60783[4:0]; // @[Modules.scala 143:103:@6874.4]
  assign _T_60785 = $signed(_T_60784); // @[Modules.scala 143:103:@6875.4]
  assign _T_60808 = $signed(-4'sh1) * $signed(io_in_226); // @[Modules.scala 143:74:@6895.4]
  assign _T_60810 = $signed(-4'sh1) * $signed(io_in_227); // @[Modules.scala 144:80:@6896.4]
  assign _T_60811 = $signed(_T_60808) + $signed(_T_60810); // @[Modules.scala 143:103:@6897.4]
  assign _T_60812 = _T_60811[4:0]; // @[Modules.scala 143:103:@6898.4]
  assign _T_60813 = $signed(_T_60812); // @[Modules.scala 143:103:@6899.4]
  assign _T_60815 = $signed(-4'sh1) * $signed(io_in_228); // @[Modules.scala 143:74:@6901.4]
  assign _T_60817 = $signed(-4'sh1) * $signed(io_in_229); // @[Modules.scala 144:80:@6902.4]
  assign _T_60818 = $signed(_T_60815) + $signed(_T_60817); // @[Modules.scala 143:103:@6903.4]
  assign _T_60819 = _T_60818[4:0]; // @[Modules.scala 143:103:@6904.4]
  assign _T_60820 = $signed(_T_60819); // @[Modules.scala 143:103:@6905.4]
  assign _T_60822 = $signed(-4'sh1) * $signed(io_in_230); // @[Modules.scala 143:74:@6907.4]
  assign _T_60825 = $signed(_T_60822) + $signed(_T_57787); // @[Modules.scala 143:103:@6909.4]
  assign _T_60826 = _T_60825[4:0]; // @[Modules.scala 143:103:@6910.4]
  assign _T_60827 = $signed(_T_60826); // @[Modules.scala 143:103:@6911.4]
  assign _T_60829 = $signed(-4'sh1) * $signed(io_in_232); // @[Modules.scala 143:74:@6913.4]
  assign _T_60831 = $signed(-4'sh1) * $signed(io_in_234); // @[Modules.scala 144:80:@6914.4]
  assign _T_60832 = $signed(_T_60829) + $signed(_T_60831); // @[Modules.scala 143:103:@6915.4]
  assign _T_60833 = _T_60832[4:0]; // @[Modules.scala 143:103:@6916.4]
  assign _T_60834 = $signed(_T_60833); // @[Modules.scala 143:103:@6917.4]
  assign _T_60838 = $signed(-4'sh1) * $signed(io_in_236); // @[Modules.scala 144:80:@6920.4]
  assign _GEN_165 = {{1{_T_60838[4]}},_T_60838}; // @[Modules.scala 143:103:@6921.4]
  assign _T_60839 = $signed(_T_54761) + $signed(_GEN_165); // @[Modules.scala 143:103:@6921.4]
  assign _T_60840 = _T_60839[5:0]; // @[Modules.scala 143:103:@6922.4]
  assign _T_60841 = $signed(_T_60840); // @[Modules.scala 143:103:@6923.4]
  assign _T_60843 = $signed(-4'sh1) * $signed(io_in_237); // @[Modules.scala 143:74:@6925.4]
  assign _T_60845 = $signed(-4'sh1) * $signed(io_in_238); // @[Modules.scala 144:80:@6926.4]
  assign _T_60846 = $signed(_T_60843) + $signed(_T_60845); // @[Modules.scala 143:103:@6927.4]
  assign _T_60847 = _T_60846[4:0]; // @[Modules.scala 143:103:@6928.4]
  assign _T_60848 = $signed(_T_60847); // @[Modules.scala 143:103:@6929.4]
  assign _T_60850 = $signed(-4'sh1) * $signed(io_in_239); // @[Modules.scala 143:74:@6931.4]
  assign _T_60853 = $signed(_T_60850) + $signed(_T_54768); // @[Modules.scala 143:103:@6933.4]
  assign _T_60854 = _T_60853[4:0]; // @[Modules.scala 143:103:@6934.4]
  assign _T_60855 = $signed(_T_60854); // @[Modules.scala 143:103:@6935.4]
  assign _T_60860 = $signed(_T_54773) + $signed(_T_54780); // @[Modules.scala 143:103:@6939.4]
  assign _T_60861 = _T_60860[4:0]; // @[Modules.scala 143:103:@6940.4]
  assign _T_60862 = $signed(_T_60861); // @[Modules.scala 143:103:@6941.4]
  assign _T_60867 = $signed(_T_54782) + $signed(_T_54787); // @[Modules.scala 143:103:@6945.4]
  assign _T_60868 = _T_60867[4:0]; // @[Modules.scala 143:103:@6946.4]
  assign _T_60869 = $signed(_T_60868); // @[Modules.scala 143:103:@6947.4]
  assign _T_60874 = $signed(_T_54789) + $signed(_T_54794); // @[Modules.scala 143:103:@6951.4]
  assign _T_60875 = _T_60874[4:0]; // @[Modules.scala 143:103:@6952.4]
  assign _T_60876 = $signed(_T_60875); // @[Modules.scala 143:103:@6953.4]
  assign _T_60881 = $signed(_T_54796) + $signed(_T_54801); // @[Modules.scala 143:103:@6957.4]
  assign _T_60882 = _T_60881[4:0]; // @[Modules.scala 143:103:@6958.4]
  assign _T_60883 = $signed(_T_60882); // @[Modules.scala 143:103:@6959.4]
  assign _T_60888 = $signed(_T_54803) + $signed(_T_57848); // @[Modules.scala 143:103:@6963.4]
  assign _T_60889 = _T_60888[4:0]; // @[Modules.scala 143:103:@6964.4]
  assign _T_60890 = $signed(_T_60889); // @[Modules.scala 143:103:@6965.4]
  assign _T_60895 = $signed(_GEN_21) + $signed(_T_54815); // @[Modules.scala 143:103:@6969.4]
  assign _T_60896 = _T_60895[5:0]; // @[Modules.scala 143:103:@6970.4]
  assign _T_60897 = $signed(_T_60896); // @[Modules.scala 143:103:@6971.4]
  assign _T_60899 = $signed(-4'sh1) * $signed(io_in_254); // @[Modules.scala 143:74:@6973.4]
  assign _T_60901 = $signed(-4'sh1) * $signed(io_in_255); // @[Modules.scala 144:80:@6974.4]
  assign _T_60902 = $signed(_T_60899) + $signed(_T_60901); // @[Modules.scala 143:103:@6975.4]
  assign _T_60903 = _T_60902[4:0]; // @[Modules.scala 143:103:@6976.4]
  assign _T_60904 = $signed(_T_60903); // @[Modules.scala 143:103:@6977.4]
  assign _T_60906 = $signed(-4'sh1) * $signed(io_in_256); // @[Modules.scala 143:74:@6979.4]
  assign _T_60908 = $signed(-4'sh1) * $signed(io_in_257); // @[Modules.scala 144:80:@6980.4]
  assign _T_60909 = $signed(_T_60906) + $signed(_T_60908); // @[Modules.scala 143:103:@6981.4]
  assign _T_60910 = _T_60909[4:0]; // @[Modules.scala 143:103:@6982.4]
  assign _T_60911 = $signed(_T_60910); // @[Modules.scala 143:103:@6983.4]
  assign _T_60913 = $signed(-4'sh1) * $signed(io_in_258); // @[Modules.scala 143:74:@6985.4]
  assign _T_60916 = $signed(_T_60913) + $signed(_T_57869); // @[Modules.scala 143:103:@6987.4]
  assign _T_60917 = _T_60916[4:0]; // @[Modules.scala 143:103:@6988.4]
  assign _T_60918 = $signed(_T_60917); // @[Modules.scala 143:103:@6989.4]
  assign _T_60920 = $signed(-4'sh1) * $signed(io_in_260); // @[Modules.scala 143:74:@6991.4]
  assign _T_60922 = $signed(4'sh1) * $signed(io_in_262); // @[Modules.scala 144:80:@6992.4]
  assign _GEN_167 = {{1{_T_60920[4]}},_T_60920}; // @[Modules.scala 143:103:@6993.4]
  assign _T_60923 = $signed(_GEN_167) + $signed(_T_60922); // @[Modules.scala 143:103:@6993.4]
  assign _T_60924 = _T_60923[5:0]; // @[Modules.scala 143:103:@6994.4]
  assign _T_60925 = $signed(_T_60924); // @[Modules.scala 143:103:@6995.4]
  assign _T_60930 = $signed(_T_54838) + $signed(_T_54843); // @[Modules.scala 143:103:@6999.4]
  assign _T_60931 = _T_60930[4:0]; // @[Modules.scala 143:103:@7000.4]
  assign _T_60932 = $signed(_T_60931); // @[Modules.scala 143:103:@7001.4]
  assign _T_60934 = $signed(-4'sh1) * $signed(io_in_266); // @[Modules.scala 143:74:@7003.4]
  assign _T_60936 = $signed(-4'sh1) * $signed(io_in_267); // @[Modules.scala 144:80:@7004.4]
  assign _T_60937 = $signed(_T_60934) + $signed(_T_60936); // @[Modules.scala 143:103:@7005.4]
  assign _T_60938 = _T_60937[4:0]; // @[Modules.scala 143:103:@7006.4]
  assign _T_60939 = $signed(_T_60938); // @[Modules.scala 143:103:@7007.4]
  assign _T_60944 = $signed(_T_54852) + $signed(_T_54857); // @[Modules.scala 143:103:@7011.4]
  assign _T_60945 = _T_60944[4:0]; // @[Modules.scala 143:103:@7012.4]
  assign _T_60946 = $signed(_T_60945); // @[Modules.scala 143:103:@7013.4]
  assign _T_60983 = $signed(-4'sh1) * $signed(io_in_282); // @[Modules.scala 143:74:@7045.4]
  assign _T_60985 = $signed(-4'sh1) * $signed(io_in_283); // @[Modules.scala 144:80:@7046.4]
  assign _T_60986 = $signed(_T_60983) + $signed(_T_60985); // @[Modules.scala 143:103:@7047.4]
  assign _T_60987 = _T_60986[4:0]; // @[Modules.scala 143:103:@7048.4]
  assign _T_60988 = $signed(_T_60987); // @[Modules.scala 143:103:@7049.4]
  assign _T_60993 = $signed(_T_54908) + $signed(_T_54913); // @[Modules.scala 143:103:@7053.4]
  assign _T_60994 = _T_60993[4:0]; // @[Modules.scala 143:103:@7054.4]
  assign _T_60995 = $signed(_T_60994); // @[Modules.scala 143:103:@7055.4]
  assign _T_61000 = $signed(_T_54915) + $signed(_T_54920); // @[Modules.scala 143:103:@7059.4]
  assign _T_61001 = _T_61000[4:0]; // @[Modules.scala 143:103:@7060.4]
  assign _T_61002 = $signed(_T_61001); // @[Modules.scala 143:103:@7061.4]
  assign _T_61004 = $signed(4'sh1) * $signed(io_in_288); // @[Modules.scala 143:74:@7063.4]
  assign _T_61006 = $signed(4'sh1) * $signed(io_in_290); // @[Modules.scala 144:80:@7064.4]
  assign _T_61007 = $signed(_T_61004) + $signed(_T_61006); // @[Modules.scala 143:103:@7065.4]
  assign _T_61008 = _T_61007[5:0]; // @[Modules.scala 143:103:@7066.4]
  assign _T_61009 = $signed(_T_61008); // @[Modules.scala 143:103:@7067.4]
  assign _T_61013 = $signed(-4'sh1) * $signed(io_in_294); // @[Modules.scala 144:80:@7070.4]
  assign _T_61014 = $signed(_T_54941) + $signed(_T_61013); // @[Modules.scala 143:103:@7071.4]
  assign _T_61015 = _T_61014[4:0]; // @[Modules.scala 143:103:@7072.4]
  assign _T_61016 = $signed(_T_61015); // @[Modules.scala 143:103:@7073.4]
  assign _T_61018 = $signed(-4'sh1) * $signed(io_in_295); // @[Modules.scala 143:74:@7075.4]
  assign _T_61020 = $signed(-4'sh1) * $signed(io_in_296); // @[Modules.scala 144:80:@7076.4]
  assign _T_61021 = $signed(_T_61018) + $signed(_T_61020); // @[Modules.scala 143:103:@7077.4]
  assign _T_61022 = _T_61021[4:0]; // @[Modules.scala 143:103:@7078.4]
  assign _T_61023 = $signed(_T_61022); // @[Modules.scala 143:103:@7079.4]
  assign _T_61025 = $signed(-4'sh1) * $signed(io_in_297); // @[Modules.scala 143:74:@7081.4]
  assign _T_61028 = $signed(_T_61025) + $signed(_T_54955); // @[Modules.scala 143:103:@7083.4]
  assign _T_61029 = _T_61028[4:0]; // @[Modules.scala 143:103:@7084.4]
  assign _T_61030 = $signed(_T_61029); // @[Modules.scala 143:103:@7085.4]
  assign _T_61035 = $signed(_T_54957) + $signed(_T_54962); // @[Modules.scala 143:103:@7089.4]
  assign _T_61036 = _T_61035[4:0]; // @[Modules.scala 143:103:@7090.4]
  assign _T_61037 = $signed(_T_61036); // @[Modules.scala 143:103:@7091.4]
  assign _T_61042 = $signed(_T_54964) + $signed(_T_54969); // @[Modules.scala 143:103:@7095.4]
  assign _T_61043 = _T_61042[4:0]; // @[Modules.scala 143:103:@7096.4]
  assign _T_61044 = $signed(_T_61043); // @[Modules.scala 143:103:@7097.4]
  assign _T_61062 = $signed(-4'sh1) * $signed(io_in_309); // @[Modules.scala 144:80:@7112.4]
  assign _GEN_168 = {{1{_T_61062[4]}},_T_61062}; // @[Modules.scala 143:103:@7113.4]
  assign _T_61063 = $signed(_T_58011) + $signed(_GEN_168); // @[Modules.scala 143:103:@7113.4]
  assign _T_61064 = _T_61063[5:0]; // @[Modules.scala 143:103:@7114.4]
  assign _T_61065 = $signed(_T_61064); // @[Modules.scala 143:103:@7115.4]
  assign _T_61069 = $signed(-4'sh1) * $signed(io_in_311); // @[Modules.scala 144:80:@7118.4]
  assign _T_61070 = $signed(_T_54992) + $signed(_T_61069); // @[Modules.scala 143:103:@7119.4]
  assign _T_61071 = _T_61070[4:0]; // @[Modules.scala 143:103:@7120.4]
  assign _T_61072 = $signed(_T_61071); // @[Modules.scala 143:103:@7121.4]
  assign _T_61077 = $signed(_T_54999) + $signed(_T_55004); // @[Modules.scala 143:103:@7125.4]
  assign _T_61078 = _T_61077[4:0]; // @[Modules.scala 143:103:@7126.4]
  assign _T_61079 = $signed(_T_61078); // @[Modules.scala 143:103:@7127.4]
  assign _T_61081 = $signed(4'sh1) * $signed(io_in_315); // @[Modules.scala 143:74:@7129.4]
  assign _T_61083 = $signed(4'sh1) * $signed(io_in_316); // @[Modules.scala 144:80:@7130.4]
  assign _T_61084 = $signed(_T_61081) + $signed(_T_61083); // @[Modules.scala 143:103:@7131.4]
  assign _T_61085 = _T_61084[5:0]; // @[Modules.scala 143:103:@7132.4]
  assign _T_61086 = $signed(_T_61085); // @[Modules.scala 143:103:@7133.4]
  assign _T_61088 = $signed(4'sh1) * $signed(io_in_317); // @[Modules.scala 143:74:@7135.4]
  assign _T_61090 = $signed(4'sh1) * $signed(io_in_318); // @[Modules.scala 144:80:@7136.4]
  assign _T_61091 = $signed(_T_61088) + $signed(_T_61090); // @[Modules.scala 143:103:@7137.4]
  assign _T_61092 = _T_61091[5:0]; // @[Modules.scala 143:103:@7138.4]
  assign _T_61093 = $signed(_T_61092); // @[Modules.scala 143:103:@7139.4]
  assign _T_61095 = $signed(4'sh1) * $signed(io_in_319); // @[Modules.scala 143:74:@7141.4]
  assign _T_61097 = $signed(4'sh1) * $signed(io_in_320); // @[Modules.scala 144:80:@7142.4]
  assign _T_61098 = $signed(_T_61095) + $signed(_T_61097); // @[Modules.scala 143:103:@7143.4]
  assign _T_61099 = _T_61098[5:0]; // @[Modules.scala 143:103:@7144.4]
  assign _T_61100 = $signed(_T_61099); // @[Modules.scala 143:103:@7145.4]
  assign _T_61104 = $signed(-4'sh1) * $signed(io_in_322); // @[Modules.scala 144:80:@7148.4]
  assign _T_61105 = $signed(_T_55032) + $signed(_T_61104); // @[Modules.scala 143:103:@7149.4]
  assign _T_61106 = _T_61105[4:0]; // @[Modules.scala 143:103:@7150.4]
  assign _T_61107 = $signed(_T_61106); // @[Modules.scala 143:103:@7151.4]
  assign _T_61109 = $signed(-4'sh1) * $signed(io_in_323); // @[Modules.scala 143:74:@7153.4]
  assign _GEN_169 = {{1{_T_61109[4]}},_T_61109}; // @[Modules.scala 143:103:@7155.4]
  assign _T_61112 = $signed(_GEN_169) + $signed(_T_58065); // @[Modules.scala 143:103:@7155.4]
  assign _T_61113 = _T_61112[5:0]; // @[Modules.scala 143:103:@7156.4]
  assign _T_61114 = $signed(_T_61113); // @[Modules.scala 143:103:@7157.4]
  assign _T_61119 = $signed(_T_58067) + $signed(_T_58072); // @[Modules.scala 143:103:@7161.4]
  assign _T_61120 = _T_61119[5:0]; // @[Modules.scala 143:103:@7162.4]
  assign _T_61121 = $signed(_T_61120); // @[Modules.scala 143:103:@7163.4]
  assign _GEN_170 = {{1{_T_58095[4]}},_T_58095}; // @[Modules.scala 143:103:@7185.4]
  assign _T_61147 = $signed(_GEN_170) + $signed(_T_58100); // @[Modules.scala 143:103:@7185.4]
  assign _T_61148 = _T_61147[5:0]; // @[Modules.scala 143:103:@7186.4]
  assign _T_61149 = $signed(_T_61148); // @[Modules.scala 143:103:@7187.4]
  assign _T_61153 = $signed(-4'sh1) * $signed(io_in_339); // @[Modules.scala 144:80:@7190.4]
  assign _T_61154 = $signed(_T_58109) + $signed(_T_61153); // @[Modules.scala 143:103:@7191.4]
  assign _T_61155 = _T_61154[4:0]; // @[Modules.scala 143:103:@7192.4]
  assign _T_61156 = $signed(_T_61155); // @[Modules.scala 143:103:@7193.4]
  assign _T_61160 = $signed(4'sh1) * $signed(io_in_342); // @[Modules.scala 144:80:@7196.4]
  assign _GEN_171 = {{1{_T_55088[4]}},_T_55088}; // @[Modules.scala 143:103:@7197.4]
  assign _T_61161 = $signed(_GEN_171) + $signed(_T_61160); // @[Modules.scala 143:103:@7197.4]
  assign _T_61162 = _T_61161[5:0]; // @[Modules.scala 143:103:@7198.4]
  assign _T_61163 = $signed(_T_61162); // @[Modules.scala 143:103:@7199.4]
  assign _T_61165 = $signed(4'sh1) * $signed(io_in_343); // @[Modules.scala 143:74:@7201.4]
  assign _T_61167 = $signed(4'sh1) * $signed(io_in_344); // @[Modules.scala 144:80:@7202.4]
  assign _T_61168 = $signed(_T_61165) + $signed(_T_61167); // @[Modules.scala 143:103:@7203.4]
  assign _T_61169 = _T_61168[5:0]; // @[Modules.scala 143:103:@7204.4]
  assign _T_61170 = $signed(_T_61169); // @[Modules.scala 143:103:@7205.4]
  assign _T_61172 = $signed(4'sh1) * $signed(io_in_345); // @[Modules.scala 143:74:@7207.4]
  assign _T_61174 = $signed(4'sh1) * $signed(io_in_346); // @[Modules.scala 144:80:@7208.4]
  assign _T_61175 = $signed(_T_61172) + $signed(_T_61174); // @[Modules.scala 143:103:@7209.4]
  assign _T_61176 = _T_61175[5:0]; // @[Modules.scala 143:103:@7210.4]
  assign _T_61177 = $signed(_T_61176); // @[Modules.scala 143:103:@7211.4]
  assign _T_61179 = $signed(4'sh1) * $signed(io_in_347); // @[Modules.scala 143:74:@7213.4]
  assign _T_61181 = $signed(4'sh1) * $signed(io_in_348); // @[Modules.scala 144:80:@7214.4]
  assign _T_61182 = $signed(_T_61179) + $signed(_T_61181); // @[Modules.scala 143:103:@7215.4]
  assign _T_61183 = _T_61182[5:0]; // @[Modules.scala 143:103:@7216.4]
  assign _T_61184 = $signed(_T_61183); // @[Modules.scala 143:103:@7217.4]
  assign _T_61188 = $signed(-4'sh1) * $signed(io_in_350); // @[Modules.scala 144:80:@7220.4]
  assign _GEN_172 = {{1{_T_61188[4]}},_T_61188}; // @[Modules.scala 143:103:@7221.4]
  assign _T_61189 = $signed(_T_58142) + $signed(_GEN_172); // @[Modules.scala 143:103:@7221.4]
  assign _T_61190 = _T_61189[5:0]; // @[Modules.scala 143:103:@7222.4]
  assign _T_61191 = $signed(_T_61190); // @[Modules.scala 143:103:@7223.4]
  assign _T_61210 = $signed(_T_58163) + $signed(_T_58170); // @[Modules.scala 143:103:@7239.4]
  assign _T_61211 = _T_61210[5:0]; // @[Modules.scala 143:103:@7240.4]
  assign _T_61212 = $signed(_T_61211); // @[Modules.scala 143:103:@7241.4]
  assign _T_61214 = $signed(4'sh1) * $signed(io_in_358); // @[Modules.scala 143:74:@7243.4]
  assign _T_61216 = $signed(4'sh1) * $signed(io_in_359); // @[Modules.scala 144:80:@7244.4]
  assign _T_61217 = $signed(_T_61214) + $signed(_T_61216); // @[Modules.scala 143:103:@7245.4]
  assign _T_61218 = _T_61217[5:0]; // @[Modules.scala 143:103:@7246.4]
  assign _T_61219 = $signed(_T_61218); // @[Modules.scala 143:103:@7247.4]
  assign _T_61224 = $signed(_T_58172) + $signed(_T_55153); // @[Modules.scala 143:103:@7251.4]
  assign _T_61225 = _T_61224[4:0]; // @[Modules.scala 143:103:@7252.4]
  assign _T_61226 = $signed(_T_61225); // @[Modules.scala 143:103:@7253.4]
  assign _T_61230 = $signed(-4'sh1) * $signed(io_in_363); // @[Modules.scala 144:80:@7256.4]
  assign _T_61231 = $signed(_T_55158) + $signed(_T_61230); // @[Modules.scala 143:103:@7257.4]
  assign _T_61232 = _T_61231[4:0]; // @[Modules.scala 143:103:@7258.4]
  assign _T_61233 = $signed(_T_61232); // @[Modules.scala 143:103:@7259.4]
  assign _T_61235 = $signed(-4'sh1) * $signed(io_in_364); // @[Modules.scala 143:74:@7261.4]
  assign _GEN_173 = {{1{_T_61235[4]}},_T_61235}; // @[Modules.scala 143:103:@7263.4]
  assign _T_61238 = $signed(_GEN_173) + $signed(_T_55167); // @[Modules.scala 143:103:@7263.4]
  assign _T_61239 = _T_61238[5:0]; // @[Modules.scala 143:103:@7264.4]
  assign _T_61240 = $signed(_T_61239); // @[Modules.scala 143:103:@7265.4]
  assign _T_61244 = $signed(-4'sh1) * $signed(io_in_367); // @[Modules.scala 144:80:@7268.4]
  assign _T_61245 = $signed(_T_58193) + $signed(_T_61244); // @[Modules.scala 143:103:@7269.4]
  assign _T_61246 = _T_61245[4:0]; // @[Modules.scala 143:103:@7270.4]
  assign _T_61247 = $signed(_T_61246); // @[Modules.scala 143:103:@7271.4]
  assign _GEN_174 = {{1{_T_55179[4]}},_T_55179}; // @[Modules.scala 143:103:@7275.4]
  assign _T_61252 = $signed(_GEN_174) + $signed(_T_58205); // @[Modules.scala 143:103:@7275.4]
  assign _T_61253 = _T_61252[5:0]; // @[Modules.scala 143:103:@7276.4]
  assign _T_61254 = $signed(_T_61253); // @[Modules.scala 143:103:@7277.4]
  assign _T_61258 = $signed(4'sh1) * $signed(io_in_371); // @[Modules.scala 144:80:@7280.4]
  assign _T_61259 = $signed(_T_58207) + $signed(_T_61258); // @[Modules.scala 143:103:@7281.4]
  assign _T_61260 = _T_61259[5:0]; // @[Modules.scala 143:103:@7282.4]
  assign _T_61261 = $signed(_T_61260); // @[Modules.scala 143:103:@7283.4]
  assign _T_61265 = $signed(4'sh1) * $signed(io_in_373); // @[Modules.scala 144:80:@7286.4]
  assign _T_61266 = $signed(_T_58212) + $signed(_T_61265); // @[Modules.scala 143:103:@7287.4]
  assign _T_61267 = _T_61266[5:0]; // @[Modules.scala 143:103:@7288.4]
  assign _T_61268 = $signed(_T_61267); // @[Modules.scala 143:103:@7289.4]
  assign _T_61270 = $signed(4'sh1) * $signed(io_in_374); // @[Modules.scala 143:74:@7291.4]
  assign _T_61272 = $signed(4'sh1) * $signed(io_in_375); // @[Modules.scala 144:80:@7292.4]
  assign _T_61273 = $signed(_T_61270) + $signed(_T_61272); // @[Modules.scala 143:103:@7293.4]
  assign _T_61274 = _T_61273[5:0]; // @[Modules.scala 143:103:@7294.4]
  assign _T_61275 = $signed(_T_61274); // @[Modules.scala 143:103:@7295.4]
  assign _T_61277 = $signed(4'sh1) * $signed(io_in_376); // @[Modules.scala 143:74:@7297.4]
  assign _T_61280 = $signed(_T_61277) + $signed(_T_58226); // @[Modules.scala 143:103:@7299.4]
  assign _T_61281 = _T_61280[5:0]; // @[Modules.scala 143:103:@7300.4]
  assign _T_61282 = $signed(_T_61281); // @[Modules.scala 143:103:@7301.4]
  assign _T_61284 = $signed(-4'sh1) * $signed(io_in_378); // @[Modules.scala 143:74:@7303.4]
  assign _GEN_175 = {{1{_T_61284[4]}},_T_61284}; // @[Modules.scala 143:103:@7305.4]
  assign _T_61287 = $signed(_GEN_175) + $signed(_T_58233); // @[Modules.scala 143:103:@7305.4]
  assign _T_61288 = _T_61287[5:0]; // @[Modules.scala 143:103:@7306.4]
  assign _T_61289 = $signed(_T_61288); // @[Modules.scala 143:103:@7307.4]
  assign _T_61294 = $signed(_T_58235) + $signed(_T_58240); // @[Modules.scala 143:103:@7311.4]
  assign _T_61295 = _T_61294[5:0]; // @[Modules.scala 143:103:@7312.4]
  assign _T_61296 = $signed(_T_61295); // @[Modules.scala 143:103:@7313.4]
  assign _T_61301 = $signed(_T_55221) + $signed(_T_58247); // @[Modules.scala 143:103:@7317.4]
  assign _T_61302 = _T_61301[5:0]; // @[Modules.scala 143:103:@7318.4]
  assign _T_61303 = $signed(_T_61302); // @[Modules.scala 143:103:@7319.4]
  assign _T_61305 = $signed(4'sh1) * $signed(io_in_385); // @[Modules.scala 143:74:@7321.4]
  assign _T_61307 = $signed(4'sh1) * $signed(io_in_386); // @[Modules.scala 144:80:@7322.4]
  assign _T_61308 = $signed(_T_61305) + $signed(_T_61307); // @[Modules.scala 143:103:@7323.4]
  assign _T_61309 = _T_61308[5:0]; // @[Modules.scala 143:103:@7324.4]
  assign _T_61310 = $signed(_T_61309); // @[Modules.scala 143:103:@7325.4]
  assign _T_61315 = $signed(_T_55230) + $signed(_T_55235); // @[Modules.scala 143:103:@7329.4]
  assign _T_61316 = _T_61315[5:0]; // @[Modules.scala 143:103:@7330.4]
  assign _T_61317 = $signed(_T_61316); // @[Modules.scala 143:103:@7331.4]
  assign _T_61322 = $signed(_T_55237) + $signed(_T_55242); // @[Modules.scala 143:103:@7335.4]
  assign _T_61323 = _T_61322[4:0]; // @[Modules.scala 143:103:@7336.4]
  assign _T_61324 = $signed(_T_61323); // @[Modules.scala 143:103:@7337.4]
  assign _T_61326 = $signed(-4'sh1) * $signed(io_in_391); // @[Modules.scala 143:74:@7339.4]
  assign _GEN_176 = {{1{_T_61326[4]}},_T_61326}; // @[Modules.scala 143:103:@7341.4]
  assign _T_61329 = $signed(_GEN_176) + $signed(_T_55249); // @[Modules.scala 143:103:@7341.4]
  assign _T_61330 = _T_61329[5:0]; // @[Modules.scala 143:103:@7342.4]
  assign _T_61331 = $signed(_T_61330); // @[Modules.scala 143:103:@7343.4]
  assign _T_61336 = $signed(_T_58282) + $signed(_T_55256); // @[Modules.scala 143:103:@7347.4]
  assign _T_61337 = _T_61336[5:0]; // @[Modules.scala 143:103:@7348.4]
  assign _T_61338 = $signed(_T_61337); // @[Modules.scala 143:103:@7349.4]
  assign _T_61343 = $signed(_T_55258) + $signed(_T_58289); // @[Modules.scala 143:103:@7353.4]
  assign _T_61344 = _T_61343[5:0]; // @[Modules.scala 143:103:@7354.4]
  assign _T_61345 = $signed(_T_61344); // @[Modules.scala 143:103:@7355.4]
  assign _T_61349 = $signed(4'sh1) * $signed(io_in_398); // @[Modules.scala 144:80:@7358.4]
  assign _T_61350 = $signed(_T_58291) + $signed(_T_61349); // @[Modules.scala 143:103:@7359.4]
  assign _T_61351 = _T_61350[5:0]; // @[Modules.scala 143:103:@7360.4]
  assign _T_61352 = $signed(_T_61351); // @[Modules.scala 143:103:@7361.4]
  assign _T_61354 = $signed(4'sh1) * $signed(io_in_399); // @[Modules.scala 143:74:@7363.4]
  assign _T_61357 = $signed(_T_61354) + $signed(_T_58296); // @[Modules.scala 143:103:@7365.4]
  assign _T_61358 = _T_61357[5:0]; // @[Modules.scala 143:103:@7366.4]
  assign _T_61359 = $signed(_T_61358); // @[Modules.scala 143:103:@7367.4]
  assign _T_61361 = $signed(4'sh1) * $signed(io_in_401); // @[Modules.scala 143:74:@7369.4]
  assign _T_61363 = $signed(4'sh1) * $signed(io_in_402); // @[Modules.scala 144:80:@7370.4]
  assign _T_61364 = $signed(_T_61361) + $signed(_T_61363); // @[Modules.scala 143:103:@7371.4]
  assign _T_61365 = _T_61364[5:0]; // @[Modules.scala 143:103:@7372.4]
  assign _T_61366 = $signed(_T_61365); // @[Modules.scala 143:103:@7373.4]
  assign _T_61368 = $signed(4'sh1) * $signed(io_in_403); // @[Modules.scala 143:74:@7375.4]
  assign _T_61370 = $signed(4'sh1) * $signed(io_in_404); // @[Modules.scala 144:80:@7376.4]
  assign _T_61371 = $signed(_T_61368) + $signed(_T_61370); // @[Modules.scala 143:103:@7377.4]
  assign _T_61372 = _T_61371[5:0]; // @[Modules.scala 143:103:@7378.4]
  assign _T_61373 = $signed(_T_61372); // @[Modules.scala 143:103:@7379.4]
  assign _T_61378 = $signed(_T_58310) + $signed(_T_55298); // @[Modules.scala 143:103:@7383.4]
  assign _T_61379 = _T_61378[5:0]; // @[Modules.scala 143:103:@7384.4]
  assign _T_61380 = $signed(_T_61379); // @[Modules.scala 143:103:@7385.4]
  assign _T_61382 = $signed(4'sh1) * $signed(io_in_408); // @[Modules.scala 143:74:@7387.4]
  assign _T_61384 = $signed(4'sh1) * $signed(io_in_409); // @[Modules.scala 144:80:@7388.4]
  assign _T_61385 = $signed(_T_61382) + $signed(_T_61384); // @[Modules.scala 143:103:@7389.4]
  assign _T_61386 = _T_61385[5:0]; // @[Modules.scala 143:103:@7390.4]
  assign _T_61387 = $signed(_T_61386); // @[Modules.scala 143:103:@7391.4]
  assign _T_61391 = $signed(4'sh1) * $signed(io_in_412); // @[Modules.scala 144:80:@7394.4]
  assign _T_61392 = $signed(_T_55307) + $signed(_T_61391); // @[Modules.scala 143:103:@7395.4]
  assign _T_61393 = _T_61392[5:0]; // @[Modules.scala 143:103:@7396.4]
  assign _T_61394 = $signed(_T_61393); // @[Modules.scala 143:103:@7397.4]
  assign _T_61398 = $signed(4'sh1) * $signed(io_in_414); // @[Modules.scala 144:80:@7400.4]
  assign _T_61399 = $signed(_T_55314) + $signed(_T_61398); // @[Modules.scala 143:103:@7401.4]
  assign _T_61400 = _T_61399[5:0]; // @[Modules.scala 143:103:@7402.4]
  assign _T_61401 = $signed(_T_61400); // @[Modules.scala 143:103:@7403.4]
  assign _T_61403 = $signed(4'sh1) * $signed(io_in_415); // @[Modules.scala 143:74:@7405.4]
  assign _T_61406 = $signed(_T_61403) + $signed(_T_55319); // @[Modules.scala 143:103:@7407.4]
  assign _T_61407 = _T_61406[5:0]; // @[Modules.scala 143:103:@7408.4]
  assign _T_61408 = $signed(_T_61407); // @[Modules.scala 143:103:@7409.4]
  assign _T_61412 = $signed(-4'sh1) * $signed(io_in_419); // @[Modules.scala 144:80:@7412.4]
  assign _T_61413 = $signed(_T_58347) + $signed(_T_61412); // @[Modules.scala 143:103:@7413.4]
  assign _T_61414 = _T_61413[4:0]; // @[Modules.scala 143:103:@7414.4]
  assign _T_61415 = $signed(_T_61414); // @[Modules.scala 143:103:@7415.4]
  assign _T_61419 = $signed(4'sh1) * $signed(io_in_421); // @[Modules.scala 144:80:@7418.4]
  assign _T_61420 = $signed(_T_55328) + $signed(_T_61419); // @[Modules.scala 143:103:@7419.4]
  assign _T_61421 = _T_61420[5:0]; // @[Modules.scala 143:103:@7420.4]
  assign _T_61422 = $signed(_T_61421); // @[Modules.scala 143:103:@7421.4]
  assign _T_61427 = $signed(_T_55335) + $signed(_T_55340); // @[Modules.scala 143:103:@7425.4]
  assign _T_61428 = _T_61427[5:0]; // @[Modules.scala 143:103:@7426.4]
  assign _T_61429 = $signed(_T_61428); // @[Modules.scala 143:103:@7427.4]
  assign _T_61431 = $signed(4'sh1) * $signed(io_in_425); // @[Modules.scala 143:74:@7429.4]
  assign _T_61433 = $signed(4'sh1) * $signed(io_in_426); // @[Modules.scala 144:80:@7430.4]
  assign _T_61434 = $signed(_T_61431) + $signed(_T_61433); // @[Modules.scala 143:103:@7431.4]
  assign _T_61435 = _T_61434[5:0]; // @[Modules.scala 143:103:@7432.4]
  assign _T_61436 = $signed(_T_61435); // @[Modules.scala 143:103:@7433.4]
  assign _T_61438 = $signed(4'sh1) * $signed(io_in_427); // @[Modules.scala 143:74:@7435.4]
  assign _T_61440 = $signed(4'sh1) * $signed(io_in_429); // @[Modules.scala 144:80:@7436.4]
  assign _T_61441 = $signed(_T_61438) + $signed(_T_61440); // @[Modules.scala 143:103:@7437.4]
  assign _T_61442 = _T_61441[5:0]; // @[Modules.scala 143:103:@7438.4]
  assign _T_61443 = $signed(_T_61442); // @[Modules.scala 143:103:@7439.4]
  assign _T_61445 = $signed(4'sh1) * $signed(io_in_430); // @[Modules.scala 143:74:@7441.4]
  assign _T_61447 = $signed(4'sh1) * $signed(io_in_431); // @[Modules.scala 144:80:@7442.4]
  assign _T_61448 = $signed(_T_61445) + $signed(_T_61447); // @[Modules.scala 143:103:@7443.4]
  assign _T_61449 = _T_61448[5:0]; // @[Modules.scala 143:103:@7444.4]
  assign _T_61450 = $signed(_T_61449); // @[Modules.scala 143:103:@7445.4]
  assign _T_61454 = $signed(-4'sh1) * $signed(io_in_433); // @[Modules.scala 144:80:@7448.4]
  assign _GEN_177 = {{1{_T_61454[4]}},_T_61454}; // @[Modules.scala 143:103:@7449.4]
  assign _T_61455 = $signed(_T_55363) + $signed(_GEN_177); // @[Modules.scala 143:103:@7449.4]
  assign _T_61456 = _T_61455[5:0]; // @[Modules.scala 143:103:@7450.4]
  assign _T_61457 = $signed(_T_61456); // @[Modules.scala 143:103:@7451.4]
  assign _T_61462 = $signed(_T_55370) + $signed(_T_55375); // @[Modules.scala 143:103:@7455.4]
  assign _T_61463 = _T_61462[5:0]; // @[Modules.scala 143:103:@7456.4]
  assign _T_61464 = $signed(_T_61463); // @[Modules.scala 143:103:@7457.4]
  assign _T_61466 = $signed(4'sh1) * $signed(io_in_436); // @[Modules.scala 143:74:@7459.4]
  assign _T_61468 = $signed(4'sh1) * $signed(io_in_437); // @[Modules.scala 144:80:@7460.4]
  assign _T_61469 = $signed(_T_61466) + $signed(_T_61468); // @[Modules.scala 143:103:@7461.4]
  assign _T_61470 = _T_61469[5:0]; // @[Modules.scala 143:103:@7462.4]
  assign _T_61471 = $signed(_T_61470); // @[Modules.scala 143:103:@7463.4]
  assign _T_61473 = $signed(-4'sh1) * $signed(io_in_438); // @[Modules.scala 143:74:@7465.4]
  assign _T_61475 = $signed(-4'sh1) * $signed(io_in_439); // @[Modules.scala 144:80:@7466.4]
  assign _T_61476 = $signed(_T_61473) + $signed(_T_61475); // @[Modules.scala 143:103:@7467.4]
  assign _T_61477 = _T_61476[4:0]; // @[Modules.scala 143:103:@7468.4]
  assign _T_61478 = $signed(_T_61477); // @[Modules.scala 143:103:@7469.4]
  assign _T_61483 = $signed(_T_55391) + $signed(_T_58403); // @[Modules.scala 143:103:@7473.4]
  assign _T_61484 = _T_61483[5:0]; // @[Modules.scala 143:103:@7474.4]
  assign _T_61485 = $signed(_T_61484); // @[Modules.scala 143:103:@7475.4]
  assign _T_61489 = $signed(4'sh1) * $signed(io_in_444); // @[Modules.scala 144:80:@7478.4]
  assign _T_61490 = $signed(_GEN_49) + $signed(_T_61489); // @[Modules.scala 143:103:@7479.4]
  assign _T_61491 = _T_61490[5:0]; // @[Modules.scala 143:103:@7480.4]
  assign _T_61492 = $signed(_T_61491); // @[Modules.scala 143:103:@7481.4]
  assign _T_61496 = $signed(-4'sh1) * $signed(io_in_447); // @[Modules.scala 144:80:@7484.4]
  assign _T_61497 = $signed(_T_58417) + $signed(_T_61496); // @[Modules.scala 143:103:@7485.4]
  assign _T_61498 = _T_61497[4:0]; // @[Modules.scala 143:103:@7486.4]
  assign _T_61499 = $signed(_T_61498); // @[Modules.scala 143:103:@7487.4]
  assign _T_61503 = $signed(4'sh1) * $signed(io_in_449); // @[Modules.scala 144:80:@7490.4]
  assign _GEN_179 = {{1{_T_55417[4]}},_T_55417}; // @[Modules.scala 143:103:@7491.4]
  assign _T_61504 = $signed(_GEN_179) + $signed(_T_61503); // @[Modules.scala 143:103:@7491.4]
  assign _T_61505 = _T_61504[5:0]; // @[Modules.scala 143:103:@7492.4]
  assign _T_61506 = $signed(_T_61505); // @[Modules.scala 143:103:@7493.4]
  assign _T_61510 = $signed(-4'sh1) * $signed(io_in_451); // @[Modules.scala 144:80:@7496.4]
  assign _GEN_180 = {{1{_T_61510[4]}},_T_61510}; // @[Modules.scala 143:103:@7497.4]
  assign _T_61511 = $signed(_T_55424) + $signed(_GEN_180); // @[Modules.scala 143:103:@7497.4]
  assign _T_61512 = _T_61511[5:0]; // @[Modules.scala 143:103:@7498.4]
  assign _T_61513 = $signed(_T_61512); // @[Modules.scala 143:103:@7499.4]
  assign _T_61522 = $signed(4'sh1) * $signed(io_in_454); // @[Modules.scala 143:74:@7507.4]
  assign _T_61525 = $signed(_T_61522) + $signed(_T_55438); // @[Modules.scala 143:103:@7509.4]
  assign _T_61526 = _T_61525[5:0]; // @[Modules.scala 143:103:@7510.4]
  assign _T_61527 = $signed(_T_61526); // @[Modules.scala 143:103:@7511.4]
  assign _GEN_181 = {{1{_T_58466[4]}},_T_58466}; // @[Modules.scala 143:103:@7515.4]
  assign _T_61532 = $signed(_T_55447) + $signed(_GEN_181); // @[Modules.scala 143:103:@7515.4]
  assign _T_61533 = _T_61532[5:0]; // @[Modules.scala 143:103:@7516.4]
  assign _T_61534 = $signed(_T_61533); // @[Modules.scala 143:103:@7517.4]
  assign _T_61536 = $signed(-4'sh1) * $signed(io_in_461); // @[Modules.scala 143:74:@7519.4]
  assign _GEN_182 = {{1{_T_61536[4]}},_T_61536}; // @[Modules.scala 143:103:@7521.4]
  assign _T_61539 = $signed(_GEN_182) + $signed(_T_55454); // @[Modules.scala 143:103:@7521.4]
  assign _T_61540 = _T_61539[5:0]; // @[Modules.scala 143:103:@7522.4]
  assign _T_61541 = $signed(_T_61540); // @[Modules.scala 143:103:@7523.4]
  assign _T_61545 = $signed(4'sh1) * $signed(io_in_464); // @[Modules.scala 144:80:@7526.4]
  assign _T_61546 = $signed(_T_55459) + $signed(_T_61545); // @[Modules.scala 143:103:@7527.4]
  assign _T_61547 = _T_61546[5:0]; // @[Modules.scala 143:103:@7528.4]
  assign _T_61548 = $signed(_T_61547); // @[Modules.scala 143:103:@7529.4]
  assign _T_61552 = $signed(-4'sh1) * $signed(io_in_467); // @[Modules.scala 144:80:@7532.4]
  assign _GEN_183 = {{1{_T_61552[4]}},_T_61552}; // @[Modules.scala 143:103:@7533.4]
  assign _T_61553 = $signed(_T_58478) + $signed(_GEN_183); // @[Modules.scala 143:103:@7533.4]
  assign _T_61554 = _T_61553[5:0]; // @[Modules.scala 143:103:@7534.4]
  assign _T_61555 = $signed(_T_61554); // @[Modules.scala 143:103:@7535.4]
  assign _T_61557 = $signed(4'sh1) * $signed(io_in_468); // @[Modules.scala 143:74:@7537.4]
  assign _T_61560 = $signed(_T_61557) + $signed(_T_55473); // @[Modules.scala 143:103:@7539.4]
  assign _T_61561 = _T_61560[5:0]; // @[Modules.scala 143:103:@7540.4]
  assign _T_61562 = $signed(_T_61561); // @[Modules.scala 143:103:@7541.4]
  assign _T_61564 = $signed(-4'sh1) * $signed(io_in_470); // @[Modules.scala 143:74:@7543.4]
  assign _T_61567 = $signed(_T_61564) + $signed(_T_55475); // @[Modules.scala 143:103:@7545.4]
  assign _T_61568 = _T_61567[4:0]; // @[Modules.scala 143:103:@7546.4]
  assign _T_61569 = $signed(_T_61568); // @[Modules.scala 143:103:@7547.4]
  assign _T_61573 = $signed(-4'sh1) * $signed(io_in_474); // @[Modules.scala 144:80:@7550.4]
  assign _T_61574 = $signed(_T_58492) + $signed(_T_61573); // @[Modules.scala 143:103:@7551.4]
  assign _T_61575 = _T_61574[4:0]; // @[Modules.scala 143:103:@7552.4]
  assign _T_61576 = $signed(_T_61575); // @[Modules.scala 143:103:@7553.4]
  assign _T_61578 = $signed(-4'sh1) * $signed(io_in_475); // @[Modules.scala 143:74:@7555.4]
  assign _T_61580 = $signed(4'sh1) * $signed(io_in_477); // @[Modules.scala 144:80:@7556.4]
  assign _GEN_184 = {{1{_T_61578[4]}},_T_61578}; // @[Modules.scala 143:103:@7557.4]
  assign _T_61581 = $signed(_GEN_184) + $signed(_T_61580); // @[Modules.scala 143:103:@7557.4]
  assign _T_61582 = _T_61581[5:0]; // @[Modules.scala 143:103:@7558.4]
  assign _T_61583 = $signed(_T_61582); // @[Modules.scala 143:103:@7559.4]
  assign _T_61585 = $signed(-4'sh1) * $signed(io_in_478); // @[Modules.scala 143:74:@7561.4]
  assign _T_61587 = $signed(-4'sh1) * $signed(io_in_479); // @[Modules.scala 144:80:@7562.4]
  assign _T_61588 = $signed(_T_61585) + $signed(_T_61587); // @[Modules.scala 143:103:@7563.4]
  assign _T_61589 = _T_61588[4:0]; // @[Modules.scala 143:103:@7564.4]
  assign _T_61590 = $signed(_T_61589); // @[Modules.scala 143:103:@7565.4]
  assign _T_61592 = $signed(-4'sh1) * $signed(io_in_480); // @[Modules.scala 143:74:@7567.4]
  assign _T_61595 = $signed(_T_61592) + $signed(_T_58520); // @[Modules.scala 143:103:@7569.4]
  assign _T_61596 = _T_61595[4:0]; // @[Modules.scala 143:103:@7570.4]
  assign _T_61597 = $signed(_T_61596); // @[Modules.scala 143:103:@7571.4]
  assign _T_61601 = $signed(4'sh1) * $signed(io_in_483); // @[Modules.scala 144:80:@7574.4]
  assign _GEN_185 = {{1{_T_58522[4]}},_T_58522}; // @[Modules.scala 143:103:@7575.4]
  assign _T_61602 = $signed(_GEN_185) + $signed(_T_61601); // @[Modules.scala 143:103:@7575.4]
  assign _T_61603 = _T_61602[5:0]; // @[Modules.scala 143:103:@7576.4]
  assign _T_61604 = $signed(_T_61603); // @[Modules.scala 143:103:@7577.4]
  assign _T_61606 = $signed(4'sh1) * $signed(io_in_484); // @[Modules.scala 143:74:@7579.4]
  assign _T_61609 = $signed(_T_61606) + $signed(_T_55508); // @[Modules.scala 143:103:@7581.4]
  assign _T_61610 = _T_61609[5:0]; // @[Modules.scala 143:103:@7582.4]
  assign _T_61611 = $signed(_T_61610); // @[Modules.scala 143:103:@7583.4]
  assign _T_61616 = $signed(_T_55517) + $signed(_T_55522); // @[Modules.scala 143:103:@7587.4]
  assign _T_61617 = _T_61616[5:0]; // @[Modules.scala 143:103:@7588.4]
  assign _T_61618 = $signed(_T_61617); // @[Modules.scala 143:103:@7589.4]
  assign _T_61622 = $signed(4'sh1) * $signed(io_in_492); // @[Modules.scala 144:80:@7592.4]
  assign _T_61623 = $signed(_T_55524) + $signed(_T_61622); // @[Modules.scala 143:103:@7593.4]
  assign _T_61624 = _T_61623[5:0]; // @[Modules.scala 143:103:@7594.4]
  assign _T_61625 = $signed(_T_61624); // @[Modules.scala 143:103:@7595.4]
  assign _T_61629 = $signed(-4'sh1) * $signed(io_in_498); // @[Modules.scala 144:80:@7598.4]
  assign _GEN_186 = {{1{_T_61629[4]}},_T_61629}; // @[Modules.scala 143:103:@7599.4]
  assign _T_61630 = $signed(_T_58557) + $signed(_GEN_186); // @[Modules.scala 143:103:@7599.4]
  assign _T_61631 = _T_61630[5:0]; // @[Modules.scala 143:103:@7600.4]
  assign _T_61632 = $signed(_T_61631); // @[Modules.scala 143:103:@7601.4]
  assign _T_61637 = $signed(_T_58571) + $signed(_T_58576); // @[Modules.scala 143:103:@7605.4]
  assign _T_61638 = _T_61637[4:0]; // @[Modules.scala 143:103:@7606.4]
  assign _T_61639 = $signed(_T_61638); // @[Modules.scala 143:103:@7607.4]
  assign _T_61643 = $signed(-4'sh1) * $signed(io_in_503); // @[Modules.scala 144:80:@7610.4]
  assign _T_61644 = $signed(_T_58578) + $signed(_T_61643); // @[Modules.scala 143:103:@7611.4]
  assign _T_61645 = _T_61644[4:0]; // @[Modules.scala 143:103:@7612.4]
  assign _T_61646 = $signed(_T_61645); // @[Modules.scala 143:103:@7613.4]
  assign _T_61651 = $signed(_GEN_56) + $signed(_T_55564); // @[Modules.scala 143:103:@7617.4]
  assign _T_61652 = _T_61651[5:0]; // @[Modules.scala 143:103:@7618.4]
  assign _T_61653 = $signed(_T_61652); // @[Modules.scala 143:103:@7619.4]
  assign _T_61657 = $signed(-4'sh1) * $signed(io_in_507); // @[Modules.scala 144:80:@7622.4]
  assign _GEN_188 = {{1{_T_61657[4]}},_T_61657}; // @[Modules.scala 143:103:@7623.4]
  assign _T_61658 = $signed(_T_55566) + $signed(_GEN_188); // @[Modules.scala 143:103:@7623.4]
  assign _T_61659 = _T_61658[5:0]; // @[Modules.scala 143:103:@7624.4]
  assign _T_61660 = $signed(_T_61659); // @[Modules.scala 143:103:@7625.4]
  assign _T_61662 = $signed(-4'sh1) * $signed(io_in_508); // @[Modules.scala 143:74:@7627.4]
  assign _T_61665 = $signed(_T_61662) + $signed(_T_58599); // @[Modules.scala 143:103:@7629.4]
  assign _T_61666 = _T_61665[4:0]; // @[Modules.scala 143:103:@7630.4]
  assign _T_61667 = $signed(_T_61666); // @[Modules.scala 143:103:@7631.4]
  assign _T_61676 = $signed(4'sh1) * $signed(io_in_512); // @[Modules.scala 143:74:@7639.4]
  assign _T_61679 = $signed(_T_61676) + $signed(_T_55587); // @[Modules.scala 143:103:@7641.4]
  assign _T_61680 = _T_61679[5:0]; // @[Modules.scala 143:103:@7642.4]
  assign _T_61681 = $signed(_T_61680); // @[Modules.scala 143:103:@7643.4]
  assign _T_61699 = $signed(-4'sh1) * $signed(io_in_521); // @[Modules.scala 144:80:@7658.4]
  assign _GEN_189 = {{1{_T_61699[4]}},_T_61699}; // @[Modules.scala 143:103:@7659.4]
  assign _T_61700 = $signed(_T_55606) + $signed(_GEN_189); // @[Modules.scala 143:103:@7659.4]
  assign _T_61701 = _T_61700[5:0]; // @[Modules.scala 143:103:@7660.4]
  assign _T_61702 = $signed(_T_61701); // @[Modules.scala 143:103:@7661.4]
  assign _T_61706 = $signed(-4'sh1) * $signed(io_in_526); // @[Modules.scala 144:80:@7664.4]
  assign _GEN_190 = {{1{_T_61706[4]}},_T_61706}; // @[Modules.scala 143:103:@7665.4]
  assign _T_61707 = $signed(_T_55622) + $signed(_GEN_190); // @[Modules.scala 143:103:@7665.4]
  assign _T_61708 = _T_61707[5:0]; // @[Modules.scala 143:103:@7666.4]
  assign _T_61709 = $signed(_T_61708); // @[Modules.scala 143:103:@7667.4]
  assign _T_61725 = $signed(-4'sh1) * $signed(io_in_531); // @[Modules.scala 143:74:@7681.4]
  assign _GEN_191 = {{1{_T_61725[4]}},_T_61725}; // @[Modules.scala 143:103:@7683.4]
  assign _T_61728 = $signed(_GEN_191) + $signed(_T_58655); // @[Modules.scala 143:103:@7683.4]
  assign _T_61729 = _T_61728[5:0]; // @[Modules.scala 143:103:@7684.4]
  assign _T_61730 = $signed(_T_61729); // @[Modules.scala 143:103:@7685.4]
  assign _T_61735 = $signed(_T_55650) + $signed(_T_55655); // @[Modules.scala 143:103:@7689.4]
  assign _T_61736 = _T_61735[5:0]; // @[Modules.scala 143:103:@7690.4]
  assign _T_61737 = $signed(_T_61736); // @[Modules.scala 143:103:@7691.4]
  assign _T_61739 = $signed(-4'sh1) * $signed(io_in_535); // @[Modules.scala 143:74:@7693.4]
  assign _T_61741 = $signed(-4'sh1) * $signed(io_in_536); // @[Modules.scala 144:80:@7694.4]
  assign _T_61742 = $signed(_T_61739) + $signed(_T_61741); // @[Modules.scala 143:103:@7695.4]
  assign _T_61743 = _T_61742[4:0]; // @[Modules.scala 143:103:@7696.4]
  assign _T_61744 = $signed(_T_61743); // @[Modules.scala 143:103:@7697.4]
  assign _T_61753 = $signed(-4'sh1) * $signed(io_in_539); // @[Modules.scala 143:74:@7705.4]
  assign _T_61756 = $signed(_T_61753) + $signed(_T_58681); // @[Modules.scala 143:103:@7707.4]
  assign _T_61757 = _T_61756[4:0]; // @[Modules.scala 143:103:@7708.4]
  assign _T_61758 = $signed(_T_61757); // @[Modules.scala 143:103:@7709.4]
  assign _GEN_192 = {{1{_T_58683[4]}},_T_58683}; // @[Modules.scala 143:103:@7713.4]
  assign _T_61763 = $signed(_GEN_192) + $signed(_T_55683); // @[Modules.scala 143:103:@7713.4]
  assign _T_61764 = _T_61763[5:0]; // @[Modules.scala 143:103:@7714.4]
  assign _T_61765 = $signed(_T_61764); // @[Modules.scala 143:103:@7715.4]
  assign _GEN_193 = {{1{_T_58697[4]}},_T_58697}; // @[Modules.scala 143:103:@7719.4]
  assign _T_61770 = $signed(_T_55685) + $signed(_GEN_193); // @[Modules.scala 143:103:@7719.4]
  assign _T_61771 = _T_61770[5:0]; // @[Modules.scala 143:103:@7720.4]
  assign _T_61772 = $signed(_T_61771); // @[Modules.scala 143:103:@7721.4]
  assign _T_61774 = $signed(-4'sh1) * $signed(io_in_546); // @[Modules.scala 143:74:@7723.4]
  assign _GEN_194 = {{1{_T_61774[4]}},_T_61774}; // @[Modules.scala 143:103:@7725.4]
  assign _T_61777 = $signed(_GEN_194) + $signed(_T_55697); // @[Modules.scala 143:103:@7725.4]
  assign _T_61778 = _T_61777[5:0]; // @[Modules.scala 143:103:@7726.4]
  assign _T_61779 = $signed(_T_61778); // @[Modules.scala 143:103:@7727.4]
  assign _GEN_195 = {{1{_T_58711[4]}},_T_58711}; // @[Modules.scala 143:103:@7731.4]
  assign _T_61784 = $signed(_T_55699) + $signed(_GEN_195); // @[Modules.scala 143:103:@7731.4]
  assign _T_61785 = _T_61784[5:0]; // @[Modules.scala 143:103:@7732.4]
  assign _T_61786 = $signed(_T_61785); // @[Modules.scala 143:103:@7733.4]
  assign _T_61809 = $signed(4'sh1) * $signed(io_in_561); // @[Modules.scala 143:74:@7753.4]
  assign _T_61812 = $signed(_T_61809) + $signed(_T_55727); // @[Modules.scala 143:103:@7755.4]
  assign _T_61813 = _T_61812[5:0]; // @[Modules.scala 143:103:@7756.4]
  assign _T_61814 = $signed(_T_61813); // @[Modules.scala 143:103:@7757.4]
  assign _T_61816 = $signed(-4'sh1) * $signed(io_in_563); // @[Modules.scala 143:74:@7759.4]
  assign _T_61818 = $signed(-4'sh1) * $signed(io_in_564); // @[Modules.scala 144:80:@7760.4]
  assign _T_61819 = $signed(_T_61816) + $signed(_T_61818); // @[Modules.scala 143:103:@7761.4]
  assign _T_61820 = _T_61819[4:0]; // @[Modules.scala 143:103:@7762.4]
  assign _T_61821 = $signed(_T_61820); // @[Modules.scala 143:103:@7763.4]
  assign _T_61826 = $signed(_T_58753) + $signed(_T_58758); // @[Modules.scala 143:103:@7767.4]
  assign _T_61827 = _T_61826[4:0]; // @[Modules.scala 143:103:@7768.4]
  assign _T_61828 = $signed(_T_61827); // @[Modules.scala 143:103:@7769.4]
  assign _T_61830 = $signed(-4'sh1) * $signed(io_in_567); // @[Modules.scala 143:74:@7771.4]
  assign _T_61832 = $signed(-4'sh1) * $signed(io_in_568); // @[Modules.scala 144:80:@7772.4]
  assign _T_61833 = $signed(_T_61830) + $signed(_T_61832); // @[Modules.scala 143:103:@7773.4]
  assign _T_61834 = _T_61833[4:0]; // @[Modules.scala 143:103:@7774.4]
  assign _T_61835 = $signed(_T_61834); // @[Modules.scala 143:103:@7775.4]
  assign _T_61837 = $signed(-4'sh1) * $signed(io_in_569); // @[Modules.scala 143:74:@7777.4]
  assign _T_61839 = $signed(-4'sh1) * $signed(io_in_570); // @[Modules.scala 144:80:@7778.4]
  assign _T_61840 = $signed(_T_61837) + $signed(_T_61839); // @[Modules.scala 143:103:@7779.4]
  assign _T_61841 = _T_61840[4:0]; // @[Modules.scala 143:103:@7780.4]
  assign _T_61842 = $signed(_T_61841); // @[Modules.scala 143:103:@7781.4]
  assign _T_61846 = $signed(4'sh1) * $signed(io_in_575); // @[Modules.scala 144:80:@7784.4]
  assign _T_61847 = $signed(_T_55762) + $signed(_T_61846); // @[Modules.scala 143:103:@7785.4]
  assign _T_61848 = _T_61847[5:0]; // @[Modules.scala 143:103:@7786.4]
  assign _T_61849 = $signed(_T_61848); // @[Modules.scala 143:103:@7787.4]
  assign _T_61851 = $signed(4'sh1) * $signed(io_in_576); // @[Modules.scala 143:74:@7789.4]
  assign _GEN_196 = {{1{_T_58781[4]}},_T_58781}; // @[Modules.scala 143:103:@7791.4]
  assign _T_61854 = $signed(_T_61851) + $signed(_GEN_196); // @[Modules.scala 143:103:@7791.4]
  assign _T_61855 = _T_61854[5:0]; // @[Modules.scala 143:103:@7792.4]
  assign _T_61856 = $signed(_T_61855); // @[Modules.scala 143:103:@7793.4]
  assign _T_61858 = $signed(-4'sh1) * $signed(io_in_579); // @[Modules.scala 143:74:@7795.4]
  assign _T_61861 = $signed(_T_61858) + $signed(_T_58793); // @[Modules.scala 143:103:@7797.4]
  assign _T_61862 = _T_61861[4:0]; // @[Modules.scala 143:103:@7798.4]
  assign _T_61863 = $signed(_T_61862); // @[Modules.scala 143:103:@7799.4]
  assign _T_61868 = $signed(_T_55774) + $signed(_T_58800); // @[Modules.scala 143:103:@7803.4]
  assign _T_61869 = _T_61868[4:0]; // @[Modules.scala 143:103:@7804.4]
  assign _T_61870 = $signed(_T_61869); // @[Modules.scala 143:103:@7805.4]
  assign _GEN_197 = {{1{_T_58802[4]}},_T_58802}; // @[Modules.scala 143:103:@7809.4]
  assign _T_61875 = $signed(_GEN_197) + $signed(_T_55783); // @[Modules.scala 143:103:@7809.4]
  assign _T_61876 = _T_61875[5:0]; // @[Modules.scala 143:103:@7810.4]
  assign _T_61877 = $signed(_T_61876); // @[Modules.scala 143:103:@7811.4]
  assign _T_61879 = $signed(-4'sh1) * $signed(io_in_586); // @[Modules.scala 143:74:@7813.4]
  assign _GEN_198 = {{1{_T_61879[4]}},_T_61879}; // @[Modules.scala 143:103:@7815.4]
  assign _T_61882 = $signed(_GEN_198) + $signed(_T_55788); // @[Modules.scala 143:103:@7815.4]
  assign _T_61883 = _T_61882[5:0]; // @[Modules.scala 143:103:@7816.4]
  assign _T_61884 = $signed(_T_61883); // @[Modules.scala 143:103:@7817.4]
  assign _T_61889 = $signed(_T_55790) + $signed(_T_55795); // @[Modules.scala 143:103:@7821.4]
  assign _T_61890 = _T_61889[5:0]; // @[Modules.scala 143:103:@7822.4]
  assign _T_61891 = $signed(_T_61890); // @[Modules.scala 143:103:@7823.4]
  assign _T_61895 = $signed(-4'sh1) * $signed(io_in_591); // @[Modules.scala 144:80:@7826.4]
  assign _GEN_199 = {{1{_T_61895[4]}},_T_61895}; // @[Modules.scala 143:103:@7827.4]
  assign _T_61896 = $signed(_T_55797) + $signed(_GEN_199); // @[Modules.scala 143:103:@7827.4]
  assign _T_61897 = _T_61896[5:0]; // @[Modules.scala 143:103:@7828.4]
  assign _T_61898 = $signed(_T_61897); // @[Modules.scala 143:103:@7829.4]
  assign _T_61900 = $signed(-4'sh1) * $signed(io_in_592); // @[Modules.scala 143:74:@7831.4]
  assign _T_61902 = $signed(-4'sh1) * $signed(io_in_593); // @[Modules.scala 144:80:@7832.4]
  assign _T_61903 = $signed(_T_61900) + $signed(_T_61902); // @[Modules.scala 143:103:@7833.4]
  assign _T_61904 = _T_61903[4:0]; // @[Modules.scala 143:103:@7834.4]
  assign _T_61905 = $signed(_T_61904); // @[Modules.scala 143:103:@7835.4]
  assign _T_61907 = $signed(-4'sh1) * $signed(io_in_594); // @[Modules.scala 143:74:@7837.4]
  assign _T_61910 = $signed(_T_61907) + $signed(_T_58837); // @[Modules.scala 143:103:@7839.4]
  assign _T_61911 = _T_61910[4:0]; // @[Modules.scala 143:103:@7840.4]
  assign _T_61912 = $signed(_T_61911); // @[Modules.scala 143:103:@7841.4]
  assign _T_61914 = $signed(-4'sh1) * $signed(io_in_596); // @[Modules.scala 143:74:@7843.4]
  assign _T_61916 = $signed(-4'sh1) * $signed(io_in_597); // @[Modules.scala 144:80:@7844.4]
  assign _T_61917 = $signed(_T_61914) + $signed(_T_61916); // @[Modules.scala 143:103:@7845.4]
  assign _T_61918 = _T_61917[4:0]; // @[Modules.scala 143:103:@7846.4]
  assign _T_61919 = $signed(_T_61918); // @[Modules.scala 143:103:@7847.4]
  assign _T_61921 = $signed(-4'sh1) * $signed(io_in_598); // @[Modules.scala 143:74:@7849.4]
  assign _T_61923 = $signed(4'sh1) * $signed(io_in_600); // @[Modules.scala 144:80:@7850.4]
  assign _GEN_200 = {{1{_T_61921[4]}},_T_61921}; // @[Modules.scala 143:103:@7851.4]
  assign _T_61924 = $signed(_GEN_200) + $signed(_T_61923); // @[Modules.scala 143:103:@7851.4]
  assign _T_61925 = _T_61924[5:0]; // @[Modules.scala 143:103:@7852.4]
  assign _T_61926 = $signed(_T_61925); // @[Modules.scala 143:103:@7853.4]
  assign _T_61931 = $signed(_T_55825) + $signed(_T_55830); // @[Modules.scala 143:103:@7857.4]
  assign _T_61932 = _T_61931[5:0]; // @[Modules.scala 143:103:@7858.4]
  assign _T_61933 = $signed(_T_61932); // @[Modules.scala 143:103:@7859.4]
  assign _T_61937 = $signed(4'sh1) * $signed(io_in_605); // @[Modules.scala 144:80:@7862.4]
  assign _T_61938 = $signed(_T_55832) + $signed(_T_61937); // @[Modules.scala 143:103:@7863.4]
  assign _T_61939 = _T_61938[5:0]; // @[Modules.scala 143:103:@7864.4]
  assign _T_61940 = $signed(_T_61939); // @[Modules.scala 143:103:@7865.4]
  assign _T_61944 = $signed(-4'sh1) * $signed(io_in_607); // @[Modules.scala 144:80:@7868.4]
  assign _T_61945 = $signed(_T_58856) + $signed(_T_61944); // @[Modules.scala 143:103:@7869.4]
  assign _T_61946 = _T_61945[4:0]; // @[Modules.scala 143:103:@7870.4]
  assign _T_61947 = $signed(_T_61946); // @[Modules.scala 143:103:@7871.4]
  assign _GEN_201 = {{1{_T_58877[4]}},_T_58877}; // @[Modules.scala 143:103:@7881.4]
  assign _T_61959 = $signed(_T_55844) + $signed(_GEN_201); // @[Modules.scala 143:103:@7881.4]
  assign _T_61960 = _T_61959[5:0]; // @[Modules.scala 143:103:@7882.4]
  assign _T_61961 = $signed(_T_61960); // @[Modules.scala 143:103:@7883.4]
  assign _GEN_202 = {{1{_T_58879[4]}},_T_58879}; // @[Modules.scala 143:103:@7887.4]
  assign _T_61966 = $signed(_GEN_202) + $signed(_T_55858); // @[Modules.scala 143:103:@7887.4]
  assign _T_61967 = _T_61966[5:0]; // @[Modules.scala 143:103:@7888.4]
  assign _T_61968 = $signed(_T_61967); // @[Modules.scala 143:103:@7889.4]
  assign _T_61973 = $signed(_T_55860) + $signed(_T_55865); // @[Modules.scala 143:103:@7893.4]
  assign _T_61974 = _T_61973[5:0]; // @[Modules.scala 143:103:@7894.4]
  assign _T_61975 = $signed(_T_61974); // @[Modules.scala 143:103:@7895.4]
  assign _T_61979 = $signed(-4'sh1) * $signed(io_in_619); // @[Modules.scala 144:80:@7898.4]
  assign _GEN_203 = {{1{_T_61979[4]}},_T_61979}; // @[Modules.scala 143:103:@7899.4]
  assign _T_61980 = $signed(_T_55867) + $signed(_GEN_203); // @[Modules.scala 143:103:@7899.4]
  assign _T_61981 = _T_61980[5:0]; // @[Modules.scala 143:103:@7900.4]
  assign _T_61982 = $signed(_T_61981); // @[Modules.scala 143:103:@7901.4]
  assign _T_61984 = $signed(-4'sh1) * $signed(io_in_620); // @[Modules.scala 143:74:@7903.4]
  assign _T_61986 = $signed(-4'sh1) * $signed(io_in_621); // @[Modules.scala 144:80:@7904.4]
  assign _T_61987 = $signed(_T_61984) + $signed(_T_61986); // @[Modules.scala 143:103:@7905.4]
  assign _T_61988 = _T_61987[4:0]; // @[Modules.scala 143:103:@7906.4]
  assign _T_61989 = $signed(_T_61988); // @[Modules.scala 143:103:@7907.4]
  assign _T_61991 = $signed(-4'sh1) * $signed(io_in_622); // @[Modules.scala 143:74:@7909.4]
  assign _T_61994 = $signed(_T_61991) + $signed(_T_55886); // @[Modules.scala 143:103:@7911.4]
  assign _T_61995 = _T_61994[4:0]; // @[Modules.scala 143:103:@7912.4]
  assign _T_61996 = $signed(_T_61995); // @[Modules.scala 143:103:@7913.4]
  assign _T_61998 = $signed(-4'sh1) * $signed(io_in_624); // @[Modules.scala 143:74:@7915.4]
  assign _T_62000 = $signed(-4'sh1) * $signed(io_in_625); // @[Modules.scala 144:80:@7916.4]
  assign _T_62001 = $signed(_T_61998) + $signed(_T_62000); // @[Modules.scala 143:103:@7917.4]
  assign _T_62002 = _T_62001[4:0]; // @[Modules.scala 143:103:@7918.4]
  assign _T_62003 = $signed(_T_62002); // @[Modules.scala 143:103:@7919.4]
  assign _T_62005 = $signed(-4'sh1) * $signed(io_in_626); // @[Modules.scala 143:74:@7921.4]
  assign _T_62008 = $signed(_T_62005) + $signed(_T_55893); // @[Modules.scala 143:103:@7923.4]
  assign _T_62009 = _T_62008[4:0]; // @[Modules.scala 143:103:@7924.4]
  assign _T_62010 = $signed(_T_62009); // @[Modules.scala 143:103:@7925.4]
  assign _T_62015 = $signed(_T_55902) + $signed(_T_55907); // @[Modules.scala 143:103:@7929.4]
  assign _T_62016 = _T_62015[4:0]; // @[Modules.scala 143:103:@7930.4]
  assign _T_62017 = $signed(_T_62016); // @[Modules.scala 143:103:@7931.4]
  assign _T_62022 = $signed(_T_55909) + $signed(_T_55914); // @[Modules.scala 143:103:@7935.4]
  assign _T_62023 = _T_62022[4:0]; // @[Modules.scala 143:103:@7936.4]
  assign _T_62024 = $signed(_T_62023); // @[Modules.scala 143:103:@7937.4]
  assign _T_62026 = $signed(4'sh1) * $signed(io_in_634); // @[Modules.scala 143:74:@7939.4]
  assign _T_62029 = $signed(_T_62026) + $signed(_T_55930); // @[Modules.scala 143:103:@7941.4]
  assign _T_62030 = _T_62029[5:0]; // @[Modules.scala 143:103:@7942.4]
  assign _T_62031 = $signed(_T_62030); // @[Modules.scala 143:103:@7943.4]
  assign _T_62036 = $signed(_T_55935) + $signed(_GEN_132); // @[Modules.scala 143:103:@7947.4]
  assign _T_62037 = _T_62036[5:0]; // @[Modules.scala 143:103:@7948.4]
  assign _T_62038 = $signed(_T_62037); // @[Modules.scala 143:103:@7949.4]
  assign _T_62049 = $signed(-4'sh1) * $signed(io_in_647); // @[Modules.scala 144:80:@7958.4]
  assign _GEN_205 = {{1{_T_62049[4]}},_T_62049}; // @[Modules.scala 143:103:@7959.4]
  assign _T_62050 = $signed(_T_55949) + $signed(_GEN_205); // @[Modules.scala 143:103:@7959.4]
  assign _T_62051 = _T_62050[5:0]; // @[Modules.scala 143:103:@7960.4]
  assign _T_62052 = $signed(_T_62051); // @[Modules.scala 143:103:@7961.4]
  assign _T_62054 = $signed(-4'sh1) * $signed(io_in_648); // @[Modules.scala 143:74:@7963.4]
  assign _T_62056 = $signed(-4'sh1) * $signed(io_in_649); // @[Modules.scala 144:80:@7964.4]
  assign _T_62057 = $signed(_T_62054) + $signed(_T_62056); // @[Modules.scala 143:103:@7965.4]
  assign _T_62058 = _T_62057[4:0]; // @[Modules.scala 143:103:@7966.4]
  assign _T_62059 = $signed(_T_62058); // @[Modules.scala 143:103:@7967.4]
  assign _T_62061 = $signed(-4'sh1) * $signed(io_in_650); // @[Modules.scala 143:74:@7969.4]
  assign _T_62063 = $signed(-4'sh1) * $signed(io_in_651); // @[Modules.scala 144:80:@7970.4]
  assign _T_62064 = $signed(_T_62061) + $signed(_T_62063); // @[Modules.scala 143:103:@7971.4]
  assign _T_62065 = _T_62064[4:0]; // @[Modules.scala 143:103:@7972.4]
  assign _T_62066 = $signed(_T_62065); // @[Modules.scala 143:103:@7973.4]
  assign _T_62103 = $signed(4'sh1) * $signed(io_in_662); // @[Modules.scala 143:74:@8005.4]
  assign _T_62106 = $signed(_T_62103) + $signed(_T_59005); // @[Modules.scala 143:103:@8007.4]
  assign _T_62107 = _T_62106[5:0]; // @[Modules.scala 143:103:@8008.4]
  assign _T_62108 = $signed(_T_62107); // @[Modules.scala 143:103:@8009.4]
  assign _T_62110 = $signed(4'sh1) * $signed(io_in_664); // @[Modules.scala 143:74:@8011.4]
  assign _T_62112 = $signed(4'sh1) * $signed(io_in_665); // @[Modules.scala 144:80:@8012.4]
  assign _T_62113 = $signed(_T_62110) + $signed(_T_62112); // @[Modules.scala 143:103:@8013.4]
  assign _T_62114 = _T_62113[5:0]; // @[Modules.scala 143:103:@8014.4]
  assign _T_62115 = $signed(_T_62114); // @[Modules.scala 143:103:@8015.4]
  assign _T_62126 = $signed(-4'sh1) * $signed(io_in_669); // @[Modules.scala 144:80:@8024.4]
  assign _T_62127 = $signed(_T_59024) + $signed(_T_62126); // @[Modules.scala 143:103:@8025.4]
  assign _T_62128 = _T_62127[4:0]; // @[Modules.scala 143:103:@8026.4]
  assign _T_62129 = $signed(_T_62128); // @[Modules.scala 143:103:@8027.4]
  assign _T_62138 = $signed(-4'sh1) * $signed(io_in_675); // @[Modules.scala 143:74:@8035.4]
  assign _T_62140 = $signed(-4'sh1) * $signed(io_in_676); // @[Modules.scala 144:80:@8036.4]
  assign _T_62141 = $signed(_T_62138) + $signed(_T_62140); // @[Modules.scala 143:103:@8037.4]
  assign _T_62142 = _T_62141[4:0]; // @[Modules.scala 143:103:@8038.4]
  assign _T_62143 = $signed(_T_62142); // @[Modules.scala 143:103:@8039.4]
  assign _T_62145 = $signed(-4'sh1) * $signed(io_in_677); // @[Modules.scala 143:74:@8041.4]
  assign _T_62147 = $signed(-4'sh1) * $signed(io_in_678); // @[Modules.scala 144:80:@8042.4]
  assign _T_62148 = $signed(_T_62145) + $signed(_T_62147); // @[Modules.scala 143:103:@8043.4]
  assign _T_62149 = _T_62148[4:0]; // @[Modules.scala 143:103:@8044.4]
  assign _T_62150 = $signed(_T_62149); // @[Modules.scala 143:103:@8045.4]
  assign _T_62155 = $signed(_T_59054) + $signed(_T_59059); // @[Modules.scala 143:103:@8049.4]
  assign _T_62156 = _T_62155[5:0]; // @[Modules.scala 143:103:@8050.4]
  assign _T_62157 = $signed(_T_62156); // @[Modules.scala 143:103:@8051.4]
  assign _T_62159 = $signed(4'sh1) * $signed(io_in_682); // @[Modules.scala 143:74:@8053.4]
  assign _GEN_206 = {{1{_T_59066[4]}},_T_59066}; // @[Modules.scala 143:103:@8055.4]
  assign _T_62162 = $signed(_T_62159) + $signed(_GEN_206); // @[Modules.scala 143:103:@8055.4]
  assign _T_62163 = _T_62162[5:0]; // @[Modules.scala 143:103:@8056.4]
  assign _T_62164 = $signed(_T_62163); // @[Modules.scala 143:103:@8057.4]
  assign _T_62183 = $signed(_T_59089) + $signed(_T_59094); // @[Modules.scala 143:103:@8073.4]
  assign _T_62184 = _T_62183[5:0]; // @[Modules.scala 143:103:@8074.4]
  assign _T_62185 = $signed(_T_62184); // @[Modules.scala 143:103:@8075.4]
  assign _T_62187 = $signed(4'sh1) * $signed(io_in_693); // @[Modules.scala 143:74:@8077.4]
  assign _T_62189 = $signed(4'sh1) * $signed(io_in_694); // @[Modules.scala 144:80:@8078.4]
  assign _T_62190 = $signed(_T_62187) + $signed(_T_62189); // @[Modules.scala 143:103:@8079.4]
  assign _T_62191 = _T_62190[5:0]; // @[Modules.scala 143:103:@8080.4]
  assign _T_62192 = $signed(_T_62191); // @[Modules.scala 143:103:@8081.4]
  assign _T_62194 = $signed(4'sh1) * $signed(io_in_695); // @[Modules.scala 143:74:@8083.4]
  assign _T_62197 = $signed(_T_62194) + $signed(_GEN_136); // @[Modules.scala 143:103:@8085.4]
  assign _T_62198 = _T_62197[5:0]; // @[Modules.scala 143:103:@8086.4]
  assign _T_62199 = $signed(_T_62198); // @[Modules.scala 143:103:@8087.4]
  assign _T_62203 = $signed(-4'sh1) * $signed(io_in_702); // @[Modules.scala 144:80:@8090.4]
  assign _GEN_208 = {{1{_T_62203[4]}},_T_62203}; // @[Modules.scala 143:103:@8091.4]
  assign _T_62204 = $signed(_T_56105) + $signed(_GEN_208); // @[Modules.scala 143:103:@8091.4]
  assign _T_62205 = _T_62204[5:0]; // @[Modules.scala 143:103:@8092.4]
  assign _T_62206 = $signed(_T_62205); // @[Modules.scala 143:103:@8093.4]
  assign _T_62210 = $signed(-4'sh1) * $signed(io_in_704); // @[Modules.scala 144:80:@8096.4]
  assign _T_62211 = $signed(_T_59122) + $signed(_T_62210); // @[Modules.scala 143:103:@8097.4]
  assign _T_62212 = _T_62211[4:0]; // @[Modules.scala 143:103:@8098.4]
  assign _T_62213 = $signed(_T_62212); // @[Modules.scala 143:103:@8099.4]
  assign _T_62215 = $signed(-4'sh1) * $signed(io_in_705); // @[Modules.scala 143:74:@8101.4]
  assign _GEN_209 = {{1{_T_62215[4]}},_T_62215}; // @[Modules.scala 143:103:@8103.4]
  assign _T_62218 = $signed(_GEN_209) + $signed(_T_59129); // @[Modules.scala 143:103:@8103.4]
  assign _T_62219 = _T_62218[5:0]; // @[Modules.scala 143:103:@8104.4]
  assign _T_62220 = $signed(_T_62219); // @[Modules.scala 143:103:@8105.4]
  assign _T_62225 = $signed(_GEN_71) + $signed(_T_56131); // @[Modules.scala 143:103:@8109.4]
  assign _T_62226 = _T_62225[5:0]; // @[Modules.scala 143:103:@8110.4]
  assign _T_62227 = $signed(_T_62226); // @[Modules.scala 143:103:@8111.4]
  assign _T_62231 = $signed(-4'sh1) * $signed(io_in_711); // @[Modules.scala 144:80:@8114.4]
  assign _GEN_211 = {{1{_T_62231[4]}},_T_62231}; // @[Modules.scala 143:103:@8115.4]
  assign _T_62232 = $signed(_T_56133) + $signed(_GEN_211); // @[Modules.scala 143:103:@8115.4]
  assign _T_62233 = _T_62232[5:0]; // @[Modules.scala 143:103:@8116.4]
  assign _T_62234 = $signed(_T_62233); // @[Modules.scala 143:103:@8117.4]
  assign _T_62239 = $signed(_T_56147) + $signed(_T_56152); // @[Modules.scala 143:103:@8121.4]
  assign _T_62240 = _T_62239[4:0]; // @[Modules.scala 143:103:@8122.4]
  assign _T_62241 = $signed(_T_62240); // @[Modules.scala 143:103:@8123.4]
  assign _T_62246 = $signed(_T_56154) + $signed(_T_56159); // @[Modules.scala 143:103:@8127.4]
  assign _T_62247 = _T_62246[4:0]; // @[Modules.scala 143:103:@8128.4]
  assign _T_62248 = $signed(_T_62247); // @[Modules.scala 143:103:@8129.4]
  assign _GEN_212 = {{1{_T_56161[4]}},_T_56161}; // @[Modules.scala 143:103:@8133.4]
  assign _T_62253 = $signed(_GEN_212) + $signed(_T_59178); // @[Modules.scala 143:103:@8133.4]
  assign _T_62254 = _T_62253[5:0]; // @[Modules.scala 143:103:@8134.4]
  assign _T_62255 = $signed(_T_62254); // @[Modules.scala 143:103:@8135.4]
  assign _GEN_213 = {{1{_T_56175[4]}},_T_56175}; // @[Modules.scala 143:103:@8139.4]
  assign _T_62260 = $signed(_T_59180) + $signed(_GEN_213); // @[Modules.scala 143:103:@8139.4]
  assign _T_62261 = _T_62260[5:0]; // @[Modules.scala 143:103:@8140.4]
  assign _T_62262 = $signed(_T_62261); // @[Modules.scala 143:103:@8141.4]
  assign _T_62273 = $signed(4'sh1) * $signed(io_in_726); // @[Modules.scala 144:80:@8150.4]
  assign _GEN_214 = {{1{_T_56187[4]}},_T_56187}; // @[Modules.scala 143:103:@8151.4]
  assign _T_62274 = $signed(_GEN_214) + $signed(_T_62273); // @[Modules.scala 143:103:@8151.4]
  assign _T_62275 = _T_62274[5:0]; // @[Modules.scala 143:103:@8152.4]
  assign _T_62276 = $signed(_T_62275); // @[Modules.scala 143:103:@8153.4]
  assign _T_62278 = $signed(4'sh1) * $signed(io_in_731); // @[Modules.scala 143:74:@8155.4]
  assign _T_62280 = $signed(4'sh1) * $signed(io_in_732); // @[Modules.scala 144:80:@8156.4]
  assign _T_62281 = $signed(_T_62278) + $signed(_T_62280); // @[Modules.scala 143:103:@8157.4]
  assign _T_62282 = _T_62281[5:0]; // @[Modules.scala 143:103:@8158.4]
  assign _T_62283 = $signed(_T_62282); // @[Modules.scala 143:103:@8159.4]
  assign _T_62285 = $signed(4'sh1) * $signed(io_in_733); // @[Modules.scala 143:74:@8161.4]
  assign _T_62288 = $signed(_T_62285) + $signed(_T_59201); // @[Modules.scala 143:103:@8163.4]
  assign _T_62289 = _T_62288[5:0]; // @[Modules.scala 143:103:@8164.4]
  assign _T_62290 = $signed(_T_62289); // @[Modules.scala 143:103:@8165.4]
  assign _T_62294 = $signed(-4'sh1) * $signed(io_in_736); // @[Modules.scala 144:80:@8168.4]
  assign _GEN_215 = {{1{_T_62294[4]}},_T_62294}; // @[Modules.scala 143:103:@8169.4]
  assign _T_62295 = $signed(_T_59206) + $signed(_GEN_215); // @[Modules.scala 143:103:@8169.4]
  assign _T_62296 = _T_62295[5:0]; // @[Modules.scala 143:103:@8170.4]
  assign _T_62297 = $signed(_T_62296); // @[Modules.scala 143:103:@8171.4]
  assign _T_62299 = $signed(-4'sh1) * $signed(io_in_737); // @[Modules.scala 143:74:@8173.4]
  assign _T_62301 = $signed(-4'sh1) * $signed(io_in_738); // @[Modules.scala 144:80:@8174.4]
  assign _T_62302 = $signed(_T_62299) + $signed(_T_62301); // @[Modules.scala 143:103:@8175.4]
  assign _T_62303 = _T_62302[4:0]; // @[Modules.scala 143:103:@8176.4]
  assign _T_62304 = $signed(_T_62303); // @[Modules.scala 143:103:@8177.4]
  assign _T_62306 = $signed(-4'sh1) * $signed(io_in_739); // @[Modules.scala 143:74:@8179.4]
  assign _T_62308 = $signed(-4'sh1) * $signed(io_in_740); // @[Modules.scala 144:80:@8180.4]
  assign _T_62309 = $signed(_T_62306) + $signed(_T_62308); // @[Modules.scala 143:103:@8181.4]
  assign _T_62310 = _T_62309[4:0]; // @[Modules.scala 143:103:@8182.4]
  assign _T_62311 = $signed(_T_62310); // @[Modules.scala 143:103:@8183.4]
  assign _T_62313 = $signed(-4'sh1) * $signed(io_in_741); // @[Modules.scala 143:74:@8185.4]
  assign _T_62316 = $signed(_T_62313) + $signed(_T_56215); // @[Modules.scala 143:103:@8187.4]
  assign _T_62317 = _T_62316[4:0]; // @[Modules.scala 143:103:@8188.4]
  assign _T_62318 = $signed(_T_62317); // @[Modules.scala 143:103:@8189.4]
  assign _T_62320 = $signed(-4'sh1) * $signed(io_in_743); // @[Modules.scala 143:74:@8191.4]
  assign _T_62322 = $signed(-4'sh1) * $signed(io_in_744); // @[Modules.scala 144:80:@8192.4]
  assign _T_62323 = $signed(_T_62320) + $signed(_T_62322); // @[Modules.scala 143:103:@8193.4]
  assign _T_62324 = _T_62323[4:0]; // @[Modules.scala 143:103:@8194.4]
  assign _T_62325 = $signed(_T_62324); // @[Modules.scala 143:103:@8195.4]
  assign _T_62327 = $signed(-4'sh1) * $signed(io_in_745); // @[Modules.scala 143:74:@8197.4]
  assign _T_62330 = $signed(_T_62327) + $signed(_T_56224); // @[Modules.scala 143:103:@8199.4]
  assign _T_62331 = _T_62330[4:0]; // @[Modules.scala 143:103:@8200.4]
  assign _T_62332 = $signed(_T_62331); // @[Modules.scala 143:103:@8201.4]
  assign _GEN_216 = {{1{_T_56229[4]}},_T_56229}; // @[Modules.scala 143:103:@8205.4]
  assign _T_62337 = $signed(_GEN_216) + $signed(_T_59250); // @[Modules.scala 143:103:@8205.4]
  assign _T_62338 = _T_62337[5:0]; // @[Modules.scala 143:103:@8206.4]
  assign _T_62339 = $signed(_T_62338); // @[Modules.scala 143:103:@8207.4]
  assign _T_62344 = $signed(_T_56238) + $signed(_T_56243); // @[Modules.scala 143:103:@8211.4]
  assign _T_62345 = _T_62344[4:0]; // @[Modules.scala 143:103:@8212.4]
  assign _T_62346 = $signed(_T_62345); // @[Modules.scala 143:103:@8213.4]
  assign _T_62348 = $signed(-4'sh1) * $signed(io_in_752); // @[Modules.scala 143:74:@8215.4]
  assign _T_62350 = $signed(-4'sh1) * $signed(io_in_753); // @[Modules.scala 144:80:@8216.4]
  assign _T_62351 = $signed(_T_62348) + $signed(_T_62350); // @[Modules.scala 143:103:@8217.4]
  assign _T_62352 = _T_62351[4:0]; // @[Modules.scala 143:103:@8218.4]
  assign _T_62353 = $signed(_T_62352); // @[Modules.scala 143:103:@8219.4]
  assign _T_62362 = $signed(-4'sh1) * $signed(io_in_762); // @[Modules.scala 143:74:@8227.4]
  assign _T_62365 = $signed(_T_62362) + $signed(_T_56257); // @[Modules.scala 143:103:@8229.4]
  assign _T_62366 = _T_62365[4:0]; // @[Modules.scala 143:103:@8230.4]
  assign _T_62367 = $signed(_T_62366); // @[Modules.scala 143:103:@8231.4]
  assign _T_62371 = $signed(-4'sh1) * $signed(io_in_765); // @[Modules.scala 144:80:@8234.4]
  assign _T_62372 = $signed(_T_56259) + $signed(_T_62371); // @[Modules.scala 143:103:@8235.4]
  assign _T_62373 = _T_62372[4:0]; // @[Modules.scala 143:103:@8236.4]
  assign _T_62374 = $signed(_T_62373); // @[Modules.scala 143:103:@8237.4]
  assign _T_62376 = $signed(-4'sh1) * $signed(io_in_766); // @[Modules.scala 143:74:@8239.4]
  assign _T_62379 = $signed(_T_62376) + $signed(_T_59290); // @[Modules.scala 143:103:@8241.4]
  assign _T_62380 = _T_62379[4:0]; // @[Modules.scala 143:103:@8242.4]
  assign _T_62381 = $signed(_T_62380); // @[Modules.scala 143:103:@8243.4]
  assign _T_62385 = $signed(-4'sh1) * $signed(io_in_769); // @[Modules.scala 144:80:@8246.4]
  assign _T_62386 = $signed(_T_59292) + $signed(_T_62385); // @[Modules.scala 143:103:@8247.4]
  assign _T_62387 = _T_62386[4:0]; // @[Modules.scala 143:103:@8248.4]
  assign _T_62388 = $signed(_T_62387); // @[Modules.scala 143:103:@8249.4]
  assign _T_62390 = $signed(-4'sh1) * $signed(io_in_770); // @[Modules.scala 143:74:@8251.4]
  assign _T_62392 = $signed(-4'sh1) * $signed(io_in_771); // @[Modules.scala 144:80:@8252.4]
  assign _T_62393 = $signed(_T_62390) + $signed(_T_62392); // @[Modules.scala 143:103:@8253.4]
  assign _T_62394 = _T_62393[4:0]; // @[Modules.scala 143:103:@8254.4]
  assign _T_62395 = $signed(_T_62394); // @[Modules.scala 143:103:@8255.4]
  assign _T_62397 = $signed(-4'sh1) * $signed(io_in_772); // @[Modules.scala 143:74:@8257.4]
  assign _T_62399 = $signed(-4'sh1) * $signed(io_in_773); // @[Modules.scala 144:80:@8258.4]
  assign _T_62400 = $signed(_T_62397) + $signed(_T_62399); // @[Modules.scala 143:103:@8259.4]
  assign _T_62401 = _T_62400[4:0]; // @[Modules.scala 143:103:@8260.4]
  assign _T_62402 = $signed(_T_62401); // @[Modules.scala 143:103:@8261.4]
  assign _T_62404 = $signed(-4'sh1) * $signed(io_in_774); // @[Modules.scala 143:74:@8263.4]
  assign _GEN_217 = {{1{_T_62404[4]}},_T_62404}; // @[Modules.scala 143:103:@8265.4]
  assign _T_62407 = $signed(_GEN_217) + $signed(_T_59318); // @[Modules.scala 143:103:@8265.4]
  assign _T_62408 = _T_62407[5:0]; // @[Modules.scala 143:103:@8266.4]
  assign _T_62409 = $signed(_T_62408); // @[Modules.scala 143:103:@8267.4]
  assign _T_62414 = $signed(_T_59320) + $signed(_T_56299); // @[Modules.scala 143:103:@8271.4]
  assign _T_62415 = _T_62414[5:0]; // @[Modules.scala 143:103:@8272.4]
  assign _T_62416 = $signed(_T_62415); // @[Modules.scala 143:103:@8273.4]
  assign buffer_2_0 = {{9{_T_60253[4]}},_T_60253}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_1 = {{9{_T_60260[4]}},_T_60260}; // @[Modules.scala 112:22:@8.4]
  assign _T_62417 = $signed(buffer_2_0) + $signed(buffer_2_1); // @[Modules.scala 160:64:@8275.4]
  assign _T_62418 = _T_62417[13:0]; // @[Modules.scala 160:64:@8276.4]
  assign buffer_2_310 = $signed(_T_62418); // @[Modules.scala 160:64:@8277.4]
  assign buffer_2_2 = {{9{_T_60267[4]}},_T_60267}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_3 = {{9{_T_60274[4]}},_T_60274}; // @[Modules.scala 112:22:@8.4]
  assign _T_62420 = $signed(buffer_2_2) + $signed(buffer_2_3); // @[Modules.scala 160:64:@8279.4]
  assign _T_62421 = _T_62420[13:0]; // @[Modules.scala 160:64:@8280.4]
  assign buffer_2_311 = $signed(_T_62421); // @[Modules.scala 160:64:@8281.4]
  assign buffer_2_4 = {{8{_T_60281[5]}},_T_60281}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_5 = {{8{_T_60288[5]}},_T_60288}; // @[Modules.scala 112:22:@8.4]
  assign _T_62423 = $signed(buffer_2_4) + $signed(buffer_2_5); // @[Modules.scala 160:64:@8283.4]
  assign _T_62424 = _T_62423[13:0]; // @[Modules.scala 160:64:@8284.4]
  assign buffer_2_312 = $signed(_T_62424); // @[Modules.scala 160:64:@8285.4]
  assign buffer_2_6 = {{9{_T_60295[4]}},_T_60295}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_7 = {{8{_T_60302[5]}},_T_60302}; // @[Modules.scala 112:22:@8.4]
  assign _T_62426 = $signed(buffer_2_6) + $signed(buffer_2_7); // @[Modules.scala 160:64:@8287.4]
  assign _T_62427 = _T_62426[13:0]; // @[Modules.scala 160:64:@8288.4]
  assign buffer_2_313 = $signed(_T_62427); // @[Modules.scala 160:64:@8289.4]
  assign buffer_2_8 = {{9{_T_60309[4]}},_T_60309}; // @[Modules.scala 112:22:@8.4]
  assign _T_62429 = $signed(buffer_2_8) + $signed(buffer_0_9); // @[Modules.scala 160:64:@8291.4]
  assign _T_62430 = _T_62429[13:0]; // @[Modules.scala 160:64:@8292.4]
  assign buffer_2_314 = $signed(_T_62430); // @[Modules.scala 160:64:@8293.4]
  assign buffer_2_11 = {{9{_T_60330[4]}},_T_60330}; // @[Modules.scala 112:22:@8.4]
  assign _T_62432 = $signed(buffer_0_10) + $signed(buffer_2_11); // @[Modules.scala 160:64:@8295.4]
  assign _T_62433 = _T_62432[13:0]; // @[Modules.scala 160:64:@8296.4]
  assign buffer_2_315 = $signed(_T_62433); // @[Modules.scala 160:64:@8297.4]
  assign buffer_2_12 = {{9{_T_60337[4]}},_T_60337}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_13 = {{9{_T_60344[4]}},_T_60344}; // @[Modules.scala 112:22:@8.4]
  assign _T_62435 = $signed(buffer_2_12) + $signed(buffer_2_13); // @[Modules.scala 160:64:@8299.4]
  assign _T_62436 = _T_62435[13:0]; // @[Modules.scala 160:64:@8300.4]
  assign buffer_2_316 = $signed(_T_62436); // @[Modules.scala 160:64:@8301.4]
  assign buffer_2_14 = {{9{_T_60351[4]}},_T_60351}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_15 = {{9{_T_60358[4]}},_T_60358}; // @[Modules.scala 112:22:@8.4]
  assign _T_62438 = $signed(buffer_2_14) + $signed(buffer_2_15); // @[Modules.scala 160:64:@8303.4]
  assign _T_62439 = _T_62438[13:0]; // @[Modules.scala 160:64:@8304.4]
  assign buffer_2_317 = $signed(_T_62439); // @[Modules.scala 160:64:@8305.4]
  assign buffer_2_16 = {{9{_T_60365[4]}},_T_60365}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_17 = {{8{_T_60372[5]}},_T_60372}; // @[Modules.scala 112:22:@8.4]
  assign _T_62441 = $signed(buffer_2_16) + $signed(buffer_2_17); // @[Modules.scala 160:64:@8307.4]
  assign _T_62442 = _T_62441[13:0]; // @[Modules.scala 160:64:@8308.4]
  assign buffer_2_318 = $signed(_T_62442); // @[Modules.scala 160:64:@8309.4]
  assign _T_62444 = $signed(buffer_1_19) + $signed(buffer_1_20); // @[Modules.scala 160:64:@8311.4]
  assign _T_62445 = _T_62444[13:0]; // @[Modules.scala 160:64:@8312.4]
  assign buffer_2_319 = $signed(_T_62445); // @[Modules.scala 160:64:@8313.4]
  assign _T_62447 = $signed(buffer_1_21) + $signed(buffer_1_22); // @[Modules.scala 160:64:@8315.4]
  assign _T_62448 = _T_62447[13:0]; // @[Modules.scala 160:64:@8316.4]
  assign buffer_2_320 = $signed(_T_62448); // @[Modules.scala 160:64:@8317.4]
  assign buffer_2_22 = {{9{_T_60407[4]}},_T_60407}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_23 = {{8{_T_60414[5]}},_T_60414}; // @[Modules.scala 112:22:@8.4]
  assign _T_62450 = $signed(buffer_2_22) + $signed(buffer_2_23); // @[Modules.scala 160:64:@8319.4]
  assign _T_62451 = _T_62450[13:0]; // @[Modules.scala 160:64:@8320.4]
  assign buffer_2_321 = $signed(_T_62451); // @[Modules.scala 160:64:@8321.4]
  assign buffer_2_24 = {{8{_T_60421[5]}},_T_60421}; // @[Modules.scala 112:22:@8.4]
  assign _T_62453 = $signed(buffer_2_24) + $signed(buffer_1_27); // @[Modules.scala 160:64:@8323.4]
  assign _T_62454 = _T_62453[13:0]; // @[Modules.scala 160:64:@8324.4]
  assign buffer_2_322 = $signed(_T_62454); // @[Modules.scala 160:64:@8325.4]
  assign buffer_2_26 = {{8{_T_60435[5]}},_T_60435}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_27 = {{8{_T_60442[5]}},_T_60442}; // @[Modules.scala 112:22:@8.4]
  assign _T_62456 = $signed(buffer_2_26) + $signed(buffer_2_27); // @[Modules.scala 160:64:@8327.4]
  assign _T_62457 = _T_62456[13:0]; // @[Modules.scala 160:64:@8328.4]
  assign buffer_2_323 = $signed(_T_62457); // @[Modules.scala 160:64:@8329.4]
  assign buffer_2_28 = {{8{_T_60449[5]}},_T_60449}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_29 = {{8{_T_60456[5]}},_T_60456}; // @[Modules.scala 112:22:@8.4]
  assign _T_62459 = $signed(buffer_2_28) + $signed(buffer_2_29); // @[Modules.scala 160:64:@8331.4]
  assign _T_62460 = _T_62459[13:0]; // @[Modules.scala 160:64:@8332.4]
  assign buffer_2_324 = $signed(_T_62460); // @[Modules.scala 160:64:@8333.4]
  assign buffer_2_30 = {{8{_T_60463[5]}},_T_60463}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_31 = {{8{_T_60470[5]}},_T_60470}; // @[Modules.scala 112:22:@8.4]
  assign _T_62462 = $signed(buffer_2_30) + $signed(buffer_2_31); // @[Modules.scala 160:64:@8335.4]
  assign _T_62463 = _T_62462[13:0]; // @[Modules.scala 160:64:@8336.4]
  assign buffer_2_325 = $signed(_T_62463); // @[Modules.scala 160:64:@8337.4]
  assign buffer_2_32 = {{9{_T_60477[4]}},_T_60477}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_33 = {{8{_T_60484[5]}},_T_60484}; // @[Modules.scala 112:22:@8.4]
  assign _T_62465 = $signed(buffer_2_32) + $signed(buffer_2_33); // @[Modules.scala 160:64:@8339.4]
  assign _T_62466 = _T_62465[13:0]; // @[Modules.scala 160:64:@8340.4]
  assign buffer_2_326 = $signed(_T_62466); // @[Modules.scala 160:64:@8341.4]
  assign buffer_2_34 = {{8{_T_60491[5]}},_T_60491}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_35 = {{8{_T_60498[5]}},_T_60498}; // @[Modules.scala 112:22:@8.4]
  assign _T_62468 = $signed(buffer_2_34) + $signed(buffer_2_35); // @[Modules.scala 160:64:@8343.4]
  assign _T_62469 = _T_62468[13:0]; // @[Modules.scala 160:64:@8344.4]
  assign buffer_2_327 = $signed(_T_62469); // @[Modules.scala 160:64:@8345.4]
  assign buffer_2_36 = {{9{_T_60505[4]}},_T_60505}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_37 = {{9{_T_60512[4]}},_T_60512}; // @[Modules.scala 112:22:@8.4]
  assign _T_62471 = $signed(buffer_2_36) + $signed(buffer_2_37); // @[Modules.scala 160:64:@8347.4]
  assign _T_62472 = _T_62471[13:0]; // @[Modules.scala 160:64:@8348.4]
  assign buffer_2_328 = $signed(_T_62472); // @[Modules.scala 160:64:@8349.4]
  assign buffer_2_38 = {{8{_T_60519[5]}},_T_60519}; // @[Modules.scala 112:22:@8.4]
  assign _T_62474 = $signed(buffer_2_38) + $signed(buffer_0_42); // @[Modules.scala 160:64:@8351.4]
  assign _T_62475 = _T_62474[13:0]; // @[Modules.scala 160:64:@8352.4]
  assign buffer_2_329 = $signed(_T_62475); // @[Modules.scala 160:64:@8353.4]
  assign _T_62477 = $signed(buffer_1_41) + $signed(buffer_1_42); // @[Modules.scala 160:64:@8355.4]
  assign _T_62478 = _T_62477[13:0]; // @[Modules.scala 160:64:@8356.4]
  assign buffer_2_330 = $signed(_T_62478); // @[Modules.scala 160:64:@8357.4]
  assign buffer_2_42 = {{8{_T_60547[5]}},_T_60547}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_43 = {{8{_T_60554[5]}},_T_60554}; // @[Modules.scala 112:22:@8.4]
  assign _T_62480 = $signed(buffer_2_42) + $signed(buffer_2_43); // @[Modules.scala 160:64:@8359.4]
  assign _T_62481 = _T_62480[13:0]; // @[Modules.scala 160:64:@8360.4]
  assign buffer_2_331 = $signed(_T_62481); // @[Modules.scala 160:64:@8361.4]
  assign buffer_2_44 = {{8{_T_60561[5]}},_T_60561}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_45 = {{9{_T_60568[4]}},_T_60568}; // @[Modules.scala 112:22:@8.4]
  assign _T_62483 = $signed(buffer_2_44) + $signed(buffer_2_45); // @[Modules.scala 160:64:@8363.4]
  assign _T_62484 = _T_62483[13:0]; // @[Modules.scala 160:64:@8364.4]
  assign buffer_2_332 = $signed(_T_62484); // @[Modules.scala 160:64:@8365.4]
  assign buffer_2_46 = {{8{_T_60575[5]}},_T_60575}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_47 = {{9{_T_60582[4]}},_T_60582}; // @[Modules.scala 112:22:@8.4]
  assign _T_62486 = $signed(buffer_2_46) + $signed(buffer_2_47); // @[Modules.scala 160:64:@8367.4]
  assign _T_62487 = _T_62486[13:0]; // @[Modules.scala 160:64:@8368.4]
  assign buffer_2_333 = $signed(_T_62487); // @[Modules.scala 160:64:@8369.4]
  assign buffer_2_48 = {{9{_T_60589[4]}},_T_60589}; // @[Modules.scala 112:22:@8.4]
  assign _T_62489 = $signed(buffer_2_48) + $signed(buffer_1_50); // @[Modules.scala 160:64:@8371.4]
  assign _T_62490 = _T_62489[13:0]; // @[Modules.scala 160:64:@8372.4]
  assign buffer_2_334 = $signed(_T_62490); // @[Modules.scala 160:64:@8373.4]
  assign buffer_2_51 = {{8{_T_60610[5]}},_T_60610}; // @[Modules.scala 112:22:@8.4]
  assign _T_62492 = $signed(buffer_1_51) + $signed(buffer_2_51); // @[Modules.scala 160:64:@8375.4]
  assign _T_62493 = _T_62492[13:0]; // @[Modules.scala 160:64:@8376.4]
  assign buffer_2_335 = $signed(_T_62493); // @[Modules.scala 160:64:@8377.4]
  assign buffer_2_52 = {{8{_T_60617[5]}},_T_60617}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_53 = {{8{_T_60624[5]}},_T_60624}; // @[Modules.scala 112:22:@8.4]
  assign _T_62495 = $signed(buffer_2_52) + $signed(buffer_2_53); // @[Modules.scala 160:64:@8379.4]
  assign _T_62496 = _T_62495[13:0]; // @[Modules.scala 160:64:@8380.4]
  assign buffer_2_336 = $signed(_T_62496); // @[Modules.scala 160:64:@8381.4]
  assign buffer_2_54 = {{8{_T_60631[5]}},_T_60631}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_55 = {{8{_T_60638[5]}},_T_60638}; // @[Modules.scala 112:22:@8.4]
  assign _T_62498 = $signed(buffer_2_54) + $signed(buffer_2_55); // @[Modules.scala 160:64:@8383.4]
  assign _T_62499 = _T_62498[13:0]; // @[Modules.scala 160:64:@8384.4]
  assign buffer_2_337 = $signed(_T_62499); // @[Modules.scala 160:64:@8385.4]
  assign buffer_2_56 = {{8{_T_60645[5]}},_T_60645}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_57 = {{8{_T_60652[5]}},_T_60652}; // @[Modules.scala 112:22:@8.4]
  assign _T_62501 = $signed(buffer_2_56) + $signed(buffer_2_57); // @[Modules.scala 160:64:@8387.4]
  assign _T_62502 = _T_62501[13:0]; // @[Modules.scala 160:64:@8388.4]
  assign buffer_2_338 = $signed(_T_62502); // @[Modules.scala 160:64:@8389.4]
  assign buffer_2_58 = {{9{_T_60659[4]}},_T_60659}; // @[Modules.scala 112:22:@8.4]
  assign _T_62504 = $signed(buffer_2_58) + $signed(buffer_0_59); // @[Modules.scala 160:64:@8391.4]
  assign _T_62505 = _T_62504[13:0]; // @[Modules.scala 160:64:@8392.4]
  assign buffer_2_339 = $signed(_T_62505); // @[Modules.scala 160:64:@8393.4]
  assign buffer_2_60 = {{9{_T_60673[4]}},_T_60673}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_61 = {{9{_T_60680[4]}},_T_60680}; // @[Modules.scala 112:22:@8.4]
  assign _T_62507 = $signed(buffer_2_60) + $signed(buffer_2_61); // @[Modules.scala 160:64:@8395.4]
  assign _T_62508 = _T_62507[13:0]; // @[Modules.scala 160:64:@8396.4]
  assign buffer_2_340 = $signed(_T_62508); // @[Modules.scala 160:64:@8397.4]
  assign buffer_2_63 = {{9{_T_60694[4]}},_T_60694}; // @[Modules.scala 112:22:@8.4]
  assign _T_62510 = $signed(buffer_1_63) + $signed(buffer_2_63); // @[Modules.scala 160:64:@8399.4]
  assign _T_62511 = _T_62510[13:0]; // @[Modules.scala 160:64:@8400.4]
  assign buffer_2_341 = $signed(_T_62511); // @[Modules.scala 160:64:@8401.4]
  assign buffer_2_64 = {{8{_T_60701[5]}},_T_60701}; // @[Modules.scala 112:22:@8.4]
  assign _T_62513 = $signed(buffer_2_64) + $signed(buffer_1_65); // @[Modules.scala 160:64:@8403.4]
  assign _T_62514 = _T_62513[13:0]; // @[Modules.scala 160:64:@8404.4]
  assign buffer_2_342 = $signed(_T_62514); // @[Modules.scala 160:64:@8405.4]
  assign buffer_2_67 = {{9{_T_60722[4]}},_T_60722}; // @[Modules.scala 112:22:@8.4]
  assign _T_62516 = $signed(buffer_1_66) + $signed(buffer_2_67); // @[Modules.scala 160:64:@8407.4]
  assign _T_62517 = _T_62516[13:0]; // @[Modules.scala 160:64:@8408.4]
  assign buffer_2_343 = $signed(_T_62517); // @[Modules.scala 160:64:@8409.4]
  assign buffer_2_68 = {{9{_T_60729[4]}},_T_60729}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_69 = {{8{_T_60736[5]}},_T_60736}; // @[Modules.scala 112:22:@8.4]
  assign _T_62519 = $signed(buffer_2_68) + $signed(buffer_2_69); // @[Modules.scala 160:64:@8411.4]
  assign _T_62520 = _T_62519[13:0]; // @[Modules.scala 160:64:@8412.4]
  assign buffer_2_344 = $signed(_T_62520); // @[Modules.scala 160:64:@8413.4]
  assign buffer_2_70 = {{9{_T_60743[4]}},_T_60743}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_71 = {{9{_T_60750[4]}},_T_60750}; // @[Modules.scala 112:22:@8.4]
  assign _T_62522 = $signed(buffer_2_70) + $signed(buffer_2_71); // @[Modules.scala 160:64:@8415.4]
  assign _T_62523 = _T_62522[13:0]; // @[Modules.scala 160:64:@8416.4]
  assign buffer_2_345 = $signed(_T_62523); // @[Modules.scala 160:64:@8417.4]
  assign buffer_2_72 = {{9{_T_60757[4]}},_T_60757}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_73 = {{9{_T_60764[4]}},_T_60764}; // @[Modules.scala 112:22:@8.4]
  assign _T_62525 = $signed(buffer_2_72) + $signed(buffer_2_73); // @[Modules.scala 160:64:@8419.4]
  assign _T_62526 = _T_62525[13:0]; // @[Modules.scala 160:64:@8420.4]
  assign buffer_2_346 = $signed(_T_62526); // @[Modules.scala 160:64:@8421.4]
  assign buffer_2_75 = {{9{_T_60778[4]}},_T_60778}; // @[Modules.scala 112:22:@8.4]
  assign _T_62528 = $signed(buffer_0_71) + $signed(buffer_2_75); // @[Modules.scala 160:64:@8423.4]
  assign _T_62529 = _T_62528[13:0]; // @[Modules.scala 160:64:@8424.4]
  assign buffer_2_347 = $signed(_T_62529); // @[Modules.scala 160:64:@8425.4]
  assign buffer_2_76 = {{9{_T_60785[4]}},_T_60785}; // @[Modules.scala 112:22:@8.4]
  assign _T_62531 = $signed(buffer_2_76) + $signed(buffer_0_74); // @[Modules.scala 160:64:@8427.4]
  assign _T_62532 = _T_62531[13:0]; // @[Modules.scala 160:64:@8428.4]
  assign buffer_2_348 = $signed(_T_62532); // @[Modules.scala 160:64:@8429.4]
  assign buffer_2_80 = {{9{_T_60813[4]}},_T_60813}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_81 = {{9{_T_60820[4]}},_T_60820}; // @[Modules.scala 112:22:@8.4]
  assign _T_62537 = $signed(buffer_2_80) + $signed(buffer_2_81); // @[Modules.scala 160:64:@8435.4]
  assign _T_62538 = _T_62537[13:0]; // @[Modules.scala 160:64:@8436.4]
  assign buffer_2_350 = $signed(_T_62538); // @[Modules.scala 160:64:@8437.4]
  assign buffer_2_82 = {{9{_T_60827[4]}},_T_60827}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_83 = {{9{_T_60834[4]}},_T_60834}; // @[Modules.scala 112:22:@8.4]
  assign _T_62540 = $signed(buffer_2_82) + $signed(buffer_2_83); // @[Modules.scala 160:64:@8439.4]
  assign _T_62541 = _T_62540[13:0]; // @[Modules.scala 160:64:@8440.4]
  assign buffer_2_351 = $signed(_T_62541); // @[Modules.scala 160:64:@8441.4]
  assign buffer_2_84 = {{8{_T_60841[5]}},_T_60841}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_85 = {{9{_T_60848[4]}},_T_60848}; // @[Modules.scala 112:22:@8.4]
  assign _T_62543 = $signed(buffer_2_84) + $signed(buffer_2_85); // @[Modules.scala 160:64:@8443.4]
  assign _T_62544 = _T_62543[13:0]; // @[Modules.scala 160:64:@8444.4]
  assign buffer_2_352 = $signed(_T_62544); // @[Modules.scala 160:64:@8445.4]
  assign buffer_2_86 = {{9{_T_60855[4]}},_T_60855}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_87 = {{9{_T_60862[4]}},_T_60862}; // @[Modules.scala 112:22:@8.4]
  assign _T_62546 = $signed(buffer_2_86) + $signed(buffer_2_87); // @[Modules.scala 160:64:@8447.4]
  assign _T_62547 = _T_62546[13:0]; // @[Modules.scala 160:64:@8448.4]
  assign buffer_2_353 = $signed(_T_62547); // @[Modules.scala 160:64:@8449.4]
  assign buffer_2_88 = {{9{_T_60869[4]}},_T_60869}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_89 = {{9{_T_60876[4]}},_T_60876}; // @[Modules.scala 112:22:@8.4]
  assign _T_62549 = $signed(buffer_2_88) + $signed(buffer_2_89); // @[Modules.scala 160:64:@8451.4]
  assign _T_62550 = _T_62549[13:0]; // @[Modules.scala 160:64:@8452.4]
  assign buffer_2_354 = $signed(_T_62550); // @[Modules.scala 160:64:@8453.4]
  assign buffer_2_90 = {{9{_T_60883[4]}},_T_60883}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_91 = {{9{_T_60890[4]}},_T_60890}; // @[Modules.scala 112:22:@8.4]
  assign _T_62552 = $signed(buffer_2_90) + $signed(buffer_2_91); // @[Modules.scala 160:64:@8455.4]
  assign _T_62553 = _T_62552[13:0]; // @[Modules.scala 160:64:@8456.4]
  assign buffer_2_355 = $signed(_T_62553); // @[Modules.scala 160:64:@8457.4]
  assign buffer_2_92 = {{8{_T_60897[5]}},_T_60897}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_93 = {{9{_T_60904[4]}},_T_60904}; // @[Modules.scala 112:22:@8.4]
  assign _T_62555 = $signed(buffer_2_92) + $signed(buffer_2_93); // @[Modules.scala 160:64:@8459.4]
  assign _T_62556 = _T_62555[13:0]; // @[Modules.scala 160:64:@8460.4]
  assign buffer_2_356 = $signed(_T_62556); // @[Modules.scala 160:64:@8461.4]
  assign buffer_2_94 = {{9{_T_60911[4]}},_T_60911}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_95 = {{9{_T_60918[4]}},_T_60918}; // @[Modules.scala 112:22:@8.4]
  assign _T_62558 = $signed(buffer_2_94) + $signed(buffer_2_95); // @[Modules.scala 160:64:@8463.4]
  assign _T_62559 = _T_62558[13:0]; // @[Modules.scala 160:64:@8464.4]
  assign buffer_2_357 = $signed(_T_62559); // @[Modules.scala 160:64:@8465.4]
  assign buffer_2_96 = {{8{_T_60925[5]}},_T_60925}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_97 = {{9{_T_60932[4]}},_T_60932}; // @[Modules.scala 112:22:@8.4]
  assign _T_62561 = $signed(buffer_2_96) + $signed(buffer_2_97); // @[Modules.scala 160:64:@8467.4]
  assign _T_62562 = _T_62561[13:0]; // @[Modules.scala 160:64:@8468.4]
  assign buffer_2_358 = $signed(_T_62562); // @[Modules.scala 160:64:@8469.4]
  assign buffer_2_98 = {{9{_T_60939[4]}},_T_60939}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_99 = {{9{_T_60946[4]}},_T_60946}; // @[Modules.scala 112:22:@8.4]
  assign _T_62564 = $signed(buffer_2_98) + $signed(buffer_2_99); // @[Modules.scala 160:64:@8471.4]
  assign _T_62565 = _T_62564[13:0]; // @[Modules.scala 160:64:@8472.4]
  assign buffer_2_359 = $signed(_T_62565); // @[Modules.scala 160:64:@8473.4]
  assign _T_62567 = $signed(buffer_0_95) + $signed(buffer_0_96); // @[Modules.scala 160:64:@8475.4]
  assign _T_62568 = _T_62567[13:0]; // @[Modules.scala 160:64:@8476.4]
  assign buffer_2_360 = $signed(_T_62568); // @[Modules.scala 160:64:@8477.4]
  assign buffer_2_105 = {{9{_T_60988[4]}},_T_60988}; // @[Modules.scala 112:22:@8.4]
  assign _T_62573 = $signed(buffer_0_99) + $signed(buffer_2_105); // @[Modules.scala 160:64:@8483.4]
  assign _T_62574 = _T_62573[13:0]; // @[Modules.scala 160:64:@8484.4]
  assign buffer_2_362 = $signed(_T_62574); // @[Modules.scala 160:64:@8485.4]
  assign buffer_2_106 = {{9{_T_60995[4]}},_T_60995}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_107 = {{9{_T_61002[4]}},_T_61002}; // @[Modules.scala 112:22:@8.4]
  assign _T_62576 = $signed(buffer_2_106) + $signed(buffer_2_107); // @[Modules.scala 160:64:@8487.4]
  assign _T_62577 = _T_62576[13:0]; // @[Modules.scala 160:64:@8488.4]
  assign buffer_2_363 = $signed(_T_62577); // @[Modules.scala 160:64:@8489.4]
  assign buffer_2_108 = {{8{_T_61009[5]}},_T_61009}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_109 = {{9{_T_61016[4]}},_T_61016}; // @[Modules.scala 112:22:@8.4]
  assign _T_62579 = $signed(buffer_2_108) + $signed(buffer_2_109); // @[Modules.scala 160:64:@8491.4]
  assign _T_62580 = _T_62579[13:0]; // @[Modules.scala 160:64:@8492.4]
  assign buffer_2_364 = $signed(_T_62580); // @[Modules.scala 160:64:@8493.4]
  assign buffer_2_110 = {{9{_T_61023[4]}},_T_61023}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_111 = {{9{_T_61030[4]}},_T_61030}; // @[Modules.scala 112:22:@8.4]
  assign _T_62582 = $signed(buffer_2_110) + $signed(buffer_2_111); // @[Modules.scala 160:64:@8495.4]
  assign _T_62583 = _T_62582[13:0]; // @[Modules.scala 160:64:@8496.4]
  assign buffer_2_365 = $signed(_T_62583); // @[Modules.scala 160:64:@8497.4]
  assign buffer_2_112 = {{9{_T_61037[4]}},_T_61037}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_113 = {{9{_T_61044[4]}},_T_61044}; // @[Modules.scala 112:22:@8.4]
  assign _T_62585 = $signed(buffer_2_112) + $signed(buffer_2_113); // @[Modules.scala 160:64:@8499.4]
  assign _T_62586 = _T_62585[13:0]; // @[Modules.scala 160:64:@8500.4]
  assign buffer_2_366 = $signed(_T_62586); // @[Modules.scala 160:64:@8501.4]
  assign buffer_2_116 = {{8{_T_61065[5]}},_T_61065}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_117 = {{9{_T_61072[4]}},_T_61072}; // @[Modules.scala 112:22:@8.4]
  assign _T_62591 = $signed(buffer_2_116) + $signed(buffer_2_117); // @[Modules.scala 160:64:@8507.4]
  assign _T_62592 = _T_62591[13:0]; // @[Modules.scala 160:64:@8508.4]
  assign buffer_2_368 = $signed(_T_62592); // @[Modules.scala 160:64:@8509.4]
  assign buffer_2_118 = {{9{_T_61079[4]}},_T_61079}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_119 = {{8{_T_61086[5]}},_T_61086}; // @[Modules.scala 112:22:@8.4]
  assign _T_62594 = $signed(buffer_2_118) + $signed(buffer_2_119); // @[Modules.scala 160:64:@8511.4]
  assign _T_62595 = _T_62594[13:0]; // @[Modules.scala 160:64:@8512.4]
  assign buffer_2_369 = $signed(_T_62595); // @[Modules.scala 160:64:@8513.4]
  assign buffer_2_120 = {{8{_T_61093[5]}},_T_61093}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_121 = {{8{_T_61100[5]}},_T_61100}; // @[Modules.scala 112:22:@8.4]
  assign _T_62597 = $signed(buffer_2_120) + $signed(buffer_2_121); // @[Modules.scala 160:64:@8515.4]
  assign _T_62598 = _T_62597[13:0]; // @[Modules.scala 160:64:@8516.4]
  assign buffer_2_370 = $signed(_T_62598); // @[Modules.scala 160:64:@8517.4]
  assign buffer_2_122 = {{9{_T_61107[4]}},_T_61107}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_123 = {{8{_T_61114[5]}},_T_61114}; // @[Modules.scala 112:22:@8.4]
  assign _T_62600 = $signed(buffer_2_122) + $signed(buffer_2_123); // @[Modules.scala 160:64:@8519.4]
  assign _T_62601 = _T_62600[13:0]; // @[Modules.scala 160:64:@8520.4]
  assign buffer_2_371 = $signed(_T_62601); // @[Modules.scala 160:64:@8521.4]
  assign buffer_2_124 = {{8{_T_61121[5]}},_T_61121}; // @[Modules.scala 112:22:@8.4]
  assign _T_62603 = $signed(buffer_2_124) + $signed(buffer_0_122); // @[Modules.scala 160:64:@8523.4]
  assign _T_62604 = _T_62603[13:0]; // @[Modules.scala 160:64:@8524.4]
  assign buffer_2_372 = $signed(_T_62604); // @[Modules.scala 160:64:@8525.4]
  assign _T_62606 = $signed(buffer_0_123) + $signed(buffer_0_124); // @[Modules.scala 160:64:@8527.4]
  assign _T_62607 = _T_62606[13:0]; // @[Modules.scala 160:64:@8528.4]
  assign buffer_2_373 = $signed(_T_62607); // @[Modules.scala 160:64:@8529.4]
  assign buffer_2_128 = {{8{_T_61149[5]}},_T_61149}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_129 = {{9{_T_61156[4]}},_T_61156}; // @[Modules.scala 112:22:@8.4]
  assign _T_62609 = $signed(buffer_2_128) + $signed(buffer_2_129); // @[Modules.scala 160:64:@8531.4]
  assign _T_62610 = _T_62609[13:0]; // @[Modules.scala 160:64:@8532.4]
  assign buffer_2_374 = $signed(_T_62610); // @[Modules.scala 160:64:@8533.4]
  assign buffer_2_130 = {{8{_T_61163[5]}},_T_61163}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_131 = {{8{_T_61170[5]}},_T_61170}; // @[Modules.scala 112:22:@8.4]
  assign _T_62612 = $signed(buffer_2_130) + $signed(buffer_2_131); // @[Modules.scala 160:64:@8535.4]
  assign _T_62613 = _T_62612[13:0]; // @[Modules.scala 160:64:@8536.4]
  assign buffer_2_375 = $signed(_T_62613); // @[Modules.scala 160:64:@8537.4]
  assign buffer_2_132 = {{8{_T_61177[5]}},_T_61177}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_133 = {{8{_T_61184[5]}},_T_61184}; // @[Modules.scala 112:22:@8.4]
  assign _T_62615 = $signed(buffer_2_132) + $signed(buffer_2_133); // @[Modules.scala 160:64:@8539.4]
  assign _T_62616 = _T_62615[13:0]; // @[Modules.scala 160:64:@8540.4]
  assign buffer_2_376 = $signed(_T_62616); // @[Modules.scala 160:64:@8541.4]
  assign buffer_2_134 = {{8{_T_61191[5]}},_T_61191}; // @[Modules.scala 112:22:@8.4]
  assign _T_62618 = $signed(buffer_2_134) + $signed(buffer_1_134); // @[Modules.scala 160:64:@8543.4]
  assign _T_62619 = _T_62618[13:0]; // @[Modules.scala 160:64:@8544.4]
  assign buffer_2_377 = $signed(_T_62619); // @[Modules.scala 160:64:@8545.4]
  assign buffer_2_137 = {{8{_T_61212[5]}},_T_61212}; // @[Modules.scala 112:22:@8.4]
  assign _T_62621 = $signed(buffer_1_135) + $signed(buffer_2_137); // @[Modules.scala 160:64:@8547.4]
  assign _T_62622 = _T_62621[13:0]; // @[Modules.scala 160:64:@8548.4]
  assign buffer_2_378 = $signed(_T_62622); // @[Modules.scala 160:64:@8549.4]
  assign buffer_2_138 = {{8{_T_61219[5]}},_T_61219}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_139 = {{9{_T_61226[4]}},_T_61226}; // @[Modules.scala 112:22:@8.4]
  assign _T_62624 = $signed(buffer_2_138) + $signed(buffer_2_139); // @[Modules.scala 160:64:@8551.4]
  assign _T_62625 = _T_62624[13:0]; // @[Modules.scala 160:64:@8552.4]
  assign buffer_2_379 = $signed(_T_62625); // @[Modules.scala 160:64:@8553.4]
  assign buffer_2_140 = {{9{_T_61233[4]}},_T_61233}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_141 = {{8{_T_61240[5]}},_T_61240}; // @[Modules.scala 112:22:@8.4]
  assign _T_62627 = $signed(buffer_2_140) + $signed(buffer_2_141); // @[Modules.scala 160:64:@8555.4]
  assign _T_62628 = _T_62627[13:0]; // @[Modules.scala 160:64:@8556.4]
  assign buffer_2_380 = $signed(_T_62628); // @[Modules.scala 160:64:@8557.4]
  assign buffer_2_142 = {{9{_T_61247[4]}},_T_61247}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_143 = {{8{_T_61254[5]}},_T_61254}; // @[Modules.scala 112:22:@8.4]
  assign _T_62630 = $signed(buffer_2_142) + $signed(buffer_2_143); // @[Modules.scala 160:64:@8559.4]
  assign _T_62631 = _T_62630[13:0]; // @[Modules.scala 160:64:@8560.4]
  assign buffer_2_381 = $signed(_T_62631); // @[Modules.scala 160:64:@8561.4]
  assign buffer_2_144 = {{8{_T_61261[5]}},_T_61261}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_145 = {{8{_T_61268[5]}},_T_61268}; // @[Modules.scala 112:22:@8.4]
  assign _T_62633 = $signed(buffer_2_144) + $signed(buffer_2_145); // @[Modules.scala 160:64:@8563.4]
  assign _T_62634 = _T_62633[13:0]; // @[Modules.scala 160:64:@8564.4]
  assign buffer_2_382 = $signed(_T_62634); // @[Modules.scala 160:64:@8565.4]
  assign buffer_2_146 = {{8{_T_61275[5]}},_T_61275}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_147 = {{8{_T_61282[5]}},_T_61282}; // @[Modules.scala 112:22:@8.4]
  assign _T_62636 = $signed(buffer_2_146) + $signed(buffer_2_147); // @[Modules.scala 160:64:@8567.4]
  assign _T_62637 = _T_62636[13:0]; // @[Modules.scala 160:64:@8568.4]
  assign buffer_2_383 = $signed(_T_62637); // @[Modules.scala 160:64:@8569.4]
  assign buffer_2_148 = {{8{_T_61289[5]}},_T_61289}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_149 = {{8{_T_61296[5]}},_T_61296}; // @[Modules.scala 112:22:@8.4]
  assign _T_62639 = $signed(buffer_2_148) + $signed(buffer_2_149); // @[Modules.scala 160:64:@8571.4]
  assign _T_62640 = _T_62639[13:0]; // @[Modules.scala 160:64:@8572.4]
  assign buffer_2_384 = $signed(_T_62640); // @[Modules.scala 160:64:@8573.4]
  assign buffer_2_150 = {{8{_T_61303[5]}},_T_61303}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_151 = {{8{_T_61310[5]}},_T_61310}; // @[Modules.scala 112:22:@8.4]
  assign _T_62642 = $signed(buffer_2_150) + $signed(buffer_2_151); // @[Modules.scala 160:64:@8575.4]
  assign _T_62643 = _T_62642[13:0]; // @[Modules.scala 160:64:@8576.4]
  assign buffer_2_385 = $signed(_T_62643); // @[Modules.scala 160:64:@8577.4]
  assign buffer_2_152 = {{8{_T_61317[5]}},_T_61317}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_153 = {{9{_T_61324[4]}},_T_61324}; // @[Modules.scala 112:22:@8.4]
  assign _T_62645 = $signed(buffer_2_152) + $signed(buffer_2_153); // @[Modules.scala 160:64:@8579.4]
  assign _T_62646 = _T_62645[13:0]; // @[Modules.scala 160:64:@8580.4]
  assign buffer_2_386 = $signed(_T_62646); // @[Modules.scala 160:64:@8581.4]
  assign buffer_2_154 = {{8{_T_61331[5]}},_T_61331}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_155 = {{8{_T_61338[5]}},_T_61338}; // @[Modules.scala 112:22:@8.4]
  assign _T_62648 = $signed(buffer_2_154) + $signed(buffer_2_155); // @[Modules.scala 160:64:@8583.4]
  assign _T_62649 = _T_62648[13:0]; // @[Modules.scala 160:64:@8584.4]
  assign buffer_2_387 = $signed(_T_62649); // @[Modules.scala 160:64:@8585.4]
  assign buffer_2_156 = {{8{_T_61345[5]}},_T_61345}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_157 = {{8{_T_61352[5]}},_T_61352}; // @[Modules.scala 112:22:@8.4]
  assign _T_62651 = $signed(buffer_2_156) + $signed(buffer_2_157); // @[Modules.scala 160:64:@8587.4]
  assign _T_62652 = _T_62651[13:0]; // @[Modules.scala 160:64:@8588.4]
  assign buffer_2_388 = $signed(_T_62652); // @[Modules.scala 160:64:@8589.4]
  assign buffer_2_158 = {{8{_T_61359[5]}},_T_61359}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_159 = {{8{_T_61366[5]}},_T_61366}; // @[Modules.scala 112:22:@8.4]
  assign _T_62654 = $signed(buffer_2_158) + $signed(buffer_2_159); // @[Modules.scala 160:64:@8591.4]
  assign _T_62655 = _T_62654[13:0]; // @[Modules.scala 160:64:@8592.4]
  assign buffer_2_389 = $signed(_T_62655); // @[Modules.scala 160:64:@8593.4]
  assign buffer_2_160 = {{8{_T_61373[5]}},_T_61373}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_161 = {{8{_T_61380[5]}},_T_61380}; // @[Modules.scala 112:22:@8.4]
  assign _T_62657 = $signed(buffer_2_160) + $signed(buffer_2_161); // @[Modules.scala 160:64:@8595.4]
  assign _T_62658 = _T_62657[13:0]; // @[Modules.scala 160:64:@8596.4]
  assign buffer_2_390 = $signed(_T_62658); // @[Modules.scala 160:64:@8597.4]
  assign buffer_2_162 = {{8{_T_61387[5]}},_T_61387}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_163 = {{8{_T_61394[5]}},_T_61394}; // @[Modules.scala 112:22:@8.4]
  assign _T_62660 = $signed(buffer_2_162) + $signed(buffer_2_163); // @[Modules.scala 160:64:@8599.4]
  assign _T_62661 = _T_62660[13:0]; // @[Modules.scala 160:64:@8600.4]
  assign buffer_2_391 = $signed(_T_62661); // @[Modules.scala 160:64:@8601.4]
  assign buffer_2_164 = {{8{_T_61401[5]}},_T_61401}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_165 = {{8{_T_61408[5]}},_T_61408}; // @[Modules.scala 112:22:@8.4]
  assign _T_62663 = $signed(buffer_2_164) + $signed(buffer_2_165); // @[Modules.scala 160:64:@8603.4]
  assign _T_62664 = _T_62663[13:0]; // @[Modules.scala 160:64:@8604.4]
  assign buffer_2_392 = $signed(_T_62664); // @[Modules.scala 160:64:@8605.4]
  assign buffer_2_166 = {{9{_T_61415[4]}},_T_61415}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_167 = {{8{_T_61422[5]}},_T_61422}; // @[Modules.scala 112:22:@8.4]
  assign _T_62666 = $signed(buffer_2_166) + $signed(buffer_2_167); // @[Modules.scala 160:64:@8607.4]
  assign _T_62667 = _T_62666[13:0]; // @[Modules.scala 160:64:@8608.4]
  assign buffer_2_393 = $signed(_T_62667); // @[Modules.scala 160:64:@8609.4]
  assign buffer_2_168 = {{8{_T_61429[5]}},_T_61429}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_169 = {{8{_T_61436[5]}},_T_61436}; // @[Modules.scala 112:22:@8.4]
  assign _T_62669 = $signed(buffer_2_168) + $signed(buffer_2_169); // @[Modules.scala 160:64:@8611.4]
  assign _T_62670 = _T_62669[13:0]; // @[Modules.scala 160:64:@8612.4]
  assign buffer_2_394 = $signed(_T_62670); // @[Modules.scala 160:64:@8613.4]
  assign buffer_2_170 = {{8{_T_61443[5]}},_T_61443}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_171 = {{8{_T_61450[5]}},_T_61450}; // @[Modules.scala 112:22:@8.4]
  assign _T_62672 = $signed(buffer_2_170) + $signed(buffer_2_171); // @[Modules.scala 160:64:@8615.4]
  assign _T_62673 = _T_62672[13:0]; // @[Modules.scala 160:64:@8616.4]
  assign buffer_2_395 = $signed(_T_62673); // @[Modules.scala 160:64:@8617.4]
  assign buffer_2_172 = {{8{_T_61457[5]}},_T_61457}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_173 = {{8{_T_61464[5]}},_T_61464}; // @[Modules.scala 112:22:@8.4]
  assign _T_62675 = $signed(buffer_2_172) + $signed(buffer_2_173); // @[Modules.scala 160:64:@8619.4]
  assign _T_62676 = _T_62675[13:0]; // @[Modules.scala 160:64:@8620.4]
  assign buffer_2_396 = $signed(_T_62676); // @[Modules.scala 160:64:@8621.4]
  assign buffer_2_174 = {{8{_T_61471[5]}},_T_61471}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_175 = {{9{_T_61478[4]}},_T_61478}; // @[Modules.scala 112:22:@8.4]
  assign _T_62678 = $signed(buffer_2_174) + $signed(buffer_2_175); // @[Modules.scala 160:64:@8623.4]
  assign _T_62679 = _T_62678[13:0]; // @[Modules.scala 160:64:@8624.4]
  assign buffer_2_397 = $signed(_T_62679); // @[Modules.scala 160:64:@8625.4]
  assign buffer_2_176 = {{8{_T_61485[5]}},_T_61485}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_177 = {{8{_T_61492[5]}},_T_61492}; // @[Modules.scala 112:22:@8.4]
  assign _T_62681 = $signed(buffer_2_176) + $signed(buffer_2_177); // @[Modules.scala 160:64:@8627.4]
  assign _T_62682 = _T_62681[13:0]; // @[Modules.scala 160:64:@8628.4]
  assign buffer_2_398 = $signed(_T_62682); // @[Modules.scala 160:64:@8629.4]
  assign buffer_2_178 = {{9{_T_61499[4]}},_T_61499}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_179 = {{8{_T_61506[5]}},_T_61506}; // @[Modules.scala 112:22:@8.4]
  assign _T_62684 = $signed(buffer_2_178) + $signed(buffer_2_179); // @[Modules.scala 160:64:@8631.4]
  assign _T_62685 = _T_62684[13:0]; // @[Modules.scala 160:64:@8632.4]
  assign buffer_2_399 = $signed(_T_62685); // @[Modules.scala 160:64:@8633.4]
  assign buffer_2_180 = {{8{_T_61513[5]}},_T_61513}; // @[Modules.scala 112:22:@8.4]
  assign _T_62687 = $signed(buffer_2_180) + $signed(buffer_0_176); // @[Modules.scala 160:64:@8635.4]
  assign _T_62688 = _T_62687[13:0]; // @[Modules.scala 160:64:@8636.4]
  assign buffer_2_400 = $signed(_T_62688); // @[Modules.scala 160:64:@8637.4]
  assign buffer_2_182 = {{8{_T_61527[5]}},_T_61527}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_183 = {{8{_T_61534[5]}},_T_61534}; // @[Modules.scala 112:22:@8.4]
  assign _T_62690 = $signed(buffer_2_182) + $signed(buffer_2_183); // @[Modules.scala 160:64:@8639.4]
  assign _T_62691 = _T_62690[13:0]; // @[Modules.scala 160:64:@8640.4]
  assign buffer_2_401 = $signed(_T_62691); // @[Modules.scala 160:64:@8641.4]
  assign buffer_2_184 = {{8{_T_61541[5]}},_T_61541}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_185 = {{8{_T_61548[5]}},_T_61548}; // @[Modules.scala 112:22:@8.4]
  assign _T_62693 = $signed(buffer_2_184) + $signed(buffer_2_185); // @[Modules.scala 160:64:@8643.4]
  assign _T_62694 = _T_62693[13:0]; // @[Modules.scala 160:64:@8644.4]
  assign buffer_2_402 = $signed(_T_62694); // @[Modules.scala 160:64:@8645.4]
  assign buffer_2_186 = {{8{_T_61555[5]}},_T_61555}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_187 = {{8{_T_61562[5]}},_T_61562}; // @[Modules.scala 112:22:@8.4]
  assign _T_62696 = $signed(buffer_2_186) + $signed(buffer_2_187); // @[Modules.scala 160:64:@8647.4]
  assign _T_62697 = _T_62696[13:0]; // @[Modules.scala 160:64:@8648.4]
  assign buffer_2_403 = $signed(_T_62697); // @[Modules.scala 160:64:@8649.4]
  assign buffer_2_188 = {{9{_T_61569[4]}},_T_61569}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_189 = {{9{_T_61576[4]}},_T_61576}; // @[Modules.scala 112:22:@8.4]
  assign _T_62699 = $signed(buffer_2_188) + $signed(buffer_2_189); // @[Modules.scala 160:64:@8651.4]
  assign _T_62700 = _T_62699[13:0]; // @[Modules.scala 160:64:@8652.4]
  assign buffer_2_404 = $signed(_T_62700); // @[Modules.scala 160:64:@8653.4]
  assign buffer_2_190 = {{8{_T_61583[5]}},_T_61583}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_191 = {{9{_T_61590[4]}},_T_61590}; // @[Modules.scala 112:22:@8.4]
  assign _T_62702 = $signed(buffer_2_190) + $signed(buffer_2_191); // @[Modules.scala 160:64:@8655.4]
  assign _T_62703 = _T_62702[13:0]; // @[Modules.scala 160:64:@8656.4]
  assign buffer_2_405 = $signed(_T_62703); // @[Modules.scala 160:64:@8657.4]
  assign buffer_2_192 = {{9{_T_61597[4]}},_T_61597}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_193 = {{8{_T_61604[5]}},_T_61604}; // @[Modules.scala 112:22:@8.4]
  assign _T_62705 = $signed(buffer_2_192) + $signed(buffer_2_193); // @[Modules.scala 160:64:@8659.4]
  assign _T_62706 = _T_62705[13:0]; // @[Modules.scala 160:64:@8660.4]
  assign buffer_2_406 = $signed(_T_62706); // @[Modules.scala 160:64:@8661.4]
  assign buffer_2_194 = {{8{_T_61611[5]}},_T_61611}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_195 = {{8{_T_61618[5]}},_T_61618}; // @[Modules.scala 112:22:@8.4]
  assign _T_62708 = $signed(buffer_2_194) + $signed(buffer_2_195); // @[Modules.scala 160:64:@8663.4]
  assign _T_62709 = _T_62708[13:0]; // @[Modules.scala 160:64:@8664.4]
  assign buffer_2_407 = $signed(_T_62709); // @[Modules.scala 160:64:@8665.4]
  assign buffer_2_196 = {{8{_T_61625[5]}},_T_61625}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_197 = {{8{_T_61632[5]}},_T_61632}; // @[Modules.scala 112:22:@8.4]
  assign _T_62711 = $signed(buffer_2_196) + $signed(buffer_2_197); // @[Modules.scala 160:64:@8667.4]
  assign _T_62712 = _T_62711[13:0]; // @[Modules.scala 160:64:@8668.4]
  assign buffer_2_408 = $signed(_T_62712); // @[Modules.scala 160:64:@8669.4]
  assign buffer_2_198 = {{9{_T_61639[4]}},_T_61639}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_199 = {{9{_T_61646[4]}},_T_61646}; // @[Modules.scala 112:22:@8.4]
  assign _T_62714 = $signed(buffer_2_198) + $signed(buffer_2_199); // @[Modules.scala 160:64:@8671.4]
  assign _T_62715 = _T_62714[13:0]; // @[Modules.scala 160:64:@8672.4]
  assign buffer_2_409 = $signed(_T_62715); // @[Modules.scala 160:64:@8673.4]
  assign buffer_2_200 = {{8{_T_61653[5]}},_T_61653}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_201 = {{8{_T_61660[5]}},_T_61660}; // @[Modules.scala 112:22:@8.4]
  assign _T_62717 = $signed(buffer_2_200) + $signed(buffer_2_201); // @[Modules.scala 160:64:@8675.4]
  assign _T_62718 = _T_62717[13:0]; // @[Modules.scala 160:64:@8676.4]
  assign buffer_2_410 = $signed(_T_62718); // @[Modules.scala 160:64:@8677.4]
  assign buffer_2_202 = {{9{_T_61667[4]}},_T_61667}; // @[Modules.scala 112:22:@8.4]
  assign _T_62720 = $signed(buffer_2_202) + $signed(buffer_1_199); // @[Modules.scala 160:64:@8679.4]
  assign _T_62721 = _T_62720[13:0]; // @[Modules.scala 160:64:@8680.4]
  assign buffer_2_411 = $signed(_T_62721); // @[Modules.scala 160:64:@8681.4]
  assign buffer_2_204 = {{8{_T_61681[5]}},_T_61681}; // @[Modules.scala 112:22:@8.4]
  assign _T_62723 = $signed(buffer_2_204) + $signed(buffer_0_199); // @[Modules.scala 160:64:@8683.4]
  assign _T_62724 = _T_62723[13:0]; // @[Modules.scala 160:64:@8684.4]
  assign buffer_2_412 = $signed(_T_62724); // @[Modules.scala 160:64:@8685.4]
  assign buffer_2_207 = {{8{_T_61702[5]}},_T_61702}; // @[Modules.scala 112:22:@8.4]
  assign _T_62726 = $signed(buffer_0_200) + $signed(buffer_2_207); // @[Modules.scala 160:64:@8687.4]
  assign _T_62727 = _T_62726[13:0]; // @[Modules.scala 160:64:@8688.4]
  assign buffer_2_413 = $signed(_T_62727); // @[Modules.scala 160:64:@8689.4]
  assign buffer_2_208 = {{8{_T_61709[5]}},_T_61709}; // @[Modules.scala 112:22:@8.4]
  assign _T_62729 = $signed(buffer_2_208) + $signed(buffer_1_204); // @[Modules.scala 160:64:@8691.4]
  assign _T_62730 = _T_62729[13:0]; // @[Modules.scala 160:64:@8692.4]
  assign buffer_2_414 = $signed(_T_62730); // @[Modules.scala 160:64:@8693.4]
  assign buffer_2_211 = {{8{_T_61730[5]}},_T_61730}; // @[Modules.scala 112:22:@8.4]
  assign _T_62732 = $signed(buffer_1_205) + $signed(buffer_2_211); // @[Modules.scala 160:64:@8695.4]
  assign _T_62733 = _T_62732[13:0]; // @[Modules.scala 160:64:@8696.4]
  assign buffer_2_415 = $signed(_T_62733); // @[Modules.scala 160:64:@8697.4]
  assign buffer_2_212 = {{8{_T_61737[5]}},_T_61737}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_213 = {{9{_T_61744[4]}},_T_61744}; // @[Modules.scala 112:22:@8.4]
  assign _T_62735 = $signed(buffer_2_212) + $signed(buffer_2_213); // @[Modules.scala 160:64:@8699.4]
  assign _T_62736 = _T_62735[13:0]; // @[Modules.scala 160:64:@8700.4]
  assign buffer_2_416 = $signed(_T_62736); // @[Modules.scala 160:64:@8701.4]
  assign buffer_2_215 = {{9{_T_61758[4]}},_T_61758}; // @[Modules.scala 112:22:@8.4]
  assign _T_62738 = $signed(buffer_1_209) + $signed(buffer_2_215); // @[Modules.scala 160:64:@8703.4]
  assign _T_62739 = _T_62738[13:0]; // @[Modules.scala 160:64:@8704.4]
  assign buffer_2_417 = $signed(_T_62739); // @[Modules.scala 160:64:@8705.4]
  assign buffer_2_216 = {{8{_T_61765[5]}},_T_61765}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_217 = {{8{_T_61772[5]}},_T_61772}; // @[Modules.scala 112:22:@8.4]
  assign _T_62741 = $signed(buffer_2_216) + $signed(buffer_2_217); // @[Modules.scala 160:64:@8707.4]
  assign _T_62742 = _T_62741[13:0]; // @[Modules.scala 160:64:@8708.4]
  assign buffer_2_418 = $signed(_T_62742); // @[Modules.scala 160:64:@8709.4]
  assign buffer_2_218 = {{8{_T_61779[5]}},_T_61779}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_219 = {{8{_T_61786[5]}},_T_61786}; // @[Modules.scala 112:22:@8.4]
  assign _T_62744 = $signed(buffer_2_218) + $signed(buffer_2_219); // @[Modules.scala 160:64:@8711.4]
  assign _T_62745 = _T_62744[13:0]; // @[Modules.scala 160:64:@8712.4]
  assign buffer_2_419 = $signed(_T_62745); // @[Modules.scala 160:64:@8713.4]
  assign buffer_2_223 = {{8{_T_61814[5]}},_T_61814}; // @[Modules.scala 112:22:@8.4]
  assign _T_62750 = $signed(buffer_1_218) + $signed(buffer_2_223); // @[Modules.scala 160:64:@8719.4]
  assign _T_62751 = _T_62750[13:0]; // @[Modules.scala 160:64:@8720.4]
  assign buffer_2_421 = $signed(_T_62751); // @[Modules.scala 160:64:@8721.4]
  assign buffer_2_224 = {{9{_T_61821[4]}},_T_61821}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_225 = {{9{_T_61828[4]}},_T_61828}; // @[Modules.scala 112:22:@8.4]
  assign _T_62753 = $signed(buffer_2_224) + $signed(buffer_2_225); // @[Modules.scala 160:64:@8723.4]
  assign _T_62754 = _T_62753[13:0]; // @[Modules.scala 160:64:@8724.4]
  assign buffer_2_422 = $signed(_T_62754); // @[Modules.scala 160:64:@8725.4]
  assign buffer_2_226 = {{9{_T_61835[4]}},_T_61835}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_227 = {{9{_T_61842[4]}},_T_61842}; // @[Modules.scala 112:22:@8.4]
  assign _T_62756 = $signed(buffer_2_226) + $signed(buffer_2_227); // @[Modules.scala 160:64:@8727.4]
  assign _T_62757 = _T_62756[13:0]; // @[Modules.scala 160:64:@8728.4]
  assign buffer_2_423 = $signed(_T_62757); // @[Modules.scala 160:64:@8729.4]
  assign buffer_2_228 = {{8{_T_61849[5]}},_T_61849}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_229 = {{8{_T_61856[5]}},_T_61856}; // @[Modules.scala 112:22:@8.4]
  assign _T_62759 = $signed(buffer_2_228) + $signed(buffer_2_229); // @[Modules.scala 160:64:@8731.4]
  assign _T_62760 = _T_62759[13:0]; // @[Modules.scala 160:64:@8732.4]
  assign buffer_2_424 = $signed(_T_62760); // @[Modules.scala 160:64:@8733.4]
  assign buffer_2_230 = {{9{_T_61863[4]}},_T_61863}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_231 = {{9{_T_61870[4]}},_T_61870}; // @[Modules.scala 112:22:@8.4]
  assign _T_62762 = $signed(buffer_2_230) + $signed(buffer_2_231); // @[Modules.scala 160:64:@8735.4]
  assign _T_62763 = _T_62762[13:0]; // @[Modules.scala 160:64:@8736.4]
  assign buffer_2_425 = $signed(_T_62763); // @[Modules.scala 160:64:@8737.4]
  assign buffer_2_232 = {{8{_T_61877[5]}},_T_61877}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_233 = {{8{_T_61884[5]}},_T_61884}; // @[Modules.scala 112:22:@8.4]
  assign _T_62765 = $signed(buffer_2_232) + $signed(buffer_2_233); // @[Modules.scala 160:64:@8739.4]
  assign _T_62766 = _T_62765[13:0]; // @[Modules.scala 160:64:@8740.4]
  assign buffer_2_426 = $signed(_T_62766); // @[Modules.scala 160:64:@8741.4]
  assign buffer_2_234 = {{8{_T_61891[5]}},_T_61891}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_235 = {{8{_T_61898[5]}},_T_61898}; // @[Modules.scala 112:22:@8.4]
  assign _T_62768 = $signed(buffer_2_234) + $signed(buffer_2_235); // @[Modules.scala 160:64:@8743.4]
  assign _T_62769 = _T_62768[13:0]; // @[Modules.scala 160:64:@8744.4]
  assign buffer_2_427 = $signed(_T_62769); // @[Modules.scala 160:64:@8745.4]
  assign buffer_2_236 = {{9{_T_61905[4]}},_T_61905}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_237 = {{9{_T_61912[4]}},_T_61912}; // @[Modules.scala 112:22:@8.4]
  assign _T_62771 = $signed(buffer_2_236) + $signed(buffer_2_237); // @[Modules.scala 160:64:@8747.4]
  assign _T_62772 = _T_62771[13:0]; // @[Modules.scala 160:64:@8748.4]
  assign buffer_2_428 = $signed(_T_62772); // @[Modules.scala 160:64:@8749.4]
  assign buffer_2_238 = {{9{_T_61919[4]}},_T_61919}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_239 = {{8{_T_61926[5]}},_T_61926}; // @[Modules.scala 112:22:@8.4]
  assign _T_62774 = $signed(buffer_2_238) + $signed(buffer_2_239); // @[Modules.scala 160:64:@8751.4]
  assign _T_62775 = _T_62774[13:0]; // @[Modules.scala 160:64:@8752.4]
  assign buffer_2_429 = $signed(_T_62775); // @[Modules.scala 160:64:@8753.4]
  assign buffer_2_240 = {{8{_T_61933[5]}},_T_61933}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_241 = {{8{_T_61940[5]}},_T_61940}; // @[Modules.scala 112:22:@8.4]
  assign _T_62777 = $signed(buffer_2_240) + $signed(buffer_2_241); // @[Modules.scala 160:64:@8755.4]
  assign _T_62778 = _T_62777[13:0]; // @[Modules.scala 160:64:@8756.4]
  assign buffer_2_430 = $signed(_T_62778); // @[Modules.scala 160:64:@8757.4]
  assign buffer_2_242 = {{9{_T_61947[4]}},_T_61947}; // @[Modules.scala 112:22:@8.4]
  assign _T_62780 = $signed(buffer_2_242) + $signed(buffer_1_236); // @[Modules.scala 160:64:@8759.4]
  assign _T_62781 = _T_62780[13:0]; // @[Modules.scala 160:64:@8760.4]
  assign buffer_2_431 = $signed(_T_62781); // @[Modules.scala 160:64:@8761.4]
  assign buffer_2_244 = {{8{_T_61961[5]}},_T_61961}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_245 = {{8{_T_61968[5]}},_T_61968}; // @[Modules.scala 112:22:@8.4]
  assign _T_62783 = $signed(buffer_2_244) + $signed(buffer_2_245); // @[Modules.scala 160:64:@8763.4]
  assign _T_62784 = _T_62783[13:0]; // @[Modules.scala 160:64:@8764.4]
  assign buffer_2_432 = $signed(_T_62784); // @[Modules.scala 160:64:@8765.4]
  assign buffer_2_246 = {{8{_T_61975[5]}},_T_61975}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_247 = {{8{_T_61982[5]}},_T_61982}; // @[Modules.scala 112:22:@8.4]
  assign _T_62786 = $signed(buffer_2_246) + $signed(buffer_2_247); // @[Modules.scala 160:64:@8767.4]
  assign _T_62787 = _T_62786[13:0]; // @[Modules.scala 160:64:@8768.4]
  assign buffer_2_433 = $signed(_T_62787); // @[Modules.scala 160:64:@8769.4]
  assign buffer_2_248 = {{9{_T_61989[4]}},_T_61989}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_249 = {{9{_T_61996[4]}},_T_61996}; // @[Modules.scala 112:22:@8.4]
  assign _T_62789 = $signed(buffer_2_248) + $signed(buffer_2_249); // @[Modules.scala 160:64:@8771.4]
  assign _T_62790 = _T_62789[13:0]; // @[Modules.scala 160:64:@8772.4]
  assign buffer_2_434 = $signed(_T_62790); // @[Modules.scala 160:64:@8773.4]
  assign buffer_2_250 = {{9{_T_62003[4]}},_T_62003}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_251 = {{9{_T_62010[4]}},_T_62010}; // @[Modules.scala 112:22:@8.4]
  assign _T_62792 = $signed(buffer_2_250) + $signed(buffer_2_251); // @[Modules.scala 160:64:@8775.4]
  assign _T_62793 = _T_62792[13:0]; // @[Modules.scala 160:64:@8776.4]
  assign buffer_2_435 = $signed(_T_62793); // @[Modules.scala 160:64:@8777.4]
  assign buffer_2_252 = {{9{_T_62017[4]}},_T_62017}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_253 = {{9{_T_62024[4]}},_T_62024}; // @[Modules.scala 112:22:@8.4]
  assign _T_62795 = $signed(buffer_2_252) + $signed(buffer_2_253); // @[Modules.scala 160:64:@8779.4]
  assign _T_62796 = _T_62795[13:0]; // @[Modules.scala 160:64:@8780.4]
  assign buffer_2_436 = $signed(_T_62796); // @[Modules.scala 160:64:@8781.4]
  assign buffer_2_254 = {{8{_T_62031[5]}},_T_62031}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_255 = {{8{_T_62038[5]}},_T_62038}; // @[Modules.scala 112:22:@8.4]
  assign _T_62798 = $signed(buffer_2_254) + $signed(buffer_2_255); // @[Modules.scala 160:64:@8783.4]
  assign _T_62799 = _T_62798[13:0]; // @[Modules.scala 160:64:@8784.4]
  assign buffer_2_437 = $signed(_T_62799); // @[Modules.scala 160:64:@8785.4]
  assign buffer_2_257 = {{8{_T_62052[5]}},_T_62052}; // @[Modules.scala 112:22:@8.4]
  assign _T_62801 = $signed(buffer_0_249) + $signed(buffer_2_257); // @[Modules.scala 160:64:@8787.4]
  assign _T_62802 = _T_62801[13:0]; // @[Modules.scala 160:64:@8788.4]
  assign buffer_2_438 = $signed(_T_62802); // @[Modules.scala 160:64:@8789.4]
  assign buffer_2_258 = {{9{_T_62059[4]}},_T_62059}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_259 = {{9{_T_62066[4]}},_T_62066}; // @[Modules.scala 112:22:@8.4]
  assign _T_62804 = $signed(buffer_2_258) + $signed(buffer_2_259); // @[Modules.scala 160:64:@8791.4]
  assign _T_62805 = _T_62804[13:0]; // @[Modules.scala 160:64:@8792.4]
  assign buffer_2_439 = $signed(_T_62805); // @[Modules.scala 160:64:@8793.4]
  assign _T_62807 = $signed(buffer_0_253) + $signed(buffer_0_254); // @[Modules.scala 160:64:@8795.4]
  assign _T_62808 = _T_62807[13:0]; // @[Modules.scala 160:64:@8796.4]
  assign buffer_2_440 = $signed(_T_62808); // @[Modules.scala 160:64:@8797.4]
  assign _T_62810 = $signed(buffer_0_255) + $signed(buffer_0_256); // @[Modules.scala 160:64:@8799.4]
  assign _T_62811 = _T_62810[13:0]; // @[Modules.scala 160:64:@8800.4]
  assign buffer_2_441 = $signed(_T_62811); // @[Modules.scala 160:64:@8801.4]
  assign buffer_2_265 = {{8{_T_62108[5]}},_T_62108}; // @[Modules.scala 112:22:@8.4]
  assign _T_62813 = $signed(buffer_0_257) + $signed(buffer_2_265); // @[Modules.scala 160:64:@8803.4]
  assign _T_62814 = _T_62813[13:0]; // @[Modules.scala 160:64:@8804.4]
  assign buffer_2_442 = $signed(_T_62814); // @[Modules.scala 160:64:@8805.4]
  assign buffer_2_266 = {{8{_T_62115[5]}},_T_62115}; // @[Modules.scala 112:22:@8.4]
  assign _T_62816 = $signed(buffer_2_266) + $signed(buffer_1_258); // @[Modules.scala 160:64:@8807.4]
  assign _T_62817 = _T_62816[13:0]; // @[Modules.scala 160:64:@8808.4]
  assign buffer_2_443 = $signed(_T_62817); // @[Modules.scala 160:64:@8809.4]
  assign buffer_2_268 = {{9{_T_62129[4]}},_T_62129}; // @[Modules.scala 112:22:@8.4]
  assign _T_62819 = $signed(buffer_2_268) + $signed(buffer_1_260); // @[Modules.scala 160:64:@8811.4]
  assign _T_62820 = _T_62819[13:0]; // @[Modules.scala 160:64:@8812.4]
  assign buffer_2_444 = $signed(_T_62820); // @[Modules.scala 160:64:@8813.4]
  assign buffer_2_270 = {{9{_T_62143[4]}},_T_62143}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_271 = {{9{_T_62150[4]}},_T_62150}; // @[Modules.scala 112:22:@8.4]
  assign _T_62822 = $signed(buffer_2_270) + $signed(buffer_2_271); // @[Modules.scala 160:64:@8815.4]
  assign _T_62823 = _T_62822[13:0]; // @[Modules.scala 160:64:@8816.4]
  assign buffer_2_445 = $signed(_T_62823); // @[Modules.scala 160:64:@8817.4]
  assign buffer_2_272 = {{8{_T_62157[5]}},_T_62157}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_273 = {{8{_T_62164[5]}},_T_62164}; // @[Modules.scala 112:22:@8.4]
  assign _T_62825 = $signed(buffer_2_272) + $signed(buffer_2_273); // @[Modules.scala 160:64:@8819.4]
  assign _T_62826 = _T_62825[13:0]; // @[Modules.scala 160:64:@8820.4]
  assign buffer_2_446 = $signed(_T_62826); // @[Modules.scala 160:64:@8821.4]
  assign _T_62828 = $signed(buffer_0_266) + $signed(buffer_0_268); // @[Modules.scala 160:64:@8823.4]
  assign _T_62829 = _T_62828[13:0]; // @[Modules.scala 160:64:@8824.4]
  assign buffer_2_447 = $signed(_T_62829); // @[Modules.scala 160:64:@8825.4]
  assign buffer_2_276 = {{8{_T_62185[5]}},_T_62185}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_277 = {{8{_T_62192[5]}},_T_62192}; // @[Modules.scala 112:22:@8.4]
  assign _T_62831 = $signed(buffer_2_276) + $signed(buffer_2_277); // @[Modules.scala 160:64:@8827.4]
  assign _T_62832 = _T_62831[13:0]; // @[Modules.scala 160:64:@8828.4]
  assign buffer_2_448 = $signed(_T_62832); // @[Modules.scala 160:64:@8829.4]
  assign buffer_2_278 = {{8{_T_62199[5]}},_T_62199}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_279 = {{8{_T_62206[5]}},_T_62206}; // @[Modules.scala 112:22:@8.4]
  assign _T_62834 = $signed(buffer_2_278) + $signed(buffer_2_279); // @[Modules.scala 160:64:@8831.4]
  assign _T_62835 = _T_62834[13:0]; // @[Modules.scala 160:64:@8832.4]
  assign buffer_2_449 = $signed(_T_62835); // @[Modules.scala 160:64:@8833.4]
  assign buffer_2_280 = {{9{_T_62213[4]}},_T_62213}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_281 = {{8{_T_62220[5]}},_T_62220}; // @[Modules.scala 112:22:@8.4]
  assign _T_62837 = $signed(buffer_2_280) + $signed(buffer_2_281); // @[Modules.scala 160:64:@8835.4]
  assign _T_62838 = _T_62837[13:0]; // @[Modules.scala 160:64:@8836.4]
  assign buffer_2_450 = $signed(_T_62838); // @[Modules.scala 160:64:@8837.4]
  assign buffer_2_282 = {{8{_T_62227[5]}},_T_62227}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_283 = {{8{_T_62234[5]}},_T_62234}; // @[Modules.scala 112:22:@8.4]
  assign _T_62840 = $signed(buffer_2_282) + $signed(buffer_2_283); // @[Modules.scala 160:64:@8839.4]
  assign _T_62841 = _T_62840[13:0]; // @[Modules.scala 160:64:@8840.4]
  assign buffer_2_451 = $signed(_T_62841); // @[Modules.scala 160:64:@8841.4]
  assign buffer_2_284 = {{9{_T_62241[4]}},_T_62241}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_285 = {{9{_T_62248[4]}},_T_62248}; // @[Modules.scala 112:22:@8.4]
  assign _T_62843 = $signed(buffer_2_284) + $signed(buffer_2_285); // @[Modules.scala 160:64:@8843.4]
  assign _T_62844 = _T_62843[13:0]; // @[Modules.scala 160:64:@8844.4]
  assign buffer_2_452 = $signed(_T_62844); // @[Modules.scala 160:64:@8845.4]
  assign buffer_2_286 = {{8{_T_62255[5]}},_T_62255}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_287 = {{8{_T_62262[5]}},_T_62262}; // @[Modules.scala 112:22:@8.4]
  assign _T_62846 = $signed(buffer_2_286) + $signed(buffer_2_287); // @[Modules.scala 160:64:@8847.4]
  assign _T_62847 = _T_62846[13:0]; // @[Modules.scala 160:64:@8848.4]
  assign buffer_2_453 = $signed(_T_62847); // @[Modules.scala 160:64:@8849.4]
  assign buffer_2_289 = {{8{_T_62276[5]}},_T_62276}; // @[Modules.scala 112:22:@8.4]
  assign _T_62849 = $signed(buffer_0_283) + $signed(buffer_2_289); // @[Modules.scala 160:64:@8851.4]
  assign _T_62850 = _T_62849[13:0]; // @[Modules.scala 160:64:@8852.4]
  assign buffer_2_454 = $signed(_T_62850); // @[Modules.scala 160:64:@8853.4]
  assign buffer_2_290 = {{8{_T_62283[5]}},_T_62283}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_291 = {{8{_T_62290[5]}},_T_62290}; // @[Modules.scala 112:22:@8.4]
  assign _T_62852 = $signed(buffer_2_290) + $signed(buffer_2_291); // @[Modules.scala 160:64:@8855.4]
  assign _T_62853 = _T_62852[13:0]; // @[Modules.scala 160:64:@8856.4]
  assign buffer_2_455 = $signed(_T_62853); // @[Modules.scala 160:64:@8857.4]
  assign buffer_2_292 = {{8{_T_62297[5]}},_T_62297}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_293 = {{9{_T_62304[4]}},_T_62304}; // @[Modules.scala 112:22:@8.4]
  assign _T_62855 = $signed(buffer_2_292) + $signed(buffer_2_293); // @[Modules.scala 160:64:@8859.4]
  assign _T_62856 = _T_62855[13:0]; // @[Modules.scala 160:64:@8860.4]
  assign buffer_2_456 = $signed(_T_62856); // @[Modules.scala 160:64:@8861.4]
  assign buffer_2_294 = {{9{_T_62311[4]}},_T_62311}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_295 = {{9{_T_62318[4]}},_T_62318}; // @[Modules.scala 112:22:@8.4]
  assign _T_62858 = $signed(buffer_2_294) + $signed(buffer_2_295); // @[Modules.scala 160:64:@8863.4]
  assign _T_62859 = _T_62858[13:0]; // @[Modules.scala 160:64:@8864.4]
  assign buffer_2_457 = $signed(_T_62859); // @[Modules.scala 160:64:@8865.4]
  assign buffer_2_296 = {{9{_T_62325[4]}},_T_62325}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_297 = {{9{_T_62332[4]}},_T_62332}; // @[Modules.scala 112:22:@8.4]
  assign _T_62861 = $signed(buffer_2_296) + $signed(buffer_2_297); // @[Modules.scala 160:64:@8867.4]
  assign _T_62862 = _T_62861[13:0]; // @[Modules.scala 160:64:@8868.4]
  assign buffer_2_458 = $signed(_T_62862); // @[Modules.scala 160:64:@8869.4]
  assign buffer_2_298 = {{8{_T_62339[5]}},_T_62339}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_299 = {{9{_T_62346[4]}},_T_62346}; // @[Modules.scala 112:22:@8.4]
  assign _T_62864 = $signed(buffer_2_298) + $signed(buffer_2_299); // @[Modules.scala 160:64:@8871.4]
  assign _T_62865 = _T_62864[13:0]; // @[Modules.scala 160:64:@8872.4]
  assign buffer_2_459 = $signed(_T_62865); // @[Modules.scala 160:64:@8873.4]
  assign buffer_2_300 = {{9{_T_62353[4]}},_T_62353}; // @[Modules.scala 112:22:@8.4]
  assign _T_62867 = $signed(buffer_2_300) + $signed(buffer_0_293); // @[Modules.scala 160:64:@8875.4]
  assign _T_62868 = _T_62867[13:0]; // @[Modules.scala 160:64:@8876.4]
  assign buffer_2_460 = $signed(_T_62868); // @[Modules.scala 160:64:@8877.4]
  assign buffer_2_302 = {{9{_T_62367[4]}},_T_62367}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_303 = {{9{_T_62374[4]}},_T_62374}; // @[Modules.scala 112:22:@8.4]
  assign _T_62870 = $signed(buffer_2_302) + $signed(buffer_2_303); // @[Modules.scala 160:64:@8879.4]
  assign _T_62871 = _T_62870[13:0]; // @[Modules.scala 160:64:@8880.4]
  assign buffer_2_461 = $signed(_T_62871); // @[Modules.scala 160:64:@8881.4]
  assign buffer_2_304 = {{9{_T_62381[4]}},_T_62381}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_305 = {{9{_T_62388[4]}},_T_62388}; // @[Modules.scala 112:22:@8.4]
  assign _T_62873 = $signed(buffer_2_304) + $signed(buffer_2_305); // @[Modules.scala 160:64:@8883.4]
  assign _T_62874 = _T_62873[13:0]; // @[Modules.scala 160:64:@8884.4]
  assign buffer_2_462 = $signed(_T_62874); // @[Modules.scala 160:64:@8885.4]
  assign buffer_2_306 = {{9{_T_62395[4]}},_T_62395}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_307 = {{9{_T_62402[4]}},_T_62402}; // @[Modules.scala 112:22:@8.4]
  assign _T_62876 = $signed(buffer_2_306) + $signed(buffer_2_307); // @[Modules.scala 160:64:@8887.4]
  assign _T_62877 = _T_62876[13:0]; // @[Modules.scala 160:64:@8888.4]
  assign buffer_2_463 = $signed(_T_62877); // @[Modules.scala 160:64:@8889.4]
  assign buffer_2_308 = {{8{_T_62409[5]}},_T_62409}; // @[Modules.scala 112:22:@8.4]
  assign buffer_2_309 = {{8{_T_62416[5]}},_T_62416}; // @[Modules.scala 112:22:@8.4]
  assign _T_62879 = $signed(buffer_2_308) + $signed(buffer_2_309); // @[Modules.scala 160:64:@8891.4]
  assign _T_62880 = _T_62879[13:0]; // @[Modules.scala 160:64:@8892.4]
  assign buffer_2_464 = $signed(_T_62880); // @[Modules.scala 160:64:@8893.4]
  assign _T_62882 = $signed(buffer_2_310) + $signed(buffer_2_311); // @[Modules.scala 166:64:@8895.4]
  assign _T_62883 = _T_62882[13:0]; // @[Modules.scala 166:64:@8896.4]
  assign buffer_2_465 = $signed(_T_62883); // @[Modules.scala 166:64:@8897.4]
  assign _T_62885 = $signed(buffer_2_312) + $signed(buffer_2_313); // @[Modules.scala 166:64:@8899.4]
  assign _T_62886 = _T_62885[13:0]; // @[Modules.scala 166:64:@8900.4]
  assign buffer_2_466 = $signed(_T_62886); // @[Modules.scala 166:64:@8901.4]
  assign _T_62888 = $signed(buffer_2_314) + $signed(buffer_2_315); // @[Modules.scala 166:64:@8903.4]
  assign _T_62889 = _T_62888[13:0]; // @[Modules.scala 166:64:@8904.4]
  assign buffer_2_467 = $signed(_T_62889); // @[Modules.scala 166:64:@8905.4]
  assign _T_62891 = $signed(buffer_2_316) + $signed(buffer_2_317); // @[Modules.scala 166:64:@8907.4]
  assign _T_62892 = _T_62891[13:0]; // @[Modules.scala 166:64:@8908.4]
  assign buffer_2_468 = $signed(_T_62892); // @[Modules.scala 166:64:@8909.4]
  assign _T_62894 = $signed(buffer_2_318) + $signed(buffer_2_319); // @[Modules.scala 166:64:@8911.4]
  assign _T_62895 = _T_62894[13:0]; // @[Modules.scala 166:64:@8912.4]
  assign buffer_2_469 = $signed(_T_62895); // @[Modules.scala 166:64:@8913.4]
  assign _T_62897 = $signed(buffer_2_320) + $signed(buffer_2_321); // @[Modules.scala 166:64:@8915.4]
  assign _T_62898 = _T_62897[13:0]; // @[Modules.scala 166:64:@8916.4]
  assign buffer_2_470 = $signed(_T_62898); // @[Modules.scala 166:64:@8917.4]
  assign _T_62900 = $signed(buffer_2_322) + $signed(buffer_2_323); // @[Modules.scala 166:64:@8919.4]
  assign _T_62901 = _T_62900[13:0]; // @[Modules.scala 166:64:@8920.4]
  assign buffer_2_471 = $signed(_T_62901); // @[Modules.scala 166:64:@8921.4]
  assign _T_62903 = $signed(buffer_2_324) + $signed(buffer_2_325); // @[Modules.scala 166:64:@8923.4]
  assign _T_62904 = _T_62903[13:0]; // @[Modules.scala 166:64:@8924.4]
  assign buffer_2_472 = $signed(_T_62904); // @[Modules.scala 166:64:@8925.4]
  assign _T_62906 = $signed(buffer_2_326) + $signed(buffer_2_327); // @[Modules.scala 166:64:@8927.4]
  assign _T_62907 = _T_62906[13:0]; // @[Modules.scala 166:64:@8928.4]
  assign buffer_2_473 = $signed(_T_62907); // @[Modules.scala 166:64:@8929.4]
  assign _T_62909 = $signed(buffer_2_328) + $signed(buffer_2_329); // @[Modules.scala 166:64:@8931.4]
  assign _T_62910 = _T_62909[13:0]; // @[Modules.scala 166:64:@8932.4]
  assign buffer_2_474 = $signed(_T_62910); // @[Modules.scala 166:64:@8933.4]
  assign _T_62912 = $signed(buffer_2_330) + $signed(buffer_2_331); // @[Modules.scala 166:64:@8935.4]
  assign _T_62913 = _T_62912[13:0]; // @[Modules.scala 166:64:@8936.4]
  assign buffer_2_475 = $signed(_T_62913); // @[Modules.scala 166:64:@8937.4]
  assign _T_62915 = $signed(buffer_2_332) + $signed(buffer_2_333); // @[Modules.scala 166:64:@8939.4]
  assign _T_62916 = _T_62915[13:0]; // @[Modules.scala 166:64:@8940.4]
  assign buffer_2_476 = $signed(_T_62916); // @[Modules.scala 166:64:@8941.4]
  assign _T_62918 = $signed(buffer_2_334) + $signed(buffer_2_335); // @[Modules.scala 166:64:@8943.4]
  assign _T_62919 = _T_62918[13:0]; // @[Modules.scala 166:64:@8944.4]
  assign buffer_2_477 = $signed(_T_62919); // @[Modules.scala 166:64:@8945.4]
  assign _T_62921 = $signed(buffer_2_336) + $signed(buffer_2_337); // @[Modules.scala 166:64:@8947.4]
  assign _T_62922 = _T_62921[13:0]; // @[Modules.scala 166:64:@8948.4]
  assign buffer_2_478 = $signed(_T_62922); // @[Modules.scala 166:64:@8949.4]
  assign _T_62924 = $signed(buffer_2_338) + $signed(buffer_2_339); // @[Modules.scala 166:64:@8951.4]
  assign _T_62925 = _T_62924[13:0]; // @[Modules.scala 166:64:@8952.4]
  assign buffer_2_479 = $signed(_T_62925); // @[Modules.scala 166:64:@8953.4]
  assign _T_62927 = $signed(buffer_2_340) + $signed(buffer_2_341); // @[Modules.scala 166:64:@8955.4]
  assign _T_62928 = _T_62927[13:0]; // @[Modules.scala 166:64:@8956.4]
  assign buffer_2_480 = $signed(_T_62928); // @[Modules.scala 166:64:@8957.4]
  assign _T_62930 = $signed(buffer_2_342) + $signed(buffer_2_343); // @[Modules.scala 166:64:@8959.4]
  assign _T_62931 = _T_62930[13:0]; // @[Modules.scala 166:64:@8960.4]
  assign buffer_2_481 = $signed(_T_62931); // @[Modules.scala 166:64:@8961.4]
  assign _T_62933 = $signed(buffer_2_344) + $signed(buffer_2_345); // @[Modules.scala 166:64:@8963.4]
  assign _T_62934 = _T_62933[13:0]; // @[Modules.scala 166:64:@8964.4]
  assign buffer_2_482 = $signed(_T_62934); // @[Modules.scala 166:64:@8965.4]
  assign _T_62936 = $signed(buffer_2_346) + $signed(buffer_2_347); // @[Modules.scala 166:64:@8967.4]
  assign _T_62937 = _T_62936[13:0]; // @[Modules.scala 166:64:@8968.4]
  assign buffer_2_483 = $signed(_T_62937); // @[Modules.scala 166:64:@8969.4]
  assign _T_62939 = $signed(buffer_2_348) + $signed(buffer_1_343); // @[Modules.scala 166:64:@8971.4]
  assign _T_62940 = _T_62939[13:0]; // @[Modules.scala 166:64:@8972.4]
  assign buffer_2_484 = $signed(_T_62940); // @[Modules.scala 166:64:@8973.4]
  assign _T_62942 = $signed(buffer_2_350) + $signed(buffer_2_351); // @[Modules.scala 166:64:@8975.4]
  assign _T_62943 = _T_62942[13:0]; // @[Modules.scala 166:64:@8976.4]
  assign buffer_2_485 = $signed(_T_62943); // @[Modules.scala 166:64:@8977.4]
  assign _T_62945 = $signed(buffer_2_352) + $signed(buffer_2_353); // @[Modules.scala 166:64:@8979.4]
  assign _T_62946 = _T_62945[13:0]; // @[Modules.scala 166:64:@8980.4]
  assign buffer_2_486 = $signed(_T_62946); // @[Modules.scala 166:64:@8981.4]
  assign _T_62948 = $signed(buffer_2_354) + $signed(buffer_2_355); // @[Modules.scala 166:64:@8983.4]
  assign _T_62949 = _T_62948[13:0]; // @[Modules.scala 166:64:@8984.4]
  assign buffer_2_487 = $signed(_T_62949); // @[Modules.scala 166:64:@8985.4]
  assign _T_62951 = $signed(buffer_2_356) + $signed(buffer_2_357); // @[Modules.scala 166:64:@8987.4]
  assign _T_62952 = _T_62951[13:0]; // @[Modules.scala 166:64:@8988.4]
  assign buffer_2_488 = $signed(_T_62952); // @[Modules.scala 166:64:@8989.4]
  assign _T_62954 = $signed(buffer_2_358) + $signed(buffer_2_359); // @[Modules.scala 166:64:@8991.4]
  assign _T_62955 = _T_62954[13:0]; // @[Modules.scala 166:64:@8992.4]
  assign buffer_2_489 = $signed(_T_62955); // @[Modules.scala 166:64:@8993.4]
  assign _T_62957 = $signed(buffer_2_360) + $signed(buffer_1_354); // @[Modules.scala 166:64:@8995.4]
  assign _T_62958 = _T_62957[13:0]; // @[Modules.scala 166:64:@8996.4]
  assign buffer_2_490 = $signed(_T_62958); // @[Modules.scala 166:64:@8997.4]
  assign _T_62960 = $signed(buffer_2_362) + $signed(buffer_2_363); // @[Modules.scala 166:64:@8999.4]
  assign _T_62961 = _T_62960[13:0]; // @[Modules.scala 166:64:@9000.4]
  assign buffer_2_491 = $signed(_T_62961); // @[Modules.scala 166:64:@9001.4]
  assign _T_62963 = $signed(buffer_2_364) + $signed(buffer_2_365); // @[Modules.scala 166:64:@9003.4]
  assign _T_62964 = _T_62963[13:0]; // @[Modules.scala 166:64:@9004.4]
  assign buffer_2_492 = $signed(_T_62964); // @[Modules.scala 166:64:@9005.4]
  assign _T_62966 = $signed(buffer_2_366) + $signed(buffer_1_360); // @[Modules.scala 166:64:@9007.4]
  assign _T_62967 = _T_62966[13:0]; // @[Modules.scala 166:64:@9008.4]
  assign buffer_2_493 = $signed(_T_62967); // @[Modules.scala 166:64:@9009.4]
  assign _T_62969 = $signed(buffer_2_368) + $signed(buffer_2_369); // @[Modules.scala 166:64:@9011.4]
  assign _T_62970 = _T_62969[13:0]; // @[Modules.scala 166:64:@9012.4]
  assign buffer_2_494 = $signed(_T_62970); // @[Modules.scala 166:64:@9013.4]
  assign _T_62972 = $signed(buffer_2_370) + $signed(buffer_2_371); // @[Modules.scala 166:64:@9015.4]
  assign _T_62973 = _T_62972[13:0]; // @[Modules.scala 166:64:@9016.4]
  assign buffer_2_495 = $signed(_T_62973); // @[Modules.scala 166:64:@9017.4]
  assign _T_62975 = $signed(buffer_2_372) + $signed(buffer_2_373); // @[Modules.scala 166:64:@9019.4]
  assign _T_62976 = _T_62975[13:0]; // @[Modules.scala 166:64:@9020.4]
  assign buffer_2_496 = $signed(_T_62976); // @[Modules.scala 166:64:@9021.4]
  assign _T_62978 = $signed(buffer_2_374) + $signed(buffer_2_375); // @[Modules.scala 166:64:@9023.4]
  assign _T_62979 = _T_62978[13:0]; // @[Modules.scala 166:64:@9024.4]
  assign buffer_2_497 = $signed(_T_62979); // @[Modules.scala 166:64:@9025.4]
  assign _T_62981 = $signed(buffer_2_376) + $signed(buffer_2_377); // @[Modules.scala 166:64:@9027.4]
  assign _T_62982 = _T_62981[13:0]; // @[Modules.scala 166:64:@9028.4]
  assign buffer_2_498 = $signed(_T_62982); // @[Modules.scala 166:64:@9029.4]
  assign _T_62984 = $signed(buffer_2_378) + $signed(buffer_2_379); // @[Modules.scala 166:64:@9031.4]
  assign _T_62985 = _T_62984[13:0]; // @[Modules.scala 166:64:@9032.4]
  assign buffer_2_499 = $signed(_T_62985); // @[Modules.scala 166:64:@9033.4]
  assign _T_62987 = $signed(buffer_2_380) + $signed(buffer_2_381); // @[Modules.scala 166:64:@9035.4]
  assign _T_62988 = _T_62987[13:0]; // @[Modules.scala 166:64:@9036.4]
  assign buffer_2_500 = $signed(_T_62988); // @[Modules.scala 166:64:@9037.4]
  assign _T_62990 = $signed(buffer_2_382) + $signed(buffer_2_383); // @[Modules.scala 166:64:@9039.4]
  assign _T_62991 = _T_62990[13:0]; // @[Modules.scala 166:64:@9040.4]
  assign buffer_2_501 = $signed(_T_62991); // @[Modules.scala 166:64:@9041.4]
  assign _T_62993 = $signed(buffer_2_384) + $signed(buffer_2_385); // @[Modules.scala 166:64:@9043.4]
  assign _T_62994 = _T_62993[13:0]; // @[Modules.scala 166:64:@9044.4]
  assign buffer_2_502 = $signed(_T_62994); // @[Modules.scala 166:64:@9045.4]
  assign _T_62996 = $signed(buffer_2_386) + $signed(buffer_2_387); // @[Modules.scala 166:64:@9047.4]
  assign _T_62997 = _T_62996[13:0]; // @[Modules.scala 166:64:@9048.4]
  assign buffer_2_503 = $signed(_T_62997); // @[Modules.scala 166:64:@9049.4]
  assign _T_62999 = $signed(buffer_2_388) + $signed(buffer_2_389); // @[Modules.scala 166:64:@9051.4]
  assign _T_63000 = _T_62999[13:0]; // @[Modules.scala 166:64:@9052.4]
  assign buffer_2_504 = $signed(_T_63000); // @[Modules.scala 166:64:@9053.4]
  assign _T_63002 = $signed(buffer_2_390) + $signed(buffer_2_391); // @[Modules.scala 166:64:@9055.4]
  assign _T_63003 = _T_63002[13:0]; // @[Modules.scala 166:64:@9056.4]
  assign buffer_2_505 = $signed(_T_63003); // @[Modules.scala 166:64:@9057.4]
  assign _T_63005 = $signed(buffer_2_392) + $signed(buffer_2_393); // @[Modules.scala 166:64:@9059.4]
  assign _T_63006 = _T_63005[13:0]; // @[Modules.scala 166:64:@9060.4]
  assign buffer_2_506 = $signed(_T_63006); // @[Modules.scala 166:64:@9061.4]
  assign _T_63008 = $signed(buffer_2_394) + $signed(buffer_2_395); // @[Modules.scala 166:64:@9063.4]
  assign _T_63009 = _T_63008[13:0]; // @[Modules.scala 166:64:@9064.4]
  assign buffer_2_507 = $signed(_T_63009); // @[Modules.scala 166:64:@9065.4]
  assign _T_63011 = $signed(buffer_2_396) + $signed(buffer_2_397); // @[Modules.scala 166:64:@9067.4]
  assign _T_63012 = _T_63011[13:0]; // @[Modules.scala 166:64:@9068.4]
  assign buffer_2_508 = $signed(_T_63012); // @[Modules.scala 166:64:@9069.4]
  assign _T_63014 = $signed(buffer_2_398) + $signed(buffer_2_399); // @[Modules.scala 166:64:@9071.4]
  assign _T_63015 = _T_63014[13:0]; // @[Modules.scala 166:64:@9072.4]
  assign buffer_2_509 = $signed(_T_63015); // @[Modules.scala 166:64:@9073.4]
  assign _T_63017 = $signed(buffer_2_400) + $signed(buffer_2_401); // @[Modules.scala 166:64:@9075.4]
  assign _T_63018 = _T_63017[13:0]; // @[Modules.scala 166:64:@9076.4]
  assign buffer_2_510 = $signed(_T_63018); // @[Modules.scala 166:64:@9077.4]
  assign _T_63020 = $signed(buffer_2_402) + $signed(buffer_2_403); // @[Modules.scala 166:64:@9079.4]
  assign _T_63021 = _T_63020[13:0]; // @[Modules.scala 166:64:@9080.4]
  assign buffer_2_511 = $signed(_T_63021); // @[Modules.scala 166:64:@9081.4]
  assign _T_63023 = $signed(buffer_2_404) + $signed(buffer_2_405); // @[Modules.scala 166:64:@9083.4]
  assign _T_63024 = _T_63023[13:0]; // @[Modules.scala 166:64:@9084.4]
  assign buffer_2_512 = $signed(_T_63024); // @[Modules.scala 166:64:@9085.4]
  assign _T_63026 = $signed(buffer_2_406) + $signed(buffer_2_407); // @[Modules.scala 166:64:@9087.4]
  assign _T_63027 = _T_63026[13:0]; // @[Modules.scala 166:64:@9088.4]
  assign buffer_2_513 = $signed(_T_63027); // @[Modules.scala 166:64:@9089.4]
  assign _T_63029 = $signed(buffer_2_408) + $signed(buffer_2_409); // @[Modules.scala 166:64:@9091.4]
  assign _T_63030 = _T_63029[13:0]; // @[Modules.scala 166:64:@9092.4]
  assign buffer_2_514 = $signed(_T_63030); // @[Modules.scala 166:64:@9093.4]
  assign _T_63032 = $signed(buffer_2_410) + $signed(buffer_2_411); // @[Modules.scala 166:64:@9095.4]
  assign _T_63033 = _T_63032[13:0]; // @[Modules.scala 166:64:@9096.4]
  assign buffer_2_515 = $signed(_T_63033); // @[Modules.scala 166:64:@9097.4]
  assign _T_63035 = $signed(buffer_2_412) + $signed(buffer_2_413); // @[Modules.scala 166:64:@9099.4]
  assign _T_63036 = _T_63035[13:0]; // @[Modules.scala 166:64:@9100.4]
  assign buffer_2_516 = $signed(_T_63036); // @[Modules.scala 166:64:@9101.4]
  assign _T_63038 = $signed(buffer_2_414) + $signed(buffer_2_415); // @[Modules.scala 166:64:@9103.4]
  assign _T_63039 = _T_63038[13:0]; // @[Modules.scala 166:64:@9104.4]
  assign buffer_2_517 = $signed(_T_63039); // @[Modules.scala 166:64:@9105.4]
  assign _T_63041 = $signed(buffer_2_416) + $signed(buffer_2_417); // @[Modules.scala 166:64:@9107.4]
  assign _T_63042 = _T_63041[13:0]; // @[Modules.scala 166:64:@9108.4]
  assign buffer_2_518 = $signed(_T_63042); // @[Modules.scala 166:64:@9109.4]
  assign _T_63044 = $signed(buffer_2_418) + $signed(buffer_2_419); // @[Modules.scala 166:64:@9111.4]
  assign _T_63045 = _T_63044[13:0]; // @[Modules.scala 166:64:@9112.4]
  assign buffer_2_519 = $signed(_T_63045); // @[Modules.scala 166:64:@9113.4]
  assign _T_63047 = $signed(buffer_1_412) + $signed(buffer_2_421); // @[Modules.scala 166:64:@9115.4]
  assign _T_63048 = _T_63047[13:0]; // @[Modules.scala 166:64:@9116.4]
  assign buffer_2_520 = $signed(_T_63048); // @[Modules.scala 166:64:@9117.4]
  assign _T_63050 = $signed(buffer_2_422) + $signed(buffer_2_423); // @[Modules.scala 166:64:@9119.4]
  assign _T_63051 = _T_63050[13:0]; // @[Modules.scala 166:64:@9120.4]
  assign buffer_2_521 = $signed(_T_63051); // @[Modules.scala 166:64:@9121.4]
  assign _T_63053 = $signed(buffer_2_424) + $signed(buffer_2_425); // @[Modules.scala 166:64:@9123.4]
  assign _T_63054 = _T_63053[13:0]; // @[Modules.scala 166:64:@9124.4]
  assign buffer_2_522 = $signed(_T_63054); // @[Modules.scala 166:64:@9125.4]
  assign _T_63056 = $signed(buffer_2_426) + $signed(buffer_2_427); // @[Modules.scala 166:64:@9127.4]
  assign _T_63057 = _T_63056[13:0]; // @[Modules.scala 166:64:@9128.4]
  assign buffer_2_523 = $signed(_T_63057); // @[Modules.scala 166:64:@9129.4]
  assign _T_63059 = $signed(buffer_2_428) + $signed(buffer_2_429); // @[Modules.scala 166:64:@9131.4]
  assign _T_63060 = _T_63059[13:0]; // @[Modules.scala 166:64:@9132.4]
  assign buffer_2_524 = $signed(_T_63060); // @[Modules.scala 166:64:@9133.4]
  assign _T_63062 = $signed(buffer_2_430) + $signed(buffer_2_431); // @[Modules.scala 166:64:@9135.4]
  assign _T_63063 = _T_63062[13:0]; // @[Modules.scala 166:64:@9136.4]
  assign buffer_2_525 = $signed(_T_63063); // @[Modules.scala 166:64:@9137.4]
  assign _T_63065 = $signed(buffer_2_432) + $signed(buffer_2_433); // @[Modules.scala 166:64:@9139.4]
  assign _T_63066 = _T_63065[13:0]; // @[Modules.scala 166:64:@9140.4]
  assign buffer_2_526 = $signed(_T_63066); // @[Modules.scala 166:64:@9141.4]
  assign _T_63068 = $signed(buffer_2_434) + $signed(buffer_2_435); // @[Modules.scala 166:64:@9143.4]
  assign _T_63069 = _T_63068[13:0]; // @[Modules.scala 166:64:@9144.4]
  assign buffer_2_527 = $signed(_T_63069); // @[Modules.scala 166:64:@9145.4]
  assign _T_63071 = $signed(buffer_2_436) + $signed(buffer_2_437); // @[Modules.scala 166:64:@9147.4]
  assign _T_63072 = _T_63071[13:0]; // @[Modules.scala 166:64:@9148.4]
  assign buffer_2_528 = $signed(_T_63072); // @[Modules.scala 166:64:@9149.4]
  assign _T_63074 = $signed(buffer_2_438) + $signed(buffer_2_439); // @[Modules.scala 166:64:@9151.4]
  assign _T_63075 = _T_63074[13:0]; // @[Modules.scala 166:64:@9152.4]
  assign buffer_2_529 = $signed(_T_63075); // @[Modules.scala 166:64:@9153.4]
  assign _T_63077 = $signed(buffer_2_440) + $signed(buffer_2_441); // @[Modules.scala 166:64:@9155.4]
  assign _T_63078 = _T_63077[13:0]; // @[Modules.scala 166:64:@9156.4]
  assign buffer_2_530 = $signed(_T_63078); // @[Modules.scala 166:64:@9157.4]
  assign _T_63080 = $signed(buffer_2_442) + $signed(buffer_2_443); // @[Modules.scala 166:64:@9159.4]
  assign _T_63081 = _T_63080[13:0]; // @[Modules.scala 166:64:@9160.4]
  assign buffer_2_531 = $signed(_T_63081); // @[Modules.scala 166:64:@9161.4]
  assign _T_63083 = $signed(buffer_2_444) + $signed(buffer_2_445); // @[Modules.scala 166:64:@9163.4]
  assign _T_63084 = _T_63083[13:0]; // @[Modules.scala 166:64:@9164.4]
  assign buffer_2_532 = $signed(_T_63084); // @[Modules.scala 166:64:@9165.4]
  assign _T_63086 = $signed(buffer_2_446) + $signed(buffer_2_447); // @[Modules.scala 166:64:@9167.4]
  assign _T_63087 = _T_63086[13:0]; // @[Modules.scala 166:64:@9168.4]
  assign buffer_2_533 = $signed(_T_63087); // @[Modules.scala 166:64:@9169.4]
  assign _T_63089 = $signed(buffer_2_448) + $signed(buffer_2_449); // @[Modules.scala 166:64:@9171.4]
  assign _T_63090 = _T_63089[13:0]; // @[Modules.scala 166:64:@9172.4]
  assign buffer_2_534 = $signed(_T_63090); // @[Modules.scala 166:64:@9173.4]
  assign _T_63092 = $signed(buffer_2_450) + $signed(buffer_2_451); // @[Modules.scala 166:64:@9175.4]
  assign _T_63093 = _T_63092[13:0]; // @[Modules.scala 166:64:@9176.4]
  assign buffer_2_535 = $signed(_T_63093); // @[Modules.scala 166:64:@9177.4]
  assign _T_63095 = $signed(buffer_2_452) + $signed(buffer_2_453); // @[Modules.scala 166:64:@9179.4]
  assign _T_63096 = _T_63095[13:0]; // @[Modules.scala 166:64:@9180.4]
  assign buffer_2_536 = $signed(_T_63096); // @[Modules.scala 166:64:@9181.4]
  assign _T_63098 = $signed(buffer_2_454) + $signed(buffer_2_455); // @[Modules.scala 166:64:@9183.4]
  assign _T_63099 = _T_63098[13:0]; // @[Modules.scala 166:64:@9184.4]
  assign buffer_2_537 = $signed(_T_63099); // @[Modules.scala 166:64:@9185.4]
  assign _T_63101 = $signed(buffer_2_456) + $signed(buffer_2_457); // @[Modules.scala 166:64:@9187.4]
  assign _T_63102 = _T_63101[13:0]; // @[Modules.scala 166:64:@9188.4]
  assign buffer_2_538 = $signed(_T_63102); // @[Modules.scala 166:64:@9189.4]
  assign _T_63104 = $signed(buffer_2_458) + $signed(buffer_2_459); // @[Modules.scala 166:64:@9191.4]
  assign _T_63105 = _T_63104[13:0]; // @[Modules.scala 166:64:@9192.4]
  assign buffer_2_539 = $signed(_T_63105); // @[Modules.scala 166:64:@9193.4]
  assign _T_63107 = $signed(buffer_2_460) + $signed(buffer_2_461); // @[Modules.scala 166:64:@9195.4]
  assign _T_63108 = _T_63107[13:0]; // @[Modules.scala 166:64:@9196.4]
  assign buffer_2_540 = $signed(_T_63108); // @[Modules.scala 166:64:@9197.4]
  assign _T_63110 = $signed(buffer_2_462) + $signed(buffer_2_463); // @[Modules.scala 166:64:@9199.4]
  assign _T_63111 = _T_63110[13:0]; // @[Modules.scala 166:64:@9200.4]
  assign buffer_2_541 = $signed(_T_63111); // @[Modules.scala 166:64:@9201.4]
  assign _T_63113 = $signed(buffer_2_465) + $signed(buffer_2_466); // @[Modules.scala 166:64:@9203.4]
  assign _T_63114 = _T_63113[13:0]; // @[Modules.scala 166:64:@9204.4]
  assign buffer_2_542 = $signed(_T_63114); // @[Modules.scala 166:64:@9205.4]
  assign _T_63116 = $signed(buffer_2_467) + $signed(buffer_2_468); // @[Modules.scala 166:64:@9207.4]
  assign _T_63117 = _T_63116[13:0]; // @[Modules.scala 166:64:@9208.4]
  assign buffer_2_543 = $signed(_T_63117); // @[Modules.scala 166:64:@9209.4]
  assign _T_63119 = $signed(buffer_2_469) + $signed(buffer_2_470); // @[Modules.scala 166:64:@9211.4]
  assign _T_63120 = _T_63119[13:0]; // @[Modules.scala 166:64:@9212.4]
  assign buffer_2_544 = $signed(_T_63120); // @[Modules.scala 166:64:@9213.4]
  assign _T_63122 = $signed(buffer_2_471) + $signed(buffer_2_472); // @[Modules.scala 166:64:@9215.4]
  assign _T_63123 = _T_63122[13:0]; // @[Modules.scala 166:64:@9216.4]
  assign buffer_2_545 = $signed(_T_63123); // @[Modules.scala 166:64:@9217.4]
  assign _T_63125 = $signed(buffer_2_473) + $signed(buffer_2_474); // @[Modules.scala 166:64:@9219.4]
  assign _T_63126 = _T_63125[13:0]; // @[Modules.scala 166:64:@9220.4]
  assign buffer_2_546 = $signed(_T_63126); // @[Modules.scala 166:64:@9221.4]
  assign _T_63128 = $signed(buffer_2_475) + $signed(buffer_2_476); // @[Modules.scala 166:64:@9223.4]
  assign _T_63129 = _T_63128[13:0]; // @[Modules.scala 166:64:@9224.4]
  assign buffer_2_547 = $signed(_T_63129); // @[Modules.scala 166:64:@9225.4]
  assign _T_63131 = $signed(buffer_2_477) + $signed(buffer_2_478); // @[Modules.scala 166:64:@9227.4]
  assign _T_63132 = _T_63131[13:0]; // @[Modules.scala 166:64:@9228.4]
  assign buffer_2_548 = $signed(_T_63132); // @[Modules.scala 166:64:@9229.4]
  assign _T_63134 = $signed(buffer_2_479) + $signed(buffer_2_480); // @[Modules.scala 166:64:@9231.4]
  assign _T_63135 = _T_63134[13:0]; // @[Modules.scala 166:64:@9232.4]
  assign buffer_2_549 = $signed(_T_63135); // @[Modules.scala 166:64:@9233.4]
  assign _T_63137 = $signed(buffer_2_481) + $signed(buffer_2_482); // @[Modules.scala 166:64:@9235.4]
  assign _T_63138 = _T_63137[13:0]; // @[Modules.scala 166:64:@9236.4]
  assign buffer_2_550 = $signed(_T_63138); // @[Modules.scala 166:64:@9237.4]
  assign _T_63140 = $signed(buffer_2_483) + $signed(buffer_2_484); // @[Modules.scala 166:64:@9239.4]
  assign _T_63141 = _T_63140[13:0]; // @[Modules.scala 166:64:@9240.4]
  assign buffer_2_551 = $signed(_T_63141); // @[Modules.scala 166:64:@9241.4]
  assign _T_63143 = $signed(buffer_2_485) + $signed(buffer_2_486); // @[Modules.scala 166:64:@9243.4]
  assign _T_63144 = _T_63143[13:0]; // @[Modules.scala 166:64:@9244.4]
  assign buffer_2_552 = $signed(_T_63144); // @[Modules.scala 166:64:@9245.4]
  assign _T_63146 = $signed(buffer_2_487) + $signed(buffer_2_488); // @[Modules.scala 166:64:@9247.4]
  assign _T_63147 = _T_63146[13:0]; // @[Modules.scala 166:64:@9248.4]
  assign buffer_2_553 = $signed(_T_63147); // @[Modules.scala 166:64:@9249.4]
  assign _T_63149 = $signed(buffer_2_489) + $signed(buffer_2_490); // @[Modules.scala 166:64:@9251.4]
  assign _T_63150 = _T_63149[13:0]; // @[Modules.scala 166:64:@9252.4]
  assign buffer_2_554 = $signed(_T_63150); // @[Modules.scala 166:64:@9253.4]
  assign _T_63152 = $signed(buffer_2_491) + $signed(buffer_2_492); // @[Modules.scala 166:64:@9255.4]
  assign _T_63153 = _T_63152[13:0]; // @[Modules.scala 166:64:@9256.4]
  assign buffer_2_555 = $signed(_T_63153); // @[Modules.scala 166:64:@9257.4]
  assign _T_63155 = $signed(buffer_2_493) + $signed(buffer_2_494); // @[Modules.scala 166:64:@9259.4]
  assign _T_63156 = _T_63155[13:0]; // @[Modules.scala 166:64:@9260.4]
  assign buffer_2_556 = $signed(_T_63156); // @[Modules.scala 166:64:@9261.4]
  assign _T_63158 = $signed(buffer_2_495) + $signed(buffer_2_496); // @[Modules.scala 166:64:@9263.4]
  assign _T_63159 = _T_63158[13:0]; // @[Modules.scala 166:64:@9264.4]
  assign buffer_2_557 = $signed(_T_63159); // @[Modules.scala 166:64:@9265.4]
  assign _T_63161 = $signed(buffer_2_497) + $signed(buffer_2_498); // @[Modules.scala 166:64:@9267.4]
  assign _T_63162 = _T_63161[13:0]; // @[Modules.scala 166:64:@9268.4]
  assign buffer_2_558 = $signed(_T_63162); // @[Modules.scala 166:64:@9269.4]
  assign _T_63164 = $signed(buffer_2_499) + $signed(buffer_2_500); // @[Modules.scala 166:64:@9271.4]
  assign _T_63165 = _T_63164[13:0]; // @[Modules.scala 166:64:@9272.4]
  assign buffer_2_559 = $signed(_T_63165); // @[Modules.scala 166:64:@9273.4]
  assign _T_63167 = $signed(buffer_2_501) + $signed(buffer_2_502); // @[Modules.scala 166:64:@9275.4]
  assign _T_63168 = _T_63167[13:0]; // @[Modules.scala 166:64:@9276.4]
  assign buffer_2_560 = $signed(_T_63168); // @[Modules.scala 166:64:@9277.4]
  assign _T_63170 = $signed(buffer_2_503) + $signed(buffer_2_504); // @[Modules.scala 166:64:@9279.4]
  assign _T_63171 = _T_63170[13:0]; // @[Modules.scala 166:64:@9280.4]
  assign buffer_2_561 = $signed(_T_63171); // @[Modules.scala 166:64:@9281.4]
  assign _T_63173 = $signed(buffer_2_505) + $signed(buffer_2_506); // @[Modules.scala 166:64:@9283.4]
  assign _T_63174 = _T_63173[13:0]; // @[Modules.scala 166:64:@9284.4]
  assign buffer_2_562 = $signed(_T_63174); // @[Modules.scala 166:64:@9285.4]
  assign _T_63176 = $signed(buffer_2_507) + $signed(buffer_2_508); // @[Modules.scala 166:64:@9287.4]
  assign _T_63177 = _T_63176[13:0]; // @[Modules.scala 166:64:@9288.4]
  assign buffer_2_563 = $signed(_T_63177); // @[Modules.scala 166:64:@9289.4]
  assign _T_63179 = $signed(buffer_2_509) + $signed(buffer_2_510); // @[Modules.scala 166:64:@9291.4]
  assign _T_63180 = _T_63179[13:0]; // @[Modules.scala 166:64:@9292.4]
  assign buffer_2_564 = $signed(_T_63180); // @[Modules.scala 166:64:@9293.4]
  assign _T_63182 = $signed(buffer_2_511) + $signed(buffer_2_512); // @[Modules.scala 166:64:@9295.4]
  assign _T_63183 = _T_63182[13:0]; // @[Modules.scala 166:64:@9296.4]
  assign buffer_2_565 = $signed(_T_63183); // @[Modules.scala 166:64:@9297.4]
  assign _T_63185 = $signed(buffer_2_513) + $signed(buffer_2_514); // @[Modules.scala 166:64:@9299.4]
  assign _T_63186 = _T_63185[13:0]; // @[Modules.scala 166:64:@9300.4]
  assign buffer_2_566 = $signed(_T_63186); // @[Modules.scala 166:64:@9301.4]
  assign _T_63188 = $signed(buffer_2_515) + $signed(buffer_2_516); // @[Modules.scala 166:64:@9303.4]
  assign _T_63189 = _T_63188[13:0]; // @[Modules.scala 166:64:@9304.4]
  assign buffer_2_567 = $signed(_T_63189); // @[Modules.scala 166:64:@9305.4]
  assign _T_63191 = $signed(buffer_2_517) + $signed(buffer_2_518); // @[Modules.scala 166:64:@9307.4]
  assign _T_63192 = _T_63191[13:0]; // @[Modules.scala 166:64:@9308.4]
  assign buffer_2_568 = $signed(_T_63192); // @[Modules.scala 166:64:@9309.4]
  assign _T_63194 = $signed(buffer_2_519) + $signed(buffer_2_520); // @[Modules.scala 166:64:@9311.4]
  assign _T_63195 = _T_63194[13:0]; // @[Modules.scala 166:64:@9312.4]
  assign buffer_2_569 = $signed(_T_63195); // @[Modules.scala 166:64:@9313.4]
  assign _T_63197 = $signed(buffer_2_521) + $signed(buffer_2_522); // @[Modules.scala 166:64:@9315.4]
  assign _T_63198 = _T_63197[13:0]; // @[Modules.scala 166:64:@9316.4]
  assign buffer_2_570 = $signed(_T_63198); // @[Modules.scala 166:64:@9317.4]
  assign _T_63200 = $signed(buffer_2_523) + $signed(buffer_2_524); // @[Modules.scala 166:64:@9319.4]
  assign _T_63201 = _T_63200[13:0]; // @[Modules.scala 166:64:@9320.4]
  assign buffer_2_571 = $signed(_T_63201); // @[Modules.scala 166:64:@9321.4]
  assign _T_63203 = $signed(buffer_2_525) + $signed(buffer_2_526); // @[Modules.scala 166:64:@9323.4]
  assign _T_63204 = _T_63203[13:0]; // @[Modules.scala 166:64:@9324.4]
  assign buffer_2_572 = $signed(_T_63204); // @[Modules.scala 166:64:@9325.4]
  assign _T_63206 = $signed(buffer_2_527) + $signed(buffer_2_528); // @[Modules.scala 166:64:@9327.4]
  assign _T_63207 = _T_63206[13:0]; // @[Modules.scala 166:64:@9328.4]
  assign buffer_2_573 = $signed(_T_63207); // @[Modules.scala 166:64:@9329.4]
  assign _T_63209 = $signed(buffer_2_529) + $signed(buffer_2_530); // @[Modules.scala 166:64:@9331.4]
  assign _T_63210 = _T_63209[13:0]; // @[Modules.scala 166:64:@9332.4]
  assign buffer_2_574 = $signed(_T_63210); // @[Modules.scala 166:64:@9333.4]
  assign _T_63212 = $signed(buffer_2_531) + $signed(buffer_2_532); // @[Modules.scala 166:64:@9335.4]
  assign _T_63213 = _T_63212[13:0]; // @[Modules.scala 166:64:@9336.4]
  assign buffer_2_575 = $signed(_T_63213); // @[Modules.scala 166:64:@9337.4]
  assign _T_63215 = $signed(buffer_2_533) + $signed(buffer_2_534); // @[Modules.scala 166:64:@9339.4]
  assign _T_63216 = _T_63215[13:0]; // @[Modules.scala 166:64:@9340.4]
  assign buffer_2_576 = $signed(_T_63216); // @[Modules.scala 166:64:@9341.4]
  assign _T_63218 = $signed(buffer_2_535) + $signed(buffer_2_536); // @[Modules.scala 166:64:@9343.4]
  assign _T_63219 = _T_63218[13:0]; // @[Modules.scala 166:64:@9344.4]
  assign buffer_2_577 = $signed(_T_63219); // @[Modules.scala 166:64:@9345.4]
  assign _T_63221 = $signed(buffer_2_537) + $signed(buffer_2_538); // @[Modules.scala 166:64:@9347.4]
  assign _T_63222 = _T_63221[13:0]; // @[Modules.scala 166:64:@9348.4]
  assign buffer_2_578 = $signed(_T_63222); // @[Modules.scala 166:64:@9349.4]
  assign _T_63224 = $signed(buffer_2_539) + $signed(buffer_2_540); // @[Modules.scala 166:64:@9351.4]
  assign _T_63225 = _T_63224[13:0]; // @[Modules.scala 166:64:@9352.4]
  assign buffer_2_579 = $signed(_T_63225); // @[Modules.scala 166:64:@9353.4]
  assign _T_63227 = $signed(buffer_2_541) + $signed(buffer_2_464); // @[Modules.scala 172:66:@9355.4]
  assign _T_63228 = _T_63227[13:0]; // @[Modules.scala 172:66:@9356.4]
  assign buffer_2_580 = $signed(_T_63228); // @[Modules.scala 172:66:@9357.4]
  assign _T_63230 = $signed(buffer_2_542) + $signed(buffer_2_543); // @[Modules.scala 166:64:@9359.4]
  assign _T_63231 = _T_63230[13:0]; // @[Modules.scala 166:64:@9360.4]
  assign buffer_2_581 = $signed(_T_63231); // @[Modules.scala 166:64:@9361.4]
  assign _T_63233 = $signed(buffer_2_544) + $signed(buffer_2_545); // @[Modules.scala 166:64:@9363.4]
  assign _T_63234 = _T_63233[13:0]; // @[Modules.scala 166:64:@9364.4]
  assign buffer_2_582 = $signed(_T_63234); // @[Modules.scala 166:64:@9365.4]
  assign _T_63236 = $signed(buffer_2_546) + $signed(buffer_2_547); // @[Modules.scala 166:64:@9367.4]
  assign _T_63237 = _T_63236[13:0]; // @[Modules.scala 166:64:@9368.4]
  assign buffer_2_583 = $signed(_T_63237); // @[Modules.scala 166:64:@9369.4]
  assign _T_63239 = $signed(buffer_2_548) + $signed(buffer_2_549); // @[Modules.scala 166:64:@9371.4]
  assign _T_63240 = _T_63239[13:0]; // @[Modules.scala 166:64:@9372.4]
  assign buffer_2_584 = $signed(_T_63240); // @[Modules.scala 166:64:@9373.4]
  assign _T_63242 = $signed(buffer_2_550) + $signed(buffer_2_551); // @[Modules.scala 166:64:@9375.4]
  assign _T_63243 = _T_63242[13:0]; // @[Modules.scala 166:64:@9376.4]
  assign buffer_2_585 = $signed(_T_63243); // @[Modules.scala 166:64:@9377.4]
  assign _T_63245 = $signed(buffer_2_552) + $signed(buffer_2_553); // @[Modules.scala 166:64:@9379.4]
  assign _T_63246 = _T_63245[13:0]; // @[Modules.scala 166:64:@9380.4]
  assign buffer_2_586 = $signed(_T_63246); // @[Modules.scala 166:64:@9381.4]
  assign _T_63248 = $signed(buffer_2_554) + $signed(buffer_2_555); // @[Modules.scala 166:64:@9383.4]
  assign _T_63249 = _T_63248[13:0]; // @[Modules.scala 166:64:@9384.4]
  assign buffer_2_587 = $signed(_T_63249); // @[Modules.scala 166:64:@9385.4]
  assign _T_63251 = $signed(buffer_2_556) + $signed(buffer_2_557); // @[Modules.scala 166:64:@9387.4]
  assign _T_63252 = _T_63251[13:0]; // @[Modules.scala 166:64:@9388.4]
  assign buffer_2_588 = $signed(_T_63252); // @[Modules.scala 166:64:@9389.4]
  assign _T_63254 = $signed(buffer_2_558) + $signed(buffer_2_559); // @[Modules.scala 166:64:@9391.4]
  assign _T_63255 = _T_63254[13:0]; // @[Modules.scala 166:64:@9392.4]
  assign buffer_2_589 = $signed(_T_63255); // @[Modules.scala 166:64:@9393.4]
  assign _T_63257 = $signed(buffer_2_560) + $signed(buffer_2_561); // @[Modules.scala 166:64:@9395.4]
  assign _T_63258 = _T_63257[13:0]; // @[Modules.scala 166:64:@9396.4]
  assign buffer_2_590 = $signed(_T_63258); // @[Modules.scala 166:64:@9397.4]
  assign _T_63260 = $signed(buffer_2_562) + $signed(buffer_2_563); // @[Modules.scala 166:64:@9399.4]
  assign _T_63261 = _T_63260[13:0]; // @[Modules.scala 166:64:@9400.4]
  assign buffer_2_591 = $signed(_T_63261); // @[Modules.scala 166:64:@9401.4]
  assign _T_63263 = $signed(buffer_2_564) + $signed(buffer_2_565); // @[Modules.scala 166:64:@9403.4]
  assign _T_63264 = _T_63263[13:0]; // @[Modules.scala 166:64:@9404.4]
  assign buffer_2_592 = $signed(_T_63264); // @[Modules.scala 166:64:@9405.4]
  assign _T_63266 = $signed(buffer_2_566) + $signed(buffer_2_567); // @[Modules.scala 166:64:@9407.4]
  assign _T_63267 = _T_63266[13:0]; // @[Modules.scala 166:64:@9408.4]
  assign buffer_2_593 = $signed(_T_63267); // @[Modules.scala 166:64:@9409.4]
  assign _T_63269 = $signed(buffer_2_568) + $signed(buffer_2_569); // @[Modules.scala 166:64:@9411.4]
  assign _T_63270 = _T_63269[13:0]; // @[Modules.scala 166:64:@9412.4]
  assign buffer_2_594 = $signed(_T_63270); // @[Modules.scala 166:64:@9413.4]
  assign _T_63272 = $signed(buffer_2_570) + $signed(buffer_2_571); // @[Modules.scala 166:64:@9415.4]
  assign _T_63273 = _T_63272[13:0]; // @[Modules.scala 166:64:@9416.4]
  assign buffer_2_595 = $signed(_T_63273); // @[Modules.scala 166:64:@9417.4]
  assign _T_63275 = $signed(buffer_2_572) + $signed(buffer_2_573); // @[Modules.scala 166:64:@9419.4]
  assign _T_63276 = _T_63275[13:0]; // @[Modules.scala 166:64:@9420.4]
  assign buffer_2_596 = $signed(_T_63276); // @[Modules.scala 166:64:@9421.4]
  assign _T_63278 = $signed(buffer_2_574) + $signed(buffer_2_575); // @[Modules.scala 166:64:@9423.4]
  assign _T_63279 = _T_63278[13:0]; // @[Modules.scala 166:64:@9424.4]
  assign buffer_2_597 = $signed(_T_63279); // @[Modules.scala 166:64:@9425.4]
  assign _T_63281 = $signed(buffer_2_576) + $signed(buffer_2_577); // @[Modules.scala 166:64:@9427.4]
  assign _T_63282 = _T_63281[13:0]; // @[Modules.scala 166:64:@9428.4]
  assign buffer_2_598 = $signed(_T_63282); // @[Modules.scala 166:64:@9429.4]
  assign _T_63284 = $signed(buffer_2_578) + $signed(buffer_2_579); // @[Modules.scala 166:64:@9431.4]
  assign _T_63285 = _T_63284[13:0]; // @[Modules.scala 166:64:@9432.4]
  assign buffer_2_599 = $signed(_T_63285); // @[Modules.scala 166:64:@9433.4]
  assign _T_63287 = $signed(buffer_2_581) + $signed(buffer_2_582); // @[Modules.scala 166:64:@9435.4]
  assign _T_63288 = _T_63287[13:0]; // @[Modules.scala 166:64:@9436.4]
  assign buffer_2_600 = $signed(_T_63288); // @[Modules.scala 166:64:@9437.4]
  assign _T_63290 = $signed(buffer_2_583) + $signed(buffer_2_584); // @[Modules.scala 166:64:@9439.4]
  assign _T_63291 = _T_63290[13:0]; // @[Modules.scala 166:64:@9440.4]
  assign buffer_2_601 = $signed(_T_63291); // @[Modules.scala 166:64:@9441.4]
  assign _T_63293 = $signed(buffer_2_585) + $signed(buffer_2_586); // @[Modules.scala 166:64:@9443.4]
  assign _T_63294 = _T_63293[13:0]; // @[Modules.scala 166:64:@9444.4]
  assign buffer_2_602 = $signed(_T_63294); // @[Modules.scala 166:64:@9445.4]
  assign _T_63296 = $signed(buffer_2_587) + $signed(buffer_2_588); // @[Modules.scala 166:64:@9447.4]
  assign _T_63297 = _T_63296[13:0]; // @[Modules.scala 166:64:@9448.4]
  assign buffer_2_603 = $signed(_T_63297); // @[Modules.scala 166:64:@9449.4]
  assign _T_63299 = $signed(buffer_2_589) + $signed(buffer_2_590); // @[Modules.scala 166:64:@9451.4]
  assign _T_63300 = _T_63299[13:0]; // @[Modules.scala 166:64:@9452.4]
  assign buffer_2_604 = $signed(_T_63300); // @[Modules.scala 166:64:@9453.4]
  assign _T_63302 = $signed(buffer_2_591) + $signed(buffer_2_592); // @[Modules.scala 166:64:@9455.4]
  assign _T_63303 = _T_63302[13:0]; // @[Modules.scala 166:64:@9456.4]
  assign buffer_2_605 = $signed(_T_63303); // @[Modules.scala 166:64:@9457.4]
  assign _T_63305 = $signed(buffer_2_593) + $signed(buffer_2_594); // @[Modules.scala 166:64:@9459.4]
  assign _T_63306 = _T_63305[13:0]; // @[Modules.scala 166:64:@9460.4]
  assign buffer_2_606 = $signed(_T_63306); // @[Modules.scala 166:64:@9461.4]
  assign _T_63308 = $signed(buffer_2_595) + $signed(buffer_2_596); // @[Modules.scala 166:64:@9463.4]
  assign _T_63309 = _T_63308[13:0]; // @[Modules.scala 166:64:@9464.4]
  assign buffer_2_607 = $signed(_T_63309); // @[Modules.scala 166:64:@9465.4]
  assign _T_63311 = $signed(buffer_2_597) + $signed(buffer_2_598); // @[Modules.scala 166:64:@9467.4]
  assign _T_63312 = _T_63311[13:0]; // @[Modules.scala 166:64:@9468.4]
  assign buffer_2_608 = $signed(_T_63312); // @[Modules.scala 166:64:@9469.4]
  assign _T_63314 = $signed(buffer_2_599) + $signed(buffer_2_580); // @[Modules.scala 172:66:@9471.4]
  assign _T_63315 = _T_63314[13:0]; // @[Modules.scala 172:66:@9472.4]
  assign buffer_2_609 = $signed(_T_63315); // @[Modules.scala 172:66:@9473.4]
  assign _T_63317 = $signed(buffer_2_600) + $signed(buffer_2_601); // @[Modules.scala 160:64:@9475.4]
  assign _T_63318 = _T_63317[13:0]; // @[Modules.scala 160:64:@9476.4]
  assign buffer_2_610 = $signed(_T_63318); // @[Modules.scala 160:64:@9477.4]
  assign _T_63320 = $signed(buffer_2_602) + $signed(buffer_2_603); // @[Modules.scala 160:64:@9479.4]
  assign _T_63321 = _T_63320[13:0]; // @[Modules.scala 160:64:@9480.4]
  assign buffer_2_611 = $signed(_T_63321); // @[Modules.scala 160:64:@9481.4]
  assign _T_63323 = $signed(buffer_2_604) + $signed(buffer_2_605); // @[Modules.scala 160:64:@9483.4]
  assign _T_63324 = _T_63323[13:0]; // @[Modules.scala 160:64:@9484.4]
  assign buffer_2_612 = $signed(_T_63324); // @[Modules.scala 160:64:@9485.4]
  assign _T_63326 = $signed(buffer_2_606) + $signed(buffer_2_607); // @[Modules.scala 160:64:@9487.4]
  assign _T_63327 = _T_63326[13:0]; // @[Modules.scala 160:64:@9488.4]
  assign buffer_2_613 = $signed(_T_63327); // @[Modules.scala 160:64:@9489.4]
  assign _T_63329 = $signed(buffer_2_608) + $signed(buffer_2_609); // @[Modules.scala 160:64:@9491.4]
  assign _T_63330 = _T_63329[13:0]; // @[Modules.scala 160:64:@9492.4]
  assign buffer_2_614 = $signed(_T_63330); // @[Modules.scala 160:64:@9493.4]
  assign _T_63332 = $signed(buffer_2_610) + $signed(buffer_2_611); // @[Modules.scala 166:64:@9495.4]
  assign _T_63333 = _T_63332[13:0]; // @[Modules.scala 166:64:@9496.4]
  assign buffer_2_615 = $signed(_T_63333); // @[Modules.scala 166:64:@9497.4]
  assign _T_63335 = $signed(buffer_2_612) + $signed(buffer_2_613); // @[Modules.scala 166:64:@9499.4]
  assign _T_63336 = _T_63335[13:0]; // @[Modules.scala 166:64:@9500.4]
  assign buffer_2_616 = $signed(_T_63336); // @[Modules.scala 166:64:@9501.4]
  assign _T_63338 = $signed(buffer_2_615) + $signed(buffer_2_616); // @[Modules.scala 160:64:@9503.4]
  assign _T_63339 = _T_63338[13:0]; // @[Modules.scala 160:64:@9504.4]
  assign buffer_2_617 = $signed(_T_63339); // @[Modules.scala 160:64:@9505.4]
  assign _T_63341 = $signed(buffer_2_617) + $signed(buffer_2_614); // @[Modules.scala 172:66:@9507.4]
  assign _T_63342 = _T_63341[13:0]; // @[Modules.scala 172:66:@9508.4]
  assign buffer_2_618 = $signed(_T_63342); // @[Modules.scala 172:66:@9509.4]
  assign _T_63362 = $signed(_T_54215) + $signed(_T_54220); // @[Modules.scala 150:103:@9690.4]
  assign _T_63363 = _T_63362[5:0]; // @[Modules.scala 150:103:@9691.4]
  assign _T_63364 = $signed(_T_63363); // @[Modules.scala 150:103:@9692.4]
  assign _T_63375 = $signed(-4'sh1) * $signed(io_in_39); // @[Modules.scala 151:80:@9701.4]
  assign _T_63376 = $signed(_T_57241) + $signed(_T_63375); // @[Modules.scala 150:103:@9702.4]
  assign _T_63377 = _T_63376[4:0]; // @[Modules.scala 150:103:@9703.4]
  assign _T_63378 = $signed(_T_63377); // @[Modules.scala 150:103:@9704.4]
  assign _GEN_218 = {{1{_T_57260[4]}},_T_57260}; // @[Modules.scala 150:103:@9714.4]
  assign _T_63390 = $signed(_T_54243) + $signed(_GEN_218); // @[Modules.scala 150:103:@9714.4]
  assign _T_63391 = _T_63390[5:0]; // @[Modules.scala 150:103:@9715.4]
  assign _T_63392 = $signed(_T_63391); // @[Modules.scala 150:103:@9716.4]
  assign _T_63397 = $signed(_T_60299) + $signed(_T_57262); // @[Modules.scala 150:103:@9720.4]
  assign _T_63398 = _T_63397[4:0]; // @[Modules.scala 150:103:@9721.4]
  assign _T_63399 = $signed(_T_63398); // @[Modules.scala 150:103:@9722.4]
  assign _T_63403 = $signed(-4'sh1) * $signed(io_in_47); // @[Modules.scala 151:80:@9725.4]
  assign _T_63404 = $signed(_T_57267) + $signed(_T_63403); // @[Modules.scala 150:103:@9726.4]
  assign _T_63405 = _T_63404[4:0]; // @[Modules.scala 150:103:@9727.4]
  assign _T_63406 = $signed(_T_63405); // @[Modules.scala 150:103:@9728.4]
  assign _T_63408 = $signed(-4'sh1) * $signed(io_in_48); // @[Modules.scala 150:74:@9730.4]
  assign _T_63411 = $signed(_T_63408) + $signed(_T_57274); // @[Modules.scala 150:103:@9732.4]
  assign _T_63412 = _T_63411[4:0]; // @[Modules.scala 150:103:@9733.4]
  assign _T_63413 = $signed(_T_63412); // @[Modules.scala 150:103:@9734.4]
  assign _T_63418 = $signed(_T_54271) + $signed(_GEN_79); // @[Modules.scala 150:103:@9738.4]
  assign _T_63419 = _T_63418[5:0]; // @[Modules.scala 150:103:@9739.4]
  assign _T_63420 = $signed(_T_63419); // @[Modules.scala 150:103:@9740.4]
  assign _T_63422 = $signed(-4'sh1) * $signed(io_in_54); // @[Modules.scala 150:74:@9742.4]
  assign _T_63425 = $signed(_T_63422) + $signed(_T_60327); // @[Modules.scala 150:103:@9744.4]
  assign _T_63426 = _T_63425[4:0]; // @[Modules.scala 150:103:@9745.4]
  assign _T_63427 = $signed(_T_63426); // @[Modules.scala 150:103:@9746.4]
  assign _T_63429 = $signed(4'sh1) * $signed(io_in_60); // @[Modules.scala 150:74:@9748.4]
  assign _T_63432 = $signed(_T_63429) + $signed(_T_54283); // @[Modules.scala 150:103:@9750.4]
  assign _T_63433 = _T_63432[5:0]; // @[Modules.scala 150:103:@9751.4]
  assign _T_63434 = $signed(_T_63433); // @[Modules.scala 150:103:@9752.4]
  assign _GEN_220 = {{1{_T_57309[4]}},_T_57309}; // @[Modules.scala 150:103:@9756.4]
  assign _T_63439 = $signed(_T_54292) + $signed(_GEN_220); // @[Modules.scala 150:103:@9756.4]
  assign _T_63440 = _T_63439[5:0]; // @[Modules.scala 150:103:@9757.4]
  assign _T_63441 = $signed(_T_63440); // @[Modules.scala 150:103:@9758.4]
  assign _T_63467 = $signed(_T_57332) + $signed(_T_57337); // @[Modules.scala 150:103:@9780.4]
  assign _T_63468 = _T_63467[4:0]; // @[Modules.scala 150:103:@9781.4]
  assign _T_63469 = $signed(_T_63468); // @[Modules.scala 150:103:@9782.4]
  assign _GEN_221 = {{1{_T_57339[4]}},_T_57339}; // @[Modules.scala 150:103:@9786.4]
  assign _T_63474 = $signed(_GEN_221) + $signed(_T_54334); // @[Modules.scala 150:103:@9786.4]
  assign _T_63475 = _T_63474[5:0]; // @[Modules.scala 150:103:@9787.4]
  assign _T_63476 = $signed(_T_63475); // @[Modules.scala 150:103:@9788.4]
  assign _T_63485 = $signed(-4'sh1) * $signed(io_in_79); // @[Modules.scala 150:74:@9796.4]
  assign _T_63487 = $signed(-4'sh1) * $signed(io_in_80); // @[Modules.scala 151:80:@9797.4]
  assign _T_63488 = $signed(_T_63485) + $signed(_T_63487); // @[Modules.scala 150:103:@9798.4]
  assign _T_63489 = _T_63488[4:0]; // @[Modules.scala 150:103:@9799.4]
  assign _T_63490 = $signed(_T_63489); // @[Modules.scala 150:103:@9800.4]
  assign _T_63492 = $signed(-4'sh1) * $signed(io_in_81); // @[Modules.scala 150:74:@9802.4]
  assign _T_63495 = $signed(_T_63492) + $signed(_T_54355); // @[Modules.scala 150:103:@9804.4]
  assign _T_63496 = _T_63495[4:0]; // @[Modules.scala 150:103:@9805.4]
  assign _T_63497 = $signed(_T_63496); // @[Modules.scala 150:103:@9806.4]
  assign _T_63499 = $signed(-4'sh1) * $signed(io_in_87); // @[Modules.scala 150:74:@9808.4]
  assign _T_63502 = $signed(_T_63499) + $signed(_T_60402); // @[Modules.scala 150:103:@9810.4]
  assign _T_63503 = _T_63502[4:0]; // @[Modules.scala 150:103:@9811.4]
  assign _T_63504 = $signed(_T_63503); // @[Modules.scala 150:103:@9812.4]
  assign _T_63509 = $signed(_T_60404) + $signed(_T_57379); // @[Modules.scala 150:103:@9816.4]
  assign _T_63510 = _T_63509[4:0]; // @[Modules.scala 150:103:@9817.4]
  assign _T_63511 = $signed(_T_63510); // @[Modules.scala 150:103:@9818.4]
  assign _T_63516 = $signed(_T_57381) + $signed(_T_57386); // @[Modules.scala 150:103:@9822.4]
  assign _T_63517 = _T_63516[4:0]; // @[Modules.scala 150:103:@9823.4]
  assign _T_63518 = $signed(_T_63517); // @[Modules.scala 150:103:@9824.4]
  assign _T_63523 = $signed(_T_57388) + $signed(_T_57393); // @[Modules.scala 150:103:@9828.4]
  assign _T_63524 = _T_63523[4:0]; // @[Modules.scala 150:103:@9829.4]
  assign _T_63525 = $signed(_T_63524); // @[Modules.scala 150:103:@9830.4]
  assign _T_63530 = $signed(_T_57395) + $signed(_T_57400); // @[Modules.scala 150:103:@9834.4]
  assign _T_63531 = _T_63530[4:0]; // @[Modules.scala 150:103:@9835.4]
  assign _T_63532 = $signed(_T_63531); // @[Modules.scala 150:103:@9836.4]
  assign _T_63537 = $signed(_T_57402) + $signed(_T_60430); // @[Modules.scala 150:103:@9840.4]
  assign _T_63538 = _T_63537[4:0]; // @[Modules.scala 150:103:@9841.4]
  assign _T_63539 = $signed(_T_63538); // @[Modules.scala 150:103:@9842.4]
  assign _T_63541 = $signed(-4'sh1) * $signed(io_in_99); // @[Modules.scala 150:74:@9844.4]
  assign _T_63543 = $signed(-4'sh1) * $signed(io_in_100); // @[Modules.scala 151:80:@9845.4]
  assign _T_63544 = $signed(_T_63541) + $signed(_T_63543); // @[Modules.scala 150:103:@9846.4]
  assign _T_63545 = _T_63544[4:0]; // @[Modules.scala 150:103:@9847.4]
  assign _T_63546 = $signed(_T_63545); // @[Modules.scala 150:103:@9848.4]
  assign _T_63551 = $signed(_T_57409) + $signed(_T_57414); // @[Modules.scala 150:103:@9852.4]
  assign _T_63552 = _T_63551[4:0]; // @[Modules.scala 150:103:@9853.4]
  assign _T_63553 = $signed(_T_63552); // @[Modules.scala 150:103:@9854.4]
  assign _T_63558 = $signed(_T_57416) + $signed(_T_57421); // @[Modules.scala 150:103:@9858.4]
  assign _T_63559 = _T_63558[4:0]; // @[Modules.scala 150:103:@9859.4]
  assign _T_63560 = $signed(_T_63559); // @[Modules.scala 150:103:@9860.4]
  assign _GEN_222 = {{1{_T_57430[4]}},_T_57430}; // @[Modules.scala 150:103:@9864.4]
  assign _T_63565 = $signed(_T_54425) + $signed(_GEN_222); // @[Modules.scala 150:103:@9864.4]
  assign _T_63566 = _T_63565[5:0]; // @[Modules.scala 150:103:@9865.4]
  assign _T_63567 = $signed(_T_63566); // @[Modules.scala 150:103:@9866.4]
  assign _T_63571 = $signed(-4'sh1) * $signed(io_in_109); // @[Modules.scala 151:80:@9869.4]
  assign _T_63572 = $signed(_T_57435) + $signed(_T_63571); // @[Modules.scala 150:103:@9870.4]
  assign _T_63573 = _T_63572[4:0]; // @[Modules.scala 150:103:@9871.4]
  assign _T_63574 = $signed(_T_63573); // @[Modules.scala 150:103:@9872.4]
  assign _T_63585 = $signed(-4'sh1) * $signed(io_in_115); // @[Modules.scala 151:80:@9881.4]
  assign _T_63586 = $signed(_T_54446) + $signed(_T_63585); // @[Modules.scala 150:103:@9882.4]
  assign _T_63587 = _T_63586[4:0]; // @[Modules.scala 150:103:@9883.4]
  assign _T_63588 = $signed(_T_63587); // @[Modules.scala 150:103:@9884.4]
  assign _T_63590 = $signed(-4'sh1) * $signed(io_in_116); // @[Modules.scala 150:74:@9886.4]
  assign _T_63593 = $signed(_T_63590) + $signed(_T_54453); // @[Modules.scala 150:103:@9888.4]
  assign _T_63594 = _T_63593[4:0]; // @[Modules.scala 150:103:@9889.4]
  assign _T_63595 = $signed(_T_63594); // @[Modules.scala 150:103:@9890.4]
  assign _T_63599 = $signed(-4'sh1) * $signed(io_in_119); // @[Modules.scala 151:80:@9893.4]
  assign _T_63600 = $signed(_T_54458) + $signed(_T_63599); // @[Modules.scala 150:103:@9894.4]
  assign _T_63601 = _T_63600[4:0]; // @[Modules.scala 150:103:@9895.4]
  assign _T_63602 = $signed(_T_63601); // @[Modules.scala 150:103:@9896.4]
  assign _T_63604 = $signed(-4'sh1) * $signed(io_in_120); // @[Modules.scala 150:74:@9898.4]
  assign _T_63606 = $signed(-4'sh1) * $signed(io_in_121); // @[Modules.scala 151:80:@9899.4]
  assign _T_63607 = $signed(_T_63604) + $signed(_T_63606); // @[Modules.scala 150:103:@9900.4]
  assign _T_63608 = _T_63607[4:0]; // @[Modules.scala 150:103:@9901.4]
  assign _T_63609 = $signed(_T_63608); // @[Modules.scala 150:103:@9902.4]
  assign _T_63614 = $signed(_T_60495) + $signed(_T_60500); // @[Modules.scala 150:103:@9906.4]
  assign _T_63615 = _T_63614[4:0]; // @[Modules.scala 150:103:@9907.4]
  assign _T_63616 = $signed(_T_63615); // @[Modules.scala 150:103:@9908.4]
  assign _T_63621 = $signed(_T_60502) + $signed(_T_60507); // @[Modules.scala 150:103:@9912.4]
  assign _T_63622 = _T_63621[4:0]; // @[Modules.scala 150:103:@9913.4]
  assign _T_63623 = $signed(_T_63622); // @[Modules.scala 150:103:@9914.4]
  assign _GEN_223 = {{1{_T_60509[4]}},_T_60509}; // @[Modules.scala 150:103:@9918.4]
  assign _T_63628 = $signed(_GEN_223) + $signed(_T_54488); // @[Modules.scala 150:103:@9918.4]
  assign _T_63629 = _T_63628[5:0]; // @[Modules.scala 150:103:@9919.4]
  assign _T_63630 = $signed(_T_63629); // @[Modules.scala 150:103:@9920.4]
  assign _T_63635 = $signed(_T_54495) + $signed(_T_57498); // @[Modules.scala 150:103:@9924.4]
  assign _T_63636 = _T_63635[5:0]; // @[Modules.scala 150:103:@9925.4]
  assign _T_63637 = $signed(_T_63636); // @[Modules.scala 150:103:@9926.4]
  assign _T_63649 = $signed(_T_57507) + $signed(_T_57512); // @[Modules.scala 150:103:@9936.4]
  assign _T_63650 = _T_63649[5:0]; // @[Modules.scala 150:103:@9937.4]
  assign _T_63651 = $signed(_T_63650); // @[Modules.scala 150:103:@9938.4]
  assign _T_63656 = $signed(_T_57514) + $signed(_T_54516); // @[Modules.scala 150:103:@9942.4]
  assign _T_63657 = _T_63656[5:0]; // @[Modules.scala 150:103:@9943.4]
  assign _T_63658 = $signed(_T_63657); // @[Modules.scala 150:103:@9944.4]
  assign _T_63663 = $signed(_T_60549) + $signed(_T_57526); // @[Modules.scala 150:103:@9948.4]
  assign _T_63664 = _T_63663[5:0]; // @[Modules.scala 150:103:@9949.4]
  assign _T_63665 = $signed(_T_63664); // @[Modules.scala 150:103:@9950.4]
  assign _T_63669 = $signed(-4'sh1) * $signed(io_in_144); // @[Modules.scala 151:80:@9953.4]
  assign _T_63670 = $signed(_T_60556) + $signed(_T_63669); // @[Modules.scala 150:103:@9954.4]
  assign _T_63671 = _T_63670[4:0]; // @[Modules.scala 150:103:@9955.4]
  assign _T_63672 = $signed(_T_63671); // @[Modules.scala 150:103:@9956.4]
  assign _T_63683 = $signed(-4'sh1) * $signed(io_in_148); // @[Modules.scala 151:80:@9965.4]
  assign _T_63684 = $signed(_T_54528) + $signed(_T_63683); // @[Modules.scala 150:103:@9966.4]
  assign _T_63685 = _T_63684[4:0]; // @[Modules.scala 150:103:@9967.4]
  assign _T_63686 = $signed(_T_63685); // @[Modules.scala 150:103:@9968.4]
  assign _T_63688 = $signed(-4'sh1) * $signed(io_in_149); // @[Modules.scala 150:74:@9970.4]
  assign _T_63691 = $signed(_T_63688) + $signed(_T_60577); // @[Modules.scala 150:103:@9972.4]
  assign _T_63692 = _T_63691[4:0]; // @[Modules.scala 150:103:@9973.4]
  assign _T_63693 = $signed(_T_63692); // @[Modules.scala 150:103:@9974.4]
  assign _T_63698 = $signed(_T_60579) + $signed(_T_60584); // @[Modules.scala 150:103:@9978.4]
  assign _T_63699 = _T_63698[4:0]; // @[Modules.scala 150:103:@9979.4]
  assign _T_63700 = $signed(_T_63699); // @[Modules.scala 150:103:@9980.4]
  assign _T_63704 = $signed(4'sh1) * $signed(io_in_154); // @[Modules.scala 151:80:@9983.4]
  assign _GEN_224 = {{1{_T_60586[4]}},_T_60586}; // @[Modules.scala 150:103:@9984.4]
  assign _T_63705 = $signed(_GEN_224) + $signed(_T_63704); // @[Modules.scala 150:103:@9984.4]
  assign _T_63706 = _T_63705[5:0]; // @[Modules.scala 150:103:@9985.4]
  assign _T_63707 = $signed(_T_63706); // @[Modules.scala 150:103:@9986.4]
  assign _T_63712 = $signed(_T_57563) + $signed(_T_54544); // @[Modules.scala 150:103:@9990.4]
  assign _T_63713 = _T_63712[4:0]; // @[Modules.scala 150:103:@9991.4]
  assign _T_63714 = $signed(_T_63713); // @[Modules.scala 150:103:@9992.4]
  assign _T_63719 = $signed(_T_54549) + $signed(_T_57575); // @[Modules.scala 150:103:@9996.4]
  assign _T_63720 = _T_63719[4:0]; // @[Modules.scala 150:103:@9997.4]
  assign _T_63721 = $signed(_T_63720); // @[Modules.scala 150:103:@9998.4]
  assign _T_63723 = $signed(4'sh1) * $signed(io_in_160); // @[Modules.scala 150:74:@10000.4]
  assign _T_63726 = $signed(_T_63723) + $signed(_T_54556); // @[Modules.scala 150:103:@10002.4]
  assign _T_63727 = _T_63726[5:0]; // @[Modules.scala 150:103:@10003.4]
  assign _T_63728 = $signed(_T_63727); // @[Modules.scala 150:103:@10004.4]
  assign _T_63730 = $signed(4'sh1) * $signed(io_in_162); // @[Modules.scala 150:74:@10006.4]
  assign _T_63733 = $signed(_T_63730) + $signed(_T_60614); // @[Modules.scala 150:103:@10008.4]
  assign _T_63734 = _T_63733[5:0]; // @[Modules.scala 150:103:@10009.4]
  assign _T_63735 = $signed(_T_63734); // @[Modules.scala 150:103:@10010.4]
  assign _T_63739 = $signed(4'sh1) * $signed(io_in_165); // @[Modules.scala 151:80:@10013.4]
  assign _T_63740 = $signed(_T_60619) + $signed(_T_63739); // @[Modules.scala 150:103:@10014.4]
  assign _T_63741 = _T_63740[5:0]; // @[Modules.scala 150:103:@10015.4]
  assign _T_63742 = $signed(_T_63741); // @[Modules.scala 150:103:@10016.4]
  assign _T_63746 = $signed(-4'sh1) * $signed(io_in_167); // @[Modules.scala 151:80:@10019.4]
  assign _GEN_225 = {{1{_T_63746[4]}},_T_63746}; // @[Modules.scala 150:103:@10020.4]
  assign _T_63747 = $signed(_T_54572) + $signed(_GEN_225); // @[Modules.scala 150:103:@10020.4]
  assign _T_63748 = _T_63747[5:0]; // @[Modules.scala 150:103:@10021.4]
  assign _T_63749 = $signed(_T_63748); // @[Modules.scala 150:103:@10022.4]
  assign _T_63754 = $signed(_T_60628) + $signed(_GEN_13); // @[Modules.scala 150:103:@10026.4]
  assign _T_63755 = _T_63754[5:0]; // @[Modules.scala 150:103:@10027.4]
  assign _T_63756 = $signed(_T_63755); // @[Modules.scala 150:103:@10028.4]
  assign _T_63760 = $signed(-4'sh1) * $signed(io_in_172); // @[Modules.scala 151:80:@10031.4]
  assign _T_63761 = $signed(_T_60635) + $signed(_T_63760); // @[Modules.scala 150:103:@10032.4]
  assign _T_63762 = _T_63761[4:0]; // @[Modules.scala 150:103:@10033.4]
  assign _T_63763 = $signed(_T_63762); // @[Modules.scala 150:103:@10034.4]
  assign _T_63768 = $signed(_T_60642) + $signed(_T_60647); // @[Modules.scala 150:103:@10038.4]
  assign _T_63769 = _T_63768[4:0]; // @[Modules.scala 150:103:@10039.4]
  assign _T_63770 = $signed(_T_63769); // @[Modules.scala 150:103:@10040.4]
  assign _T_63772 = $signed(-4'sh1) * $signed(io_in_175); // @[Modules.scala 150:74:@10042.4]
  assign _T_63774 = $signed(-4'sh1) * $signed(io_in_176); // @[Modules.scala 151:80:@10043.4]
  assign _T_63775 = $signed(_T_63772) + $signed(_T_63774); // @[Modules.scala 150:103:@10044.4]
  assign _T_63776 = _T_63775[4:0]; // @[Modules.scala 150:103:@10045.4]
  assign _T_63777 = $signed(_T_63776); // @[Modules.scala 150:103:@10046.4]
  assign _T_63782 = $signed(_T_57619) + $signed(_T_54607); // @[Modules.scala 150:103:@10050.4]
  assign _T_63783 = _T_63782[4:0]; // @[Modules.scala 150:103:@10051.4]
  assign _T_63784 = $signed(_T_63783); // @[Modules.scala 150:103:@10052.4]
  assign _GEN_227 = {{1{_T_60656[4]}},_T_60656}; // @[Modules.scala 150:103:@10056.4]
  assign _T_63789 = $signed(_GEN_227) + $signed(_T_57631); // @[Modules.scala 150:103:@10056.4]
  assign _T_63790 = _T_63789[5:0]; // @[Modules.scala 150:103:@10057.4]
  assign _T_63791 = $signed(_T_63790); // @[Modules.scala 150:103:@10058.4]
  assign _T_63796 = $signed(_T_54614) + $signed(_T_60668); // @[Modules.scala 150:103:@10062.4]
  assign _T_63797 = _T_63796[4:0]; // @[Modules.scala 150:103:@10063.4]
  assign _T_63798 = $signed(_T_63797); // @[Modules.scala 150:103:@10064.4]
  assign _T_63810 = $signed(_T_54628) + $signed(_T_60691); // @[Modules.scala 150:103:@10074.4]
  assign _T_63811 = _T_63810[4:0]; // @[Modules.scala 150:103:@10075.4]
  assign _T_63812 = $signed(_T_63811); // @[Modules.scala 150:103:@10076.4]
  assign _T_63814 = $signed(4'sh1) * $signed(io_in_190); // @[Modules.scala 150:74:@10078.4]
  assign _T_63817 = $signed(_T_63814) + $signed(_T_60698); // @[Modules.scala 150:103:@10080.4]
  assign _T_63818 = _T_63817[5:0]; // @[Modules.scala 150:103:@10081.4]
  assign _T_63819 = $signed(_T_63818); // @[Modules.scala 150:103:@10082.4]
  assign _T_63821 = $signed(4'sh1) * $signed(io_in_192); // @[Modules.scala 150:74:@10084.4]
  assign _T_63823 = $signed(4'sh1) * $signed(io_in_193); // @[Modules.scala 151:80:@10085.4]
  assign _T_63824 = $signed(_T_63821) + $signed(_T_63823); // @[Modules.scala 150:103:@10086.4]
  assign _T_63825 = _T_63824[5:0]; // @[Modules.scala 150:103:@10087.4]
  assign _T_63826 = $signed(_T_63825); // @[Modules.scala 150:103:@10088.4]
  assign _T_63828 = $signed(-4'sh1) * $signed(io_in_195); // @[Modules.scala 150:74:@10090.4]
  assign _GEN_228 = {{1{_T_63828[4]}},_T_63828}; // @[Modules.scala 150:103:@10092.4]
  assign _T_63831 = $signed(_GEN_228) + $signed(_T_57675); // @[Modules.scala 150:103:@10092.4]
  assign _T_63832 = _T_63831[5:0]; // @[Modules.scala 150:103:@10093.4]
  assign _T_63833 = $signed(_T_63832); // @[Modules.scala 150:103:@10094.4]
  assign _T_63835 = $signed(-4'sh1) * $signed(io_in_198); // @[Modules.scala 150:74:@10096.4]
  assign _T_63838 = $signed(_T_63835) + $signed(_T_60717); // @[Modules.scala 150:103:@10098.4]
  assign _T_63839 = _T_63838[4:0]; // @[Modules.scala 150:103:@10099.4]
  assign _T_63840 = $signed(_T_63839); // @[Modules.scala 150:103:@10100.4]
  assign _T_63845 = $signed(_T_60719) + $signed(_T_60724); // @[Modules.scala 150:103:@10104.4]
  assign _T_63846 = _T_63845[4:0]; // @[Modules.scala 150:103:@10105.4]
  assign _T_63847 = $signed(_T_63846); // @[Modules.scala 150:103:@10106.4]
  assign _T_63852 = $signed(_T_60726) + $signed(_T_57701); // @[Modules.scala 150:103:@10110.4]
  assign _T_63853 = _T_63852[4:0]; // @[Modules.scala 150:103:@10111.4]
  assign _T_63854 = $signed(_T_63853); // @[Modules.scala 150:103:@10112.4]
  assign _T_63859 = $signed(_T_60733) + $signed(_T_54684); // @[Modules.scala 150:103:@10116.4]
  assign _T_63860 = _T_63859[4:0]; // @[Modules.scala 150:103:@10117.4]
  assign _T_63861 = $signed(_T_63860); // @[Modules.scala 150:103:@10118.4]
  assign _T_63866 = $signed(_T_60740) + $signed(_T_60747); // @[Modules.scala 150:103:@10122.4]
  assign _T_63867 = _T_63866[4:0]; // @[Modules.scala 150:103:@10123.4]
  assign _T_63868 = $signed(_T_63867); // @[Modules.scala 150:103:@10124.4]
  assign _GEN_229 = {{1{_T_60752[4]}},_T_60752}; // @[Modules.scala 150:103:@10128.4]
  assign _T_63873 = $signed(_GEN_229) + $signed(_T_57722); // @[Modules.scala 150:103:@10128.4]
  assign _T_63874 = _T_63873[5:0]; // @[Modules.scala 150:103:@10129.4]
  assign _T_63875 = $signed(_T_63874); // @[Modules.scala 150:103:@10130.4]
  assign _T_63880 = $signed(_T_57724) + $signed(_T_57729); // @[Modules.scala 150:103:@10134.4]
  assign _T_63881 = _T_63880[5:0]; // @[Modules.scala 150:103:@10135.4]
  assign _T_63882 = $signed(_T_63881); // @[Modules.scala 150:103:@10136.4]
  assign _T_63884 = $signed(4'sh1) * $signed(io_in_214); // @[Modules.scala 150:74:@10138.4]
  assign _GEN_230 = {{1{_T_60773[4]}},_T_60773}; // @[Modules.scala 150:103:@10140.4]
  assign _T_63887 = $signed(_T_63884) + $signed(_GEN_230); // @[Modules.scala 150:103:@10140.4]
  assign _T_63888 = _T_63887[5:0]; // @[Modules.scala 150:103:@10141.4]
  assign _T_63889 = $signed(_T_63888); // @[Modules.scala 150:103:@10142.4]
  assign _T_63893 = $signed(4'sh1) * $signed(io_in_218); // @[Modules.scala 151:80:@10145.4]
  assign _GEN_231 = {{1{_T_54703[4]}},_T_54703}; // @[Modules.scala 150:103:@10146.4]
  assign _T_63894 = $signed(_GEN_231) + $signed(_T_63893); // @[Modules.scala 150:103:@10146.4]
  assign _T_63895 = _T_63894[5:0]; // @[Modules.scala 150:103:@10147.4]
  assign _T_63896 = $signed(_T_63895); // @[Modules.scala 150:103:@10148.4]
  assign _T_63898 = $signed(4'sh1) * $signed(io_in_219); // @[Modules.scala 150:74:@10150.4]
  assign _T_63900 = $signed(4'sh1) * $signed(io_in_220); // @[Modules.scala 151:80:@10151.4]
  assign _T_63901 = $signed(_T_63898) + $signed(_T_63900); // @[Modules.scala 150:103:@10152.4]
  assign _T_63902 = _T_63901[5:0]; // @[Modules.scala 150:103:@10153.4]
  assign _T_63903 = $signed(_T_63902); // @[Modules.scala 150:103:@10154.4]
  assign _T_63905 = $signed(4'sh1) * $signed(io_in_221); // @[Modules.scala 150:74:@10156.4]
  assign _T_63907 = $signed(4'sh1) * $signed(io_in_222); // @[Modules.scala 151:80:@10157.4]
  assign _T_63908 = $signed(_T_63905) + $signed(_T_63907); // @[Modules.scala 150:103:@10158.4]
  assign _T_63909 = _T_63908[5:0]; // @[Modules.scala 150:103:@10159.4]
  assign _T_63910 = $signed(_T_63909); // @[Modules.scala 150:103:@10160.4]
  assign _T_63915 = $signed(_T_57759) + $signed(_T_54726); // @[Modules.scala 150:103:@10164.4]
  assign _T_63916 = _T_63915[4:0]; // @[Modules.scala 150:103:@10165.4]
  assign _T_63917 = $signed(_T_63916); // @[Modules.scala 150:103:@10166.4]
  assign _T_63943 = $signed(_T_60831) + $signed(_T_57794); // @[Modules.scala 150:103:@10188.4]
  assign _T_63944 = _T_63943[4:0]; // @[Modules.scala 150:103:@10189.4]
  assign _T_63945 = $signed(_T_63944); // @[Modules.scala 150:103:@10190.4]
  assign _T_63950 = $signed(_T_60838) + $signed(_T_60845); // @[Modules.scala 150:103:@10194.4]
  assign _T_63951 = _T_63950[4:0]; // @[Modules.scala 150:103:@10195.4]
  assign _T_63952 = $signed(_T_63951); // @[Modules.scala 150:103:@10196.4]
  assign _T_63968 = $signed(4'sh1) * $signed(io_in_243); // @[Modules.scala 150:74:@10210.4]
  assign _T_63970 = $signed(4'sh1) * $signed(io_in_244); // @[Modules.scala 151:80:@10211.4]
  assign _T_63971 = $signed(_T_63968) + $signed(_T_63970); // @[Modules.scala 150:103:@10212.4]
  assign _T_63972 = _T_63971[5:0]; // @[Modules.scala 150:103:@10213.4]
  assign _T_63973 = $signed(_T_63972); // @[Modules.scala 150:103:@10214.4]
  assign _T_63975 = $signed(4'sh1) * $signed(io_in_246); // @[Modules.scala 150:74:@10216.4]
  assign _T_63977 = $signed(4'sh1) * $signed(io_in_247); // @[Modules.scala 151:80:@10217.4]
  assign _T_63978 = $signed(_T_63975) + $signed(_T_63977); // @[Modules.scala 150:103:@10218.4]
  assign _T_63979 = _T_63978[5:0]; // @[Modules.scala 150:103:@10219.4]
  assign _T_63980 = $signed(_T_63979); // @[Modules.scala 150:103:@10220.4]
  assign _T_63982 = $signed(4'sh1) * $signed(io_in_248); // @[Modules.scala 150:74:@10222.4]
  assign _T_63984 = $signed(4'sh1) * $signed(io_in_249); // @[Modules.scala 151:80:@10223.4]
  assign _T_63985 = $signed(_T_63982) + $signed(_T_63984); // @[Modules.scala 150:103:@10224.4]
  assign _T_63986 = _T_63985[5:0]; // @[Modules.scala 150:103:@10225.4]
  assign _T_63987 = $signed(_T_63986); // @[Modules.scala 150:103:@10226.4]
  assign _T_63989 = $signed(4'sh1) * $signed(io_in_250); // @[Modules.scala 150:74:@10228.4]
  assign _T_63992 = $signed(_T_63989) + $signed(_GEN_96); // @[Modules.scala 150:103:@10230.4]
  assign _T_63993 = _T_63992[5:0]; // @[Modules.scala 150:103:@10231.4]
  assign _T_63994 = $signed(_T_63993); // @[Modules.scala 150:103:@10232.4]
  assign _T_63996 = $signed(-4'sh1) * $signed(io_in_253); // @[Modules.scala 150:74:@10234.4]
  assign _T_63999 = $signed(_T_63996) + $signed(_T_60899); // @[Modules.scala 150:103:@10236.4]
  assign _T_64000 = _T_63999[4:0]; // @[Modules.scala 150:103:@10237.4]
  assign _T_64001 = $signed(_T_64000); // @[Modules.scala 150:103:@10238.4]
  assign _T_64006 = $signed(_T_60901) + $signed(_T_60906); // @[Modules.scala 150:103:@10242.4]
  assign _T_64007 = _T_64006[4:0]; // @[Modules.scala 150:103:@10243.4]
  assign _T_64008 = $signed(_T_64007); // @[Modules.scala 150:103:@10244.4]
  assign _T_64013 = $signed(_T_60908) + $signed(_T_60913); // @[Modules.scala 150:103:@10248.4]
  assign _T_64014 = _T_64013[4:0]; // @[Modules.scala 150:103:@10249.4]
  assign _T_64015 = $signed(_T_64014); // @[Modules.scala 150:103:@10250.4]
  assign _T_64019 = $signed(4'sh1) * $signed(io_in_261); // @[Modules.scala 151:80:@10253.4]
  assign _T_64020 = $signed(_T_54824) + $signed(_T_64019); // @[Modules.scala 150:103:@10254.4]
  assign _T_64021 = _T_64020[5:0]; // @[Modules.scala 150:103:@10255.4]
  assign _T_64022 = $signed(_T_64021); // @[Modules.scala 150:103:@10256.4]
  assign _T_64026 = $signed(4'sh1) * $signed(io_in_263); // @[Modules.scala 151:80:@10259.4]
  assign _T_64027 = $signed(_T_60922) + $signed(_T_64026); // @[Modules.scala 150:103:@10260.4]
  assign _T_64028 = _T_64027[5:0]; // @[Modules.scala 150:103:@10261.4]
  assign _T_64029 = $signed(_T_64028); // @[Modules.scala 150:103:@10262.4]
  assign _T_64034 = $signed(_T_54843) + $signed(_T_60934); // @[Modules.scala 150:103:@10266.4]
  assign _T_64035 = _T_64034[4:0]; // @[Modules.scala 150:103:@10267.4]
  assign _T_64036 = $signed(_T_64035); // @[Modules.scala 150:103:@10268.4]
  assign _T_64041 = $signed(_T_60936) + $signed(_T_54852); // @[Modules.scala 150:103:@10272.4]
  assign _T_64042 = _T_64041[4:0]; // @[Modules.scala 150:103:@10273.4]
  assign _T_64043 = $signed(_T_64042); // @[Modules.scala 150:103:@10274.4]
  assign _T_64061 = $signed(4'sh1) * $signed(io_in_274); // @[Modules.scala 151:80:@10289.4]
  assign _GEN_233 = {{1{_T_54871[4]}},_T_54871}; // @[Modules.scala 150:103:@10290.4]
  assign _T_64062 = $signed(_GEN_233) + $signed(_T_64061); // @[Modules.scala 150:103:@10290.4]
  assign _T_64063 = _T_64062[5:0]; // @[Modules.scala 150:103:@10291.4]
  assign _T_64064 = $signed(_T_64063); // @[Modules.scala 150:103:@10292.4]
  assign _T_64066 = $signed(4'sh1) * $signed(io_in_275); // @[Modules.scala 150:74:@10294.4]
  assign _T_64068 = $signed(4'sh1) * $signed(io_in_276); // @[Modules.scala 151:80:@10295.4]
  assign _T_64069 = $signed(_T_64066) + $signed(_T_64068); // @[Modules.scala 150:103:@10296.4]
  assign _T_64070 = _T_64069[5:0]; // @[Modules.scala 150:103:@10297.4]
  assign _T_64071 = $signed(_T_64070); // @[Modules.scala 150:103:@10298.4]
  assign _T_64073 = $signed(4'sh1) * $signed(io_in_277); // @[Modules.scala 150:74:@10300.4]
  assign _T_64075 = $signed(4'sh1) * $signed(io_in_278); // @[Modules.scala 151:80:@10301.4]
  assign _T_64076 = $signed(_T_64073) + $signed(_T_64075); // @[Modules.scala 150:103:@10302.4]
  assign _T_64077 = _T_64076[5:0]; // @[Modules.scala 150:103:@10303.4]
  assign _T_64078 = $signed(_T_64077); // @[Modules.scala 150:103:@10304.4]
  assign _GEN_234 = {{1{_T_60983[4]}},_T_60983}; // @[Modules.scala 150:103:@10314.4]
  assign _T_64090 = $signed(_T_54899) + $signed(_GEN_234); // @[Modules.scala 150:103:@10314.4]
  assign _T_64091 = _T_64090[5:0]; // @[Modules.scala 150:103:@10315.4]
  assign _T_64092 = $signed(_T_64091); // @[Modules.scala 150:103:@10316.4]
  assign _T_64097 = $signed(_T_60985) + $signed(_T_54908); // @[Modules.scala 150:103:@10320.4]
  assign _T_64098 = _T_64097[4:0]; // @[Modules.scala 150:103:@10321.4]
  assign _T_64099 = $signed(_T_64098); // @[Modules.scala 150:103:@10322.4]
  assign _T_64103 = $signed(4'sh1) * $signed(io_in_286); // @[Modules.scala 151:80:@10325.4]
  assign _GEN_235 = {{1{_T_54913[4]}},_T_54913}; // @[Modules.scala 150:103:@10326.4]
  assign _T_64104 = $signed(_GEN_235) + $signed(_T_64103); // @[Modules.scala 150:103:@10326.4]
  assign _T_64105 = _T_64104[5:0]; // @[Modules.scala 150:103:@10327.4]
  assign _T_64106 = $signed(_T_64105); // @[Modules.scala 150:103:@10328.4]
  assign _T_64108 = $signed(4'sh1) * $signed(io_in_287); // @[Modules.scala 150:74:@10330.4]
  assign _T_64111 = $signed(_T_64108) + $signed(_T_61004); // @[Modules.scala 150:103:@10332.4]
  assign _T_64112 = _T_64111[5:0]; // @[Modules.scala 150:103:@10333.4]
  assign _T_64113 = $signed(_T_64112); // @[Modules.scala 150:103:@10334.4]
  assign _T_64115 = $signed(4'sh1) * $signed(io_in_289); // @[Modules.scala 150:74:@10336.4]
  assign _T_64118 = $signed(_T_64115) + $signed(_T_61006); // @[Modules.scala 150:103:@10338.4]
  assign _T_64119 = _T_64118[5:0]; // @[Modules.scala 150:103:@10339.4]
  assign _T_64120 = $signed(_T_64119); // @[Modules.scala 150:103:@10340.4]
  assign _T_64122 = $signed(4'sh1) * $signed(io_in_291); // @[Modules.scala 150:74:@10342.4]
  assign _T_64124 = $signed(4'sh1) * $signed(io_in_292); // @[Modules.scala 151:80:@10343.4]
  assign _T_64125 = $signed(_T_64122) + $signed(_T_64124); // @[Modules.scala 150:103:@10344.4]
  assign _T_64126 = _T_64125[5:0]; // @[Modules.scala 150:103:@10345.4]
  assign _T_64127 = $signed(_T_64126); // @[Modules.scala 150:103:@10346.4]
  assign _T_64132 = $signed(_T_61013) + $signed(_T_61018); // @[Modules.scala 150:103:@10350.4]
  assign _T_64133 = _T_64132[4:0]; // @[Modules.scala 150:103:@10351.4]
  assign _T_64134 = $signed(_T_64133); // @[Modules.scala 150:103:@10352.4]
  assign _T_64139 = $signed(_T_61020) + $signed(_T_61025); // @[Modules.scala 150:103:@10356.4]
  assign _T_64140 = _T_64139[4:0]; // @[Modules.scala 150:103:@10357.4]
  assign _T_64141 = $signed(_T_64140); // @[Modules.scala 150:103:@10358.4]
  assign _T_64164 = $signed(4'sh1) * $signed(io_in_304); // @[Modules.scala 150:74:@10378.4]
  assign _T_64166 = $signed(4'sh1) * $signed(io_in_305); // @[Modules.scala 151:80:@10379.4]
  assign _T_64167 = $signed(_T_64164) + $signed(_T_64166); // @[Modules.scala 150:103:@10380.4]
  assign _T_64168 = _T_64167[5:0]; // @[Modules.scala 150:103:@10381.4]
  assign _T_64169 = $signed(_T_64168); // @[Modules.scala 150:103:@10382.4]
  assign _T_64171 = $signed(4'sh1) * $signed(io_in_306); // @[Modules.scala 150:74:@10384.4]
  assign _T_64173 = $signed(-4'sh1) * $signed(io_in_307); // @[Modules.scala 151:80:@10385.4]
  assign _GEN_236 = {{1{_T_64173[4]}},_T_64173}; // @[Modules.scala 150:103:@10386.4]
  assign _T_64174 = $signed(_T_64171) + $signed(_GEN_236); // @[Modules.scala 150:103:@10386.4]
  assign _T_64175 = _T_64174[5:0]; // @[Modules.scala 150:103:@10387.4]
  assign _T_64176 = $signed(_T_64175); // @[Modules.scala 150:103:@10388.4]
  assign _T_64181 = $signed(_T_54985) + $signed(_T_61062); // @[Modules.scala 150:103:@10392.4]
  assign _T_64182 = _T_64181[4:0]; // @[Modules.scala 150:103:@10393.4]
  assign _T_64183 = $signed(_T_64182); // @[Modules.scala 150:103:@10394.4]
  assign _T_64194 = $signed(4'sh1) * $signed(io_in_313); // @[Modules.scala 151:80:@10403.4]
  assign _T_64195 = $signed(_T_58025) + $signed(_T_64194); // @[Modules.scala 150:103:@10404.4]
  assign _T_64196 = _T_64195[5:0]; // @[Modules.scala 150:103:@10405.4]
  assign _T_64197 = $signed(_T_64196); // @[Modules.scala 150:103:@10406.4]
  assign _T_64202 = $signed(_T_58032) + $signed(_T_61081); // @[Modules.scala 150:103:@10410.4]
  assign _T_64203 = _T_64202[5:0]; // @[Modules.scala 150:103:@10411.4]
  assign _T_64204 = $signed(_T_64203); // @[Modules.scala 150:103:@10412.4]
  assign _T_64209 = $signed(_T_61083) + $signed(_T_61088); // @[Modules.scala 150:103:@10416.4]
  assign _T_64210 = _T_64209[5:0]; // @[Modules.scala 150:103:@10417.4]
  assign _T_64211 = $signed(_T_64210); // @[Modules.scala 150:103:@10418.4]
  assign _T_64216 = $signed(_T_61090) + $signed(_T_61095); // @[Modules.scala 150:103:@10422.4]
  assign _T_64217 = _T_64216[5:0]; // @[Modules.scala 150:103:@10423.4]
  assign _T_64218 = $signed(_T_64217); // @[Modules.scala 150:103:@10424.4]
  assign _T_64223 = $signed(_T_61097) + $signed(_T_58053); // @[Modules.scala 150:103:@10428.4]
  assign _T_64224 = _T_64223[5:0]; // @[Modules.scala 150:103:@10429.4]
  assign _T_64225 = $signed(_T_64224); // @[Modules.scala 150:103:@10430.4]
  assign _T_64230 = $signed(_T_58058) + $signed(_GEN_169); // @[Modules.scala 150:103:@10434.4]
  assign _T_64231 = _T_64230[5:0]; // @[Modules.scala 150:103:@10435.4]
  assign _T_64232 = $signed(_T_64231); // @[Modules.scala 150:103:@10436.4]
  assign _T_64262 = $signed(4'sh1) * $signed(io_in_333); // @[Modules.scala 150:74:@10462.4]
  assign _T_64264 = $signed(4'sh1) * $signed(io_in_334); // @[Modules.scala 151:80:@10463.4]
  assign _T_64265 = $signed(_T_64262) + $signed(_T_64264); // @[Modules.scala 150:103:@10464.4]
  assign _T_64266 = _T_64265[5:0]; // @[Modules.scala 150:103:@10465.4]
  assign _T_64267 = $signed(_T_64266); // @[Modules.scala 150:103:@10466.4]
  assign _T_64272 = $signed(_T_58100) + $signed(_GEN_29); // @[Modules.scala 150:103:@10470.4]
  assign _T_64273 = _T_64272[5:0]; // @[Modules.scala 150:103:@10471.4]
  assign _T_64274 = $signed(_T_64273); // @[Modules.scala 150:103:@10472.4]
  assign _GEN_239 = {{1{_T_61153[4]}},_T_61153}; // @[Modules.scala 150:103:@10482.4]
  assign _T_64286 = $signed(_GEN_239) + $signed(_T_58116); // @[Modules.scala 150:103:@10482.4]
  assign _T_64287 = _T_64286[5:0]; // @[Modules.scala 150:103:@10483.4]
  assign _T_64288 = $signed(_T_64287); // @[Modules.scala 150:103:@10484.4]
  assign _T_64293 = $signed(_T_58121) + $signed(_T_61160); // @[Modules.scala 150:103:@10488.4]
  assign _T_64294 = _T_64293[5:0]; // @[Modules.scala 150:103:@10489.4]
  assign _T_64295 = $signed(_T_64294); // @[Modules.scala 150:103:@10490.4]
  assign _T_64334 = $signed(-4'sh1) * $signed(io_in_356); // @[Modules.scala 151:80:@10523.4]
  assign _T_64335 = $signed(_T_55132) + $signed(_T_64334); // @[Modules.scala 150:103:@10524.4]
  assign _T_64336 = _T_64335[4:0]; // @[Modules.scala 150:103:@10525.4]
  assign _T_64337 = $signed(_T_64336); // @[Modules.scala 150:103:@10526.4]
  assign _T_64342 = $signed(_T_55139) + $signed(_T_55144); // @[Modules.scala 150:103:@10530.4]
  assign _T_64343 = _T_64342[4:0]; // @[Modules.scala 150:103:@10531.4]
  assign _T_64344 = $signed(_T_64343); // @[Modules.scala 150:103:@10532.4]
  assign _T_64349 = $signed(_T_55146) + $signed(_T_58172); // @[Modules.scala 150:103:@10536.4]
  assign _T_64350 = _T_64349[4:0]; // @[Modules.scala 150:103:@10537.4]
  assign _T_64351 = $signed(_T_64350); // @[Modules.scala 150:103:@10538.4]
  assign _T_64355 = $signed(4'sh1) * $signed(io_in_362); // @[Modules.scala 151:80:@10541.4]
  assign _T_64356 = $signed(_T_58177) + $signed(_T_64355); // @[Modules.scala 150:103:@10542.4]
  assign _T_64357 = _T_64356[5:0]; // @[Modules.scala 150:103:@10543.4]
  assign _T_64358 = $signed(_T_64357); // @[Modules.scala 150:103:@10544.4]
  assign _GEN_240 = {{1{_T_61230[4]}},_T_61230}; // @[Modules.scala 150:103:@10548.4]
  assign _T_64363 = $signed(_GEN_240) + $signed(_T_55165); // @[Modules.scala 150:103:@10548.4]
  assign _T_64364 = _T_64363[5:0]; // @[Modules.scala 150:103:@10549.4]
  assign _T_64365 = $signed(_T_64364); // @[Modules.scala 150:103:@10550.4]
  assign _T_64377 = $signed(_T_58200) + $signed(_T_58205); // @[Modules.scala 150:103:@10560.4]
  assign _T_64378 = _T_64377[5:0]; // @[Modules.scala 150:103:@10561.4]
  assign _T_64379 = $signed(_T_64378); // @[Modules.scala 150:103:@10562.4]
  assign _T_64412 = $signed(_T_55214) + $signed(_T_58233); // @[Modules.scala 150:103:@10590.4]
  assign _T_64413 = _T_64412[5:0]; // @[Modules.scala 150:103:@10591.4]
  assign _T_64414 = $signed(_T_64413); // @[Modules.scala 150:103:@10592.4]
  assign _T_64433 = $signed(_T_58249) + $signed(_T_61305); // @[Modules.scala 150:103:@10608.4]
  assign _T_64434 = _T_64433[5:0]; // @[Modules.scala 150:103:@10609.4]
  assign _T_64435 = $signed(_T_64434); // @[Modules.scala 150:103:@10610.4]
  assign _T_64440 = $signed(_T_55228) + $signed(_T_58261); // @[Modules.scala 150:103:@10614.4]
  assign _T_64441 = _T_64440[4:0]; // @[Modules.scala 150:103:@10615.4]
  assign _T_64442 = $signed(_T_64441); // @[Modules.scala 150:103:@10616.4]
  assign _T_64447 = $signed(_T_58263) + $signed(_T_55237); // @[Modules.scala 150:103:@10620.4]
  assign _T_64448 = _T_64447[4:0]; // @[Modules.scala 150:103:@10621.4]
  assign _T_64449 = $signed(_T_64448); // @[Modules.scala 150:103:@10622.4]
  assign _T_64454 = $signed(_GEN_37) + $signed(_T_55249); // @[Modules.scala 150:103:@10626.4]
  assign _T_64455 = _T_64454[5:0]; // @[Modules.scala 150:103:@10627.4]
  assign _T_64456 = $signed(_T_64455); // @[Modules.scala 150:103:@10628.4]
  assign _T_64458 = $signed(-4'sh1) * $signed(io_in_394); // @[Modules.scala 150:74:@10630.4]
  assign _GEN_242 = {{1{_T_64458[4]}},_T_64458}; // @[Modules.scala 150:103:@10632.4]
  assign _T_64461 = $signed(_GEN_242) + $signed(_T_58289); // @[Modules.scala 150:103:@10632.4]
  assign _T_64462 = _T_64461[5:0]; // @[Modules.scala 150:103:@10633.4]
  assign _T_64463 = $signed(_T_64462); // @[Modules.scala 150:103:@10634.4]
  assign _T_64489 = $signed(_T_61370) + $signed(_T_58310); // @[Modules.scala 150:103:@10656.4]
  assign _T_64490 = _T_64489[5:0]; // @[Modules.scala 150:103:@10657.4]
  assign _T_64491 = $signed(_T_64490); // @[Modules.scala 150:103:@10658.4]
  assign _T_64496 = $signed(_T_55293) + $signed(_T_55298); // @[Modules.scala 150:103:@10662.4]
  assign _T_64497 = _T_64496[5:0]; // @[Modules.scala 150:103:@10663.4]
  assign _T_64498 = $signed(_T_64497); // @[Modules.scala 150:103:@10664.4]
  assign _GEN_243 = {{1{_T_58333[4]}},_T_58333}; // @[Modules.scala 150:103:@10674.4]
  assign _T_64510 = $signed(_T_61391) + $signed(_GEN_243); // @[Modules.scala 150:103:@10674.4]
  assign _T_64511 = _T_64510[5:0]; // @[Modules.scala 150:103:@10675.4]
  assign _T_64512 = $signed(_T_64511); // @[Modules.scala 150:103:@10676.4]
  assign _T_64531 = $signed(_T_55328) + $signed(_T_55335); // @[Modules.scala 150:103:@10692.4]
  assign _T_64532 = _T_64531[5:0]; // @[Modules.scala 150:103:@10693.4]
  assign _T_64533 = $signed(_T_64532); // @[Modules.scala 150:103:@10694.4]
  assign _GEN_245 = {{1{_T_55347[4]}},_T_55347}; // @[Modules.scala 150:103:@10704.4]
  assign _T_64545 = $signed(_GEN_245) + $signed(_T_61438); // @[Modules.scala 150:103:@10704.4]
  assign _T_64546 = _T_64545[5:0]; // @[Modules.scala 150:103:@10705.4]
  assign _T_64547 = $signed(_T_64546); // @[Modules.scala 150:103:@10706.4]
  assign _T_64549 = $signed(4'sh1) * $signed(io_in_428); // @[Modules.scala 150:74:@10708.4]
  assign _T_64552 = $signed(_T_64549) + $signed(_T_55363); // @[Modules.scala 150:103:@10710.4]
  assign _T_64553 = _T_64552[5:0]; // @[Modules.scala 150:103:@10711.4]
  assign _T_64554 = $signed(_T_64553); // @[Modules.scala 150:103:@10712.4]
  assign _T_64573 = $signed(_T_55382) + $signed(_T_61473); // @[Modules.scala 150:103:@10728.4]
  assign _T_64574 = _T_64573[4:0]; // @[Modules.scala 150:103:@10729.4]
  assign _T_64575 = $signed(_T_64574); // @[Modules.scala 150:103:@10730.4]
  assign _T_64579 = $signed(-4'sh1) * $signed(io_in_440); // @[Modules.scala 151:80:@10733.4]
  assign _T_64580 = $signed(_T_61475) + $signed(_T_64579); // @[Modules.scala 150:103:@10734.4]
  assign _T_64581 = _T_64580[4:0]; // @[Modules.scala 150:103:@10735.4]
  assign _T_64582 = $signed(_T_64581); // @[Modules.scala 150:103:@10736.4]
  assign _T_64587 = $signed(_T_58401) + $signed(_T_55398); // @[Modules.scala 150:103:@10740.4]
  assign _T_64588 = _T_64587[4:0]; // @[Modules.scala 150:103:@10741.4]
  assign _T_64589 = $signed(_T_64588); // @[Modules.scala 150:103:@10742.4]
  assign _T_64608 = $signed(_T_61496) + $signed(_T_55417); // @[Modules.scala 150:103:@10758.4]
  assign _T_64609 = _T_64608[4:0]; // @[Modules.scala 150:103:@10759.4]
  assign _T_64610 = $signed(_T_64609); // @[Modules.scala 150:103:@10760.4]
  assign _T_64614 = $signed(-4'sh1) * $signed(io_in_450); // @[Modules.scala 151:80:@10763.4]
  assign _T_64615 = $signed(_T_55419) + $signed(_T_64614); // @[Modules.scala 150:103:@10764.4]
  assign _T_64616 = _T_64615[4:0]; // @[Modules.scala 150:103:@10765.4]
  assign _T_64617 = $signed(_T_64616); // @[Modules.scala 150:103:@10766.4]
  assign _T_64622 = $signed(_T_61510) + $signed(_T_55431); // @[Modules.scala 150:103:@10770.4]
  assign _T_64623 = _T_64622[4:0]; // @[Modules.scala 150:103:@10771.4]
  assign _T_64624 = $signed(_T_64623); // @[Modules.scala 150:103:@10772.4]
  assign _T_64635 = $signed(4'sh1) * $signed(io_in_456); // @[Modules.scala 151:80:@10781.4]
  assign _GEN_247 = {{1{_T_58450[4]}},_T_58450}; // @[Modules.scala 150:103:@10782.4]
  assign _T_64636 = $signed(_GEN_247) + $signed(_T_64635); // @[Modules.scala 150:103:@10782.4]
  assign _T_64637 = _T_64636[5:0]; // @[Modules.scala 150:103:@10783.4]
  assign _T_64638 = $signed(_T_64637); // @[Modules.scala 150:103:@10784.4]
  assign _T_64643 = $signed(_T_55440) + $signed(_T_55445); // @[Modules.scala 150:103:@10788.4]
  assign _T_64644 = _T_64643[5:0]; // @[Modules.scala 150:103:@10789.4]
  assign _T_64645 = $signed(_T_64644); // @[Modules.scala 150:103:@10790.4]
  assign _T_64649 = $signed(4'sh1) * $signed(io_in_460); // @[Modules.scala 151:80:@10793.4]
  assign _T_64650 = $signed(_T_55447) + $signed(_T_64649); // @[Modules.scala 150:103:@10794.4]
  assign _T_64651 = _T_64650[5:0]; // @[Modules.scala 150:103:@10795.4]
  assign _T_64652 = $signed(_T_64651); // @[Modules.scala 150:103:@10796.4]
  assign _T_64671 = $signed(_T_55466) + $signed(_T_61552); // @[Modules.scala 150:103:@10812.4]
  assign _T_64672 = _T_64671[4:0]; // @[Modules.scala 150:103:@10813.4]
  assign _T_64673 = $signed(_T_64672); // @[Modules.scala 150:103:@10814.4]
  assign _T_64675 = $signed(-4'sh1) * $signed(io_in_468); // @[Modules.scala 150:74:@10816.4]
  assign _T_64677 = $signed(-4'sh1) * $signed(io_in_469); // @[Modules.scala 151:80:@10817.4]
  assign _T_64678 = $signed(_T_64675) + $signed(_T_64677); // @[Modules.scala 150:103:@10818.4]
  assign _T_64679 = _T_64678[4:0]; // @[Modules.scala 150:103:@10819.4]
  assign _T_64680 = $signed(_T_64679); // @[Modules.scala 150:103:@10820.4]
  assign _T_64699 = $signed(_T_61573) + $signed(_T_61578); // @[Modules.scala 150:103:@10836.4]
  assign _T_64700 = _T_64699[4:0]; // @[Modules.scala 150:103:@10837.4]
  assign _T_64701 = $signed(_T_64700); // @[Modules.scala 150:103:@10838.4]
  assign _GEN_249 = {{1{_T_61585[4]}},_T_61585}; // @[Modules.scala 150:103:@10842.4]
  assign _T_64706 = $signed(_T_61580) + $signed(_GEN_249); // @[Modules.scala 150:103:@10842.4]
  assign _T_64707 = _T_64706[5:0]; // @[Modules.scala 150:103:@10843.4]
  assign _T_64708 = $signed(_T_64707); // @[Modules.scala 150:103:@10844.4]
  assign _T_64713 = $signed(_T_61587) + $signed(_T_61592); // @[Modules.scala 150:103:@10848.4]
  assign _T_64714 = _T_64713[4:0]; // @[Modules.scala 150:103:@10849.4]
  assign _T_64715 = $signed(_T_64714); // @[Modules.scala 150:103:@10850.4]
  assign _T_64720 = $signed(_T_58520) + $signed(_T_58527); // @[Modules.scala 150:103:@10854.4]
  assign _T_64721 = _T_64720[4:0]; // @[Modules.scala 150:103:@10855.4]
  assign _T_64722 = $signed(_T_64721); // @[Modules.scala 150:103:@10856.4]
  assign _T_64726 = $signed(4'sh1) * $signed(io_in_485); // @[Modules.scala 151:80:@10859.4]
  assign _T_64727 = $signed(_T_61606) + $signed(_T_64726); // @[Modules.scala 150:103:@10860.4]
  assign _T_64728 = _T_64727[5:0]; // @[Modules.scala 150:103:@10861.4]
  assign _T_64729 = $signed(_T_64728); // @[Modules.scala 150:103:@10862.4]
  assign _T_64748 = $signed(_T_55522) + $signed(_GEN_115); // @[Modules.scala 150:103:@10878.4]
  assign _T_64749 = _T_64748[5:0]; // @[Modules.scala 150:103:@10879.4]
  assign _T_64750 = $signed(_T_64749); // @[Modules.scala 150:103:@10880.4]
  assign _T_64754 = $signed(-4'sh1) * $signed(io_in_497); // @[Modules.scala 151:80:@10883.4]
  assign _T_64755 = $signed(_T_58562) + $signed(_T_64754); // @[Modules.scala 150:103:@10884.4]
  assign _T_64756 = _T_64755[4:0]; // @[Modules.scala 150:103:@10885.4]
  assign _T_64757 = $signed(_T_64756); // @[Modules.scala 150:103:@10886.4]
  assign _T_64768 = $signed(-4'sh1) * $signed(io_in_502); // @[Modules.scala 151:80:@10895.4]
  assign _T_64769 = $signed(_T_58578) + $signed(_T_64768); // @[Modules.scala 150:103:@10896.4]
  assign _T_64770 = _T_64769[4:0]; // @[Modules.scala 150:103:@10897.4]
  assign _T_64771 = $signed(_T_64770); // @[Modules.scala 150:103:@10898.4]
  assign _GEN_251 = {{1{_T_61643[4]}},_T_61643}; // @[Modules.scala 150:103:@10902.4]
  assign _T_64776 = $signed(_GEN_251) + $signed(_T_58590); // @[Modules.scala 150:103:@10902.4]
  assign _T_64777 = _T_64776[5:0]; // @[Modules.scala 150:103:@10903.4]
  assign _T_64778 = $signed(_T_64777); // @[Modules.scala 150:103:@10904.4]
  assign _T_64782 = $signed(-4'sh1) * $signed(io_in_506); // @[Modules.scala 151:80:@10907.4]
  assign _GEN_252 = {{1{_T_64782[4]}},_T_64782}; // @[Modules.scala 150:103:@10908.4]
  assign _T_64783 = $signed(_T_55564) + $signed(_GEN_252); // @[Modules.scala 150:103:@10908.4]
  assign _T_64784 = _T_64783[5:0]; // @[Modules.scala 150:103:@10909.4]
  assign _T_64785 = $signed(_T_64784); // @[Modules.scala 150:103:@10910.4]
  assign _T_64790 = $signed(_T_61657) + $signed(_T_61662); // @[Modules.scala 150:103:@10914.4]
  assign _T_64791 = _T_64790[4:0]; // @[Modules.scala 150:103:@10915.4]
  assign _T_64792 = $signed(_T_64791); // @[Modules.scala 150:103:@10916.4]
  assign _T_64796 = $signed(4'sh1) * $signed(io_in_510); // @[Modules.scala 151:80:@10919.4]
  assign _T_64797 = $signed(_GEN_117) + $signed(_T_64796); // @[Modules.scala 150:103:@10920.4]
  assign _T_64798 = _T_64797[5:0]; // @[Modules.scala 150:103:@10921.4]
  assign _T_64799 = $signed(_T_64798); // @[Modules.scala 150:103:@10922.4]
  assign _GEN_254 = {{1{_T_58606[4]}},_T_58606}; // @[Modules.scala 150:103:@10926.4]
  assign _T_64804 = $signed(_GEN_254) + $signed(_T_55587); // @[Modules.scala 150:103:@10926.4]
  assign _T_64805 = _T_64804[5:0]; // @[Modules.scala 150:103:@10927.4]
  assign _T_64806 = $signed(_T_64805); // @[Modules.scala 150:103:@10928.4]
  assign _T_64825 = $signed(_T_58632) + $signed(_GEN_189); // @[Modules.scala 150:103:@10944.4]
  assign _T_64826 = _T_64825[5:0]; // @[Modules.scala 150:103:@10945.4]
  assign _T_64827 = $signed(_T_64826); // @[Modules.scala 150:103:@10946.4]
  assign _T_64829 = $signed(-4'sh1) * $signed(io_in_522); // @[Modules.scala 150:74:@10948.4]
  assign _T_64831 = $signed(-4'sh1) * $signed(io_in_523); // @[Modules.scala 151:80:@10949.4]
  assign _T_64832 = $signed(_T_64829) + $signed(_T_64831); // @[Modules.scala 150:103:@10950.4]
  assign _T_64833 = _T_64832[4:0]; // @[Modules.scala 150:103:@10951.4]
  assign _T_64834 = $signed(_T_64833); // @[Modules.scala 150:103:@10952.4]
  assign _T_64838 = $signed(-4'sh1) * $signed(io_in_525); // @[Modules.scala 151:80:@10955.4]
  assign _GEN_256 = {{1{_T_64838[4]}},_T_64838}; // @[Modules.scala 150:103:@10956.4]
  assign _T_64839 = $signed(_T_55622) + $signed(_GEN_256); // @[Modules.scala 150:103:@10956.4]
  assign _T_64840 = _T_64839[5:0]; // @[Modules.scala 150:103:@10957.4]
  assign _T_64841 = $signed(_T_64840); // @[Modules.scala 150:103:@10958.4]
  assign _T_64846 = $signed(_T_61706) + $signed(_T_58639); // @[Modules.scala 150:103:@10962.4]
  assign _T_64847 = _T_64846[4:0]; // @[Modules.scala 150:103:@10963.4]
  assign _T_64848 = $signed(_T_64847); // @[Modules.scala 150:103:@10964.4]
  assign _T_64853 = $signed(_T_58641) + $signed(_T_58646); // @[Modules.scala 150:103:@10968.4]
  assign _T_64854 = _T_64853[4:0]; // @[Modules.scala 150:103:@10969.4]
  assign _T_64855 = $signed(_T_64854); // @[Modules.scala 150:103:@10970.4]
  assign _GEN_257 = {{1{_T_58648[4]}},_T_58648}; // @[Modules.scala 150:103:@10974.4]
  assign _T_64860 = $signed(_GEN_257) + $signed(_T_55643); // @[Modules.scala 150:103:@10974.4]
  assign _T_64861 = _T_64860[5:0]; // @[Modules.scala 150:103:@10975.4]
  assign _T_64862 = $signed(_T_64861); // @[Modules.scala 150:103:@10976.4]
  assign _T_64867 = $signed(_T_58655) + $signed(_GEN_119); // @[Modules.scala 150:103:@10980.4]
  assign _T_64868 = _T_64867[5:0]; // @[Modules.scala 150:103:@10981.4]
  assign _T_64869 = $signed(_T_64868); // @[Modules.scala 150:103:@10982.4]
  assign _T_64871 = $signed(-4'sh1) * $signed(io_in_534); // @[Modules.scala 150:74:@10984.4]
  assign _T_64874 = $signed(_T_64871) + $signed(_T_61739); // @[Modules.scala 150:103:@10986.4]
  assign _T_64875 = _T_64874[4:0]; // @[Modules.scala 150:103:@10987.4]
  assign _T_64876 = $signed(_T_64875); // @[Modules.scala 150:103:@10988.4]
  assign _T_64881 = $signed(_T_61741) + $signed(_T_58674); // @[Modules.scala 150:103:@10992.4]
  assign _T_64882 = _T_64881[4:0]; // @[Modules.scala 150:103:@10993.4]
  assign _T_64883 = $signed(_T_64882); // @[Modules.scala 150:103:@10994.4]
  assign _T_64888 = $signed(_T_58676) + $signed(_T_58683); // @[Modules.scala 150:103:@10998.4]
  assign _T_64889 = _T_64888[4:0]; // @[Modules.scala 150:103:@10999.4]
  assign _T_64890 = $signed(_T_64889); // @[Modules.scala 150:103:@11000.4]
  assign _T_64906 = $signed(-4'sh1) * $signed(io_in_547); // @[Modules.scala 150:74:@11014.4]
  assign _T_64909 = $signed(_T_64906) + $signed(_T_58704); // @[Modules.scala 150:103:@11016.4]
  assign _T_64910 = _T_64909[4:0]; // @[Modules.scala 150:103:@11017.4]
  assign _T_64911 = $signed(_T_64910); // @[Modules.scala 150:103:@11018.4]
  assign _T_64920 = $signed(-4'sh1) * $signed(io_in_551); // @[Modules.scala 150:74:@11026.4]
  assign _GEN_259 = {{1{_T_64920[4]}},_T_64920}; // @[Modules.scala 150:103:@11028.4]
  assign _T_64923 = $signed(_GEN_259) + $signed(_T_55711); // @[Modules.scala 150:103:@11028.4]
  assign _T_64924 = _T_64923[5:0]; // @[Modules.scala 150:103:@11029.4]
  assign _T_64925 = $signed(_T_64924); // @[Modules.scala 150:103:@11030.4]
  assign _T_64930 = $signed(_T_58718) + $signed(_T_58723); // @[Modules.scala 150:103:@11034.4]
  assign _T_64931 = _T_64930[4:0]; // @[Modules.scala 150:103:@11035.4]
  assign _T_64932 = $signed(_T_64931); // @[Modules.scala 150:103:@11036.4]
  assign _GEN_260 = {{1{_T_58732[4]}},_T_58732}; // @[Modules.scala 150:103:@11040.4]
  assign _T_64937 = $signed(_T_55713) + $signed(_GEN_260); // @[Modules.scala 150:103:@11040.4]
  assign _T_64938 = _T_64937[5:0]; // @[Modules.scala 150:103:@11041.4]
  assign _T_64939 = $signed(_T_64938); // @[Modules.scala 150:103:@11042.4]
  assign _T_64943 = $signed(4'sh1) * $signed(io_in_559); // @[Modules.scala 151:80:@11045.4]
  assign _GEN_261 = {{1{_T_58737[4]}},_T_58737}; // @[Modules.scala 150:103:@11046.4]
  assign _T_64944 = $signed(_GEN_261) + $signed(_T_64943); // @[Modules.scala 150:103:@11046.4]
  assign _T_64945 = _T_64944[5:0]; // @[Modules.scala 150:103:@11047.4]
  assign _T_64946 = $signed(_T_64945); // @[Modules.scala 150:103:@11048.4]
  assign _T_64948 = $signed(-4'sh1) * $signed(io_in_561); // @[Modules.scala 150:74:@11050.4]
  assign _T_64950 = $signed(-4'sh1) * $signed(io_in_562); // @[Modules.scala 151:80:@11051.4]
  assign _T_64951 = $signed(_T_64948) + $signed(_T_64950); // @[Modules.scala 150:103:@11052.4]
  assign _T_64952 = _T_64951[4:0]; // @[Modules.scala 150:103:@11053.4]
  assign _T_64953 = $signed(_T_64952); // @[Modules.scala 150:103:@11054.4]
  assign _T_64969 = $signed(4'sh1) * $signed(io_in_568); // @[Modules.scala 150:74:@11068.4]
  assign _GEN_262 = {{1{_T_61839[4]}},_T_61839}; // @[Modules.scala 150:103:@11070.4]
  assign _T_64972 = $signed(_T_64969) + $signed(_GEN_262); // @[Modules.scala 150:103:@11070.4]
  assign _T_64973 = _T_64972[5:0]; // @[Modules.scala 150:103:@11071.4]
  assign _T_64974 = $signed(_T_64973); // @[Modules.scala 150:103:@11072.4]
  assign _T_64979 = $signed(_T_58760) + $signed(_T_58765); // @[Modules.scala 150:103:@11076.4]
  assign _T_64980 = _T_64979[4:0]; // @[Modules.scala 150:103:@11077.4]
  assign _T_64981 = $signed(_T_64980); // @[Modules.scala 150:103:@11078.4]
  assign _T_64985 = $signed(-4'sh1) * $signed(io_in_574); // @[Modules.scala 151:80:@11081.4]
  assign _T_64986 = $signed(_T_58767) + $signed(_T_64985); // @[Modules.scala 150:103:@11082.4]
  assign _T_64987 = _T_64986[4:0]; // @[Modules.scala 150:103:@11083.4]
  assign _T_64988 = $signed(_T_64987); // @[Modules.scala 150:103:@11084.4]
  assign _T_65004 = $signed(4'sh1) * $signed(io_in_582); // @[Modules.scala 150:74:@11098.4]
  assign _T_65007 = $signed(_T_65004) + $signed(_GEN_124); // @[Modules.scala 150:103:@11100.4]
  assign _T_65008 = _T_65007[5:0]; // @[Modules.scala 150:103:@11101.4]
  assign _T_65009 = $signed(_T_65008); // @[Modules.scala 150:103:@11102.4]
  assign _T_65028 = $signed(_T_61895) + $signed(_T_61900); // @[Modules.scala 150:103:@11118.4]
  assign _T_65029 = _T_65028[4:0]; // @[Modules.scala 150:103:@11119.4]
  assign _T_65030 = $signed(_T_65029); // @[Modules.scala 150:103:@11120.4]
  assign _T_65035 = $signed(_T_61902) + $signed(_T_61907); // @[Modules.scala 150:103:@11124.4]
  assign _T_65036 = _T_65035[4:0]; // @[Modules.scala 150:103:@11125.4]
  assign _T_65037 = $signed(_T_65036); // @[Modules.scala 150:103:@11126.4]
  assign _T_65048 = $signed(-4'sh1) * $signed(io_in_604); // @[Modules.scala 151:80:@11135.4]
  assign _GEN_265 = {{1{_T_65048[4]}},_T_65048}; // @[Modules.scala 150:103:@11136.4]
  assign _T_65049 = $signed(_T_55825) + $signed(_GEN_265); // @[Modules.scala 150:103:@11136.4]
  assign _T_65050 = _T_65049[5:0]; // @[Modules.scala 150:103:@11137.4]
  assign _T_65051 = $signed(_T_65050); // @[Modules.scala 150:103:@11138.4]
  assign _T_65056 = $signed(_T_58851) + $signed(_T_61944); // @[Modules.scala 150:103:@11142.4]
  assign _T_65057 = _T_65056[4:0]; // @[Modules.scala 150:103:@11143.4]
  assign _T_65058 = $signed(_T_65057); // @[Modules.scala 150:103:@11144.4]
  assign _T_65063 = $signed(_GEN_65) + $signed(_T_55844); // @[Modules.scala 150:103:@11148.4]
  assign _T_65064 = _T_65063[5:0]; // @[Modules.scala 150:103:@11149.4]
  assign _T_65065 = $signed(_T_65064); // @[Modules.scala 150:103:@11150.4]
  assign _T_65074 = $signed(-4'sh1) * $signed(io_in_614); // @[Modules.scala 150:74:@11158.4]
  assign _GEN_267 = {{1{_T_65074[4]}},_T_65074}; // @[Modules.scala 150:103:@11160.4]
  assign _T_65077 = $signed(_GEN_267) + $signed(_T_55860); // @[Modules.scala 150:103:@11160.4]
  assign _T_65078 = _T_65077[5:0]; // @[Modules.scala 150:103:@11161.4]
  assign _T_65079 = $signed(_T_65078); // @[Modules.scala 150:103:@11162.4]
  assign _T_65083 = $signed(-4'sh1) * $signed(io_in_618); // @[Modules.scala 151:80:@11165.4]
  assign _GEN_268 = {{1{_T_65083[4]}},_T_65083}; // @[Modules.scala 150:103:@11166.4]
  assign _T_65084 = $signed(_T_55865) + $signed(_GEN_268); // @[Modules.scala 150:103:@11166.4]
  assign _T_65085 = _T_65084[5:0]; // @[Modules.scala 150:103:@11167.4]
  assign _T_65086 = $signed(_T_65085); // @[Modules.scala 150:103:@11168.4]
  assign _T_65091 = $signed(_T_61979) + $signed(_T_61984); // @[Modules.scala 150:103:@11172.4]
  assign _T_65092 = _T_65091[4:0]; // @[Modules.scala 150:103:@11173.4]
  assign _T_65093 = $signed(_T_65092); // @[Modules.scala 150:103:@11174.4]
  assign _T_65098 = $signed(_T_61986) + $signed(_T_61991); // @[Modules.scala 150:103:@11178.4]
  assign _T_65099 = _T_65098[4:0]; // @[Modules.scala 150:103:@11179.4]
  assign _T_65100 = $signed(_T_65099); // @[Modules.scala 150:103:@11180.4]
  assign _T_65105 = $signed(_T_55886) + $signed(_T_61998); // @[Modules.scala 150:103:@11184.4]
  assign _T_65106 = _T_65105[4:0]; // @[Modules.scala 150:103:@11185.4]
  assign _T_65107 = $signed(_T_65106); // @[Modules.scala 150:103:@11186.4]
  assign _T_65112 = $signed(_T_62000) + $signed(_T_62005); // @[Modules.scala 150:103:@11190.4]
  assign _T_65113 = _T_65112[4:0]; // @[Modules.scala 150:103:@11191.4]
  assign _T_65114 = $signed(_T_65113); // @[Modules.scala 150:103:@11192.4]
  assign _T_65125 = $signed(4'sh1) * $signed(io_in_631); // @[Modules.scala 151:80:@11201.4]
  assign _GEN_269 = {{1{_T_55900[4]}},_T_55900}; // @[Modules.scala 150:103:@11202.4]
  assign _T_65126 = $signed(_GEN_269) + $signed(_T_65125); // @[Modules.scala 150:103:@11202.4]
  assign _T_65127 = _T_65126[5:0]; // @[Modules.scala 150:103:@11203.4]
  assign _T_65128 = $signed(_T_65127); // @[Modules.scala 150:103:@11204.4]
  assign _T_65130 = $signed(4'sh1) * $signed(io_in_632); // @[Modules.scala 150:74:@11206.4]
  assign _T_65133 = $signed(_T_65130) + $signed(_T_58933); // @[Modules.scala 150:103:@11208.4]
  assign _T_65134 = _T_65133[5:0]; // @[Modules.scala 150:103:@11209.4]
  assign _T_65135 = $signed(_T_65134); // @[Modules.scala 150:103:@11210.4]
  assign _T_65140 = $signed(_T_62026) + $signed(_T_55921); // @[Modules.scala 150:103:@11214.4]
  assign _T_65141 = _T_65140[5:0]; // @[Modules.scala 150:103:@11215.4]
  assign _T_65142 = $signed(_T_65141); // @[Modules.scala 150:103:@11216.4]
  assign _GEN_270 = {{1{_T_58940[4]}},_T_58940}; // @[Modules.scala 150:103:@11220.4]
  assign _T_65147 = $signed(_GEN_270) + $signed(_T_55928); // @[Modules.scala 150:103:@11220.4]
  assign _T_65148 = _T_65147[5:0]; // @[Modules.scala 150:103:@11221.4]
  assign _T_65149 = $signed(_T_65148); // @[Modules.scala 150:103:@11222.4]
  assign _GEN_271 = {{1{_T_58949[4]}},_T_58949}; // @[Modules.scala 150:103:@11226.4]
  assign _T_65154 = $signed(_T_55930) + $signed(_GEN_271); // @[Modules.scala 150:103:@11226.4]
  assign _T_65155 = _T_65154[5:0]; // @[Modules.scala 150:103:@11227.4]
  assign _T_65156 = $signed(_T_65155); // @[Modules.scala 150:103:@11228.4]
  assign _T_65160 = $signed(-4'sh1) * $signed(io_in_641); // @[Modules.scala 151:80:@11231.4]
  assign _T_65161 = $signed(_T_58954) + $signed(_T_65160); // @[Modules.scala 150:103:@11232.4]
  assign _T_65162 = _T_65161[4:0]; // @[Modules.scala 150:103:@11233.4]
  assign _T_65163 = $signed(_T_65162); // @[Modules.scala 150:103:@11234.4]
  assign _T_65165 = $signed(-4'sh1) * $signed(io_in_642); // @[Modules.scala 150:74:@11236.4]
  assign _T_65168 = $signed(_T_65165) + $signed(_T_62049); // @[Modules.scala 150:103:@11238.4]
  assign _T_65169 = _T_65168[4:0]; // @[Modules.scala 150:103:@11239.4]
  assign _T_65170 = $signed(_T_65169); // @[Modules.scala 150:103:@11240.4]
  assign _T_65188 = $signed(4'sh1) * $signed(io_in_656); // @[Modules.scala 151:80:@11255.4]
  assign _T_65189 = $signed(_T_58984) + $signed(_T_65188); // @[Modules.scala 150:103:@11256.4]
  assign _T_65190 = _T_65189[5:0]; // @[Modules.scala 150:103:@11257.4]
  assign _T_65191 = $signed(_T_65190); // @[Modules.scala 150:103:@11258.4]
  assign _T_65193 = $signed(4'sh1) * $signed(io_in_658); // @[Modules.scala 150:74:@11260.4]
  assign _T_65195 = $signed(4'sh1) * $signed(io_in_659); // @[Modules.scala 151:80:@11261.4]
  assign _T_65196 = $signed(_T_65193) + $signed(_T_65195); // @[Modules.scala 150:103:@11262.4]
  assign _T_65197 = _T_65196[5:0]; // @[Modules.scala 150:103:@11263.4]
  assign _T_65198 = $signed(_T_65197); // @[Modules.scala 150:103:@11264.4]
  assign _T_65200 = $signed(4'sh1) * $signed(io_in_660); // @[Modules.scala 150:74:@11266.4]
  assign _T_65203 = $signed(_T_65200) + $signed(_T_59003); // @[Modules.scala 150:103:@11268.4]
  assign _T_65204 = _T_65203[5:0]; // @[Modules.scala 150:103:@11269.4]
  assign _T_65205 = $signed(_T_65204); // @[Modules.scala 150:103:@11270.4]
  assign _T_65221 = $signed(4'sh1) * $signed(io_in_666); // @[Modules.scala 150:74:@11284.4]
  assign _T_65224 = $signed(_T_65221) + $signed(_GEN_133); // @[Modules.scala 150:103:@11286.4]
  assign _T_65225 = _T_65224[5:0]; // @[Modules.scala 150:103:@11287.4]
  assign _T_65226 = $signed(_T_65225); // @[Modules.scala 150:103:@11288.4]
  assign _T_65230 = $signed(-4'sh1) * $signed(io_in_670); // @[Modules.scala 151:80:@11291.4]
  assign _T_65231 = $signed(_T_62126) + $signed(_T_65230); // @[Modules.scala 150:103:@11292.4]
  assign _T_65232 = _T_65231[4:0]; // @[Modules.scala 150:103:@11293.4]
  assign _T_65233 = $signed(_T_65232); // @[Modules.scala 150:103:@11294.4]
  assign _GEN_273 = {{1{_T_62138[4]}},_T_62138}; // @[Modules.scala 150:103:@11298.4]
  assign _T_65238 = $signed(_T_59033) + $signed(_GEN_273); // @[Modules.scala 150:103:@11298.4]
  assign _T_65239 = _T_65238[5:0]; // @[Modules.scala 150:103:@11299.4]
  assign _T_65240 = $signed(_T_65239); // @[Modules.scala 150:103:@11300.4]
  assign _T_65245 = $signed(_T_62140) + $signed(_T_62145); // @[Modules.scala 150:103:@11304.4]
  assign _T_65246 = _T_65245[4:0]; // @[Modules.scala 150:103:@11305.4]
  assign _T_65247 = $signed(_T_65246); // @[Modules.scala 150:103:@11306.4]
  assign _T_65251 = $signed(-4'sh1) * $signed(io_in_679); // @[Modules.scala 151:80:@11309.4]
  assign _T_65252 = $signed(_T_62147) + $signed(_T_65251); // @[Modules.scala 150:103:@11310.4]
  assign _T_65253 = _T_65252[4:0]; // @[Modules.scala 150:103:@11311.4]
  assign _T_65254 = $signed(_T_65253); // @[Modules.scala 150:103:@11312.4]
  assign _T_65259 = $signed(_T_56049) + $signed(_T_56054); // @[Modules.scala 150:103:@11316.4]
  assign _T_65260 = _T_65259[4:0]; // @[Modules.scala 150:103:@11317.4]
  assign _T_65261 = $signed(_T_65260); // @[Modules.scala 150:103:@11318.4]
  assign _T_65265 = $signed(-4'sh1) * $signed(io_in_683); // @[Modules.scala 151:80:@11321.4]
  assign _T_65266 = $signed(_T_56056) + $signed(_T_65265); // @[Modules.scala 150:103:@11322.4]
  assign _T_65267 = _T_65266[4:0]; // @[Modules.scala 150:103:@11323.4]
  assign _T_65268 = $signed(_T_65267); // @[Modules.scala 150:103:@11324.4]
  assign _T_65280 = $signed(_T_56063) + $signed(_T_56068); // @[Modules.scala 150:103:@11334.4]
  assign _T_65281 = _T_65280[4:0]; // @[Modules.scala 150:103:@11335.4]
  assign _T_65282 = $signed(_T_65281); // @[Modules.scala 150:103:@11336.4]
  assign _GEN_274 = {{1{_T_56070[4]}},_T_56070}; // @[Modules.scala 150:103:@11340.4]
  assign _T_65287 = $signed(_GEN_274) + $signed(_T_59082); // @[Modules.scala 150:103:@11340.4]
  assign _T_65288 = _T_65287[5:0]; // @[Modules.scala 150:103:@11341.4]
  assign _T_65289 = $signed(_T_65288); // @[Modules.scala 150:103:@11342.4]
  assign _T_65301 = $signed(_T_59094) + $signed(_T_62187); // @[Modules.scala 150:103:@11352.4]
  assign _T_65302 = _T_65301[5:0]; // @[Modules.scala 150:103:@11353.4]
  assign _T_65303 = $signed(_T_65302); // @[Modules.scala 150:103:@11354.4]
  assign _T_65308 = $signed(_T_62189) + $signed(_T_62194); // @[Modules.scala 150:103:@11358.4]
  assign _T_65309 = _T_65308[5:0]; // @[Modules.scala 150:103:@11359.4]
  assign _T_65310 = $signed(_T_65309); // @[Modules.scala 150:103:@11360.4]
  assign _T_65314 = $signed(-4'sh1) * $signed(io_in_697); // @[Modules.scala 151:80:@11363.4]
  assign _GEN_275 = {{1{_T_65314[4]}},_T_65314}; // @[Modules.scala 150:103:@11364.4]
  assign _T_65315 = $signed(_T_56098) + $signed(_GEN_275); // @[Modules.scala 150:103:@11364.4]
  assign _T_65316 = _T_65315[5:0]; // @[Modules.scala 150:103:@11365.4]
  assign _T_65317 = $signed(_T_65316); // @[Modules.scala 150:103:@11366.4]
  assign _T_65329 = $signed(_T_56117) + $signed(_GEN_209); // @[Modules.scala 150:103:@11376.4]
  assign _T_65330 = _T_65329[5:0]; // @[Modules.scala 150:103:@11377.4]
  assign _T_65331 = $signed(_T_65330); // @[Modules.scala 150:103:@11378.4]
  assign _T_65336 = $signed(_T_56119) + $signed(_T_56124); // @[Modules.scala 150:103:@11382.4]
  assign _T_65337 = _T_65336[4:0]; // @[Modules.scala 150:103:@11383.4]
  assign _T_65338 = $signed(_T_65337); // @[Modules.scala 150:103:@11384.4]
  assign _T_65340 = $signed(-4'sh1) * $signed(io_in_708); // @[Modules.scala 150:74:@11386.4]
  assign _T_65342 = $signed(-4'sh1) * $signed(io_in_709); // @[Modules.scala 151:80:@11387.4]
  assign _T_65343 = $signed(_T_65340) + $signed(_T_65342); // @[Modules.scala 150:103:@11388.4]
  assign _T_65344 = _T_65343[4:0]; // @[Modules.scala 150:103:@11389.4]
  assign _T_65345 = $signed(_T_65344); // @[Modules.scala 150:103:@11390.4]
  assign _T_65347 = $signed(-4'sh1) * $signed(io_in_710); // @[Modules.scala 150:74:@11392.4]
  assign _T_65350 = $signed(_T_65347) + $signed(_T_62231); // @[Modules.scala 150:103:@11394.4]
  assign _T_65351 = _T_65350[4:0]; // @[Modules.scala 150:103:@11395.4]
  assign _T_65352 = $signed(_T_65351); // @[Modules.scala 150:103:@11396.4]
  assign _T_65354 = $signed(-4'sh1) * $signed(io_in_712); // @[Modules.scala 150:74:@11398.4]
  assign _T_65357 = $signed(_T_65354) + $signed(_T_56145); // @[Modules.scala 150:103:@11400.4]
  assign _T_65358 = _T_65357[4:0]; // @[Modules.scala 150:103:@11401.4]
  assign _T_65359 = $signed(_T_65358); // @[Modules.scala 150:103:@11402.4]
  assign _GEN_277 = {{1{_T_56159[4]}},_T_56159}; // @[Modules.scala 150:103:@11412.4]
  assign _T_65371 = $signed(_GEN_277) + $signed(_T_59173); // @[Modules.scala 150:103:@11412.4]
  assign _T_65372 = _T_65371[5:0]; // @[Modules.scala 150:103:@11413.4]
  assign _T_65373 = $signed(_T_65372); // @[Modules.scala 150:103:@11414.4]
  assign _T_65382 = $signed(4'sh1) * $signed(io_in_722); // @[Modules.scala 150:74:@11422.4]
  assign _T_65384 = $signed(4'sh1) * $signed(io_in_723); // @[Modules.scala 151:80:@11423.4]
  assign _T_65385 = $signed(_T_65382) + $signed(_T_65384); // @[Modules.scala 150:103:@11424.4]
  assign _T_65386 = _T_65385[5:0]; // @[Modules.scala 150:103:@11425.4]
  assign _T_65387 = $signed(_T_65386); // @[Modules.scala 150:103:@11426.4]
  assign _T_65392 = $signed(_T_56182) + $signed(_T_56187); // @[Modules.scala 150:103:@11430.4]
  assign _T_65393 = _T_65392[4:0]; // @[Modules.scala 150:103:@11431.4]
  assign _T_65394 = $signed(_T_65393); // @[Modules.scala 150:103:@11432.4]
  assign _T_65399 = $signed(_T_62273) + $signed(_T_62278); // @[Modules.scala 150:103:@11436.4]
  assign _T_65400 = _T_65399[5:0]; // @[Modules.scala 150:103:@11437.4]
  assign _T_65401 = $signed(_T_65400); // @[Modules.scala 150:103:@11438.4]
  assign _T_65406 = $signed(_T_62280) + $signed(_T_62285); // @[Modules.scala 150:103:@11442.4]
  assign _T_65407 = _T_65406[5:0]; // @[Modules.scala 150:103:@11443.4]
  assign _T_65408 = $signed(_T_65407); // @[Modules.scala 150:103:@11444.4]
  assign _T_65410 = $signed(-4'sh1) * $signed(io_in_735); // @[Modules.scala 150:74:@11446.4]
  assign _T_65413 = $signed(_T_65410) + $signed(_T_62294); // @[Modules.scala 150:103:@11448.4]
  assign _T_65414 = _T_65413[4:0]; // @[Modules.scala 150:103:@11449.4]
  assign _T_65415 = $signed(_T_65414); // @[Modules.scala 150:103:@11450.4]
  assign _T_65455 = $signed(_T_56229) + $signed(_T_56236); // @[Modules.scala 150:103:@11484.4]
  assign _T_65456 = _T_65455[4:0]; // @[Modules.scala 150:103:@11485.4]
  assign _T_65457 = $signed(_T_65456); // @[Modules.scala 150:103:@11486.4]
  assign _GEN_278 = {{1{_T_62350[4]}},_T_62350}; // @[Modules.scala 150:103:@11496.4]
  assign _T_65469 = $signed(_T_56245) + $signed(_GEN_278); // @[Modules.scala 150:103:@11496.4]
  assign _T_65470 = _T_65469[5:0]; // @[Modules.scala 150:103:@11497.4]
  assign _T_65471 = $signed(_T_65470); // @[Modules.scala 150:103:@11498.4]
  assign _T_65475 = $signed(-4'sh1) * $signed(io_in_761); // @[Modules.scala 151:80:@11501.4]
  assign _T_65476 = $signed(_T_59269) + $signed(_T_65475); // @[Modules.scala 150:103:@11502.4]
  assign _T_65477 = _T_65476[4:0]; // @[Modules.scala 150:103:@11503.4]
  assign _T_65478 = $signed(_T_65477); // @[Modules.scala 150:103:@11504.4]
  assign _T_65525 = $signed(_T_62404) + $signed(_T_56292); // @[Modules.scala 150:103:@11544.4]
  assign _T_65526 = _T_65525[4:0]; // @[Modules.scala 150:103:@11545.4]
  assign _T_65527 = $signed(_T_65526); // @[Modules.scala 150:103:@11546.4]
  assign _T_65529 = $signed(-4'sh1) * $signed(io_in_777); // @[Modules.scala 150:74:@11548.4]
  assign _T_65532 = $signed(_T_65529) + $signed(_T_59327); // @[Modules.scala 150:103:@11550.4]
  assign _T_65533 = _T_65532[4:0]; // @[Modules.scala 150:103:@11551.4]
  assign _T_65534 = $signed(_T_65533); // @[Modules.scala 150:103:@11552.4]
  assign buffer_3_2 = {{8{_T_63364[5]}},_T_63364}; // @[Modules.scala 112:22:@8.4]
  assign _T_65540 = $signed(buffer_3_2) + $signed(buffer_2_3); // @[Modules.scala 160:64:@11560.4]
  assign _T_65541 = _T_65540[13:0]; // @[Modules.scala 160:64:@11561.4]
  assign buffer_3_315 = $signed(_T_65541); // @[Modules.scala 160:64:@11562.4]
  assign buffer_3_4 = {{9{_T_63378[4]}},_T_63378}; // @[Modules.scala 112:22:@8.4]
  assign _T_65543 = $signed(buffer_3_4) + $signed(buffer_2_6); // @[Modules.scala 160:64:@11564.4]
  assign _T_65544 = _T_65543[13:0]; // @[Modules.scala 160:64:@11565.4]
  assign buffer_3_316 = $signed(_T_65544); // @[Modules.scala 160:64:@11566.4]
  assign buffer_3_6 = {{8{_T_63392[5]}},_T_63392}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_7 = {{9{_T_63399[4]}},_T_63399}; // @[Modules.scala 112:22:@8.4]
  assign _T_65546 = $signed(buffer_3_6) + $signed(buffer_3_7); // @[Modules.scala 160:64:@11568.4]
  assign _T_65547 = _T_65546[13:0]; // @[Modules.scala 160:64:@11569.4]
  assign buffer_3_317 = $signed(_T_65547); // @[Modules.scala 160:64:@11570.4]
  assign buffer_3_8 = {{9{_T_63406[4]}},_T_63406}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_9 = {{9{_T_63413[4]}},_T_63413}; // @[Modules.scala 112:22:@8.4]
  assign _T_65549 = $signed(buffer_3_8) + $signed(buffer_3_9); // @[Modules.scala 160:64:@11572.4]
  assign _T_65550 = _T_65549[13:0]; // @[Modules.scala 160:64:@11573.4]
  assign buffer_3_318 = $signed(_T_65550); // @[Modules.scala 160:64:@11574.4]
  assign buffer_3_10 = {{8{_T_63420[5]}},_T_63420}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_11 = {{9{_T_63427[4]}},_T_63427}; // @[Modules.scala 112:22:@8.4]
  assign _T_65552 = $signed(buffer_3_10) + $signed(buffer_3_11); // @[Modules.scala 160:64:@11576.4]
  assign _T_65553 = _T_65552[13:0]; // @[Modules.scala 160:64:@11577.4]
  assign buffer_3_319 = $signed(_T_65553); // @[Modules.scala 160:64:@11578.4]
  assign buffer_3_12 = {{8{_T_63434[5]}},_T_63434}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_13 = {{8{_T_63441[5]}},_T_63441}; // @[Modules.scala 112:22:@8.4]
  assign _T_65555 = $signed(buffer_3_12) + $signed(buffer_3_13); // @[Modules.scala 160:64:@11580.4]
  assign _T_65556 = _T_65555[13:0]; // @[Modules.scala 160:64:@11581.4]
  assign buffer_3_320 = $signed(_T_65556); // @[Modules.scala 160:64:@11582.4]
  assign buffer_3_17 = {{9{_T_63469[4]}},_T_63469}; // @[Modules.scala 112:22:@8.4]
  assign _T_65561 = $signed(buffer_2_16) + $signed(buffer_3_17); // @[Modules.scala 160:64:@11588.4]
  assign _T_65562 = _T_65561[13:0]; // @[Modules.scala 160:64:@11589.4]
  assign buffer_3_322 = $signed(_T_65562); // @[Modules.scala 160:64:@11590.4]
  assign buffer_3_18 = {{8{_T_63476[5]}},_T_63476}; // @[Modules.scala 112:22:@8.4]
  assign _T_65564 = $signed(buffer_3_18) + $signed(buffer_0_20); // @[Modules.scala 160:64:@11592.4]
  assign _T_65565 = _T_65564[13:0]; // @[Modules.scala 160:64:@11593.4]
  assign buffer_3_323 = $signed(_T_65565); // @[Modules.scala 160:64:@11594.4]
  assign buffer_3_20 = {{9{_T_63490[4]}},_T_63490}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_21 = {{9{_T_63497[4]}},_T_63497}; // @[Modules.scala 112:22:@8.4]
  assign _T_65567 = $signed(buffer_3_20) + $signed(buffer_3_21); // @[Modules.scala 160:64:@11596.4]
  assign _T_65568 = _T_65567[13:0]; // @[Modules.scala 160:64:@11597.4]
  assign buffer_3_324 = $signed(_T_65568); // @[Modules.scala 160:64:@11598.4]
  assign buffer_3_22 = {{9{_T_63504[4]}},_T_63504}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_23 = {{9{_T_63511[4]}},_T_63511}; // @[Modules.scala 112:22:@8.4]
  assign _T_65570 = $signed(buffer_3_22) + $signed(buffer_3_23); // @[Modules.scala 160:64:@11600.4]
  assign _T_65571 = _T_65570[13:0]; // @[Modules.scala 160:64:@11601.4]
  assign buffer_3_325 = $signed(_T_65571); // @[Modules.scala 160:64:@11602.4]
  assign buffer_3_24 = {{9{_T_63518[4]}},_T_63518}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_25 = {{9{_T_63525[4]}},_T_63525}; // @[Modules.scala 112:22:@8.4]
  assign _T_65573 = $signed(buffer_3_24) + $signed(buffer_3_25); // @[Modules.scala 160:64:@11604.4]
  assign _T_65574 = _T_65573[13:0]; // @[Modules.scala 160:64:@11605.4]
  assign buffer_3_326 = $signed(_T_65574); // @[Modules.scala 160:64:@11606.4]
  assign buffer_3_26 = {{9{_T_63532[4]}},_T_63532}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_27 = {{9{_T_63539[4]}},_T_63539}; // @[Modules.scala 112:22:@8.4]
  assign _T_65576 = $signed(buffer_3_26) + $signed(buffer_3_27); // @[Modules.scala 160:64:@11608.4]
  assign _T_65577 = _T_65576[13:0]; // @[Modules.scala 160:64:@11609.4]
  assign buffer_3_327 = $signed(_T_65577); // @[Modules.scala 160:64:@11610.4]
  assign buffer_3_28 = {{9{_T_63546[4]}},_T_63546}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_29 = {{9{_T_63553[4]}},_T_63553}; // @[Modules.scala 112:22:@8.4]
  assign _T_65579 = $signed(buffer_3_28) + $signed(buffer_3_29); // @[Modules.scala 160:64:@11612.4]
  assign _T_65580 = _T_65579[13:0]; // @[Modules.scala 160:64:@11613.4]
  assign buffer_3_328 = $signed(_T_65580); // @[Modules.scala 160:64:@11614.4]
  assign buffer_3_30 = {{9{_T_63560[4]}},_T_63560}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_31 = {{8{_T_63567[5]}},_T_63567}; // @[Modules.scala 112:22:@8.4]
  assign _T_65582 = $signed(buffer_3_30) + $signed(buffer_3_31); // @[Modules.scala 160:64:@11616.4]
  assign _T_65583 = _T_65582[13:0]; // @[Modules.scala 160:64:@11617.4]
  assign buffer_3_329 = $signed(_T_65583); // @[Modules.scala 160:64:@11618.4]
  assign buffer_3_32 = {{9{_T_63574[4]}},_T_63574}; // @[Modules.scala 112:22:@8.4]
  assign _T_65585 = $signed(buffer_3_32) + $signed(buffer_1_33); // @[Modules.scala 160:64:@11620.4]
  assign _T_65586 = _T_65585[13:0]; // @[Modules.scala 160:64:@11621.4]
  assign buffer_3_330 = $signed(_T_65586); // @[Modules.scala 160:64:@11622.4]
  assign buffer_3_34 = {{9{_T_63588[4]}},_T_63588}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_35 = {{9{_T_63595[4]}},_T_63595}; // @[Modules.scala 112:22:@8.4]
  assign _T_65588 = $signed(buffer_3_34) + $signed(buffer_3_35); // @[Modules.scala 160:64:@11624.4]
  assign _T_65589 = _T_65588[13:0]; // @[Modules.scala 160:64:@11625.4]
  assign buffer_3_331 = $signed(_T_65589); // @[Modules.scala 160:64:@11626.4]
  assign buffer_3_36 = {{9{_T_63602[4]}},_T_63602}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_37 = {{9{_T_63609[4]}},_T_63609}; // @[Modules.scala 112:22:@8.4]
  assign _T_65591 = $signed(buffer_3_36) + $signed(buffer_3_37); // @[Modules.scala 160:64:@11628.4]
  assign _T_65592 = _T_65591[13:0]; // @[Modules.scala 160:64:@11629.4]
  assign buffer_3_332 = $signed(_T_65592); // @[Modules.scala 160:64:@11630.4]
  assign buffer_3_38 = {{9{_T_63616[4]}},_T_63616}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_39 = {{9{_T_63623[4]}},_T_63623}; // @[Modules.scala 112:22:@8.4]
  assign _T_65594 = $signed(buffer_3_38) + $signed(buffer_3_39); // @[Modules.scala 160:64:@11632.4]
  assign _T_65595 = _T_65594[13:0]; // @[Modules.scala 160:64:@11633.4]
  assign buffer_3_333 = $signed(_T_65595); // @[Modules.scala 160:64:@11634.4]
  assign buffer_3_40 = {{8{_T_63630[5]}},_T_63630}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_41 = {{8{_T_63637[5]}},_T_63637}; // @[Modules.scala 112:22:@8.4]
  assign _T_65597 = $signed(buffer_3_40) + $signed(buffer_3_41); // @[Modules.scala 160:64:@11636.4]
  assign _T_65598 = _T_65597[13:0]; // @[Modules.scala 160:64:@11637.4]
  assign buffer_3_334 = $signed(_T_65598); // @[Modules.scala 160:64:@11638.4]
  assign buffer_3_43 = {{8{_T_63651[5]}},_T_63651}; // @[Modules.scala 112:22:@8.4]
  assign _T_65600 = $signed(buffer_0_43) + $signed(buffer_3_43); // @[Modules.scala 160:64:@11640.4]
  assign _T_65601 = _T_65600[13:0]; // @[Modules.scala 160:64:@11641.4]
  assign buffer_3_335 = $signed(_T_65601); // @[Modules.scala 160:64:@11642.4]
  assign buffer_3_44 = {{8{_T_63658[5]}},_T_63658}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_45 = {{8{_T_63665[5]}},_T_63665}; // @[Modules.scala 112:22:@8.4]
  assign _T_65603 = $signed(buffer_3_44) + $signed(buffer_3_45); // @[Modules.scala 160:64:@11644.4]
  assign _T_65604 = _T_65603[13:0]; // @[Modules.scala 160:64:@11645.4]
  assign buffer_3_336 = $signed(_T_65604); // @[Modules.scala 160:64:@11646.4]
  assign buffer_3_46 = {{9{_T_63672[4]}},_T_63672}; // @[Modules.scala 112:22:@8.4]
  assign _T_65606 = $signed(buffer_3_46) + $signed(buffer_2_45); // @[Modules.scala 160:64:@11648.4]
  assign _T_65607 = _T_65606[13:0]; // @[Modules.scala 160:64:@11649.4]
  assign buffer_3_337 = $signed(_T_65607); // @[Modules.scala 160:64:@11650.4]
  assign buffer_3_48 = {{9{_T_63686[4]}},_T_63686}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_49 = {{9{_T_63693[4]}},_T_63693}; // @[Modules.scala 112:22:@8.4]
  assign _T_65609 = $signed(buffer_3_48) + $signed(buffer_3_49); // @[Modules.scala 160:64:@11652.4]
  assign _T_65610 = _T_65609[13:0]; // @[Modules.scala 160:64:@11653.4]
  assign buffer_3_338 = $signed(_T_65610); // @[Modules.scala 160:64:@11654.4]
  assign buffer_3_50 = {{9{_T_63700[4]}},_T_63700}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_51 = {{8{_T_63707[5]}},_T_63707}; // @[Modules.scala 112:22:@8.4]
  assign _T_65612 = $signed(buffer_3_50) + $signed(buffer_3_51); // @[Modules.scala 160:64:@11656.4]
  assign _T_65613 = _T_65612[13:0]; // @[Modules.scala 160:64:@11657.4]
  assign buffer_3_339 = $signed(_T_65613); // @[Modules.scala 160:64:@11658.4]
  assign buffer_3_52 = {{9{_T_63714[4]}},_T_63714}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_53 = {{9{_T_63721[4]}},_T_63721}; // @[Modules.scala 112:22:@8.4]
  assign _T_65615 = $signed(buffer_3_52) + $signed(buffer_3_53); // @[Modules.scala 160:64:@11660.4]
  assign _T_65616 = _T_65615[13:0]; // @[Modules.scala 160:64:@11661.4]
  assign buffer_3_340 = $signed(_T_65616); // @[Modules.scala 160:64:@11662.4]
  assign buffer_3_54 = {{8{_T_63728[5]}},_T_63728}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_55 = {{8{_T_63735[5]}},_T_63735}; // @[Modules.scala 112:22:@8.4]
  assign _T_65618 = $signed(buffer_3_54) + $signed(buffer_3_55); // @[Modules.scala 160:64:@11664.4]
  assign _T_65619 = _T_65618[13:0]; // @[Modules.scala 160:64:@11665.4]
  assign buffer_3_341 = $signed(_T_65619); // @[Modules.scala 160:64:@11666.4]
  assign buffer_3_56 = {{8{_T_63742[5]}},_T_63742}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_57 = {{8{_T_63749[5]}},_T_63749}; // @[Modules.scala 112:22:@8.4]
  assign _T_65621 = $signed(buffer_3_56) + $signed(buffer_3_57); // @[Modules.scala 160:64:@11668.4]
  assign _T_65622 = _T_65621[13:0]; // @[Modules.scala 160:64:@11669.4]
  assign buffer_3_342 = $signed(_T_65622); // @[Modules.scala 160:64:@11670.4]
  assign buffer_3_58 = {{8{_T_63756[5]}},_T_63756}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_59 = {{9{_T_63763[4]}},_T_63763}; // @[Modules.scala 112:22:@8.4]
  assign _T_65624 = $signed(buffer_3_58) + $signed(buffer_3_59); // @[Modules.scala 160:64:@11672.4]
  assign _T_65625 = _T_65624[13:0]; // @[Modules.scala 160:64:@11673.4]
  assign buffer_3_343 = $signed(_T_65625); // @[Modules.scala 160:64:@11674.4]
  assign buffer_3_60 = {{9{_T_63770[4]}},_T_63770}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_61 = {{9{_T_63777[4]}},_T_63777}; // @[Modules.scala 112:22:@8.4]
  assign _T_65627 = $signed(buffer_3_60) + $signed(buffer_3_61); // @[Modules.scala 160:64:@11676.4]
  assign _T_65628 = _T_65627[13:0]; // @[Modules.scala 160:64:@11677.4]
  assign buffer_3_344 = $signed(_T_65628); // @[Modules.scala 160:64:@11678.4]
  assign buffer_3_62 = {{9{_T_63784[4]}},_T_63784}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_63 = {{8{_T_63791[5]}},_T_63791}; // @[Modules.scala 112:22:@8.4]
  assign _T_65630 = $signed(buffer_3_62) + $signed(buffer_3_63); // @[Modules.scala 160:64:@11680.4]
  assign _T_65631 = _T_65630[13:0]; // @[Modules.scala 160:64:@11681.4]
  assign buffer_3_345 = $signed(_T_65631); // @[Modules.scala 160:64:@11682.4]
  assign buffer_3_64 = {{9{_T_63798[4]}},_T_63798}; // @[Modules.scala 112:22:@8.4]
  assign _T_65633 = $signed(buffer_3_64) + $signed(buffer_0_60); // @[Modules.scala 160:64:@11684.4]
  assign _T_65634 = _T_65633[13:0]; // @[Modules.scala 160:64:@11685.4]
  assign buffer_3_346 = $signed(_T_65634); // @[Modules.scala 160:64:@11686.4]
  assign buffer_3_66 = {{9{_T_63812[4]}},_T_63812}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_67 = {{8{_T_63819[5]}},_T_63819}; // @[Modules.scala 112:22:@8.4]
  assign _T_65636 = $signed(buffer_3_66) + $signed(buffer_3_67); // @[Modules.scala 160:64:@11688.4]
  assign _T_65637 = _T_65636[13:0]; // @[Modules.scala 160:64:@11689.4]
  assign buffer_3_347 = $signed(_T_65637); // @[Modules.scala 160:64:@11690.4]
  assign buffer_3_68 = {{8{_T_63826[5]}},_T_63826}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_69 = {{8{_T_63833[5]}},_T_63833}; // @[Modules.scala 112:22:@8.4]
  assign _T_65639 = $signed(buffer_3_68) + $signed(buffer_3_69); // @[Modules.scala 160:64:@11692.4]
  assign _T_65640 = _T_65639[13:0]; // @[Modules.scala 160:64:@11693.4]
  assign buffer_3_348 = $signed(_T_65640); // @[Modules.scala 160:64:@11694.4]
  assign buffer_3_70 = {{9{_T_63840[4]}},_T_63840}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_71 = {{9{_T_63847[4]}},_T_63847}; // @[Modules.scala 112:22:@8.4]
  assign _T_65642 = $signed(buffer_3_70) + $signed(buffer_3_71); // @[Modules.scala 160:64:@11696.4]
  assign _T_65643 = _T_65642[13:0]; // @[Modules.scala 160:64:@11697.4]
  assign buffer_3_349 = $signed(_T_65643); // @[Modules.scala 160:64:@11698.4]
  assign buffer_3_72 = {{9{_T_63854[4]}},_T_63854}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_73 = {{9{_T_63861[4]}},_T_63861}; // @[Modules.scala 112:22:@8.4]
  assign _T_65645 = $signed(buffer_3_72) + $signed(buffer_3_73); // @[Modules.scala 160:64:@11700.4]
  assign _T_65646 = _T_65645[13:0]; // @[Modules.scala 160:64:@11701.4]
  assign buffer_3_350 = $signed(_T_65646); // @[Modules.scala 160:64:@11702.4]
  assign buffer_3_74 = {{9{_T_63868[4]}},_T_63868}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_75 = {{8{_T_63875[5]}},_T_63875}; // @[Modules.scala 112:22:@8.4]
  assign _T_65648 = $signed(buffer_3_74) + $signed(buffer_3_75); // @[Modules.scala 160:64:@11704.4]
  assign _T_65649 = _T_65648[13:0]; // @[Modules.scala 160:64:@11705.4]
  assign buffer_3_351 = $signed(_T_65649); // @[Modules.scala 160:64:@11706.4]
  assign buffer_3_76 = {{8{_T_63882[5]}},_T_63882}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_77 = {{8{_T_63889[5]}},_T_63889}; // @[Modules.scala 112:22:@8.4]
  assign _T_65651 = $signed(buffer_3_76) + $signed(buffer_3_77); // @[Modules.scala 160:64:@11708.4]
  assign _T_65652 = _T_65651[13:0]; // @[Modules.scala 160:64:@11709.4]
  assign buffer_3_352 = $signed(_T_65652); // @[Modules.scala 160:64:@11710.4]
  assign buffer_3_78 = {{8{_T_63896[5]}},_T_63896}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_79 = {{8{_T_63903[5]}},_T_63903}; // @[Modules.scala 112:22:@8.4]
  assign _T_65654 = $signed(buffer_3_78) + $signed(buffer_3_79); // @[Modules.scala 160:64:@11712.4]
  assign _T_65655 = _T_65654[13:0]; // @[Modules.scala 160:64:@11713.4]
  assign buffer_3_353 = $signed(_T_65655); // @[Modules.scala 160:64:@11714.4]
  assign buffer_3_80 = {{8{_T_63910[5]}},_T_63910}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_81 = {{9{_T_63917[4]}},_T_63917}; // @[Modules.scala 112:22:@8.4]
  assign _T_65657 = $signed(buffer_3_80) + $signed(buffer_3_81); // @[Modules.scala 160:64:@11716.4]
  assign _T_65658 = _T_65657[13:0]; // @[Modules.scala 160:64:@11717.4]
  assign buffer_3_354 = $signed(_T_65658); // @[Modules.scala 160:64:@11718.4]
  assign buffer_3_85 = {{9{_T_63945[4]}},_T_63945}; // @[Modules.scala 112:22:@8.4]
  assign _T_65663 = $signed(buffer_2_82) + $signed(buffer_3_85); // @[Modules.scala 160:64:@11724.4]
  assign _T_65664 = _T_65663[13:0]; // @[Modules.scala 160:64:@11725.4]
  assign buffer_3_356 = $signed(_T_65664); // @[Modules.scala 160:64:@11726.4]
  assign buffer_3_86 = {{9{_T_63952[4]}},_T_63952}; // @[Modules.scala 112:22:@8.4]
  assign _T_65666 = $signed(buffer_3_86) + $signed(buffer_2_86); // @[Modules.scala 160:64:@11728.4]
  assign _T_65667 = _T_65666[13:0]; // @[Modules.scala 160:64:@11729.4]
  assign buffer_3_357 = $signed(_T_65667); // @[Modules.scala 160:64:@11730.4]
  assign buffer_3_89 = {{8{_T_63973[5]}},_T_63973}; // @[Modules.scala 112:22:@8.4]
  assign _T_65669 = $signed(buffer_1_86) + $signed(buffer_3_89); // @[Modules.scala 160:64:@11732.4]
  assign _T_65670 = _T_65669[13:0]; // @[Modules.scala 160:64:@11733.4]
  assign buffer_3_358 = $signed(_T_65670); // @[Modules.scala 160:64:@11734.4]
  assign buffer_3_90 = {{8{_T_63980[5]}},_T_63980}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_91 = {{8{_T_63987[5]}},_T_63987}; // @[Modules.scala 112:22:@8.4]
  assign _T_65672 = $signed(buffer_3_90) + $signed(buffer_3_91); // @[Modules.scala 160:64:@11736.4]
  assign _T_65673 = _T_65672[13:0]; // @[Modules.scala 160:64:@11737.4]
  assign buffer_3_359 = $signed(_T_65673); // @[Modules.scala 160:64:@11738.4]
  assign buffer_3_92 = {{8{_T_63994[5]}},_T_63994}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_93 = {{9{_T_64001[4]}},_T_64001}; // @[Modules.scala 112:22:@8.4]
  assign _T_65675 = $signed(buffer_3_92) + $signed(buffer_3_93); // @[Modules.scala 160:64:@11740.4]
  assign _T_65676 = _T_65675[13:0]; // @[Modules.scala 160:64:@11741.4]
  assign buffer_3_360 = $signed(_T_65676); // @[Modules.scala 160:64:@11742.4]
  assign buffer_3_94 = {{9{_T_64008[4]}},_T_64008}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_95 = {{9{_T_64015[4]}},_T_64015}; // @[Modules.scala 112:22:@8.4]
  assign _T_65678 = $signed(buffer_3_94) + $signed(buffer_3_95); // @[Modules.scala 160:64:@11744.4]
  assign _T_65679 = _T_65678[13:0]; // @[Modules.scala 160:64:@11745.4]
  assign buffer_3_361 = $signed(_T_65679); // @[Modules.scala 160:64:@11746.4]
  assign buffer_3_96 = {{8{_T_64022[5]}},_T_64022}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_97 = {{8{_T_64029[5]}},_T_64029}; // @[Modules.scala 112:22:@8.4]
  assign _T_65681 = $signed(buffer_3_96) + $signed(buffer_3_97); // @[Modules.scala 160:64:@11748.4]
  assign _T_65682 = _T_65681[13:0]; // @[Modules.scala 160:64:@11749.4]
  assign buffer_3_362 = $signed(_T_65682); // @[Modules.scala 160:64:@11750.4]
  assign buffer_3_98 = {{9{_T_64036[4]}},_T_64036}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_99 = {{9{_T_64043[4]}},_T_64043}; // @[Modules.scala 112:22:@8.4]
  assign _T_65684 = $signed(buffer_3_98) + $signed(buffer_3_99); // @[Modules.scala 160:64:@11752.4]
  assign _T_65685 = _T_65684[13:0]; // @[Modules.scala 160:64:@11753.4]
  assign buffer_3_363 = $signed(_T_65685); // @[Modules.scala 160:64:@11754.4]
  assign buffer_3_102 = {{8{_T_64064[5]}},_T_64064}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_103 = {{8{_T_64071[5]}},_T_64071}; // @[Modules.scala 112:22:@8.4]
  assign _T_65690 = $signed(buffer_3_102) + $signed(buffer_3_103); // @[Modules.scala 160:64:@11760.4]
  assign _T_65691 = _T_65690[13:0]; // @[Modules.scala 160:64:@11761.4]
  assign buffer_3_365 = $signed(_T_65691); // @[Modules.scala 160:64:@11762.4]
  assign buffer_3_104 = {{8{_T_64078[5]}},_T_64078}; // @[Modules.scala 112:22:@8.4]
  assign _T_65693 = $signed(buffer_3_104) + $signed(buffer_0_99); // @[Modules.scala 160:64:@11764.4]
  assign _T_65694 = _T_65693[13:0]; // @[Modules.scala 160:64:@11765.4]
  assign buffer_3_366 = $signed(_T_65694); // @[Modules.scala 160:64:@11766.4]
  assign buffer_3_106 = {{8{_T_64092[5]}},_T_64092}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_107 = {{9{_T_64099[4]}},_T_64099}; // @[Modules.scala 112:22:@8.4]
  assign _T_65696 = $signed(buffer_3_106) + $signed(buffer_3_107); // @[Modules.scala 160:64:@11768.4]
  assign _T_65697 = _T_65696[13:0]; // @[Modules.scala 160:64:@11769.4]
  assign buffer_3_367 = $signed(_T_65697); // @[Modules.scala 160:64:@11770.4]
  assign buffer_3_108 = {{8{_T_64106[5]}},_T_64106}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_109 = {{8{_T_64113[5]}},_T_64113}; // @[Modules.scala 112:22:@8.4]
  assign _T_65699 = $signed(buffer_3_108) + $signed(buffer_3_109); // @[Modules.scala 160:64:@11772.4]
  assign _T_65700 = _T_65699[13:0]; // @[Modules.scala 160:64:@11773.4]
  assign buffer_3_368 = $signed(_T_65700); // @[Modules.scala 160:64:@11774.4]
  assign buffer_3_110 = {{8{_T_64120[5]}},_T_64120}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_111 = {{8{_T_64127[5]}},_T_64127}; // @[Modules.scala 112:22:@8.4]
  assign _T_65702 = $signed(buffer_3_110) + $signed(buffer_3_111); // @[Modules.scala 160:64:@11776.4]
  assign _T_65703 = _T_65702[13:0]; // @[Modules.scala 160:64:@11777.4]
  assign buffer_3_369 = $signed(_T_65703); // @[Modules.scala 160:64:@11778.4]
  assign buffer_3_112 = {{9{_T_64134[4]}},_T_64134}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_113 = {{9{_T_64141[4]}},_T_64141}; // @[Modules.scala 112:22:@8.4]
  assign _T_65705 = $signed(buffer_3_112) + $signed(buffer_3_113); // @[Modules.scala 160:64:@11780.4]
  assign _T_65706 = _T_65705[13:0]; // @[Modules.scala 160:64:@11781.4]
  assign buffer_3_370 = $signed(_T_65706); // @[Modules.scala 160:64:@11782.4]
  assign buffer_3_117 = {{8{_T_64169[5]}},_T_64169}; // @[Modules.scala 112:22:@8.4]
  assign _T_65711 = $signed(buffer_0_110) + $signed(buffer_3_117); // @[Modules.scala 160:64:@11788.4]
  assign _T_65712 = _T_65711[13:0]; // @[Modules.scala 160:64:@11789.4]
  assign buffer_3_372 = $signed(_T_65712); // @[Modules.scala 160:64:@11790.4]
  assign buffer_3_118 = {{8{_T_64176[5]}},_T_64176}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_119 = {{9{_T_64183[4]}},_T_64183}; // @[Modules.scala 112:22:@8.4]
  assign _T_65714 = $signed(buffer_3_118) + $signed(buffer_3_119); // @[Modules.scala 160:64:@11792.4]
  assign _T_65715 = _T_65714[13:0]; // @[Modules.scala 160:64:@11793.4]
  assign buffer_3_373 = $signed(_T_65715); // @[Modules.scala 160:64:@11794.4]
  assign buffer_3_121 = {{8{_T_64197[5]}},_T_64197}; // @[Modules.scala 112:22:@8.4]
  assign _T_65717 = $signed(buffer_2_117) + $signed(buffer_3_121); // @[Modules.scala 160:64:@11796.4]
  assign _T_65718 = _T_65717[13:0]; // @[Modules.scala 160:64:@11797.4]
  assign buffer_3_374 = $signed(_T_65718); // @[Modules.scala 160:64:@11798.4]
  assign buffer_3_122 = {{8{_T_64204[5]}},_T_64204}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_123 = {{8{_T_64211[5]}},_T_64211}; // @[Modules.scala 112:22:@8.4]
  assign _T_65720 = $signed(buffer_3_122) + $signed(buffer_3_123); // @[Modules.scala 160:64:@11800.4]
  assign _T_65721 = _T_65720[13:0]; // @[Modules.scala 160:64:@11801.4]
  assign buffer_3_375 = $signed(_T_65721); // @[Modules.scala 160:64:@11802.4]
  assign buffer_3_124 = {{8{_T_64218[5]}},_T_64218}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_125 = {{8{_T_64225[5]}},_T_64225}; // @[Modules.scala 112:22:@8.4]
  assign _T_65723 = $signed(buffer_3_124) + $signed(buffer_3_125); // @[Modules.scala 160:64:@11804.4]
  assign _T_65724 = _T_65723[13:0]; // @[Modules.scala 160:64:@11805.4]
  assign buffer_3_376 = $signed(_T_65724); // @[Modules.scala 160:64:@11806.4]
  assign buffer_3_126 = {{8{_T_64232[5]}},_T_64232}; // @[Modules.scala 112:22:@8.4]
  assign _T_65726 = $signed(buffer_3_126) + $signed(buffer_0_120); // @[Modules.scala 160:64:@11808.4]
  assign _T_65727 = _T_65726[13:0]; // @[Modules.scala 160:64:@11809.4]
  assign buffer_3_377 = $signed(_T_65727); // @[Modules.scala 160:64:@11810.4]
  assign _T_65729 = $signed(buffer_0_121) + $signed(buffer_0_122); // @[Modules.scala 160:64:@11812.4]
  assign _T_65730 = _T_65729[13:0]; // @[Modules.scala 160:64:@11813.4]
  assign buffer_3_378 = $signed(_T_65730); // @[Modules.scala 160:64:@11814.4]
  assign buffer_3_131 = {{8{_T_64267[5]}},_T_64267}; // @[Modules.scala 112:22:@8.4]
  assign _T_65732 = $signed(buffer_0_123) + $signed(buffer_3_131); // @[Modules.scala 160:64:@11816.4]
  assign _T_65733 = _T_65732[13:0]; // @[Modules.scala 160:64:@11817.4]
  assign buffer_3_379 = $signed(_T_65733); // @[Modules.scala 160:64:@11818.4]
  assign buffer_3_132 = {{8{_T_64274[5]}},_T_64274}; // @[Modules.scala 112:22:@8.4]
  assign _T_65735 = $signed(buffer_3_132) + $signed(buffer_1_128); // @[Modules.scala 160:64:@11820.4]
  assign _T_65736 = _T_65735[13:0]; // @[Modules.scala 160:64:@11821.4]
  assign buffer_3_380 = $signed(_T_65736); // @[Modules.scala 160:64:@11822.4]
  assign buffer_3_134 = {{8{_T_64288[5]}},_T_64288}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_135 = {{8{_T_64295[5]}},_T_64295}; // @[Modules.scala 112:22:@8.4]
  assign _T_65738 = $signed(buffer_3_134) + $signed(buffer_3_135); // @[Modules.scala 160:64:@11824.4]
  assign _T_65739 = _T_65738[13:0]; // @[Modules.scala 160:64:@11825.4]
  assign buffer_3_381 = $signed(_T_65739); // @[Modules.scala 160:64:@11826.4]
  assign _T_65741 = $signed(buffer_2_131) + $signed(buffer_2_132); // @[Modules.scala 160:64:@11828.4]
  assign _T_65742 = _T_65741[13:0]; // @[Modules.scala 160:64:@11829.4]
  assign buffer_3_382 = $signed(_T_65742); // @[Modules.scala 160:64:@11830.4]
  assign _T_65744 = $signed(buffer_2_133) + $signed(buffer_1_133); // @[Modules.scala 160:64:@11832.4]
  assign _T_65745 = _T_65744[13:0]; // @[Modules.scala 160:64:@11833.4]
  assign buffer_3_383 = $signed(_T_65745); // @[Modules.scala 160:64:@11834.4]
  assign buffer_3_141 = {{9{_T_64337[4]}},_T_64337}; // @[Modules.scala 112:22:@8.4]
  assign _T_65747 = $signed(buffer_1_134) + $signed(buffer_3_141); // @[Modules.scala 160:64:@11836.4]
  assign _T_65748 = _T_65747[13:0]; // @[Modules.scala 160:64:@11837.4]
  assign buffer_3_384 = $signed(_T_65748); // @[Modules.scala 160:64:@11838.4]
  assign buffer_3_142 = {{9{_T_64344[4]}},_T_64344}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_143 = {{9{_T_64351[4]}},_T_64351}; // @[Modules.scala 112:22:@8.4]
  assign _T_65750 = $signed(buffer_3_142) + $signed(buffer_3_143); // @[Modules.scala 160:64:@11840.4]
  assign _T_65751 = _T_65750[13:0]; // @[Modules.scala 160:64:@11841.4]
  assign buffer_3_385 = $signed(_T_65751); // @[Modules.scala 160:64:@11842.4]
  assign buffer_3_144 = {{8{_T_64358[5]}},_T_64358}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_145 = {{8{_T_64365[5]}},_T_64365}; // @[Modules.scala 112:22:@8.4]
  assign _T_65753 = $signed(buffer_3_144) + $signed(buffer_3_145); // @[Modules.scala 160:64:@11844.4]
  assign _T_65754 = _T_65753[13:0]; // @[Modules.scala 160:64:@11845.4]
  assign buffer_3_386 = $signed(_T_65754); // @[Modules.scala 160:64:@11846.4]
  assign buffer_3_147 = {{8{_T_64379[5]}},_T_64379}; // @[Modules.scala 112:22:@8.4]
  assign _T_65756 = $signed(buffer_2_142) + $signed(buffer_3_147); // @[Modules.scala 160:64:@11848.4]
  assign _T_65757 = _T_65756[13:0]; // @[Modules.scala 160:64:@11849.4]
  assign buffer_3_387 = $signed(_T_65757); // @[Modules.scala 160:64:@11850.4]
  assign buffer_3_152 = {{8{_T_64414[5]}},_T_64414}; // @[Modules.scala 112:22:@8.4]
  assign _T_65765 = $signed(buffer_3_152) + $signed(buffer_2_149); // @[Modules.scala 160:64:@11860.4]
  assign _T_65766 = _T_65765[13:0]; // @[Modules.scala 160:64:@11861.4]
  assign buffer_3_390 = $signed(_T_65766); // @[Modules.scala 160:64:@11862.4]
  assign buffer_3_155 = {{8{_T_64435[5]}},_T_64435}; // @[Modules.scala 112:22:@8.4]
  assign _T_65768 = $signed(buffer_2_150) + $signed(buffer_3_155); // @[Modules.scala 160:64:@11864.4]
  assign _T_65769 = _T_65768[13:0]; // @[Modules.scala 160:64:@11865.4]
  assign buffer_3_391 = $signed(_T_65769); // @[Modules.scala 160:64:@11866.4]
  assign buffer_3_156 = {{9{_T_64442[4]}},_T_64442}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_157 = {{9{_T_64449[4]}},_T_64449}; // @[Modules.scala 112:22:@8.4]
  assign _T_65771 = $signed(buffer_3_156) + $signed(buffer_3_157); // @[Modules.scala 160:64:@11868.4]
  assign _T_65772 = _T_65771[13:0]; // @[Modules.scala 160:64:@11869.4]
  assign buffer_3_392 = $signed(_T_65772); // @[Modules.scala 160:64:@11870.4]
  assign buffer_3_158 = {{8{_T_64456[5]}},_T_64456}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_159 = {{8{_T_64463[5]}},_T_64463}; // @[Modules.scala 112:22:@8.4]
  assign _T_65774 = $signed(buffer_3_158) + $signed(buffer_3_159); // @[Modules.scala 160:64:@11872.4]
  assign _T_65775 = _T_65774[13:0]; // @[Modules.scala 160:64:@11873.4]
  assign buffer_3_393 = $signed(_T_65775); // @[Modules.scala 160:64:@11874.4]
  assign _T_65777 = $signed(buffer_2_157) + $signed(buffer_2_158); // @[Modules.scala 160:64:@11876.4]
  assign _T_65778 = _T_65777[13:0]; // @[Modules.scala 160:64:@11877.4]
  assign buffer_3_394 = $signed(_T_65778); // @[Modules.scala 160:64:@11878.4]
  assign buffer_3_163 = {{8{_T_64491[5]}},_T_64491}; // @[Modules.scala 112:22:@8.4]
  assign _T_65780 = $signed(buffer_2_159) + $signed(buffer_3_163); // @[Modules.scala 160:64:@11880.4]
  assign _T_65781 = _T_65780[13:0]; // @[Modules.scala 160:64:@11881.4]
  assign buffer_3_395 = $signed(_T_65781); // @[Modules.scala 160:64:@11882.4]
  assign buffer_3_164 = {{8{_T_64498[5]}},_T_64498}; // @[Modules.scala 112:22:@8.4]
  assign _T_65783 = $signed(buffer_3_164) + $signed(buffer_2_162); // @[Modules.scala 160:64:@11884.4]
  assign _T_65784 = _T_65783[13:0]; // @[Modules.scala 160:64:@11885.4]
  assign buffer_3_396 = $signed(_T_65784); // @[Modules.scala 160:64:@11886.4]
  assign buffer_3_166 = {{8{_T_64512[5]}},_T_64512}; // @[Modules.scala 112:22:@8.4]
  assign _T_65786 = $signed(buffer_3_166) + $signed(buffer_1_161); // @[Modules.scala 160:64:@11888.4]
  assign _T_65787 = _T_65786[13:0]; // @[Modules.scala 160:64:@11889.4]
  assign buffer_3_397 = $signed(_T_65787); // @[Modules.scala 160:64:@11890.4]
  assign buffer_3_169 = {{8{_T_64533[5]}},_T_64533}; // @[Modules.scala 112:22:@8.4]
  assign _T_65789 = $signed(buffer_1_162) + $signed(buffer_3_169); // @[Modules.scala 160:64:@11892.4]
  assign _T_65790 = _T_65789[13:0]; // @[Modules.scala 160:64:@11893.4]
  assign buffer_3_398 = $signed(_T_65790); // @[Modules.scala 160:64:@11894.4]
  assign buffer_3_171 = {{8{_T_64547[5]}},_T_64547}; // @[Modules.scala 112:22:@8.4]
  assign _T_65792 = $signed(buffer_0_163) + $signed(buffer_3_171); // @[Modules.scala 160:64:@11896.4]
  assign _T_65793 = _T_65792[13:0]; // @[Modules.scala 160:64:@11897.4]
  assign buffer_3_399 = $signed(_T_65793); // @[Modules.scala 160:64:@11898.4]
  assign buffer_3_172 = {{8{_T_64554[5]}},_T_64554}; // @[Modules.scala 112:22:@8.4]
  assign _T_65795 = $signed(buffer_3_172) + $signed(buffer_0_167); // @[Modules.scala 160:64:@11900.4]
  assign _T_65796 = _T_65795[13:0]; // @[Modules.scala 160:64:@11901.4]
  assign buffer_3_400 = $signed(_T_65796); // @[Modules.scala 160:64:@11902.4]
  assign buffer_3_175 = {{9{_T_64575[4]}},_T_64575}; // @[Modules.scala 112:22:@8.4]
  assign _T_65798 = $signed(buffer_0_168) + $signed(buffer_3_175); // @[Modules.scala 160:64:@11904.4]
  assign _T_65799 = _T_65798[13:0]; // @[Modules.scala 160:64:@11905.4]
  assign buffer_3_401 = $signed(_T_65799); // @[Modules.scala 160:64:@11906.4]
  assign buffer_3_176 = {{9{_T_64582[4]}},_T_64582}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_177 = {{9{_T_64589[4]}},_T_64589}; // @[Modules.scala 112:22:@8.4]
  assign _T_65801 = $signed(buffer_3_176) + $signed(buffer_3_177); // @[Modules.scala 160:64:@11908.4]
  assign _T_65802 = _T_65801[13:0]; // @[Modules.scala 160:64:@11909.4]
  assign buffer_3_402 = $signed(_T_65802); // @[Modules.scala 160:64:@11910.4]
  assign _T_65804 = $signed(buffer_1_171) + $signed(buffer_1_172); // @[Modules.scala 160:64:@11912.4]
  assign _T_65805 = _T_65804[13:0]; // @[Modules.scala 160:64:@11913.4]
  assign buffer_3_403 = $signed(_T_65805); // @[Modules.scala 160:64:@11914.4]
  assign buffer_3_180 = {{9{_T_64610[4]}},_T_64610}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_181 = {{9{_T_64617[4]}},_T_64617}; // @[Modules.scala 112:22:@8.4]
  assign _T_65807 = $signed(buffer_3_180) + $signed(buffer_3_181); // @[Modules.scala 160:64:@11916.4]
  assign _T_65808 = _T_65807[13:0]; // @[Modules.scala 160:64:@11917.4]
  assign buffer_3_404 = $signed(_T_65808); // @[Modules.scala 160:64:@11918.4]
  assign buffer_3_182 = {{9{_T_64624[4]}},_T_64624}; // @[Modules.scala 112:22:@8.4]
  assign _T_65810 = $signed(buffer_3_182) + $signed(buffer_1_176); // @[Modules.scala 160:64:@11920.4]
  assign _T_65811 = _T_65810[13:0]; // @[Modules.scala 160:64:@11921.4]
  assign buffer_3_405 = $signed(_T_65811); // @[Modules.scala 160:64:@11922.4]
  assign buffer_3_184 = {{8{_T_64638[5]}},_T_64638}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_185 = {{8{_T_64645[5]}},_T_64645}; // @[Modules.scala 112:22:@8.4]
  assign _T_65813 = $signed(buffer_3_184) + $signed(buffer_3_185); // @[Modules.scala 160:64:@11924.4]
  assign _T_65814 = _T_65813[13:0]; // @[Modules.scala 160:64:@11925.4]
  assign buffer_3_406 = $signed(_T_65814); // @[Modules.scala 160:64:@11926.4]
  assign buffer_3_186 = {{8{_T_64652[5]}},_T_64652}; // @[Modules.scala 112:22:@8.4]
  assign _T_65816 = $signed(buffer_3_186) + $signed(buffer_0_179); // @[Modules.scala 160:64:@11928.4]
  assign _T_65817 = _T_65816[13:0]; // @[Modules.scala 160:64:@11929.4]
  assign buffer_3_407 = $signed(_T_65817); // @[Modules.scala 160:64:@11930.4]
  assign buffer_3_189 = {{9{_T_64673[4]}},_T_64673}; // @[Modules.scala 112:22:@8.4]
  assign _T_65819 = $signed(buffer_0_180) + $signed(buffer_3_189); // @[Modules.scala 160:64:@11932.4]
  assign _T_65820 = _T_65819[13:0]; // @[Modules.scala 160:64:@11933.4]
  assign buffer_3_408 = $signed(_T_65820); // @[Modules.scala 160:64:@11934.4]
  assign buffer_3_190 = {{9{_T_64680[4]}},_T_64680}; // @[Modules.scala 112:22:@8.4]
  assign _T_65822 = $signed(buffer_3_190) + $signed(buffer_2_188); // @[Modules.scala 160:64:@11936.4]
  assign _T_65823 = _T_65822[13:0]; // @[Modules.scala 160:64:@11937.4]
  assign buffer_3_409 = $signed(_T_65823); // @[Modules.scala 160:64:@11938.4]
  assign buffer_3_193 = {{9{_T_64701[4]}},_T_64701}; // @[Modules.scala 112:22:@8.4]
  assign _T_65825 = $signed(buffer_1_183) + $signed(buffer_3_193); // @[Modules.scala 160:64:@11940.4]
  assign _T_65826 = _T_65825[13:0]; // @[Modules.scala 160:64:@11941.4]
  assign buffer_3_410 = $signed(_T_65826); // @[Modules.scala 160:64:@11942.4]
  assign buffer_3_194 = {{8{_T_64708[5]}},_T_64708}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_195 = {{9{_T_64715[4]}},_T_64715}; // @[Modules.scala 112:22:@8.4]
  assign _T_65828 = $signed(buffer_3_194) + $signed(buffer_3_195); // @[Modules.scala 160:64:@11944.4]
  assign _T_65829 = _T_65828[13:0]; // @[Modules.scala 160:64:@11945.4]
  assign buffer_3_411 = $signed(_T_65829); // @[Modules.scala 160:64:@11946.4]
  assign buffer_3_196 = {{9{_T_64722[4]}},_T_64722}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_197 = {{8{_T_64729[5]}},_T_64729}; // @[Modules.scala 112:22:@8.4]
  assign _T_65831 = $signed(buffer_3_196) + $signed(buffer_3_197); // @[Modules.scala 160:64:@11948.4]
  assign _T_65832 = _T_65831[13:0]; // @[Modules.scala 160:64:@11949.4]
  assign buffer_3_412 = $signed(_T_65832); // @[Modules.scala 160:64:@11950.4]
  assign _T_65834 = $signed(buffer_0_187) + $signed(buffer_0_188); // @[Modules.scala 160:64:@11952.4]
  assign _T_65835 = _T_65834[13:0]; // @[Modules.scala 160:64:@11953.4]
  assign buffer_3_413 = $signed(_T_65835); // @[Modules.scala 160:64:@11954.4]
  assign buffer_3_200 = {{8{_T_64750[5]}},_T_64750}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_201 = {{9{_T_64757[4]}},_T_64757}; // @[Modules.scala 112:22:@8.4]
  assign _T_65837 = $signed(buffer_3_200) + $signed(buffer_3_201); // @[Modules.scala 160:64:@11956.4]
  assign _T_65838 = _T_65837[13:0]; // @[Modules.scala 160:64:@11957.4]
  assign buffer_3_414 = $signed(_T_65838); // @[Modules.scala 160:64:@11958.4]
  assign buffer_3_203 = {{9{_T_64771[4]}},_T_64771}; // @[Modules.scala 112:22:@8.4]
  assign _T_65840 = $signed(buffer_2_198) + $signed(buffer_3_203); // @[Modules.scala 160:64:@11960.4]
  assign _T_65841 = _T_65840[13:0]; // @[Modules.scala 160:64:@11961.4]
  assign buffer_3_415 = $signed(_T_65841); // @[Modules.scala 160:64:@11962.4]
  assign buffer_3_204 = {{8{_T_64778[5]}},_T_64778}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_205 = {{8{_T_64785[5]}},_T_64785}; // @[Modules.scala 112:22:@8.4]
  assign _T_65843 = $signed(buffer_3_204) + $signed(buffer_3_205); // @[Modules.scala 160:64:@11964.4]
  assign _T_65844 = _T_65843[13:0]; // @[Modules.scala 160:64:@11965.4]
  assign buffer_3_416 = $signed(_T_65844); // @[Modules.scala 160:64:@11966.4]
  assign buffer_3_206 = {{9{_T_64792[4]}},_T_64792}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_207 = {{8{_T_64799[5]}},_T_64799}; // @[Modules.scala 112:22:@8.4]
  assign _T_65846 = $signed(buffer_3_206) + $signed(buffer_3_207); // @[Modules.scala 160:64:@11968.4]
  assign _T_65847 = _T_65846[13:0]; // @[Modules.scala 160:64:@11969.4]
  assign buffer_3_417 = $signed(_T_65847); // @[Modules.scala 160:64:@11970.4]
  assign buffer_3_208 = {{8{_T_64806[5]}},_T_64806}; // @[Modules.scala 112:22:@8.4]
  assign _T_65849 = $signed(buffer_3_208) + $signed(buffer_0_199); // @[Modules.scala 160:64:@11972.4]
  assign _T_65850 = _T_65849[13:0]; // @[Modules.scala 160:64:@11973.4]
  assign buffer_3_418 = $signed(_T_65850); // @[Modules.scala 160:64:@11974.4]
  assign buffer_3_211 = {{8{_T_64827[5]}},_T_64827}; // @[Modules.scala 112:22:@8.4]
  assign _T_65852 = $signed(buffer_0_200) + $signed(buffer_3_211); // @[Modules.scala 160:64:@11976.4]
  assign _T_65853 = _T_65852[13:0]; // @[Modules.scala 160:64:@11977.4]
  assign buffer_3_419 = $signed(_T_65853); // @[Modules.scala 160:64:@11978.4]
  assign buffer_3_212 = {{9{_T_64834[4]}},_T_64834}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_213 = {{8{_T_64841[5]}},_T_64841}; // @[Modules.scala 112:22:@8.4]
  assign _T_65855 = $signed(buffer_3_212) + $signed(buffer_3_213); // @[Modules.scala 160:64:@11980.4]
  assign _T_65856 = _T_65855[13:0]; // @[Modules.scala 160:64:@11981.4]
  assign buffer_3_420 = $signed(_T_65856); // @[Modules.scala 160:64:@11982.4]
  assign buffer_3_214 = {{9{_T_64848[4]}},_T_64848}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_215 = {{9{_T_64855[4]}},_T_64855}; // @[Modules.scala 112:22:@8.4]
  assign _T_65858 = $signed(buffer_3_214) + $signed(buffer_3_215); // @[Modules.scala 160:64:@11984.4]
  assign _T_65859 = _T_65858[13:0]; // @[Modules.scala 160:64:@11985.4]
  assign buffer_3_421 = $signed(_T_65859); // @[Modules.scala 160:64:@11986.4]
  assign buffer_3_216 = {{8{_T_64862[5]}},_T_64862}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_217 = {{8{_T_64869[5]}},_T_64869}; // @[Modules.scala 112:22:@8.4]
  assign _T_65861 = $signed(buffer_3_216) + $signed(buffer_3_217); // @[Modules.scala 160:64:@11988.4]
  assign _T_65862 = _T_65861[13:0]; // @[Modules.scala 160:64:@11989.4]
  assign buffer_3_422 = $signed(_T_65862); // @[Modules.scala 160:64:@11990.4]
  assign buffer_3_218 = {{9{_T_64876[4]}},_T_64876}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_219 = {{9{_T_64883[4]}},_T_64883}; // @[Modules.scala 112:22:@8.4]
  assign _T_65864 = $signed(buffer_3_218) + $signed(buffer_3_219); // @[Modules.scala 160:64:@11992.4]
  assign _T_65865 = _T_65864[13:0]; // @[Modules.scala 160:64:@11993.4]
  assign buffer_3_423 = $signed(_T_65865); // @[Modules.scala 160:64:@11994.4]
  assign buffer_3_220 = {{9{_T_64890[4]}},_T_64890}; // @[Modules.scala 112:22:@8.4]
  assign _T_65867 = $signed(buffer_3_220) + $signed(buffer_1_211); // @[Modules.scala 160:64:@11996.4]
  assign _T_65868 = _T_65867[13:0]; // @[Modules.scala 160:64:@11997.4]
  assign buffer_3_424 = $signed(_T_65868); // @[Modules.scala 160:64:@11998.4]
  assign buffer_3_223 = {{9{_T_64911[4]}},_T_64911}; // @[Modules.scala 112:22:@8.4]
  assign _T_65870 = $signed(buffer_1_212) + $signed(buffer_3_223); // @[Modules.scala 160:64:@12000.4]
  assign _T_65871 = _T_65870[13:0]; // @[Modules.scala 160:64:@12001.4]
  assign buffer_3_425 = $signed(_T_65871); // @[Modules.scala 160:64:@12002.4]
  assign buffer_3_225 = {{8{_T_64925[5]}},_T_64925}; // @[Modules.scala 112:22:@8.4]
  assign _T_65873 = $signed(buffer_1_214) + $signed(buffer_3_225); // @[Modules.scala 160:64:@12004.4]
  assign _T_65874 = _T_65873[13:0]; // @[Modules.scala 160:64:@12005.4]
  assign buffer_3_426 = $signed(_T_65874); // @[Modules.scala 160:64:@12006.4]
  assign buffer_3_226 = {{9{_T_64932[4]}},_T_64932}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_227 = {{8{_T_64939[5]}},_T_64939}; // @[Modules.scala 112:22:@8.4]
  assign _T_65876 = $signed(buffer_3_226) + $signed(buffer_3_227); // @[Modules.scala 160:64:@12008.4]
  assign _T_65877 = _T_65876[13:0]; // @[Modules.scala 160:64:@12009.4]
  assign buffer_3_427 = $signed(_T_65877); // @[Modules.scala 160:64:@12010.4]
  assign buffer_3_228 = {{8{_T_64946[5]}},_T_64946}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_229 = {{9{_T_64953[4]}},_T_64953}; // @[Modules.scala 112:22:@8.4]
  assign _T_65879 = $signed(buffer_3_228) + $signed(buffer_3_229); // @[Modules.scala 160:64:@12012.4]
  assign _T_65880 = _T_65879[13:0]; // @[Modules.scala 160:64:@12013.4]
  assign buffer_3_428 = $signed(_T_65880); // @[Modules.scala 160:64:@12014.4]
  assign buffer_3_232 = {{8{_T_64974[5]}},_T_64974}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_233 = {{9{_T_64981[4]}},_T_64981}; // @[Modules.scala 112:22:@8.4]
  assign _T_65885 = $signed(buffer_3_232) + $signed(buffer_3_233); // @[Modules.scala 160:64:@12020.4]
  assign _T_65886 = _T_65885[13:0]; // @[Modules.scala 160:64:@12021.4]
  assign buffer_3_430 = $signed(_T_65886); // @[Modules.scala 160:64:@12022.4]
  assign buffer_3_234 = {{9{_T_64988[4]}},_T_64988}; // @[Modules.scala 112:22:@8.4]
  assign _T_65888 = $signed(buffer_3_234) + $signed(buffer_1_224); // @[Modules.scala 160:64:@12024.4]
  assign _T_65889 = _T_65888[13:0]; // @[Modules.scala 160:64:@12025.4]
  assign buffer_3_431 = $signed(_T_65889); // @[Modules.scala 160:64:@12026.4]
  assign buffer_3_237 = {{8{_T_65009[5]}},_T_65009}; // @[Modules.scala 112:22:@8.4]
  assign _T_65891 = $signed(buffer_2_230) + $signed(buffer_3_237); // @[Modules.scala 160:64:@12028.4]
  assign _T_65892 = _T_65891[13:0]; // @[Modules.scala 160:64:@12029.4]
  assign buffer_3_432 = $signed(_T_65892); // @[Modules.scala 160:64:@12030.4]
  assign _T_65894 = $signed(buffer_2_233) + $signed(buffer_2_234); // @[Modules.scala 160:64:@12032.4]
  assign _T_65895 = _T_65894[13:0]; // @[Modules.scala 160:64:@12033.4]
  assign buffer_3_433 = $signed(_T_65895); // @[Modules.scala 160:64:@12034.4]
  assign buffer_3_240 = {{9{_T_65030[4]}},_T_65030}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_241 = {{9{_T_65037[4]}},_T_65037}; // @[Modules.scala 112:22:@8.4]
  assign _T_65897 = $signed(buffer_3_240) + $signed(buffer_3_241); // @[Modules.scala 160:64:@12036.4]
  assign _T_65898 = _T_65897[13:0]; // @[Modules.scala 160:64:@12037.4]
  assign buffer_3_434 = $signed(_T_65898); // @[Modules.scala 160:64:@12038.4]
  assign buffer_3_243 = {{8{_T_65051[5]}},_T_65051}; // @[Modules.scala 112:22:@8.4]
  assign _T_65900 = $signed(buffer_0_231) + $signed(buffer_3_243); // @[Modules.scala 160:64:@12040.4]
  assign _T_65901 = _T_65900[13:0]; // @[Modules.scala 160:64:@12041.4]
  assign buffer_3_435 = $signed(_T_65901); // @[Modules.scala 160:64:@12042.4]
  assign buffer_3_244 = {{9{_T_65058[4]}},_T_65058}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_245 = {{8{_T_65065[5]}},_T_65065}; // @[Modules.scala 112:22:@8.4]
  assign _T_65903 = $signed(buffer_3_244) + $signed(buffer_3_245); // @[Modules.scala 160:64:@12044.4]
  assign _T_65904 = _T_65903[13:0]; // @[Modules.scala 160:64:@12045.4]
  assign buffer_3_436 = $signed(_T_65904); // @[Modules.scala 160:64:@12046.4]
  assign buffer_3_247 = {{8{_T_65079[5]}},_T_65079}; // @[Modules.scala 112:22:@8.4]
  assign _T_65906 = $signed(buffer_1_238) + $signed(buffer_3_247); // @[Modules.scala 160:64:@12048.4]
  assign _T_65907 = _T_65906[13:0]; // @[Modules.scala 160:64:@12049.4]
  assign buffer_3_437 = $signed(_T_65907); // @[Modules.scala 160:64:@12050.4]
  assign buffer_3_248 = {{8{_T_65086[5]}},_T_65086}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_249 = {{9{_T_65093[4]}},_T_65093}; // @[Modules.scala 112:22:@8.4]
  assign _T_65909 = $signed(buffer_3_248) + $signed(buffer_3_249); // @[Modules.scala 160:64:@12052.4]
  assign _T_65910 = _T_65909[13:0]; // @[Modules.scala 160:64:@12053.4]
  assign buffer_3_438 = $signed(_T_65910); // @[Modules.scala 160:64:@12054.4]
  assign buffer_3_250 = {{9{_T_65100[4]}},_T_65100}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_251 = {{9{_T_65107[4]}},_T_65107}; // @[Modules.scala 112:22:@8.4]
  assign _T_65912 = $signed(buffer_3_250) + $signed(buffer_3_251); // @[Modules.scala 160:64:@12056.4]
  assign _T_65913 = _T_65912[13:0]; // @[Modules.scala 160:64:@12057.4]
  assign buffer_3_439 = $signed(_T_65913); // @[Modules.scala 160:64:@12058.4]
  assign buffer_3_252 = {{9{_T_65114[4]}},_T_65114}; // @[Modules.scala 112:22:@8.4]
  assign _T_65915 = $signed(buffer_3_252) + $signed(buffer_0_242); // @[Modules.scala 160:64:@12060.4]
  assign _T_65916 = _T_65915[13:0]; // @[Modules.scala 160:64:@12061.4]
  assign buffer_3_440 = $signed(_T_65916); // @[Modules.scala 160:64:@12062.4]
  assign buffer_3_254 = {{8{_T_65128[5]}},_T_65128}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_255 = {{8{_T_65135[5]}},_T_65135}; // @[Modules.scala 112:22:@8.4]
  assign _T_65918 = $signed(buffer_3_254) + $signed(buffer_3_255); // @[Modules.scala 160:64:@12064.4]
  assign _T_65919 = _T_65918[13:0]; // @[Modules.scala 160:64:@12065.4]
  assign buffer_3_441 = $signed(_T_65919); // @[Modules.scala 160:64:@12066.4]
  assign buffer_3_256 = {{8{_T_65142[5]}},_T_65142}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_257 = {{8{_T_65149[5]}},_T_65149}; // @[Modules.scala 112:22:@8.4]
  assign _T_65921 = $signed(buffer_3_256) + $signed(buffer_3_257); // @[Modules.scala 160:64:@12068.4]
  assign _T_65922 = _T_65921[13:0]; // @[Modules.scala 160:64:@12069.4]
  assign buffer_3_442 = $signed(_T_65922); // @[Modules.scala 160:64:@12070.4]
  assign buffer_3_258 = {{8{_T_65156[5]}},_T_65156}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_259 = {{9{_T_65163[4]}},_T_65163}; // @[Modules.scala 112:22:@8.4]
  assign _T_65924 = $signed(buffer_3_258) + $signed(buffer_3_259); // @[Modules.scala 160:64:@12072.4]
  assign _T_65925 = _T_65924[13:0]; // @[Modules.scala 160:64:@12073.4]
  assign buffer_3_443 = $signed(_T_65925); // @[Modules.scala 160:64:@12074.4]
  assign buffer_3_260 = {{9{_T_65170[4]}},_T_65170}; // @[Modules.scala 112:22:@8.4]
  assign _T_65927 = $signed(buffer_3_260) + $signed(buffer_2_258); // @[Modules.scala 160:64:@12076.4]
  assign _T_65928 = _T_65927[13:0]; // @[Modules.scala 160:64:@12077.4]
  assign buffer_3_444 = $signed(_T_65928); // @[Modules.scala 160:64:@12078.4]
  assign buffer_3_263 = {{8{_T_65191[5]}},_T_65191}; // @[Modules.scala 112:22:@8.4]
  assign _T_65930 = $signed(buffer_2_259) + $signed(buffer_3_263); // @[Modules.scala 160:64:@12080.4]
  assign _T_65931 = _T_65930[13:0]; // @[Modules.scala 160:64:@12081.4]
  assign buffer_3_445 = $signed(_T_65931); // @[Modules.scala 160:64:@12082.4]
  assign buffer_3_264 = {{8{_T_65198[5]}},_T_65198}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_265 = {{8{_T_65205[5]}},_T_65205}; // @[Modules.scala 112:22:@8.4]
  assign _T_65933 = $signed(buffer_3_264) + $signed(buffer_3_265); // @[Modules.scala 160:64:@12084.4]
  assign _T_65934 = _T_65933[13:0]; // @[Modules.scala 160:64:@12085.4]
  assign buffer_3_446 = $signed(_T_65934); // @[Modules.scala 160:64:@12086.4]
  assign _T_65936 = $signed(buffer_2_265) + $signed(buffer_2_266); // @[Modules.scala 160:64:@12088.4]
  assign _T_65937 = _T_65936[13:0]; // @[Modules.scala 160:64:@12089.4]
  assign buffer_3_447 = $signed(_T_65937); // @[Modules.scala 160:64:@12090.4]
  assign buffer_3_268 = {{8{_T_65226[5]}},_T_65226}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_269 = {{9{_T_65233[4]}},_T_65233}; // @[Modules.scala 112:22:@8.4]
  assign _T_65939 = $signed(buffer_3_268) + $signed(buffer_3_269); // @[Modules.scala 160:64:@12092.4]
  assign _T_65940 = _T_65939[13:0]; // @[Modules.scala 160:64:@12093.4]
  assign buffer_3_448 = $signed(_T_65940); // @[Modules.scala 160:64:@12094.4]
  assign buffer_3_270 = {{8{_T_65240[5]}},_T_65240}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_271 = {{9{_T_65247[4]}},_T_65247}; // @[Modules.scala 112:22:@8.4]
  assign _T_65942 = $signed(buffer_3_270) + $signed(buffer_3_271); // @[Modules.scala 160:64:@12096.4]
  assign _T_65943 = _T_65942[13:0]; // @[Modules.scala 160:64:@12097.4]
  assign buffer_3_449 = $signed(_T_65943); // @[Modules.scala 160:64:@12098.4]
  assign buffer_3_272 = {{9{_T_65254[4]}},_T_65254}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_273 = {{9{_T_65261[4]}},_T_65261}; // @[Modules.scala 112:22:@8.4]
  assign _T_65945 = $signed(buffer_3_272) + $signed(buffer_3_273); // @[Modules.scala 160:64:@12100.4]
  assign _T_65946 = _T_65945[13:0]; // @[Modules.scala 160:64:@12101.4]
  assign buffer_3_450 = $signed(_T_65946); // @[Modules.scala 160:64:@12102.4]
  assign buffer_3_274 = {{9{_T_65268[4]}},_T_65268}; // @[Modules.scala 112:22:@8.4]
  assign _T_65948 = $signed(buffer_3_274) + $signed(buffer_1_265); // @[Modules.scala 160:64:@12104.4]
  assign _T_65949 = _T_65948[13:0]; // @[Modules.scala 160:64:@12105.4]
  assign buffer_3_451 = $signed(_T_65949); // @[Modules.scala 160:64:@12106.4]
  assign buffer_3_276 = {{9{_T_65282[4]}},_T_65282}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_277 = {{8{_T_65289[5]}},_T_65289}; // @[Modules.scala 112:22:@8.4]
  assign _T_65951 = $signed(buffer_3_276) + $signed(buffer_3_277); // @[Modules.scala 160:64:@12108.4]
  assign _T_65952 = _T_65951[13:0]; // @[Modules.scala 160:64:@12109.4]
  assign buffer_3_452 = $signed(_T_65952); // @[Modules.scala 160:64:@12110.4]
  assign buffer_3_279 = {{8{_T_65303[5]}},_T_65303}; // @[Modules.scala 112:22:@8.4]
  assign _T_65954 = $signed(buffer_1_268) + $signed(buffer_3_279); // @[Modules.scala 160:64:@12112.4]
  assign _T_65955 = _T_65954[13:0]; // @[Modules.scala 160:64:@12113.4]
  assign buffer_3_453 = $signed(_T_65955); // @[Modules.scala 160:64:@12114.4]
  assign buffer_3_280 = {{8{_T_65310[5]}},_T_65310}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_281 = {{8{_T_65317[5]}},_T_65317}; // @[Modules.scala 112:22:@8.4]
  assign _T_65957 = $signed(buffer_3_280) + $signed(buffer_3_281); // @[Modules.scala 160:64:@12116.4]
  assign _T_65958 = _T_65957[13:0]; // @[Modules.scala 160:64:@12117.4]
  assign buffer_3_454 = $signed(_T_65958); // @[Modules.scala 160:64:@12118.4]
  assign buffer_3_283 = {{8{_T_65331[5]}},_T_65331}; // @[Modules.scala 112:22:@8.4]
  assign _T_65960 = $signed(buffer_0_273) + $signed(buffer_3_283); // @[Modules.scala 160:64:@12120.4]
  assign _T_65961 = _T_65960[13:0]; // @[Modules.scala 160:64:@12121.4]
  assign buffer_3_455 = $signed(_T_65961); // @[Modules.scala 160:64:@12122.4]
  assign buffer_3_284 = {{9{_T_65338[4]}},_T_65338}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_285 = {{9{_T_65345[4]}},_T_65345}; // @[Modules.scala 112:22:@8.4]
  assign _T_65963 = $signed(buffer_3_284) + $signed(buffer_3_285); // @[Modules.scala 160:64:@12124.4]
  assign _T_65964 = _T_65963[13:0]; // @[Modules.scala 160:64:@12125.4]
  assign buffer_3_456 = $signed(_T_65964); // @[Modules.scala 160:64:@12126.4]
  assign buffer_3_286 = {{9{_T_65352[4]}},_T_65352}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_287 = {{9{_T_65359[4]}},_T_65359}; // @[Modules.scala 112:22:@8.4]
  assign _T_65966 = $signed(buffer_3_286) + $signed(buffer_3_287); // @[Modules.scala 160:64:@12128.4]
  assign _T_65967 = _T_65966[13:0]; // @[Modules.scala 160:64:@12129.4]
  assign buffer_3_457 = $signed(_T_65967); // @[Modules.scala 160:64:@12130.4]
  assign buffer_3_289 = {{8{_T_65373[5]}},_T_65373}; // @[Modules.scala 112:22:@8.4]
  assign _T_65969 = $signed(buffer_2_284) + $signed(buffer_3_289); // @[Modules.scala 160:64:@12132.4]
  assign _T_65970 = _T_65969[13:0]; // @[Modules.scala 160:64:@12133.4]
  assign buffer_3_458 = $signed(_T_65970); // @[Modules.scala 160:64:@12134.4]
  assign buffer_3_291 = {{8{_T_65387[5]}},_T_65387}; // @[Modules.scala 112:22:@8.4]
  assign _T_65972 = $signed(buffer_1_281) + $signed(buffer_3_291); // @[Modules.scala 160:64:@12136.4]
  assign _T_65973 = _T_65972[13:0]; // @[Modules.scala 160:64:@12137.4]
  assign buffer_3_459 = $signed(_T_65973); // @[Modules.scala 160:64:@12138.4]
  assign buffer_3_292 = {{9{_T_65394[4]}},_T_65394}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_293 = {{8{_T_65401[5]}},_T_65401}; // @[Modules.scala 112:22:@8.4]
  assign _T_65975 = $signed(buffer_3_292) + $signed(buffer_3_293); // @[Modules.scala 160:64:@12140.4]
  assign _T_65976 = _T_65975[13:0]; // @[Modules.scala 160:64:@12141.4]
  assign buffer_3_460 = $signed(_T_65976); // @[Modules.scala 160:64:@12142.4]
  assign buffer_3_294 = {{8{_T_65408[5]}},_T_65408}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_295 = {{9{_T_65415[4]}},_T_65415}; // @[Modules.scala 112:22:@8.4]
  assign _T_65978 = $signed(buffer_3_294) + $signed(buffer_3_295); // @[Modules.scala 160:64:@12144.4]
  assign _T_65979 = _T_65978[13:0]; // @[Modules.scala 160:64:@12145.4]
  assign buffer_3_461 = $signed(_T_65979); // @[Modules.scala 160:64:@12146.4]
  assign _T_65981 = $signed(buffer_2_293) + $signed(buffer_2_294); // @[Modules.scala 160:64:@12148.4]
  assign _T_65982 = _T_65981[13:0]; // @[Modules.scala 160:64:@12149.4]
  assign buffer_3_462 = $signed(_T_65982); // @[Modules.scala 160:64:@12150.4]
  assign _T_65984 = $signed(buffer_2_295) + $signed(buffer_2_296); // @[Modules.scala 160:64:@12152.4]
  assign _T_65985 = _T_65984[13:0]; // @[Modules.scala 160:64:@12153.4]
  assign buffer_3_463 = $signed(_T_65985); // @[Modules.scala 160:64:@12154.4]
  assign buffer_3_301 = {{9{_T_65457[4]}},_T_65457}; // @[Modules.scala 112:22:@8.4]
  assign _T_65987 = $signed(buffer_2_297) + $signed(buffer_3_301); // @[Modules.scala 160:64:@12156.4]
  assign _T_65988 = _T_65987[13:0]; // @[Modules.scala 160:64:@12157.4]
  assign buffer_3_464 = $signed(_T_65988); // @[Modules.scala 160:64:@12158.4]
  assign buffer_3_303 = {{8{_T_65471[5]}},_T_65471}; // @[Modules.scala 112:22:@8.4]
  assign _T_65990 = $signed(buffer_2_299) + $signed(buffer_3_303); // @[Modules.scala 160:64:@12160.4]
  assign _T_65991 = _T_65990[13:0]; // @[Modules.scala 160:64:@12161.4]
  assign buffer_3_465 = $signed(_T_65991); // @[Modules.scala 160:64:@12162.4]
  assign buffer_3_304 = {{9{_T_65478[4]}},_T_65478}; // @[Modules.scala 112:22:@8.4]
  assign _T_65993 = $signed(buffer_3_304) + $signed(buffer_2_302); // @[Modules.scala 160:64:@12164.4]
  assign _T_65994 = _T_65993[13:0]; // @[Modules.scala 160:64:@12165.4]
  assign buffer_3_466 = $signed(_T_65994); // @[Modules.scala 160:64:@12166.4]
  assign _T_65996 = $signed(buffer_2_303) + $signed(buffer_2_304); // @[Modules.scala 160:64:@12168.4]
  assign _T_65997 = _T_65996[13:0]; // @[Modules.scala 160:64:@12169.4]
  assign buffer_3_467 = $signed(_T_65997); // @[Modules.scala 160:64:@12170.4]
  assign _T_65999 = $signed(buffer_2_305) + $signed(buffer_2_306); // @[Modules.scala 160:64:@12172.4]
  assign _T_66000 = _T_65999[13:0]; // @[Modules.scala 160:64:@12173.4]
  assign buffer_3_468 = $signed(_T_66000); // @[Modules.scala 160:64:@12174.4]
  assign buffer_3_311 = {{9{_T_65527[4]}},_T_65527}; // @[Modules.scala 112:22:@8.4]
  assign _T_66002 = $signed(buffer_2_307) + $signed(buffer_3_311); // @[Modules.scala 160:64:@12176.4]
  assign _T_66003 = _T_66002[13:0]; // @[Modules.scala 160:64:@12177.4]
  assign buffer_3_469 = $signed(_T_66003); // @[Modules.scala 160:64:@12178.4]
  assign buffer_3_312 = {{9{_T_65534[4]}},_T_65534}; // @[Modules.scala 112:22:@8.4]
  assign buffer_3_313 = {{9{_T_59332[4]}},_T_59332}; // @[Modules.scala 112:22:@8.4]
  assign _T_66005 = $signed(buffer_3_312) + $signed(buffer_3_313); // @[Modules.scala 160:64:@12180.4]
  assign _T_66006 = _T_66005[13:0]; // @[Modules.scala 160:64:@12181.4]
  assign buffer_3_470 = $signed(_T_66006); // @[Modules.scala 160:64:@12182.4]
  assign _T_66008 = $signed(buffer_2_310) + $signed(buffer_3_315); // @[Modules.scala 166:64:@12184.4]
  assign _T_66009 = _T_66008[13:0]; // @[Modules.scala 166:64:@12185.4]
  assign buffer_3_471 = $signed(_T_66009); // @[Modules.scala 166:64:@12186.4]
  assign _T_66011 = $signed(buffer_3_316) + $signed(buffer_3_317); // @[Modules.scala 166:64:@12188.4]
  assign _T_66012 = _T_66011[13:0]; // @[Modules.scala 166:64:@12189.4]
  assign buffer_3_472 = $signed(_T_66012); // @[Modules.scala 166:64:@12190.4]
  assign _T_66014 = $signed(buffer_3_318) + $signed(buffer_3_319); // @[Modules.scala 166:64:@12192.4]
  assign _T_66015 = _T_66014[13:0]; // @[Modules.scala 166:64:@12193.4]
  assign buffer_3_473 = $signed(_T_66015); // @[Modules.scala 166:64:@12194.4]
  assign _T_66017 = $signed(buffer_3_320) + $signed(buffer_2_317); // @[Modules.scala 166:64:@12196.4]
  assign _T_66018 = _T_66017[13:0]; // @[Modules.scala 166:64:@12197.4]
  assign buffer_3_474 = $signed(_T_66018); // @[Modules.scala 166:64:@12198.4]
  assign _T_66020 = $signed(buffer_3_322) + $signed(buffer_3_323); // @[Modules.scala 166:64:@12200.4]
  assign _T_66021 = _T_66020[13:0]; // @[Modules.scala 166:64:@12201.4]
  assign buffer_3_475 = $signed(_T_66021); // @[Modules.scala 166:64:@12202.4]
  assign _T_66023 = $signed(buffer_3_324) + $signed(buffer_3_325); // @[Modules.scala 166:64:@12204.4]
  assign _T_66024 = _T_66023[13:0]; // @[Modules.scala 166:64:@12205.4]
  assign buffer_3_476 = $signed(_T_66024); // @[Modules.scala 166:64:@12206.4]
  assign _T_66026 = $signed(buffer_3_326) + $signed(buffer_3_327); // @[Modules.scala 166:64:@12208.4]
  assign _T_66027 = _T_66026[13:0]; // @[Modules.scala 166:64:@12209.4]
  assign buffer_3_477 = $signed(_T_66027); // @[Modules.scala 166:64:@12210.4]
  assign _T_66029 = $signed(buffer_3_328) + $signed(buffer_3_329); // @[Modules.scala 166:64:@12212.4]
  assign _T_66030 = _T_66029[13:0]; // @[Modules.scala 166:64:@12213.4]
  assign buffer_3_478 = $signed(_T_66030); // @[Modules.scala 166:64:@12214.4]
  assign _T_66032 = $signed(buffer_3_330) + $signed(buffer_3_331); // @[Modules.scala 166:64:@12216.4]
  assign _T_66033 = _T_66032[13:0]; // @[Modules.scala 166:64:@12217.4]
  assign buffer_3_479 = $signed(_T_66033); // @[Modules.scala 166:64:@12218.4]
  assign _T_66035 = $signed(buffer_3_332) + $signed(buffer_3_333); // @[Modules.scala 166:64:@12220.4]
  assign _T_66036 = _T_66035[13:0]; // @[Modules.scala 166:64:@12221.4]
  assign buffer_3_480 = $signed(_T_66036); // @[Modules.scala 166:64:@12222.4]
  assign _T_66038 = $signed(buffer_3_334) + $signed(buffer_3_335); // @[Modules.scala 166:64:@12224.4]
  assign _T_66039 = _T_66038[13:0]; // @[Modules.scala 166:64:@12225.4]
  assign buffer_3_481 = $signed(_T_66039); // @[Modules.scala 166:64:@12226.4]
  assign _T_66041 = $signed(buffer_3_336) + $signed(buffer_3_337); // @[Modules.scala 166:64:@12228.4]
  assign _T_66042 = _T_66041[13:0]; // @[Modules.scala 166:64:@12229.4]
  assign buffer_3_482 = $signed(_T_66042); // @[Modules.scala 166:64:@12230.4]
  assign _T_66044 = $signed(buffer_3_338) + $signed(buffer_3_339); // @[Modules.scala 166:64:@12232.4]
  assign _T_66045 = _T_66044[13:0]; // @[Modules.scala 166:64:@12233.4]
  assign buffer_3_483 = $signed(_T_66045); // @[Modules.scala 166:64:@12234.4]
  assign _T_66047 = $signed(buffer_3_340) + $signed(buffer_3_341); // @[Modules.scala 166:64:@12236.4]
  assign _T_66048 = _T_66047[13:0]; // @[Modules.scala 166:64:@12237.4]
  assign buffer_3_484 = $signed(_T_66048); // @[Modules.scala 166:64:@12238.4]
  assign _T_66050 = $signed(buffer_3_342) + $signed(buffer_3_343); // @[Modules.scala 166:64:@12240.4]
  assign _T_66051 = _T_66050[13:0]; // @[Modules.scala 166:64:@12241.4]
  assign buffer_3_485 = $signed(_T_66051); // @[Modules.scala 166:64:@12242.4]
  assign _T_66053 = $signed(buffer_3_344) + $signed(buffer_3_345); // @[Modules.scala 166:64:@12244.4]
  assign _T_66054 = _T_66053[13:0]; // @[Modules.scala 166:64:@12245.4]
  assign buffer_3_486 = $signed(_T_66054); // @[Modules.scala 166:64:@12246.4]
  assign _T_66056 = $signed(buffer_3_346) + $signed(buffer_3_347); // @[Modules.scala 166:64:@12248.4]
  assign _T_66057 = _T_66056[13:0]; // @[Modules.scala 166:64:@12249.4]
  assign buffer_3_487 = $signed(_T_66057); // @[Modules.scala 166:64:@12250.4]
  assign _T_66059 = $signed(buffer_3_348) + $signed(buffer_3_349); // @[Modules.scala 166:64:@12252.4]
  assign _T_66060 = _T_66059[13:0]; // @[Modules.scala 166:64:@12253.4]
  assign buffer_3_488 = $signed(_T_66060); // @[Modules.scala 166:64:@12254.4]
  assign _T_66062 = $signed(buffer_3_350) + $signed(buffer_3_351); // @[Modules.scala 166:64:@12256.4]
  assign _T_66063 = _T_66062[13:0]; // @[Modules.scala 166:64:@12257.4]
  assign buffer_3_489 = $signed(_T_66063); // @[Modules.scala 166:64:@12258.4]
  assign _T_66065 = $signed(buffer_3_352) + $signed(buffer_3_353); // @[Modules.scala 166:64:@12260.4]
  assign _T_66066 = _T_66065[13:0]; // @[Modules.scala 166:64:@12261.4]
  assign buffer_3_490 = $signed(_T_66066); // @[Modules.scala 166:64:@12262.4]
  assign _T_66068 = $signed(buffer_3_354) + $signed(buffer_2_350); // @[Modules.scala 166:64:@12264.4]
  assign _T_66069 = _T_66068[13:0]; // @[Modules.scala 166:64:@12265.4]
  assign buffer_3_491 = $signed(_T_66069); // @[Modules.scala 166:64:@12266.4]
  assign _T_66071 = $signed(buffer_3_356) + $signed(buffer_3_357); // @[Modules.scala 166:64:@12268.4]
  assign _T_66072 = _T_66071[13:0]; // @[Modules.scala 166:64:@12269.4]
  assign buffer_3_492 = $signed(_T_66072); // @[Modules.scala 166:64:@12270.4]
  assign _T_66074 = $signed(buffer_3_358) + $signed(buffer_3_359); // @[Modules.scala 166:64:@12272.4]
  assign _T_66075 = _T_66074[13:0]; // @[Modules.scala 166:64:@12273.4]
  assign buffer_3_493 = $signed(_T_66075); // @[Modules.scala 166:64:@12274.4]
  assign _T_66077 = $signed(buffer_3_360) + $signed(buffer_3_361); // @[Modules.scala 166:64:@12276.4]
  assign _T_66078 = _T_66077[13:0]; // @[Modules.scala 166:64:@12277.4]
  assign buffer_3_494 = $signed(_T_66078); // @[Modules.scala 166:64:@12278.4]
  assign _T_66080 = $signed(buffer_3_362) + $signed(buffer_3_363); // @[Modules.scala 166:64:@12280.4]
  assign _T_66081 = _T_66080[13:0]; // @[Modules.scala 166:64:@12281.4]
  assign buffer_3_495 = $signed(_T_66081); // @[Modules.scala 166:64:@12282.4]
  assign _T_66083 = $signed(buffer_0_349) + $signed(buffer_3_365); // @[Modules.scala 166:64:@12284.4]
  assign _T_66084 = _T_66083[13:0]; // @[Modules.scala 166:64:@12285.4]
  assign buffer_3_496 = $signed(_T_66084); // @[Modules.scala 166:64:@12286.4]
  assign _T_66086 = $signed(buffer_3_366) + $signed(buffer_3_367); // @[Modules.scala 166:64:@12288.4]
  assign _T_66087 = _T_66086[13:0]; // @[Modules.scala 166:64:@12289.4]
  assign buffer_3_497 = $signed(_T_66087); // @[Modules.scala 166:64:@12290.4]
  assign _T_66089 = $signed(buffer_3_368) + $signed(buffer_3_369); // @[Modules.scala 166:64:@12292.4]
  assign _T_66090 = _T_66089[13:0]; // @[Modules.scala 166:64:@12293.4]
  assign buffer_3_498 = $signed(_T_66090); // @[Modules.scala 166:64:@12294.4]
  assign _T_66092 = $signed(buffer_3_370) + $signed(buffer_0_356); // @[Modules.scala 166:64:@12296.4]
  assign _T_66093 = _T_66092[13:0]; // @[Modules.scala 166:64:@12297.4]
  assign buffer_3_499 = $signed(_T_66093); // @[Modules.scala 166:64:@12298.4]
  assign _T_66095 = $signed(buffer_3_372) + $signed(buffer_3_373); // @[Modules.scala 166:64:@12300.4]
  assign _T_66096 = _T_66095[13:0]; // @[Modules.scala 166:64:@12301.4]
  assign buffer_3_500 = $signed(_T_66096); // @[Modules.scala 166:64:@12302.4]
  assign _T_66098 = $signed(buffer_3_374) + $signed(buffer_3_375); // @[Modules.scala 166:64:@12304.4]
  assign _T_66099 = _T_66098[13:0]; // @[Modules.scala 166:64:@12305.4]
  assign buffer_3_501 = $signed(_T_66099); // @[Modules.scala 166:64:@12306.4]
  assign _T_66101 = $signed(buffer_3_376) + $signed(buffer_3_377); // @[Modules.scala 166:64:@12308.4]
  assign _T_66102 = _T_66101[13:0]; // @[Modules.scala 166:64:@12309.4]
  assign buffer_3_502 = $signed(_T_66102); // @[Modules.scala 166:64:@12310.4]
  assign _T_66104 = $signed(buffer_3_378) + $signed(buffer_3_379); // @[Modules.scala 166:64:@12312.4]
  assign _T_66105 = _T_66104[13:0]; // @[Modules.scala 166:64:@12313.4]
  assign buffer_3_503 = $signed(_T_66105); // @[Modules.scala 166:64:@12314.4]
  assign _T_66107 = $signed(buffer_3_380) + $signed(buffer_3_381); // @[Modules.scala 166:64:@12316.4]
  assign _T_66108 = _T_66107[13:0]; // @[Modules.scala 166:64:@12317.4]
  assign buffer_3_504 = $signed(_T_66108); // @[Modules.scala 166:64:@12318.4]
  assign _T_66110 = $signed(buffer_3_382) + $signed(buffer_3_383); // @[Modules.scala 166:64:@12320.4]
  assign _T_66111 = _T_66110[13:0]; // @[Modules.scala 166:64:@12321.4]
  assign buffer_3_505 = $signed(_T_66111); // @[Modules.scala 166:64:@12322.4]
  assign _T_66113 = $signed(buffer_3_384) + $signed(buffer_3_385); // @[Modules.scala 166:64:@12324.4]
  assign _T_66114 = _T_66113[13:0]; // @[Modules.scala 166:64:@12325.4]
  assign buffer_3_506 = $signed(_T_66114); // @[Modules.scala 166:64:@12326.4]
  assign _T_66116 = $signed(buffer_3_386) + $signed(buffer_3_387); // @[Modules.scala 166:64:@12328.4]
  assign _T_66117 = _T_66116[13:0]; // @[Modules.scala 166:64:@12329.4]
  assign buffer_3_507 = $signed(_T_66117); // @[Modules.scala 166:64:@12330.4]
  assign _T_66122 = $signed(buffer_3_390) + $signed(buffer_3_391); // @[Modules.scala 166:64:@12336.4]
  assign _T_66123 = _T_66122[13:0]; // @[Modules.scala 166:64:@12337.4]
  assign buffer_3_509 = $signed(_T_66123); // @[Modules.scala 166:64:@12338.4]
  assign _T_66125 = $signed(buffer_3_392) + $signed(buffer_3_393); // @[Modules.scala 166:64:@12340.4]
  assign _T_66126 = _T_66125[13:0]; // @[Modules.scala 166:64:@12341.4]
  assign buffer_3_510 = $signed(_T_66126); // @[Modules.scala 166:64:@12342.4]
  assign _T_66128 = $signed(buffer_3_394) + $signed(buffer_3_395); // @[Modules.scala 166:64:@12344.4]
  assign _T_66129 = _T_66128[13:0]; // @[Modules.scala 166:64:@12345.4]
  assign buffer_3_511 = $signed(_T_66129); // @[Modules.scala 166:64:@12346.4]
  assign _T_66131 = $signed(buffer_3_396) + $signed(buffer_3_397); // @[Modules.scala 166:64:@12348.4]
  assign _T_66132 = _T_66131[13:0]; // @[Modules.scala 166:64:@12349.4]
  assign buffer_3_512 = $signed(_T_66132); // @[Modules.scala 166:64:@12350.4]
  assign _T_66134 = $signed(buffer_3_398) + $signed(buffer_3_399); // @[Modules.scala 166:64:@12352.4]
  assign _T_66135 = _T_66134[13:0]; // @[Modules.scala 166:64:@12353.4]
  assign buffer_3_513 = $signed(_T_66135); // @[Modules.scala 166:64:@12354.4]
  assign _T_66137 = $signed(buffer_3_400) + $signed(buffer_3_401); // @[Modules.scala 166:64:@12356.4]
  assign _T_66138 = _T_66137[13:0]; // @[Modules.scala 166:64:@12357.4]
  assign buffer_3_514 = $signed(_T_66138); // @[Modules.scala 166:64:@12358.4]
  assign _T_66140 = $signed(buffer_3_402) + $signed(buffer_3_403); // @[Modules.scala 166:64:@12360.4]
  assign _T_66141 = _T_66140[13:0]; // @[Modules.scala 166:64:@12361.4]
  assign buffer_3_515 = $signed(_T_66141); // @[Modules.scala 166:64:@12362.4]
  assign _T_66143 = $signed(buffer_3_404) + $signed(buffer_3_405); // @[Modules.scala 166:64:@12364.4]
  assign _T_66144 = _T_66143[13:0]; // @[Modules.scala 166:64:@12365.4]
  assign buffer_3_516 = $signed(_T_66144); // @[Modules.scala 166:64:@12366.4]
  assign _T_66146 = $signed(buffer_3_406) + $signed(buffer_3_407); // @[Modules.scala 166:64:@12368.4]
  assign _T_66147 = _T_66146[13:0]; // @[Modules.scala 166:64:@12369.4]
  assign buffer_3_517 = $signed(_T_66147); // @[Modules.scala 166:64:@12370.4]
  assign _T_66149 = $signed(buffer_3_408) + $signed(buffer_3_409); // @[Modules.scala 166:64:@12372.4]
  assign _T_66150 = _T_66149[13:0]; // @[Modules.scala 166:64:@12373.4]
  assign buffer_3_518 = $signed(_T_66150); // @[Modules.scala 166:64:@12374.4]
  assign _T_66152 = $signed(buffer_3_410) + $signed(buffer_3_411); // @[Modules.scala 166:64:@12376.4]
  assign _T_66153 = _T_66152[13:0]; // @[Modules.scala 166:64:@12377.4]
  assign buffer_3_519 = $signed(_T_66153); // @[Modules.scala 166:64:@12378.4]
  assign _T_66155 = $signed(buffer_3_412) + $signed(buffer_3_413); // @[Modules.scala 166:64:@12380.4]
  assign _T_66156 = _T_66155[13:0]; // @[Modules.scala 166:64:@12381.4]
  assign buffer_3_520 = $signed(_T_66156); // @[Modules.scala 166:64:@12382.4]
  assign _T_66158 = $signed(buffer_3_414) + $signed(buffer_3_415); // @[Modules.scala 166:64:@12384.4]
  assign _T_66159 = _T_66158[13:0]; // @[Modules.scala 166:64:@12385.4]
  assign buffer_3_521 = $signed(_T_66159); // @[Modules.scala 166:64:@12386.4]
  assign _T_66161 = $signed(buffer_3_416) + $signed(buffer_3_417); // @[Modules.scala 166:64:@12388.4]
  assign _T_66162 = _T_66161[13:0]; // @[Modules.scala 166:64:@12389.4]
  assign buffer_3_522 = $signed(_T_66162); // @[Modules.scala 166:64:@12390.4]
  assign _T_66164 = $signed(buffer_3_418) + $signed(buffer_3_419); // @[Modules.scala 166:64:@12392.4]
  assign _T_66165 = _T_66164[13:0]; // @[Modules.scala 166:64:@12393.4]
  assign buffer_3_523 = $signed(_T_66165); // @[Modules.scala 166:64:@12394.4]
  assign _T_66167 = $signed(buffer_3_420) + $signed(buffer_3_421); // @[Modules.scala 166:64:@12396.4]
  assign _T_66168 = _T_66167[13:0]; // @[Modules.scala 166:64:@12397.4]
  assign buffer_3_524 = $signed(_T_66168); // @[Modules.scala 166:64:@12398.4]
  assign _T_66170 = $signed(buffer_3_422) + $signed(buffer_3_423); // @[Modules.scala 166:64:@12400.4]
  assign _T_66171 = _T_66170[13:0]; // @[Modules.scala 166:64:@12401.4]
  assign buffer_3_525 = $signed(_T_66171); // @[Modules.scala 166:64:@12402.4]
  assign _T_66173 = $signed(buffer_3_424) + $signed(buffer_3_425); // @[Modules.scala 166:64:@12404.4]
  assign _T_66174 = _T_66173[13:0]; // @[Modules.scala 166:64:@12405.4]
  assign buffer_3_526 = $signed(_T_66174); // @[Modules.scala 166:64:@12406.4]
  assign _T_66176 = $signed(buffer_3_426) + $signed(buffer_3_427); // @[Modules.scala 166:64:@12408.4]
  assign _T_66177 = _T_66176[13:0]; // @[Modules.scala 166:64:@12409.4]
  assign buffer_3_527 = $signed(_T_66177); // @[Modules.scala 166:64:@12410.4]
  assign _T_66179 = $signed(buffer_3_428) + $signed(buffer_2_422); // @[Modules.scala 166:64:@12412.4]
  assign _T_66180 = _T_66179[13:0]; // @[Modules.scala 166:64:@12413.4]
  assign buffer_3_528 = $signed(_T_66180); // @[Modules.scala 166:64:@12414.4]
  assign _T_66182 = $signed(buffer_3_430) + $signed(buffer_3_431); // @[Modules.scala 166:64:@12416.4]
  assign _T_66183 = _T_66182[13:0]; // @[Modules.scala 166:64:@12417.4]
  assign buffer_3_529 = $signed(_T_66183); // @[Modules.scala 166:64:@12418.4]
  assign _T_66185 = $signed(buffer_3_432) + $signed(buffer_3_433); // @[Modules.scala 166:64:@12420.4]
  assign _T_66186 = _T_66185[13:0]; // @[Modules.scala 166:64:@12421.4]
  assign buffer_3_530 = $signed(_T_66186); // @[Modules.scala 166:64:@12422.4]
  assign _T_66188 = $signed(buffer_3_434) + $signed(buffer_3_435); // @[Modules.scala 166:64:@12424.4]
  assign _T_66189 = _T_66188[13:0]; // @[Modules.scala 166:64:@12425.4]
  assign buffer_3_531 = $signed(_T_66189); // @[Modules.scala 166:64:@12426.4]
  assign _T_66191 = $signed(buffer_3_436) + $signed(buffer_3_437); // @[Modules.scala 166:64:@12428.4]
  assign _T_66192 = _T_66191[13:0]; // @[Modules.scala 166:64:@12429.4]
  assign buffer_3_532 = $signed(_T_66192); // @[Modules.scala 166:64:@12430.4]
  assign _T_66194 = $signed(buffer_3_438) + $signed(buffer_3_439); // @[Modules.scala 166:64:@12432.4]
  assign _T_66195 = _T_66194[13:0]; // @[Modules.scala 166:64:@12433.4]
  assign buffer_3_533 = $signed(_T_66195); // @[Modules.scala 166:64:@12434.4]
  assign _T_66197 = $signed(buffer_3_440) + $signed(buffer_3_441); // @[Modules.scala 166:64:@12436.4]
  assign _T_66198 = _T_66197[13:0]; // @[Modules.scala 166:64:@12437.4]
  assign buffer_3_534 = $signed(_T_66198); // @[Modules.scala 166:64:@12438.4]
  assign _T_66200 = $signed(buffer_3_442) + $signed(buffer_3_443); // @[Modules.scala 166:64:@12440.4]
  assign _T_66201 = _T_66200[13:0]; // @[Modules.scala 166:64:@12441.4]
  assign buffer_3_535 = $signed(_T_66201); // @[Modules.scala 166:64:@12442.4]
  assign _T_66203 = $signed(buffer_3_444) + $signed(buffer_3_445); // @[Modules.scala 166:64:@12444.4]
  assign _T_66204 = _T_66203[13:0]; // @[Modules.scala 166:64:@12445.4]
  assign buffer_3_536 = $signed(_T_66204); // @[Modules.scala 166:64:@12446.4]
  assign _T_66206 = $signed(buffer_3_446) + $signed(buffer_3_447); // @[Modules.scala 166:64:@12448.4]
  assign _T_66207 = _T_66206[13:0]; // @[Modules.scala 166:64:@12449.4]
  assign buffer_3_537 = $signed(_T_66207); // @[Modules.scala 166:64:@12450.4]
  assign _T_66209 = $signed(buffer_3_448) + $signed(buffer_3_449); // @[Modules.scala 166:64:@12452.4]
  assign _T_66210 = _T_66209[13:0]; // @[Modules.scala 166:64:@12453.4]
  assign buffer_3_538 = $signed(_T_66210); // @[Modules.scala 166:64:@12454.4]
  assign _T_66212 = $signed(buffer_3_450) + $signed(buffer_3_451); // @[Modules.scala 166:64:@12456.4]
  assign _T_66213 = _T_66212[13:0]; // @[Modules.scala 166:64:@12457.4]
  assign buffer_3_539 = $signed(_T_66213); // @[Modules.scala 166:64:@12458.4]
  assign _T_66215 = $signed(buffer_3_452) + $signed(buffer_3_453); // @[Modules.scala 166:64:@12460.4]
  assign _T_66216 = _T_66215[13:0]; // @[Modules.scala 166:64:@12461.4]
  assign buffer_3_540 = $signed(_T_66216); // @[Modules.scala 166:64:@12462.4]
  assign _T_66218 = $signed(buffer_3_454) + $signed(buffer_3_455); // @[Modules.scala 166:64:@12464.4]
  assign _T_66219 = _T_66218[13:0]; // @[Modules.scala 166:64:@12465.4]
  assign buffer_3_541 = $signed(_T_66219); // @[Modules.scala 166:64:@12466.4]
  assign _T_66221 = $signed(buffer_3_456) + $signed(buffer_3_457); // @[Modules.scala 166:64:@12468.4]
  assign _T_66222 = _T_66221[13:0]; // @[Modules.scala 166:64:@12469.4]
  assign buffer_3_542 = $signed(_T_66222); // @[Modules.scala 166:64:@12470.4]
  assign _T_66224 = $signed(buffer_3_458) + $signed(buffer_3_459); // @[Modules.scala 166:64:@12472.4]
  assign _T_66225 = _T_66224[13:0]; // @[Modules.scala 166:64:@12473.4]
  assign buffer_3_543 = $signed(_T_66225); // @[Modules.scala 166:64:@12474.4]
  assign _T_66227 = $signed(buffer_3_460) + $signed(buffer_3_461); // @[Modules.scala 166:64:@12476.4]
  assign _T_66228 = _T_66227[13:0]; // @[Modules.scala 166:64:@12477.4]
  assign buffer_3_544 = $signed(_T_66228); // @[Modules.scala 166:64:@12478.4]
  assign _T_66230 = $signed(buffer_3_462) + $signed(buffer_3_463); // @[Modules.scala 166:64:@12480.4]
  assign _T_66231 = _T_66230[13:0]; // @[Modules.scala 166:64:@12481.4]
  assign buffer_3_545 = $signed(_T_66231); // @[Modules.scala 166:64:@12482.4]
  assign _T_66233 = $signed(buffer_3_464) + $signed(buffer_3_465); // @[Modules.scala 166:64:@12484.4]
  assign _T_66234 = _T_66233[13:0]; // @[Modules.scala 166:64:@12485.4]
  assign buffer_3_546 = $signed(_T_66234); // @[Modules.scala 166:64:@12486.4]
  assign _T_66236 = $signed(buffer_3_466) + $signed(buffer_3_467); // @[Modules.scala 166:64:@12488.4]
  assign _T_66237 = _T_66236[13:0]; // @[Modules.scala 166:64:@12489.4]
  assign buffer_3_547 = $signed(_T_66237); // @[Modules.scala 166:64:@12490.4]
  assign _T_66239 = $signed(buffer_3_468) + $signed(buffer_3_469); // @[Modules.scala 166:64:@12492.4]
  assign _T_66240 = _T_66239[13:0]; // @[Modules.scala 166:64:@12493.4]
  assign buffer_3_548 = $signed(_T_66240); // @[Modules.scala 166:64:@12494.4]
  assign _T_66242 = $signed(buffer_3_471) + $signed(buffer_3_472); // @[Modules.scala 160:64:@12496.4]
  assign _T_66243 = _T_66242[13:0]; // @[Modules.scala 160:64:@12497.4]
  assign buffer_3_549 = $signed(_T_66243); // @[Modules.scala 160:64:@12498.4]
  assign _T_66245 = $signed(buffer_3_473) + $signed(buffer_3_474); // @[Modules.scala 160:64:@12500.4]
  assign _T_66246 = _T_66245[13:0]; // @[Modules.scala 160:64:@12501.4]
  assign buffer_3_550 = $signed(_T_66246); // @[Modules.scala 160:64:@12502.4]
  assign _T_66248 = $signed(buffer_3_475) + $signed(buffer_3_476); // @[Modules.scala 160:64:@12504.4]
  assign _T_66249 = _T_66248[13:0]; // @[Modules.scala 160:64:@12505.4]
  assign buffer_3_551 = $signed(_T_66249); // @[Modules.scala 160:64:@12506.4]
  assign _T_66251 = $signed(buffer_3_477) + $signed(buffer_3_478); // @[Modules.scala 160:64:@12508.4]
  assign _T_66252 = _T_66251[13:0]; // @[Modules.scala 160:64:@12509.4]
  assign buffer_3_552 = $signed(_T_66252); // @[Modules.scala 160:64:@12510.4]
  assign _T_66254 = $signed(buffer_3_479) + $signed(buffer_3_480); // @[Modules.scala 160:64:@12512.4]
  assign _T_66255 = _T_66254[13:0]; // @[Modules.scala 160:64:@12513.4]
  assign buffer_3_553 = $signed(_T_66255); // @[Modules.scala 160:64:@12514.4]
  assign _T_66257 = $signed(buffer_3_481) + $signed(buffer_3_482); // @[Modules.scala 160:64:@12516.4]
  assign _T_66258 = _T_66257[13:0]; // @[Modules.scala 160:64:@12517.4]
  assign buffer_3_554 = $signed(_T_66258); // @[Modules.scala 160:64:@12518.4]
  assign _T_66260 = $signed(buffer_3_483) + $signed(buffer_3_484); // @[Modules.scala 160:64:@12520.4]
  assign _T_66261 = _T_66260[13:0]; // @[Modules.scala 160:64:@12521.4]
  assign buffer_3_555 = $signed(_T_66261); // @[Modules.scala 160:64:@12522.4]
  assign _T_66263 = $signed(buffer_3_485) + $signed(buffer_3_486); // @[Modules.scala 160:64:@12524.4]
  assign _T_66264 = _T_66263[13:0]; // @[Modules.scala 160:64:@12525.4]
  assign buffer_3_556 = $signed(_T_66264); // @[Modules.scala 160:64:@12526.4]
  assign _T_66266 = $signed(buffer_3_487) + $signed(buffer_3_488); // @[Modules.scala 160:64:@12528.4]
  assign _T_66267 = _T_66266[13:0]; // @[Modules.scala 160:64:@12529.4]
  assign buffer_3_557 = $signed(_T_66267); // @[Modules.scala 160:64:@12530.4]
  assign _T_66269 = $signed(buffer_3_489) + $signed(buffer_3_490); // @[Modules.scala 160:64:@12532.4]
  assign _T_66270 = _T_66269[13:0]; // @[Modules.scala 160:64:@12533.4]
  assign buffer_3_558 = $signed(_T_66270); // @[Modules.scala 160:64:@12534.4]
  assign _T_66272 = $signed(buffer_3_491) + $signed(buffer_3_492); // @[Modules.scala 160:64:@12536.4]
  assign _T_66273 = _T_66272[13:0]; // @[Modules.scala 160:64:@12537.4]
  assign buffer_3_559 = $signed(_T_66273); // @[Modules.scala 160:64:@12538.4]
  assign _T_66275 = $signed(buffer_3_493) + $signed(buffer_3_494); // @[Modules.scala 160:64:@12540.4]
  assign _T_66276 = _T_66275[13:0]; // @[Modules.scala 160:64:@12541.4]
  assign buffer_3_560 = $signed(_T_66276); // @[Modules.scala 160:64:@12542.4]
  assign _T_66278 = $signed(buffer_3_495) + $signed(buffer_3_496); // @[Modules.scala 160:64:@12544.4]
  assign _T_66279 = _T_66278[13:0]; // @[Modules.scala 160:64:@12545.4]
  assign buffer_3_561 = $signed(_T_66279); // @[Modules.scala 160:64:@12546.4]
  assign _T_66281 = $signed(buffer_3_497) + $signed(buffer_3_498); // @[Modules.scala 160:64:@12548.4]
  assign _T_66282 = _T_66281[13:0]; // @[Modules.scala 160:64:@12549.4]
  assign buffer_3_562 = $signed(_T_66282); // @[Modules.scala 160:64:@12550.4]
  assign _T_66284 = $signed(buffer_3_499) + $signed(buffer_3_500); // @[Modules.scala 160:64:@12552.4]
  assign _T_66285 = _T_66284[13:0]; // @[Modules.scala 160:64:@12553.4]
  assign buffer_3_563 = $signed(_T_66285); // @[Modules.scala 160:64:@12554.4]
  assign _T_66287 = $signed(buffer_3_501) + $signed(buffer_3_502); // @[Modules.scala 160:64:@12556.4]
  assign _T_66288 = _T_66287[13:0]; // @[Modules.scala 160:64:@12557.4]
  assign buffer_3_564 = $signed(_T_66288); // @[Modules.scala 160:64:@12558.4]
  assign _T_66290 = $signed(buffer_3_503) + $signed(buffer_3_504); // @[Modules.scala 160:64:@12560.4]
  assign _T_66291 = _T_66290[13:0]; // @[Modules.scala 160:64:@12561.4]
  assign buffer_3_565 = $signed(_T_66291); // @[Modules.scala 160:64:@12562.4]
  assign _T_66293 = $signed(buffer_3_505) + $signed(buffer_3_506); // @[Modules.scala 160:64:@12564.4]
  assign _T_66294 = _T_66293[13:0]; // @[Modules.scala 160:64:@12565.4]
  assign buffer_3_566 = $signed(_T_66294); // @[Modules.scala 160:64:@12566.4]
  assign _T_66296 = $signed(buffer_3_507) + $signed(buffer_2_501); // @[Modules.scala 160:64:@12568.4]
  assign _T_66297 = _T_66296[13:0]; // @[Modules.scala 160:64:@12569.4]
  assign buffer_3_567 = $signed(_T_66297); // @[Modules.scala 160:64:@12570.4]
  assign _T_66299 = $signed(buffer_3_509) + $signed(buffer_3_510); // @[Modules.scala 160:64:@12572.4]
  assign _T_66300 = _T_66299[13:0]; // @[Modules.scala 160:64:@12573.4]
  assign buffer_3_568 = $signed(_T_66300); // @[Modules.scala 160:64:@12574.4]
  assign _T_66302 = $signed(buffer_3_511) + $signed(buffer_3_512); // @[Modules.scala 160:64:@12576.4]
  assign _T_66303 = _T_66302[13:0]; // @[Modules.scala 160:64:@12577.4]
  assign buffer_3_569 = $signed(_T_66303); // @[Modules.scala 160:64:@12578.4]
  assign _T_66305 = $signed(buffer_3_513) + $signed(buffer_3_514); // @[Modules.scala 160:64:@12580.4]
  assign _T_66306 = _T_66305[13:0]; // @[Modules.scala 160:64:@12581.4]
  assign buffer_3_570 = $signed(_T_66306); // @[Modules.scala 160:64:@12582.4]
  assign _T_66308 = $signed(buffer_3_515) + $signed(buffer_3_516); // @[Modules.scala 160:64:@12584.4]
  assign _T_66309 = _T_66308[13:0]; // @[Modules.scala 160:64:@12585.4]
  assign buffer_3_571 = $signed(_T_66309); // @[Modules.scala 160:64:@12586.4]
  assign _T_66311 = $signed(buffer_3_517) + $signed(buffer_3_518); // @[Modules.scala 160:64:@12588.4]
  assign _T_66312 = _T_66311[13:0]; // @[Modules.scala 160:64:@12589.4]
  assign buffer_3_572 = $signed(_T_66312); // @[Modules.scala 160:64:@12590.4]
  assign _T_66314 = $signed(buffer_3_519) + $signed(buffer_3_520); // @[Modules.scala 160:64:@12592.4]
  assign _T_66315 = _T_66314[13:0]; // @[Modules.scala 160:64:@12593.4]
  assign buffer_3_573 = $signed(_T_66315); // @[Modules.scala 160:64:@12594.4]
  assign _T_66317 = $signed(buffer_3_521) + $signed(buffer_3_522); // @[Modules.scala 160:64:@12596.4]
  assign _T_66318 = _T_66317[13:0]; // @[Modules.scala 160:64:@12597.4]
  assign buffer_3_574 = $signed(_T_66318); // @[Modules.scala 160:64:@12598.4]
  assign _T_66320 = $signed(buffer_3_523) + $signed(buffer_3_524); // @[Modules.scala 160:64:@12600.4]
  assign _T_66321 = _T_66320[13:0]; // @[Modules.scala 160:64:@12601.4]
  assign buffer_3_575 = $signed(_T_66321); // @[Modules.scala 160:64:@12602.4]
  assign _T_66323 = $signed(buffer_3_525) + $signed(buffer_3_526); // @[Modules.scala 160:64:@12604.4]
  assign _T_66324 = _T_66323[13:0]; // @[Modules.scala 160:64:@12605.4]
  assign buffer_3_576 = $signed(_T_66324); // @[Modules.scala 160:64:@12606.4]
  assign _T_66326 = $signed(buffer_3_527) + $signed(buffer_3_528); // @[Modules.scala 160:64:@12608.4]
  assign _T_66327 = _T_66326[13:0]; // @[Modules.scala 160:64:@12609.4]
  assign buffer_3_577 = $signed(_T_66327); // @[Modules.scala 160:64:@12610.4]
  assign _T_66329 = $signed(buffer_3_529) + $signed(buffer_3_530); // @[Modules.scala 160:64:@12612.4]
  assign _T_66330 = _T_66329[13:0]; // @[Modules.scala 160:64:@12613.4]
  assign buffer_3_578 = $signed(_T_66330); // @[Modules.scala 160:64:@12614.4]
  assign _T_66332 = $signed(buffer_3_531) + $signed(buffer_3_532); // @[Modules.scala 160:64:@12616.4]
  assign _T_66333 = _T_66332[13:0]; // @[Modules.scala 160:64:@12617.4]
  assign buffer_3_579 = $signed(_T_66333); // @[Modules.scala 160:64:@12618.4]
  assign _T_66335 = $signed(buffer_3_533) + $signed(buffer_3_534); // @[Modules.scala 160:64:@12620.4]
  assign _T_66336 = _T_66335[13:0]; // @[Modules.scala 160:64:@12621.4]
  assign buffer_3_580 = $signed(_T_66336); // @[Modules.scala 160:64:@12622.4]
  assign _T_66338 = $signed(buffer_3_535) + $signed(buffer_3_536); // @[Modules.scala 160:64:@12624.4]
  assign _T_66339 = _T_66338[13:0]; // @[Modules.scala 160:64:@12625.4]
  assign buffer_3_581 = $signed(_T_66339); // @[Modules.scala 160:64:@12626.4]
  assign _T_66341 = $signed(buffer_3_537) + $signed(buffer_3_538); // @[Modules.scala 160:64:@12628.4]
  assign _T_66342 = _T_66341[13:0]; // @[Modules.scala 160:64:@12629.4]
  assign buffer_3_582 = $signed(_T_66342); // @[Modules.scala 160:64:@12630.4]
  assign _T_66344 = $signed(buffer_3_539) + $signed(buffer_3_540); // @[Modules.scala 160:64:@12632.4]
  assign _T_66345 = _T_66344[13:0]; // @[Modules.scala 160:64:@12633.4]
  assign buffer_3_583 = $signed(_T_66345); // @[Modules.scala 160:64:@12634.4]
  assign _T_66347 = $signed(buffer_3_541) + $signed(buffer_3_542); // @[Modules.scala 160:64:@12636.4]
  assign _T_66348 = _T_66347[13:0]; // @[Modules.scala 160:64:@12637.4]
  assign buffer_3_584 = $signed(_T_66348); // @[Modules.scala 160:64:@12638.4]
  assign _T_66350 = $signed(buffer_3_543) + $signed(buffer_3_544); // @[Modules.scala 160:64:@12640.4]
  assign _T_66351 = _T_66350[13:0]; // @[Modules.scala 160:64:@12641.4]
  assign buffer_3_585 = $signed(_T_66351); // @[Modules.scala 160:64:@12642.4]
  assign _T_66353 = $signed(buffer_3_545) + $signed(buffer_3_546); // @[Modules.scala 160:64:@12644.4]
  assign _T_66354 = _T_66353[13:0]; // @[Modules.scala 160:64:@12645.4]
  assign buffer_3_586 = $signed(_T_66354); // @[Modules.scala 160:64:@12646.4]
  assign _T_66356 = $signed(buffer_3_547) + $signed(buffer_3_548); // @[Modules.scala 160:64:@12648.4]
  assign _T_66357 = _T_66356[13:0]; // @[Modules.scala 160:64:@12649.4]
  assign buffer_3_587 = $signed(_T_66357); // @[Modules.scala 160:64:@12650.4]
  assign _T_66359 = $signed(buffer_3_549) + $signed(buffer_3_550); // @[Modules.scala 166:64:@12652.4]
  assign _T_66360 = _T_66359[13:0]; // @[Modules.scala 166:64:@12653.4]
  assign buffer_3_588 = $signed(_T_66360); // @[Modules.scala 166:64:@12654.4]
  assign _T_66362 = $signed(buffer_3_551) + $signed(buffer_3_552); // @[Modules.scala 166:64:@12656.4]
  assign _T_66363 = _T_66362[13:0]; // @[Modules.scala 166:64:@12657.4]
  assign buffer_3_589 = $signed(_T_66363); // @[Modules.scala 166:64:@12658.4]
  assign _T_66365 = $signed(buffer_3_553) + $signed(buffer_3_554); // @[Modules.scala 166:64:@12660.4]
  assign _T_66366 = _T_66365[13:0]; // @[Modules.scala 166:64:@12661.4]
  assign buffer_3_590 = $signed(_T_66366); // @[Modules.scala 166:64:@12662.4]
  assign _T_66368 = $signed(buffer_3_555) + $signed(buffer_3_556); // @[Modules.scala 166:64:@12664.4]
  assign _T_66369 = _T_66368[13:0]; // @[Modules.scala 166:64:@12665.4]
  assign buffer_3_591 = $signed(_T_66369); // @[Modules.scala 166:64:@12666.4]
  assign _T_66371 = $signed(buffer_3_557) + $signed(buffer_3_558); // @[Modules.scala 166:64:@12668.4]
  assign _T_66372 = _T_66371[13:0]; // @[Modules.scala 166:64:@12669.4]
  assign buffer_3_592 = $signed(_T_66372); // @[Modules.scala 166:64:@12670.4]
  assign _T_66374 = $signed(buffer_3_559) + $signed(buffer_3_560); // @[Modules.scala 166:64:@12672.4]
  assign _T_66375 = _T_66374[13:0]; // @[Modules.scala 166:64:@12673.4]
  assign buffer_3_593 = $signed(_T_66375); // @[Modules.scala 166:64:@12674.4]
  assign _T_66377 = $signed(buffer_3_561) + $signed(buffer_3_562); // @[Modules.scala 166:64:@12676.4]
  assign _T_66378 = _T_66377[13:0]; // @[Modules.scala 166:64:@12677.4]
  assign buffer_3_594 = $signed(_T_66378); // @[Modules.scala 166:64:@12678.4]
  assign _T_66380 = $signed(buffer_3_563) + $signed(buffer_3_564); // @[Modules.scala 166:64:@12680.4]
  assign _T_66381 = _T_66380[13:0]; // @[Modules.scala 166:64:@12681.4]
  assign buffer_3_595 = $signed(_T_66381); // @[Modules.scala 166:64:@12682.4]
  assign _T_66383 = $signed(buffer_3_565) + $signed(buffer_3_566); // @[Modules.scala 166:64:@12684.4]
  assign _T_66384 = _T_66383[13:0]; // @[Modules.scala 166:64:@12685.4]
  assign buffer_3_596 = $signed(_T_66384); // @[Modules.scala 166:64:@12686.4]
  assign _T_66386 = $signed(buffer_3_567) + $signed(buffer_3_568); // @[Modules.scala 166:64:@12688.4]
  assign _T_66387 = _T_66386[13:0]; // @[Modules.scala 166:64:@12689.4]
  assign buffer_3_597 = $signed(_T_66387); // @[Modules.scala 166:64:@12690.4]
  assign _T_66389 = $signed(buffer_3_569) + $signed(buffer_3_570); // @[Modules.scala 166:64:@12692.4]
  assign _T_66390 = _T_66389[13:0]; // @[Modules.scala 166:64:@12693.4]
  assign buffer_3_598 = $signed(_T_66390); // @[Modules.scala 166:64:@12694.4]
  assign _T_66392 = $signed(buffer_3_571) + $signed(buffer_3_572); // @[Modules.scala 166:64:@12696.4]
  assign _T_66393 = _T_66392[13:0]; // @[Modules.scala 166:64:@12697.4]
  assign buffer_3_599 = $signed(_T_66393); // @[Modules.scala 166:64:@12698.4]
  assign _T_66395 = $signed(buffer_3_573) + $signed(buffer_3_574); // @[Modules.scala 166:64:@12700.4]
  assign _T_66396 = _T_66395[13:0]; // @[Modules.scala 166:64:@12701.4]
  assign buffer_3_600 = $signed(_T_66396); // @[Modules.scala 166:64:@12702.4]
  assign _T_66398 = $signed(buffer_3_575) + $signed(buffer_3_576); // @[Modules.scala 166:64:@12704.4]
  assign _T_66399 = _T_66398[13:0]; // @[Modules.scala 166:64:@12705.4]
  assign buffer_3_601 = $signed(_T_66399); // @[Modules.scala 166:64:@12706.4]
  assign _T_66401 = $signed(buffer_3_577) + $signed(buffer_3_578); // @[Modules.scala 166:64:@12708.4]
  assign _T_66402 = _T_66401[13:0]; // @[Modules.scala 166:64:@12709.4]
  assign buffer_3_602 = $signed(_T_66402); // @[Modules.scala 166:64:@12710.4]
  assign _T_66404 = $signed(buffer_3_579) + $signed(buffer_3_580); // @[Modules.scala 166:64:@12712.4]
  assign _T_66405 = _T_66404[13:0]; // @[Modules.scala 166:64:@12713.4]
  assign buffer_3_603 = $signed(_T_66405); // @[Modules.scala 166:64:@12714.4]
  assign _T_66407 = $signed(buffer_3_581) + $signed(buffer_3_582); // @[Modules.scala 166:64:@12716.4]
  assign _T_66408 = _T_66407[13:0]; // @[Modules.scala 166:64:@12717.4]
  assign buffer_3_604 = $signed(_T_66408); // @[Modules.scala 166:64:@12718.4]
  assign _T_66410 = $signed(buffer_3_583) + $signed(buffer_3_584); // @[Modules.scala 166:64:@12720.4]
  assign _T_66411 = _T_66410[13:0]; // @[Modules.scala 166:64:@12721.4]
  assign buffer_3_605 = $signed(_T_66411); // @[Modules.scala 166:64:@12722.4]
  assign _T_66413 = $signed(buffer_3_585) + $signed(buffer_3_586); // @[Modules.scala 166:64:@12724.4]
  assign _T_66414 = _T_66413[13:0]; // @[Modules.scala 166:64:@12725.4]
  assign buffer_3_606 = $signed(_T_66414); // @[Modules.scala 166:64:@12726.4]
  assign _T_66416 = $signed(buffer_3_587) + $signed(buffer_3_470); // @[Modules.scala 172:66:@12728.4]
  assign _T_66417 = _T_66416[13:0]; // @[Modules.scala 172:66:@12729.4]
  assign buffer_3_607 = $signed(_T_66417); // @[Modules.scala 172:66:@12730.4]
  assign _T_66419 = $signed(buffer_3_588) + $signed(buffer_3_589); // @[Modules.scala 160:64:@12732.4]
  assign _T_66420 = _T_66419[13:0]; // @[Modules.scala 160:64:@12733.4]
  assign buffer_3_608 = $signed(_T_66420); // @[Modules.scala 160:64:@12734.4]
  assign _T_66422 = $signed(buffer_3_590) + $signed(buffer_3_591); // @[Modules.scala 160:64:@12736.4]
  assign _T_66423 = _T_66422[13:0]; // @[Modules.scala 160:64:@12737.4]
  assign buffer_3_609 = $signed(_T_66423); // @[Modules.scala 160:64:@12738.4]
  assign _T_66425 = $signed(buffer_3_592) + $signed(buffer_3_593); // @[Modules.scala 160:64:@12740.4]
  assign _T_66426 = _T_66425[13:0]; // @[Modules.scala 160:64:@12741.4]
  assign buffer_3_610 = $signed(_T_66426); // @[Modules.scala 160:64:@12742.4]
  assign _T_66428 = $signed(buffer_3_594) + $signed(buffer_3_595); // @[Modules.scala 160:64:@12744.4]
  assign _T_66429 = _T_66428[13:0]; // @[Modules.scala 160:64:@12745.4]
  assign buffer_3_611 = $signed(_T_66429); // @[Modules.scala 160:64:@12746.4]
  assign _T_66431 = $signed(buffer_3_596) + $signed(buffer_3_597); // @[Modules.scala 160:64:@12748.4]
  assign _T_66432 = _T_66431[13:0]; // @[Modules.scala 160:64:@12749.4]
  assign buffer_3_612 = $signed(_T_66432); // @[Modules.scala 160:64:@12750.4]
  assign _T_66434 = $signed(buffer_3_598) + $signed(buffer_3_599); // @[Modules.scala 160:64:@12752.4]
  assign _T_66435 = _T_66434[13:0]; // @[Modules.scala 160:64:@12753.4]
  assign buffer_3_613 = $signed(_T_66435); // @[Modules.scala 160:64:@12754.4]
  assign _T_66437 = $signed(buffer_3_600) + $signed(buffer_3_601); // @[Modules.scala 160:64:@12756.4]
  assign _T_66438 = _T_66437[13:0]; // @[Modules.scala 160:64:@12757.4]
  assign buffer_3_614 = $signed(_T_66438); // @[Modules.scala 160:64:@12758.4]
  assign _T_66440 = $signed(buffer_3_602) + $signed(buffer_3_603); // @[Modules.scala 160:64:@12760.4]
  assign _T_66441 = _T_66440[13:0]; // @[Modules.scala 160:64:@12761.4]
  assign buffer_3_615 = $signed(_T_66441); // @[Modules.scala 160:64:@12762.4]
  assign _T_66443 = $signed(buffer_3_604) + $signed(buffer_3_605); // @[Modules.scala 160:64:@12764.4]
  assign _T_66444 = _T_66443[13:0]; // @[Modules.scala 160:64:@12765.4]
  assign buffer_3_616 = $signed(_T_66444); // @[Modules.scala 160:64:@12766.4]
  assign _T_66446 = $signed(buffer_3_606) + $signed(buffer_3_607); // @[Modules.scala 160:64:@12768.4]
  assign _T_66447 = _T_66446[13:0]; // @[Modules.scala 160:64:@12769.4]
  assign buffer_3_617 = $signed(_T_66447); // @[Modules.scala 160:64:@12770.4]
  assign _T_66449 = $signed(buffer_3_608) + $signed(buffer_3_609); // @[Modules.scala 160:64:@12772.4]
  assign _T_66450 = _T_66449[13:0]; // @[Modules.scala 160:64:@12773.4]
  assign buffer_3_618 = $signed(_T_66450); // @[Modules.scala 160:64:@12774.4]
  assign _T_66452 = $signed(buffer_3_610) + $signed(buffer_3_611); // @[Modules.scala 160:64:@12776.4]
  assign _T_66453 = _T_66452[13:0]; // @[Modules.scala 160:64:@12777.4]
  assign buffer_3_619 = $signed(_T_66453); // @[Modules.scala 160:64:@12778.4]
  assign _T_66455 = $signed(buffer_3_612) + $signed(buffer_3_613); // @[Modules.scala 160:64:@12780.4]
  assign _T_66456 = _T_66455[13:0]; // @[Modules.scala 160:64:@12781.4]
  assign buffer_3_620 = $signed(_T_66456); // @[Modules.scala 160:64:@12782.4]
  assign _T_66458 = $signed(buffer_3_614) + $signed(buffer_3_615); // @[Modules.scala 160:64:@12784.4]
  assign _T_66459 = _T_66458[13:0]; // @[Modules.scala 160:64:@12785.4]
  assign buffer_3_621 = $signed(_T_66459); // @[Modules.scala 160:64:@12786.4]
  assign _T_66461 = $signed(buffer_3_616) + $signed(buffer_3_617); // @[Modules.scala 160:64:@12788.4]
  assign _T_66462 = _T_66461[13:0]; // @[Modules.scala 160:64:@12789.4]
  assign buffer_3_622 = $signed(_T_66462); // @[Modules.scala 160:64:@12790.4]
  assign _T_66464 = $signed(buffer_3_618) + $signed(buffer_3_619); // @[Modules.scala 166:64:@12792.4]
  assign _T_66465 = _T_66464[13:0]; // @[Modules.scala 166:64:@12793.4]
  assign buffer_3_623 = $signed(_T_66465); // @[Modules.scala 166:64:@12794.4]
  assign _T_66467 = $signed(buffer_3_620) + $signed(buffer_3_621); // @[Modules.scala 166:64:@12796.4]
  assign _T_66468 = _T_66467[13:0]; // @[Modules.scala 166:64:@12797.4]
  assign buffer_3_624 = $signed(_T_66468); // @[Modules.scala 166:64:@12798.4]
  assign _T_66470 = $signed(buffer_3_623) + $signed(buffer_3_624); // @[Modules.scala 160:64:@12800.4]
  assign _T_66471 = _T_66470[13:0]; // @[Modules.scala 160:64:@12801.4]
  assign buffer_3_625 = $signed(_T_66471); // @[Modules.scala 160:64:@12802.4]
  assign _T_66473 = $signed(buffer_3_625) + $signed(buffer_3_622); // @[Modules.scala 172:66:@12804.4]
  assign _T_66474 = _T_66473[13:0]; // @[Modules.scala 172:66:@12805.4]
  assign buffer_3_626 = $signed(_T_66474); // @[Modules.scala 172:66:@12806.4]
  assign _T_66491 = $signed(4'sh1) * $signed(io_in_30); // @[Modules.scala 150:74:@12977.4]
  assign _GEN_279 = {{1{_T_60271[4]}},_T_60271}; // @[Modules.scala 150:103:@12979.4]
  assign _T_66494 = $signed(_T_66491) + $signed(_GEN_279); // @[Modules.scala 150:103:@12979.4]
  assign _T_66495 = _T_66494[5:0]; // @[Modules.scala 150:103:@12980.4]
  assign _T_66496 = $signed(_T_66495); // @[Modules.scala 150:103:@12981.4]
  assign _T_66500 = $signed(-4'sh1) * $signed(io_in_38); // @[Modules.scala 151:80:@12984.4]
  assign _T_66501 = $signed(_T_57241) + $signed(_T_66500); // @[Modules.scala 150:103:@12985.4]
  assign _T_66502 = _T_66501[4:0]; // @[Modules.scala 150:103:@12986.4]
  assign _T_66503 = $signed(_T_66502); // @[Modules.scala 150:103:@12987.4]
  assign _T_66508 = $signed(_T_63375) + $signed(_T_57248); // @[Modules.scala 150:103:@12991.4]
  assign _T_66509 = _T_66508[4:0]; // @[Modules.scala 150:103:@12992.4]
  assign _T_66510 = $signed(_T_66509); // @[Modules.scala 150:103:@12993.4]
  assign _T_66522 = $signed(_GEN_144) + $signed(_T_54255); // @[Modules.scala 150:103:@13003.4]
  assign _T_66523 = _T_66522[5:0]; // @[Modules.scala 150:103:@13004.4]
  assign _T_66524 = $signed(_T_66523); // @[Modules.scala 150:103:@13005.4]
  assign _T_66529 = $signed(_T_54257) + $signed(_T_54262); // @[Modules.scala 150:103:@13009.4]
  assign _T_66530 = _T_66529[5:0]; // @[Modules.scala 150:103:@13010.4]
  assign _T_66531 = $signed(_T_66530); // @[Modules.scala 150:103:@13011.4]
  assign _T_66543 = $signed(_T_57276) + $signed(_T_57281); // @[Modules.scala 150:103:@13021.4]
  assign _T_66544 = _T_66543[4:0]; // @[Modules.scala 150:103:@13022.4]
  assign _T_66545 = $signed(_T_66544); // @[Modules.scala 150:103:@13023.4]
  assign _GEN_281 = {{1{_T_60327[4]}},_T_60327}; // @[Modules.scala 150:103:@13027.4]
  assign _T_66550 = $signed(_GEN_281) + $signed(_T_63429); // @[Modules.scala 150:103:@13027.4]
  assign _T_66551 = _T_66550[5:0]; // @[Modules.scala 150:103:@13028.4]
  assign _T_66552 = $signed(_T_66551); // @[Modules.scala 150:103:@13029.4]
  assign _T_66564 = $signed(_T_57297) + $signed(_T_57302); // @[Modules.scala 150:103:@13039.4]
  assign _T_66565 = _T_66564[4:0]; // @[Modules.scala 150:103:@13040.4]
  assign _T_66566 = $signed(_T_66565); // @[Modules.scala 150:103:@13041.4]
  assign _T_66571 = $signed(_T_57304) + $signed(_T_57309); // @[Modules.scala 150:103:@13045.4]
  assign _T_66572 = _T_66571[4:0]; // @[Modules.scala 150:103:@13046.4]
  assign _T_66573 = $signed(_T_66572); // @[Modules.scala 150:103:@13047.4]
  assign _T_66603 = $signed(-4'sh1) * $signed(io_in_76); // @[Modules.scala 150:74:@13073.4]
  assign _T_66605 = $signed(-4'sh1) * $signed(io_in_77); // @[Modules.scala 151:80:@13074.4]
  assign _T_66606 = $signed(_T_66603) + $signed(_T_66605); // @[Modules.scala 150:103:@13075.4]
  assign _T_66607 = _T_66606[4:0]; // @[Modules.scala 150:103:@13076.4]
  assign _T_66608 = $signed(_T_66607); // @[Modules.scala 150:103:@13077.4]
  assign _T_66610 = $signed(-4'sh1) * $signed(io_in_78); // @[Modules.scala 150:74:@13079.4]
  assign _GEN_282 = {{1{_T_66610[4]}},_T_66610}; // @[Modules.scala 150:103:@13081.4]
  assign _T_66613 = $signed(_GEN_282) + $signed(_T_54346); // @[Modules.scala 150:103:@13081.4]
  assign _T_66614 = _T_66613[5:0]; // @[Modules.scala 150:103:@13082.4]
  assign _T_66615 = $signed(_T_66614); // @[Modules.scala 150:103:@13083.4]
  assign _T_66624 = $signed(4'sh1) * $signed(io_in_86); // @[Modules.scala 150:74:@13091.4]
  assign _GEN_283 = {{1{_T_63499[4]}},_T_63499}; // @[Modules.scala 150:103:@13093.4]
  assign _T_66627 = $signed(_T_66624) + $signed(_GEN_283); // @[Modules.scala 150:103:@13093.4]
  assign _T_66628 = _T_66627[5:0]; // @[Modules.scala 150:103:@13094.4]
  assign _T_66629 = $signed(_T_66628); // @[Modules.scala 150:103:@13095.4]
  assign _GEN_284 = {{1{_T_57423[4]}},_T_57423}; // @[Modules.scala 150:103:@13147.4]
  assign _T_66690 = $signed(_GEN_284) + $signed(_T_54425); // @[Modules.scala 150:103:@13147.4]
  assign _T_66691 = _T_66690[5:0]; // @[Modules.scala 150:103:@13148.4]
  assign _T_66692 = $signed(_T_66691); // @[Modules.scala 150:103:@13149.4]
  assign _T_66697 = $signed(_T_54430) + $signed(_GEN_84); // @[Modules.scala 150:103:@13153.4]
  assign _T_66698 = _T_66697[5:0]; // @[Modules.scala 150:103:@13154.4]
  assign _T_66699 = $signed(_T_66698); // @[Modules.scala 150:103:@13155.4]
  assign _T_66711 = $signed(_T_54444) + $signed(_T_57449); // @[Modules.scala 150:103:@13165.4]
  assign _T_66712 = _T_66711[5:0]; // @[Modules.scala 150:103:@13166.4]
  assign _T_66713 = $signed(_T_66712); // @[Modules.scala 150:103:@13167.4]
  assign _T_66718 = $signed(_T_57451) + $signed(_T_54451); // @[Modules.scala 150:103:@13171.4]
  assign _T_66719 = _T_66718[5:0]; // @[Modules.scala 150:103:@13172.4]
  assign _T_66720 = $signed(_T_66719); // @[Modules.scala 150:103:@13173.4]
  assign _T_66725 = $signed(_T_54453) + $signed(_T_54458); // @[Modules.scala 150:103:@13177.4]
  assign _T_66726 = _T_66725[4:0]; // @[Modules.scala 150:103:@13178.4]
  assign _T_66727 = $signed(_T_66726); // @[Modules.scala 150:103:@13179.4]
  assign _T_66732 = $signed(_T_63599) + $signed(_T_63604); // @[Modules.scala 150:103:@13183.4]
  assign _T_66733 = _T_66732[4:0]; // @[Modules.scala 150:103:@13184.4]
  assign _T_66734 = $signed(_T_66733); // @[Modules.scala 150:103:@13185.4]
  assign _T_66739 = $signed(_T_63606) + $signed(_T_60495); // @[Modules.scala 150:103:@13189.4]
  assign _T_66740 = _T_66739[4:0]; // @[Modules.scala 150:103:@13190.4]
  assign _T_66741 = $signed(_T_66740); // @[Modules.scala 150:103:@13191.4]
  assign _T_66750 = $signed(-4'sh1) * $signed(io_in_129); // @[Modules.scala 150:74:@13199.4]
  assign _GEN_287 = {{1{_T_66750[4]}},_T_66750}; // @[Modules.scala 150:103:@13201.4]
  assign _T_66753 = $signed(_GEN_287) + $signed(_T_54495); // @[Modules.scala 150:103:@13201.4]
  assign _T_66754 = _T_66753[5:0]; // @[Modules.scala 150:103:@13202.4]
  assign _T_66755 = $signed(_T_66754); // @[Modules.scala 150:103:@13203.4]
  assign _GEN_288 = {{1{_T_54507[4]}},_T_54507}; // @[Modules.scala 150:103:@13213.4]
  assign _T_66767 = $signed(_T_54502) + $signed(_GEN_288); // @[Modules.scala 150:103:@13213.4]
  assign _T_66768 = _T_66767[5:0]; // @[Modules.scala 150:103:@13214.4]
  assign _T_66769 = $signed(_T_66768); // @[Modules.scala 150:103:@13215.4]
  assign _T_66774 = $signed(_T_54509) + $signed(_T_54514); // @[Modules.scala 150:103:@13219.4]
  assign _T_66775 = _T_66774[4:0]; // @[Modules.scala 150:103:@13220.4]
  assign _T_66776 = $signed(_T_66775); // @[Modules.scala 150:103:@13221.4]
  assign _T_66781 = $signed(_GEN_152) + $signed(_T_60549); // @[Modules.scala 150:103:@13225.4]
  assign _T_66782 = _T_66781[5:0]; // @[Modules.scala 150:103:@13226.4]
  assign _T_66783 = $signed(_T_66782); // @[Modules.scala 150:103:@13227.4]
  assign _GEN_290 = {{1{_T_63669[4]}},_T_63669}; // @[Modules.scala 150:103:@13231.4]
  assign _T_66788 = $signed(_T_57526) + $signed(_GEN_290); // @[Modules.scala 150:103:@13231.4]
  assign _T_66789 = _T_66788[5:0]; // @[Modules.scala 150:103:@13232.4]
  assign _T_66790 = $signed(_T_66789); // @[Modules.scala 150:103:@13233.4]
  assign _T_66823 = $signed(_T_60586) + $signed(_T_57561); // @[Modules.scala 150:103:@13261.4]
  assign _T_66824 = _T_66823[4:0]; // @[Modules.scala 150:103:@13262.4]
  assign _T_66825 = $signed(_T_66824); // @[Modules.scala 150:103:@13263.4]
  assign _T_66841 = $signed(-4'sh1) * $signed(io_in_159); // @[Modules.scala 150:74:@13277.4]
  assign _T_66844 = $signed(_T_66841) + $signed(_T_54551); // @[Modules.scala 150:103:@13279.4]
  assign _T_66845 = _T_66844[4:0]; // @[Modules.scala 150:103:@13280.4]
  assign _T_66846 = $signed(_T_66845); // @[Modules.scala 150:103:@13281.4]
  assign _T_66851 = $signed(_T_60607) + $signed(_T_54558); // @[Modules.scala 150:103:@13285.4]
  assign _T_66852 = _T_66851[4:0]; // @[Modules.scala 150:103:@13286.4]
  assign _T_66853 = $signed(_T_66852); // @[Modules.scala 150:103:@13287.4]
  assign _T_66865 = $signed(_T_54570) + $signed(_T_57596); // @[Modules.scala 150:103:@13297.4]
  assign _T_66866 = _T_66865[4:0]; // @[Modules.scala 150:103:@13298.4]
  assign _T_66867 = $signed(_T_66866); // @[Modules.scala 150:103:@13299.4]
  assign _T_66872 = $signed(_T_54577) + $signed(_GEN_13); // @[Modules.scala 150:103:@13303.4]
  assign _T_66873 = _T_66872[5:0]; // @[Modules.scala 150:103:@13304.4]
  assign _T_66874 = $signed(_T_66873); // @[Modules.scala 150:103:@13305.4]
  assign _T_66879 = $signed(_GEN_159) + $signed(_T_54591); // @[Modules.scala 150:103:@13309.4]
  assign _T_66880 = _T_66879[5:0]; // @[Modules.scala 150:103:@13310.4]
  assign _T_66881 = $signed(_T_66880); // @[Modules.scala 150:103:@13311.4]
  assign _T_66907 = $signed(_T_60656) + $signed(_T_54612); // @[Modules.scala 150:103:@13333.4]
  assign _T_66908 = _T_66907[4:0]; // @[Modules.scala 150:103:@13334.4]
  assign _T_66909 = $signed(_T_66908); // @[Modules.scala 150:103:@13335.4]
  assign _T_66914 = $signed(_T_57633) + $signed(_T_57638); // @[Modules.scala 150:103:@13339.4]
  assign _T_66915 = _T_66914[5:0]; // @[Modules.scala 150:103:@13340.4]
  assign _T_66916 = $signed(_T_66915); // @[Modules.scala 150:103:@13341.4]
  assign _T_66920 = $signed(4'sh1) * $signed(io_in_185); // @[Modules.scala 151:80:@13344.4]
  assign _T_66921 = $signed(_T_57640) + $signed(_T_66920); // @[Modules.scala 150:103:@13345.4]
  assign _T_66922 = _T_66921[5:0]; // @[Modules.scala 150:103:@13346.4]
  assign _T_66923 = $signed(_T_66922); // @[Modules.scala 150:103:@13347.4]
  assign _T_66925 = $signed(4'sh1) * $signed(io_in_186); // @[Modules.scala 150:74:@13349.4]
  assign _GEN_293 = {{1{_T_60691[4]}},_T_60691}; // @[Modules.scala 150:103:@13351.4]
  assign _T_66928 = $signed(_T_66925) + $signed(_GEN_293); // @[Modules.scala 150:103:@13351.4]
  assign _T_66929 = _T_66928[5:0]; // @[Modules.scala 150:103:@13352.4]
  assign _T_66930 = $signed(_T_66929); // @[Modules.scala 150:103:@13353.4]
  assign _T_66977 = $signed(_T_57701) + $signed(_T_60740); // @[Modules.scala 150:103:@13393.4]
  assign _T_66978 = _T_66977[4:0]; // @[Modules.scala 150:103:@13394.4]
  assign _T_66979 = $signed(_T_66978); // @[Modules.scala 150:103:@13395.4]
  assign _T_66984 = $signed(_T_57710) + $signed(_T_57715); // @[Modules.scala 150:103:@13399.4]
  assign _T_66985 = _T_66984[5:0]; // @[Modules.scala 150:103:@13400.4]
  assign _T_66986 = $signed(_T_66985); // @[Modules.scala 150:103:@13401.4]
  assign _T_66991 = $signed(_T_57717) + $signed(_T_57722); // @[Modules.scala 150:103:@13405.4]
  assign _T_66992 = _T_66991[5:0]; // @[Modules.scala 150:103:@13406.4]
  assign _T_66993 = $signed(_T_66992); // @[Modules.scala 150:103:@13407.4]
  assign _GEN_295 = {{1{_T_54705[4]}},_T_54705}; // @[Modules.scala 150:103:@13417.4]
  assign _T_67005 = $signed(_T_57738) + $signed(_GEN_295); // @[Modules.scala 150:103:@13417.4]
  assign _T_67006 = _T_67005[5:0]; // @[Modules.scala 150:103:@13418.4]
  assign _T_67007 = $signed(_T_67006); // @[Modules.scala 150:103:@13419.4]
  assign _GEN_296 = {{1{_T_57757[4]}},_T_57757}; // @[Modules.scala 150:103:@13435.4]
  assign _T_67026 = $signed(_GEN_296) + $signed(_T_54724); // @[Modules.scala 150:103:@13435.4]
  assign _T_67027 = _T_67026[5:0]; // @[Modules.scala 150:103:@13436.4]
  assign _T_67028 = $signed(_T_67027); // @[Modules.scala 150:103:@13437.4]
  assign _T_67033 = $signed(_T_57764) + $signed(_T_54738); // @[Modules.scala 150:103:@13441.4]
  assign _T_67034 = _T_67033[5:0]; // @[Modules.scala 150:103:@13442.4]
  assign _T_67035 = $signed(_T_67034); // @[Modules.scala 150:103:@13443.4]
  assign _GEN_297 = {{1{_T_60822[4]}},_T_60822}; // @[Modules.scala 150:103:@13447.4]
  assign _T_67040 = $signed(_T_54740) + $signed(_GEN_297); // @[Modules.scala 150:103:@13447.4]
  assign _T_67041 = _T_67040[5:0]; // @[Modules.scala 150:103:@13448.4]
  assign _T_67042 = $signed(_T_67041); // @[Modules.scala 150:103:@13449.4]
  assign _T_67053 = $signed(4'sh1) * $signed(io_in_236); // @[Modules.scala 151:80:@13458.4]
  assign _GEN_298 = {{1{_T_60831[4]}},_T_60831}; // @[Modules.scala 150:103:@13459.4]
  assign _T_67054 = $signed(_GEN_298) + $signed(_T_67053); // @[Modules.scala 150:103:@13459.4]
  assign _T_67055 = _T_67054[5:0]; // @[Modules.scala 150:103:@13460.4]
  assign _T_67056 = $signed(_T_67055); // @[Modules.scala 150:103:@13461.4]
  assign _GEN_299 = {{1{_T_54780[4]}},_T_54780}; // @[Modules.scala 150:103:@13477.4]
  assign _T_67075 = $signed(_T_57813) + $signed(_GEN_299); // @[Modules.scala 150:103:@13477.4]
  assign _T_67076 = _T_67075[5:0]; // @[Modules.scala 150:103:@13478.4]
  assign _T_67077 = $signed(_T_67076); // @[Modules.scala 150:103:@13479.4]
  assign _T_67110 = $signed(_T_57850) + $signed(_T_54815); // @[Modules.scala 150:103:@13507.4]
  assign _T_67111 = _T_67110[5:0]; // @[Modules.scala 150:103:@13508.4]
  assign _T_67112 = $signed(_T_67111); // @[Modules.scala 150:103:@13509.4]
  assign _GEN_300 = {{1{_T_60906[4]}},_T_60906}; // @[Modules.scala 150:103:@13513.4]
  assign _T_67117 = $signed(_T_57857) + $signed(_GEN_300); // @[Modules.scala 150:103:@13513.4]
  assign _T_67118 = _T_67117[5:0]; // @[Modules.scala 150:103:@13514.4]
  assign _T_67119 = $signed(_T_67118); // @[Modules.scala 150:103:@13515.4]
  assign _T_67124 = $signed(_T_60913) + $signed(_T_54831); // @[Modules.scala 150:103:@13519.4]
  assign _T_67125 = _T_67124[4:0]; // @[Modules.scala 150:103:@13520.4]
  assign _T_67126 = $signed(_T_67125); // @[Modules.scala 150:103:@13521.4]
  assign _T_67130 = $signed(4'sh1) * $signed(io_in_264); // @[Modules.scala 151:80:@13524.4]
  assign _T_67131 = $signed(_T_64026) + $signed(_T_67130); // @[Modules.scala 150:103:@13525.4]
  assign _T_67132 = _T_67131[5:0]; // @[Modules.scala 150:103:@13526.4]
  assign _T_67133 = $signed(_T_67132); // @[Modules.scala 150:103:@13527.4]
  assign _T_67135 = $signed(4'sh1) * $signed(io_in_265); // @[Modules.scala 150:74:@13529.4]
  assign _T_67138 = $signed(_T_67135) + $signed(_T_54845); // @[Modules.scala 150:103:@13531.4]
  assign _T_67139 = _T_67138[5:0]; // @[Modules.scala 150:103:@13532.4]
  assign _T_67140 = $signed(_T_67139); // @[Modules.scala 150:103:@13533.4]
  assign _T_67145 = $signed(_T_54850) + $signed(_T_57890); // @[Modules.scala 150:103:@13537.4]
  assign _T_67146 = _T_67145[5:0]; // @[Modules.scala 150:103:@13538.4]
  assign _T_67147 = $signed(_T_67146); // @[Modules.scala 150:103:@13539.4]
  assign _T_67152 = $signed(_T_57892) + $signed(_T_57897); // @[Modules.scala 150:103:@13543.4]
  assign _T_67153 = _T_67152[5:0]; // @[Modules.scala 150:103:@13544.4]
  assign _T_67154 = $signed(_T_67153); // @[Modules.scala 150:103:@13545.4]
  assign _T_67187 = $signed(_T_57927) + $signed(_T_54899); // @[Modules.scala 150:103:@13573.4]
  assign _T_67188 = _T_67187[5:0]; // @[Modules.scala 150:103:@13574.4]
  assign _T_67189 = $signed(_T_67188); // @[Modules.scala 150:103:@13575.4]
  assign _T_67200 = $signed(4'sh1) * $signed(io_in_285); // @[Modules.scala 151:80:@13584.4]
  assign _T_67201 = $signed(_GEN_24) + $signed(_T_67200); // @[Modules.scala 150:103:@13585.4]
  assign _T_67202 = _T_67201[5:0]; // @[Modules.scala 150:103:@13586.4]
  assign _T_67203 = $signed(_T_67202); // @[Modules.scala 150:103:@13587.4]
  assign _GEN_302 = {{1{_T_54927[4]}},_T_54927}; // @[Modules.scala 150:103:@13591.4]
  assign _T_67208 = $signed(_T_61004) + $signed(_GEN_302); // @[Modules.scala 150:103:@13591.4]
  assign _T_67209 = _T_67208[5:0]; // @[Modules.scala 150:103:@13592.4]
  assign _T_67210 = $signed(_T_67209); // @[Modules.scala 150:103:@13593.4]
  assign _T_67215 = $signed(_T_64122) + $signed(_GEN_99); // @[Modules.scala 150:103:@13597.4]
  assign _T_67216 = _T_67215[5:0]; // @[Modules.scala 150:103:@13598.4]
  assign _T_67217 = $signed(_T_67216); // @[Modules.scala 150:103:@13599.4]
  assign _T_67222 = $signed(_T_57962) + $signed(_T_54943); // @[Modules.scala 150:103:@13603.4]
  assign _T_67223 = _T_67222[5:0]; // @[Modules.scala 150:103:@13604.4]
  assign _T_67224 = $signed(_T_67223); // @[Modules.scala 150:103:@13605.4]
  assign _T_67247 = $signed(4'sh1) * $signed(io_in_302); // @[Modules.scala 150:74:@13625.4]
  assign _GEN_304 = {{1{_T_54971[4]}},_T_54971}; // @[Modules.scala 150:103:@13627.4]
  assign _T_67250 = $signed(_T_67247) + $signed(_GEN_304); // @[Modules.scala 150:103:@13627.4]
  assign _T_67251 = _T_67250[5:0]; // @[Modules.scala 150:103:@13628.4]
  assign _T_67252 = $signed(_T_67251); // @[Modules.scala 150:103:@13629.4]
  assign _T_67264 = $signed(_T_54983) + $signed(_T_64173); // @[Modules.scala 150:103:@13639.4]
  assign _T_67265 = _T_67264[4:0]; // @[Modules.scala 150:103:@13640.4]
  assign _T_67266 = $signed(_T_67265); // @[Modules.scala 150:103:@13641.4]
  assign _T_67271 = $signed(_T_58011) + $signed(_T_54990); // @[Modules.scala 150:103:@13645.4]
  assign _T_67272 = _T_67271[5:0]; // @[Modules.scala 150:103:@13646.4]
  assign _T_67273 = $signed(_T_67272); // @[Modules.scala 150:103:@13647.4]
  assign _T_67278 = $signed(_T_58018) + $signed(_T_58025); // @[Modules.scala 150:103:@13651.4]
  assign _T_67279 = _T_67278[5:0]; // @[Modules.scala 150:103:@13652.4]
  assign _T_67280 = $signed(_T_67279); // @[Modules.scala 150:103:@13653.4]
  assign _T_67285 = $signed(_T_64194) + $signed(_T_58032); // @[Modules.scala 150:103:@13657.4]
  assign _T_67286 = _T_67285[5:0]; // @[Modules.scala 150:103:@13658.4]
  assign _T_67287 = $signed(_T_67286); // @[Modules.scala 150:103:@13659.4]
  assign _T_67299 = $signed(_GEN_101) + $signed(_T_58058); // @[Modules.scala 150:103:@13669.4]
  assign _T_67300 = _T_67299[5:0]; // @[Modules.scala 150:103:@13670.4]
  assign _T_67301 = $signed(_T_67300); // @[Modules.scala 150:103:@13671.4]
  assign _T_67306 = $signed(_T_55034) + $signed(_T_58065); // @[Modules.scala 150:103:@13675.4]
  assign _T_67307 = _T_67306[5:0]; // @[Modules.scala 150:103:@13676.4]
  assign _T_67308 = $signed(_T_67307); // @[Modules.scala 150:103:@13677.4]
  assign _GEN_306 = {{1{_T_55041[4]}},_T_55041}; // @[Modules.scala 150:103:@13681.4]
  assign _T_67313 = $signed(_GEN_306) + $signed(_T_58074); // @[Modules.scala 150:103:@13681.4]
  assign _T_67314 = _T_67313[5:0]; // @[Modules.scala 150:103:@13682.4]
  assign _T_67315 = $signed(_T_67314); // @[Modules.scala 150:103:@13683.4]
  assign _T_67324 = $signed(4'sh1) * $signed(io_in_330); // @[Modules.scala 150:74:@13691.4]
  assign _GEN_307 = {{1{_T_55062[4]}},_T_55062}; // @[Modules.scala 150:103:@13693.4]
  assign _T_67327 = $signed(_T_67324) + $signed(_GEN_307); // @[Modules.scala 150:103:@13693.4]
  assign _T_67328 = _T_67327[5:0]; // @[Modules.scala 150:103:@13694.4]
  assign _T_67329 = $signed(_T_67328); // @[Modules.scala 150:103:@13695.4]
  assign _T_67340 = $signed(-4'sh1) * $signed(io_in_335); // @[Modules.scala 151:80:@13704.4]
  assign _T_67341 = $signed(_T_58095) + $signed(_T_67340); // @[Modules.scala 150:103:@13705.4]
  assign _T_67342 = _T_67341[4:0]; // @[Modules.scala 150:103:@13706.4]
  assign _T_67343 = $signed(_T_67342); // @[Modules.scala 150:103:@13707.4]
  assign _GEN_308 = {{1{_T_58109[4]}},_T_58109}; // @[Modules.scala 150:103:@13711.4]
  assign _T_67348 = $signed(_T_55076) + $signed(_GEN_308); // @[Modules.scala 150:103:@13711.4]
  assign _T_67349 = _T_67348[5:0]; // @[Modules.scala 150:103:@13712.4]
  assign _T_67350 = $signed(_T_67349); // @[Modules.scala 150:103:@13713.4]
  assign _GEN_309 = {{1{_T_55109[4]}},_T_55109}; // @[Modules.scala 150:103:@13729.4]
  assign _T_67369 = $signed(_T_61167) + $signed(_GEN_309); // @[Modules.scala 150:103:@13729.4]
  assign _T_67370 = _T_67369[5:0]; // @[Modules.scala 150:103:@13730.4]
  assign _T_67371 = $signed(_T_67370); // @[Modules.scala 150:103:@13731.4]
  assign _GEN_310 = {{1{_T_55118[4]}},_T_55118}; // @[Modules.scala 150:103:@13741.4]
  assign _T_67383 = $signed(_GEN_310) + $signed(_T_55123); // @[Modules.scala 150:103:@13741.4]
  assign _T_67384 = _T_67383[5:0]; // @[Modules.scala 150:103:@13742.4]
  assign _T_67385 = $signed(_T_67384); // @[Modules.scala 150:103:@13743.4]
  assign _GEN_311 = {{1{_T_55130[4]}},_T_55130}; // @[Modules.scala 150:103:@13747.4]
  assign _T_67390 = $signed(_T_55125) + $signed(_GEN_311); // @[Modules.scala 150:103:@13747.4]
  assign _T_67391 = _T_67390[5:0]; // @[Modules.scala 150:103:@13748.4]
  assign _T_67392 = $signed(_T_67391); // @[Modules.scala 150:103:@13749.4]
  assign _GEN_312 = {{1{_T_55132[4]}},_T_55132}; // @[Modules.scala 150:103:@13753.4]
  assign _T_67397 = $signed(_GEN_312) + $signed(_T_58158); // @[Modules.scala 150:103:@13753.4]
  assign _T_67398 = _T_67397[5:0]; // @[Modules.scala 150:103:@13754.4]
  assign _T_67399 = $signed(_T_67398); // @[Modules.scala 150:103:@13755.4]
  assign _T_67411 = $signed(_T_58170) + $signed(_T_61214); // @[Modules.scala 150:103:@13765.4]
  assign _T_67412 = _T_67411[5:0]; // @[Modules.scala 150:103:@13766.4]
  assign _T_67413 = $signed(_T_67412); // @[Modules.scala 150:103:@13767.4]
  assign _T_67425 = $signed(_T_55153) + $signed(_T_55158); // @[Modules.scala 150:103:@13777.4]
  assign _T_67426 = _T_67425[4:0]; // @[Modules.scala 150:103:@13778.4]
  assign _T_67427 = $signed(_T_67426); // @[Modules.scala 150:103:@13779.4]
  assign _GEN_314 = {{1{_T_58193[4]}},_T_58193}; // @[Modules.scala 150:103:@13789.4]
  assign _T_67439 = $signed(_GEN_314) + $signed(_T_55174); // @[Modules.scala 150:103:@13789.4]
  assign _T_67440 = _T_67439[5:0]; // @[Modules.scala 150:103:@13790.4]
  assign _T_67441 = $signed(_T_67440); // @[Modules.scala 150:103:@13791.4]
  assign _GEN_316 = {{1{_T_55209[4]}},_T_55209}; // @[Modules.scala 150:103:@13813.4]
  assign _T_67467 = $signed(_GEN_316) + $signed(_T_55214); // @[Modules.scala 150:103:@13813.4]
  assign _T_67468 = _T_67467[5:0]; // @[Modules.scala 150:103:@13814.4]
  assign _T_67469 = $signed(_T_67468); // @[Modules.scala 150:103:@13815.4]
  assign _T_67474 = $signed(_T_58233) + $signed(_T_55221); // @[Modules.scala 150:103:@13819.4]
  assign _T_67475 = _T_67474[5:0]; // @[Modules.scala 150:103:@13820.4]
  assign _T_67476 = $signed(_T_67475); // @[Modules.scala 150:103:@13821.4]
  assign _GEN_317 = {{1{_T_58261[4]}},_T_58261}; // @[Modules.scala 150:103:@13831.4]
  assign _T_67488 = $signed(_T_61305) + $signed(_GEN_317); // @[Modules.scala 150:103:@13831.4]
  assign _T_67489 = _T_67488[5:0]; // @[Modules.scala 150:103:@13832.4]
  assign _T_67490 = $signed(_T_67489); // @[Modules.scala 150:103:@13833.4]
  assign _T_67502 = $signed(_T_55242) + $signed(_T_61326); // @[Modules.scala 150:103:@13843.4]
  assign _T_67503 = _T_67502[4:0]; // @[Modules.scala 150:103:@13844.4]
  assign _T_67504 = $signed(_T_67503); // @[Modules.scala 150:103:@13845.4]
  assign _T_67509 = $signed(_GEN_106) + $signed(_T_58282); // @[Modules.scala 150:103:@13849.4]
  assign _T_67510 = _T_67509[5:0]; // @[Modules.scala 150:103:@13850.4]
  assign _T_67511 = $signed(_T_67510); // @[Modules.scala 150:103:@13851.4]
  assign _T_67516 = $signed(_GEN_242) + $signed(_T_55258); // @[Modules.scala 150:103:@13855.4]
  assign _T_67517 = _T_67516[5:0]; // @[Modules.scala 150:103:@13856.4]
  assign _T_67518 = $signed(_T_67517); // @[Modules.scala 150:103:@13857.4]
  assign _T_67550 = $signed(-4'sh1) * $signed(io_in_405); // @[Modules.scala 151:80:@13884.4]
  assign _T_67551 = $signed(_T_55291) + $signed(_T_67550); // @[Modules.scala 150:103:@13885.4]
  assign _T_67552 = _T_67551[4:0]; // @[Modules.scala 150:103:@13886.4]
  assign _T_67553 = $signed(_T_67552); // @[Modules.scala 150:103:@13887.4]
  assign _T_67565 = $signed(_T_55307) + $signed(_T_55312); // @[Modules.scala 150:103:@13897.4]
  assign _T_67566 = _T_67565[5:0]; // @[Modules.scala 150:103:@13898.4]
  assign _T_67567 = $signed(_T_67566); // @[Modules.scala 150:103:@13899.4]
  assign _T_67585 = $signed(4'sh1) * $signed(io_in_419); // @[Modules.scala 151:80:@13914.4]
  assign _T_67586 = $signed(_GEN_42) + $signed(_T_67585); // @[Modules.scala 150:103:@13915.4]
  assign _T_67587 = _T_67586[5:0]; // @[Modules.scala 150:103:@13916.4]
  assign _T_67588 = $signed(_T_67587); // @[Modules.scala 150:103:@13917.4]
  assign _T_67597 = $signed(-4'sh1) * $signed(io_in_422); // @[Modules.scala 150:74:@13925.4]
  assign _GEN_321 = {{1{_T_67597[4]}},_T_67597}; // @[Modules.scala 150:103:@13927.4]
  assign _T_67600 = $signed(_GEN_321) + $signed(_T_58361); // @[Modules.scala 150:103:@13927.4]
  assign _T_67601 = _T_67600[5:0]; // @[Modules.scala 150:103:@13928.4]
  assign _T_67602 = $signed(_T_67601); // @[Modules.scala 150:103:@13929.4]
  assign _T_67614 = $signed(_T_55354) + $signed(_T_55361); // @[Modules.scala 150:103:@13939.4]
  assign _T_67615 = _T_67614[4:0]; // @[Modules.scala 150:103:@13940.4]
  assign _T_67616 = $signed(_T_67615); // @[Modules.scala 150:103:@13941.4]
  assign _T_67621 = $signed(_T_58382) + $signed(_T_58387); // @[Modules.scala 150:103:@13945.4]
  assign _T_67622 = _T_67621[4:0]; // @[Modules.scala 150:103:@13946.4]
  assign _T_67623 = $signed(_T_67622); // @[Modules.scala 150:103:@13947.4]
  assign _T_67628 = $signed(_GEN_177) + $signed(_T_55370); // @[Modules.scala 150:103:@13951.4]
  assign _T_67629 = _T_67628[5:0]; // @[Modules.scala 150:103:@13952.4]
  assign _T_67630 = $signed(_T_67629); // @[Modules.scala 150:103:@13953.4]
  assign _T_67635 = $signed(_T_61468) + $signed(_T_55384); // @[Modules.scala 150:103:@13957.4]
  assign _T_67636 = _T_67635[5:0]; // @[Modules.scala 150:103:@13958.4]
  assign _T_67637 = $signed(_T_67636); // @[Modules.scala 150:103:@13959.4]
  assign _GEN_323 = {{1{_T_64579[4]}},_T_64579}; // @[Modules.scala 150:103:@13963.4]
  assign _T_67642 = $signed(_GEN_323) + $signed(_T_55396); // @[Modules.scala 150:103:@13963.4]
  assign _T_67643 = _T_67642[5:0]; // @[Modules.scala 150:103:@13964.4]
  assign _T_67644 = $signed(_T_67643); // @[Modules.scala 150:103:@13965.4]
  assign _GEN_324 = {{1{_T_61496[4]}},_T_61496}; // @[Modules.scala 150:103:@13981.4]
  assign _T_67663 = $signed(_GEN_324) + $signed(_T_58424); // @[Modules.scala 150:103:@13981.4]
  assign _T_67664 = _T_67663[5:0]; // @[Modules.scala 150:103:@13982.4]
  assign _T_67665 = $signed(_T_67664); // @[Modules.scala 150:103:@13983.4]
  assign _T_67670 = $signed(_T_64614) + $signed(_T_55433); // @[Modules.scala 150:103:@13987.4]
  assign _T_67671 = _T_67670[4:0]; // @[Modules.scala 150:103:@13988.4]
  assign _T_67672 = $signed(_T_67671); // @[Modules.scala 150:103:@13989.4]
  assign _GEN_325 = {{1{_T_58445[4]}},_T_58445}; // @[Modules.scala 150:103:@13993.4]
  assign _T_67677 = $signed(_GEN_325) + $signed(_T_64635); // @[Modules.scala 150:103:@13993.4]
  assign _T_67678 = _T_67677[5:0]; // @[Modules.scala 150:103:@13994.4]
  assign _T_67679 = $signed(_T_67678); // @[Modules.scala 150:103:@13995.4]
  assign _T_67684 = $signed(_T_58459) + $signed(_T_58464); // @[Modules.scala 150:103:@13999.4]
  assign _T_67685 = _T_67684[4:0]; // @[Modules.scala 150:103:@14000.4]
  assign _T_67686 = $signed(_T_67685); // @[Modules.scala 150:103:@14001.4]
  assign _T_67691 = $signed(_T_58466) + $signed(_T_61536); // @[Modules.scala 150:103:@14005.4]
  assign _T_67692 = _T_67691[4:0]; // @[Modules.scala 150:103:@14006.4]
  assign _T_67693 = $signed(_T_67692); // @[Modules.scala 150:103:@14007.4]
  assign _T_67695 = $signed(-4'sh1) * $signed(io_in_462); // @[Modules.scala 150:74:@14009.4]
  assign _T_67698 = $signed(_T_67695) + $signed(_T_58471); // @[Modules.scala 150:103:@14011.4]
  assign _T_67699 = _T_67698[4:0]; // @[Modules.scala 150:103:@14012.4]
  assign _T_67700 = $signed(_T_67699); // @[Modules.scala 150:103:@14013.4]
  assign _T_67705 = $signed(_T_58480) + $signed(_GEN_52); // @[Modules.scala 150:103:@14017.4]
  assign _T_67706 = _T_67705[5:0]; // @[Modules.scala 150:103:@14018.4]
  assign _T_67707 = $signed(_T_67706); // @[Modules.scala 150:103:@14019.4]
  assign _T_67747 = $signed(_T_61606) + $signed(_GEN_54); // @[Modules.scala 150:103:@14053.4]
  assign _T_67748 = _T_67747[5:0]; // @[Modules.scala 150:103:@14054.4]
  assign _T_67749 = $signed(_T_67748); // @[Modules.scala 150:103:@14055.4]
  assign _GEN_330 = {{1{_T_58536[4]}},_T_58536}; // @[Modules.scala 150:103:@14059.4]
  assign _T_67754 = $signed(_GEN_330) + $signed(_T_55517); // @[Modules.scala 150:103:@14059.4]
  assign _T_67755 = _T_67754[5:0]; // @[Modules.scala 150:103:@14060.4]
  assign _T_67756 = $signed(_T_67755); // @[Modules.scala 150:103:@14061.4]
  assign _GEN_331 = {{1{_T_55531[4]}},_T_55531}; // @[Modules.scala 150:103:@14065.4]
  assign _T_67761 = $signed(_T_61622) + $signed(_GEN_331); // @[Modules.scala 150:103:@14065.4]
  assign _T_67762 = _T_67761[5:0]; // @[Modules.scala 150:103:@14066.4]
  assign _T_67763 = $signed(_T_67762); // @[Modules.scala 150:103:@14067.4]
  assign _T_67765 = $signed(4'sh1) * $signed(io_in_495); // @[Modules.scala 150:74:@14069.4]
  assign _T_67767 = $signed(4'sh1) * $signed(io_in_496); // @[Modules.scala 151:80:@14070.4]
  assign _T_67768 = $signed(_T_67765) + $signed(_T_67767); // @[Modules.scala 150:103:@14071.4]
  assign _T_67769 = _T_67768[5:0]; // @[Modules.scala 150:103:@14072.4]
  assign _T_67770 = $signed(_T_67769); // @[Modules.scala 150:103:@14073.4]
  assign _T_67775 = $signed(_T_55538) + $signed(_GEN_186); // @[Modules.scala 150:103:@14077.4]
  assign _T_67776 = _T_67775[5:0]; // @[Modules.scala 150:103:@14078.4]
  assign _T_67777 = $signed(_T_67776); // @[Modules.scala 150:103:@14079.4]
  assign _T_67796 = $signed(_T_55557) + $signed(_T_58590); // @[Modules.scala 150:103:@14095.4]
  assign _T_67797 = _T_67796[5:0]; // @[Modules.scala 150:103:@14096.4]
  assign _T_67798 = $signed(_T_67797); // @[Modules.scala 150:103:@14097.4]
  assign _T_67817 = $signed(_T_58599) + $signed(_T_55580); // @[Modules.scala 150:103:@14113.4]
  assign _T_67818 = _T_67817[4:0]; // @[Modules.scala 150:103:@14114.4]
  assign _T_67819 = $signed(_T_67818); // @[Modules.scala 150:103:@14115.4]
  assign _T_67824 = $signed(_T_58606) + $signed(_T_55585); // @[Modules.scala 150:103:@14119.4]
  assign _T_67825 = _T_67824[4:0]; // @[Modules.scala 150:103:@14120.4]
  assign _T_67826 = $signed(_T_67825); // @[Modules.scala 150:103:@14121.4]
  assign _T_67831 = $signed(_T_58613) + $signed(_T_58618); // @[Modules.scala 150:103:@14125.4]
  assign _T_67832 = _T_67831[4:0]; // @[Modules.scala 150:103:@14126.4]
  assign _T_67833 = $signed(_T_67832); // @[Modules.scala 150:103:@14127.4]
  assign _T_67845 = $signed(_T_55606) + $signed(_GEN_256); // @[Modules.scala 150:103:@14137.4]
  assign _T_67846 = _T_67845[5:0]; // @[Modules.scala 150:103:@14138.4]
  assign _T_67847 = $signed(_T_67846); // @[Modules.scala 150:103:@14139.4]
  assign _GEN_335 = {{1{_T_64871[4]}},_T_64871}; // @[Modules.scala 150:103:@14161.4]
  assign _T_67873 = $signed(_T_58655) + $signed(_GEN_335); // @[Modules.scala 150:103:@14161.4]
  assign _T_67874 = _T_67873[5:0]; // @[Modules.scala 150:103:@14162.4]
  assign _T_67875 = $signed(_T_67874); // @[Modules.scala 150:103:@14163.4]
  assign _T_67901 = $signed(_T_58683) + $signed(_T_58688); // @[Modules.scala 150:103:@14185.4]
  assign _T_67902 = _T_67901[4:0]; // @[Modules.scala 150:103:@14186.4]
  assign _T_67903 = $signed(_T_67902); // @[Modules.scala 150:103:@14187.4]
  assign _GEN_336 = {{1{_T_58690[4]}},_T_58690}; // @[Modules.scala 150:103:@14191.4]
  assign _T_67908 = $signed(_GEN_336) + $signed(_T_55690); // @[Modules.scala 150:103:@14191.4]
  assign _T_67909 = _T_67908[5:0]; // @[Modules.scala 150:103:@14192.4]
  assign _T_67910 = $signed(_T_67909); // @[Modules.scala 150:103:@14193.4]
  assign _T_67928 = $signed(-4'sh1) * $signed(io_in_552); // @[Modules.scala 151:80:@14208.4]
  assign _T_67929 = $signed(_T_64920) + $signed(_T_67928); // @[Modules.scala 150:103:@14209.4]
  assign _T_67930 = _T_67929[4:0]; // @[Modules.scala 150:103:@14210.4]
  assign _T_67931 = $signed(_T_67930); // @[Modules.scala 150:103:@14211.4]
  assign _T_67943 = $signed(_T_58725) + $signed(_T_58730); // @[Modules.scala 150:103:@14221.4]
  assign _T_67944 = _T_67943[4:0]; // @[Modules.scala 150:103:@14222.4]
  assign _T_67945 = $signed(_T_67944); // @[Modules.scala 150:103:@14223.4]
  assign _T_67950 = $signed(_GEN_260) + $signed(_T_55720); // @[Modules.scala 150:103:@14227.4]
  assign _T_67951 = _T_67950[5:0]; // @[Modules.scala 150:103:@14228.4]
  assign _T_67952 = $signed(_T_67951); // @[Modules.scala 150:103:@14229.4]
  assign _GEN_338 = {{1{_T_64950[4]}},_T_64950}; // @[Modules.scala 150:103:@14233.4]
  assign _T_67957 = $signed(_T_64943) + $signed(_GEN_338); // @[Modules.scala 150:103:@14233.4]
  assign _T_67958 = _T_67957[5:0]; // @[Modules.scala 150:103:@14234.4]
  assign _T_67959 = $signed(_T_67958); // @[Modules.scala 150:103:@14235.4]
  assign _T_67991 = $signed(-4'sh1) * $signed(io_in_575); // @[Modules.scala 151:80:@14262.4]
  assign _GEN_339 = {{1{_T_67991[4]}},_T_67991}; // @[Modules.scala 150:103:@14263.4]
  assign _T_67992 = $signed(_T_55755) + $signed(_GEN_339); // @[Modules.scala 150:103:@14263.4]
  assign _T_67993 = _T_67992[5:0]; // @[Modules.scala 150:103:@14264.4]
  assign _T_67994 = $signed(_T_67993); // @[Modules.scala 150:103:@14265.4]
  assign _T_67999 = $signed(_T_58774) + $signed(_T_58781); // @[Modules.scala 150:103:@14269.4]
  assign _T_68000 = _T_67999[4:0]; // @[Modules.scala 150:103:@14270.4]
  assign _T_68001 = $signed(_T_68000); // @[Modules.scala 150:103:@14271.4]
  assign _T_68006 = $signed(_T_61858) + $signed(_T_55769); // @[Modules.scala 150:103:@14275.4]
  assign _T_68007 = _T_68006[4:0]; // @[Modules.scala 150:103:@14276.4]
  assign _T_68008 = $signed(_T_68007); // @[Modules.scala 150:103:@14277.4]
  assign _GEN_340 = {{1{_T_58800[4]}},_T_58800}; // @[Modules.scala 150:103:@14287.4]
  assign _T_68020 = $signed(_GEN_340) + $signed(_T_55781); // @[Modules.scala 150:103:@14287.4]
  assign _T_68021 = _T_68020[5:0]; // @[Modules.scala 150:103:@14288.4]
  assign _T_68022 = $signed(_T_68021); // @[Modules.scala 150:103:@14289.4]
  assign _GEN_341 = {{1{_T_58814[4]}},_T_58814}; // @[Modules.scala 150:103:@14293.4]
  assign _T_68027 = $signed(_T_58809) + $signed(_GEN_341); // @[Modules.scala 150:103:@14293.4]
  assign _T_68028 = _T_68027[5:0]; // @[Modules.scala 150:103:@14294.4]
  assign _T_68029 = $signed(_T_68028); // @[Modules.scala 150:103:@14295.4]
  assign _GEN_342 = {{1{_T_58816[4]}},_T_58816}; // @[Modules.scala 150:103:@14299.4]
  assign _T_68034 = $signed(_GEN_342) + $signed(_T_55795); // @[Modules.scala 150:103:@14299.4]
  assign _T_68035 = _T_68034[5:0]; // @[Modules.scala 150:103:@14300.4]
  assign _T_68036 = $signed(_T_68035); // @[Modules.scala 150:103:@14301.4]
  assign _T_68038 = $signed(-4'sh1) * $signed(io_in_590); // @[Modules.scala 150:74:@14303.4]
  assign _T_68041 = $signed(_T_68038) + $signed(_T_61895); // @[Modules.scala 150:103:@14305.4]
  assign _T_68042 = _T_68041[4:0]; // @[Modules.scala 150:103:@14306.4]
  assign _T_68043 = $signed(_T_68042); // @[Modules.scala 150:103:@14307.4]
  assign _T_68069 = $signed(_T_55823) + $signed(_GEN_126); // @[Modules.scala 150:103:@14329.4]
  assign _T_68070 = _T_68069[5:0]; // @[Modules.scala 150:103:@14330.4]
  assign _T_68071 = $signed(_T_68070); // @[Modules.scala 150:103:@14331.4]
  assign _T_68075 = $signed(-4'sh1) * $signed(io_in_603); // @[Modules.scala 151:80:@14334.4]
  assign _T_68076 = $signed(_T_58849) + $signed(_T_68075); // @[Modules.scala 150:103:@14335.4]
  assign _T_68077 = _T_68076[4:0]; // @[Modules.scala 150:103:@14336.4]
  assign _T_68078 = $signed(_T_68077); // @[Modules.scala 150:103:@14337.4]
  assign _T_68083 = $signed(_T_65048) + $signed(_T_58856); // @[Modules.scala 150:103:@14341.4]
  assign _T_68084 = _T_68083[4:0]; // @[Modules.scala 150:103:@14342.4]
  assign _T_68085 = $signed(_T_68084); // @[Modules.scala 150:103:@14343.4]
  assign _T_68090 = $signed(_T_61944) + $signed(_T_58865); // @[Modules.scala 150:103:@14347.4]
  assign _T_68091 = _T_68090[4:0]; // @[Modules.scala 150:103:@14348.4]
  assign _T_68092 = $signed(_T_68091); // @[Modules.scala 150:103:@14349.4]
  assign _T_68111 = $signed(_T_65074) + $signed(_T_58886); // @[Modules.scala 150:103:@14365.4]
  assign _T_68112 = _T_68111[4:0]; // @[Modules.scala 150:103:@14366.4]
  assign _T_68113 = $signed(_T_68112); // @[Modules.scala 150:103:@14367.4]
  assign _T_68118 = $signed(_T_58891) + $signed(_T_65083); // @[Modules.scala 150:103:@14371.4]
  assign _T_68119 = _T_68118[4:0]; // @[Modules.scala 150:103:@14372.4]
  assign _T_68120 = $signed(_T_68119); // @[Modules.scala 150:103:@14373.4]
  assign _T_68153 = $signed(_T_55895) + $signed(_T_55900); // @[Modules.scala 150:103:@14401.4]
  assign _T_68154 = _T_68153[4:0]; // @[Modules.scala 150:103:@14402.4]
  assign _T_68155 = $signed(_T_68154); // @[Modules.scala 150:103:@14403.4]
  assign _T_68171 = $signed(-4'sh1) * $signed(io_in_635); // @[Modules.scala 150:74:@14417.4]
  assign _T_68174 = $signed(_T_68171) + $signed(_T_58940); // @[Modules.scala 150:103:@14419.4]
  assign _T_68175 = _T_68174[4:0]; // @[Modules.scala 150:103:@14420.4]
  assign _T_68176 = $signed(_T_68175); // @[Modules.scala 150:103:@14421.4]
  assign _T_68181 = $signed(_T_58942) + $signed(_T_58947); // @[Modules.scala 150:103:@14425.4]
  assign _T_68182 = _T_68181[4:0]; // @[Modules.scala 150:103:@14426.4]
  assign _T_68183 = $signed(_T_68182); // @[Modules.scala 150:103:@14427.4]
  assign _GEN_344 = {{1{_T_65160[4]}},_T_65160}; // @[Modules.scala 150:103:@14431.4]
  assign _T_68188 = $signed(_T_55937) + $signed(_GEN_344); // @[Modules.scala 150:103:@14431.4]
  assign _T_68189 = _T_68188[5:0]; // @[Modules.scala 150:103:@14432.4]
  assign _T_68190 = $signed(_T_68189); // @[Modules.scala 150:103:@14433.4]
  assign _T_68194 = $signed(-4'sh1) * $signed(io_in_646); // @[Modules.scala 151:80:@14436.4]
  assign _GEN_345 = {{1{_T_68194[4]}},_T_68194}; // @[Modules.scala 150:103:@14437.4]
  assign _T_68195 = $signed(_T_55944) + $signed(_GEN_345); // @[Modules.scala 150:103:@14437.4]
  assign _T_68196 = _T_68195[5:0]; // @[Modules.scala 150:103:@14438.4]
  assign _T_68197 = $signed(_T_68196); // @[Modules.scala 150:103:@14439.4]
  assign _T_68202 = $signed(_T_62049) + $signed(_T_62054); // @[Modules.scala 150:103:@14443.4]
  assign _T_68203 = _T_68202[4:0]; // @[Modules.scala 150:103:@14444.4]
  assign _T_68204 = $signed(_T_68203); // @[Modules.scala 150:103:@14445.4]
  assign _T_68209 = $signed(_T_62056) + $signed(_T_62061); // @[Modules.scala 150:103:@14449.4]
  assign _T_68210 = _T_68209[4:0]; // @[Modules.scala 150:103:@14450.4]
  assign _T_68211 = $signed(_T_68210); // @[Modules.scala 150:103:@14451.4]
  assign _GEN_346 = {{1{_T_62063[4]}},_T_62063}; // @[Modules.scala 150:103:@14455.4]
  assign _T_68216 = $signed(_GEN_346) + $signed(_T_58982); // @[Modules.scala 150:103:@14455.4]
  assign _T_68217 = _T_68216[5:0]; // @[Modules.scala 150:103:@14456.4]
  assign _T_68218 = $signed(_T_68217); // @[Modules.scala 150:103:@14457.4]
  assign _T_68220 = $signed(4'sh1) * $signed(io_in_654); // @[Modules.scala 150:74:@14459.4]
  assign _GEN_347 = {{1{_T_55979[4]}},_T_55979}; // @[Modules.scala 150:103:@14461.4]
  assign _T_68223 = $signed(_T_68220) + $signed(_GEN_347); // @[Modules.scala 150:103:@14461.4]
  assign _T_68224 = _T_68223[5:0]; // @[Modules.scala 150:103:@14462.4]
  assign _T_68225 = $signed(_T_68224); // @[Modules.scala 150:103:@14463.4]
  assign _GEN_348 = {{1{_T_56005[4]}},_T_56005}; // @[Modules.scala 150:103:@14479.4]
  assign _T_68244 = $signed(_T_65200) + $signed(_GEN_348); // @[Modules.scala 150:103:@14479.4]
  assign _T_68245 = _T_68244[5:0]; // @[Modules.scala 150:103:@14480.4]
  assign _T_68246 = $signed(_T_68245); // @[Modules.scala 150:103:@14481.4]
  assign _T_68251 = $signed(_T_56007) + $signed(_T_56012); // @[Modules.scala 150:103:@14485.4]
  assign _T_68252 = _T_68251[4:0]; // @[Modules.scala 150:103:@14486.4]
  assign _T_68253 = $signed(_T_68252); // @[Modules.scala 150:103:@14487.4]
  assign _T_68257 = $signed(4'sh1) * $signed(io_in_668); // @[Modules.scala 151:80:@14490.4]
  assign _GEN_349 = {{1{_T_56014[4]}},_T_56014}; // @[Modules.scala 150:103:@14491.4]
  assign _T_68258 = $signed(_GEN_349) + $signed(_T_68257); // @[Modules.scala 150:103:@14491.4]
  assign _T_68259 = _T_68258[5:0]; // @[Modules.scala 150:103:@14492.4]
  assign _T_68260 = $signed(_T_68259); // @[Modules.scala 150:103:@14493.4]
  assign _GEN_351 = {{1{_T_62140[4]}},_T_62140}; // @[Modules.scala 150:103:@14509.4]
  assign _T_68279 = $signed(_GEN_351) + $signed(_T_56040); // @[Modules.scala 150:103:@14509.4]
  assign _T_68280 = _T_68279[5:0]; // @[Modules.scala 150:103:@14510.4]
  assign _T_68281 = $signed(_T_68280); // @[Modules.scala 150:103:@14511.4]
  assign _GEN_352 = {{1{_T_65251[4]}},_T_65251}; // @[Modules.scala 150:103:@14515.4]
  assign _T_68286 = $signed(_T_56042) + $signed(_GEN_352); // @[Modules.scala 150:103:@14515.4]
  assign _T_68287 = _T_68286[5:0]; // @[Modules.scala 150:103:@14516.4]
  assign _T_68288 = $signed(_T_68287); // @[Modules.scala 150:103:@14517.4]
  assign _T_68293 = $signed(_T_56049) + $signed(_T_56056); // @[Modules.scala 150:103:@14521.4]
  assign _T_68294 = _T_68293[4:0]; // @[Modules.scala 150:103:@14522.4]
  assign _T_68295 = $signed(_T_68294); // @[Modules.scala 150:103:@14523.4]
  assign _T_68300 = $signed(_T_65265) + $signed(_T_59066); // @[Modules.scala 150:103:@14527.4]
  assign _T_68301 = _T_68300[4:0]; // @[Modules.scala 150:103:@14528.4]
  assign _T_68302 = $signed(_T_68301); // @[Modules.scala 150:103:@14529.4]
  assign _GEN_353 = {{1{_T_56075[4]}},_T_56075}; // @[Modules.scala 150:103:@14545.4]
  assign _T_68321 = $signed(_GEN_353) + $signed(_T_59094); // @[Modules.scala 150:103:@14545.4]
  assign _T_68322 = _T_68321[5:0]; // @[Modules.scala 150:103:@14546.4]
  assign _T_68323 = $signed(_T_68322); // @[Modules.scala 150:103:@14547.4]
  assign _T_68335 = $signed(_T_62194) + $signed(_T_56098); // @[Modules.scala 150:103:@14557.4]
  assign _T_68336 = _T_68335[5:0]; // @[Modules.scala 150:103:@14558.4]
  assign _T_68337 = $signed(_T_68336); // @[Modules.scala 150:103:@14559.4]
  assign _T_68341 = $signed(-4'sh1) * $signed(io_in_698); // @[Modules.scala 151:80:@14562.4]
  assign _T_68342 = $signed(_T_65314) + $signed(_T_68341); // @[Modules.scala 150:103:@14563.4]
  assign _T_68343 = _T_68342[4:0]; // @[Modules.scala 150:103:@14564.4]
  assign _T_68344 = $signed(_T_68343); // @[Modules.scala 150:103:@14565.4]
  assign _T_68349 = $signed(_T_62203) + $signed(_T_59122); // @[Modules.scala 150:103:@14569.4]
  assign _T_68350 = _T_68349[4:0]; // @[Modules.scala 150:103:@14570.4]
  assign _T_68351 = $signed(_T_68350); // @[Modules.scala 150:103:@14571.4]
  assign _GEN_354 = {{1{_T_62210[4]}},_T_62210}; // @[Modules.scala 150:103:@14575.4]
  assign _T_68356 = $signed(_GEN_354) + $signed(_T_59124); // @[Modules.scala 150:103:@14575.4]
  assign _T_68357 = _T_68356[5:0]; // @[Modules.scala 150:103:@14576.4]
  assign _T_68358 = $signed(_T_68357); // @[Modules.scala 150:103:@14577.4]
  assign _T_68423 = $signed(4'sh1) * $signed(io_in_724); // @[Modules.scala 150:74:@14633.4]
  assign _T_68426 = $signed(_T_68423) + $signed(_T_59185); // @[Modules.scala 150:103:@14635.4]
  assign _T_68427 = _T_68426[5:0]; // @[Modules.scala 150:103:@14636.4]
  assign _T_68428 = $signed(_T_68427); // @[Modules.scala 150:103:@14637.4]
  assign _T_68433 = $signed(_GEN_139) + $signed(_T_62278); // @[Modules.scala 150:103:@14641.4]
  assign _T_68434 = _T_68433[5:0]; // @[Modules.scala 150:103:@14642.4]
  assign _T_68435 = $signed(_T_68434); // @[Modules.scala 150:103:@14643.4]
  assign _T_68447 = $signed(_T_59201) + $signed(_T_59206); // @[Modules.scala 150:103:@14653.4]
  assign _T_68448 = _T_68447[5:0]; // @[Modules.scala 150:103:@14654.4]
  assign _T_68449 = $signed(_T_68448); // @[Modules.scala 150:103:@14655.4]
  assign _T_68454 = $signed(_T_56196) + $signed(_T_56201); // @[Modules.scala 150:103:@14659.4]
  assign _T_68455 = _T_68454[5:0]; // @[Modules.scala 150:103:@14660.4]
  assign _T_68456 = $signed(_T_68455); // @[Modules.scala 150:103:@14661.4]
  assign _T_68461 = $signed(_T_56203) + $signed(_T_56208); // @[Modules.scala 150:103:@14665.4]
  assign _T_68462 = _T_68461[5:0]; // @[Modules.scala 150:103:@14666.4]
  assign _T_68463 = $signed(_T_68462); // @[Modules.scala 150:103:@14667.4]
  assign _T_68468 = $signed(_T_56210) + $signed(_T_59227); // @[Modules.scala 150:103:@14671.4]
  assign _T_68469 = _T_68468[5:0]; // @[Modules.scala 150:103:@14672.4]
  assign _T_68470 = $signed(_T_68469); // @[Modules.scala 150:103:@14673.4]
  assign _T_68475 = $signed(_T_59229) + $signed(_T_59234); // @[Modules.scala 150:103:@14677.4]
  assign _T_68476 = _T_68475[5:0]; // @[Modules.scala 150:103:@14678.4]
  assign _T_68477 = $signed(_T_68476); // @[Modules.scala 150:103:@14679.4]
  assign _T_68482 = $signed(_T_56217) + $signed(_T_56222); // @[Modules.scala 150:103:@14683.4]
  assign _T_68483 = _T_68482[5:0]; // @[Modules.scala 150:103:@14684.4]
  assign _T_68484 = $signed(_T_68483); // @[Modules.scala 150:103:@14685.4]
  assign _T_68489 = $signed(_T_59243) + $signed(_T_59248); // @[Modules.scala 150:103:@14689.4]
  assign _T_68490 = _T_68489[5:0]; // @[Modules.scala 150:103:@14690.4]
  assign _T_68491 = $signed(_T_68490); // @[Modules.scala 150:103:@14691.4]
  assign _T_68496 = $signed(_T_59250) + $signed(_T_59255); // @[Modules.scala 150:103:@14695.4]
  assign _T_68497 = _T_68496[5:0]; // @[Modules.scala 150:103:@14696.4]
  assign _T_68498 = $signed(_T_68497); // @[Modules.scala 150:103:@14697.4]
  assign _T_68500 = $signed(4'sh1) * $signed(io_in_750); // @[Modules.scala 150:74:@14699.4]
  assign _T_68502 = $signed(4'sh1) * $signed(io_in_751); // @[Modules.scala 151:80:@14700.4]
  assign _T_68503 = $signed(_T_68500) + $signed(_T_68502); // @[Modules.scala 150:103:@14701.4]
  assign _T_68504 = _T_68503[5:0]; // @[Modules.scala 150:103:@14702.4]
  assign _T_68505 = $signed(_T_68504); // @[Modules.scala 150:103:@14703.4]
  assign _T_68523 = $signed(4'sh1) * $signed(io_in_763); // @[Modules.scala 151:80:@14718.4]
  assign _T_68524 = $signed(_T_59276) + $signed(_T_68523); // @[Modules.scala 150:103:@14719.4]
  assign _T_68525 = _T_68524[5:0]; // @[Modules.scala 150:103:@14720.4]
  assign _T_68526 = $signed(_T_68525); // @[Modules.scala 150:103:@14721.4]
  assign _GEN_356 = {{1{_T_62399[4]}},_T_62399}; // @[Modules.scala 150:103:@14743.4]
  assign _T_68552 = $signed(_GEN_356) + $signed(_T_59313); // @[Modules.scala 150:103:@14743.4]
  assign _T_68553 = _T_68552[5:0]; // @[Modules.scala 150:103:@14744.4]
  assign _T_68554 = $signed(_T_68553); // @[Modules.scala 150:103:@14745.4]
  assign buffer_4_2 = {{8{_T_66496[5]}},_T_66496}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_3 = {{9{_T_66503[4]}},_T_66503}; // @[Modules.scala 112:22:@8.4]
  assign _T_68574 = $signed(buffer_4_2) + $signed(buffer_4_3); // @[Modules.scala 160:64:@14765.4]
  assign _T_68575 = _T_68574[13:0]; // @[Modules.scala 160:64:@14766.4]
  assign buffer_4_301 = $signed(_T_68575); // @[Modules.scala 160:64:@14767.4]
  assign buffer_4_4 = {{9{_T_66510[4]}},_T_66510}; // @[Modules.scala 112:22:@8.4]
  assign _T_68577 = $signed(buffer_4_4) + $signed(buffer_1_6); // @[Modules.scala 160:64:@14769.4]
  assign _T_68578 = _T_68577[13:0]; // @[Modules.scala 160:64:@14770.4]
  assign buffer_4_302 = $signed(_T_68578); // @[Modules.scala 160:64:@14771.4]
  assign buffer_4_6 = {{8{_T_66524[5]}},_T_66524}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_7 = {{8{_T_66531[5]}},_T_66531}; // @[Modules.scala 112:22:@8.4]
  assign _T_68580 = $signed(buffer_4_6) + $signed(buffer_4_7); // @[Modules.scala 160:64:@14773.4]
  assign _T_68581 = _T_68580[13:0]; // @[Modules.scala 160:64:@14774.4]
  assign buffer_4_303 = $signed(_T_68581); // @[Modules.scala 160:64:@14775.4]
  assign buffer_4_9 = {{9{_T_66545[4]}},_T_66545}; // @[Modules.scala 112:22:@8.4]
  assign _T_68583 = $signed(buffer_3_9) + $signed(buffer_4_9); // @[Modules.scala 160:64:@14777.4]
  assign _T_68584 = _T_68583[13:0]; // @[Modules.scala 160:64:@14778.4]
  assign buffer_4_304 = $signed(_T_68584); // @[Modules.scala 160:64:@14779.4]
  assign buffer_4_10 = {{8{_T_66552[5]}},_T_66552}; // @[Modules.scala 112:22:@8.4]
  assign _T_68586 = $signed(buffer_4_10) + $signed(buffer_0_12); // @[Modules.scala 160:64:@14781.4]
  assign _T_68587 = _T_68586[13:0]; // @[Modules.scala 160:64:@14782.4]
  assign buffer_4_305 = $signed(_T_68587); // @[Modules.scala 160:64:@14783.4]
  assign buffer_4_12 = {{9{_T_66566[4]}},_T_66566}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_13 = {{9{_T_66573[4]}},_T_66573}; // @[Modules.scala 112:22:@8.4]
  assign _T_68589 = $signed(buffer_4_12) + $signed(buffer_4_13); // @[Modules.scala 160:64:@14785.4]
  assign _T_68590 = _T_68589[13:0]; // @[Modules.scala 160:64:@14786.4]
  assign buffer_4_306 = $signed(_T_68590); // @[Modules.scala 160:64:@14787.4]
  assign _T_68595 = $signed(buffer_2_16) + $signed(buffer_1_18); // @[Modules.scala 160:64:@14793.4]
  assign _T_68596 = _T_68595[13:0]; // @[Modules.scala 160:64:@14794.4]
  assign buffer_4_308 = $signed(_T_68596); // @[Modules.scala 160:64:@14795.4]
  assign buffer_4_18 = {{9{_T_66608[4]}},_T_66608}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_19 = {{8{_T_66615[5]}},_T_66615}; // @[Modules.scala 112:22:@8.4]
  assign _T_68598 = $signed(buffer_4_18) + $signed(buffer_4_19); // @[Modules.scala 160:64:@14797.4]
  assign _T_68599 = _T_68598[13:0]; // @[Modules.scala 160:64:@14798.4]
  assign buffer_4_309 = $signed(_T_68599); // @[Modules.scala 160:64:@14799.4]
  assign buffer_4_21 = {{8{_T_66629[5]}},_T_66629}; // @[Modules.scala 112:22:@8.4]
  assign _T_68601 = $signed(buffer_1_21) + $signed(buffer_4_21); // @[Modules.scala 160:64:@14801.4]
  assign _T_68602 = _T_68601[13:0]; // @[Modules.scala 160:64:@14802.4]
  assign buffer_4_310 = $signed(_T_68602); // @[Modules.scala 160:64:@14803.4]
  assign _T_68604 = $signed(buffer_3_23) + $signed(buffer_3_24); // @[Modules.scala 160:64:@14805.4]
  assign _T_68605 = _T_68604[13:0]; // @[Modules.scala 160:64:@14806.4]
  assign buffer_4_311 = $signed(_T_68605); // @[Modules.scala 160:64:@14807.4]
  assign _T_68607 = $signed(buffer_3_25) + $signed(buffer_3_26); // @[Modules.scala 160:64:@14809.4]
  assign _T_68608 = _T_68607[13:0]; // @[Modules.scala 160:64:@14810.4]
  assign buffer_4_312 = $signed(_T_68608); // @[Modules.scala 160:64:@14811.4]
  assign _T_68610 = $signed(buffer_3_27) + $signed(buffer_3_28); // @[Modules.scala 160:64:@14813.4]
  assign _T_68611 = _T_68610[13:0]; // @[Modules.scala 160:64:@14814.4]
  assign buffer_4_313 = $signed(_T_68611); // @[Modules.scala 160:64:@14815.4]
  assign _T_68613 = $signed(buffer_3_29) + $signed(buffer_3_30); // @[Modules.scala 160:64:@14817.4]
  assign _T_68614 = _T_68613[13:0]; // @[Modules.scala 160:64:@14818.4]
  assign buffer_4_314 = $signed(_T_68614); // @[Modules.scala 160:64:@14819.4]
  assign buffer_4_30 = {{8{_T_66692[5]}},_T_66692}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_31 = {{8{_T_66699[5]}},_T_66699}; // @[Modules.scala 112:22:@8.4]
  assign _T_68616 = $signed(buffer_4_30) + $signed(buffer_4_31); // @[Modules.scala 160:64:@14821.4]
  assign _T_68617 = _T_68616[13:0]; // @[Modules.scala 160:64:@14822.4]
  assign buffer_4_315 = $signed(_T_68617); // @[Modules.scala 160:64:@14823.4]
  assign buffer_4_33 = {{8{_T_66713[5]}},_T_66713}; // @[Modules.scala 112:22:@8.4]
  assign _T_68619 = $signed(buffer_0_34) + $signed(buffer_4_33); // @[Modules.scala 160:64:@14825.4]
  assign _T_68620 = _T_68619[13:0]; // @[Modules.scala 160:64:@14826.4]
  assign buffer_4_316 = $signed(_T_68620); // @[Modules.scala 160:64:@14827.4]
  assign buffer_4_34 = {{8{_T_66720[5]}},_T_66720}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_35 = {{9{_T_66727[4]}},_T_66727}; // @[Modules.scala 112:22:@8.4]
  assign _T_68622 = $signed(buffer_4_34) + $signed(buffer_4_35); // @[Modules.scala 160:64:@14829.4]
  assign _T_68623 = _T_68622[13:0]; // @[Modules.scala 160:64:@14830.4]
  assign buffer_4_317 = $signed(_T_68623); // @[Modules.scala 160:64:@14831.4]
  assign buffer_4_36 = {{9{_T_66734[4]}},_T_66734}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_37 = {{9{_T_66741[4]}},_T_66741}; // @[Modules.scala 112:22:@8.4]
  assign _T_68625 = $signed(buffer_4_36) + $signed(buffer_4_37); // @[Modules.scala 160:64:@14833.4]
  assign _T_68626 = _T_68625[13:0]; // @[Modules.scala 160:64:@14834.4]
  assign buffer_4_318 = $signed(_T_68626); // @[Modules.scala 160:64:@14835.4]
  assign buffer_4_39 = {{8{_T_66755[5]}},_T_66755}; // @[Modules.scala 112:22:@8.4]
  assign _T_68628 = $signed(buffer_2_36) + $signed(buffer_4_39); // @[Modules.scala 160:64:@14837.4]
  assign _T_68629 = _T_68628[13:0]; // @[Modules.scala 160:64:@14838.4]
  assign buffer_4_319 = $signed(_T_68629); // @[Modules.scala 160:64:@14839.4]
  assign buffer_4_41 = {{8{_T_66769[5]}},_T_66769}; // @[Modules.scala 112:22:@8.4]
  assign _T_68631 = $signed(buffer_1_41) + $signed(buffer_4_41); // @[Modules.scala 160:64:@14841.4]
  assign _T_68632 = _T_68631[13:0]; // @[Modules.scala 160:64:@14842.4]
  assign buffer_4_320 = $signed(_T_68632); // @[Modules.scala 160:64:@14843.4]
  assign buffer_4_42 = {{9{_T_66776[4]}},_T_66776}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_43 = {{8{_T_66783[5]}},_T_66783}; // @[Modules.scala 112:22:@8.4]
  assign _T_68634 = $signed(buffer_4_42) + $signed(buffer_4_43); // @[Modules.scala 160:64:@14845.4]
  assign _T_68635 = _T_68634[13:0]; // @[Modules.scala 160:64:@14846.4]
  assign buffer_4_321 = $signed(_T_68635); // @[Modules.scala 160:64:@14847.4]
  assign buffer_4_44 = {{8{_T_66790[5]}},_T_66790}; // @[Modules.scala 112:22:@8.4]
  assign _T_68637 = $signed(buffer_4_44) + $signed(buffer_2_45); // @[Modules.scala 160:64:@14849.4]
  assign _T_68638 = _T_68637[13:0]; // @[Modules.scala 160:64:@14850.4]
  assign buffer_4_322 = $signed(_T_68638); // @[Modules.scala 160:64:@14851.4]
  assign buffer_4_49 = {{9{_T_66825[4]}},_T_66825}; // @[Modules.scala 112:22:@8.4]
  assign _T_68643 = $signed(buffer_3_50) + $signed(buffer_4_49); // @[Modules.scala 160:64:@14857.4]
  assign _T_68644 = _T_68643[13:0]; // @[Modules.scala 160:64:@14858.4]
  assign buffer_4_324 = $signed(_T_68644); // @[Modules.scala 160:64:@14859.4]
  assign buffer_4_52 = {{9{_T_66846[4]}},_T_66846}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_53 = {{9{_T_66853[4]}},_T_66853}; // @[Modules.scala 112:22:@8.4]
  assign _T_68649 = $signed(buffer_4_52) + $signed(buffer_4_53); // @[Modules.scala 160:64:@14865.4]
  assign _T_68650 = _T_68649[13:0]; // @[Modules.scala 160:64:@14866.4]
  assign buffer_4_326 = $signed(_T_68650); // @[Modules.scala 160:64:@14867.4]
  assign buffer_4_55 = {{9{_T_66867[4]}},_T_66867}; // @[Modules.scala 112:22:@8.4]
  assign _T_68652 = $signed(buffer_0_52) + $signed(buffer_4_55); // @[Modules.scala 160:64:@14869.4]
  assign _T_68653 = _T_68652[13:0]; // @[Modules.scala 160:64:@14870.4]
  assign buffer_4_327 = $signed(_T_68653); // @[Modules.scala 160:64:@14871.4]
  assign buffer_4_56 = {{8{_T_66874[5]}},_T_66874}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_57 = {{8{_T_66881[5]}},_T_66881}; // @[Modules.scala 112:22:@8.4]
  assign _T_68655 = $signed(buffer_4_56) + $signed(buffer_4_57); // @[Modules.scala 160:64:@14873.4]
  assign _T_68656 = _T_68655[13:0]; // @[Modules.scala 160:64:@14874.4]
  assign buffer_4_328 = $signed(_T_68656); // @[Modules.scala 160:64:@14875.4]
  assign buffer_4_61 = {{9{_T_66909[4]}},_T_66909}; // @[Modules.scala 112:22:@8.4]
  assign _T_68661 = $signed(buffer_3_62) + $signed(buffer_4_61); // @[Modules.scala 160:64:@14881.4]
  assign _T_68662 = _T_68661[13:0]; // @[Modules.scala 160:64:@14882.4]
  assign buffer_4_330 = $signed(_T_68662); // @[Modules.scala 160:64:@14883.4]
  assign buffer_4_62 = {{8{_T_66916[5]}},_T_66916}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_63 = {{8{_T_66923[5]}},_T_66923}; // @[Modules.scala 112:22:@8.4]
  assign _T_68664 = $signed(buffer_4_62) + $signed(buffer_4_63); // @[Modules.scala 160:64:@14885.4]
  assign _T_68665 = _T_68664[13:0]; // @[Modules.scala 160:64:@14886.4]
  assign buffer_4_331 = $signed(_T_68665); // @[Modules.scala 160:64:@14887.4]
  assign buffer_4_64 = {{8{_T_66930[5]}},_T_66930}; // @[Modules.scala 112:22:@8.4]
  assign _T_68667 = $signed(buffer_4_64) + $signed(buffer_1_64); // @[Modules.scala 160:64:@14889.4]
  assign _T_68668 = _T_68667[13:0]; // @[Modules.scala 160:64:@14890.4]
  assign buffer_4_332 = $signed(_T_68668); // @[Modules.scala 160:64:@14891.4]
  assign _T_68670 = $signed(buffer_1_65) + $signed(buffer_1_66); // @[Modules.scala 160:64:@14893.4]
  assign _T_68671 = _T_68670[13:0]; // @[Modules.scala 160:64:@14894.4]
  assign buffer_4_333 = $signed(_T_68671); // @[Modules.scala 160:64:@14895.4]
  assign buffer_4_71 = {{9{_T_66979[4]}},_T_66979}; // @[Modules.scala 112:22:@8.4]
  assign _T_68676 = $signed(buffer_2_68) + $signed(buffer_4_71); // @[Modules.scala 160:64:@14901.4]
  assign _T_68677 = _T_68676[13:0]; // @[Modules.scala 160:64:@14902.4]
  assign buffer_4_335 = $signed(_T_68677); // @[Modules.scala 160:64:@14903.4]
  assign buffer_4_72 = {{8{_T_66986[5]}},_T_66986}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_73 = {{8{_T_66993[5]}},_T_66993}; // @[Modules.scala 112:22:@8.4]
  assign _T_68679 = $signed(buffer_4_72) + $signed(buffer_4_73); // @[Modules.scala 160:64:@14905.4]
  assign _T_68680 = _T_68679[13:0]; // @[Modules.scala 160:64:@14906.4]
  assign buffer_4_336 = $signed(_T_68680); // @[Modules.scala 160:64:@14907.4]
  assign buffer_4_75 = {{8{_T_67007[5]}},_T_67007}; // @[Modules.scala 112:22:@8.4]
  assign _T_68682 = $signed(buffer_3_76) + $signed(buffer_4_75); // @[Modules.scala 160:64:@14909.4]
  assign _T_68683 = _T_68682[13:0]; // @[Modules.scala 160:64:@14910.4]
  assign buffer_4_337 = $signed(_T_68683); // @[Modules.scala 160:64:@14911.4]
  assign buffer_4_78 = {{8{_T_67028[5]}},_T_67028}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_79 = {{8{_T_67035[5]}},_T_67035}; // @[Modules.scala 112:22:@8.4]
  assign _T_68688 = $signed(buffer_4_78) + $signed(buffer_4_79); // @[Modules.scala 160:64:@14917.4]
  assign _T_68689 = _T_68688[13:0]; // @[Modules.scala 160:64:@14918.4]
  assign buffer_4_339 = $signed(_T_68689); // @[Modules.scala 160:64:@14919.4]
  assign buffer_4_80 = {{8{_T_67042[5]}},_T_67042}; // @[Modules.scala 112:22:@8.4]
  assign _T_68691 = $signed(buffer_4_80) + $signed(buffer_0_79); // @[Modules.scala 160:64:@14921.4]
  assign _T_68692 = _T_68691[13:0]; // @[Modules.scala 160:64:@14922.4]
  assign buffer_4_340 = $signed(_T_68692); // @[Modules.scala 160:64:@14923.4]
  assign buffer_4_82 = {{8{_T_67056[5]}},_T_67056}; // @[Modules.scala 112:22:@8.4]
  assign _T_68694 = $signed(buffer_4_82) + $signed(buffer_1_84); // @[Modules.scala 160:64:@14925.4]
  assign _T_68695 = _T_68694[13:0]; // @[Modules.scala 160:64:@14926.4]
  assign buffer_4_341 = $signed(_T_68695); // @[Modules.scala 160:64:@14927.4]
  assign buffer_4_85 = {{8{_T_67077[5]}},_T_67077}; // @[Modules.scala 112:22:@8.4]
  assign _T_68697 = $signed(buffer_1_85) + $signed(buffer_4_85); // @[Modules.scala 160:64:@14929.4]
  assign _T_68698 = _T_68697[13:0]; // @[Modules.scala 160:64:@14930.4]
  assign buffer_4_342 = $signed(_T_68698); // @[Modules.scala 160:64:@14931.4]
  assign buffer_4_90 = {{8{_T_67112[5]}},_T_67112}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_91 = {{8{_T_67119[5]}},_T_67119}; // @[Modules.scala 112:22:@8.4]
  assign _T_68706 = $signed(buffer_4_90) + $signed(buffer_4_91); // @[Modules.scala 160:64:@14941.4]
  assign _T_68707 = _T_68706[13:0]; // @[Modules.scala 160:64:@14942.4]
  assign buffer_4_345 = $signed(_T_68707); // @[Modules.scala 160:64:@14943.4]
  assign buffer_4_92 = {{9{_T_67126[4]}},_T_67126}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_93 = {{8{_T_67133[5]}},_T_67133}; // @[Modules.scala 112:22:@8.4]
  assign _T_68709 = $signed(buffer_4_92) + $signed(buffer_4_93); // @[Modules.scala 160:64:@14945.4]
  assign _T_68710 = _T_68709[13:0]; // @[Modules.scala 160:64:@14946.4]
  assign buffer_4_346 = $signed(_T_68710); // @[Modules.scala 160:64:@14947.4]
  assign buffer_4_94 = {{8{_T_67140[5]}},_T_67140}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_95 = {{8{_T_67147[5]}},_T_67147}; // @[Modules.scala 112:22:@8.4]
  assign _T_68712 = $signed(buffer_4_94) + $signed(buffer_4_95); // @[Modules.scala 160:64:@14949.4]
  assign _T_68713 = _T_68712[13:0]; // @[Modules.scala 160:64:@14950.4]
  assign buffer_4_347 = $signed(_T_68713); // @[Modules.scala 160:64:@14951.4]
  assign buffer_4_96 = {{8{_T_67154[5]}},_T_67154}; // @[Modules.scala 112:22:@8.4]
  assign _T_68715 = $signed(buffer_4_96) + $signed(buffer_0_95); // @[Modules.scala 160:64:@14953.4]
  assign _T_68716 = _T_68715[13:0]; // @[Modules.scala 160:64:@14954.4]
  assign buffer_4_348 = $signed(_T_68716); // @[Modules.scala 160:64:@14955.4]
  assign buffer_4_101 = {{8{_T_67189[5]}},_T_67189}; // @[Modules.scala 112:22:@8.4]
  assign _T_68721 = $signed(buffer_0_98) + $signed(buffer_4_101); // @[Modules.scala 160:64:@14961.4]
  assign _T_68722 = _T_68721[13:0]; // @[Modules.scala 160:64:@14962.4]
  assign buffer_4_350 = $signed(_T_68722); // @[Modules.scala 160:64:@14963.4]
  assign buffer_4_103 = {{8{_T_67203[5]}},_T_67203}; // @[Modules.scala 112:22:@8.4]
  assign _T_68724 = $signed(buffer_2_105) + $signed(buffer_4_103); // @[Modules.scala 160:64:@14965.4]
  assign _T_68725 = _T_68724[13:0]; // @[Modules.scala 160:64:@14966.4]
  assign buffer_4_351 = $signed(_T_68725); // @[Modules.scala 160:64:@14967.4]
  assign buffer_4_104 = {{8{_T_67210[5]}},_T_67210}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_105 = {{8{_T_67217[5]}},_T_67217}; // @[Modules.scala 112:22:@8.4]
  assign _T_68727 = $signed(buffer_4_104) + $signed(buffer_4_105); // @[Modules.scala 160:64:@14969.4]
  assign _T_68728 = _T_68727[13:0]; // @[Modules.scala 160:64:@14970.4]
  assign buffer_4_352 = $signed(_T_68728); // @[Modules.scala 160:64:@14971.4]
  assign buffer_4_106 = {{8{_T_67224[5]}},_T_67224}; // @[Modules.scala 112:22:@8.4]
  assign _T_68730 = $signed(buffer_4_106) + $signed(buffer_0_107); // @[Modules.scala 160:64:@14973.4]
  assign _T_68731 = _T_68730[13:0]; // @[Modules.scala 160:64:@14974.4]
  assign buffer_4_353 = $signed(_T_68731); // @[Modules.scala 160:64:@14975.4]
  assign _T_68733 = $signed(buffer_2_111) + $signed(buffer_1_111); // @[Modules.scala 160:64:@14977.4]
  assign _T_68734 = _T_68733[13:0]; // @[Modules.scala 160:64:@14978.4]
  assign buffer_4_354 = $signed(_T_68734); // @[Modules.scala 160:64:@14979.4]
  assign buffer_4_110 = {{8{_T_67252[5]}},_T_67252}; // @[Modules.scala 112:22:@8.4]
  assign _T_68736 = $signed(buffer_4_110) + $signed(buffer_0_111); // @[Modules.scala 160:64:@14981.4]
  assign _T_68737 = _T_68736[13:0]; // @[Modules.scala 160:64:@14982.4]
  assign buffer_4_355 = $signed(_T_68737); // @[Modules.scala 160:64:@14983.4]
  assign buffer_4_112 = {{9{_T_67266[4]}},_T_67266}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_113 = {{8{_T_67273[5]}},_T_67273}; // @[Modules.scala 112:22:@8.4]
  assign _T_68739 = $signed(buffer_4_112) + $signed(buffer_4_113); // @[Modules.scala 160:64:@14985.4]
  assign _T_68740 = _T_68739[13:0]; // @[Modules.scala 160:64:@14986.4]
  assign buffer_4_356 = $signed(_T_68740); // @[Modules.scala 160:64:@14987.4]
  assign buffer_4_114 = {{8{_T_67280[5]}},_T_67280}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_115 = {{8{_T_67287[5]}},_T_67287}; // @[Modules.scala 112:22:@8.4]
  assign _T_68742 = $signed(buffer_4_114) + $signed(buffer_4_115); // @[Modules.scala 160:64:@14989.4]
  assign _T_68743 = _T_68742[13:0]; // @[Modules.scala 160:64:@14990.4]
  assign buffer_4_357 = $signed(_T_68743); // @[Modules.scala 160:64:@14991.4]
  assign buffer_4_117 = {{8{_T_67301[5]}},_T_67301}; // @[Modules.scala 112:22:@8.4]
  assign _T_68745 = $signed(buffer_2_120) + $signed(buffer_4_117); // @[Modules.scala 160:64:@14993.4]
  assign _T_68746 = _T_68745[13:0]; // @[Modules.scala 160:64:@14994.4]
  assign buffer_4_358 = $signed(_T_68746); // @[Modules.scala 160:64:@14995.4]
  assign buffer_4_118 = {{8{_T_67308[5]}},_T_67308}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_119 = {{8{_T_67315[5]}},_T_67315}; // @[Modules.scala 112:22:@8.4]
  assign _T_68748 = $signed(buffer_4_118) + $signed(buffer_4_119); // @[Modules.scala 160:64:@14997.4]
  assign _T_68749 = _T_68748[13:0]; // @[Modules.scala 160:64:@14998.4]
  assign buffer_4_359 = $signed(_T_68749); // @[Modules.scala 160:64:@14999.4]
  assign buffer_4_121 = {{8{_T_67329[5]}},_T_67329}; // @[Modules.scala 112:22:@8.4]
  assign _T_68751 = $signed(buffer_1_124) + $signed(buffer_4_121); // @[Modules.scala 160:64:@15001.4]
  assign _T_68752 = _T_68751[13:0]; // @[Modules.scala 160:64:@15002.4]
  assign buffer_4_360 = $signed(_T_68752); // @[Modules.scala 160:64:@15003.4]
  assign buffer_4_123 = {{9{_T_67343[4]}},_T_67343}; // @[Modules.scala 112:22:@8.4]
  assign _T_68754 = $signed(buffer_0_124) + $signed(buffer_4_123); // @[Modules.scala 160:64:@15005.4]
  assign _T_68755 = _T_68754[13:0]; // @[Modules.scala 160:64:@15006.4]
  assign buffer_4_361 = $signed(_T_68755); // @[Modules.scala 160:64:@15007.4]
  assign buffer_4_124 = {{8{_T_67350[5]}},_T_67350}; // @[Modules.scala 112:22:@8.4]
  assign _T_68757 = $signed(buffer_4_124) + $signed(buffer_1_129); // @[Modules.scala 160:64:@15009.4]
  assign _T_68758 = _T_68757[13:0]; // @[Modules.scala 160:64:@15010.4]
  assign buffer_4_362 = $signed(_T_68758); // @[Modules.scala 160:64:@15011.4]
  assign buffer_4_127 = {{8{_T_67371[5]}},_T_67371}; // @[Modules.scala 112:22:@8.4]
  assign _T_68760 = $signed(buffer_3_135) + $signed(buffer_4_127); // @[Modules.scala 160:64:@15013.4]
  assign _T_68761 = _T_68760[13:0]; // @[Modules.scala 160:64:@15014.4]
  assign buffer_4_363 = $signed(_T_68761); // @[Modules.scala 160:64:@15015.4]
  assign buffer_4_129 = {{8{_T_67385[5]}},_T_67385}; // @[Modules.scala 112:22:@8.4]
  assign _T_68763 = $signed(buffer_1_132) + $signed(buffer_4_129); // @[Modules.scala 160:64:@15017.4]
  assign _T_68764 = _T_68763[13:0]; // @[Modules.scala 160:64:@15018.4]
  assign buffer_4_364 = $signed(_T_68764); // @[Modules.scala 160:64:@15019.4]
  assign buffer_4_130 = {{8{_T_67392[5]}},_T_67392}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_131 = {{8{_T_67399[5]}},_T_67399}; // @[Modules.scala 112:22:@8.4]
  assign _T_68766 = $signed(buffer_4_130) + $signed(buffer_4_131); // @[Modules.scala 160:64:@15021.4]
  assign _T_68767 = _T_68766[13:0]; // @[Modules.scala 160:64:@15022.4]
  assign buffer_4_365 = $signed(_T_68767); // @[Modules.scala 160:64:@15023.4]
  assign buffer_4_133 = {{8{_T_67413[5]}},_T_67413}; // @[Modules.scala 112:22:@8.4]
  assign _T_68769 = $signed(buffer_1_136) + $signed(buffer_4_133); // @[Modules.scala 160:64:@15025.4]
  assign _T_68770 = _T_68769[13:0]; // @[Modules.scala 160:64:@15026.4]
  assign buffer_4_366 = $signed(_T_68770); // @[Modules.scala 160:64:@15027.4]
  assign buffer_4_135 = {{9{_T_67427[4]}},_T_67427}; // @[Modules.scala 112:22:@8.4]
  assign _T_68772 = $signed(buffer_3_143) + $signed(buffer_4_135); // @[Modules.scala 160:64:@15029.4]
  assign _T_68773 = _T_68772[13:0]; // @[Modules.scala 160:64:@15030.4]
  assign buffer_4_367 = $signed(_T_68773); // @[Modules.scala 160:64:@15031.4]
  assign buffer_4_137 = {{8{_T_67441[5]}},_T_67441}; // @[Modules.scala 112:22:@8.4]
  assign _T_68775 = $signed(buffer_2_141) + $signed(buffer_4_137); // @[Modules.scala 160:64:@15033.4]
  assign _T_68776 = _T_68775[13:0]; // @[Modules.scala 160:64:@15034.4]
  assign buffer_4_368 = $signed(_T_68776); // @[Modules.scala 160:64:@15035.4]
  assign _T_68778 = $signed(buffer_3_147) + $signed(buffer_1_143); // @[Modules.scala 160:64:@15037.4]
  assign _T_68779 = _T_68778[13:0]; // @[Modules.scala 160:64:@15038.4]
  assign buffer_4_369 = $signed(_T_68779); // @[Modules.scala 160:64:@15039.4]
  assign buffer_4_141 = {{8{_T_67469[5]}},_T_67469}; // @[Modules.scala 112:22:@8.4]
  assign _T_68781 = $signed(buffer_1_144) + $signed(buffer_4_141); // @[Modules.scala 160:64:@15041.4]
  assign _T_68782 = _T_68781[13:0]; // @[Modules.scala 160:64:@15042.4]
  assign buffer_4_370 = $signed(_T_68782); // @[Modules.scala 160:64:@15043.4]
  assign buffer_4_142 = {{8{_T_67476[5]}},_T_67476}; // @[Modules.scala 112:22:@8.4]
  assign _T_68784 = $signed(buffer_4_142) + $signed(buffer_1_148); // @[Modules.scala 160:64:@15045.4]
  assign _T_68785 = _T_68784[13:0]; // @[Modules.scala 160:64:@15046.4]
  assign buffer_4_371 = $signed(_T_68785); // @[Modules.scala 160:64:@15047.4]
  assign buffer_4_144 = {{8{_T_67490[5]}},_T_67490}; // @[Modules.scala 112:22:@8.4]
  assign _T_68787 = $signed(buffer_4_144) + $signed(buffer_3_157); // @[Modules.scala 160:64:@15049.4]
  assign _T_68788 = _T_68787[13:0]; // @[Modules.scala 160:64:@15050.4]
  assign buffer_4_372 = $signed(_T_68788); // @[Modules.scala 160:64:@15051.4]
  assign buffer_4_146 = {{9{_T_67504[4]}},_T_67504}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_147 = {{8{_T_67511[5]}},_T_67511}; // @[Modules.scala 112:22:@8.4]
  assign _T_68790 = $signed(buffer_4_146) + $signed(buffer_4_147); // @[Modules.scala 160:64:@15053.4]
  assign _T_68791 = _T_68790[13:0]; // @[Modules.scala 160:64:@15054.4]
  assign buffer_4_373 = $signed(_T_68791); // @[Modules.scala 160:64:@15055.4]
  assign buffer_4_148 = {{8{_T_67518[5]}},_T_67518}; // @[Modules.scala 112:22:@8.4]
  assign _T_68793 = $signed(buffer_4_148) + $signed(buffer_1_154); // @[Modules.scala 160:64:@15057.4]
  assign _T_68794 = _T_68793[13:0]; // @[Modules.scala 160:64:@15058.4]
  assign buffer_4_374 = $signed(_T_68794); // @[Modules.scala 160:64:@15059.4]
  assign _T_68796 = $signed(buffer_0_153) + $signed(buffer_0_154); // @[Modules.scala 160:64:@15061.4]
  assign _T_68797 = _T_68796[13:0]; // @[Modules.scala 160:64:@15062.4]
  assign buffer_4_375 = $signed(_T_68797); // @[Modules.scala 160:64:@15063.4]
  assign buffer_4_153 = {{9{_T_67553[4]}},_T_67553}; // @[Modules.scala 112:22:@8.4]
  assign _T_68799 = $signed(buffer_0_155) + $signed(buffer_4_153); // @[Modules.scala 160:64:@15065.4]
  assign _T_68800 = _T_68799[13:0]; // @[Modules.scala 160:64:@15066.4]
  assign buffer_4_376 = $signed(_T_68800); // @[Modules.scala 160:64:@15067.4]
  assign buffer_4_155 = {{8{_T_67567[5]}},_T_67567}; // @[Modules.scala 112:22:@8.4]
  assign _T_68802 = $signed(buffer_3_164) + $signed(buffer_4_155); // @[Modules.scala 160:64:@15069.4]
  assign _T_68803 = _T_68802[13:0]; // @[Modules.scala 160:64:@15070.4]
  assign buffer_4_377 = $signed(_T_68803); // @[Modules.scala 160:64:@15071.4]
  assign _T_68805 = $signed(buffer_2_164) + $signed(buffer_1_161); // @[Modules.scala 160:64:@15073.4]
  assign _T_68806 = _T_68805[13:0]; // @[Modules.scala 160:64:@15074.4]
  assign buffer_4_378 = $signed(_T_68806); // @[Modules.scala 160:64:@15075.4]
  assign buffer_4_158 = {{8{_T_67588[5]}},_T_67588}; // @[Modules.scala 112:22:@8.4]
  assign _T_68808 = $signed(buffer_4_158) + $signed(buffer_1_163); // @[Modules.scala 160:64:@15077.4]
  assign _T_68809 = _T_68808[13:0]; // @[Modules.scala 160:64:@15078.4]
  assign buffer_4_379 = $signed(_T_68809); // @[Modules.scala 160:64:@15079.4]
  assign buffer_4_160 = {{8{_T_67602[5]}},_T_67602}; // @[Modules.scala 112:22:@8.4]
  assign _T_68811 = $signed(buffer_4_160) + $signed(buffer_0_164); // @[Modules.scala 160:64:@15081.4]
  assign _T_68812 = _T_68811[13:0]; // @[Modules.scala 160:64:@15082.4]
  assign buffer_4_380 = $signed(_T_68812); // @[Modules.scala 160:64:@15083.4]
  assign buffer_4_162 = {{9{_T_67616[4]}},_T_67616}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_163 = {{9{_T_67623[4]}},_T_67623}; // @[Modules.scala 112:22:@8.4]
  assign _T_68814 = $signed(buffer_4_162) + $signed(buffer_4_163); // @[Modules.scala 160:64:@15085.4]
  assign _T_68815 = _T_68814[13:0]; // @[Modules.scala 160:64:@15086.4]
  assign buffer_4_381 = $signed(_T_68815); // @[Modules.scala 160:64:@15087.4]
  assign buffer_4_164 = {{8{_T_67630[5]}},_T_67630}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_165 = {{8{_T_67637[5]}},_T_67637}; // @[Modules.scala 112:22:@8.4]
  assign _T_68817 = $signed(buffer_4_164) + $signed(buffer_4_165); // @[Modules.scala 160:64:@15089.4]
  assign _T_68818 = _T_68817[13:0]; // @[Modules.scala 160:64:@15090.4]
  assign buffer_4_382 = $signed(_T_68818); // @[Modules.scala 160:64:@15091.4]
  assign buffer_4_166 = {{8{_T_67644[5]}},_T_67644}; // @[Modules.scala 112:22:@8.4]
  assign _T_68820 = $signed(buffer_4_166) + $signed(buffer_1_171); // @[Modules.scala 160:64:@15093.4]
  assign _T_68821 = _T_68820[13:0]; // @[Modules.scala 160:64:@15094.4]
  assign buffer_4_383 = $signed(_T_68821); // @[Modules.scala 160:64:@15095.4]
  assign buffer_4_169 = {{8{_T_67665[5]}},_T_67665}; // @[Modules.scala 112:22:@8.4]
  assign _T_68823 = $signed(buffer_1_172) + $signed(buffer_4_169); // @[Modules.scala 160:64:@15097.4]
  assign _T_68824 = _T_68823[13:0]; // @[Modules.scala 160:64:@15098.4]
  assign buffer_4_384 = $signed(_T_68824); // @[Modules.scala 160:64:@15099.4]
  assign buffer_4_170 = {{9{_T_67672[4]}},_T_67672}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_171 = {{8{_T_67679[5]}},_T_67679}; // @[Modules.scala 112:22:@8.4]
  assign _T_68826 = $signed(buffer_4_170) + $signed(buffer_4_171); // @[Modules.scala 160:64:@15101.4]
  assign _T_68827 = _T_68826[13:0]; // @[Modules.scala 160:64:@15102.4]
  assign buffer_4_385 = $signed(_T_68827); // @[Modules.scala 160:64:@15103.4]
  assign buffer_4_172 = {{9{_T_67686[4]}},_T_67686}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_173 = {{9{_T_67693[4]}},_T_67693}; // @[Modules.scala 112:22:@8.4]
  assign _T_68829 = $signed(buffer_4_172) + $signed(buffer_4_173); // @[Modules.scala 160:64:@15105.4]
  assign _T_68830 = _T_68829[13:0]; // @[Modules.scala 160:64:@15106.4]
  assign buffer_4_386 = $signed(_T_68830); // @[Modules.scala 160:64:@15107.4]
  assign buffer_4_174 = {{9{_T_67700[4]}},_T_67700}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_175 = {{8{_T_67707[5]}},_T_67707}; // @[Modules.scala 112:22:@8.4]
  assign _T_68832 = $signed(buffer_4_174) + $signed(buffer_4_175); // @[Modules.scala 160:64:@15109.4]
  assign _T_68833 = _T_68832[13:0]; // @[Modules.scala 160:64:@15110.4]
  assign buffer_4_387 = $signed(_T_68833); // @[Modules.scala 160:64:@15111.4]
  assign _T_68838 = $signed(buffer_3_194) + $signed(buffer_2_192); // @[Modules.scala 160:64:@15117.4]
  assign _T_68839 = _T_68838[13:0]; // @[Modules.scala 160:64:@15118.4]
  assign buffer_4_389 = $signed(_T_68839); // @[Modules.scala 160:64:@15119.4]
  assign buffer_4_181 = {{8{_T_67749[5]}},_T_67749}; // @[Modules.scala 112:22:@8.4]
  assign _T_68841 = $signed(buffer_2_193) + $signed(buffer_4_181); // @[Modules.scala 160:64:@15121.4]
  assign _T_68842 = _T_68841[13:0]; // @[Modules.scala 160:64:@15122.4]
  assign buffer_4_390 = $signed(_T_68842); // @[Modules.scala 160:64:@15123.4]
  assign buffer_4_182 = {{8{_T_67756[5]}},_T_67756}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_183 = {{8{_T_67763[5]}},_T_67763}; // @[Modules.scala 112:22:@8.4]
  assign _T_68844 = $signed(buffer_4_182) + $signed(buffer_4_183); // @[Modules.scala 160:64:@15125.4]
  assign _T_68845 = _T_68844[13:0]; // @[Modules.scala 160:64:@15126.4]
  assign buffer_4_391 = $signed(_T_68845); // @[Modules.scala 160:64:@15127.4]
  assign buffer_4_184 = {{8{_T_67770[5]}},_T_67770}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_185 = {{8{_T_67777[5]}},_T_67777}; // @[Modules.scala 112:22:@8.4]
  assign _T_68847 = $signed(buffer_4_184) + $signed(buffer_4_185); // @[Modules.scala 160:64:@15129.4]
  assign _T_68848 = _T_68847[13:0]; // @[Modules.scala 160:64:@15130.4]
  assign buffer_4_392 = $signed(_T_68848); // @[Modules.scala 160:64:@15131.4]
  assign buffer_4_188 = {{8{_T_67798[5]}},_T_67798}; // @[Modules.scala 112:22:@8.4]
  assign _T_68853 = $signed(buffer_4_188) + $signed(buffer_3_205); // @[Modules.scala 160:64:@15137.4]
  assign _T_68854 = _T_68853[13:0]; // @[Modules.scala 160:64:@15138.4]
  assign buffer_4_394 = $signed(_T_68854); // @[Modules.scala 160:64:@15139.4]
  assign buffer_4_191 = {{9{_T_67819[4]}},_T_67819}; // @[Modules.scala 112:22:@8.4]
  assign _T_68856 = $signed(buffer_3_206) + $signed(buffer_4_191); // @[Modules.scala 160:64:@15141.4]
  assign _T_68857 = _T_68856[13:0]; // @[Modules.scala 160:64:@15142.4]
  assign buffer_4_395 = $signed(_T_68857); // @[Modules.scala 160:64:@15143.4]
  assign buffer_4_192 = {{9{_T_67826[4]}},_T_67826}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_193 = {{9{_T_67833[4]}},_T_67833}; // @[Modules.scala 112:22:@8.4]
  assign _T_68859 = $signed(buffer_4_192) + $signed(buffer_4_193); // @[Modules.scala 160:64:@15145.4]
  assign _T_68860 = _T_68859[13:0]; // @[Modules.scala 160:64:@15146.4]
  assign buffer_4_396 = $signed(_T_68860); // @[Modules.scala 160:64:@15147.4]
  assign buffer_4_195 = {{8{_T_67847[5]}},_T_67847}; // @[Modules.scala 112:22:@8.4]
  assign _T_68862 = $signed(buffer_0_200) + $signed(buffer_4_195); // @[Modules.scala 160:64:@15149.4]
  assign _T_68863 = _T_68862[13:0]; // @[Modules.scala 160:64:@15150.4]
  assign buffer_4_397 = $signed(_T_68863); // @[Modules.scala 160:64:@15151.4]
  assign buffer_4_199 = {{8{_T_67875[5]}},_T_67875}; // @[Modules.scala 112:22:@8.4]
  assign _T_68868 = $signed(buffer_0_206) + $signed(buffer_4_199); // @[Modules.scala 160:64:@15157.4]
  assign _T_68869 = _T_68868[13:0]; // @[Modules.scala 160:64:@15158.4]
  assign buffer_4_399 = $signed(_T_68869); // @[Modules.scala 160:64:@15159.4]
  assign _T_68871 = $signed(buffer_2_213) + $signed(buffer_1_209); // @[Modules.scala 160:64:@15161.4]
  assign _T_68872 = _T_68871[13:0]; // @[Modules.scala 160:64:@15162.4]
  assign buffer_4_400 = $signed(_T_68872); // @[Modules.scala 160:64:@15163.4]
  assign buffer_4_203 = {{9{_T_67903[4]}},_T_67903}; // @[Modules.scala 112:22:@8.4]
  assign _T_68874 = $signed(buffer_2_215) + $signed(buffer_4_203); // @[Modules.scala 160:64:@15165.4]
  assign _T_68875 = _T_68874[13:0]; // @[Modules.scala 160:64:@15166.4]
  assign buffer_4_401 = $signed(_T_68875); // @[Modules.scala 160:64:@15167.4]
  assign buffer_4_204 = {{8{_T_67910[5]}},_T_67910}; // @[Modules.scala 112:22:@8.4]
  assign _T_68877 = $signed(buffer_4_204) + $signed(buffer_3_223); // @[Modules.scala 160:64:@15169.4]
  assign _T_68878 = _T_68877[13:0]; // @[Modules.scala 160:64:@15170.4]
  assign buffer_4_402 = $signed(_T_68878); // @[Modules.scala 160:64:@15171.4]
  assign buffer_4_207 = {{9{_T_67931[4]}},_T_67931}; // @[Modules.scala 112:22:@8.4]
  assign _T_68880 = $signed(buffer_1_214) + $signed(buffer_4_207); // @[Modules.scala 160:64:@15173.4]
  assign _T_68881 = _T_68880[13:0]; // @[Modules.scala 160:64:@15174.4]
  assign buffer_4_403 = $signed(_T_68881); // @[Modules.scala 160:64:@15175.4]
  assign buffer_4_209 = {{9{_T_67945[4]}},_T_67945}; // @[Modules.scala 112:22:@8.4]
  assign _T_68883 = $signed(buffer_3_226) + $signed(buffer_4_209); // @[Modules.scala 160:64:@15177.4]
  assign _T_68884 = _T_68883[13:0]; // @[Modules.scala 160:64:@15178.4]
  assign buffer_4_404 = $signed(_T_68884); // @[Modules.scala 160:64:@15179.4]
  assign buffer_4_210 = {{8{_T_67952[5]}},_T_67952}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_211 = {{8{_T_67959[5]}},_T_67959}; // @[Modules.scala 112:22:@8.4]
  assign _T_68886 = $signed(buffer_4_210) + $signed(buffer_4_211); // @[Modules.scala 160:64:@15181.4]
  assign _T_68887 = _T_68886[13:0]; // @[Modules.scala 160:64:@15182.4]
  assign buffer_4_405 = $signed(_T_68887); // @[Modules.scala 160:64:@15183.4]
  assign buffer_4_216 = {{8{_T_67994[5]}},_T_67994}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_217 = {{9{_T_68001[4]}},_T_68001}; // @[Modules.scala 112:22:@8.4]
  assign _T_68895 = $signed(buffer_4_216) + $signed(buffer_4_217); // @[Modules.scala 160:64:@15193.4]
  assign _T_68896 = _T_68895[13:0]; // @[Modules.scala 160:64:@15194.4]
  assign buffer_4_408 = $signed(_T_68896); // @[Modules.scala 160:64:@15195.4]
  assign buffer_4_218 = {{9{_T_68008[4]}},_T_68008}; // @[Modules.scala 112:22:@8.4]
  assign _T_68898 = $signed(buffer_4_218) + $signed(buffer_1_226); // @[Modules.scala 160:64:@15197.4]
  assign _T_68899 = _T_68898[13:0]; // @[Modules.scala 160:64:@15198.4]
  assign buffer_4_409 = $signed(_T_68899); // @[Modules.scala 160:64:@15199.4]
  assign buffer_4_220 = {{8{_T_68022[5]}},_T_68022}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_221 = {{8{_T_68029[5]}},_T_68029}; // @[Modules.scala 112:22:@8.4]
  assign _T_68901 = $signed(buffer_4_220) + $signed(buffer_4_221); // @[Modules.scala 160:64:@15201.4]
  assign _T_68902 = _T_68901[13:0]; // @[Modules.scala 160:64:@15202.4]
  assign buffer_4_410 = $signed(_T_68902); // @[Modules.scala 160:64:@15203.4]
  assign buffer_4_222 = {{8{_T_68036[5]}},_T_68036}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_223 = {{9{_T_68043[4]}},_T_68043}; // @[Modules.scala 112:22:@8.4]
  assign _T_68904 = $signed(buffer_4_222) + $signed(buffer_4_223); // @[Modules.scala 160:64:@15205.4]
  assign _T_68905 = _T_68904[13:0]; // @[Modules.scala 160:64:@15206.4]
  assign buffer_4_411 = $signed(_T_68905); // @[Modules.scala 160:64:@15207.4]
  assign buffer_4_227 = {{8{_T_68071[5]}},_T_68071}; // @[Modules.scala 112:22:@8.4]
  assign _T_68910 = $signed(buffer_2_238) + $signed(buffer_4_227); // @[Modules.scala 160:64:@15213.4]
  assign _T_68911 = _T_68910[13:0]; // @[Modules.scala 160:64:@15214.4]
  assign buffer_4_413 = $signed(_T_68911); // @[Modules.scala 160:64:@15215.4]
  assign buffer_4_228 = {{9{_T_68078[4]}},_T_68078}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_229 = {{9{_T_68085[4]}},_T_68085}; // @[Modules.scala 112:22:@8.4]
  assign _T_68913 = $signed(buffer_4_228) + $signed(buffer_4_229); // @[Modules.scala 160:64:@15217.4]
  assign _T_68914 = _T_68913[13:0]; // @[Modules.scala 160:64:@15218.4]
  assign buffer_4_414 = $signed(_T_68914); // @[Modules.scala 160:64:@15219.4]
  assign buffer_4_230 = {{9{_T_68092[4]}},_T_68092}; // @[Modules.scala 112:22:@8.4]
  assign _T_68916 = $signed(buffer_4_230) + $signed(buffer_1_237); // @[Modules.scala 160:64:@15221.4]
  assign _T_68917 = _T_68916[13:0]; // @[Modules.scala 160:64:@15222.4]
  assign buffer_4_415 = $signed(_T_68917); // @[Modules.scala 160:64:@15223.4]
  assign buffer_4_233 = {{9{_T_68113[4]}},_T_68113}; // @[Modules.scala 112:22:@8.4]
  assign _T_68919 = $signed(buffer_0_236) + $signed(buffer_4_233); // @[Modules.scala 160:64:@15225.4]
  assign _T_68920 = _T_68919[13:0]; // @[Modules.scala 160:64:@15226.4]
  assign buffer_4_416 = $signed(_T_68920); // @[Modules.scala 160:64:@15227.4]
  assign buffer_4_234 = {{9{_T_68120[4]}},_T_68120}; // @[Modules.scala 112:22:@8.4]
  assign _T_68922 = $signed(buffer_4_234) + $signed(buffer_3_249); // @[Modules.scala 160:64:@15229.4]
  assign _T_68923 = _T_68922[13:0]; // @[Modules.scala 160:64:@15230.4]
  assign buffer_4_417 = $signed(_T_68923); // @[Modules.scala 160:64:@15231.4]
  assign buffer_4_239 = {{9{_T_68155[4]}},_T_68155}; // @[Modules.scala 112:22:@8.4]
  assign _T_68928 = $signed(buffer_2_251) + $signed(buffer_4_239); // @[Modules.scala 160:64:@15237.4]
  assign _T_68929 = _T_68928[13:0]; // @[Modules.scala 160:64:@15238.4]
  assign buffer_4_419 = $signed(_T_68929); // @[Modules.scala 160:64:@15239.4]
  assign _T_68931 = $signed(buffer_2_252) + $signed(buffer_0_245); // @[Modules.scala 160:64:@15241.4]
  assign _T_68932 = _T_68931[13:0]; // @[Modules.scala 160:64:@15242.4]
  assign buffer_4_420 = $signed(_T_68932); // @[Modules.scala 160:64:@15243.4]
  assign buffer_4_242 = {{9{_T_68176[4]}},_T_68176}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_243 = {{9{_T_68183[4]}},_T_68183}; // @[Modules.scala 112:22:@8.4]
  assign _T_68934 = $signed(buffer_4_242) + $signed(buffer_4_243); // @[Modules.scala 160:64:@15245.4]
  assign _T_68935 = _T_68934[13:0]; // @[Modules.scala 160:64:@15246.4]
  assign buffer_4_421 = $signed(_T_68935); // @[Modules.scala 160:64:@15247.4]
  assign buffer_4_244 = {{8{_T_68190[5]}},_T_68190}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_245 = {{8{_T_68197[5]}},_T_68197}; // @[Modules.scala 112:22:@8.4]
  assign _T_68937 = $signed(buffer_4_244) + $signed(buffer_4_245); // @[Modules.scala 160:64:@15249.4]
  assign _T_68938 = _T_68937[13:0]; // @[Modules.scala 160:64:@15250.4]
  assign buffer_4_422 = $signed(_T_68938); // @[Modules.scala 160:64:@15251.4]
  assign buffer_4_246 = {{9{_T_68204[4]}},_T_68204}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_247 = {{9{_T_68211[4]}},_T_68211}; // @[Modules.scala 112:22:@8.4]
  assign _T_68940 = $signed(buffer_4_246) + $signed(buffer_4_247); // @[Modules.scala 160:64:@15253.4]
  assign _T_68941 = _T_68940[13:0]; // @[Modules.scala 160:64:@15254.4]
  assign buffer_4_423 = $signed(_T_68941); // @[Modules.scala 160:64:@15255.4]
  assign buffer_4_248 = {{8{_T_68218[5]}},_T_68218}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_249 = {{8{_T_68225[5]}},_T_68225}; // @[Modules.scala 112:22:@8.4]
  assign _T_68943 = $signed(buffer_4_248) + $signed(buffer_4_249); // @[Modules.scala 160:64:@15257.4]
  assign _T_68944 = _T_68943[13:0]; // @[Modules.scala 160:64:@15258.4]
  assign buffer_4_424 = $signed(_T_68944); // @[Modules.scala 160:64:@15259.4]
  assign buffer_4_252 = {{8{_T_68246[5]}},_T_68246}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_253 = {{9{_T_68253[4]}},_T_68253}; // @[Modules.scala 112:22:@8.4]
  assign _T_68949 = $signed(buffer_4_252) + $signed(buffer_4_253); // @[Modules.scala 160:64:@15265.4]
  assign _T_68950 = _T_68949[13:0]; // @[Modules.scala 160:64:@15266.4]
  assign buffer_4_426 = $signed(_T_68950); // @[Modules.scala 160:64:@15267.4]
  assign buffer_4_254 = {{8{_T_68260[5]}},_T_68260}; // @[Modules.scala 112:22:@8.4]
  assign _T_68952 = $signed(buffer_4_254) + $signed(buffer_3_269); // @[Modules.scala 160:64:@15269.4]
  assign _T_68953 = _T_68952[13:0]; // @[Modules.scala 160:64:@15270.4]
  assign buffer_4_427 = $signed(_T_68953); // @[Modules.scala 160:64:@15271.4]
  assign buffer_4_257 = {{8{_T_68281[5]}},_T_68281}; // @[Modules.scala 112:22:@8.4]
  assign _T_68955 = $signed(buffer_3_270) + $signed(buffer_4_257); // @[Modules.scala 160:64:@15273.4]
  assign _T_68956 = _T_68955[13:0]; // @[Modules.scala 160:64:@15274.4]
  assign buffer_4_428 = $signed(_T_68956); // @[Modules.scala 160:64:@15275.4]
  assign buffer_4_258 = {{8{_T_68288[5]}},_T_68288}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_259 = {{9{_T_68295[4]}},_T_68295}; // @[Modules.scala 112:22:@8.4]
  assign _T_68958 = $signed(buffer_4_258) + $signed(buffer_4_259); // @[Modules.scala 160:64:@15277.4]
  assign _T_68959 = _T_68958[13:0]; // @[Modules.scala 160:64:@15278.4]
  assign buffer_4_429 = $signed(_T_68959); // @[Modules.scala 160:64:@15279.4]
  assign buffer_4_260 = {{9{_T_68302[4]}},_T_68302}; // @[Modules.scala 112:22:@8.4]
  assign _T_68961 = $signed(buffer_4_260) + $signed(buffer_0_266); // @[Modules.scala 160:64:@15281.4]
  assign _T_68962 = _T_68961[13:0]; // @[Modules.scala 160:64:@15282.4]
  assign buffer_4_430 = $signed(_T_68962); // @[Modules.scala 160:64:@15283.4]
  assign buffer_4_263 = {{8{_T_68323[5]}},_T_68323}; // @[Modules.scala 112:22:@8.4]
  assign _T_68964 = $signed(buffer_0_267) + $signed(buffer_4_263); // @[Modules.scala 160:64:@15285.4]
  assign _T_68965 = _T_68964[13:0]; // @[Modules.scala 160:64:@15286.4]
  assign buffer_4_431 = $signed(_T_68965); // @[Modules.scala 160:64:@15287.4]
  assign buffer_4_265 = {{8{_T_68337[5]}},_T_68337}; // @[Modules.scala 112:22:@8.4]
  assign _T_68967 = $signed(buffer_2_277) + $signed(buffer_4_265); // @[Modules.scala 160:64:@15289.4]
  assign _T_68968 = _T_68967[13:0]; // @[Modules.scala 160:64:@15290.4]
  assign buffer_4_432 = $signed(_T_68968); // @[Modules.scala 160:64:@15291.4]
  assign buffer_4_266 = {{9{_T_68344[4]}},_T_68344}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_267 = {{9{_T_68351[4]}},_T_68351}; // @[Modules.scala 112:22:@8.4]
  assign _T_68970 = $signed(buffer_4_266) + $signed(buffer_4_267); // @[Modules.scala 160:64:@15293.4]
  assign _T_68971 = _T_68970[13:0]; // @[Modules.scala 160:64:@15294.4]
  assign buffer_4_433 = $signed(_T_68971); // @[Modules.scala 160:64:@15295.4]
  assign buffer_4_268 = {{8{_T_68358[5]}},_T_68358}; // @[Modules.scala 112:22:@8.4]
  assign _T_68973 = $signed(buffer_4_268) + $signed(buffer_1_274); // @[Modules.scala 160:64:@15297.4]
  assign _T_68974 = _T_68973[13:0]; // @[Modules.scala 160:64:@15298.4]
  assign buffer_4_434 = $signed(_T_68974); // @[Modules.scala 160:64:@15299.4]
  assign _T_68976 = $signed(buffer_1_275) + $signed(buffer_1_276); // @[Modules.scala 160:64:@15301.4]
  assign _T_68977 = _T_68976[13:0]; // @[Modules.scala 160:64:@15302.4]
  assign buffer_4_435 = $signed(_T_68977); // @[Modules.scala 160:64:@15303.4]
  assign _T_68979 = $signed(buffer_1_277) + $signed(buffer_1_278); // @[Modules.scala 160:64:@15305.4]
  assign _T_68980 = _T_68979[13:0]; // @[Modules.scala 160:64:@15306.4]
  assign buffer_4_436 = $signed(_T_68980); // @[Modules.scala 160:64:@15307.4]
  assign _T_68982 = $signed(buffer_1_279) + $signed(buffer_1_280); // @[Modules.scala 160:64:@15309.4]
  assign _T_68983 = _T_68982[13:0]; // @[Modules.scala 160:64:@15310.4]
  assign buffer_4_437 = $signed(_T_68983); // @[Modules.scala 160:64:@15311.4]
  assign buffer_4_278 = {{8{_T_68428[5]}},_T_68428}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_279 = {{8{_T_68435[5]}},_T_68435}; // @[Modules.scala 112:22:@8.4]
  assign _T_68988 = $signed(buffer_4_278) + $signed(buffer_4_279); // @[Modules.scala 160:64:@15317.4]
  assign _T_68989 = _T_68988[13:0]; // @[Modules.scala 160:64:@15318.4]
  assign buffer_4_439 = $signed(_T_68989); // @[Modules.scala 160:64:@15319.4]
  assign buffer_4_281 = {{8{_T_68449[5]}},_T_68449}; // @[Modules.scala 112:22:@8.4]
  assign _T_68991 = $signed(buffer_3_294) + $signed(buffer_4_281); // @[Modules.scala 160:64:@15321.4]
  assign _T_68992 = _T_68991[13:0]; // @[Modules.scala 160:64:@15322.4]
  assign buffer_4_440 = $signed(_T_68992); // @[Modules.scala 160:64:@15323.4]
  assign buffer_4_282 = {{8{_T_68456[5]}},_T_68456}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_283 = {{8{_T_68463[5]}},_T_68463}; // @[Modules.scala 112:22:@8.4]
  assign _T_68994 = $signed(buffer_4_282) + $signed(buffer_4_283); // @[Modules.scala 160:64:@15325.4]
  assign _T_68995 = _T_68994[13:0]; // @[Modules.scala 160:64:@15326.4]
  assign buffer_4_441 = $signed(_T_68995); // @[Modules.scala 160:64:@15327.4]
  assign buffer_4_284 = {{8{_T_68470[5]}},_T_68470}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_285 = {{8{_T_68477[5]}},_T_68477}; // @[Modules.scala 112:22:@8.4]
  assign _T_68997 = $signed(buffer_4_284) + $signed(buffer_4_285); // @[Modules.scala 160:64:@15329.4]
  assign _T_68998 = _T_68997[13:0]; // @[Modules.scala 160:64:@15330.4]
  assign buffer_4_442 = $signed(_T_68998); // @[Modules.scala 160:64:@15331.4]
  assign buffer_4_286 = {{8{_T_68484[5]}},_T_68484}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_287 = {{8{_T_68491[5]}},_T_68491}; // @[Modules.scala 112:22:@8.4]
  assign _T_69000 = $signed(buffer_4_286) + $signed(buffer_4_287); // @[Modules.scala 160:64:@15333.4]
  assign _T_69001 = _T_69000[13:0]; // @[Modules.scala 160:64:@15334.4]
  assign buffer_4_443 = $signed(_T_69001); // @[Modules.scala 160:64:@15335.4]
  assign buffer_4_288 = {{8{_T_68498[5]}},_T_68498}; // @[Modules.scala 112:22:@8.4]
  assign buffer_4_289 = {{8{_T_68505[5]}},_T_68505}; // @[Modules.scala 112:22:@8.4]
  assign _T_69003 = $signed(buffer_4_288) + $signed(buffer_4_289); // @[Modules.scala 160:64:@15337.4]
  assign _T_69004 = _T_69003[13:0]; // @[Modules.scala 160:64:@15338.4]
  assign buffer_4_444 = $signed(_T_69004); // @[Modules.scala 160:64:@15339.4]
  assign _T_69006 = $signed(buffer_1_293) + $signed(buffer_3_304); // @[Modules.scala 160:64:@15341.4]
  assign _T_69007 = _T_69006[13:0]; // @[Modules.scala 160:64:@15342.4]
  assign buffer_4_445 = $signed(_T_69007); // @[Modules.scala 160:64:@15343.4]
  assign buffer_4_292 = {{8{_T_68526[5]}},_T_68526}; // @[Modules.scala 112:22:@8.4]
  assign _T_69009 = $signed(buffer_4_292) + $signed(buffer_0_295); // @[Modules.scala 160:64:@15345.4]
  assign _T_69010 = _T_69009[13:0]; // @[Modules.scala 160:64:@15346.4]
  assign buffer_4_446 = $signed(_T_69010); // @[Modules.scala 160:64:@15347.4]
  assign buffer_4_296 = {{8{_T_68554[5]}},_T_68554}; // @[Modules.scala 112:22:@8.4]
  assign _T_69015 = $signed(buffer_4_296) + $signed(buffer_1_301); // @[Modules.scala 160:64:@15353.4]
  assign _T_69016 = _T_69015[13:0]; // @[Modules.scala 160:64:@15354.4]
  assign buffer_4_448 = $signed(_T_69016); // @[Modules.scala 160:64:@15355.4]
  assign _T_69021 = $signed(buffer_0_302) + $signed(buffer_4_301); // @[Modules.scala 160:64:@15361.4]
  assign _T_69022 = _T_69021[13:0]; // @[Modules.scala 160:64:@15362.4]
  assign buffer_4_450 = $signed(_T_69022); // @[Modules.scala 160:64:@15363.4]
  assign _T_69024 = $signed(buffer_4_302) + $signed(buffer_4_303); // @[Modules.scala 160:64:@15365.4]
  assign _T_69025 = _T_69024[13:0]; // @[Modules.scala 160:64:@15366.4]
  assign buffer_4_451 = $signed(_T_69025); // @[Modules.scala 160:64:@15367.4]
  assign _T_69027 = $signed(buffer_4_304) + $signed(buffer_4_305); // @[Modules.scala 160:64:@15369.4]
  assign _T_69028 = _T_69027[13:0]; // @[Modules.scala 160:64:@15370.4]
  assign buffer_4_452 = $signed(_T_69028); // @[Modules.scala 160:64:@15371.4]
  assign _T_69030 = $signed(buffer_4_306) + $signed(buffer_2_317); // @[Modules.scala 160:64:@15373.4]
  assign _T_69031 = _T_69030[13:0]; // @[Modules.scala 160:64:@15374.4]
  assign buffer_4_453 = $signed(_T_69031); // @[Modules.scala 160:64:@15375.4]
  assign _T_69033 = $signed(buffer_4_308) + $signed(buffer_4_309); // @[Modules.scala 160:64:@15377.4]
  assign _T_69034 = _T_69033[13:0]; // @[Modules.scala 160:64:@15378.4]
  assign buffer_4_454 = $signed(_T_69034); // @[Modules.scala 160:64:@15379.4]
  assign _T_69036 = $signed(buffer_4_310) + $signed(buffer_4_311); // @[Modules.scala 160:64:@15381.4]
  assign _T_69037 = _T_69036[13:0]; // @[Modules.scala 160:64:@15382.4]
  assign buffer_4_455 = $signed(_T_69037); // @[Modules.scala 160:64:@15383.4]
  assign _T_69039 = $signed(buffer_4_312) + $signed(buffer_4_313); // @[Modules.scala 160:64:@15385.4]
  assign _T_69040 = _T_69039[13:0]; // @[Modules.scala 160:64:@15386.4]
  assign buffer_4_456 = $signed(_T_69040); // @[Modules.scala 160:64:@15387.4]
  assign _T_69042 = $signed(buffer_4_314) + $signed(buffer_4_315); // @[Modules.scala 160:64:@15389.4]
  assign _T_69043 = _T_69042[13:0]; // @[Modules.scala 160:64:@15390.4]
  assign buffer_4_457 = $signed(_T_69043); // @[Modules.scala 160:64:@15391.4]
  assign _T_69045 = $signed(buffer_4_316) + $signed(buffer_4_317); // @[Modules.scala 160:64:@15393.4]
  assign _T_69046 = _T_69045[13:0]; // @[Modules.scala 160:64:@15394.4]
  assign buffer_4_458 = $signed(_T_69046); // @[Modules.scala 160:64:@15395.4]
  assign _T_69048 = $signed(buffer_4_318) + $signed(buffer_4_319); // @[Modules.scala 160:64:@15397.4]
  assign _T_69049 = _T_69048[13:0]; // @[Modules.scala 160:64:@15398.4]
  assign buffer_4_459 = $signed(_T_69049); // @[Modules.scala 160:64:@15399.4]
  assign _T_69051 = $signed(buffer_4_320) + $signed(buffer_4_321); // @[Modules.scala 160:64:@15401.4]
  assign _T_69052 = _T_69051[13:0]; // @[Modules.scala 160:64:@15402.4]
  assign buffer_4_460 = $signed(_T_69052); // @[Modules.scala 160:64:@15403.4]
  assign _T_69054 = $signed(buffer_4_322) + $signed(buffer_3_338); // @[Modules.scala 160:64:@15405.4]
  assign _T_69055 = _T_69054[13:0]; // @[Modules.scala 160:64:@15406.4]
  assign buffer_4_461 = $signed(_T_69055); // @[Modules.scala 160:64:@15407.4]
  assign _T_69057 = $signed(buffer_4_324) + $signed(buffer_3_340); // @[Modules.scala 160:64:@15409.4]
  assign _T_69058 = _T_69057[13:0]; // @[Modules.scala 160:64:@15410.4]
  assign buffer_4_462 = $signed(_T_69058); // @[Modules.scala 160:64:@15411.4]
  assign _T_69060 = $signed(buffer_4_326) + $signed(buffer_4_327); // @[Modules.scala 160:64:@15413.4]
  assign _T_69061 = _T_69060[13:0]; // @[Modules.scala 160:64:@15414.4]
  assign buffer_4_463 = $signed(_T_69061); // @[Modules.scala 160:64:@15415.4]
  assign _T_69063 = $signed(buffer_4_328) + $signed(buffer_3_344); // @[Modules.scala 160:64:@15417.4]
  assign _T_69064 = _T_69063[13:0]; // @[Modules.scala 160:64:@15418.4]
  assign buffer_4_464 = $signed(_T_69064); // @[Modules.scala 160:64:@15419.4]
  assign _T_69066 = $signed(buffer_4_330) + $signed(buffer_4_331); // @[Modules.scala 160:64:@15421.4]
  assign _T_69067 = _T_69066[13:0]; // @[Modules.scala 160:64:@15422.4]
  assign buffer_4_465 = $signed(_T_69067); // @[Modules.scala 160:64:@15423.4]
  assign _T_69069 = $signed(buffer_4_332) + $signed(buffer_4_333); // @[Modules.scala 160:64:@15425.4]
  assign _T_69070 = _T_69069[13:0]; // @[Modules.scala 160:64:@15426.4]
  assign buffer_4_466 = $signed(_T_69070); // @[Modules.scala 160:64:@15427.4]
  assign _T_69072 = $signed(buffer_0_335) + $signed(buffer_4_335); // @[Modules.scala 160:64:@15429.4]
  assign _T_69073 = _T_69072[13:0]; // @[Modules.scala 160:64:@15430.4]
  assign buffer_4_467 = $signed(_T_69073); // @[Modules.scala 160:64:@15431.4]
  assign _T_69075 = $signed(buffer_4_336) + $signed(buffer_4_337); // @[Modules.scala 160:64:@15433.4]
  assign _T_69076 = _T_69075[13:0]; // @[Modules.scala 160:64:@15434.4]
  assign buffer_4_468 = $signed(_T_69076); // @[Modules.scala 160:64:@15435.4]
  assign _T_69078 = $signed(buffer_1_342) + $signed(buffer_4_339); // @[Modules.scala 160:64:@15437.4]
  assign _T_69079 = _T_69078[13:0]; // @[Modules.scala 160:64:@15438.4]
  assign buffer_4_469 = $signed(_T_69079); // @[Modules.scala 160:64:@15439.4]
  assign _T_69081 = $signed(buffer_4_340) + $signed(buffer_4_341); // @[Modules.scala 160:64:@15441.4]
  assign _T_69082 = _T_69081[13:0]; // @[Modules.scala 160:64:@15442.4]
  assign buffer_4_470 = $signed(_T_69082); // @[Modules.scala 160:64:@15443.4]
  assign _T_69084 = $signed(buffer_4_342) + $signed(buffer_2_354); // @[Modules.scala 160:64:@15445.4]
  assign _T_69085 = _T_69084[13:0]; // @[Modules.scala 160:64:@15446.4]
  assign buffer_4_471 = $signed(_T_69085); // @[Modules.scala 160:64:@15447.4]
  assign _T_69087 = $signed(buffer_2_355) + $signed(buffer_4_345); // @[Modules.scala 160:64:@15449.4]
  assign _T_69088 = _T_69087[13:0]; // @[Modules.scala 160:64:@15450.4]
  assign buffer_4_472 = $signed(_T_69088); // @[Modules.scala 160:64:@15451.4]
  assign _T_69090 = $signed(buffer_4_346) + $signed(buffer_4_347); // @[Modules.scala 160:64:@15453.4]
  assign _T_69091 = _T_69090[13:0]; // @[Modules.scala 160:64:@15454.4]
  assign buffer_4_473 = $signed(_T_69091); // @[Modules.scala 160:64:@15455.4]
  assign _T_69093 = $signed(buffer_4_348) + $signed(buffer_0_350); // @[Modules.scala 160:64:@15457.4]
  assign _T_69094 = _T_69093[13:0]; // @[Modules.scala 160:64:@15458.4]
  assign buffer_4_474 = $signed(_T_69094); // @[Modules.scala 160:64:@15459.4]
  assign _T_69096 = $signed(buffer_4_350) + $signed(buffer_4_351); // @[Modules.scala 160:64:@15461.4]
  assign _T_69097 = _T_69096[13:0]; // @[Modules.scala 160:64:@15462.4]
  assign buffer_4_475 = $signed(_T_69097); // @[Modules.scala 160:64:@15463.4]
  assign _T_69099 = $signed(buffer_4_352) + $signed(buffer_4_353); // @[Modules.scala 160:64:@15465.4]
  assign _T_69100 = _T_69099[13:0]; // @[Modules.scala 160:64:@15466.4]
  assign buffer_4_476 = $signed(_T_69100); // @[Modules.scala 160:64:@15467.4]
  assign _T_69102 = $signed(buffer_4_354) + $signed(buffer_4_355); // @[Modules.scala 160:64:@15469.4]
  assign _T_69103 = _T_69102[13:0]; // @[Modules.scala 160:64:@15470.4]
  assign buffer_4_477 = $signed(_T_69103); // @[Modules.scala 160:64:@15471.4]
  assign _T_69105 = $signed(buffer_4_356) + $signed(buffer_4_357); // @[Modules.scala 160:64:@15473.4]
  assign _T_69106 = _T_69105[13:0]; // @[Modules.scala 160:64:@15474.4]
  assign buffer_4_478 = $signed(_T_69106); // @[Modules.scala 160:64:@15475.4]
  assign _T_69108 = $signed(buffer_4_358) + $signed(buffer_4_359); // @[Modules.scala 160:64:@15477.4]
  assign _T_69109 = _T_69108[13:0]; // @[Modules.scala 160:64:@15478.4]
  assign buffer_4_479 = $signed(_T_69109); // @[Modules.scala 160:64:@15479.4]
  assign _T_69111 = $signed(buffer_4_360) + $signed(buffer_4_361); // @[Modules.scala 160:64:@15481.4]
  assign _T_69112 = _T_69111[13:0]; // @[Modules.scala 160:64:@15482.4]
  assign buffer_4_480 = $signed(_T_69112); // @[Modules.scala 160:64:@15483.4]
  assign _T_69114 = $signed(buffer_4_362) + $signed(buffer_4_363); // @[Modules.scala 160:64:@15485.4]
  assign _T_69115 = _T_69114[13:0]; // @[Modules.scala 160:64:@15486.4]
  assign buffer_4_481 = $signed(_T_69115); // @[Modules.scala 160:64:@15487.4]
  assign _T_69117 = $signed(buffer_4_364) + $signed(buffer_4_365); // @[Modules.scala 160:64:@15489.4]
  assign _T_69118 = _T_69117[13:0]; // @[Modules.scala 160:64:@15490.4]
  assign buffer_4_482 = $signed(_T_69118); // @[Modules.scala 160:64:@15491.4]
  assign _T_69120 = $signed(buffer_4_366) + $signed(buffer_4_367); // @[Modules.scala 160:64:@15493.4]
  assign _T_69121 = _T_69120[13:0]; // @[Modules.scala 160:64:@15494.4]
  assign buffer_4_483 = $signed(_T_69121); // @[Modules.scala 160:64:@15495.4]
  assign _T_69123 = $signed(buffer_4_368) + $signed(buffer_4_369); // @[Modules.scala 160:64:@15497.4]
  assign _T_69124 = _T_69123[13:0]; // @[Modules.scala 160:64:@15498.4]
  assign buffer_4_484 = $signed(_T_69124); // @[Modules.scala 160:64:@15499.4]
  assign _T_69126 = $signed(buffer_4_370) + $signed(buffer_4_371); // @[Modules.scala 160:64:@15501.4]
  assign _T_69127 = _T_69126[13:0]; // @[Modules.scala 160:64:@15502.4]
  assign buffer_4_485 = $signed(_T_69127); // @[Modules.scala 160:64:@15503.4]
  assign _T_69129 = $signed(buffer_4_372) + $signed(buffer_4_373); // @[Modules.scala 160:64:@15505.4]
  assign _T_69130 = _T_69129[13:0]; // @[Modules.scala 160:64:@15506.4]
  assign buffer_4_486 = $signed(_T_69130); // @[Modules.scala 160:64:@15507.4]
  assign _T_69132 = $signed(buffer_4_374) + $signed(buffer_4_375); // @[Modules.scala 160:64:@15509.4]
  assign _T_69133 = _T_69132[13:0]; // @[Modules.scala 160:64:@15510.4]
  assign buffer_4_487 = $signed(_T_69133); // @[Modules.scala 160:64:@15511.4]
  assign _T_69135 = $signed(buffer_4_376) + $signed(buffer_4_377); // @[Modules.scala 160:64:@15513.4]
  assign _T_69136 = _T_69135[13:0]; // @[Modules.scala 160:64:@15514.4]
  assign buffer_4_488 = $signed(_T_69136); // @[Modules.scala 160:64:@15515.4]
  assign _T_69138 = $signed(buffer_4_378) + $signed(buffer_4_379); // @[Modules.scala 160:64:@15517.4]
  assign _T_69139 = _T_69138[13:0]; // @[Modules.scala 160:64:@15518.4]
  assign buffer_4_489 = $signed(_T_69139); // @[Modules.scala 160:64:@15519.4]
  assign _T_69141 = $signed(buffer_4_380) + $signed(buffer_4_381); // @[Modules.scala 160:64:@15521.4]
  assign _T_69142 = _T_69141[13:0]; // @[Modules.scala 160:64:@15522.4]
  assign buffer_4_490 = $signed(_T_69142); // @[Modules.scala 160:64:@15523.4]
  assign _T_69144 = $signed(buffer_4_382) + $signed(buffer_4_383); // @[Modules.scala 160:64:@15525.4]
  assign _T_69145 = _T_69144[13:0]; // @[Modules.scala 160:64:@15526.4]
  assign buffer_4_491 = $signed(_T_69145); // @[Modules.scala 160:64:@15527.4]
  assign _T_69147 = $signed(buffer_4_384) + $signed(buffer_4_385); // @[Modules.scala 160:64:@15529.4]
  assign _T_69148 = _T_69147[13:0]; // @[Modules.scala 160:64:@15530.4]
  assign buffer_4_492 = $signed(_T_69148); // @[Modules.scala 160:64:@15531.4]
  assign _T_69150 = $signed(buffer_4_386) + $signed(buffer_4_387); // @[Modules.scala 160:64:@15533.4]
  assign _T_69151 = _T_69150[13:0]; // @[Modules.scala 160:64:@15534.4]
  assign buffer_4_493 = $signed(_T_69151); // @[Modules.scala 160:64:@15535.4]
  assign _T_69153 = $signed(buffer_3_410) + $signed(buffer_4_389); // @[Modules.scala 160:64:@15537.4]
  assign _T_69154 = _T_69153[13:0]; // @[Modules.scala 160:64:@15538.4]
  assign buffer_4_494 = $signed(_T_69154); // @[Modules.scala 160:64:@15539.4]
  assign _T_69156 = $signed(buffer_4_390) + $signed(buffer_4_391); // @[Modules.scala 160:64:@15541.4]
  assign _T_69157 = _T_69156[13:0]; // @[Modules.scala 160:64:@15542.4]
  assign buffer_4_495 = $signed(_T_69157); // @[Modules.scala 160:64:@15543.4]
  assign _T_69159 = $signed(buffer_4_392) + $signed(buffer_3_415); // @[Modules.scala 160:64:@15545.4]
  assign _T_69160 = _T_69159[13:0]; // @[Modules.scala 160:64:@15546.4]
  assign buffer_4_496 = $signed(_T_69160); // @[Modules.scala 160:64:@15547.4]
  assign _T_69162 = $signed(buffer_4_394) + $signed(buffer_4_395); // @[Modules.scala 160:64:@15549.4]
  assign _T_69163 = _T_69162[13:0]; // @[Modules.scala 160:64:@15550.4]
  assign buffer_4_497 = $signed(_T_69163); // @[Modules.scala 160:64:@15551.4]
  assign _T_69165 = $signed(buffer_4_396) + $signed(buffer_4_397); // @[Modules.scala 160:64:@15553.4]
  assign _T_69166 = _T_69165[13:0]; // @[Modules.scala 160:64:@15554.4]
  assign buffer_4_498 = $signed(_T_69166); // @[Modules.scala 160:64:@15555.4]
  assign _T_69168 = $signed(buffer_3_421) + $signed(buffer_4_399); // @[Modules.scala 160:64:@15557.4]
  assign _T_69169 = _T_69168[13:0]; // @[Modules.scala 160:64:@15558.4]
  assign buffer_4_499 = $signed(_T_69169); // @[Modules.scala 160:64:@15559.4]
  assign _T_69171 = $signed(buffer_4_400) + $signed(buffer_4_401); // @[Modules.scala 160:64:@15561.4]
  assign _T_69172 = _T_69171[13:0]; // @[Modules.scala 160:64:@15562.4]
  assign buffer_4_500 = $signed(_T_69172); // @[Modules.scala 160:64:@15563.4]
  assign _T_69174 = $signed(buffer_4_402) + $signed(buffer_4_403); // @[Modules.scala 160:64:@15565.4]
  assign _T_69175 = _T_69174[13:0]; // @[Modules.scala 160:64:@15566.4]
  assign buffer_4_501 = $signed(_T_69175); // @[Modules.scala 160:64:@15567.4]
  assign _T_69177 = $signed(buffer_4_404) + $signed(buffer_4_405); // @[Modules.scala 160:64:@15569.4]
  assign _T_69178 = _T_69177[13:0]; // @[Modules.scala 160:64:@15570.4]
  assign buffer_4_502 = $signed(_T_69178); // @[Modules.scala 160:64:@15571.4]
  assign _T_69183 = $signed(buffer_4_408) + $signed(buffer_4_409); // @[Modules.scala 160:64:@15577.4]
  assign _T_69184 = _T_69183[13:0]; // @[Modules.scala 160:64:@15578.4]
  assign buffer_4_504 = $signed(_T_69184); // @[Modules.scala 160:64:@15579.4]
  assign _T_69186 = $signed(buffer_4_410) + $signed(buffer_4_411); // @[Modules.scala 160:64:@15581.4]
  assign _T_69187 = _T_69186[13:0]; // @[Modules.scala 160:64:@15582.4]
  assign buffer_4_505 = $signed(_T_69187); // @[Modules.scala 160:64:@15583.4]
  assign _T_69189 = $signed(buffer_2_428) + $signed(buffer_4_413); // @[Modules.scala 160:64:@15585.4]
  assign _T_69190 = _T_69189[13:0]; // @[Modules.scala 160:64:@15586.4]
  assign buffer_4_506 = $signed(_T_69190); // @[Modules.scala 160:64:@15587.4]
  assign _T_69192 = $signed(buffer_4_414) + $signed(buffer_4_415); // @[Modules.scala 160:64:@15589.4]
  assign _T_69193 = _T_69192[13:0]; // @[Modules.scala 160:64:@15590.4]
  assign buffer_4_507 = $signed(_T_69193); // @[Modules.scala 160:64:@15591.4]
  assign _T_69195 = $signed(buffer_4_416) + $signed(buffer_4_417); // @[Modules.scala 160:64:@15593.4]
  assign _T_69196 = _T_69195[13:0]; // @[Modules.scala 160:64:@15594.4]
  assign buffer_4_508 = $signed(_T_69196); // @[Modules.scala 160:64:@15595.4]
  assign _T_69198 = $signed(buffer_3_439) + $signed(buffer_4_419); // @[Modules.scala 160:64:@15597.4]
  assign _T_69199 = _T_69198[13:0]; // @[Modules.scala 160:64:@15598.4]
  assign buffer_4_509 = $signed(_T_69199); // @[Modules.scala 160:64:@15599.4]
  assign _T_69201 = $signed(buffer_4_420) + $signed(buffer_4_421); // @[Modules.scala 160:64:@15601.4]
  assign _T_69202 = _T_69201[13:0]; // @[Modules.scala 160:64:@15602.4]
  assign buffer_4_510 = $signed(_T_69202); // @[Modules.scala 160:64:@15603.4]
  assign _T_69204 = $signed(buffer_4_422) + $signed(buffer_4_423); // @[Modules.scala 160:64:@15605.4]
  assign _T_69205 = _T_69204[13:0]; // @[Modules.scala 160:64:@15606.4]
  assign buffer_4_511 = $signed(_T_69205); // @[Modules.scala 160:64:@15607.4]
  assign _T_69207 = $signed(buffer_4_424) + $signed(buffer_2_441); // @[Modules.scala 160:64:@15609.4]
  assign _T_69208 = _T_69207[13:0]; // @[Modules.scala 160:64:@15610.4]
  assign buffer_4_512 = $signed(_T_69208); // @[Modules.scala 160:64:@15611.4]
  assign _T_69210 = $signed(buffer_4_426) + $signed(buffer_4_427); // @[Modules.scala 160:64:@15613.4]
  assign _T_69211 = _T_69210[13:0]; // @[Modules.scala 160:64:@15614.4]
  assign buffer_4_513 = $signed(_T_69211); // @[Modules.scala 160:64:@15615.4]
  assign _T_69213 = $signed(buffer_4_428) + $signed(buffer_4_429); // @[Modules.scala 160:64:@15617.4]
  assign _T_69214 = _T_69213[13:0]; // @[Modules.scala 160:64:@15618.4]
  assign buffer_4_514 = $signed(_T_69214); // @[Modules.scala 160:64:@15619.4]
  assign _T_69216 = $signed(buffer_4_430) + $signed(buffer_4_431); // @[Modules.scala 160:64:@15621.4]
  assign _T_69217 = _T_69216[13:0]; // @[Modules.scala 160:64:@15622.4]
  assign buffer_4_515 = $signed(_T_69217); // @[Modules.scala 160:64:@15623.4]
  assign _T_69219 = $signed(buffer_4_432) + $signed(buffer_4_433); // @[Modules.scala 160:64:@15625.4]
  assign _T_69220 = _T_69219[13:0]; // @[Modules.scala 160:64:@15626.4]
  assign buffer_4_516 = $signed(_T_69220); // @[Modules.scala 160:64:@15627.4]
  assign _T_69222 = $signed(buffer_4_434) + $signed(buffer_4_435); // @[Modules.scala 160:64:@15629.4]
  assign _T_69223 = _T_69222[13:0]; // @[Modules.scala 160:64:@15630.4]
  assign buffer_4_517 = $signed(_T_69223); // @[Modules.scala 160:64:@15631.4]
  assign _T_69225 = $signed(buffer_4_436) + $signed(buffer_4_437); // @[Modules.scala 160:64:@15633.4]
  assign _T_69226 = _T_69225[13:0]; // @[Modules.scala 160:64:@15634.4]
  assign buffer_4_518 = $signed(_T_69226); // @[Modules.scala 160:64:@15635.4]
  assign _T_69228 = $signed(buffer_3_459) + $signed(buffer_4_439); // @[Modules.scala 160:64:@15637.4]
  assign _T_69229 = _T_69228[13:0]; // @[Modules.scala 160:64:@15638.4]
  assign buffer_4_519 = $signed(_T_69229); // @[Modules.scala 160:64:@15639.4]
  assign _T_69231 = $signed(buffer_4_440) + $signed(buffer_4_441); // @[Modules.scala 160:64:@15641.4]
  assign _T_69232 = _T_69231[13:0]; // @[Modules.scala 160:64:@15642.4]
  assign buffer_4_520 = $signed(_T_69232); // @[Modules.scala 160:64:@15643.4]
  assign _T_69234 = $signed(buffer_4_442) + $signed(buffer_4_443); // @[Modules.scala 160:64:@15645.4]
  assign _T_69235 = _T_69234[13:0]; // @[Modules.scala 160:64:@15646.4]
  assign buffer_4_521 = $signed(_T_69235); // @[Modules.scala 160:64:@15647.4]
  assign _T_69237 = $signed(buffer_4_444) + $signed(buffer_4_445); // @[Modules.scala 160:64:@15649.4]
  assign _T_69238 = _T_69237[13:0]; // @[Modules.scala 160:64:@15650.4]
  assign buffer_4_522 = $signed(_T_69238); // @[Modules.scala 160:64:@15651.4]
  assign _T_69240 = $signed(buffer_4_446) + $signed(buffer_1_453); // @[Modules.scala 160:64:@15653.4]
  assign _T_69241 = _T_69240[13:0]; // @[Modules.scala 160:64:@15654.4]
  assign buffer_4_523 = $signed(_T_69241); // @[Modules.scala 160:64:@15655.4]
  assign _T_69243 = $signed(buffer_4_448) + $signed(buffer_0_452); // @[Modules.scala 160:64:@15657.4]
  assign _T_69244 = _T_69243[13:0]; // @[Modules.scala 160:64:@15658.4]
  assign buffer_4_524 = $signed(_T_69244); // @[Modules.scala 160:64:@15659.4]
  assign _T_69246 = $signed(buffer_4_450) + $signed(buffer_4_451); // @[Modules.scala 166:64:@15661.4]
  assign _T_69247 = _T_69246[13:0]; // @[Modules.scala 166:64:@15662.4]
  assign buffer_4_525 = $signed(_T_69247); // @[Modules.scala 166:64:@15663.4]
  assign _T_69249 = $signed(buffer_4_452) + $signed(buffer_4_453); // @[Modules.scala 166:64:@15665.4]
  assign _T_69250 = _T_69249[13:0]; // @[Modules.scala 166:64:@15666.4]
  assign buffer_4_526 = $signed(_T_69250); // @[Modules.scala 166:64:@15667.4]
  assign _T_69252 = $signed(buffer_4_454) + $signed(buffer_4_455); // @[Modules.scala 166:64:@15669.4]
  assign _T_69253 = _T_69252[13:0]; // @[Modules.scala 166:64:@15670.4]
  assign buffer_4_527 = $signed(_T_69253); // @[Modules.scala 166:64:@15671.4]
  assign _T_69255 = $signed(buffer_4_456) + $signed(buffer_4_457); // @[Modules.scala 166:64:@15673.4]
  assign _T_69256 = _T_69255[13:0]; // @[Modules.scala 166:64:@15674.4]
  assign buffer_4_528 = $signed(_T_69256); // @[Modules.scala 166:64:@15675.4]
  assign _T_69258 = $signed(buffer_4_458) + $signed(buffer_4_459); // @[Modules.scala 166:64:@15677.4]
  assign _T_69259 = _T_69258[13:0]; // @[Modules.scala 166:64:@15678.4]
  assign buffer_4_529 = $signed(_T_69259); // @[Modules.scala 166:64:@15679.4]
  assign _T_69261 = $signed(buffer_4_460) + $signed(buffer_4_461); // @[Modules.scala 166:64:@15681.4]
  assign _T_69262 = _T_69261[13:0]; // @[Modules.scala 166:64:@15682.4]
  assign buffer_4_530 = $signed(_T_69262); // @[Modules.scala 166:64:@15683.4]
  assign _T_69264 = $signed(buffer_4_462) + $signed(buffer_4_463); // @[Modules.scala 166:64:@15685.4]
  assign _T_69265 = _T_69264[13:0]; // @[Modules.scala 166:64:@15686.4]
  assign buffer_4_531 = $signed(_T_69265); // @[Modules.scala 166:64:@15687.4]
  assign _T_69267 = $signed(buffer_4_464) + $signed(buffer_4_465); // @[Modules.scala 166:64:@15689.4]
  assign _T_69268 = _T_69267[13:0]; // @[Modules.scala 166:64:@15690.4]
  assign buffer_4_532 = $signed(_T_69268); // @[Modules.scala 166:64:@15691.4]
  assign _T_69270 = $signed(buffer_4_466) + $signed(buffer_4_467); // @[Modules.scala 166:64:@15693.4]
  assign _T_69271 = _T_69270[13:0]; // @[Modules.scala 166:64:@15694.4]
  assign buffer_4_533 = $signed(_T_69271); // @[Modules.scala 166:64:@15695.4]
  assign _T_69273 = $signed(buffer_4_468) + $signed(buffer_4_469); // @[Modules.scala 166:64:@15697.4]
  assign _T_69274 = _T_69273[13:0]; // @[Modules.scala 166:64:@15698.4]
  assign buffer_4_534 = $signed(_T_69274); // @[Modules.scala 166:64:@15699.4]
  assign _T_69276 = $signed(buffer_4_470) + $signed(buffer_4_471); // @[Modules.scala 166:64:@15701.4]
  assign _T_69277 = _T_69276[13:0]; // @[Modules.scala 166:64:@15702.4]
  assign buffer_4_535 = $signed(_T_69277); // @[Modules.scala 166:64:@15703.4]
  assign _T_69279 = $signed(buffer_4_472) + $signed(buffer_4_473); // @[Modules.scala 166:64:@15705.4]
  assign _T_69280 = _T_69279[13:0]; // @[Modules.scala 166:64:@15706.4]
  assign buffer_4_536 = $signed(_T_69280); // @[Modules.scala 166:64:@15707.4]
  assign _T_69282 = $signed(buffer_4_474) + $signed(buffer_4_475); // @[Modules.scala 166:64:@15709.4]
  assign _T_69283 = _T_69282[13:0]; // @[Modules.scala 166:64:@15710.4]
  assign buffer_4_537 = $signed(_T_69283); // @[Modules.scala 166:64:@15711.4]
  assign _T_69285 = $signed(buffer_4_476) + $signed(buffer_4_477); // @[Modules.scala 166:64:@15713.4]
  assign _T_69286 = _T_69285[13:0]; // @[Modules.scala 166:64:@15714.4]
  assign buffer_4_538 = $signed(_T_69286); // @[Modules.scala 166:64:@15715.4]
  assign _T_69288 = $signed(buffer_4_478) + $signed(buffer_4_479); // @[Modules.scala 166:64:@15717.4]
  assign _T_69289 = _T_69288[13:0]; // @[Modules.scala 166:64:@15718.4]
  assign buffer_4_539 = $signed(_T_69289); // @[Modules.scala 166:64:@15719.4]
  assign _T_69291 = $signed(buffer_4_480) + $signed(buffer_4_481); // @[Modules.scala 166:64:@15721.4]
  assign _T_69292 = _T_69291[13:0]; // @[Modules.scala 166:64:@15722.4]
  assign buffer_4_540 = $signed(_T_69292); // @[Modules.scala 166:64:@15723.4]
  assign _T_69294 = $signed(buffer_4_482) + $signed(buffer_4_483); // @[Modules.scala 166:64:@15725.4]
  assign _T_69295 = _T_69294[13:0]; // @[Modules.scala 166:64:@15726.4]
  assign buffer_4_541 = $signed(_T_69295); // @[Modules.scala 166:64:@15727.4]
  assign _T_69297 = $signed(buffer_4_484) + $signed(buffer_4_485); // @[Modules.scala 166:64:@15729.4]
  assign _T_69298 = _T_69297[13:0]; // @[Modules.scala 166:64:@15730.4]
  assign buffer_4_542 = $signed(_T_69298); // @[Modules.scala 166:64:@15731.4]
  assign _T_69300 = $signed(buffer_4_486) + $signed(buffer_4_487); // @[Modules.scala 166:64:@15733.4]
  assign _T_69301 = _T_69300[13:0]; // @[Modules.scala 166:64:@15734.4]
  assign buffer_4_543 = $signed(_T_69301); // @[Modules.scala 166:64:@15735.4]
  assign _T_69303 = $signed(buffer_4_488) + $signed(buffer_4_489); // @[Modules.scala 166:64:@15737.4]
  assign _T_69304 = _T_69303[13:0]; // @[Modules.scala 166:64:@15738.4]
  assign buffer_4_544 = $signed(_T_69304); // @[Modules.scala 166:64:@15739.4]
  assign _T_69306 = $signed(buffer_4_490) + $signed(buffer_4_491); // @[Modules.scala 166:64:@15741.4]
  assign _T_69307 = _T_69306[13:0]; // @[Modules.scala 166:64:@15742.4]
  assign buffer_4_545 = $signed(_T_69307); // @[Modules.scala 166:64:@15743.4]
  assign _T_69309 = $signed(buffer_4_492) + $signed(buffer_4_493); // @[Modules.scala 166:64:@15745.4]
  assign _T_69310 = _T_69309[13:0]; // @[Modules.scala 166:64:@15746.4]
  assign buffer_4_546 = $signed(_T_69310); // @[Modules.scala 166:64:@15747.4]
  assign _T_69312 = $signed(buffer_4_494) + $signed(buffer_4_495); // @[Modules.scala 166:64:@15749.4]
  assign _T_69313 = _T_69312[13:0]; // @[Modules.scala 166:64:@15750.4]
  assign buffer_4_547 = $signed(_T_69313); // @[Modules.scala 166:64:@15751.4]
  assign _T_69315 = $signed(buffer_4_496) + $signed(buffer_4_497); // @[Modules.scala 166:64:@15753.4]
  assign _T_69316 = _T_69315[13:0]; // @[Modules.scala 166:64:@15754.4]
  assign buffer_4_548 = $signed(_T_69316); // @[Modules.scala 166:64:@15755.4]
  assign _T_69318 = $signed(buffer_4_498) + $signed(buffer_4_499); // @[Modules.scala 166:64:@15757.4]
  assign _T_69319 = _T_69318[13:0]; // @[Modules.scala 166:64:@15758.4]
  assign buffer_4_549 = $signed(_T_69319); // @[Modules.scala 166:64:@15759.4]
  assign _T_69321 = $signed(buffer_4_500) + $signed(buffer_4_501); // @[Modules.scala 166:64:@15761.4]
  assign _T_69322 = _T_69321[13:0]; // @[Modules.scala 166:64:@15762.4]
  assign buffer_4_550 = $signed(_T_69322); // @[Modules.scala 166:64:@15763.4]
  assign _T_69324 = $signed(buffer_4_502) + $signed(buffer_2_521); // @[Modules.scala 166:64:@15765.4]
  assign _T_69325 = _T_69324[13:0]; // @[Modules.scala 166:64:@15766.4]
  assign buffer_4_551 = $signed(_T_69325); // @[Modules.scala 166:64:@15767.4]
  assign _T_69327 = $signed(buffer_4_504) + $signed(buffer_4_505); // @[Modules.scala 166:64:@15769.4]
  assign _T_69328 = _T_69327[13:0]; // @[Modules.scala 166:64:@15770.4]
  assign buffer_4_552 = $signed(_T_69328); // @[Modules.scala 166:64:@15771.4]
  assign _T_69330 = $signed(buffer_4_506) + $signed(buffer_4_507); // @[Modules.scala 166:64:@15773.4]
  assign _T_69331 = _T_69330[13:0]; // @[Modules.scala 166:64:@15774.4]
  assign buffer_4_553 = $signed(_T_69331); // @[Modules.scala 166:64:@15775.4]
  assign _T_69333 = $signed(buffer_4_508) + $signed(buffer_4_509); // @[Modules.scala 166:64:@15777.4]
  assign _T_69334 = _T_69333[13:0]; // @[Modules.scala 166:64:@15778.4]
  assign buffer_4_554 = $signed(_T_69334); // @[Modules.scala 166:64:@15779.4]
  assign _T_69336 = $signed(buffer_4_510) + $signed(buffer_4_511); // @[Modules.scala 166:64:@15781.4]
  assign _T_69337 = _T_69336[13:0]; // @[Modules.scala 166:64:@15782.4]
  assign buffer_4_555 = $signed(_T_69337); // @[Modules.scala 166:64:@15783.4]
  assign _T_69339 = $signed(buffer_4_512) + $signed(buffer_4_513); // @[Modules.scala 166:64:@15785.4]
  assign _T_69340 = _T_69339[13:0]; // @[Modules.scala 166:64:@15786.4]
  assign buffer_4_556 = $signed(_T_69340); // @[Modules.scala 166:64:@15787.4]
  assign _T_69342 = $signed(buffer_4_514) + $signed(buffer_4_515); // @[Modules.scala 166:64:@15789.4]
  assign _T_69343 = _T_69342[13:0]; // @[Modules.scala 166:64:@15790.4]
  assign buffer_4_557 = $signed(_T_69343); // @[Modules.scala 166:64:@15791.4]
  assign _T_69345 = $signed(buffer_4_516) + $signed(buffer_4_517); // @[Modules.scala 166:64:@15793.4]
  assign _T_69346 = _T_69345[13:0]; // @[Modules.scala 166:64:@15794.4]
  assign buffer_4_558 = $signed(_T_69346); // @[Modules.scala 166:64:@15795.4]
  assign _T_69348 = $signed(buffer_4_518) + $signed(buffer_4_519); // @[Modules.scala 166:64:@15797.4]
  assign _T_69349 = _T_69348[13:0]; // @[Modules.scala 166:64:@15798.4]
  assign buffer_4_559 = $signed(_T_69349); // @[Modules.scala 166:64:@15799.4]
  assign _T_69351 = $signed(buffer_4_520) + $signed(buffer_4_521); // @[Modules.scala 166:64:@15801.4]
  assign _T_69352 = _T_69351[13:0]; // @[Modules.scala 166:64:@15802.4]
  assign buffer_4_560 = $signed(_T_69352); // @[Modules.scala 166:64:@15803.4]
  assign _T_69354 = $signed(buffer_4_522) + $signed(buffer_4_523); // @[Modules.scala 166:64:@15805.4]
  assign _T_69355 = _T_69354[13:0]; // @[Modules.scala 166:64:@15806.4]
  assign buffer_4_561 = $signed(_T_69355); // @[Modules.scala 166:64:@15807.4]
  assign _T_69357 = $signed(buffer_4_525) + $signed(buffer_4_526); // @[Modules.scala 166:64:@15809.4]
  assign _T_69358 = _T_69357[13:0]; // @[Modules.scala 166:64:@15810.4]
  assign buffer_4_562 = $signed(_T_69358); // @[Modules.scala 166:64:@15811.4]
  assign _T_69360 = $signed(buffer_4_527) + $signed(buffer_4_528); // @[Modules.scala 166:64:@15813.4]
  assign _T_69361 = _T_69360[13:0]; // @[Modules.scala 166:64:@15814.4]
  assign buffer_4_563 = $signed(_T_69361); // @[Modules.scala 166:64:@15815.4]
  assign _T_69363 = $signed(buffer_4_529) + $signed(buffer_4_530); // @[Modules.scala 166:64:@15817.4]
  assign _T_69364 = _T_69363[13:0]; // @[Modules.scala 166:64:@15818.4]
  assign buffer_4_564 = $signed(_T_69364); // @[Modules.scala 166:64:@15819.4]
  assign _T_69366 = $signed(buffer_4_531) + $signed(buffer_4_532); // @[Modules.scala 166:64:@15821.4]
  assign _T_69367 = _T_69366[13:0]; // @[Modules.scala 166:64:@15822.4]
  assign buffer_4_565 = $signed(_T_69367); // @[Modules.scala 166:64:@15823.4]
  assign _T_69369 = $signed(buffer_4_533) + $signed(buffer_4_534); // @[Modules.scala 166:64:@15825.4]
  assign _T_69370 = _T_69369[13:0]; // @[Modules.scala 166:64:@15826.4]
  assign buffer_4_566 = $signed(_T_69370); // @[Modules.scala 166:64:@15827.4]
  assign _T_69372 = $signed(buffer_4_535) + $signed(buffer_4_536); // @[Modules.scala 166:64:@15829.4]
  assign _T_69373 = _T_69372[13:0]; // @[Modules.scala 166:64:@15830.4]
  assign buffer_4_567 = $signed(_T_69373); // @[Modules.scala 166:64:@15831.4]
  assign _T_69375 = $signed(buffer_4_537) + $signed(buffer_4_538); // @[Modules.scala 166:64:@15833.4]
  assign _T_69376 = _T_69375[13:0]; // @[Modules.scala 166:64:@15834.4]
  assign buffer_4_568 = $signed(_T_69376); // @[Modules.scala 166:64:@15835.4]
  assign _T_69378 = $signed(buffer_4_539) + $signed(buffer_4_540); // @[Modules.scala 166:64:@15837.4]
  assign _T_69379 = _T_69378[13:0]; // @[Modules.scala 166:64:@15838.4]
  assign buffer_4_569 = $signed(_T_69379); // @[Modules.scala 166:64:@15839.4]
  assign _T_69381 = $signed(buffer_4_541) + $signed(buffer_4_542); // @[Modules.scala 166:64:@15841.4]
  assign _T_69382 = _T_69381[13:0]; // @[Modules.scala 166:64:@15842.4]
  assign buffer_4_570 = $signed(_T_69382); // @[Modules.scala 166:64:@15843.4]
  assign _T_69384 = $signed(buffer_4_543) + $signed(buffer_4_544); // @[Modules.scala 166:64:@15845.4]
  assign _T_69385 = _T_69384[13:0]; // @[Modules.scala 166:64:@15846.4]
  assign buffer_4_571 = $signed(_T_69385); // @[Modules.scala 166:64:@15847.4]
  assign _T_69387 = $signed(buffer_4_545) + $signed(buffer_4_546); // @[Modules.scala 166:64:@15849.4]
  assign _T_69388 = _T_69387[13:0]; // @[Modules.scala 166:64:@15850.4]
  assign buffer_4_572 = $signed(_T_69388); // @[Modules.scala 166:64:@15851.4]
  assign _T_69390 = $signed(buffer_4_547) + $signed(buffer_4_548); // @[Modules.scala 166:64:@15853.4]
  assign _T_69391 = _T_69390[13:0]; // @[Modules.scala 166:64:@15854.4]
  assign buffer_4_573 = $signed(_T_69391); // @[Modules.scala 166:64:@15855.4]
  assign _T_69393 = $signed(buffer_4_549) + $signed(buffer_4_550); // @[Modules.scala 166:64:@15857.4]
  assign _T_69394 = _T_69393[13:0]; // @[Modules.scala 166:64:@15858.4]
  assign buffer_4_574 = $signed(_T_69394); // @[Modules.scala 166:64:@15859.4]
  assign _T_69396 = $signed(buffer_4_551) + $signed(buffer_4_552); // @[Modules.scala 166:64:@15861.4]
  assign _T_69397 = _T_69396[13:0]; // @[Modules.scala 166:64:@15862.4]
  assign buffer_4_575 = $signed(_T_69397); // @[Modules.scala 166:64:@15863.4]
  assign _T_69399 = $signed(buffer_4_553) + $signed(buffer_4_554); // @[Modules.scala 166:64:@15865.4]
  assign _T_69400 = _T_69399[13:0]; // @[Modules.scala 166:64:@15866.4]
  assign buffer_4_576 = $signed(_T_69400); // @[Modules.scala 166:64:@15867.4]
  assign _T_69402 = $signed(buffer_4_555) + $signed(buffer_4_556); // @[Modules.scala 166:64:@15869.4]
  assign _T_69403 = _T_69402[13:0]; // @[Modules.scala 166:64:@15870.4]
  assign buffer_4_577 = $signed(_T_69403); // @[Modules.scala 166:64:@15871.4]
  assign _T_69405 = $signed(buffer_4_557) + $signed(buffer_4_558); // @[Modules.scala 166:64:@15873.4]
  assign _T_69406 = _T_69405[13:0]; // @[Modules.scala 166:64:@15874.4]
  assign buffer_4_578 = $signed(_T_69406); // @[Modules.scala 166:64:@15875.4]
  assign _T_69408 = $signed(buffer_4_559) + $signed(buffer_4_560); // @[Modules.scala 166:64:@15877.4]
  assign _T_69409 = _T_69408[13:0]; // @[Modules.scala 166:64:@15878.4]
  assign buffer_4_579 = $signed(_T_69409); // @[Modules.scala 166:64:@15879.4]
  assign _T_69411 = $signed(buffer_4_561) + $signed(buffer_4_524); // @[Modules.scala 172:66:@15881.4]
  assign _T_69412 = _T_69411[13:0]; // @[Modules.scala 172:66:@15882.4]
  assign buffer_4_580 = $signed(_T_69412); // @[Modules.scala 172:66:@15883.4]
  assign _T_69414 = $signed(buffer_4_562) + $signed(buffer_4_563); // @[Modules.scala 166:64:@15885.4]
  assign _T_69415 = _T_69414[13:0]; // @[Modules.scala 166:64:@15886.4]
  assign buffer_4_581 = $signed(_T_69415); // @[Modules.scala 166:64:@15887.4]
  assign _T_69417 = $signed(buffer_4_564) + $signed(buffer_4_565); // @[Modules.scala 166:64:@15889.4]
  assign _T_69418 = _T_69417[13:0]; // @[Modules.scala 166:64:@15890.4]
  assign buffer_4_582 = $signed(_T_69418); // @[Modules.scala 166:64:@15891.4]
  assign _T_69420 = $signed(buffer_4_566) + $signed(buffer_4_567); // @[Modules.scala 166:64:@15893.4]
  assign _T_69421 = _T_69420[13:0]; // @[Modules.scala 166:64:@15894.4]
  assign buffer_4_583 = $signed(_T_69421); // @[Modules.scala 166:64:@15895.4]
  assign _T_69423 = $signed(buffer_4_568) + $signed(buffer_4_569); // @[Modules.scala 166:64:@15897.4]
  assign _T_69424 = _T_69423[13:0]; // @[Modules.scala 166:64:@15898.4]
  assign buffer_4_584 = $signed(_T_69424); // @[Modules.scala 166:64:@15899.4]
  assign _T_69426 = $signed(buffer_4_570) + $signed(buffer_4_571); // @[Modules.scala 166:64:@15901.4]
  assign _T_69427 = _T_69426[13:0]; // @[Modules.scala 166:64:@15902.4]
  assign buffer_4_585 = $signed(_T_69427); // @[Modules.scala 166:64:@15903.4]
  assign _T_69429 = $signed(buffer_4_572) + $signed(buffer_4_573); // @[Modules.scala 166:64:@15905.4]
  assign _T_69430 = _T_69429[13:0]; // @[Modules.scala 166:64:@15906.4]
  assign buffer_4_586 = $signed(_T_69430); // @[Modules.scala 166:64:@15907.4]
  assign _T_69432 = $signed(buffer_4_574) + $signed(buffer_4_575); // @[Modules.scala 166:64:@15909.4]
  assign _T_69433 = _T_69432[13:0]; // @[Modules.scala 166:64:@15910.4]
  assign buffer_4_587 = $signed(_T_69433); // @[Modules.scala 166:64:@15911.4]
  assign _T_69435 = $signed(buffer_4_576) + $signed(buffer_4_577); // @[Modules.scala 166:64:@15913.4]
  assign _T_69436 = _T_69435[13:0]; // @[Modules.scala 166:64:@15914.4]
  assign buffer_4_588 = $signed(_T_69436); // @[Modules.scala 166:64:@15915.4]
  assign _T_69438 = $signed(buffer_4_578) + $signed(buffer_4_579); // @[Modules.scala 166:64:@15917.4]
  assign _T_69439 = _T_69438[13:0]; // @[Modules.scala 166:64:@15918.4]
  assign buffer_4_589 = $signed(_T_69439); // @[Modules.scala 166:64:@15919.4]
  assign _T_69441 = $signed(buffer_4_581) + $signed(buffer_4_582); // @[Modules.scala 166:64:@15921.4]
  assign _T_69442 = _T_69441[13:0]; // @[Modules.scala 166:64:@15922.4]
  assign buffer_4_590 = $signed(_T_69442); // @[Modules.scala 166:64:@15923.4]
  assign _T_69444 = $signed(buffer_4_583) + $signed(buffer_4_584); // @[Modules.scala 166:64:@15925.4]
  assign _T_69445 = _T_69444[13:0]; // @[Modules.scala 166:64:@15926.4]
  assign buffer_4_591 = $signed(_T_69445); // @[Modules.scala 166:64:@15927.4]
  assign _T_69447 = $signed(buffer_4_585) + $signed(buffer_4_586); // @[Modules.scala 166:64:@15929.4]
  assign _T_69448 = _T_69447[13:0]; // @[Modules.scala 166:64:@15930.4]
  assign buffer_4_592 = $signed(_T_69448); // @[Modules.scala 166:64:@15931.4]
  assign _T_69450 = $signed(buffer_4_587) + $signed(buffer_4_588); // @[Modules.scala 166:64:@15933.4]
  assign _T_69451 = _T_69450[13:0]; // @[Modules.scala 166:64:@15934.4]
  assign buffer_4_593 = $signed(_T_69451); // @[Modules.scala 166:64:@15935.4]
  assign _T_69453 = $signed(buffer_4_589) + $signed(buffer_4_580); // @[Modules.scala 172:66:@15937.4]
  assign _T_69454 = _T_69453[13:0]; // @[Modules.scala 172:66:@15938.4]
  assign buffer_4_594 = $signed(_T_69454); // @[Modules.scala 172:66:@15939.4]
  assign _T_69456 = $signed(buffer_4_590) + $signed(buffer_4_591); // @[Modules.scala 166:64:@15941.4]
  assign _T_69457 = _T_69456[13:0]; // @[Modules.scala 166:64:@15942.4]
  assign buffer_4_595 = $signed(_T_69457); // @[Modules.scala 166:64:@15943.4]
  assign _T_69459 = $signed(buffer_4_592) + $signed(buffer_4_593); // @[Modules.scala 166:64:@15945.4]
  assign _T_69460 = _T_69459[13:0]; // @[Modules.scala 166:64:@15946.4]
  assign buffer_4_596 = $signed(_T_69460); // @[Modules.scala 166:64:@15947.4]
  assign _T_69462 = $signed(buffer_4_595) + $signed(buffer_4_596); // @[Modules.scala 160:64:@15949.4]
  assign _T_69463 = _T_69462[13:0]; // @[Modules.scala 160:64:@15950.4]
  assign buffer_4_597 = $signed(_T_69463); // @[Modules.scala 160:64:@15951.4]
  assign _T_69465 = $signed(buffer_4_597) + $signed(buffer_4_594); // @[Modules.scala 172:66:@15953.4]
  assign _T_69466 = _T_69465[13:0]; // @[Modules.scala 172:66:@15954.4]
  assign buffer_4_598 = $signed(_T_69466); // @[Modules.scala 172:66:@15955.4]
  assign _T_69469 = $signed(4'sh1) * $signed(io_in_0); // @[Modules.scala 143:74:@16142.4]
  assign _T_69471 = $signed(-4'sh1) * $signed(io_in_5); // @[Modules.scala 144:80:@16143.4]
  assign _GEN_357 = {{1{_T_69471[4]}},_T_69471}; // @[Modules.scala 143:103:@16144.4]
  assign _T_69472 = $signed(_T_69469) + $signed(_GEN_357); // @[Modules.scala 143:103:@16144.4]
  assign _T_69473 = _T_69472[5:0]; // @[Modules.scala 143:103:@16145.4]
  assign _T_69474 = $signed(_T_69473); // @[Modules.scala 143:103:@16146.4]
  assign _T_69500 = $signed(_T_57232) + $signed(_GEN_279); // @[Modules.scala 143:103:@16168.4]
  assign _T_69501 = _T_69500[5:0]; // @[Modules.scala 143:103:@16169.4]
  assign _T_69502 = $signed(_T_69501); // @[Modules.scala 143:103:@16170.4]
  assign _T_69514 = $signed(_T_66500) + $signed(_T_63375); // @[Modules.scala 143:103:@16180.4]
  assign _T_69515 = _T_69514[4:0]; // @[Modules.scala 143:103:@16181.4]
  assign _T_69516 = $signed(_T_69515); // @[Modules.scala 143:103:@16182.4]
  assign _GEN_359 = {{1{_T_63403[4]}},_T_63403}; // @[Modules.scala 143:103:@16198.4]
  assign _T_69535 = $signed(_T_54257) + $signed(_GEN_359); // @[Modules.scala 143:103:@16198.4]
  assign _T_69536 = _T_69535[5:0]; // @[Modules.scala 143:103:@16199.4]
  assign _T_69537 = $signed(_T_69536); // @[Modules.scala 143:103:@16200.4]
  assign _T_69548 = $signed(-4'sh1) * $signed(io_in_52); // @[Modules.scala 144:80:@16209.4]
  assign _GEN_360 = {{1{_T_69548[4]}},_T_69548}; // @[Modules.scala 143:103:@16210.4]
  assign _T_69549 = $signed(_T_54276) + $signed(_GEN_360); // @[Modules.scala 143:103:@16210.4]
  assign _T_69550 = _T_69549[5:0]; // @[Modules.scala 143:103:@16211.4]
  assign _T_69551 = $signed(_T_69550); // @[Modules.scala 143:103:@16212.4]
  assign _T_69556 = $signed(_T_54278) + $signed(_GEN_80); // @[Modules.scala 143:103:@16216.4]
  assign _T_69557 = _T_69556[5:0]; // @[Modules.scala 143:103:@16217.4]
  assign _T_69558 = $signed(_T_69557); // @[Modules.scala 143:103:@16218.4]
  assign _T_69619 = $signed(_GEN_282) + $signed(_T_54348); // @[Modules.scala 143:103:@16270.4]
  assign _T_69620 = _T_69619[5:0]; // @[Modules.scala 143:103:@16271.4]
  assign _T_69621 = $signed(_T_69620); // @[Modules.scala 143:103:@16272.4]
  assign _GEN_364 = {{1{_T_57386[4]}},_T_57386}; // @[Modules.scala 143:103:@16288.4]
  assign _T_69640 = $signed(_T_54369) + $signed(_GEN_364); // @[Modules.scala 143:103:@16288.4]
  assign _T_69641 = _T_69640[5:0]; // @[Modules.scala 143:103:@16289.4]
  assign _T_69642 = $signed(_T_69641); // @[Modules.scala 143:103:@16290.4]
  assign _T_69661 = $signed(_T_60430) + $signed(_T_63541); // @[Modules.scala 143:103:@16306.4]
  assign _T_69662 = _T_69661[4:0]; // @[Modules.scala 143:103:@16307.4]
  assign _T_69663 = $signed(_T_69662); // @[Modules.scala 143:103:@16308.4]
  assign _T_69668 = $signed(_T_63543) + $signed(_T_57409); // @[Modules.scala 143:103:@16312.4]
  assign _T_69669 = _T_69668[4:0]; // @[Modules.scala 143:103:@16313.4]
  assign _T_69670 = $signed(_T_69669); // @[Modules.scala 143:103:@16314.4]
  assign _T_69696 = $signed(_T_63571) + $signed(_T_54439); // @[Modules.scala 143:103:@16336.4]
  assign _T_69697 = _T_69696[4:0]; // @[Modules.scala 143:103:@16337.4]
  assign _T_69698 = $signed(_T_69697); // @[Modules.scala 143:103:@16338.4]
  assign _T_69703 = $signed(_T_60474) + $signed(_T_54446); // @[Modules.scala 143:103:@16342.4]
  assign _T_69704 = _T_69703[4:0]; // @[Modules.scala 143:103:@16343.4]
  assign _T_69705 = $signed(_T_69704); // @[Modules.scala 143:103:@16344.4]
  assign _GEN_365 = {{1{_T_63590[4]}},_T_63590}; // @[Modules.scala 143:103:@16348.4]
  assign _T_69710 = $signed(_T_57451) + $signed(_GEN_365); // @[Modules.scala 143:103:@16348.4]
  assign _T_69711 = _T_69710[5:0]; // @[Modules.scala 143:103:@16349.4]
  assign _T_69712 = $signed(_T_69711); // @[Modules.scala 143:103:@16350.4]
  assign _T_69724 = $signed(_T_60488) + $signed(_T_54460); // @[Modules.scala 143:103:@16360.4]
  assign _T_69725 = _T_69724[5:0]; // @[Modules.scala 143:103:@16361.4]
  assign _T_69726 = $signed(_T_69725); // @[Modules.scala 143:103:@16362.4]
  assign _T_69749 = $signed(4'sh1) * $signed(io_in_127); // @[Modules.scala 143:74:@16382.4]
  assign _T_69752 = $signed(_T_69749) + $signed(_T_54486); // @[Modules.scala 143:103:@16384.4]
  assign _T_69753 = _T_69752[5:0]; // @[Modules.scala 143:103:@16385.4]
  assign _T_69754 = $signed(_T_69753); // @[Modules.scala 143:103:@16386.4]
  assign _T_69763 = $signed(-4'sh1) * $signed(io_in_132); // @[Modules.scala 143:74:@16394.4]
  assign _T_69765 = $signed(-4'sh1) * $signed(io_in_133); // @[Modules.scala 144:80:@16395.4]
  assign _T_69766 = $signed(_T_69763) + $signed(_T_69765); // @[Modules.scala 143:103:@16396.4]
  assign _T_69767 = _T_69766[4:0]; // @[Modules.scala 143:103:@16397.4]
  assign _T_69768 = $signed(_T_69767); // @[Modules.scala 143:103:@16398.4]
  assign _T_69770 = $signed(-4'sh1) * $signed(io_in_134); // @[Modules.scala 143:74:@16400.4]
  assign _T_69773 = $signed(_T_69770) + $signed(_T_54507); // @[Modules.scala 143:103:@16402.4]
  assign _T_69774 = _T_69773[4:0]; // @[Modules.scala 143:103:@16403.4]
  assign _T_69775 = $signed(_T_69774); // @[Modules.scala 143:103:@16404.4]
  assign _GEN_366 = {{1{_T_54509[4]}},_T_54509}; // @[Modules.scala 143:103:@16408.4]
  assign _T_69780 = $signed(_GEN_366) + $signed(_T_57514); // @[Modules.scala 143:103:@16408.4]
  assign _T_69781 = _T_69780[5:0]; // @[Modules.scala 143:103:@16409.4]
  assign _T_69782 = $signed(_T_69781); // @[Modules.scala 143:103:@16410.4]
  assign _T_69794 = $signed(_GEN_290) + $signed(_T_57540); // @[Modules.scala 143:103:@16420.4]
  assign _T_69795 = _T_69794[5:0]; // @[Modules.scala 143:103:@16421.4]
  assign _T_69796 = $signed(_T_69795); // @[Modules.scala 143:103:@16422.4]
  assign _T_69819 = $signed(4'sh1) * $signed(io_in_153); // @[Modules.scala 143:74:@16442.4]
  assign _T_69822 = $signed(_T_69819) + $signed(_T_63704); // @[Modules.scala 143:103:@16444.4]
  assign _T_69823 = _T_69822[5:0]; // @[Modules.scala 143:103:@16445.4]
  assign _T_69824 = $signed(_T_69823); // @[Modules.scala 143:103:@16446.4]
  assign _T_69826 = $signed(4'sh1) * $signed(io_in_155); // @[Modules.scala 143:74:@16448.4]
  assign _T_69828 = $signed(4'sh1) * $signed(io_in_156); // @[Modules.scala 144:80:@16449.4]
  assign _T_69829 = $signed(_T_69826) + $signed(_T_69828); // @[Modules.scala 143:103:@16450.4]
  assign _T_69830 = _T_69829[5:0]; // @[Modules.scala 143:103:@16451.4]
  assign _T_69831 = $signed(_T_69830); // @[Modules.scala 143:103:@16452.4]
  assign _T_69833 = $signed(4'sh1) * $signed(io_in_157); // @[Modules.scala 143:74:@16454.4]
  assign _GEN_369 = {{1{_T_66841[4]}},_T_66841}; // @[Modules.scala 143:103:@16456.4]
  assign _T_69836 = $signed(_T_69833) + $signed(_GEN_369); // @[Modules.scala 143:103:@16456.4]
  assign _T_69837 = _T_69836[5:0]; // @[Modules.scala 143:103:@16457.4]
  assign _T_69838 = $signed(_T_69837); // @[Modules.scala 143:103:@16458.4]
  assign _T_69843 = $signed(_T_54551) + $signed(_T_60607); // @[Modules.scala 143:103:@16462.4]
  assign _T_69844 = _T_69843[4:0]; // @[Modules.scala 143:103:@16463.4]
  assign _T_69845 = $signed(_T_69844); // @[Modules.scala 143:103:@16464.4]
  assign _GEN_370 = {{1{_T_54565[4]}},_T_54565}; // @[Modules.scala 143:103:@16474.4]
  assign _T_69857 = $signed(_GEN_370) + $signed(_T_63739); // @[Modules.scala 143:103:@16474.4]
  assign _T_69858 = _T_69857[5:0]; // @[Modules.scala 143:103:@16475.4]
  assign _T_69859 = $signed(_T_69858); // @[Modules.scala 143:103:@16476.4]
  assign _T_69878 = $signed(_T_63760) + $signed(_T_60642); // @[Modules.scala 143:103:@16492.4]
  assign _T_69879 = _T_69878[4:0]; // @[Modules.scala 143:103:@16493.4]
  assign _T_69880 = $signed(_T_69879); // @[Modules.scala 143:103:@16494.4]
  assign _GEN_373 = {{1{_T_63772[4]}},_T_63772}; // @[Modules.scala 143:103:@16498.4]
  assign _T_69885 = $signed(_T_54598) + $signed(_GEN_373); // @[Modules.scala 143:103:@16498.4]
  assign _T_69886 = _T_69885[5:0]; // @[Modules.scala 143:103:@16499.4]
  assign _T_69887 = $signed(_T_69886); // @[Modules.scala 143:103:@16500.4]
  assign _T_69891 = $signed(4'sh1) * $signed(io_in_177); // @[Modules.scala 144:80:@16503.4]
  assign _T_69892 = $signed(_T_54605) + $signed(_T_69891); // @[Modules.scala 143:103:@16504.4]
  assign _T_69893 = _T_69892[5:0]; // @[Modules.scala 143:103:@16505.4]
  assign _T_69894 = $signed(_T_69893); // @[Modules.scala 143:103:@16506.4]
  assign _T_69899 = $signed(_T_57626) + $signed(_T_57631); // @[Modules.scala 143:103:@16510.4]
  assign _T_69900 = _T_69899[5:0]; // @[Modules.scala 143:103:@16511.4]
  assign _T_69901 = $signed(_T_69900); // @[Modules.scala 143:103:@16512.4]
  assign _T_69913 = $signed(_T_57640) + $signed(_T_57645); // @[Modules.scala 143:103:@16522.4]
  assign _T_69914 = _T_69913[5:0]; // @[Modules.scala 143:103:@16523.4]
  assign _T_69915 = $signed(_T_69914); // @[Modules.scala 143:103:@16524.4]
  assign _T_69920 = $signed(_T_66920) + $signed(_T_66925); // @[Modules.scala 143:103:@16528.4]
  assign _T_69921 = _T_69920[5:0]; // @[Modules.scala 143:103:@16529.4]
  assign _T_69922 = $signed(_T_69921); // @[Modules.scala 143:103:@16530.4]
  assign _T_69924 = $signed(4'sh1) * $signed(io_in_188); // @[Modules.scala 143:74:@16532.4]
  assign _T_69927 = $signed(_T_69924) + $signed(_GEN_162); // @[Modules.scala 143:103:@16534.4]
  assign _T_69928 = _T_69927[5:0]; // @[Modules.scala 143:103:@16535.4]
  assign _T_69929 = $signed(_T_69928); // @[Modules.scala 143:103:@16536.4]
  assign _GEN_375 = {{1{_T_54640[4]}},_T_54640}; // @[Modules.scala 143:103:@16540.4]
  assign _T_69934 = $signed(_GEN_375) + $signed(_T_63823); // @[Modules.scala 143:103:@16540.4]
  assign _T_69935 = _T_69934[5:0]; // @[Modules.scala 143:103:@16541.4]
  assign _T_69936 = $signed(_T_69935); // @[Modules.scala 143:103:@16542.4]
  assign _T_69938 = $signed(4'sh1) * $signed(io_in_194); // @[Modules.scala 143:74:@16544.4]
  assign _T_69941 = $signed(_T_69938) + $signed(_GEN_228); // @[Modules.scala 143:103:@16546.4]
  assign _T_69942 = _T_69941[5:0]; // @[Modules.scala 143:103:@16547.4]
  assign _T_69943 = $signed(_T_69942); // @[Modules.scala 143:103:@16548.4]
  assign _T_69947 = $signed(-4'sh1) * $signed(io_in_197); // @[Modules.scala 144:80:@16551.4]
  assign _T_69948 = $signed(_T_54656) + $signed(_T_69947); // @[Modules.scala 143:103:@16552.4]
  assign _T_69949 = _T_69948[4:0]; // @[Modules.scala 143:103:@16553.4]
  assign _T_69950 = $signed(_T_69949); // @[Modules.scala 143:103:@16554.4]
  assign _T_69955 = $signed(_T_54663) + $signed(_T_54668); // @[Modules.scala 143:103:@16558.4]
  assign _T_69956 = _T_69955[5:0]; // @[Modules.scala 143:103:@16559.4]
  assign _T_69957 = $signed(_T_69956); // @[Modules.scala 143:103:@16560.4]
  assign _GEN_377 = {{1{_T_60719[4]}},_T_60719}; // @[Modules.scala 143:103:@16564.4]
  assign _T_69962 = $signed(_GEN_377) + $signed(_T_54677); // @[Modules.scala 143:103:@16564.4]
  assign _T_69963 = _T_69962[5:0]; // @[Modules.scala 143:103:@16565.4]
  assign _T_69964 = $signed(_T_69963); // @[Modules.scala 143:103:@16566.4]
  assign _T_69968 = $signed(4'sh1) * $signed(io_in_204); // @[Modules.scala 144:80:@16569.4]
  assign _T_69969 = $signed(_T_54682) + $signed(_T_69968); // @[Modules.scala 143:103:@16570.4]
  assign _T_69970 = _T_69969[5:0]; // @[Modules.scala 143:103:@16571.4]
  assign _T_69971 = $signed(_T_69970); // @[Modules.scala 143:103:@16572.4]
  assign _T_69973 = $signed(4'sh1) * $signed(io_in_205); // @[Modules.scala 143:74:@16574.4]
  assign _T_69976 = $signed(_T_69973) + $signed(_T_54689); // @[Modules.scala 143:103:@16576.4]
  assign _T_69977 = _T_69976[5:0]; // @[Modules.scala 143:103:@16577.4]
  assign _T_69978 = $signed(_T_69977); // @[Modules.scala 143:103:@16578.4]
  assign _T_70004 = $signed(_T_57729) + $signed(_T_63884); // @[Modules.scala 143:103:@16600.4]
  assign _T_70005 = _T_70004[5:0]; // @[Modules.scala 143:103:@16601.4]
  assign _T_70006 = $signed(_T_70005); // @[Modules.scala 143:103:@16602.4]
  assign _T_70010 = $signed(4'sh1) * $signed(io_in_217); // @[Modules.scala 144:80:@16605.4]
  assign _T_70011 = $signed(_T_57738) + $signed(_T_70010); // @[Modules.scala 143:103:@16606.4]
  assign _T_70012 = _T_70011[5:0]; // @[Modules.scala 143:103:@16607.4]
  assign _T_70013 = $signed(_T_70012); // @[Modules.scala 143:103:@16608.4]
  assign _GEN_378 = {{1{_T_57759[4]}},_T_57759}; // @[Modules.scala 143:103:@16624.4]
  assign _T_70032 = $signed(_GEN_378) + $signed(_T_57764); // @[Modules.scala 143:103:@16624.4]
  assign _T_70033 = _T_70032[5:0]; // @[Modules.scala 143:103:@16625.4]
  assign _T_70034 = $signed(_T_70033); // @[Modules.scala 143:103:@16626.4]
  assign _T_70036 = $signed(-4'sh1) * $signed(io_in_225); // @[Modules.scala 143:74:@16628.4]
  assign _GEN_379 = {{1{_T_70036[4]}},_T_70036}; // @[Modules.scala 143:103:@16630.4]
  assign _T_70039 = $signed(_GEN_379) + $signed(_T_54733); // @[Modules.scala 143:103:@16630.4]
  assign _T_70040 = _T_70039[5:0]; // @[Modules.scala 143:103:@16631.4]
  assign _T_70041 = $signed(_T_70040); // @[Modules.scala 143:103:@16632.4]
  assign _T_70057 = $signed(4'sh1) * $signed(io_in_233); // @[Modules.scala 143:74:@16646.4]
  assign _T_70059 = $signed(4'sh1) * $signed(io_in_234); // @[Modules.scala 144:80:@16647.4]
  assign _T_70060 = $signed(_T_70057) + $signed(_T_70059); // @[Modules.scala 143:103:@16648.4]
  assign _T_70061 = _T_70060[5:0]; // @[Modules.scala 143:103:@16649.4]
  assign _T_70062 = $signed(_T_70061); // @[Modules.scala 143:103:@16650.4]
  assign _T_70067 = $signed(_T_54761) + $signed(_T_67053); // @[Modules.scala 143:103:@16654.4]
  assign _T_70068 = _T_70067[5:0]; // @[Modules.scala 143:103:@16655.4]
  assign _T_70069 = $signed(_T_70068); // @[Modules.scala 143:103:@16656.4]
  assign _T_70099 = $signed(4'sh1) * $signed(io_in_245); // @[Modules.scala 143:74:@16682.4]
  assign _T_70102 = $signed(_T_70099) + $signed(_T_63975); // @[Modules.scala 143:103:@16684.4]
  assign _T_70103 = _T_70102[5:0]; // @[Modules.scala 143:103:@16685.4]
  assign _T_70104 = $signed(_T_70103); // @[Modules.scala 143:103:@16686.4]
  assign _T_70109 = $signed(_T_63977) + $signed(_T_63982); // @[Modules.scala 143:103:@16690.4]
  assign _T_70110 = _T_70109[5:0]; // @[Modules.scala 143:103:@16691.4]
  assign _T_70111 = $signed(_T_70110); // @[Modules.scala 143:103:@16692.4]
  assign _T_70116 = $signed(_T_63984) + $signed(_T_63989); // @[Modules.scala 143:103:@16696.4]
  assign _T_70117 = _T_70116[5:0]; // @[Modules.scala 143:103:@16697.4]
  assign _T_70118 = $signed(_T_70117); // @[Modules.scala 143:103:@16698.4]
  assign _T_70123 = $signed(_T_54808) + $signed(_T_57850); // @[Modules.scala 143:103:@16702.4]
  assign _T_70124 = _T_70123[5:0]; // @[Modules.scala 143:103:@16703.4]
  assign _T_70125 = $signed(_T_70124); // @[Modules.scala 143:103:@16704.4]
  assign _T_70137 = $signed(_T_57857) + $signed(_T_54822); // @[Modules.scala 143:103:@16714.4]
  assign _T_70138 = _T_70137[5:0]; // @[Modules.scala 143:103:@16715.4]
  assign _T_70139 = $signed(_T_70138); // @[Modules.scala 143:103:@16716.4]
  assign _T_70143 = $signed(4'sh1) * $signed(io_in_258); // @[Modules.scala 144:80:@16719.4]
  assign _T_70144 = $signed(_T_57864) + $signed(_T_70143); // @[Modules.scala 143:103:@16720.4]
  assign _T_70145 = _T_70144[5:0]; // @[Modules.scala 143:103:@16721.4]
  assign _T_70146 = $signed(_T_70145); // @[Modules.scala 143:103:@16722.4]
  assign _T_70148 = $signed(4'sh1) * $signed(io_in_259); // @[Modules.scala 143:74:@16724.4]
  assign _T_70151 = $signed(_T_70148) + $signed(_T_54824); // @[Modules.scala 143:103:@16726.4]
  assign _T_70152 = _T_70151[5:0]; // @[Modules.scala 143:103:@16727.4]
  assign _T_70153 = $signed(_T_70152); // @[Modules.scala 143:103:@16728.4]
  assign _T_70158 = $signed(_T_64019) + $signed(_T_60922); // @[Modules.scala 143:103:@16732.4]
  assign _T_70159 = _T_70158[5:0]; // @[Modules.scala 143:103:@16733.4]
  assign _T_70160 = $signed(_T_70159); // @[Modules.scala 143:103:@16734.4]
  assign _T_70186 = $signed(_T_57892) + $signed(_T_57899); // @[Modules.scala 143:103:@16756.4]
  assign _T_70187 = _T_70186[5:0]; // @[Modules.scala 143:103:@16757.4]
  assign _T_70188 = $signed(_T_70187); // @[Modules.scala 143:103:@16758.4]
  assign _T_70192 = $signed(4'sh1) * $signed(io_in_273); // @[Modules.scala 144:80:@16761.4]
  assign _T_70193 = $signed(_T_57904) + $signed(_T_70192); // @[Modules.scala 143:103:@16762.4]
  assign _T_70194 = _T_70193[5:0]; // @[Modules.scala 143:103:@16763.4]
  assign _T_70195 = $signed(_T_70194); // @[Modules.scala 143:103:@16764.4]
  assign _T_70200 = $signed(_T_64061) + $signed(_T_64066); // @[Modules.scala 143:103:@16768.4]
  assign _T_70201 = _T_70200[5:0]; // @[Modules.scala 143:103:@16769.4]
  assign _T_70202 = $signed(_T_70201); // @[Modules.scala 143:103:@16770.4]
  assign _T_70207 = $signed(_T_64068) + $signed(_T_64073); // @[Modules.scala 143:103:@16774.4]
  assign _T_70208 = _T_70207[5:0]; // @[Modules.scala 143:103:@16775.4]
  assign _T_70209 = $signed(_T_70208); // @[Modules.scala 143:103:@16776.4]
  assign _T_70213 = $signed(4'sh1) * $signed(io_in_279); // @[Modules.scala 144:80:@16779.4]
  assign _T_70214 = $signed(_T_64075) + $signed(_T_70213); // @[Modules.scala 143:103:@16780.4]
  assign _T_70215 = _T_70214[5:0]; // @[Modules.scala 143:103:@16781.4]
  assign _T_70216 = $signed(_T_70215); // @[Modules.scala 143:103:@16782.4]
  assign _T_70220 = $signed(-4'sh1) * $signed(io_in_281); // @[Modules.scala 144:80:@16785.4]
  assign _GEN_380 = {{1{_T_70220[4]}},_T_70220}; // @[Modules.scala 143:103:@16786.4]
  assign _T_70221 = $signed(_T_57927) + $signed(_GEN_380); // @[Modules.scala 143:103:@16786.4]
  assign _T_70222 = _T_70221[5:0]; // @[Modules.scala 143:103:@16787.4]
  assign _T_70223 = $signed(_T_70222); // @[Modules.scala 143:103:@16788.4]
  assign _T_70235 = $signed(_T_67200) + $signed(_T_64108); // @[Modules.scala 143:103:@16798.4]
  assign _T_70236 = _T_70235[5:0]; // @[Modules.scala 143:103:@16799.4]
  assign _T_70237 = $signed(_T_70236); // @[Modules.scala 143:103:@16800.4]
  assign _T_70242 = $signed(_T_61004) + $signed(_T_64115); // @[Modules.scala 143:103:@16804.4]
  assign _T_70243 = _T_70242[5:0]; // @[Modules.scala 143:103:@16805.4]
  assign _T_70244 = $signed(_T_70243); // @[Modules.scala 143:103:@16806.4]
  assign _T_70249 = $signed(_T_61006) + $signed(_T_64122); // @[Modules.scala 143:103:@16810.4]
  assign _T_70250 = _T_70249[5:0]; // @[Modules.scala 143:103:@16811.4]
  assign _T_70251 = $signed(_T_70250); // @[Modules.scala 143:103:@16812.4]
  assign _T_70256 = $signed(_T_64124) + $signed(_GEN_25); // @[Modules.scala 143:103:@16816.4]
  assign _T_70257 = _T_70256[5:0]; // @[Modules.scala 143:103:@16817.4]
  assign _T_70258 = $signed(_T_70257); // @[Modules.scala 143:103:@16818.4]
  assign _T_70270 = $signed(_T_57983) + $signed(_T_57988); // @[Modules.scala 143:103:@16828.4]
  assign _T_70271 = _T_70270[5:0]; // @[Modules.scala 143:103:@16829.4]
  assign _T_70272 = $signed(_T_70271); // @[Modules.scala 143:103:@16830.4]
  assign _T_70277 = $signed(_T_57990) + $signed(_T_67247); // @[Modules.scala 143:103:@16834.4]
  assign _T_70278 = _T_70277[5:0]; // @[Modules.scala 143:103:@16835.4]
  assign _T_70279 = $signed(_T_70278); // @[Modules.scala 143:103:@16836.4]
  assign _T_70281 = $signed(4'sh1) * $signed(io_in_303); // @[Modules.scala 143:74:@16838.4]
  assign _T_70284 = $signed(_T_70281) + $signed(_T_64164); // @[Modules.scala 143:103:@16840.4]
  assign _T_70285 = _T_70284[5:0]; // @[Modules.scala 143:103:@16841.4]
  assign _T_70286 = $signed(_T_70285); // @[Modules.scala 143:103:@16842.4]
  assign _T_70291 = $signed(_T_64166) + $signed(_T_64171); // @[Modules.scala 143:103:@16846.4]
  assign _T_70292 = _T_70291[5:0]; // @[Modules.scala 143:103:@16847.4]
  assign _T_70293 = $signed(_T_70292); // @[Modules.scala 143:103:@16848.4]
  assign _T_70319 = $signed(_T_55006) + $signed(_T_55013); // @[Modules.scala 143:103:@16870.4]
  assign _T_70320 = _T_70319[4:0]; // @[Modules.scala 143:103:@16871.4]
  assign _T_70321 = $signed(_T_70320); // @[Modules.scala 143:103:@16872.4]
  assign _GEN_382 = {{1{_T_61104[4]}},_T_61104}; // @[Modules.scala 143:103:@16876.4]
  assign _T_70326 = $signed(_T_61088) + $signed(_GEN_382); // @[Modules.scala 143:103:@16876.4]
  assign _T_70327 = _T_70326[5:0]; // @[Modules.scala 143:103:@16877.4]
  assign _T_70328 = $signed(_T_70327); // @[Modules.scala 143:103:@16878.4]
  assign _T_70333 = $signed(_GEN_169) + $signed(_T_58072); // @[Modules.scala 143:103:@16882.4]
  assign _T_70334 = _T_70333[5:0]; // @[Modules.scala 143:103:@16883.4]
  assign _T_70335 = $signed(_T_70334); // @[Modules.scala 143:103:@16884.4]
  assign _T_70340 = $signed(_T_58074) + $signed(_T_58079); // @[Modules.scala 143:103:@16888.4]
  assign _T_70341 = _T_70340[5:0]; // @[Modules.scala 143:103:@16889.4]
  assign _T_70342 = $signed(_T_70341); // @[Modules.scala 143:103:@16890.4]
  assign _T_70347 = $signed(_T_55055) + $signed(_T_55060); // @[Modules.scala 143:103:@16894.4]
  assign _T_70348 = _T_70347[4:0]; // @[Modules.scala 143:103:@16895.4]
  assign _T_70349 = $signed(_T_70348); // @[Modules.scala 143:103:@16896.4]
  assign _T_70351 = $signed(4'sh1) * $signed(io_in_331); // @[Modules.scala 143:74:@16898.4]
  assign _T_70353 = $signed(4'sh1) * $signed(io_in_332); // @[Modules.scala 144:80:@16899.4]
  assign _T_70354 = $signed(_T_70351) + $signed(_T_70353); // @[Modules.scala 143:103:@16900.4]
  assign _T_70355 = _T_70354[5:0]; // @[Modules.scala 143:103:@16901.4]
  assign _T_70356 = $signed(_T_70355); // @[Modules.scala 143:103:@16902.4]
  assign _T_70368 = $signed(_T_67340) + $signed(_T_55074); // @[Modules.scala 143:103:@16912.4]
  assign _T_70369 = _T_70368[4:0]; // @[Modules.scala 143:103:@16913.4]
  assign _T_70370 = $signed(_T_70369); // @[Modules.scala 143:103:@16914.4]
  assign _T_70382 = $signed(_T_58116) + $signed(_T_58121); // @[Modules.scala 143:103:@16924.4]
  assign _T_70383 = _T_70382[5:0]; // @[Modules.scala 143:103:@16925.4]
  assign _T_70384 = $signed(_T_70383); // @[Modules.scala 143:103:@16926.4]
  assign _GEN_384 = {{1{_T_55111[4]}},_T_55111}; // @[Modules.scala 143:103:@16942.4]
  assign _T_70403 = $signed(_GEN_384) + $signed(_T_61181); // @[Modules.scala 143:103:@16942.4]
  assign _T_70404 = _T_70403[5:0]; // @[Modules.scala 143:103:@16943.4]
  assign _T_70405 = $signed(_T_70404); // @[Modules.scala 143:103:@16944.4]
  assign _T_70410 = $signed(_T_55118) + $signed(_T_61188); // @[Modules.scala 143:103:@16948.4]
  assign _T_70411 = _T_70410[4:0]; // @[Modules.scala 143:103:@16949.4]
  assign _T_70412 = $signed(_T_70411); // @[Modules.scala 143:103:@16950.4]
  assign _T_70414 = $signed(-4'sh1) * $signed(io_in_351); // @[Modules.scala 143:74:@16952.4]
  assign _T_70417 = $signed(_T_70414) + $signed(_T_55130); // @[Modules.scala 143:103:@16954.4]
  assign _T_70418 = _T_70417[4:0]; // @[Modules.scala 143:103:@16955.4]
  assign _T_70419 = $signed(_T_70418); // @[Modules.scala 143:103:@16956.4]
  assign _T_70466 = $signed(_T_55172) + $signed(_T_58200); // @[Modules.scala 143:103:@16996.4]
  assign _T_70467 = _T_70466[5:0]; // @[Modules.scala 143:103:@16997.4]
  assign _T_70468 = $signed(_T_70467); // @[Modules.scala 143:103:@16998.4]
  assign _T_70473 = $signed(_T_55181) + $signed(_T_55186); // @[Modules.scala 143:103:@17002.4]
  assign _T_70474 = _T_70473[4:0]; // @[Modules.scala 143:103:@17003.4]
  assign _T_70475 = $signed(_T_70474); // @[Modules.scala 143:103:@17004.4]
  assign _T_70480 = $signed(_T_55188) + $signed(_T_55193); // @[Modules.scala 143:103:@17008.4]
  assign _T_70481 = _T_70480[4:0]; // @[Modules.scala 143:103:@17009.4]
  assign _T_70482 = $signed(_T_70481); // @[Modules.scala 143:103:@17010.4]
  assign _T_70487 = $signed(_T_61277) + $signed(_GEN_175); // @[Modules.scala 143:103:@17014.4]
  assign _T_70488 = _T_70487[5:0]; // @[Modules.scala 143:103:@17015.4]
  assign _T_70489 = $signed(_T_70488); // @[Modules.scala 143:103:@17016.4]
  assign _T_70491 = $signed(-4'sh1) * $signed(io_in_379); // @[Modules.scala 143:74:@17018.4]
  assign _GEN_387 = {{1{_T_70491[4]}},_T_70491}; // @[Modules.scala 143:103:@17020.4]
  assign _T_70494 = $signed(_GEN_387) + $signed(_T_55221); // @[Modules.scala 143:103:@17020.4]
  assign _T_70495 = _T_70494[5:0]; // @[Modules.scala 143:103:@17021.4]
  assign _T_70496 = $signed(_T_70495); // @[Modules.scala 143:103:@17022.4]
  assign _GEN_388 = {{1{_T_58254[4]}},_T_58254}; // @[Modules.scala 143:103:@17026.4]
  assign _T_70501 = $signed(_T_58249) + $signed(_GEN_388); // @[Modules.scala 143:103:@17026.4]
  assign _T_70502 = _T_70501[5:0]; // @[Modules.scala 143:103:@17027.4]
  assign _T_70503 = $signed(_T_70502); // @[Modules.scala 143:103:@17028.4]
  assign _GEN_389 = {{1{_T_58263[4]}},_T_58263}; // @[Modules.scala 143:103:@17038.4]
  assign _T_70515 = $signed(_GEN_389) + $signed(_T_58268); // @[Modules.scala 143:103:@17038.4]
  assign _T_70516 = _T_70515[5:0]; // @[Modules.scala 143:103:@17039.4]
  assign _T_70517 = $signed(_T_70516); // @[Modules.scala 143:103:@17040.4]
  assign _T_70522 = $signed(_T_58270) + $signed(_T_55244); // @[Modules.scala 143:103:@17044.4]
  assign _T_70523 = _T_70522[5:0]; // @[Modules.scala 143:103:@17045.4]
  assign _T_70524 = $signed(_T_70523); // @[Modules.scala 143:103:@17046.4]
  assign _T_70529 = $signed(_T_58277) + $signed(_T_55251); // @[Modules.scala 143:103:@17050.4]
  assign _T_70530 = _T_70529[4:0]; // @[Modules.scala 143:103:@17051.4]
  assign _T_70531 = $signed(_T_70530); // @[Modules.scala 143:103:@17052.4]
  assign _T_70533 = $signed(-4'sh1) * $signed(io_in_395); // @[Modules.scala 143:74:@17054.4]
  assign _T_70536 = $signed(_T_70533) + $signed(_T_55263); // @[Modules.scala 143:103:@17056.4]
  assign _T_70537 = _T_70536[4:0]; // @[Modules.scala 143:103:@17057.4]
  assign _T_70538 = $signed(_T_70537); // @[Modules.scala 143:103:@17058.4]
  assign _T_70543 = $signed(_T_55265) + $signed(_T_55270); // @[Modules.scala 143:103:@17062.4]
  assign _T_70544 = _T_70543[4:0]; // @[Modules.scala 143:103:@17063.4]
  assign _T_70545 = $signed(_T_70544); // @[Modules.scala 143:103:@17064.4]
  assign _T_70550 = $signed(_T_55272) + $signed(_T_55277); // @[Modules.scala 143:103:@17068.4]
  assign _T_70551 = _T_70550[4:0]; // @[Modules.scala 143:103:@17069.4]
  assign _T_70552 = $signed(_T_70551); // @[Modules.scala 143:103:@17070.4]
  assign _T_70557 = $signed(_T_55279) + $signed(_T_55284); // @[Modules.scala 143:103:@17074.4]
  assign _T_70558 = _T_70557[4:0]; // @[Modules.scala 143:103:@17075.4]
  assign _T_70559 = $signed(_T_70558); // @[Modules.scala 143:103:@17076.4]
  assign _T_70570 = $signed(-4'sh1) * $signed(io_in_406); // @[Modules.scala 144:80:@17085.4]
  assign _T_70571 = $signed(_T_67550) + $signed(_T_70570); // @[Modules.scala 143:103:@17086.4]
  assign _T_70572 = _T_70571[4:0]; // @[Modules.scala 143:103:@17087.4]
  assign _T_70573 = $signed(_T_70572); // @[Modules.scala 143:103:@17088.4]
  assign _T_70575 = $signed(-4'sh1) * $signed(io_in_407); // @[Modules.scala 143:74:@17090.4]
  assign _GEN_390 = {{1{_T_70575[4]}},_T_70575}; // @[Modules.scala 143:103:@17092.4]
  assign _T_70578 = $signed(_GEN_390) + $signed(_T_61382); // @[Modules.scala 143:103:@17092.4]
  assign _T_70579 = _T_70578[5:0]; // @[Modules.scala 143:103:@17093.4]
  assign _T_70580 = $signed(_T_70579); // @[Modules.scala 143:103:@17094.4]
  assign _T_70584 = $signed(-4'sh1) * $signed(io_in_410); // @[Modules.scala 144:80:@17097.4]
  assign _GEN_391 = {{1{_T_70584[4]}},_T_70584}; // @[Modules.scala 143:103:@17098.4]
  assign _T_70585 = $signed(_T_61384) + $signed(_GEN_391); // @[Modules.scala 143:103:@17098.4]
  assign _T_70586 = _T_70585[5:0]; // @[Modules.scala 143:103:@17099.4]
  assign _T_70587 = $signed(_T_70586); // @[Modules.scala 143:103:@17100.4]
  assign _T_70589 = $signed(-4'sh1) * $signed(io_in_411); // @[Modules.scala 143:74:@17102.4]
  assign _T_70592 = $signed(_T_70589) + $signed(_T_58331); // @[Modules.scala 143:103:@17104.4]
  assign _T_70593 = _T_70592[4:0]; // @[Modules.scala 143:103:@17105.4]
  assign _T_70594 = $signed(_T_70593); // @[Modules.scala 143:103:@17106.4]
  assign _T_70599 = $signed(_T_58333) + $signed(_T_58338); // @[Modules.scala 143:103:@17110.4]
  assign _T_70600 = _T_70599[4:0]; // @[Modules.scala 143:103:@17111.4]
  assign _T_70601 = $signed(_T_70600); // @[Modules.scala 143:103:@17112.4]
  assign _T_70605 = $signed(4'sh1) * $signed(io_in_417); // @[Modules.scala 144:80:@17115.4]
  assign _GEN_392 = {{1{_T_58340[4]}},_T_58340}; // @[Modules.scala 143:103:@17116.4]
  assign _T_70606 = $signed(_GEN_392) + $signed(_T_70605); // @[Modules.scala 143:103:@17116.4]
  assign _T_70607 = _T_70606[5:0]; // @[Modules.scala 143:103:@17117.4]
  assign _T_70608 = $signed(_T_70607); // @[Modules.scala 143:103:@17118.4]
  assign _T_70613 = $signed(_T_55326) + $signed(_T_67585); // @[Modules.scala 143:103:@17122.4]
  assign _T_70614 = _T_70613[5:0]; // @[Modules.scala 143:103:@17123.4]
  assign _T_70615 = $signed(_T_70614); // @[Modules.scala 143:103:@17124.4]
  assign _T_70620 = $signed(_T_55328) + $signed(_GEN_43); // @[Modules.scala 143:103:@17128.4]
  assign _T_70621 = _T_70620[5:0]; // @[Modules.scala 143:103:@17129.4]
  assign _T_70622 = $signed(_T_70621); // @[Modules.scala 143:103:@17130.4]
  assign _T_70626 = $signed(-4'sh1) * $signed(io_in_423); // @[Modules.scala 144:80:@17133.4]
  assign _T_70627 = $signed(_T_67597) + $signed(_T_70626); // @[Modules.scala 143:103:@17134.4]
  assign _T_70628 = _T_70627[4:0]; // @[Modules.scala 143:103:@17135.4]
  assign _T_70629 = $signed(_T_70628); // @[Modules.scala 143:103:@17136.4]
  assign _T_70634 = $signed(_T_55342) + $signed(_T_55347); // @[Modules.scala 143:103:@17140.4]
  assign _T_70635 = _T_70634[4:0]; // @[Modules.scala 143:103:@17141.4]
  assign _T_70636 = $signed(_T_70635); // @[Modules.scala 143:103:@17142.4]
  assign _T_70641 = $signed(_T_55349) + $signed(_T_55354); // @[Modules.scala 143:103:@17146.4]
  assign _T_70642 = _T_70641[4:0]; // @[Modules.scala 143:103:@17147.4]
  assign _T_70643 = $signed(_T_70642); // @[Modules.scala 143:103:@17148.4]
  assign _GEN_394 = {{1{_T_58375[4]}},_T_58375}; // @[Modules.scala 143:103:@17152.4]
  assign _T_70648 = $signed(_GEN_394) + $signed(_T_61445); // @[Modules.scala 143:103:@17152.4]
  assign _T_70649 = _T_70648[5:0]; // @[Modules.scala 143:103:@17153.4]
  assign _T_70650 = $signed(_T_70649); // @[Modules.scala 143:103:@17154.4]
  assign _T_70661 = $signed(-4'sh1) * $signed(io_in_434); // @[Modules.scala 144:80:@17163.4]
  assign _T_70662 = $signed(_T_61454) + $signed(_T_70661); // @[Modules.scala 143:103:@17164.4]
  assign _T_70663 = _T_70662[4:0]; // @[Modules.scala 143:103:@17165.4]
  assign _T_70664 = $signed(_T_70663); // @[Modules.scala 143:103:@17166.4]
  assign _T_70666 = $signed(-4'sh1) * $signed(io_in_435); // @[Modules.scala 143:74:@17168.4]
  assign _GEN_395 = {{1{_T_70666[4]}},_T_70666}; // @[Modules.scala 143:103:@17170.4]
  assign _T_70669 = $signed(_GEN_395) + $signed(_T_61468); // @[Modules.scala 143:103:@17170.4]
  assign _T_70670 = _T_70669[5:0]; // @[Modules.scala 143:103:@17171.4]
  assign _T_70671 = $signed(_T_70670); // @[Modules.scala 143:103:@17172.4]
  assign _T_70704 = $signed(_T_58424) + $signed(_GEN_112); // @[Modules.scala 143:103:@17200.4]
  assign _T_70705 = _T_70704[5:0]; // @[Modules.scala 143:103:@17201.4]
  assign _T_70706 = $signed(_T_70705); // @[Modules.scala 143:103:@17202.4]
  assign _T_70718 = $signed(_T_58438) + $signed(_GEN_325); // @[Modules.scala 143:103:@17212.4]
  assign _T_70719 = _T_70718[5:0]; // @[Modules.scala 143:103:@17213.4]
  assign _T_70720 = $signed(_T_70719); // @[Modules.scala 143:103:@17214.4]
  assign _T_70725 = $signed(_GEN_247) + $signed(_T_55440); // @[Modules.scala 143:103:@17218.4]
  assign _T_70726 = _T_70725[5:0]; // @[Modules.scala 143:103:@17219.4]
  assign _T_70727 = $signed(_T_70726); // @[Modules.scala 143:103:@17220.4]
  assign _GEN_400 = {{1{_T_58464[4]}},_T_58464}; // @[Modules.scala 143:103:@17224.4]
  assign _T_70732 = $signed(_GEN_400) + $signed(_T_64649); // @[Modules.scala 143:103:@17224.4]
  assign _T_70733 = _T_70732[5:0]; // @[Modules.scala 143:103:@17225.4]
  assign _T_70734 = $signed(_T_70733); // @[Modules.scala 143:103:@17226.4]
  assign _T_70739 = $signed(_T_61536) + $signed(_T_67695); // @[Modules.scala 143:103:@17230.4]
  assign _T_70740 = _T_70739[4:0]; // @[Modules.scala 143:103:@17231.4]
  assign _T_70741 = $signed(_T_70740); // @[Modules.scala 143:103:@17232.4]
  assign _GEN_402 = {{1{_T_64675[4]}},_T_64675}; // @[Modules.scala 143:103:@17248.4]
  assign _T_70760 = $signed(_GEN_402) + $signed(_T_55473); // @[Modules.scala 143:103:@17248.4]
  assign _T_70761 = _T_70760[5:0]; // @[Modules.scala 143:103:@17249.4]
  assign _T_70762 = $signed(_T_70761); // @[Modules.scala 143:103:@17250.4]
  assign _T_70766 = $signed(4'sh1) * $signed(io_in_472); // @[Modules.scala 144:80:@17253.4]
  assign _T_70767 = $signed(_GEN_52) + $signed(_T_70766); // @[Modules.scala 143:103:@17254.4]
  assign _T_70768 = _T_70767[5:0]; // @[Modules.scala 143:103:@17255.4]
  assign _T_70769 = $signed(_T_70768); // @[Modules.scala 143:103:@17256.4]
  assign _T_70780 = $signed(-4'sh1) * $signed(io_in_476); // @[Modules.scala 144:80:@17265.4]
  assign _GEN_404 = {{1{_T_70780[4]}},_T_70780}; // @[Modules.scala 143:103:@17266.4]
  assign _T_70781 = $signed(_T_58501) + $signed(_GEN_404); // @[Modules.scala 143:103:@17266.4]
  assign _T_70782 = _T_70781[5:0]; // @[Modules.scala 143:103:@17267.4]
  assign _T_70783 = $signed(_T_70782); // @[Modules.scala 143:103:@17268.4]
  assign _T_70799 = $signed(4'sh1) * $signed(io_in_481); // @[Modules.scala 143:74:@17282.4]
  assign _T_70802 = $signed(_T_70799) + $signed(_T_55501); // @[Modules.scala 143:103:@17284.4]
  assign _T_70803 = _T_70802[5:0]; // @[Modules.scala 143:103:@17285.4]
  assign _T_70804 = $signed(_T_70803); // @[Modules.scala 143:103:@17286.4]
  assign _T_70809 = $signed(_T_58527) + $signed(_T_58536); // @[Modules.scala 143:103:@17290.4]
  assign _T_70810 = _T_70809[4:0]; // @[Modules.scala 143:103:@17291.4]
  assign _T_70811 = $signed(_T_70810); // @[Modules.scala 143:103:@17292.4]
  assign _T_70815 = $signed(-4'sh1) * $signed(io_in_489); // @[Modules.scala 144:80:@17295.4]
  assign _T_70816 = $signed(_T_58541) + $signed(_T_70815); // @[Modules.scala 143:103:@17296.4]
  assign _T_70817 = _T_70816[4:0]; // @[Modules.scala 143:103:@17297.4]
  assign _T_70818 = $signed(_T_70817); // @[Modules.scala 143:103:@17298.4]
  assign _T_70829 = $signed(4'sh1) * $signed(io_in_493); // @[Modules.scala 144:80:@17307.4]
  assign _T_70830 = $signed(_T_61622) + $signed(_T_70829); // @[Modules.scala 143:103:@17308.4]
  assign _T_70831 = _T_70830[5:0]; // @[Modules.scala 143:103:@17309.4]
  assign _T_70832 = $signed(_T_70831); // @[Modules.scala 143:103:@17310.4]
  assign _T_70837 = $signed(_T_58557) + $signed(_T_55543); // @[Modules.scala 143:103:@17314.4]
  assign _T_70838 = _T_70837[5:0]; // @[Modules.scala 143:103:@17315.4]
  assign _T_70839 = $signed(_T_70838); // @[Modules.scala 143:103:@17316.4]
  assign _T_70844 = $signed(_T_55545) + $signed(_T_55550); // @[Modules.scala 143:103:@17320.4]
  assign _T_70845 = _T_70844[5:0]; // @[Modules.scala 143:103:@17321.4]
  assign _T_70846 = $signed(_T_70845); // @[Modules.scala 143:103:@17322.4]
  assign _T_70855 = $signed(-4'sh1) * $signed(io_in_505); // @[Modules.scala 143:74:@17330.4]
  assign _GEN_406 = {{1{_T_70855[4]}},_T_70855}; // @[Modules.scala 143:103:@17332.4]
  assign _T_70858 = $signed(_GEN_406) + $signed(_T_55566); // @[Modules.scala 143:103:@17332.4]
  assign _T_70859 = _T_70858[5:0]; // @[Modules.scala 143:103:@17333.4]
  assign _T_70860 = $signed(_T_70859); // @[Modules.scala 143:103:@17334.4]
  assign _T_70872 = $signed(_T_55578) + $signed(_T_64796); // @[Modules.scala 143:103:@17344.4]
  assign _T_70873 = _T_70872[5:0]; // @[Modules.scala 143:103:@17345.4]
  assign _T_70874 = $signed(_T_70873); // @[Modules.scala 143:103:@17346.4]
  assign _T_70876 = $signed(4'sh1) * $signed(io_in_511); // @[Modules.scala 143:74:@17348.4]
  assign _T_70879 = $signed(_T_70876) + $signed(_GEN_58); // @[Modules.scala 143:103:@17350.4]
  assign _T_70880 = _T_70879[5:0]; // @[Modules.scala 143:103:@17351.4]
  assign _T_70881 = $signed(_T_70880); // @[Modules.scala 143:103:@17352.4]
  assign _T_70897 = $signed(-4'sh1) * $signed(io_in_518); // @[Modules.scala 143:74:@17366.4]
  assign _GEN_408 = {{1{_T_70897[4]}},_T_70897}; // @[Modules.scala 143:103:@17368.4]
  assign _T_70900 = $signed(_GEN_408) + $signed(_T_58632); // @[Modules.scala 143:103:@17368.4]
  assign _T_70901 = _T_70900[5:0]; // @[Modules.scala 143:103:@17369.4]
  assign _T_70902 = $signed(_T_70901); // @[Modules.scala 143:103:@17370.4]
  assign _T_70904 = $signed(4'sh1) * $signed(io_in_520); // @[Modules.scala 143:74:@17372.4]
  assign _T_70907 = $signed(_T_70904) + $signed(_T_55615); // @[Modules.scala 143:103:@17374.4]
  assign _T_70908 = _T_70907[5:0]; // @[Modules.scala 143:103:@17375.4]
  assign _T_70909 = $signed(_T_70908); // @[Modules.scala 143:103:@17376.4]
  assign _T_70911 = $signed(4'sh1) * $signed(io_in_522); // @[Modules.scala 143:74:@17378.4]
  assign _GEN_409 = {{1{_T_64831[4]}},_T_64831}; // @[Modules.scala 143:103:@17380.4]
  assign _T_70914 = $signed(_T_70911) + $signed(_GEN_409); // @[Modules.scala 143:103:@17380.4]
  assign _T_70915 = _T_70914[5:0]; // @[Modules.scala 143:103:@17381.4]
  assign _T_70916 = $signed(_T_70915); // @[Modules.scala 143:103:@17382.4]
  assign _T_70918 = $signed(4'sh1) * $signed(io_in_525); // @[Modules.scala 143:74:@17384.4]
  assign _T_70921 = $signed(_T_70918) + $signed(_T_55627); // @[Modules.scala 143:103:@17386.4]
  assign _T_70922 = _T_70921[5:0]; // @[Modules.scala 143:103:@17387.4]
  assign _T_70923 = $signed(_T_70922); // @[Modules.scala 143:103:@17388.4]
  assign _T_70928 = $signed(_T_55629) + $signed(_T_55634); // @[Modules.scala 143:103:@17392.4]
  assign _T_70929 = _T_70928[5:0]; // @[Modules.scala 143:103:@17393.4]
  assign _T_70930 = $signed(_T_70929); // @[Modules.scala 143:103:@17394.4]
  assign _T_70935 = $signed(_T_55636) + $signed(_T_55641); // @[Modules.scala 143:103:@17398.4]
  assign _T_70936 = _T_70935[5:0]; // @[Modules.scala 143:103:@17399.4]
  assign _T_70937 = $signed(_T_70936); // @[Modules.scala 143:103:@17400.4]
  assign _T_70960 = $signed(4'sh1) * $signed(io_in_538); // @[Modules.scala 143:74:@17420.4]
  assign _T_70963 = $signed(_T_70960) + $signed(_T_55669); // @[Modules.scala 143:103:@17422.4]
  assign _T_70964 = _T_70963[5:0]; // @[Modules.scala 143:103:@17423.4]
  assign _T_70965 = $signed(_T_70964); // @[Modules.scala 143:103:@17424.4]
  assign _GEN_411 = {{1{_T_58688[4]}},_T_58688}; // @[Modules.scala 143:103:@17428.4]
  assign _T_70970 = $signed(_T_55671) + $signed(_GEN_411); // @[Modules.scala 143:103:@17428.4]
  assign _T_70971 = _T_70970[5:0]; // @[Modules.scala 143:103:@17429.4]
  assign _T_70972 = $signed(_T_70971); // @[Modules.scala 143:103:@17430.4]
  assign _T_70977 = $signed(_T_58690) + $signed(_T_58695); // @[Modules.scala 143:103:@17434.4]
  assign _T_70978 = _T_70977[4:0]; // @[Modules.scala 143:103:@17435.4]
  assign _T_70979 = $signed(_T_70978); // @[Modules.scala 143:103:@17436.4]
  assign _T_70984 = $signed(_T_58697) + $signed(_T_64906); // @[Modules.scala 143:103:@17440.4]
  assign _T_70985 = _T_70984[4:0]; // @[Modules.scala 143:103:@17441.4]
  assign _T_70986 = $signed(_T_70985); // @[Modules.scala 143:103:@17442.4]
  assign _T_70990 = $signed(4'sh1) * $signed(io_in_550); // @[Modules.scala 144:80:@17445.4]
  assign _T_70991 = $signed(_T_55704) + $signed(_T_70990); // @[Modules.scala 143:103:@17446.4]
  assign _T_70992 = _T_70991[5:0]; // @[Modules.scala 143:103:@17447.4]
  assign _T_70993 = $signed(_T_70992); // @[Modules.scala 143:103:@17448.4]
  assign _T_71002 = $signed(4'sh1) * $signed(io_in_553); // @[Modules.scala 143:74:@17456.4]
  assign _T_71004 = $signed(4'sh1) * $signed(io_in_554); // @[Modules.scala 144:80:@17457.4]
  assign _T_71005 = $signed(_T_71002) + $signed(_T_71004); // @[Modules.scala 143:103:@17458.4]
  assign _T_71006 = _T_71005[5:0]; // @[Modules.scala 143:103:@17459.4]
  assign _T_71007 = $signed(_T_71006); // @[Modules.scala 143:103:@17460.4]
  assign _T_71009 = $signed(4'sh1) * $signed(io_in_555); // @[Modules.scala 143:74:@17462.4]
  assign _T_71012 = $signed(_T_71009) + $signed(_T_55713); // @[Modules.scala 143:103:@17464.4]
  assign _T_71013 = _T_71012[5:0]; // @[Modules.scala 143:103:@17465.4]
  assign _T_71014 = $signed(_T_71013); // @[Modules.scala 143:103:@17466.4]
  assign _T_71026 = $signed(_T_55725) + $signed(_T_64948); // @[Modules.scala 143:103:@17476.4]
  assign _T_71027 = _T_71026[4:0]; // @[Modules.scala 143:103:@17477.4]
  assign _T_71028 = $signed(_T_71027); // @[Modules.scala 143:103:@17478.4]
  assign _T_71040 = $signed(_T_55734) + $signed(_T_55739); // @[Modules.scala 143:103:@17488.4]
  assign _T_71041 = _T_71040[5:0]; // @[Modules.scala 143:103:@17489.4]
  assign _T_71042 = $signed(_T_71041); // @[Modules.scala 143:103:@17490.4]
  assign _T_71047 = $signed(_T_55741) + $signed(_T_55746); // @[Modules.scala 143:103:@17494.4]
  assign _T_71048 = _T_71047[5:0]; // @[Modules.scala 143:103:@17495.4]
  assign _T_71049 = $signed(_T_71048); // @[Modules.scala 143:103:@17496.4]
  assign _GEN_414 = {{1{_T_58760[4]}},_T_58760}; // @[Modules.scala 143:103:@17506.4]
  assign _T_71061 = $signed(_GEN_414) + $signed(_T_55760); // @[Modules.scala 143:103:@17506.4]
  assign _T_71062 = _T_71061[5:0]; // @[Modules.scala 143:103:@17507.4]
  assign _T_71063 = $signed(_T_71062); // @[Modules.scala 143:103:@17508.4]
  assign _T_71068 = $signed(_T_64985) + $signed(_T_67991); // @[Modules.scala 143:103:@17512.4]
  assign _T_71069 = _T_71068[4:0]; // @[Modules.scala 143:103:@17513.4]
  assign _T_71070 = $signed(_T_71069); // @[Modules.scala 143:103:@17514.4]
  assign _T_71075 = $signed(_T_58774) + $signed(_T_58779); // @[Modules.scala 143:103:@17518.4]
  assign _T_71076 = _T_71075[4:0]; // @[Modules.scala 143:103:@17519.4]
  assign _T_71077 = $signed(_T_71076); // @[Modules.scala 143:103:@17520.4]
  assign _T_71082 = $signed(_T_55767) + $signed(_T_58786); // @[Modules.scala 143:103:@17524.4]
  assign _T_71083 = _T_71082[5:0]; // @[Modules.scala 143:103:@17525.4]
  assign _T_71084 = $signed(_T_71083); // @[Modules.scala 143:103:@17526.4]
  assign _T_71088 = $signed(4'sh1) * $signed(io_in_581); // @[Modules.scala 144:80:@17529.4]
  assign _T_71089 = $signed(_T_58788) + $signed(_T_71088); // @[Modules.scala 143:103:@17530.4]
  assign _T_71090 = _T_71089[5:0]; // @[Modules.scala 143:103:@17531.4]
  assign _T_71091 = $signed(_T_71090); // @[Modules.scala 143:103:@17532.4]
  assign _T_71096 = $signed(_T_65004) + $signed(_T_55776); // @[Modules.scala 143:103:@17536.4]
  assign _T_71097 = _T_71096[5:0]; // @[Modules.scala 143:103:@17537.4]
  assign _T_71098 = $signed(_T_71097); // @[Modules.scala 143:103:@17538.4]
  assign _T_71116 = $signed(-4'sh1) * $signed(io_in_589); // @[Modules.scala 144:80:@17553.4]
  assign _GEN_416 = {{1{_T_71116[4]}},_T_71116}; // @[Modules.scala 143:103:@17554.4]
  assign _T_71117 = $signed(_T_55790) + $signed(_GEN_416); // @[Modules.scala 143:103:@17554.4]
  assign _T_71118 = _T_71117[5:0]; // @[Modules.scala 143:103:@17555.4]
  assign _T_71119 = $signed(_T_71118); // @[Modules.scala 143:103:@17556.4]
  assign _T_71124 = $signed(_T_55797) + $signed(_T_55802); // @[Modules.scala 143:103:@17560.4]
  assign _T_71125 = _T_71124[5:0]; // @[Modules.scala 143:103:@17561.4]
  assign _T_71126 = $signed(_T_71125); // @[Modules.scala 143:103:@17562.4]
  assign _T_71131 = $signed(_T_55804) + $signed(_T_55809); // @[Modules.scala 143:103:@17566.4]
  assign _T_71132 = _T_71131[5:0]; // @[Modules.scala 143:103:@17567.4]
  assign _T_71133 = $signed(_T_71132); // @[Modules.scala 143:103:@17568.4]
  assign _T_71137 = $signed(4'sh1) * $signed(io_in_595); // @[Modules.scala 144:80:@17571.4]
  assign _T_71138 = $signed(_T_55811) + $signed(_T_71137); // @[Modules.scala 143:103:@17572.4]
  assign _T_71139 = _T_71138[5:0]; // @[Modules.scala 143:103:@17573.4]
  assign _T_71140 = $signed(_T_71139); // @[Modules.scala 143:103:@17574.4]
  assign _GEN_417 = {{1{_T_61916[4]}},_T_61916}; // @[Modules.scala 143:103:@17578.4]
  assign _T_71145 = $signed(_T_55816) + $signed(_GEN_417); // @[Modules.scala 143:103:@17578.4]
  assign _T_71146 = _T_71145[5:0]; // @[Modules.scala 143:103:@17579.4]
  assign _T_71147 = $signed(_T_71146); // @[Modules.scala 143:103:@17580.4]
  assign _T_71151 = $signed(-4'sh1) * $signed(io_in_599); // @[Modules.scala 144:80:@17583.4]
  assign _T_71152 = $signed(_T_61921) + $signed(_T_71151); // @[Modules.scala 143:103:@17584.4]
  assign _T_71153 = _T_71152[4:0]; // @[Modules.scala 143:103:@17585.4]
  assign _T_71154 = $signed(_T_71153); // @[Modules.scala 143:103:@17586.4]
  assign _T_71159 = $signed(_T_58844) + $signed(_T_58849); // @[Modules.scala 143:103:@17590.4]
  assign _T_71160 = _T_71159[4:0]; // @[Modules.scala 143:103:@17591.4]
  assign _T_71161 = $signed(_T_71160); // @[Modules.scala 143:103:@17592.4]
  assign _T_71163 = $signed(-4'sh1) * $signed(io_in_602); // @[Modules.scala 143:74:@17594.4]
  assign _T_71166 = $signed(_T_71163) + $signed(_T_68075); // @[Modules.scala 143:103:@17596.4]
  assign _T_71167 = _T_71166[4:0]; // @[Modules.scala 143:103:@17597.4]
  assign _T_71168 = $signed(_T_71167); // @[Modules.scala 143:103:@17598.4]
  assign _T_71173 = $signed(_T_65048) + $signed(_T_58851); // @[Modules.scala 143:103:@17602.4]
  assign _T_71174 = _T_71173[4:0]; // @[Modules.scala 143:103:@17603.4]
  assign _T_71175 = $signed(_T_71174); // @[Modules.scala 143:103:@17604.4]
  assign _T_71179 = $signed(4'sh1) * $signed(io_in_608); // @[Modules.scala 144:80:@17607.4]
  assign _T_71180 = $signed(_T_58858) + $signed(_T_71179); // @[Modules.scala 143:103:@17608.4]
  assign _T_71181 = _T_71180[5:0]; // @[Modules.scala 143:103:@17609.4]
  assign _T_71182 = $signed(_T_71181); // @[Modules.scala 143:103:@17610.4]
  assign _T_71187 = $signed(_T_55839) + $signed(_T_55844); // @[Modules.scala 143:103:@17614.4]
  assign _T_71188 = _T_71187[5:0]; // @[Modules.scala 143:103:@17615.4]
  assign _T_71189 = $signed(_T_71188); // @[Modules.scala 143:103:@17616.4]
  assign _T_71194 = $signed(_T_55846) + $signed(_T_55851); // @[Modules.scala 143:103:@17620.4]
  assign _T_71195 = _T_71194[5:0]; // @[Modules.scala 143:103:@17621.4]
  assign _T_71196 = $signed(_T_71195); // @[Modules.scala 143:103:@17622.4]
  assign _T_71201 = $signed(_T_58879) + $signed(_T_65074); // @[Modules.scala 143:103:@17626.4]
  assign _T_71202 = _T_71201[4:0]; // @[Modules.scala 143:103:@17627.4]
  assign _T_71203 = $signed(_T_71202); // @[Modules.scala 143:103:@17628.4]
  assign _T_71208 = $signed(_T_55860) + $signed(_T_55867); // @[Modules.scala 143:103:@17632.4]
  assign _T_71209 = _T_71208[5:0]; // @[Modules.scala 143:103:@17633.4]
  assign _T_71210 = $signed(_T_71209); // @[Modules.scala 143:103:@17634.4]
  assign _T_71221 = $signed(4'sh1) * $signed(io_in_623); // @[Modules.scala 144:80:@17643.4]
  assign _GEN_418 = {{1{_T_61986[4]}},_T_61986}; // @[Modules.scala 143:103:@17644.4]
  assign _T_71222 = $signed(_GEN_418) + $signed(_T_71221); // @[Modules.scala 143:103:@17644.4]
  assign _T_71223 = _T_71222[5:0]; // @[Modules.scala 143:103:@17645.4]
  assign _T_71224 = $signed(_T_71223); // @[Modules.scala 143:103:@17646.4]
  assign _T_71235 = $signed(4'sh1) * $signed(io_in_627); // @[Modules.scala 144:80:@17655.4]
  assign _T_71236 = $signed(_T_58919) + $signed(_T_71235); // @[Modules.scala 143:103:@17656.4]
  assign _T_71237 = _T_71236[5:0]; // @[Modules.scala 143:103:@17657.4]
  assign _T_71238 = $signed(_T_71237); // @[Modules.scala 143:103:@17658.4]
  assign _T_71240 = $signed(4'sh1) * $signed(io_in_628); // @[Modules.scala 143:74:@17660.4]
  assign _T_71242 = $signed(4'sh1) * $signed(io_in_629); // @[Modules.scala 144:80:@17661.4]
  assign _T_71243 = $signed(_T_71240) + $signed(_T_71242); // @[Modules.scala 143:103:@17662.4]
  assign _T_71244 = _T_71243[5:0]; // @[Modules.scala 143:103:@17663.4]
  assign _T_71245 = $signed(_T_71244); // @[Modules.scala 143:103:@17664.4]
  assign _T_71247 = $signed(4'sh1) * $signed(io_in_630); // @[Modules.scala 143:74:@17666.4]
  assign _T_71250 = $signed(_T_71247) + $signed(_T_65125); // @[Modules.scala 143:103:@17668.4]
  assign _T_71251 = _T_71250[5:0]; // @[Modules.scala 143:103:@17669.4]
  assign _T_71252 = $signed(_T_71251); // @[Modules.scala 143:103:@17670.4]
  assign _GEN_419 = {{1{_T_55914[4]}},_T_55914}; // @[Modules.scala 143:103:@17674.4]
  assign _T_71257 = $signed(_GEN_419) + $signed(_T_62026); // @[Modules.scala 143:103:@17674.4]
  assign _T_71258 = _T_71257[5:0]; // @[Modules.scala 143:103:@17675.4]
  assign _T_71259 = $signed(_T_71258); // @[Modules.scala 143:103:@17676.4]
  assign _T_71264 = $signed(_T_55921) + $signed(_T_55930); // @[Modules.scala 143:103:@17680.4]
  assign _T_71265 = _T_71264[5:0]; // @[Modules.scala 143:103:@17681.4]
  assign _T_71266 = $signed(_T_71265); // @[Modules.scala 143:103:@17682.4]
  assign _T_71271 = $signed(_T_55935) + $signed(_GEN_344); // @[Modules.scala 143:103:@17686.4]
  assign _T_71272 = _T_71271[5:0]; // @[Modules.scala 143:103:@17687.4]
  assign _T_71273 = $signed(_T_71272); // @[Modules.scala 143:103:@17688.4]
  assign _T_71278 = $signed(_T_65165) + $signed(_T_68194); // @[Modules.scala 143:103:@17692.4]
  assign _T_71279 = _T_71278[4:0]; // @[Modules.scala 143:103:@17693.4]
  assign _T_71280 = $signed(_T_71279); // @[Modules.scala 143:103:@17694.4]
  assign _T_71285 = $signed(_T_55951) + $signed(_T_55956); // @[Modules.scala 143:103:@17698.4]
  assign _T_71286 = _T_71285[5:0]; // @[Modules.scala 143:103:@17699.4]
  assign _T_71287 = $signed(_T_71286); // @[Modules.scala 143:103:@17700.4]
  assign _T_71299 = $signed(_T_62063) + $signed(_T_55970); // @[Modules.scala 143:103:@17710.4]
  assign _T_71300 = _T_71299[4:0]; // @[Modules.scala 143:103:@17711.4]
  assign _T_71301 = $signed(_T_71300); // @[Modules.scala 143:103:@17712.4]
  assign _T_71303 = $signed(4'sh1) * $signed(io_in_653); // @[Modules.scala 143:74:@17714.4]
  assign _T_71306 = $signed(_T_71303) + $signed(_T_68220); // @[Modules.scala 143:103:@17716.4]
  assign _T_71307 = _T_71306[5:0]; // @[Modules.scala 143:103:@17717.4]
  assign _T_71308 = $signed(_T_71307); // @[Modules.scala 143:103:@17718.4]
  assign _T_71317 = $signed(4'sh1) * $signed(io_in_657); // @[Modules.scala 143:74:@17726.4]
  assign _T_71320 = $signed(_T_71317) + $signed(_T_65193); // @[Modules.scala 143:103:@17728.4]
  assign _T_71321 = _T_71320[5:0]; // @[Modules.scala 143:103:@17729.4]
  assign _T_71322 = $signed(_T_71321); // @[Modules.scala 143:103:@17730.4]
  assign _T_71327 = $signed(_T_65195) + $signed(_T_65200); // @[Modules.scala 143:103:@17734.4]
  assign _T_71328 = _T_71327[5:0]; // @[Modules.scala 143:103:@17735.4]
  assign _T_71329 = $signed(_T_71328); // @[Modules.scala 143:103:@17736.4]
  assign _T_71334 = $signed(_T_59003) + $signed(_GEN_348); // @[Modules.scala 143:103:@17740.4]
  assign _T_71335 = _T_71334[5:0]; // @[Modules.scala 143:103:@17741.4]
  assign _T_71336 = $signed(_T_71335); // @[Modules.scala 143:103:@17742.4]
  assign _T_71348 = $signed(_T_56014) + $signed(_T_62126); // @[Modules.scala 143:103:@17752.4]
  assign _T_71349 = _T_71348[4:0]; // @[Modules.scala 143:103:@17753.4]
  assign _T_71350 = $signed(_T_71349); // @[Modules.scala 143:103:@17754.4]
  assign _T_71354 = $signed(-4'sh1) * $signed(io_in_673); // @[Modules.scala 144:80:@17757.4]
  assign _T_71355 = $signed(_T_65230) + $signed(_T_71354); // @[Modules.scala 143:103:@17758.4]
  assign _T_71356 = _T_71355[4:0]; // @[Modules.scala 143:103:@17759.4]
  assign _T_71357 = $signed(_T_71356); // @[Modules.scala 143:103:@17760.4]
  assign _T_71362 = $signed(_GEN_67) + $signed(_T_56033); // @[Modules.scala 143:103:@17764.4]
  assign _T_71363 = _T_71362[5:0]; // @[Modules.scala 143:103:@17765.4]
  assign _T_71364 = $signed(_T_71363); // @[Modules.scala 143:103:@17766.4]
  assign _T_71369 = $signed(_T_56035) + $signed(_T_56042); // @[Modules.scala 143:103:@17770.4]
  assign _T_71370 = _T_71369[5:0]; // @[Modules.scala 143:103:@17771.4]
  assign _T_71371 = $signed(_T_71370); // @[Modules.scala 143:103:@17772.4]
  assign _T_71383 = $signed(_T_59059) + $signed(_T_62159); // @[Modules.scala 143:103:@17782.4]
  assign _T_71384 = _T_71383[5:0]; // @[Modules.scala 143:103:@17783.4]
  assign _T_71385 = $signed(_T_71384); // @[Modules.scala 143:103:@17784.4]
  assign _T_71389 = $signed(4'sh1) * $signed(io_in_684); // @[Modules.scala 144:80:@17787.4]
  assign _T_71390 = $signed(_T_59061) + $signed(_T_71389); // @[Modules.scala 143:103:@17788.4]
  assign _T_71391 = _T_71390[5:0]; // @[Modules.scala 143:103:@17789.4]
  assign _T_71392 = $signed(_T_71391); // @[Modules.scala 143:103:@17790.4]
  assign _T_71394 = $signed(4'sh1) * $signed(io_in_685); // @[Modules.scala 143:74:@17792.4]
  assign _T_71396 = $signed(4'sh1) * $signed(io_in_686); // @[Modules.scala 144:80:@17793.4]
  assign _T_71397 = $signed(_T_71394) + $signed(_T_71396); // @[Modules.scala 143:103:@17794.4]
  assign _T_71398 = _T_71397[5:0]; // @[Modules.scala 143:103:@17795.4]
  assign _T_71399 = $signed(_T_71398); // @[Modules.scala 143:103:@17796.4]
  assign _T_71404 = $signed(_T_59075) + $signed(_T_59080); // @[Modules.scala 143:103:@17800.4]
  assign _T_71405 = _T_71404[5:0]; // @[Modules.scala 143:103:@17801.4]
  assign _T_71406 = $signed(_T_71405); // @[Modules.scala 143:103:@17802.4]
  assign _T_71411 = $signed(_T_59082) + $signed(_T_59087); // @[Modules.scala 143:103:@17806.4]
  assign _T_71412 = _T_71411[5:0]; // @[Modules.scala 143:103:@17807.4]
  assign _T_71413 = $signed(_T_71412); // @[Modules.scala 143:103:@17808.4]
  assign _GEN_423 = {{1{_T_68341[4]}},_T_68341}; // @[Modules.scala 143:103:@17824.4]
  assign _T_71432 = $signed(_T_56098) + $signed(_GEN_423); // @[Modules.scala 143:103:@17824.4]
  assign _T_71433 = _T_71432[5:0]; // @[Modules.scala 143:103:@17825.4]
  assign _T_71434 = $signed(_T_71433); // @[Modules.scala 143:103:@17826.4]
  assign _T_71446 = $signed(_T_56117) + $signed(_T_59124); // @[Modules.scala 143:103:@17836.4]
  assign _T_71447 = _T_71446[5:0]; // @[Modules.scala 143:103:@17837.4]
  assign _T_71448 = $signed(_T_71447); // @[Modules.scala 143:103:@17838.4]
  assign _T_71509 = $signed(_T_65382) + $signed(_T_59185); // @[Modules.scala 143:103:@17890.4]
  assign _T_71510 = _T_71509[5:0]; // @[Modules.scala 143:103:@17891.4]
  assign _T_71511 = $signed(_T_71510); // @[Modules.scala 143:103:@17892.4]
  assign _T_71515 = $signed(-4'sh1) * $signed(io_in_728); // @[Modules.scala 144:80:@17895.4]
  assign _T_71516 = $signed(_T_56189) + $signed(_T_71515); // @[Modules.scala 143:103:@17896.4]
  assign _T_71517 = _T_71516[4:0]; // @[Modules.scala 143:103:@17897.4]
  assign _T_71518 = $signed(_T_71517); // @[Modules.scala 143:103:@17898.4]
  assign _T_71520 = $signed(-4'sh1) * $signed(io_in_729); // @[Modules.scala 143:74:@17900.4]
  assign _GEN_424 = {{1{_T_71520[4]}},_T_71520}; // @[Modules.scala 143:103:@17902.4]
  assign _T_71523 = $signed(_GEN_424) + $signed(_T_62278); // @[Modules.scala 143:103:@17902.4]
  assign _T_71524 = _T_71523[5:0]; // @[Modules.scala 143:103:@17903.4]
  assign _T_71525 = $signed(_T_71524); // @[Modules.scala 143:103:@17904.4]
  assign _T_71586 = $signed(_T_59255) + $signed(_T_68500); // @[Modules.scala 143:103:@17956.4]
  assign _T_71587 = _T_71586[5:0]; // @[Modules.scala 143:103:@17957.4]
  assign _T_71588 = $signed(_T_71587); // @[Modules.scala 143:103:@17958.4]
  assign _T_71593 = $signed(_T_68502) + $signed(_T_56245); // @[Modules.scala 143:103:@17962.4]
  assign _T_71594 = _T_71593[5:0]; // @[Modules.scala 143:103:@17963.4]
  assign _T_71595 = $signed(_T_71594); // @[Modules.scala 143:103:@17964.4]
  assign _T_71600 = $signed(_T_62350) + $signed(_T_59269); // @[Modules.scala 143:103:@17968.4]
  assign _T_71601 = _T_71600[4:0]; // @[Modules.scala 143:103:@17969.4]
  assign _T_71602 = $signed(_T_71601); // @[Modules.scala 143:103:@17970.4]
  assign _T_71607 = $signed(_T_56252) + $signed(_T_59276); // @[Modules.scala 143:103:@17974.4]
  assign _T_71608 = _T_71607[5:0]; // @[Modules.scala 143:103:@17975.4]
  assign _T_71609 = $signed(_T_71608); // @[Modules.scala 143:103:@17976.4]
  assign _T_71614 = $signed(_T_59278) + $signed(_T_56264); // @[Modules.scala 143:103:@17980.4]
  assign _T_71615 = _T_71614[5:0]; // @[Modules.scala 143:103:@17981.4]
  assign _T_71616 = $signed(_T_71615); // @[Modules.scala 143:103:@17982.4]
  assign _T_71621 = $signed(_T_56266) + $signed(_T_56271); // @[Modules.scala 143:103:@17986.4]
  assign _T_71622 = _T_71621[5:0]; // @[Modules.scala 143:103:@17987.4]
  assign _T_71623 = $signed(_T_71622); // @[Modules.scala 143:103:@17988.4]
  assign _T_71625 = $signed(4'sh1) * $signed(io_in_768); // @[Modules.scala 143:74:@17990.4]
  assign _T_71628 = $signed(_T_71625) + $signed(_T_56273); // @[Modules.scala 143:103:@17992.4]
  assign _T_71629 = _T_71628[5:0]; // @[Modules.scala 143:103:@17993.4]
  assign _T_71630 = $signed(_T_71629); // @[Modules.scala 143:103:@17994.4]
  assign _T_71649 = $signed(_T_59313) + $signed(_T_59318); // @[Modules.scala 143:103:@18010.4]
  assign _T_71650 = _T_71649[5:0]; // @[Modules.scala 143:103:@18011.4]
  assign _T_71651 = $signed(_T_71650); // @[Modules.scala 143:103:@18012.4]
  assign _GEN_425 = {{1{_T_59332[4]}},_T_59332}; // @[Modules.scala 143:103:@18022.4]
  assign _T_71663 = $signed(_T_56301) + $signed(_GEN_425); // @[Modules.scala 143:103:@18022.4]
  assign _T_71664 = _T_71663[5:0]; // @[Modules.scala 143:103:@18023.4]
  assign _T_71665 = $signed(_T_71664); // @[Modules.scala 143:103:@18024.4]
  assign buffer_5_0 = {{8{_T_69474[5]}},_T_69474}; // @[Modules.scala 112:22:@8.4]
  assign _T_71666 = $signed(buffer_5_0) + $signed(buffer_2_0); // @[Modules.scala 160:64:@18026.4]
  assign _T_71667 = _T_71666[13:0]; // @[Modules.scala 160:64:@18027.4]
  assign buffer_5_314 = $signed(_T_71667); // @[Modules.scala 160:64:@18028.4]
  assign _T_71669 = $signed(buffer_2_1) + $signed(buffer_3_2); // @[Modules.scala 160:64:@18030.4]
  assign _T_71670 = _T_71669[13:0]; // @[Modules.scala 160:64:@18031.4]
  assign buffer_5_315 = $signed(_T_71670); // @[Modules.scala 160:64:@18032.4]
  assign buffer_5_4 = {{8{_T_69502[5]}},_T_69502}; // @[Modules.scala 112:22:@8.4]
  assign _T_71672 = $signed(buffer_5_4) + $signed(buffer_1_4); // @[Modules.scala 160:64:@18034.4]
  assign _T_71673 = _T_71672[13:0]; // @[Modules.scala 160:64:@18035.4]
  assign buffer_5_316 = $signed(_T_71673); // @[Modules.scala 160:64:@18036.4]
  assign buffer_5_6 = {{9{_T_69516[4]}},_T_69516}; // @[Modules.scala 112:22:@8.4]
  assign _T_71675 = $signed(buffer_5_6) + $signed(buffer_1_6); // @[Modules.scala 160:64:@18038.4]
  assign _T_71676 = _T_71675[13:0]; // @[Modules.scala 160:64:@18039.4]
  assign buffer_5_317 = $signed(_T_71676); // @[Modules.scala 160:64:@18040.4]
  assign buffer_5_9 = {{8{_T_69537[5]}},_T_69537}; // @[Modules.scala 112:22:@8.4]
  assign _T_71678 = $signed(buffer_0_7) + $signed(buffer_5_9); // @[Modules.scala 160:64:@18042.4]
  assign _T_71679 = _T_71678[13:0]; // @[Modules.scala 160:64:@18043.4]
  assign buffer_5_318 = $signed(_T_71679); // @[Modules.scala 160:64:@18044.4]
  assign buffer_5_11 = {{8{_T_69551[5]}},_T_69551}; // @[Modules.scala 112:22:@8.4]
  assign _T_71681 = $signed(buffer_1_9) + $signed(buffer_5_11); // @[Modules.scala 160:64:@18046.4]
  assign _T_71682 = _T_71681[13:0]; // @[Modules.scala 160:64:@18047.4]
  assign buffer_5_319 = $signed(_T_71682); // @[Modules.scala 160:64:@18048.4]
  assign buffer_5_12 = {{8{_T_69558[5]}},_T_69558}; // @[Modules.scala 112:22:@8.4]
  assign _T_71684 = $signed(buffer_5_12) + $signed(buffer_0_12); // @[Modules.scala 160:64:@18050.4]
  assign _T_71685 = _T_71684[13:0]; // @[Modules.scala 160:64:@18051.4]
  assign buffer_5_320 = $signed(_T_71685); // @[Modules.scala 160:64:@18052.4]
  assign buffer_5_21 = {{8{_T_69621[5]}},_T_69621}; // @[Modules.scala 112:22:@8.4]
  assign _T_71696 = $signed(buffer_4_18) + $signed(buffer_5_21); // @[Modules.scala 160:64:@18066.4]
  assign _T_71697 = _T_71696[13:0]; // @[Modules.scala 160:64:@18067.4]
  assign buffer_5_324 = $signed(_T_71697); // @[Modules.scala 160:64:@18068.4]
  assign buffer_5_24 = {{8{_T_69642[5]}},_T_69642}; // @[Modules.scala 112:22:@8.4]
  assign _T_71702 = $signed(buffer_5_24) + $signed(buffer_0_26); // @[Modules.scala 160:64:@18074.4]
  assign _T_71703 = _T_71702[13:0]; // @[Modules.scala 160:64:@18075.4]
  assign buffer_5_326 = $signed(_T_71703); // @[Modules.scala 160:64:@18076.4]
  assign buffer_5_27 = {{9{_T_69663[4]}},_T_69663}; // @[Modules.scala 112:22:@8.4]
  assign _T_71705 = $signed(buffer_0_27) + $signed(buffer_5_27); // @[Modules.scala 160:64:@18078.4]
  assign _T_71706 = _T_71705[13:0]; // @[Modules.scala 160:64:@18079.4]
  assign buffer_5_327 = $signed(_T_71706); // @[Modules.scala 160:64:@18080.4]
  assign buffer_5_28 = {{9{_T_69670[4]}},_T_69670}; // @[Modules.scala 112:22:@8.4]
  assign _T_71708 = $signed(buffer_5_28) + $signed(buffer_1_29); // @[Modules.scala 160:64:@18082.4]
  assign _T_71709 = _T_71708[13:0]; // @[Modules.scala 160:64:@18083.4]
  assign buffer_5_328 = $signed(_T_71709); // @[Modules.scala 160:64:@18084.4]
  assign buffer_5_32 = {{9{_T_69698[4]}},_T_69698}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_33 = {{9{_T_69705[4]}},_T_69705}; // @[Modules.scala 112:22:@8.4]
  assign _T_71714 = $signed(buffer_5_32) + $signed(buffer_5_33); // @[Modules.scala 160:64:@18090.4]
  assign _T_71715 = _T_71714[13:0]; // @[Modules.scala 160:64:@18091.4]
  assign buffer_5_330 = $signed(_T_71715); // @[Modules.scala 160:64:@18092.4]
  assign buffer_5_34 = {{8{_T_69712[5]}},_T_69712}; // @[Modules.scala 112:22:@8.4]
  assign _T_71717 = $signed(buffer_5_34) + $signed(buffer_1_35); // @[Modules.scala 160:64:@18094.4]
  assign _T_71718 = _T_71717[13:0]; // @[Modules.scala 160:64:@18095.4]
  assign buffer_5_331 = $signed(_T_71718); // @[Modules.scala 160:64:@18096.4]
  assign buffer_5_36 = {{8{_T_69726[5]}},_T_69726}; // @[Modules.scala 112:22:@8.4]
  assign _T_71720 = $signed(buffer_5_36) + $signed(buffer_0_38); // @[Modules.scala 160:64:@18098.4]
  assign _T_71721 = _T_71720[13:0]; // @[Modules.scala 160:64:@18099.4]
  assign buffer_5_332 = $signed(_T_71721); // @[Modules.scala 160:64:@18100.4]
  assign _T_71723 = $signed(buffer_0_39) + $signed(buffer_0_40); // @[Modules.scala 160:64:@18102.4]
  assign _T_71724 = _T_71723[13:0]; // @[Modules.scala 160:64:@18103.4]
  assign buffer_5_333 = $signed(_T_71724); // @[Modules.scala 160:64:@18104.4]
  assign buffer_5_40 = {{8{_T_69754[5]}},_T_69754}; // @[Modules.scala 112:22:@8.4]
  assign _T_71726 = $signed(buffer_5_40) + $signed(buffer_0_42); // @[Modules.scala 160:64:@18106.4]
  assign _T_71727 = _T_71726[13:0]; // @[Modules.scala 160:64:@18107.4]
  assign buffer_5_334 = $signed(_T_71727); // @[Modules.scala 160:64:@18108.4]
  assign buffer_5_42 = {{9{_T_69768[4]}},_T_69768}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_43 = {{9{_T_69775[4]}},_T_69775}; // @[Modules.scala 112:22:@8.4]
  assign _T_71729 = $signed(buffer_5_42) + $signed(buffer_5_43); // @[Modules.scala 160:64:@18110.4]
  assign _T_71730 = _T_71729[13:0]; // @[Modules.scala 160:64:@18111.4]
  assign buffer_5_335 = $signed(_T_71730); // @[Modules.scala 160:64:@18112.4]
  assign buffer_5_44 = {{8{_T_69782[5]}},_T_69782}; // @[Modules.scala 112:22:@8.4]
  assign _T_71732 = $signed(buffer_5_44) + $signed(buffer_1_44); // @[Modules.scala 160:64:@18114.4]
  assign _T_71733 = _T_71732[13:0]; // @[Modules.scala 160:64:@18115.4]
  assign buffer_5_336 = $signed(_T_71733); // @[Modules.scala 160:64:@18116.4]
  assign buffer_5_46 = {{8{_T_69796[5]}},_T_69796}; // @[Modules.scala 112:22:@8.4]
  assign _T_71735 = $signed(buffer_5_46) + $signed(buffer_2_46); // @[Modules.scala 160:64:@18118.4]
  assign _T_71736 = _T_71735[13:0]; // @[Modules.scala 160:64:@18119.4]
  assign buffer_5_337 = $signed(_T_71736); // @[Modules.scala 160:64:@18120.4]
  assign buffer_5_50 = {{8{_T_69824[5]}},_T_69824}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_51 = {{8{_T_69831[5]}},_T_69831}; // @[Modules.scala 112:22:@8.4]
  assign _T_71741 = $signed(buffer_5_50) + $signed(buffer_5_51); // @[Modules.scala 160:64:@18126.4]
  assign _T_71742 = _T_71741[13:0]; // @[Modules.scala 160:64:@18127.4]
  assign buffer_5_339 = $signed(_T_71742); // @[Modules.scala 160:64:@18128.4]
  assign buffer_5_52 = {{8{_T_69838[5]}},_T_69838}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_53 = {{9{_T_69845[4]}},_T_69845}; // @[Modules.scala 112:22:@8.4]
  assign _T_71744 = $signed(buffer_5_52) + $signed(buffer_5_53); // @[Modules.scala 160:64:@18130.4]
  assign _T_71745 = _T_71744[13:0]; // @[Modules.scala 160:64:@18131.4]
  assign buffer_5_340 = $signed(_T_71745); // @[Modules.scala 160:64:@18132.4]
  assign buffer_5_55 = {{8{_T_69859[5]}},_T_69859}; // @[Modules.scala 112:22:@8.4]
  assign _T_71747 = $signed(buffer_1_53) + $signed(buffer_5_55); // @[Modules.scala 160:64:@18134.4]
  assign _T_71748 = _T_71747[13:0]; // @[Modules.scala 160:64:@18135.4]
  assign buffer_5_341 = $signed(_T_71748); // @[Modules.scala 160:64:@18136.4]
  assign _T_71750 = $signed(buffer_3_57) + $signed(buffer_0_55); // @[Modules.scala 160:64:@18138.4]
  assign _T_71751 = _T_71750[13:0]; // @[Modules.scala 160:64:@18139.4]
  assign buffer_5_342 = $signed(_T_71751); // @[Modules.scala 160:64:@18140.4]
  assign buffer_5_58 = {{9{_T_69880[4]}},_T_69880}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_59 = {{8{_T_69887[5]}},_T_69887}; // @[Modules.scala 112:22:@8.4]
  assign _T_71753 = $signed(buffer_5_58) + $signed(buffer_5_59); // @[Modules.scala 160:64:@18142.4]
  assign _T_71754 = _T_71753[13:0]; // @[Modules.scala 160:64:@18143.4]
  assign buffer_5_343 = $signed(_T_71754); // @[Modules.scala 160:64:@18144.4]
  assign buffer_5_60 = {{8{_T_69894[5]}},_T_69894}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_61 = {{8{_T_69901[5]}},_T_69901}; // @[Modules.scala 112:22:@8.4]
  assign _T_71756 = $signed(buffer_5_60) + $signed(buffer_5_61); // @[Modules.scala 160:64:@18146.4]
  assign _T_71757 = _T_71756[13:0]; // @[Modules.scala 160:64:@18147.4]
  assign buffer_5_344 = $signed(_T_71757); // @[Modules.scala 160:64:@18148.4]
  assign buffer_5_63 = {{8{_T_69915[5]}},_T_69915}; // @[Modules.scala 112:22:@8.4]
  assign _T_71759 = $signed(buffer_4_62) + $signed(buffer_5_63); // @[Modules.scala 160:64:@18150.4]
  assign _T_71760 = _T_71759[13:0]; // @[Modules.scala 160:64:@18151.4]
  assign buffer_5_345 = $signed(_T_71760); // @[Modules.scala 160:64:@18152.4]
  assign buffer_5_64 = {{8{_T_69922[5]}},_T_69922}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_65 = {{8{_T_69929[5]}},_T_69929}; // @[Modules.scala 112:22:@8.4]
  assign _T_71762 = $signed(buffer_5_64) + $signed(buffer_5_65); // @[Modules.scala 160:64:@18154.4]
  assign _T_71763 = _T_71762[13:0]; // @[Modules.scala 160:64:@18155.4]
  assign buffer_5_346 = $signed(_T_71763); // @[Modules.scala 160:64:@18156.4]
  assign buffer_5_66 = {{8{_T_69936[5]}},_T_69936}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_67 = {{8{_T_69943[5]}},_T_69943}; // @[Modules.scala 112:22:@8.4]
  assign _T_71765 = $signed(buffer_5_66) + $signed(buffer_5_67); // @[Modules.scala 160:64:@18158.4]
  assign _T_71766 = _T_71765[13:0]; // @[Modules.scala 160:64:@18159.4]
  assign buffer_5_347 = $signed(_T_71766); // @[Modules.scala 160:64:@18160.4]
  assign buffer_5_68 = {{9{_T_69950[4]}},_T_69950}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_69 = {{8{_T_69957[5]}},_T_69957}; // @[Modules.scala 112:22:@8.4]
  assign _T_71768 = $signed(buffer_5_68) + $signed(buffer_5_69); // @[Modules.scala 160:64:@18162.4]
  assign _T_71769 = _T_71768[13:0]; // @[Modules.scala 160:64:@18163.4]
  assign buffer_5_348 = $signed(_T_71769); // @[Modules.scala 160:64:@18164.4]
  assign buffer_5_70 = {{8{_T_69964[5]}},_T_69964}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_71 = {{8{_T_69971[5]}},_T_69971}; // @[Modules.scala 112:22:@8.4]
  assign _T_71771 = $signed(buffer_5_70) + $signed(buffer_5_71); // @[Modules.scala 160:64:@18166.4]
  assign _T_71772 = _T_71771[13:0]; // @[Modules.scala 160:64:@18167.4]
  assign buffer_5_349 = $signed(_T_71772); // @[Modules.scala 160:64:@18168.4]
  assign buffer_5_72 = {{8{_T_69978[5]}},_T_69978}; // @[Modules.scala 112:22:@8.4]
  assign _T_71774 = $signed(buffer_5_72) + $signed(buffer_1_71); // @[Modules.scala 160:64:@18170.4]
  assign _T_71775 = _T_71774[13:0]; // @[Modules.scala 160:64:@18171.4]
  assign buffer_5_350 = $signed(_T_71775); // @[Modules.scala 160:64:@18172.4]
  assign buffer_5_76 = {{8{_T_70006[5]}},_T_70006}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_77 = {{8{_T_70013[5]}},_T_70013}; // @[Modules.scala 112:22:@8.4]
  assign _T_71780 = $signed(buffer_5_76) + $signed(buffer_5_77); // @[Modules.scala 160:64:@18178.4]
  assign _T_71781 = _T_71780[13:0]; // @[Modules.scala 160:64:@18179.4]
  assign buffer_5_352 = $signed(_T_71781); // @[Modules.scala 160:64:@18180.4]
  assign _T_71783 = $signed(buffer_3_79) + $signed(buffer_3_80); // @[Modules.scala 160:64:@18182.4]
  assign _T_71784 = _T_71783[13:0]; // @[Modules.scala 160:64:@18183.4]
  assign buffer_5_353 = $signed(_T_71784); // @[Modules.scala 160:64:@18184.4]
  assign buffer_5_80 = {{8{_T_70034[5]}},_T_70034}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_81 = {{8{_T_70041[5]}},_T_70041}; // @[Modules.scala 112:22:@8.4]
  assign _T_71786 = $signed(buffer_5_80) + $signed(buffer_5_81); // @[Modules.scala 160:64:@18186.4]
  assign _T_71787 = _T_71786[13:0]; // @[Modules.scala 160:64:@18187.4]
  assign buffer_5_354 = $signed(_T_71787); // @[Modules.scala 160:64:@18188.4]
  assign buffer_5_84 = {{8{_T_70062[5]}},_T_70062}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_85 = {{8{_T_70069[5]}},_T_70069}; // @[Modules.scala 112:22:@8.4]
  assign _T_71792 = $signed(buffer_5_84) + $signed(buffer_5_85); // @[Modules.scala 160:64:@18194.4]
  assign _T_71793 = _T_71792[13:0]; // @[Modules.scala 160:64:@18195.4]
  assign buffer_5_356 = $signed(_T_71793); // @[Modules.scala 160:64:@18196.4]
  assign buffer_5_90 = {{8{_T_70104[5]}},_T_70104}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_91 = {{8{_T_70111[5]}},_T_70111}; // @[Modules.scala 112:22:@8.4]
  assign _T_71801 = $signed(buffer_5_90) + $signed(buffer_5_91); // @[Modules.scala 160:64:@18206.4]
  assign _T_71802 = _T_71801[13:0]; // @[Modules.scala 160:64:@18207.4]
  assign buffer_5_359 = $signed(_T_71802); // @[Modules.scala 160:64:@18208.4]
  assign buffer_5_92 = {{8{_T_70118[5]}},_T_70118}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_93 = {{8{_T_70125[5]}},_T_70125}; // @[Modules.scala 112:22:@8.4]
  assign _T_71804 = $signed(buffer_5_92) + $signed(buffer_5_93); // @[Modules.scala 160:64:@18210.4]
  assign _T_71805 = _T_71804[13:0]; // @[Modules.scala 160:64:@18211.4]
  assign buffer_5_360 = $signed(_T_71805); // @[Modules.scala 160:64:@18212.4]
  assign buffer_5_95 = {{8{_T_70139[5]}},_T_70139}; // @[Modules.scala 112:22:@8.4]
  assign _T_71807 = $signed(buffer_0_88) + $signed(buffer_5_95); // @[Modules.scala 160:64:@18214.4]
  assign _T_71808 = _T_71807[13:0]; // @[Modules.scala 160:64:@18215.4]
  assign buffer_5_361 = $signed(_T_71808); // @[Modules.scala 160:64:@18216.4]
  assign buffer_5_96 = {{8{_T_70146[5]}},_T_70146}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_97 = {{8{_T_70153[5]}},_T_70153}; // @[Modules.scala 112:22:@8.4]
  assign _T_71810 = $signed(buffer_5_96) + $signed(buffer_5_97); // @[Modules.scala 160:64:@18218.4]
  assign _T_71811 = _T_71810[13:0]; // @[Modules.scala 160:64:@18219.4]
  assign buffer_5_362 = $signed(_T_71811); // @[Modules.scala 160:64:@18220.4]
  assign buffer_5_98 = {{8{_T_70160[5]}},_T_70160}; // @[Modules.scala 112:22:@8.4]
  assign _T_71813 = $signed(buffer_5_98) + $signed(buffer_4_93); // @[Modules.scala 160:64:@18222.4]
  assign _T_71814 = _T_71813[13:0]; // @[Modules.scala 160:64:@18223.4]
  assign buffer_5_363 = $signed(_T_71814); // @[Modules.scala 160:64:@18224.4]
  assign buffer_5_102 = {{8{_T_70188[5]}},_T_70188}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_103 = {{8{_T_70195[5]}},_T_70195}; // @[Modules.scala 112:22:@8.4]
  assign _T_71819 = $signed(buffer_5_102) + $signed(buffer_5_103); // @[Modules.scala 160:64:@18230.4]
  assign _T_71820 = _T_71819[13:0]; // @[Modules.scala 160:64:@18231.4]
  assign buffer_5_365 = $signed(_T_71820); // @[Modules.scala 160:64:@18232.4]
  assign buffer_5_104 = {{8{_T_70202[5]}},_T_70202}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_105 = {{8{_T_70209[5]}},_T_70209}; // @[Modules.scala 112:22:@8.4]
  assign _T_71822 = $signed(buffer_5_104) + $signed(buffer_5_105); // @[Modules.scala 160:64:@18234.4]
  assign _T_71823 = _T_71822[13:0]; // @[Modules.scala 160:64:@18235.4]
  assign buffer_5_366 = $signed(_T_71823); // @[Modules.scala 160:64:@18236.4]
  assign buffer_5_106 = {{8{_T_70216[5]}},_T_70216}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_107 = {{8{_T_70223[5]}},_T_70223}; // @[Modules.scala 112:22:@8.4]
  assign _T_71825 = $signed(buffer_5_106) + $signed(buffer_5_107); // @[Modules.scala 160:64:@18238.4]
  assign _T_71826 = _T_71825[13:0]; // @[Modules.scala 160:64:@18239.4]
  assign buffer_5_367 = $signed(_T_71826); // @[Modules.scala 160:64:@18240.4]
  assign buffer_5_109 = {{8{_T_70237[5]}},_T_70237}; // @[Modules.scala 112:22:@8.4]
  assign _T_71828 = $signed(buffer_2_105) + $signed(buffer_5_109); // @[Modules.scala 160:64:@18242.4]
  assign _T_71829 = _T_71828[13:0]; // @[Modules.scala 160:64:@18243.4]
  assign buffer_5_368 = $signed(_T_71829); // @[Modules.scala 160:64:@18244.4]
  assign buffer_5_110 = {{8{_T_70244[5]}},_T_70244}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_111 = {{8{_T_70251[5]}},_T_70251}; // @[Modules.scala 112:22:@8.4]
  assign _T_71831 = $signed(buffer_5_110) + $signed(buffer_5_111); // @[Modules.scala 160:64:@18246.4]
  assign _T_71832 = _T_71831[13:0]; // @[Modules.scala 160:64:@18247.4]
  assign buffer_5_369 = $signed(_T_71832); // @[Modules.scala 160:64:@18248.4]
  assign buffer_5_112 = {{8{_T_70258[5]}},_T_70258}; // @[Modules.scala 112:22:@8.4]
  assign _T_71834 = $signed(buffer_5_112) + $signed(buffer_1_109); // @[Modules.scala 160:64:@18250.4]
  assign _T_71835 = _T_71834[13:0]; // @[Modules.scala 160:64:@18251.4]
  assign buffer_5_370 = $signed(_T_71835); // @[Modules.scala 160:64:@18252.4]
  assign buffer_5_114 = {{8{_T_70272[5]}},_T_70272}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_115 = {{8{_T_70279[5]}},_T_70279}; // @[Modules.scala 112:22:@8.4]
  assign _T_71837 = $signed(buffer_5_114) + $signed(buffer_5_115); // @[Modules.scala 160:64:@18254.4]
  assign _T_71838 = _T_71837[13:0]; // @[Modules.scala 160:64:@18255.4]
  assign buffer_5_371 = $signed(_T_71838); // @[Modules.scala 160:64:@18256.4]
  assign buffer_5_116 = {{8{_T_70286[5]}},_T_70286}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_117 = {{8{_T_70293[5]}},_T_70293}; // @[Modules.scala 112:22:@8.4]
  assign _T_71840 = $signed(buffer_5_116) + $signed(buffer_5_117); // @[Modules.scala 160:64:@18258.4]
  assign _T_71841 = _T_71840[13:0]; // @[Modules.scala 160:64:@18259.4]
  assign buffer_5_372 = $signed(_T_71841); // @[Modules.scala 160:64:@18260.4]
  assign buffer_5_121 = {{9{_T_70321[4]}},_T_70321}; // @[Modules.scala 112:22:@8.4]
  assign _T_71846 = $signed(buffer_3_121) + $signed(buffer_5_121); // @[Modules.scala 160:64:@18266.4]
  assign _T_71847 = _T_71846[13:0]; // @[Modules.scala 160:64:@18267.4]
  assign buffer_5_374 = $signed(_T_71847); // @[Modules.scala 160:64:@18268.4]
  assign buffer_5_122 = {{8{_T_70328[5]}},_T_70328}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_123 = {{8{_T_70335[5]}},_T_70335}; // @[Modules.scala 112:22:@8.4]
  assign _T_71849 = $signed(buffer_5_122) + $signed(buffer_5_123); // @[Modules.scala 160:64:@18270.4]
  assign _T_71850 = _T_71849[13:0]; // @[Modules.scala 160:64:@18271.4]
  assign buffer_5_375 = $signed(_T_71850); // @[Modules.scala 160:64:@18272.4]
  assign buffer_5_124 = {{8{_T_70342[5]}},_T_70342}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_125 = {{9{_T_70349[4]}},_T_70349}; // @[Modules.scala 112:22:@8.4]
  assign _T_71852 = $signed(buffer_5_124) + $signed(buffer_5_125); // @[Modules.scala 160:64:@18274.4]
  assign _T_71853 = _T_71852[13:0]; // @[Modules.scala 160:64:@18275.4]
  assign buffer_5_376 = $signed(_T_71853); // @[Modules.scala 160:64:@18276.4]
  assign buffer_5_126 = {{8{_T_70356[5]}},_T_70356}; // @[Modules.scala 112:22:@8.4]
  assign _T_71855 = $signed(buffer_5_126) + $signed(buffer_3_131); // @[Modules.scala 160:64:@18278.4]
  assign _T_71856 = _T_71855[13:0]; // @[Modules.scala 160:64:@18279.4]
  assign buffer_5_377 = $signed(_T_71856); // @[Modules.scala 160:64:@18280.4]
  assign buffer_5_128 = {{9{_T_70370[4]}},_T_70370}; // @[Modules.scala 112:22:@8.4]
  assign _T_71858 = $signed(buffer_5_128) + $signed(buffer_0_126); // @[Modules.scala 160:64:@18282.4]
  assign _T_71859 = _T_71858[13:0]; // @[Modules.scala 160:64:@18283.4]
  assign buffer_5_378 = $signed(_T_71859); // @[Modules.scala 160:64:@18284.4]
  assign buffer_5_130 = {{8{_T_70384[5]}},_T_70384}; // @[Modules.scala 112:22:@8.4]
  assign _T_71861 = $signed(buffer_5_130) + $signed(buffer_0_128); // @[Modules.scala 160:64:@18286.4]
  assign _T_71862 = _T_71861[13:0]; // @[Modules.scala 160:64:@18287.4]
  assign buffer_5_379 = $signed(_T_71862); // @[Modules.scala 160:64:@18288.4]
  assign buffer_5_133 = {{8{_T_70405[5]}},_T_70405}; // @[Modules.scala 112:22:@8.4]
  assign _T_71864 = $signed(buffer_0_129) + $signed(buffer_5_133); // @[Modules.scala 160:64:@18290.4]
  assign _T_71865 = _T_71864[13:0]; // @[Modules.scala 160:64:@18291.4]
  assign buffer_5_380 = $signed(_T_71865); // @[Modules.scala 160:64:@18292.4]
  assign buffer_5_134 = {{9{_T_70412[4]}},_T_70412}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_135 = {{9{_T_70419[4]}},_T_70419}; // @[Modules.scala 112:22:@8.4]
  assign _T_71867 = $signed(buffer_5_134) + $signed(buffer_5_135); // @[Modules.scala 160:64:@18294.4]
  assign _T_71868 = _T_71867[13:0]; // @[Modules.scala 160:64:@18295.4]
  assign buffer_5_381 = $signed(_T_71868); // @[Modules.scala 160:64:@18296.4]
  assign _T_71870 = $signed(buffer_4_131) + $signed(buffer_1_136); // @[Modules.scala 160:64:@18298.4]
  assign _T_71871 = _T_71870[13:0]; // @[Modules.scala 160:64:@18299.4]
  assign buffer_5_382 = $signed(_T_71871); // @[Modules.scala 160:64:@18300.4]
  assign _T_71876 = $signed(buffer_3_144) + $signed(buffer_1_139); // @[Modules.scala 160:64:@18306.4]
  assign _T_71877 = _T_71876[13:0]; // @[Modules.scala 160:64:@18307.4]
  assign buffer_5_384 = $signed(_T_71877); // @[Modules.scala 160:64:@18308.4]
  assign buffer_5_142 = {{8{_T_70468[5]}},_T_70468}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_143 = {{9{_T_70475[4]}},_T_70475}; // @[Modules.scala 112:22:@8.4]
  assign _T_71879 = $signed(buffer_5_142) + $signed(buffer_5_143); // @[Modules.scala 160:64:@18310.4]
  assign _T_71880 = _T_71879[13:0]; // @[Modules.scala 160:64:@18311.4]
  assign buffer_5_385 = $signed(_T_71880); // @[Modules.scala 160:64:@18312.4]
  assign buffer_5_144 = {{9{_T_70482[4]}},_T_70482}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_145 = {{8{_T_70489[5]}},_T_70489}; // @[Modules.scala 112:22:@8.4]
  assign _T_71882 = $signed(buffer_5_144) + $signed(buffer_5_145); // @[Modules.scala 160:64:@18314.4]
  assign _T_71883 = _T_71882[13:0]; // @[Modules.scala 160:64:@18315.4]
  assign buffer_5_386 = $signed(_T_71883); // @[Modules.scala 160:64:@18316.4]
  assign buffer_5_146 = {{8{_T_70496[5]}},_T_70496}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_147 = {{8{_T_70503[5]}},_T_70503}; // @[Modules.scala 112:22:@8.4]
  assign _T_71885 = $signed(buffer_5_146) + $signed(buffer_5_147); // @[Modules.scala 160:64:@18318.4]
  assign _T_71886 = _T_71885[13:0]; // @[Modules.scala 160:64:@18319.4]
  assign buffer_5_387 = $signed(_T_71886); // @[Modules.scala 160:64:@18320.4]
  assign buffer_5_149 = {{8{_T_70517[5]}},_T_70517}; // @[Modules.scala 112:22:@8.4]
  assign _T_71888 = $signed(buffer_3_156) + $signed(buffer_5_149); // @[Modules.scala 160:64:@18322.4]
  assign _T_71889 = _T_71888[13:0]; // @[Modules.scala 160:64:@18323.4]
  assign buffer_5_388 = $signed(_T_71889); // @[Modules.scala 160:64:@18324.4]
  assign buffer_5_150 = {{8{_T_70524[5]}},_T_70524}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_151 = {{9{_T_70531[4]}},_T_70531}; // @[Modules.scala 112:22:@8.4]
  assign _T_71891 = $signed(buffer_5_150) + $signed(buffer_5_151); // @[Modules.scala 160:64:@18326.4]
  assign _T_71892 = _T_71891[13:0]; // @[Modules.scala 160:64:@18327.4]
  assign buffer_5_389 = $signed(_T_71892); // @[Modules.scala 160:64:@18328.4]
  assign buffer_5_152 = {{9{_T_70538[4]}},_T_70538}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_153 = {{9{_T_70545[4]}},_T_70545}; // @[Modules.scala 112:22:@8.4]
  assign _T_71894 = $signed(buffer_5_152) + $signed(buffer_5_153); // @[Modules.scala 160:64:@18330.4]
  assign _T_71895 = _T_71894[13:0]; // @[Modules.scala 160:64:@18331.4]
  assign buffer_5_390 = $signed(_T_71895); // @[Modules.scala 160:64:@18332.4]
  assign buffer_5_154 = {{9{_T_70552[4]}},_T_70552}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_155 = {{9{_T_70559[4]}},_T_70559}; // @[Modules.scala 112:22:@8.4]
  assign _T_71897 = $signed(buffer_5_154) + $signed(buffer_5_155); // @[Modules.scala 160:64:@18334.4]
  assign _T_71898 = _T_71897[13:0]; // @[Modules.scala 160:64:@18335.4]
  assign buffer_5_391 = $signed(_T_71898); // @[Modules.scala 160:64:@18336.4]
  assign buffer_5_157 = {{9{_T_70573[4]}},_T_70573}; // @[Modules.scala 112:22:@8.4]
  assign _T_71900 = $signed(buffer_2_160) + $signed(buffer_5_157); // @[Modules.scala 160:64:@18338.4]
  assign _T_71901 = _T_71900[13:0]; // @[Modules.scala 160:64:@18339.4]
  assign buffer_5_392 = $signed(_T_71901); // @[Modules.scala 160:64:@18340.4]
  assign buffer_5_158 = {{8{_T_70580[5]}},_T_70580}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_159 = {{8{_T_70587[5]}},_T_70587}; // @[Modules.scala 112:22:@8.4]
  assign _T_71903 = $signed(buffer_5_158) + $signed(buffer_5_159); // @[Modules.scala 160:64:@18342.4]
  assign _T_71904 = _T_71903[13:0]; // @[Modules.scala 160:64:@18343.4]
  assign buffer_5_393 = $signed(_T_71904); // @[Modules.scala 160:64:@18344.4]
  assign buffer_5_160 = {{9{_T_70594[4]}},_T_70594}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_161 = {{9{_T_70601[4]}},_T_70601}; // @[Modules.scala 112:22:@8.4]
  assign _T_71906 = $signed(buffer_5_160) + $signed(buffer_5_161); // @[Modules.scala 160:64:@18346.4]
  assign _T_71907 = _T_71906[13:0]; // @[Modules.scala 160:64:@18347.4]
  assign buffer_5_394 = $signed(_T_71907); // @[Modules.scala 160:64:@18348.4]
  assign buffer_5_162 = {{8{_T_70608[5]}},_T_70608}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_163 = {{8{_T_70615[5]}},_T_70615}; // @[Modules.scala 112:22:@8.4]
  assign _T_71909 = $signed(buffer_5_162) + $signed(buffer_5_163); // @[Modules.scala 160:64:@18350.4]
  assign _T_71910 = _T_71909[13:0]; // @[Modules.scala 160:64:@18351.4]
  assign buffer_5_395 = $signed(_T_71910); // @[Modules.scala 160:64:@18352.4]
  assign buffer_5_164 = {{8{_T_70622[5]}},_T_70622}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_165 = {{9{_T_70629[4]}},_T_70629}; // @[Modules.scala 112:22:@8.4]
  assign _T_71912 = $signed(buffer_5_164) + $signed(buffer_5_165); // @[Modules.scala 160:64:@18354.4]
  assign _T_71913 = _T_71912[13:0]; // @[Modules.scala 160:64:@18355.4]
  assign buffer_5_396 = $signed(_T_71913); // @[Modules.scala 160:64:@18356.4]
  assign buffer_5_166 = {{9{_T_70636[4]}},_T_70636}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_167 = {{9{_T_70643[4]}},_T_70643}; // @[Modules.scala 112:22:@8.4]
  assign _T_71915 = $signed(buffer_5_166) + $signed(buffer_5_167); // @[Modules.scala 160:64:@18358.4]
  assign _T_71916 = _T_71915[13:0]; // @[Modules.scala 160:64:@18359.4]
  assign buffer_5_397 = $signed(_T_71916); // @[Modules.scala 160:64:@18360.4]
  assign buffer_5_168 = {{8{_T_70650[5]}},_T_70650}; // @[Modules.scala 112:22:@8.4]
  assign _T_71918 = $signed(buffer_5_168) + $signed(buffer_4_163); // @[Modules.scala 160:64:@18362.4]
  assign _T_71919 = _T_71918[13:0]; // @[Modules.scala 160:64:@18363.4]
  assign buffer_5_398 = $signed(_T_71919); // @[Modules.scala 160:64:@18364.4]
  assign buffer_5_170 = {{9{_T_70664[4]}},_T_70664}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_171 = {{8{_T_70671[5]}},_T_70671}; // @[Modules.scala 112:22:@8.4]
  assign _T_71921 = $signed(buffer_5_170) + $signed(buffer_5_171); // @[Modules.scala 160:64:@18366.4]
  assign _T_71922 = _T_71921[13:0]; // @[Modules.scala 160:64:@18367.4]
  assign buffer_5_399 = $signed(_T_71922); // @[Modules.scala 160:64:@18368.4]
  assign buffer_5_176 = {{8{_T_70706[5]}},_T_70706}; // @[Modules.scala 112:22:@8.4]
  assign _T_71930 = $signed(buffer_5_176) + $signed(buffer_0_175); // @[Modules.scala 160:64:@18378.4]
  assign _T_71931 = _T_71930[13:0]; // @[Modules.scala 160:64:@18379.4]
  assign buffer_5_402 = $signed(_T_71931); // @[Modules.scala 160:64:@18380.4]
  assign buffer_5_178 = {{8{_T_70720[5]}},_T_70720}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_179 = {{8{_T_70727[5]}},_T_70727}; // @[Modules.scala 112:22:@8.4]
  assign _T_71933 = $signed(buffer_5_178) + $signed(buffer_5_179); // @[Modules.scala 160:64:@18382.4]
  assign _T_71934 = _T_71933[13:0]; // @[Modules.scala 160:64:@18383.4]
  assign buffer_5_403 = $signed(_T_71934); // @[Modules.scala 160:64:@18384.4]
  assign buffer_5_180 = {{8{_T_70734[5]}},_T_70734}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_181 = {{9{_T_70741[4]}},_T_70741}; // @[Modules.scala 112:22:@8.4]
  assign _T_71936 = $signed(buffer_5_180) + $signed(buffer_5_181); // @[Modules.scala 160:64:@18386.4]
  assign _T_71937 = _T_71936[13:0]; // @[Modules.scala 160:64:@18387.4]
  assign buffer_5_404 = $signed(_T_71937); // @[Modules.scala 160:64:@18388.4]
  assign _T_71939 = $signed(buffer_1_180) + $signed(buffer_2_186); // @[Modules.scala 160:64:@18390.4]
  assign _T_71940 = _T_71939[13:0]; // @[Modules.scala 160:64:@18391.4]
  assign buffer_5_405 = $signed(_T_71940); // @[Modules.scala 160:64:@18392.4]
  assign buffer_5_184 = {{8{_T_70762[5]}},_T_70762}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_185 = {{8{_T_70769[5]}},_T_70769}; // @[Modules.scala 112:22:@8.4]
  assign _T_71942 = $signed(buffer_5_184) + $signed(buffer_5_185); // @[Modules.scala 160:64:@18394.4]
  assign _T_71943 = _T_71942[13:0]; // @[Modules.scala 160:64:@18395.4]
  assign buffer_5_406 = $signed(_T_71943); // @[Modules.scala 160:64:@18396.4]
  assign buffer_5_187 = {{8{_T_70783[5]}},_T_70783}; // @[Modules.scala 112:22:@8.4]
  assign _T_71945 = $signed(buffer_0_183) + $signed(buffer_5_187); // @[Modules.scala 160:64:@18398.4]
  assign _T_71946 = _T_71945[13:0]; // @[Modules.scala 160:64:@18399.4]
  assign buffer_5_407 = $signed(_T_71946); // @[Modules.scala 160:64:@18400.4]
  assign buffer_5_190 = {{8{_T_70804[5]}},_T_70804}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_191 = {{9{_T_70811[4]}},_T_70811}; // @[Modules.scala 112:22:@8.4]
  assign _T_71951 = $signed(buffer_5_190) + $signed(buffer_5_191); // @[Modules.scala 160:64:@18406.4]
  assign _T_71952 = _T_71951[13:0]; // @[Modules.scala 160:64:@18407.4]
  assign buffer_5_409 = $signed(_T_71952); // @[Modules.scala 160:64:@18408.4]
  assign buffer_5_192 = {{9{_T_70818[4]}},_T_70818}; // @[Modules.scala 112:22:@8.4]
  assign _T_71954 = $signed(buffer_5_192) + $signed(buffer_1_191); // @[Modules.scala 160:64:@18410.4]
  assign _T_71955 = _T_71954[13:0]; // @[Modules.scala 160:64:@18411.4]
  assign buffer_5_410 = $signed(_T_71955); // @[Modules.scala 160:64:@18412.4]
  assign buffer_5_194 = {{8{_T_70832[5]}},_T_70832}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_195 = {{8{_T_70839[5]}},_T_70839}; // @[Modules.scala 112:22:@8.4]
  assign _T_71957 = $signed(buffer_5_194) + $signed(buffer_5_195); // @[Modules.scala 160:64:@18414.4]
  assign _T_71958 = _T_71957[13:0]; // @[Modules.scala 160:64:@18415.4]
  assign buffer_5_411 = $signed(_T_71958); // @[Modules.scala 160:64:@18416.4]
  assign buffer_5_196 = {{8{_T_70846[5]}},_T_70846}; // @[Modules.scala 112:22:@8.4]
  assign _T_71960 = $signed(buffer_5_196) + $signed(buffer_1_196); // @[Modules.scala 160:64:@18418.4]
  assign _T_71961 = _T_71960[13:0]; // @[Modules.scala 160:64:@18419.4]
  assign buffer_5_412 = $signed(_T_71961); // @[Modules.scala 160:64:@18420.4]
  assign buffer_5_198 = {{8{_T_70860[5]}},_T_70860}; // @[Modules.scala 112:22:@8.4]
  assign _T_71963 = $signed(buffer_5_198) + $signed(buffer_0_196); // @[Modules.scala 160:64:@18422.4]
  assign _T_71964 = _T_71963[13:0]; // @[Modules.scala 160:64:@18423.4]
  assign buffer_5_413 = $signed(_T_71964); // @[Modules.scala 160:64:@18424.4]
  assign buffer_5_200 = {{8{_T_70874[5]}},_T_70874}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_201 = {{8{_T_70881[5]}},_T_70881}; // @[Modules.scala 112:22:@8.4]
  assign _T_71966 = $signed(buffer_5_200) + $signed(buffer_5_201); // @[Modules.scala 160:64:@18426.4]
  assign _T_71967 = _T_71966[13:0]; // @[Modules.scala 160:64:@18427.4]
  assign buffer_5_414 = $signed(_T_71967); // @[Modules.scala 160:64:@18428.4]
  assign _T_71969 = $signed(buffer_1_201) + $signed(buffer_1_202); // @[Modules.scala 160:64:@18430.4]
  assign _T_71970 = _T_71969[13:0]; // @[Modules.scala 160:64:@18431.4]
  assign buffer_5_415 = $signed(_T_71970); // @[Modules.scala 160:64:@18432.4]
  assign buffer_5_204 = {{8{_T_70902[5]}},_T_70902}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_205 = {{8{_T_70909[5]}},_T_70909}; // @[Modules.scala 112:22:@8.4]
  assign _T_71972 = $signed(buffer_5_204) + $signed(buffer_5_205); // @[Modules.scala 160:64:@18434.4]
  assign _T_71973 = _T_71972[13:0]; // @[Modules.scala 160:64:@18435.4]
  assign buffer_5_416 = $signed(_T_71973); // @[Modules.scala 160:64:@18436.4]
  assign buffer_5_206 = {{8{_T_70916[5]}},_T_70916}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_207 = {{8{_T_70923[5]}},_T_70923}; // @[Modules.scala 112:22:@8.4]
  assign _T_71975 = $signed(buffer_5_206) + $signed(buffer_5_207); // @[Modules.scala 160:64:@18438.4]
  assign _T_71976 = _T_71975[13:0]; // @[Modules.scala 160:64:@18439.4]
  assign buffer_5_417 = $signed(_T_71976); // @[Modules.scala 160:64:@18440.4]
  assign buffer_5_208 = {{8{_T_70930[5]}},_T_70930}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_209 = {{8{_T_70937[5]}},_T_70937}; // @[Modules.scala 112:22:@8.4]
  assign _T_71978 = $signed(buffer_5_208) + $signed(buffer_5_209); // @[Modules.scala 160:64:@18442.4]
  assign _T_71979 = _T_71978[13:0]; // @[Modules.scala 160:64:@18443.4]
  assign buffer_5_418 = $signed(_T_71979); // @[Modules.scala 160:64:@18444.4]
  assign _T_71981 = $signed(buffer_0_207) + $signed(buffer_0_208); // @[Modules.scala 160:64:@18446.4]
  assign _T_71982 = _T_71981[13:0]; // @[Modules.scala 160:64:@18447.4]
  assign buffer_5_419 = $signed(_T_71982); // @[Modules.scala 160:64:@18448.4]
  assign buffer_5_213 = {{8{_T_70965[5]}},_T_70965}; // @[Modules.scala 112:22:@8.4]
  assign _T_71984 = $signed(buffer_0_209) + $signed(buffer_5_213); // @[Modules.scala 160:64:@18450.4]
  assign _T_71985 = _T_71984[13:0]; // @[Modules.scala 160:64:@18451.4]
  assign buffer_5_420 = $signed(_T_71985); // @[Modules.scala 160:64:@18452.4]
  assign buffer_5_214 = {{8{_T_70972[5]}},_T_70972}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_215 = {{9{_T_70979[4]}},_T_70979}; // @[Modules.scala 112:22:@8.4]
  assign _T_71987 = $signed(buffer_5_214) + $signed(buffer_5_215); // @[Modules.scala 160:64:@18454.4]
  assign _T_71988 = _T_71987[13:0]; // @[Modules.scala 160:64:@18455.4]
  assign buffer_5_421 = $signed(_T_71988); // @[Modules.scala 160:64:@18456.4]
  assign buffer_5_216 = {{9{_T_70986[4]}},_T_70986}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_217 = {{8{_T_70993[5]}},_T_70993}; // @[Modules.scala 112:22:@8.4]
  assign _T_71990 = $signed(buffer_5_216) + $signed(buffer_5_217); // @[Modules.scala 160:64:@18458.4]
  assign _T_71991 = _T_71990[13:0]; // @[Modules.scala 160:64:@18459.4]
  assign buffer_5_422 = $signed(_T_71991); // @[Modules.scala 160:64:@18460.4]
  assign buffer_5_219 = {{8{_T_71007[5]}},_T_71007}; // @[Modules.scala 112:22:@8.4]
  assign _T_71993 = $signed(buffer_3_225) + $signed(buffer_5_219); // @[Modules.scala 160:64:@18462.4]
  assign _T_71994 = _T_71993[13:0]; // @[Modules.scala 160:64:@18463.4]
  assign buffer_5_423 = $signed(_T_71994); // @[Modules.scala 160:64:@18464.4]
  assign buffer_5_220 = {{8{_T_71014[5]}},_T_71014}; // @[Modules.scala 112:22:@8.4]
  assign _T_71996 = $signed(buffer_5_220) + $signed(buffer_0_217); // @[Modules.scala 160:64:@18466.4]
  assign _T_71997 = _T_71996[13:0]; // @[Modules.scala 160:64:@18467.4]
  assign buffer_5_424 = $signed(_T_71997); // @[Modules.scala 160:64:@18468.4]
  assign buffer_5_222 = {{9{_T_71028[4]}},_T_71028}; // @[Modules.scala 112:22:@8.4]
  assign _T_71999 = $signed(buffer_5_222) + $signed(buffer_1_219); // @[Modules.scala 160:64:@18470.4]
  assign _T_72000 = _T_71999[13:0]; // @[Modules.scala 160:64:@18471.4]
  assign buffer_5_425 = $signed(_T_72000); // @[Modules.scala 160:64:@18472.4]
  assign buffer_5_224 = {{8{_T_71042[5]}},_T_71042}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_225 = {{8{_T_71049[5]}},_T_71049}; // @[Modules.scala 112:22:@8.4]
  assign _T_72002 = $signed(buffer_5_224) + $signed(buffer_5_225); // @[Modules.scala 160:64:@18474.4]
  assign _T_72003 = _T_72002[13:0]; // @[Modules.scala 160:64:@18475.4]
  assign buffer_5_426 = $signed(_T_72003); // @[Modules.scala 160:64:@18476.4]
  assign buffer_5_227 = {{8{_T_71063[5]}},_T_71063}; // @[Modules.scala 112:22:@8.4]
  assign _T_72005 = $signed(buffer_3_232) + $signed(buffer_5_227); // @[Modules.scala 160:64:@18478.4]
  assign _T_72006 = _T_72005[13:0]; // @[Modules.scala 160:64:@18479.4]
  assign buffer_5_427 = $signed(_T_72006); // @[Modules.scala 160:64:@18480.4]
  assign buffer_5_228 = {{9{_T_71070[4]}},_T_71070}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_229 = {{9{_T_71077[4]}},_T_71077}; // @[Modules.scala 112:22:@8.4]
  assign _T_72008 = $signed(buffer_5_228) + $signed(buffer_5_229); // @[Modules.scala 160:64:@18482.4]
  assign _T_72009 = _T_72008[13:0]; // @[Modules.scala 160:64:@18483.4]
  assign buffer_5_428 = $signed(_T_72009); // @[Modules.scala 160:64:@18484.4]
  assign buffer_5_230 = {{8{_T_71084[5]}},_T_71084}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_231 = {{8{_T_71091[5]}},_T_71091}; // @[Modules.scala 112:22:@8.4]
  assign _T_72011 = $signed(buffer_5_230) + $signed(buffer_5_231); // @[Modules.scala 160:64:@18486.4]
  assign _T_72012 = _T_72011[13:0]; // @[Modules.scala 160:64:@18487.4]
  assign buffer_5_429 = $signed(_T_72012); // @[Modules.scala 160:64:@18488.4]
  assign buffer_5_232 = {{8{_T_71098[5]}},_T_71098}; // @[Modules.scala 112:22:@8.4]
  assign _T_72014 = $signed(buffer_5_232) + $signed(buffer_0_226); // @[Modules.scala 160:64:@18490.4]
  assign _T_72015 = _T_72014[13:0]; // @[Modules.scala 160:64:@18491.4]
  assign buffer_5_430 = $signed(_T_72015); // @[Modules.scala 160:64:@18492.4]
  assign buffer_5_235 = {{8{_T_71119[5]}},_T_71119}; // @[Modules.scala 112:22:@8.4]
  assign _T_72017 = $signed(buffer_2_233) + $signed(buffer_5_235); // @[Modules.scala 160:64:@18494.4]
  assign _T_72018 = _T_72017[13:0]; // @[Modules.scala 160:64:@18495.4]
  assign buffer_5_431 = $signed(_T_72018); // @[Modules.scala 160:64:@18496.4]
  assign buffer_5_236 = {{8{_T_71126[5]}},_T_71126}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_237 = {{8{_T_71133[5]}},_T_71133}; // @[Modules.scala 112:22:@8.4]
  assign _T_72020 = $signed(buffer_5_236) + $signed(buffer_5_237); // @[Modules.scala 160:64:@18498.4]
  assign _T_72021 = _T_72020[13:0]; // @[Modules.scala 160:64:@18499.4]
  assign buffer_5_432 = $signed(_T_72021); // @[Modules.scala 160:64:@18500.4]
  assign buffer_5_238 = {{8{_T_71140[5]}},_T_71140}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_239 = {{8{_T_71147[5]}},_T_71147}; // @[Modules.scala 112:22:@8.4]
  assign _T_72023 = $signed(buffer_5_238) + $signed(buffer_5_239); // @[Modules.scala 160:64:@18502.4]
  assign _T_72024 = _T_72023[13:0]; // @[Modules.scala 160:64:@18503.4]
  assign buffer_5_433 = $signed(_T_72024); // @[Modules.scala 160:64:@18504.4]
  assign buffer_5_240 = {{9{_T_71154[4]}},_T_71154}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_241 = {{9{_T_71161[4]}},_T_71161}; // @[Modules.scala 112:22:@8.4]
  assign _T_72026 = $signed(buffer_5_240) + $signed(buffer_5_241); // @[Modules.scala 160:64:@18506.4]
  assign _T_72027 = _T_72026[13:0]; // @[Modules.scala 160:64:@18507.4]
  assign buffer_5_434 = $signed(_T_72027); // @[Modules.scala 160:64:@18508.4]
  assign buffer_5_242 = {{9{_T_71168[4]}},_T_71168}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_243 = {{9{_T_71175[4]}},_T_71175}; // @[Modules.scala 112:22:@8.4]
  assign _T_72029 = $signed(buffer_5_242) + $signed(buffer_5_243); // @[Modules.scala 160:64:@18510.4]
  assign _T_72030 = _T_72029[13:0]; // @[Modules.scala 160:64:@18511.4]
  assign buffer_5_435 = $signed(_T_72030); // @[Modules.scala 160:64:@18512.4]
  assign buffer_5_244 = {{8{_T_71182[5]}},_T_71182}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_245 = {{8{_T_71189[5]}},_T_71189}; // @[Modules.scala 112:22:@8.4]
  assign _T_72032 = $signed(buffer_5_244) + $signed(buffer_5_245); // @[Modules.scala 160:64:@18514.4]
  assign _T_72033 = _T_72032[13:0]; // @[Modules.scala 160:64:@18515.4]
  assign buffer_5_436 = $signed(_T_72033); // @[Modules.scala 160:64:@18516.4]
  assign buffer_5_246 = {{8{_T_71196[5]}},_T_71196}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_247 = {{9{_T_71203[4]}},_T_71203}; // @[Modules.scala 112:22:@8.4]
  assign _T_72035 = $signed(buffer_5_246) + $signed(buffer_5_247); // @[Modules.scala 160:64:@18518.4]
  assign _T_72036 = _T_72035[13:0]; // @[Modules.scala 160:64:@18519.4]
  assign buffer_5_437 = $signed(_T_72036); // @[Modules.scala 160:64:@18520.4]
  assign buffer_5_248 = {{8{_T_71210[5]}},_T_71210}; // @[Modules.scala 112:22:@8.4]
  assign _T_72038 = $signed(buffer_5_248) + $signed(buffer_0_239); // @[Modules.scala 160:64:@18522.4]
  assign _T_72039 = _T_72038[13:0]; // @[Modules.scala 160:64:@18523.4]
  assign buffer_5_438 = $signed(_T_72039); // @[Modules.scala 160:64:@18524.4]
  assign buffer_5_250 = {{8{_T_71224[5]}},_T_71224}; // @[Modules.scala 112:22:@8.4]
  assign _T_72041 = $signed(buffer_5_250) + $signed(buffer_1_243); // @[Modules.scala 160:64:@18526.4]
  assign _T_72042 = _T_72041[13:0]; // @[Modules.scala 160:64:@18527.4]
  assign buffer_5_439 = $signed(_T_72042); // @[Modules.scala 160:64:@18528.4]
  assign buffer_5_252 = {{8{_T_71238[5]}},_T_71238}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_253 = {{8{_T_71245[5]}},_T_71245}; // @[Modules.scala 112:22:@8.4]
  assign _T_72044 = $signed(buffer_5_252) + $signed(buffer_5_253); // @[Modules.scala 160:64:@18530.4]
  assign _T_72045 = _T_72044[13:0]; // @[Modules.scala 160:64:@18531.4]
  assign buffer_5_440 = $signed(_T_72045); // @[Modules.scala 160:64:@18532.4]
  assign buffer_5_254 = {{8{_T_71252[5]}},_T_71252}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_255 = {{8{_T_71259[5]}},_T_71259}; // @[Modules.scala 112:22:@8.4]
  assign _T_72047 = $signed(buffer_5_254) + $signed(buffer_5_255); // @[Modules.scala 160:64:@18534.4]
  assign _T_72048 = _T_72047[13:0]; // @[Modules.scala 160:64:@18535.4]
  assign buffer_5_441 = $signed(_T_72048); // @[Modules.scala 160:64:@18536.4]
  assign buffer_5_256 = {{8{_T_71266[5]}},_T_71266}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_257 = {{8{_T_71273[5]}},_T_71273}; // @[Modules.scala 112:22:@8.4]
  assign _T_72050 = $signed(buffer_5_256) + $signed(buffer_5_257); // @[Modules.scala 160:64:@18538.4]
  assign _T_72051 = _T_72050[13:0]; // @[Modules.scala 160:64:@18539.4]
  assign buffer_5_442 = $signed(_T_72051); // @[Modules.scala 160:64:@18540.4]
  assign buffer_5_258 = {{9{_T_71280[4]}},_T_71280}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_259 = {{8{_T_71287[5]}},_T_71287}; // @[Modules.scala 112:22:@8.4]
  assign _T_72053 = $signed(buffer_5_258) + $signed(buffer_5_259); // @[Modules.scala 160:64:@18542.4]
  assign _T_72054 = _T_72053[13:0]; // @[Modules.scala 160:64:@18543.4]
  assign buffer_5_443 = $signed(_T_72054); // @[Modules.scala 160:64:@18544.4]
  assign buffer_5_261 = {{9{_T_71301[4]}},_T_71301}; // @[Modules.scala 112:22:@8.4]
  assign _T_72056 = $signed(buffer_4_247) + $signed(buffer_5_261); // @[Modules.scala 160:64:@18546.4]
  assign _T_72057 = _T_72056[13:0]; // @[Modules.scala 160:64:@18547.4]
  assign buffer_5_444 = $signed(_T_72057); // @[Modules.scala 160:64:@18548.4]
  assign buffer_5_262 = {{8{_T_71308[5]}},_T_71308}; // @[Modules.scala 112:22:@8.4]
  assign _T_72059 = $signed(buffer_5_262) + $signed(buffer_3_263); // @[Modules.scala 160:64:@18550.4]
  assign _T_72060 = _T_72059[13:0]; // @[Modules.scala 160:64:@18551.4]
  assign buffer_5_445 = $signed(_T_72060); // @[Modules.scala 160:64:@18552.4]
  assign buffer_5_264 = {{8{_T_71322[5]}},_T_71322}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_265 = {{8{_T_71329[5]}},_T_71329}; // @[Modules.scala 112:22:@8.4]
  assign _T_72062 = $signed(buffer_5_264) + $signed(buffer_5_265); // @[Modules.scala 160:64:@18554.4]
  assign _T_72063 = _T_72062[13:0]; // @[Modules.scala 160:64:@18555.4]
  assign buffer_5_446 = $signed(_T_72063); // @[Modules.scala 160:64:@18556.4]
  assign buffer_5_266 = {{8{_T_71336[5]}},_T_71336}; // @[Modules.scala 112:22:@8.4]
  assign _T_72065 = $signed(buffer_5_266) + $signed(buffer_4_253); // @[Modules.scala 160:64:@18558.4]
  assign _T_72066 = _T_72065[13:0]; // @[Modules.scala 160:64:@18559.4]
  assign buffer_5_447 = $signed(_T_72066); // @[Modules.scala 160:64:@18560.4]
  assign buffer_5_268 = {{9{_T_71350[4]}},_T_71350}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_269 = {{9{_T_71357[4]}},_T_71357}; // @[Modules.scala 112:22:@8.4]
  assign _T_72068 = $signed(buffer_5_268) + $signed(buffer_5_269); // @[Modules.scala 160:64:@18562.4]
  assign _T_72069 = _T_72068[13:0]; // @[Modules.scala 160:64:@18563.4]
  assign buffer_5_448 = $signed(_T_72069); // @[Modules.scala 160:64:@18564.4]
  assign buffer_5_270 = {{8{_T_71364[5]}},_T_71364}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_271 = {{8{_T_71371[5]}},_T_71371}; // @[Modules.scala 112:22:@8.4]
  assign _T_72071 = $signed(buffer_5_270) + $signed(buffer_5_271); // @[Modules.scala 160:64:@18566.4]
  assign _T_72072 = _T_72071[13:0]; // @[Modules.scala 160:64:@18567.4]
  assign buffer_5_449 = $signed(_T_72072); // @[Modules.scala 160:64:@18568.4]
  assign buffer_5_273 = {{8{_T_71385[5]}},_T_71385}; // @[Modules.scala 112:22:@8.4]
  assign _T_72074 = $signed(buffer_1_263) + $signed(buffer_5_273); // @[Modules.scala 160:64:@18570.4]
  assign _T_72075 = _T_72074[13:0]; // @[Modules.scala 160:64:@18571.4]
  assign buffer_5_450 = $signed(_T_72075); // @[Modules.scala 160:64:@18572.4]
  assign buffer_5_274 = {{8{_T_71392[5]}},_T_71392}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_275 = {{8{_T_71399[5]}},_T_71399}; // @[Modules.scala 112:22:@8.4]
  assign _T_72077 = $signed(buffer_5_274) + $signed(buffer_5_275); // @[Modules.scala 160:64:@18574.4]
  assign _T_72078 = _T_72077[13:0]; // @[Modules.scala 160:64:@18575.4]
  assign buffer_5_451 = $signed(_T_72078); // @[Modules.scala 160:64:@18576.4]
  assign buffer_5_276 = {{8{_T_71406[5]}},_T_71406}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_277 = {{8{_T_71413[5]}},_T_71413}; // @[Modules.scala 112:22:@8.4]
  assign _T_72080 = $signed(buffer_5_276) + $signed(buffer_5_277); // @[Modules.scala 160:64:@18578.4]
  assign _T_72081 = _T_72080[13:0]; // @[Modules.scala 160:64:@18579.4]
  assign buffer_5_452 = $signed(_T_72081); // @[Modules.scala 160:64:@18580.4]
  assign buffer_5_280 = {{8{_T_71434[5]}},_T_71434}; // @[Modules.scala 112:22:@8.4]
  assign _T_72086 = $signed(buffer_5_280) + $signed(buffer_4_267); // @[Modules.scala 160:64:@18586.4]
  assign _T_72087 = _T_72086[13:0]; // @[Modules.scala 160:64:@18587.4]
  assign buffer_5_454 = $signed(_T_72087); // @[Modules.scala 160:64:@18588.4]
  assign buffer_5_282 = {{8{_T_71448[5]}},_T_71448}; // @[Modules.scala 112:22:@8.4]
  assign _T_72089 = $signed(buffer_5_282) + $signed(buffer_1_274); // @[Modules.scala 160:64:@18590.4]
  assign _T_72090 = _T_72089[13:0]; // @[Modules.scala 160:64:@18591.4]
  assign buffer_5_455 = $signed(_T_72090); // @[Modules.scala 160:64:@18592.4]
  assign buffer_5_291 = {{8{_T_71511[5]}},_T_71511}; // @[Modules.scala 112:22:@8.4]
  assign _T_72101 = $signed(buffer_1_281) + $signed(buffer_5_291); // @[Modules.scala 160:64:@18606.4]
  assign _T_72102 = _T_72101[13:0]; // @[Modules.scala 160:64:@18607.4]
  assign buffer_5_459 = $signed(_T_72102); // @[Modules.scala 160:64:@18608.4]
  assign buffer_5_292 = {{9{_T_71518[4]}},_T_71518}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_293 = {{8{_T_71525[5]}},_T_71525}; // @[Modules.scala 112:22:@8.4]
  assign _T_72104 = $signed(buffer_5_292) + $signed(buffer_5_293); // @[Modules.scala 160:64:@18610.4]
  assign _T_72105 = _T_72104[13:0]; // @[Modules.scala 160:64:@18611.4]
  assign buffer_5_460 = $signed(_T_72105); // @[Modules.scala 160:64:@18612.4]
  assign _T_72110 = $signed(buffer_4_282) + $signed(buffer_0_287); // @[Modules.scala 160:64:@18618.4]
  assign _T_72111 = _T_72110[13:0]; // @[Modules.scala 160:64:@18619.4]
  assign buffer_5_462 = $signed(_T_72111); // @[Modules.scala 160:64:@18620.4]
  assign buffer_5_302 = {{8{_T_71588[5]}},_T_71588}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_303 = {{8{_T_71595[5]}},_T_71595}; // @[Modules.scala 112:22:@8.4]
  assign _T_72119 = $signed(buffer_5_302) + $signed(buffer_5_303); // @[Modules.scala 160:64:@18630.4]
  assign _T_72120 = _T_72119[13:0]; // @[Modules.scala 160:64:@18631.4]
  assign buffer_5_465 = $signed(_T_72120); // @[Modules.scala 160:64:@18632.4]
  assign buffer_5_304 = {{9{_T_71602[4]}},_T_71602}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_305 = {{8{_T_71609[5]}},_T_71609}; // @[Modules.scala 112:22:@8.4]
  assign _T_72122 = $signed(buffer_5_304) + $signed(buffer_5_305); // @[Modules.scala 160:64:@18634.4]
  assign _T_72123 = _T_72122[13:0]; // @[Modules.scala 160:64:@18635.4]
  assign buffer_5_466 = $signed(_T_72123); // @[Modules.scala 160:64:@18636.4]
  assign buffer_5_306 = {{8{_T_71616[5]}},_T_71616}; // @[Modules.scala 112:22:@8.4]
  assign buffer_5_307 = {{8{_T_71623[5]}},_T_71623}; // @[Modules.scala 112:22:@8.4]
  assign _T_72125 = $signed(buffer_5_306) + $signed(buffer_5_307); // @[Modules.scala 160:64:@18638.4]
  assign _T_72126 = _T_72125[13:0]; // @[Modules.scala 160:64:@18639.4]
  assign buffer_5_467 = $signed(_T_72126); // @[Modules.scala 160:64:@18640.4]
  assign buffer_5_308 = {{8{_T_71630[5]}},_T_71630}; // @[Modules.scala 112:22:@8.4]
  assign _T_72128 = $signed(buffer_5_308) + $signed(buffer_0_297); // @[Modules.scala 160:64:@18642.4]
  assign _T_72129 = _T_72128[13:0]; // @[Modules.scala 160:64:@18643.4]
  assign buffer_5_468 = $signed(_T_72129); // @[Modules.scala 160:64:@18644.4]
  assign buffer_5_311 = {{8{_T_71651[5]}},_T_71651}; // @[Modules.scala 112:22:@8.4]
  assign _T_72131 = $signed(buffer_0_298) + $signed(buffer_5_311); // @[Modules.scala 160:64:@18646.4]
  assign _T_72132 = _T_72131[13:0]; // @[Modules.scala 160:64:@18647.4]
  assign buffer_5_469 = $signed(_T_72132); // @[Modules.scala 160:64:@18648.4]
  assign buffer_5_313 = {{8{_T_71665[5]}},_T_71665}; // @[Modules.scala 112:22:@8.4]
  assign _T_72134 = $signed(buffer_2_309) + $signed(buffer_5_313); // @[Modules.scala 160:64:@18650.4]
  assign _T_72135 = _T_72134[13:0]; // @[Modules.scala 160:64:@18651.4]
  assign buffer_5_470 = $signed(_T_72135); // @[Modules.scala 160:64:@18652.4]
  assign _T_72137 = $signed(buffer_5_314) + $signed(buffer_5_315); // @[Modules.scala 166:64:@18654.4]
  assign _T_72138 = _T_72137[13:0]; // @[Modules.scala 166:64:@18655.4]
  assign buffer_5_471 = $signed(_T_72138); // @[Modules.scala 166:64:@18656.4]
  assign _T_72140 = $signed(buffer_5_316) + $signed(buffer_5_317); // @[Modules.scala 166:64:@18658.4]
  assign _T_72141 = _T_72140[13:0]; // @[Modules.scala 166:64:@18659.4]
  assign buffer_5_472 = $signed(_T_72141); // @[Modules.scala 166:64:@18660.4]
  assign _T_72143 = $signed(buffer_5_318) + $signed(buffer_5_319); // @[Modules.scala 166:64:@18662.4]
  assign _T_72144 = _T_72143[13:0]; // @[Modules.scala 166:64:@18663.4]
  assign buffer_5_473 = $signed(_T_72144); // @[Modules.scala 166:64:@18664.4]
  assign _T_72146 = $signed(buffer_5_320) + $signed(buffer_4_306); // @[Modules.scala 166:64:@18666.4]
  assign _T_72147 = _T_72146[13:0]; // @[Modules.scala 166:64:@18667.4]
  assign buffer_5_474 = $signed(_T_72147); // @[Modules.scala 166:64:@18668.4]
  assign _T_72149 = $signed(buffer_2_317) + $signed(buffer_3_322); // @[Modules.scala 166:64:@18670.4]
  assign _T_72150 = _T_72149[13:0]; // @[Modules.scala 166:64:@18671.4]
  assign buffer_5_475 = $signed(_T_72150); // @[Modules.scala 166:64:@18672.4]
  assign _T_72152 = $signed(buffer_5_324) + $signed(buffer_1_315); // @[Modules.scala 166:64:@18674.4]
  assign _T_72153 = _T_72152[13:0]; // @[Modules.scala 166:64:@18675.4]
  assign buffer_5_476 = $signed(_T_72153); // @[Modules.scala 166:64:@18676.4]
  assign _T_72155 = $signed(buffer_5_326) + $signed(buffer_5_327); // @[Modules.scala 166:64:@18678.4]
  assign _T_72156 = _T_72155[13:0]; // @[Modules.scala 166:64:@18679.4]
  assign buffer_5_477 = $signed(_T_72156); // @[Modules.scala 166:64:@18680.4]
  assign _T_72158 = $signed(buffer_5_328) + $signed(buffer_1_319); // @[Modules.scala 166:64:@18682.4]
  assign _T_72159 = _T_72158[13:0]; // @[Modules.scala 166:64:@18683.4]
  assign buffer_5_478 = $signed(_T_72159); // @[Modules.scala 166:64:@18684.4]
  assign _T_72161 = $signed(buffer_5_330) + $signed(buffer_5_331); // @[Modules.scala 166:64:@18686.4]
  assign _T_72162 = _T_72161[13:0]; // @[Modules.scala 166:64:@18687.4]
  assign buffer_5_479 = $signed(_T_72162); // @[Modules.scala 166:64:@18688.4]
  assign _T_72164 = $signed(buffer_5_332) + $signed(buffer_5_333); // @[Modules.scala 166:64:@18690.4]
  assign _T_72165 = _T_72164[13:0]; // @[Modules.scala 166:64:@18691.4]
  assign buffer_5_480 = $signed(_T_72165); // @[Modules.scala 166:64:@18692.4]
  assign _T_72167 = $signed(buffer_5_334) + $signed(buffer_5_335); // @[Modules.scala 166:64:@18694.4]
  assign _T_72168 = _T_72167[13:0]; // @[Modules.scala 166:64:@18695.4]
  assign buffer_5_481 = $signed(_T_72168); // @[Modules.scala 166:64:@18696.4]
  assign _T_72170 = $signed(buffer_5_336) + $signed(buffer_5_337); // @[Modules.scala 166:64:@18698.4]
  assign _T_72171 = _T_72170[13:0]; // @[Modules.scala 166:64:@18699.4]
  assign buffer_5_482 = $signed(_T_72171); // @[Modules.scala 166:64:@18700.4]
  assign _T_72173 = $signed(buffer_1_328) + $signed(buffer_5_339); // @[Modules.scala 166:64:@18702.4]
  assign _T_72174 = _T_72173[13:0]; // @[Modules.scala 166:64:@18703.4]
  assign buffer_5_483 = $signed(_T_72174); // @[Modules.scala 166:64:@18704.4]
  assign _T_72176 = $signed(buffer_5_340) + $signed(buffer_5_341); // @[Modules.scala 166:64:@18706.4]
  assign _T_72177 = _T_72176[13:0]; // @[Modules.scala 166:64:@18707.4]
  assign buffer_5_484 = $signed(_T_72177); // @[Modules.scala 166:64:@18708.4]
  assign _T_72179 = $signed(buffer_5_342) + $signed(buffer_5_343); // @[Modules.scala 166:64:@18710.4]
  assign _T_72180 = _T_72179[13:0]; // @[Modules.scala 166:64:@18711.4]
  assign buffer_5_485 = $signed(_T_72180); // @[Modules.scala 166:64:@18712.4]
  assign _T_72182 = $signed(buffer_5_344) + $signed(buffer_5_345); // @[Modules.scala 166:64:@18714.4]
  assign _T_72183 = _T_72182[13:0]; // @[Modules.scala 166:64:@18715.4]
  assign buffer_5_486 = $signed(_T_72183); // @[Modules.scala 166:64:@18716.4]
  assign _T_72185 = $signed(buffer_5_346) + $signed(buffer_5_347); // @[Modules.scala 166:64:@18718.4]
  assign _T_72186 = _T_72185[13:0]; // @[Modules.scala 166:64:@18719.4]
  assign buffer_5_487 = $signed(_T_72186); // @[Modules.scala 166:64:@18720.4]
  assign _T_72188 = $signed(buffer_5_348) + $signed(buffer_5_349); // @[Modules.scala 166:64:@18722.4]
  assign _T_72189 = _T_72188[13:0]; // @[Modules.scala 166:64:@18723.4]
  assign buffer_5_488 = $signed(_T_72189); // @[Modules.scala 166:64:@18724.4]
  assign _T_72191 = $signed(buffer_5_350) + $signed(buffer_1_340); // @[Modules.scala 166:64:@18726.4]
  assign _T_72192 = _T_72191[13:0]; // @[Modules.scala 166:64:@18727.4]
  assign buffer_5_489 = $signed(_T_72192); // @[Modules.scala 166:64:@18728.4]
  assign _T_72194 = $signed(buffer_5_352) + $signed(buffer_5_353); // @[Modules.scala 166:64:@18730.4]
  assign _T_72195 = _T_72194[13:0]; // @[Modules.scala 166:64:@18731.4]
  assign buffer_5_490 = $signed(_T_72195); // @[Modules.scala 166:64:@18732.4]
  assign _T_72197 = $signed(buffer_5_354) + $signed(buffer_0_341); // @[Modules.scala 166:64:@18734.4]
  assign _T_72198 = _T_72197[13:0]; // @[Modules.scala 166:64:@18735.4]
  assign buffer_5_491 = $signed(_T_72198); // @[Modules.scala 166:64:@18736.4]
  assign _T_72200 = $signed(buffer_5_356) + $signed(buffer_1_346); // @[Modules.scala 166:64:@18738.4]
  assign _T_72201 = _T_72200[13:0]; // @[Modules.scala 166:64:@18739.4]
  assign buffer_5_492 = $signed(_T_72201); // @[Modules.scala 166:64:@18740.4]
  assign _T_72203 = $signed(buffer_3_358) + $signed(buffer_5_359); // @[Modules.scala 166:64:@18742.4]
  assign _T_72204 = _T_72203[13:0]; // @[Modules.scala 166:64:@18743.4]
  assign buffer_5_493 = $signed(_T_72204); // @[Modules.scala 166:64:@18744.4]
  assign _T_72206 = $signed(buffer_5_360) + $signed(buffer_5_361); // @[Modules.scala 166:64:@18746.4]
  assign _T_72207 = _T_72206[13:0]; // @[Modules.scala 166:64:@18747.4]
  assign buffer_5_494 = $signed(_T_72207); // @[Modules.scala 166:64:@18748.4]
  assign _T_72209 = $signed(buffer_5_362) + $signed(buffer_5_363); // @[Modules.scala 166:64:@18750.4]
  assign _T_72210 = _T_72209[13:0]; // @[Modules.scala 166:64:@18751.4]
  assign buffer_5_495 = $signed(_T_72210); // @[Modules.scala 166:64:@18752.4]
  assign _T_72212 = $signed(buffer_4_347) + $signed(buffer_5_365); // @[Modules.scala 166:64:@18754.4]
  assign _T_72213 = _T_72212[13:0]; // @[Modules.scala 166:64:@18755.4]
  assign buffer_5_496 = $signed(_T_72213); // @[Modules.scala 166:64:@18756.4]
  assign _T_72215 = $signed(buffer_5_366) + $signed(buffer_5_367); // @[Modules.scala 166:64:@18758.4]
  assign _T_72216 = _T_72215[13:0]; // @[Modules.scala 166:64:@18759.4]
  assign buffer_5_497 = $signed(_T_72216); // @[Modules.scala 166:64:@18760.4]
  assign _T_72218 = $signed(buffer_5_368) + $signed(buffer_5_369); // @[Modules.scala 166:64:@18762.4]
  assign _T_72219 = _T_72218[13:0]; // @[Modules.scala 166:64:@18763.4]
  assign buffer_5_498 = $signed(_T_72219); // @[Modules.scala 166:64:@18764.4]
  assign _T_72221 = $signed(buffer_5_370) + $signed(buffer_5_371); // @[Modules.scala 166:64:@18766.4]
  assign _T_72222 = _T_72221[13:0]; // @[Modules.scala 166:64:@18767.4]
  assign buffer_5_499 = $signed(_T_72222); // @[Modules.scala 166:64:@18768.4]
  assign _T_72224 = $signed(buffer_5_372) + $signed(buffer_1_361); // @[Modules.scala 166:64:@18770.4]
  assign _T_72225 = _T_72224[13:0]; // @[Modules.scala 166:64:@18771.4]
  assign buffer_5_500 = $signed(_T_72225); // @[Modules.scala 166:64:@18772.4]
  assign _T_72227 = $signed(buffer_5_374) + $signed(buffer_5_375); // @[Modules.scala 166:64:@18774.4]
  assign _T_72228 = _T_72227[13:0]; // @[Modules.scala 166:64:@18775.4]
  assign buffer_5_501 = $signed(_T_72228); // @[Modules.scala 166:64:@18776.4]
  assign _T_72230 = $signed(buffer_5_376) + $signed(buffer_5_377); // @[Modules.scala 166:64:@18778.4]
  assign _T_72231 = _T_72230[13:0]; // @[Modules.scala 166:64:@18779.4]
  assign buffer_5_502 = $signed(_T_72231); // @[Modules.scala 166:64:@18780.4]
  assign _T_72233 = $signed(buffer_5_378) + $signed(buffer_5_379); // @[Modules.scala 166:64:@18782.4]
  assign _T_72234 = _T_72233[13:0]; // @[Modules.scala 166:64:@18783.4]
  assign buffer_5_503 = $signed(_T_72234); // @[Modules.scala 166:64:@18784.4]
  assign _T_72236 = $signed(buffer_5_380) + $signed(buffer_5_381); // @[Modules.scala 166:64:@18786.4]
  assign _T_72237 = _T_72236[13:0]; // @[Modules.scala 166:64:@18787.4]
  assign buffer_5_504 = $signed(_T_72237); // @[Modules.scala 166:64:@18788.4]
  assign _T_72239 = $signed(buffer_5_382) + $signed(buffer_3_385); // @[Modules.scala 166:64:@18790.4]
  assign _T_72240 = _T_72239[13:0]; // @[Modules.scala 166:64:@18791.4]
  assign buffer_5_505 = $signed(_T_72240); // @[Modules.scala 166:64:@18792.4]
  assign _T_72242 = $signed(buffer_5_384) + $signed(buffer_5_385); // @[Modules.scala 166:64:@18794.4]
  assign _T_72243 = _T_72242[13:0]; // @[Modules.scala 166:64:@18795.4]
  assign buffer_5_506 = $signed(_T_72243); // @[Modules.scala 166:64:@18796.4]
  assign _T_72245 = $signed(buffer_5_386) + $signed(buffer_5_387); // @[Modules.scala 166:64:@18798.4]
  assign _T_72246 = _T_72245[13:0]; // @[Modules.scala 166:64:@18799.4]
  assign buffer_5_507 = $signed(_T_72246); // @[Modules.scala 166:64:@18800.4]
  assign _T_72248 = $signed(buffer_5_388) + $signed(buffer_5_389); // @[Modules.scala 166:64:@18802.4]
  assign _T_72249 = _T_72248[13:0]; // @[Modules.scala 166:64:@18803.4]
  assign buffer_5_508 = $signed(_T_72249); // @[Modules.scala 166:64:@18804.4]
  assign _T_72251 = $signed(buffer_5_390) + $signed(buffer_5_391); // @[Modules.scala 166:64:@18806.4]
  assign _T_72252 = _T_72251[13:0]; // @[Modules.scala 166:64:@18807.4]
  assign buffer_5_509 = $signed(_T_72252); // @[Modules.scala 166:64:@18808.4]
  assign _T_72254 = $signed(buffer_5_392) + $signed(buffer_5_393); // @[Modules.scala 166:64:@18810.4]
  assign _T_72255 = _T_72254[13:0]; // @[Modules.scala 166:64:@18811.4]
  assign buffer_5_510 = $signed(_T_72255); // @[Modules.scala 166:64:@18812.4]
  assign _T_72257 = $signed(buffer_5_394) + $signed(buffer_5_395); // @[Modules.scala 166:64:@18814.4]
  assign _T_72258 = _T_72257[13:0]; // @[Modules.scala 166:64:@18815.4]
  assign buffer_5_511 = $signed(_T_72258); // @[Modules.scala 166:64:@18816.4]
  assign _T_72260 = $signed(buffer_5_396) + $signed(buffer_5_397); // @[Modules.scala 166:64:@18818.4]
  assign _T_72261 = _T_72260[13:0]; // @[Modules.scala 166:64:@18819.4]
  assign buffer_5_512 = $signed(_T_72261); // @[Modules.scala 166:64:@18820.4]
  assign _T_72263 = $signed(buffer_5_398) + $signed(buffer_5_399); // @[Modules.scala 166:64:@18822.4]
  assign _T_72264 = _T_72263[13:0]; // @[Modules.scala 166:64:@18823.4]
  assign buffer_5_513 = $signed(_T_72264); // @[Modules.scala 166:64:@18824.4]
  assign _T_72266 = $signed(buffer_3_402) + $signed(buffer_0_388); // @[Modules.scala 166:64:@18826.4]
  assign _T_72267 = _T_72266[13:0]; // @[Modules.scala 166:64:@18827.4]
  assign buffer_5_514 = $signed(_T_72267); // @[Modules.scala 166:64:@18828.4]
  assign _T_72269 = $signed(buffer_5_402) + $signed(buffer_5_403); // @[Modules.scala 166:64:@18830.4]
  assign _T_72270 = _T_72269[13:0]; // @[Modules.scala 166:64:@18831.4]
  assign buffer_5_515 = $signed(_T_72270); // @[Modules.scala 166:64:@18832.4]
  assign _T_72272 = $signed(buffer_5_404) + $signed(buffer_5_405); // @[Modules.scala 166:64:@18834.4]
  assign _T_72273 = _T_72272[13:0]; // @[Modules.scala 166:64:@18835.4]
  assign buffer_5_516 = $signed(_T_72273); // @[Modules.scala 166:64:@18836.4]
  assign _T_72275 = $signed(buffer_5_406) + $signed(buffer_5_407); // @[Modules.scala 166:64:@18838.4]
  assign _T_72276 = _T_72275[13:0]; // @[Modules.scala 166:64:@18839.4]
  assign buffer_5_517 = $signed(_T_72276); // @[Modules.scala 166:64:@18840.4]
  assign _T_72278 = $signed(buffer_0_394) + $signed(buffer_5_409); // @[Modules.scala 166:64:@18842.4]
  assign _T_72279 = _T_72278[13:0]; // @[Modules.scala 166:64:@18843.4]
  assign buffer_5_518 = $signed(_T_72279); // @[Modules.scala 166:64:@18844.4]
  assign _T_72281 = $signed(buffer_5_410) + $signed(buffer_5_411); // @[Modules.scala 166:64:@18846.4]
  assign _T_72282 = _T_72281[13:0]; // @[Modules.scala 166:64:@18847.4]
  assign buffer_5_519 = $signed(_T_72282); // @[Modules.scala 166:64:@18848.4]
  assign _T_72284 = $signed(buffer_5_412) + $signed(buffer_5_413); // @[Modules.scala 166:64:@18850.4]
  assign _T_72285 = _T_72284[13:0]; // @[Modules.scala 166:64:@18851.4]
  assign buffer_5_520 = $signed(_T_72285); // @[Modules.scala 166:64:@18852.4]
  assign _T_72287 = $signed(buffer_5_414) + $signed(buffer_5_415); // @[Modules.scala 166:64:@18854.4]
  assign _T_72288 = _T_72287[13:0]; // @[Modules.scala 166:64:@18855.4]
  assign buffer_5_521 = $signed(_T_72288); // @[Modules.scala 166:64:@18856.4]
  assign _T_72290 = $signed(buffer_5_416) + $signed(buffer_5_417); // @[Modules.scala 166:64:@18858.4]
  assign _T_72291 = _T_72290[13:0]; // @[Modules.scala 166:64:@18859.4]
  assign buffer_5_522 = $signed(_T_72291); // @[Modules.scala 166:64:@18860.4]
  assign _T_72293 = $signed(buffer_5_418) + $signed(buffer_5_419); // @[Modules.scala 166:64:@18862.4]
  assign _T_72294 = _T_72293[13:0]; // @[Modules.scala 166:64:@18863.4]
  assign buffer_5_523 = $signed(_T_72294); // @[Modules.scala 166:64:@18864.4]
  assign _T_72296 = $signed(buffer_5_420) + $signed(buffer_5_421); // @[Modules.scala 166:64:@18866.4]
  assign _T_72297 = _T_72296[13:0]; // @[Modules.scala 166:64:@18867.4]
  assign buffer_5_524 = $signed(_T_72297); // @[Modules.scala 166:64:@18868.4]
  assign _T_72299 = $signed(buffer_5_422) + $signed(buffer_5_423); // @[Modules.scala 166:64:@18870.4]
  assign _T_72300 = _T_72299[13:0]; // @[Modules.scala 166:64:@18871.4]
  assign buffer_5_525 = $signed(_T_72300); // @[Modules.scala 166:64:@18872.4]
  assign _T_72302 = $signed(buffer_5_424) + $signed(buffer_5_425); // @[Modules.scala 166:64:@18874.4]
  assign _T_72303 = _T_72302[13:0]; // @[Modules.scala 166:64:@18875.4]
  assign buffer_5_526 = $signed(_T_72303); // @[Modules.scala 166:64:@18876.4]
  assign _T_72305 = $signed(buffer_5_426) + $signed(buffer_5_427); // @[Modules.scala 166:64:@18878.4]
  assign _T_72306 = _T_72305[13:0]; // @[Modules.scala 166:64:@18879.4]
  assign buffer_5_527 = $signed(_T_72306); // @[Modules.scala 166:64:@18880.4]
  assign _T_72308 = $signed(buffer_5_428) + $signed(buffer_5_429); // @[Modules.scala 166:64:@18882.4]
  assign _T_72309 = _T_72308[13:0]; // @[Modules.scala 166:64:@18883.4]
  assign buffer_5_528 = $signed(_T_72309); // @[Modules.scala 166:64:@18884.4]
  assign _T_72311 = $signed(buffer_5_430) + $signed(buffer_5_431); // @[Modules.scala 166:64:@18886.4]
  assign _T_72312 = _T_72311[13:0]; // @[Modules.scala 166:64:@18887.4]
  assign buffer_5_529 = $signed(_T_72312); // @[Modules.scala 166:64:@18888.4]
  assign _T_72314 = $signed(buffer_5_432) + $signed(buffer_5_433); // @[Modules.scala 166:64:@18890.4]
  assign _T_72315 = _T_72314[13:0]; // @[Modules.scala 166:64:@18891.4]
  assign buffer_5_530 = $signed(_T_72315); // @[Modules.scala 166:64:@18892.4]
  assign _T_72317 = $signed(buffer_5_434) + $signed(buffer_5_435); // @[Modules.scala 166:64:@18894.4]
  assign _T_72318 = _T_72317[13:0]; // @[Modules.scala 166:64:@18895.4]
  assign buffer_5_531 = $signed(_T_72318); // @[Modules.scala 166:64:@18896.4]
  assign _T_72320 = $signed(buffer_5_436) + $signed(buffer_5_437); // @[Modules.scala 166:64:@18898.4]
  assign _T_72321 = _T_72320[13:0]; // @[Modules.scala 166:64:@18899.4]
  assign buffer_5_532 = $signed(_T_72321); // @[Modules.scala 166:64:@18900.4]
  assign _T_72323 = $signed(buffer_5_438) + $signed(buffer_5_439); // @[Modules.scala 166:64:@18902.4]
  assign _T_72324 = _T_72323[13:0]; // @[Modules.scala 166:64:@18903.4]
  assign buffer_5_533 = $signed(_T_72324); // @[Modules.scala 166:64:@18904.4]
  assign _T_72326 = $signed(buffer_5_440) + $signed(buffer_5_441); // @[Modules.scala 166:64:@18906.4]
  assign _T_72327 = _T_72326[13:0]; // @[Modules.scala 166:64:@18907.4]
  assign buffer_5_534 = $signed(_T_72327); // @[Modules.scala 166:64:@18908.4]
  assign _T_72329 = $signed(buffer_5_442) + $signed(buffer_5_443); // @[Modules.scala 166:64:@18910.4]
  assign _T_72330 = _T_72329[13:0]; // @[Modules.scala 166:64:@18911.4]
  assign buffer_5_535 = $signed(_T_72330); // @[Modules.scala 166:64:@18912.4]
  assign _T_72332 = $signed(buffer_5_444) + $signed(buffer_5_445); // @[Modules.scala 166:64:@18914.4]
  assign _T_72333 = _T_72332[13:0]; // @[Modules.scala 166:64:@18915.4]
  assign buffer_5_536 = $signed(_T_72333); // @[Modules.scala 166:64:@18916.4]
  assign _T_72335 = $signed(buffer_5_446) + $signed(buffer_5_447); // @[Modules.scala 166:64:@18918.4]
  assign _T_72336 = _T_72335[13:0]; // @[Modules.scala 166:64:@18919.4]
  assign buffer_5_537 = $signed(_T_72336); // @[Modules.scala 166:64:@18920.4]
  assign _T_72338 = $signed(buffer_5_448) + $signed(buffer_5_449); // @[Modules.scala 166:64:@18922.4]
  assign _T_72339 = _T_72338[13:0]; // @[Modules.scala 166:64:@18923.4]
  assign buffer_5_538 = $signed(_T_72339); // @[Modules.scala 166:64:@18924.4]
  assign _T_72341 = $signed(buffer_5_450) + $signed(buffer_5_451); // @[Modules.scala 166:64:@18926.4]
  assign _T_72342 = _T_72341[13:0]; // @[Modules.scala 166:64:@18927.4]
  assign buffer_5_539 = $signed(_T_72342); // @[Modules.scala 166:64:@18928.4]
  assign _T_72344 = $signed(buffer_5_452) + $signed(buffer_2_448); // @[Modules.scala 166:64:@18930.4]
  assign _T_72345 = _T_72344[13:0]; // @[Modules.scala 166:64:@18931.4]
  assign buffer_5_540 = $signed(_T_72345); // @[Modules.scala 166:64:@18932.4]
  assign _T_72347 = $signed(buffer_5_454) + $signed(buffer_5_455); // @[Modules.scala 166:64:@18934.4]
  assign _T_72348 = _T_72347[13:0]; // @[Modules.scala 166:64:@18935.4]
  assign buffer_5_541 = $signed(_T_72348); // @[Modules.scala 166:64:@18936.4]
  assign _T_72350 = $signed(buffer_4_435) + $signed(buffer_4_436); // @[Modules.scala 166:64:@18938.4]
  assign _T_72351 = _T_72350[13:0]; // @[Modules.scala 166:64:@18939.4]
  assign buffer_5_542 = $signed(_T_72351); // @[Modules.scala 166:64:@18940.4]
  assign _T_72353 = $signed(buffer_4_437) + $signed(buffer_5_459); // @[Modules.scala 166:64:@18942.4]
  assign _T_72354 = _T_72353[13:0]; // @[Modules.scala 166:64:@18943.4]
  assign buffer_5_543 = $signed(_T_72354); // @[Modules.scala 166:64:@18944.4]
  assign _T_72356 = $signed(buffer_5_460) + $signed(buffer_4_440); // @[Modules.scala 166:64:@18946.4]
  assign _T_72357 = _T_72356[13:0]; // @[Modules.scala 166:64:@18947.4]
  assign buffer_5_544 = $signed(_T_72357); // @[Modules.scala 166:64:@18948.4]
  assign _T_72359 = $signed(buffer_5_462) + $signed(buffer_1_448); // @[Modules.scala 166:64:@18950.4]
  assign _T_72360 = _T_72359[13:0]; // @[Modules.scala 166:64:@18951.4]
  assign buffer_5_545 = $signed(_T_72360); // @[Modules.scala 166:64:@18952.4]
  assign _T_72362 = $signed(buffer_1_449) + $signed(buffer_5_465); // @[Modules.scala 166:64:@18954.4]
  assign _T_72363 = _T_72362[13:0]; // @[Modules.scala 166:64:@18955.4]
  assign buffer_5_546 = $signed(_T_72363); // @[Modules.scala 166:64:@18956.4]
  assign _T_72365 = $signed(buffer_5_466) + $signed(buffer_5_467); // @[Modules.scala 166:64:@18958.4]
  assign _T_72366 = _T_72365[13:0]; // @[Modules.scala 166:64:@18959.4]
  assign buffer_5_547 = $signed(_T_72366); // @[Modules.scala 166:64:@18960.4]
  assign _T_72368 = $signed(buffer_5_468) + $signed(buffer_5_469); // @[Modules.scala 166:64:@18962.4]
  assign _T_72369 = _T_72368[13:0]; // @[Modules.scala 166:64:@18963.4]
  assign buffer_5_548 = $signed(_T_72369); // @[Modules.scala 166:64:@18964.4]
  assign _T_72371 = $signed(buffer_5_471) + $signed(buffer_5_472); // @[Modules.scala 160:64:@18966.4]
  assign _T_72372 = _T_72371[13:0]; // @[Modules.scala 160:64:@18967.4]
  assign buffer_5_549 = $signed(_T_72372); // @[Modules.scala 160:64:@18968.4]
  assign _T_72374 = $signed(buffer_5_473) + $signed(buffer_5_474); // @[Modules.scala 160:64:@18970.4]
  assign _T_72375 = _T_72374[13:0]; // @[Modules.scala 160:64:@18971.4]
  assign buffer_5_550 = $signed(_T_72375); // @[Modules.scala 160:64:@18972.4]
  assign _T_72377 = $signed(buffer_5_475) + $signed(buffer_5_476); // @[Modules.scala 160:64:@18974.4]
  assign _T_72378 = _T_72377[13:0]; // @[Modules.scala 160:64:@18975.4]
  assign buffer_5_551 = $signed(_T_72378); // @[Modules.scala 160:64:@18976.4]
  assign _T_72380 = $signed(buffer_5_477) + $signed(buffer_5_478); // @[Modules.scala 160:64:@18978.4]
  assign _T_72381 = _T_72380[13:0]; // @[Modules.scala 160:64:@18979.4]
  assign buffer_5_552 = $signed(_T_72381); // @[Modules.scala 160:64:@18980.4]
  assign _T_72383 = $signed(buffer_5_479) + $signed(buffer_5_480); // @[Modules.scala 160:64:@18982.4]
  assign _T_72384 = _T_72383[13:0]; // @[Modules.scala 160:64:@18983.4]
  assign buffer_5_553 = $signed(_T_72384); // @[Modules.scala 160:64:@18984.4]
  assign _T_72386 = $signed(buffer_5_481) + $signed(buffer_5_482); // @[Modules.scala 160:64:@18986.4]
  assign _T_72387 = _T_72386[13:0]; // @[Modules.scala 160:64:@18987.4]
  assign buffer_5_554 = $signed(_T_72387); // @[Modules.scala 160:64:@18988.4]
  assign _T_72389 = $signed(buffer_5_483) + $signed(buffer_5_484); // @[Modules.scala 160:64:@18990.4]
  assign _T_72390 = _T_72389[13:0]; // @[Modules.scala 160:64:@18991.4]
  assign buffer_5_555 = $signed(_T_72390); // @[Modules.scala 160:64:@18992.4]
  assign _T_72392 = $signed(buffer_5_485) + $signed(buffer_5_486); // @[Modules.scala 160:64:@18994.4]
  assign _T_72393 = _T_72392[13:0]; // @[Modules.scala 160:64:@18995.4]
  assign buffer_5_556 = $signed(_T_72393); // @[Modules.scala 160:64:@18996.4]
  assign _T_72395 = $signed(buffer_5_487) + $signed(buffer_5_488); // @[Modules.scala 160:64:@18998.4]
  assign _T_72396 = _T_72395[13:0]; // @[Modules.scala 160:64:@18999.4]
  assign buffer_5_557 = $signed(_T_72396); // @[Modules.scala 160:64:@19000.4]
  assign _T_72398 = $signed(buffer_5_489) + $signed(buffer_5_490); // @[Modules.scala 160:64:@19002.4]
  assign _T_72399 = _T_72398[13:0]; // @[Modules.scala 160:64:@19003.4]
  assign buffer_5_558 = $signed(_T_72399); // @[Modules.scala 160:64:@19004.4]
  assign _T_72401 = $signed(buffer_5_491) + $signed(buffer_5_492); // @[Modules.scala 160:64:@19006.4]
  assign _T_72402 = _T_72401[13:0]; // @[Modules.scala 160:64:@19007.4]
  assign buffer_5_559 = $signed(_T_72402); // @[Modules.scala 160:64:@19008.4]
  assign _T_72404 = $signed(buffer_5_493) + $signed(buffer_5_494); // @[Modules.scala 160:64:@19010.4]
  assign _T_72405 = _T_72404[13:0]; // @[Modules.scala 160:64:@19011.4]
  assign buffer_5_560 = $signed(_T_72405); // @[Modules.scala 160:64:@19012.4]
  assign _T_72407 = $signed(buffer_5_495) + $signed(buffer_5_496); // @[Modules.scala 160:64:@19014.4]
  assign _T_72408 = _T_72407[13:0]; // @[Modules.scala 160:64:@19015.4]
  assign buffer_5_561 = $signed(_T_72408); // @[Modules.scala 160:64:@19016.4]
  assign _T_72410 = $signed(buffer_5_497) + $signed(buffer_5_498); // @[Modules.scala 160:64:@19018.4]
  assign _T_72411 = _T_72410[13:0]; // @[Modules.scala 160:64:@19019.4]
  assign buffer_5_562 = $signed(_T_72411); // @[Modules.scala 160:64:@19020.4]
  assign _T_72413 = $signed(buffer_5_499) + $signed(buffer_5_500); // @[Modules.scala 160:64:@19022.4]
  assign _T_72414 = _T_72413[13:0]; // @[Modules.scala 160:64:@19023.4]
  assign buffer_5_563 = $signed(_T_72414); // @[Modules.scala 160:64:@19024.4]
  assign _T_72416 = $signed(buffer_5_501) + $signed(buffer_5_502); // @[Modules.scala 160:64:@19026.4]
  assign _T_72417 = _T_72416[13:0]; // @[Modules.scala 160:64:@19027.4]
  assign buffer_5_564 = $signed(_T_72417); // @[Modules.scala 160:64:@19028.4]
  assign _T_72419 = $signed(buffer_5_503) + $signed(buffer_5_504); // @[Modules.scala 160:64:@19030.4]
  assign _T_72420 = _T_72419[13:0]; // @[Modules.scala 160:64:@19031.4]
  assign buffer_5_565 = $signed(_T_72420); // @[Modules.scala 160:64:@19032.4]
  assign _T_72422 = $signed(buffer_5_505) + $signed(buffer_5_506); // @[Modules.scala 160:64:@19034.4]
  assign _T_72423 = _T_72422[13:0]; // @[Modules.scala 160:64:@19035.4]
  assign buffer_5_566 = $signed(_T_72423); // @[Modules.scala 160:64:@19036.4]
  assign _T_72425 = $signed(buffer_5_507) + $signed(buffer_5_508); // @[Modules.scala 160:64:@19038.4]
  assign _T_72426 = _T_72425[13:0]; // @[Modules.scala 160:64:@19039.4]
  assign buffer_5_567 = $signed(_T_72426); // @[Modules.scala 160:64:@19040.4]
  assign _T_72428 = $signed(buffer_5_509) + $signed(buffer_5_510); // @[Modules.scala 160:64:@19042.4]
  assign _T_72429 = _T_72428[13:0]; // @[Modules.scala 160:64:@19043.4]
  assign buffer_5_568 = $signed(_T_72429); // @[Modules.scala 160:64:@19044.4]
  assign _T_72431 = $signed(buffer_5_511) + $signed(buffer_5_512); // @[Modules.scala 160:64:@19046.4]
  assign _T_72432 = _T_72431[13:0]; // @[Modules.scala 160:64:@19047.4]
  assign buffer_5_569 = $signed(_T_72432); // @[Modules.scala 160:64:@19048.4]
  assign _T_72434 = $signed(buffer_5_513) + $signed(buffer_5_514); // @[Modules.scala 160:64:@19050.4]
  assign _T_72435 = _T_72434[13:0]; // @[Modules.scala 160:64:@19051.4]
  assign buffer_5_570 = $signed(_T_72435); // @[Modules.scala 160:64:@19052.4]
  assign _T_72437 = $signed(buffer_5_515) + $signed(buffer_5_516); // @[Modules.scala 160:64:@19054.4]
  assign _T_72438 = _T_72437[13:0]; // @[Modules.scala 160:64:@19055.4]
  assign buffer_5_571 = $signed(_T_72438); // @[Modules.scala 160:64:@19056.4]
  assign _T_72440 = $signed(buffer_5_517) + $signed(buffer_5_518); // @[Modules.scala 160:64:@19058.4]
  assign _T_72441 = _T_72440[13:0]; // @[Modules.scala 160:64:@19059.4]
  assign buffer_5_572 = $signed(_T_72441); // @[Modules.scala 160:64:@19060.4]
  assign _T_72443 = $signed(buffer_5_519) + $signed(buffer_5_520); // @[Modules.scala 160:64:@19062.4]
  assign _T_72444 = _T_72443[13:0]; // @[Modules.scala 160:64:@19063.4]
  assign buffer_5_573 = $signed(_T_72444); // @[Modules.scala 160:64:@19064.4]
  assign _T_72446 = $signed(buffer_5_521) + $signed(buffer_5_522); // @[Modules.scala 160:64:@19066.4]
  assign _T_72447 = _T_72446[13:0]; // @[Modules.scala 160:64:@19067.4]
  assign buffer_5_574 = $signed(_T_72447); // @[Modules.scala 160:64:@19068.4]
  assign _T_72449 = $signed(buffer_5_523) + $signed(buffer_5_524); // @[Modules.scala 160:64:@19070.4]
  assign _T_72450 = _T_72449[13:0]; // @[Modules.scala 160:64:@19071.4]
  assign buffer_5_575 = $signed(_T_72450); // @[Modules.scala 160:64:@19072.4]
  assign _T_72452 = $signed(buffer_5_525) + $signed(buffer_5_526); // @[Modules.scala 160:64:@19074.4]
  assign _T_72453 = _T_72452[13:0]; // @[Modules.scala 160:64:@19075.4]
  assign buffer_5_576 = $signed(_T_72453); // @[Modules.scala 160:64:@19076.4]
  assign _T_72455 = $signed(buffer_5_527) + $signed(buffer_5_528); // @[Modules.scala 160:64:@19078.4]
  assign _T_72456 = _T_72455[13:0]; // @[Modules.scala 160:64:@19079.4]
  assign buffer_5_577 = $signed(_T_72456); // @[Modules.scala 160:64:@19080.4]
  assign _T_72458 = $signed(buffer_5_529) + $signed(buffer_5_530); // @[Modules.scala 160:64:@19082.4]
  assign _T_72459 = _T_72458[13:0]; // @[Modules.scala 160:64:@19083.4]
  assign buffer_5_578 = $signed(_T_72459); // @[Modules.scala 160:64:@19084.4]
  assign _T_72461 = $signed(buffer_5_531) + $signed(buffer_5_532); // @[Modules.scala 160:64:@19086.4]
  assign _T_72462 = _T_72461[13:0]; // @[Modules.scala 160:64:@19087.4]
  assign buffer_5_579 = $signed(_T_72462); // @[Modules.scala 160:64:@19088.4]
  assign _T_72464 = $signed(buffer_5_533) + $signed(buffer_5_534); // @[Modules.scala 160:64:@19090.4]
  assign _T_72465 = _T_72464[13:0]; // @[Modules.scala 160:64:@19091.4]
  assign buffer_5_580 = $signed(_T_72465); // @[Modules.scala 160:64:@19092.4]
  assign _T_72467 = $signed(buffer_5_535) + $signed(buffer_5_536); // @[Modules.scala 160:64:@19094.4]
  assign _T_72468 = _T_72467[13:0]; // @[Modules.scala 160:64:@19095.4]
  assign buffer_5_581 = $signed(_T_72468); // @[Modules.scala 160:64:@19096.4]
  assign _T_72470 = $signed(buffer_5_537) + $signed(buffer_5_538); // @[Modules.scala 160:64:@19098.4]
  assign _T_72471 = _T_72470[13:0]; // @[Modules.scala 160:64:@19099.4]
  assign buffer_5_582 = $signed(_T_72471); // @[Modules.scala 160:64:@19100.4]
  assign _T_72473 = $signed(buffer_5_539) + $signed(buffer_5_540); // @[Modules.scala 160:64:@19102.4]
  assign _T_72474 = _T_72473[13:0]; // @[Modules.scala 160:64:@19103.4]
  assign buffer_5_583 = $signed(_T_72474); // @[Modules.scala 160:64:@19104.4]
  assign _T_72476 = $signed(buffer_5_541) + $signed(buffer_5_542); // @[Modules.scala 160:64:@19106.4]
  assign _T_72477 = _T_72476[13:0]; // @[Modules.scala 160:64:@19107.4]
  assign buffer_5_584 = $signed(_T_72477); // @[Modules.scala 160:64:@19108.4]
  assign _T_72479 = $signed(buffer_5_543) + $signed(buffer_5_544); // @[Modules.scala 160:64:@19110.4]
  assign _T_72480 = _T_72479[13:0]; // @[Modules.scala 160:64:@19111.4]
  assign buffer_5_585 = $signed(_T_72480); // @[Modules.scala 160:64:@19112.4]
  assign _T_72482 = $signed(buffer_5_545) + $signed(buffer_5_546); // @[Modules.scala 160:64:@19114.4]
  assign _T_72483 = _T_72482[13:0]; // @[Modules.scala 160:64:@19115.4]
  assign buffer_5_586 = $signed(_T_72483); // @[Modules.scala 160:64:@19116.4]
  assign _T_72485 = $signed(buffer_5_547) + $signed(buffer_5_548); // @[Modules.scala 160:64:@19118.4]
  assign _T_72486 = _T_72485[13:0]; // @[Modules.scala 160:64:@19119.4]
  assign buffer_5_587 = $signed(_T_72486); // @[Modules.scala 160:64:@19120.4]
  assign _T_72488 = $signed(buffer_5_549) + $signed(buffer_5_550); // @[Modules.scala 166:64:@19122.4]
  assign _T_72489 = _T_72488[13:0]; // @[Modules.scala 166:64:@19123.4]
  assign buffer_5_588 = $signed(_T_72489); // @[Modules.scala 166:64:@19124.4]
  assign _T_72491 = $signed(buffer_5_551) + $signed(buffer_5_552); // @[Modules.scala 166:64:@19126.4]
  assign _T_72492 = _T_72491[13:0]; // @[Modules.scala 166:64:@19127.4]
  assign buffer_5_589 = $signed(_T_72492); // @[Modules.scala 166:64:@19128.4]
  assign _T_72494 = $signed(buffer_5_553) + $signed(buffer_5_554); // @[Modules.scala 166:64:@19130.4]
  assign _T_72495 = _T_72494[13:0]; // @[Modules.scala 166:64:@19131.4]
  assign buffer_5_590 = $signed(_T_72495); // @[Modules.scala 166:64:@19132.4]
  assign _T_72497 = $signed(buffer_5_555) + $signed(buffer_5_556); // @[Modules.scala 166:64:@19134.4]
  assign _T_72498 = _T_72497[13:0]; // @[Modules.scala 166:64:@19135.4]
  assign buffer_5_591 = $signed(_T_72498); // @[Modules.scala 166:64:@19136.4]
  assign _T_72500 = $signed(buffer_5_557) + $signed(buffer_5_558); // @[Modules.scala 166:64:@19138.4]
  assign _T_72501 = _T_72500[13:0]; // @[Modules.scala 166:64:@19139.4]
  assign buffer_5_592 = $signed(_T_72501); // @[Modules.scala 166:64:@19140.4]
  assign _T_72503 = $signed(buffer_5_559) + $signed(buffer_5_560); // @[Modules.scala 166:64:@19142.4]
  assign _T_72504 = _T_72503[13:0]; // @[Modules.scala 166:64:@19143.4]
  assign buffer_5_593 = $signed(_T_72504); // @[Modules.scala 166:64:@19144.4]
  assign _T_72506 = $signed(buffer_5_561) + $signed(buffer_5_562); // @[Modules.scala 166:64:@19146.4]
  assign _T_72507 = _T_72506[13:0]; // @[Modules.scala 166:64:@19147.4]
  assign buffer_5_594 = $signed(_T_72507); // @[Modules.scala 166:64:@19148.4]
  assign _T_72509 = $signed(buffer_5_563) + $signed(buffer_5_564); // @[Modules.scala 166:64:@19150.4]
  assign _T_72510 = _T_72509[13:0]; // @[Modules.scala 166:64:@19151.4]
  assign buffer_5_595 = $signed(_T_72510); // @[Modules.scala 166:64:@19152.4]
  assign _T_72512 = $signed(buffer_5_565) + $signed(buffer_5_566); // @[Modules.scala 166:64:@19154.4]
  assign _T_72513 = _T_72512[13:0]; // @[Modules.scala 166:64:@19155.4]
  assign buffer_5_596 = $signed(_T_72513); // @[Modules.scala 166:64:@19156.4]
  assign _T_72515 = $signed(buffer_5_567) + $signed(buffer_5_568); // @[Modules.scala 166:64:@19158.4]
  assign _T_72516 = _T_72515[13:0]; // @[Modules.scala 166:64:@19159.4]
  assign buffer_5_597 = $signed(_T_72516); // @[Modules.scala 166:64:@19160.4]
  assign _T_72518 = $signed(buffer_5_569) + $signed(buffer_5_570); // @[Modules.scala 166:64:@19162.4]
  assign _T_72519 = _T_72518[13:0]; // @[Modules.scala 166:64:@19163.4]
  assign buffer_5_598 = $signed(_T_72519); // @[Modules.scala 166:64:@19164.4]
  assign _T_72521 = $signed(buffer_5_571) + $signed(buffer_5_572); // @[Modules.scala 166:64:@19166.4]
  assign _T_72522 = _T_72521[13:0]; // @[Modules.scala 166:64:@19167.4]
  assign buffer_5_599 = $signed(_T_72522); // @[Modules.scala 166:64:@19168.4]
  assign _T_72524 = $signed(buffer_5_573) + $signed(buffer_5_574); // @[Modules.scala 166:64:@19170.4]
  assign _T_72525 = _T_72524[13:0]; // @[Modules.scala 166:64:@19171.4]
  assign buffer_5_600 = $signed(_T_72525); // @[Modules.scala 166:64:@19172.4]
  assign _T_72527 = $signed(buffer_5_575) + $signed(buffer_5_576); // @[Modules.scala 166:64:@19174.4]
  assign _T_72528 = _T_72527[13:0]; // @[Modules.scala 166:64:@19175.4]
  assign buffer_5_601 = $signed(_T_72528); // @[Modules.scala 166:64:@19176.4]
  assign _T_72530 = $signed(buffer_5_577) + $signed(buffer_5_578); // @[Modules.scala 166:64:@19178.4]
  assign _T_72531 = _T_72530[13:0]; // @[Modules.scala 166:64:@19179.4]
  assign buffer_5_602 = $signed(_T_72531); // @[Modules.scala 166:64:@19180.4]
  assign _T_72533 = $signed(buffer_5_579) + $signed(buffer_5_580); // @[Modules.scala 166:64:@19182.4]
  assign _T_72534 = _T_72533[13:0]; // @[Modules.scala 166:64:@19183.4]
  assign buffer_5_603 = $signed(_T_72534); // @[Modules.scala 166:64:@19184.4]
  assign _T_72536 = $signed(buffer_5_581) + $signed(buffer_5_582); // @[Modules.scala 166:64:@19186.4]
  assign _T_72537 = _T_72536[13:0]; // @[Modules.scala 166:64:@19187.4]
  assign buffer_5_604 = $signed(_T_72537); // @[Modules.scala 166:64:@19188.4]
  assign _T_72539 = $signed(buffer_5_583) + $signed(buffer_5_584); // @[Modules.scala 166:64:@19190.4]
  assign _T_72540 = _T_72539[13:0]; // @[Modules.scala 166:64:@19191.4]
  assign buffer_5_605 = $signed(_T_72540); // @[Modules.scala 166:64:@19192.4]
  assign _T_72542 = $signed(buffer_5_585) + $signed(buffer_5_586); // @[Modules.scala 166:64:@19194.4]
  assign _T_72543 = _T_72542[13:0]; // @[Modules.scala 166:64:@19195.4]
  assign buffer_5_606 = $signed(_T_72543); // @[Modules.scala 166:64:@19196.4]
  assign _T_72545 = $signed(buffer_5_587) + $signed(buffer_5_470); // @[Modules.scala 172:66:@19198.4]
  assign _T_72546 = _T_72545[13:0]; // @[Modules.scala 172:66:@19199.4]
  assign buffer_5_607 = $signed(_T_72546); // @[Modules.scala 172:66:@19200.4]
  assign _T_72548 = $signed(buffer_5_588) + $signed(buffer_5_589); // @[Modules.scala 160:64:@19202.4]
  assign _T_72549 = _T_72548[13:0]; // @[Modules.scala 160:64:@19203.4]
  assign buffer_5_608 = $signed(_T_72549); // @[Modules.scala 160:64:@19204.4]
  assign _T_72551 = $signed(buffer_5_590) + $signed(buffer_5_591); // @[Modules.scala 160:64:@19206.4]
  assign _T_72552 = _T_72551[13:0]; // @[Modules.scala 160:64:@19207.4]
  assign buffer_5_609 = $signed(_T_72552); // @[Modules.scala 160:64:@19208.4]
  assign _T_72554 = $signed(buffer_5_592) + $signed(buffer_5_593); // @[Modules.scala 160:64:@19210.4]
  assign _T_72555 = _T_72554[13:0]; // @[Modules.scala 160:64:@19211.4]
  assign buffer_5_610 = $signed(_T_72555); // @[Modules.scala 160:64:@19212.4]
  assign _T_72557 = $signed(buffer_5_594) + $signed(buffer_5_595); // @[Modules.scala 160:64:@19214.4]
  assign _T_72558 = _T_72557[13:0]; // @[Modules.scala 160:64:@19215.4]
  assign buffer_5_611 = $signed(_T_72558); // @[Modules.scala 160:64:@19216.4]
  assign _T_72560 = $signed(buffer_5_596) + $signed(buffer_5_597); // @[Modules.scala 160:64:@19218.4]
  assign _T_72561 = _T_72560[13:0]; // @[Modules.scala 160:64:@19219.4]
  assign buffer_5_612 = $signed(_T_72561); // @[Modules.scala 160:64:@19220.4]
  assign _T_72563 = $signed(buffer_5_598) + $signed(buffer_5_599); // @[Modules.scala 160:64:@19222.4]
  assign _T_72564 = _T_72563[13:0]; // @[Modules.scala 160:64:@19223.4]
  assign buffer_5_613 = $signed(_T_72564); // @[Modules.scala 160:64:@19224.4]
  assign _T_72566 = $signed(buffer_5_600) + $signed(buffer_5_601); // @[Modules.scala 160:64:@19226.4]
  assign _T_72567 = _T_72566[13:0]; // @[Modules.scala 160:64:@19227.4]
  assign buffer_5_614 = $signed(_T_72567); // @[Modules.scala 160:64:@19228.4]
  assign _T_72569 = $signed(buffer_5_602) + $signed(buffer_5_603); // @[Modules.scala 160:64:@19230.4]
  assign _T_72570 = _T_72569[13:0]; // @[Modules.scala 160:64:@19231.4]
  assign buffer_5_615 = $signed(_T_72570); // @[Modules.scala 160:64:@19232.4]
  assign _T_72572 = $signed(buffer_5_604) + $signed(buffer_5_605); // @[Modules.scala 160:64:@19234.4]
  assign _T_72573 = _T_72572[13:0]; // @[Modules.scala 160:64:@19235.4]
  assign buffer_5_616 = $signed(_T_72573); // @[Modules.scala 160:64:@19236.4]
  assign _T_72575 = $signed(buffer_5_606) + $signed(buffer_5_607); // @[Modules.scala 160:64:@19238.4]
  assign _T_72576 = _T_72575[13:0]; // @[Modules.scala 160:64:@19239.4]
  assign buffer_5_617 = $signed(_T_72576); // @[Modules.scala 160:64:@19240.4]
  assign _T_72578 = $signed(buffer_5_608) + $signed(buffer_5_609); // @[Modules.scala 160:64:@19242.4]
  assign _T_72579 = _T_72578[13:0]; // @[Modules.scala 160:64:@19243.4]
  assign buffer_5_618 = $signed(_T_72579); // @[Modules.scala 160:64:@19244.4]
  assign _T_72581 = $signed(buffer_5_610) + $signed(buffer_5_611); // @[Modules.scala 160:64:@19246.4]
  assign _T_72582 = _T_72581[13:0]; // @[Modules.scala 160:64:@19247.4]
  assign buffer_5_619 = $signed(_T_72582); // @[Modules.scala 160:64:@19248.4]
  assign _T_72584 = $signed(buffer_5_612) + $signed(buffer_5_613); // @[Modules.scala 160:64:@19250.4]
  assign _T_72585 = _T_72584[13:0]; // @[Modules.scala 160:64:@19251.4]
  assign buffer_5_620 = $signed(_T_72585); // @[Modules.scala 160:64:@19252.4]
  assign _T_72587 = $signed(buffer_5_614) + $signed(buffer_5_615); // @[Modules.scala 160:64:@19254.4]
  assign _T_72588 = _T_72587[13:0]; // @[Modules.scala 160:64:@19255.4]
  assign buffer_5_621 = $signed(_T_72588); // @[Modules.scala 160:64:@19256.4]
  assign _T_72590 = $signed(buffer_5_616) + $signed(buffer_5_617); // @[Modules.scala 160:64:@19258.4]
  assign _T_72591 = _T_72590[13:0]; // @[Modules.scala 160:64:@19259.4]
  assign buffer_5_622 = $signed(_T_72591); // @[Modules.scala 160:64:@19260.4]
  assign _T_72593 = $signed(buffer_5_618) + $signed(buffer_5_619); // @[Modules.scala 166:64:@19262.4]
  assign _T_72594 = _T_72593[13:0]; // @[Modules.scala 166:64:@19263.4]
  assign buffer_5_623 = $signed(_T_72594); // @[Modules.scala 166:64:@19264.4]
  assign _T_72596 = $signed(buffer_5_620) + $signed(buffer_5_621); // @[Modules.scala 166:64:@19266.4]
  assign _T_72597 = _T_72596[13:0]; // @[Modules.scala 166:64:@19267.4]
  assign buffer_5_624 = $signed(_T_72597); // @[Modules.scala 166:64:@19268.4]
  assign _T_72599 = $signed(buffer_5_623) + $signed(buffer_5_624); // @[Modules.scala 160:64:@19270.4]
  assign _T_72600 = _T_72599[13:0]; // @[Modules.scala 160:64:@19271.4]
  assign buffer_5_625 = $signed(_T_72600); // @[Modules.scala 160:64:@19272.4]
  assign _T_72602 = $signed(buffer_5_625) + $signed(buffer_5_622); // @[Modules.scala 172:66:@19274.4]
  assign _T_72603 = _T_72602[13:0]; // @[Modules.scala 172:66:@19275.4]
  assign buffer_5_626 = $signed(_T_72603); // @[Modules.scala 172:66:@19276.4]
  assign _T_72620 = $signed(-4'sh1) * $signed(io_in_21); // @[Modules.scala 143:74:@19447.4]
  assign _GEN_426 = {{1{_T_72620[4]}},_T_72620}; // @[Modules.scala 143:103:@19449.4]
  assign _T_72623 = $signed(_GEN_426) + $signed(_T_54215); // @[Modules.scala 143:103:@19449.4]
  assign _T_72624 = _T_72623[5:0]; // @[Modules.scala 143:103:@19450.4]
  assign _T_72625 = $signed(_T_72624); // @[Modules.scala 143:103:@19451.4]
  assign _T_72630 = $signed(_T_60264) + $signed(_T_60269); // @[Modules.scala 143:103:@19455.4]
  assign _T_72631 = _T_72630[4:0]; // @[Modules.scala 143:103:@19456.4]
  assign _T_72632 = $signed(_T_72631); // @[Modules.scala 143:103:@19457.4]
  assign _T_72637 = $signed(_T_60271) + $signed(_T_57239); // @[Modules.scala 143:103:@19461.4]
  assign _T_72638 = _T_72637[4:0]; // @[Modules.scala 143:103:@19462.4]
  assign _T_72639 = $signed(_T_72638); // @[Modules.scala 143:103:@19463.4]
  assign _T_72665 = $signed(_GEN_218) + $signed(_T_54250); // @[Modules.scala 143:103:@19485.4]
  assign _T_72666 = _T_72665[5:0]; // @[Modules.scala 143:103:@19486.4]
  assign _T_72667 = $signed(_T_72666); // @[Modules.scala 143:103:@19487.4]
  assign _T_72672 = $signed(_T_54255) + $signed(_GEN_78); // @[Modules.scala 143:103:@19491.4]
  assign _T_72673 = _T_72672[5:0]; // @[Modules.scala 143:103:@19492.4]
  assign _T_72674 = $signed(_T_72673); // @[Modules.scala 143:103:@19493.4]
  assign _T_72679 = $signed(_GEN_359) + $signed(_T_54269); // @[Modules.scala 143:103:@19497.4]
  assign _T_72680 = _T_72679[5:0]; // @[Modules.scala 143:103:@19498.4]
  assign _T_72681 = $signed(_T_72680); // @[Modules.scala 143:103:@19499.4]
  assign _T_72686 = $signed(_T_54271) + $signed(_T_54276); // @[Modules.scala 143:103:@19503.4]
  assign _T_72687 = _T_72686[5:0]; // @[Modules.scala 143:103:@19504.4]
  assign _T_72688 = $signed(_T_72687); // @[Modules.scala 143:103:@19505.4]
  assign _T_72749 = $signed(_T_57339) + $signed(_T_66603); // @[Modules.scala 143:103:@19557.4]
  assign _T_72750 = _T_72749[4:0]; // @[Modules.scala 143:103:@19558.4]
  assign _T_72751 = $signed(_T_72750); // @[Modules.scala 143:103:@19559.4]
  assign _T_72756 = $signed(_T_66605) + $signed(_T_66610); // @[Modules.scala 143:103:@19563.4]
  assign _T_72757 = _T_72756[4:0]; // @[Modules.scala 143:103:@19564.4]
  assign _T_72758 = $signed(_T_72757); // @[Modules.scala 143:103:@19565.4]
  assign _GEN_431 = {{1{_T_63487[4]}},_T_63487}; // @[Modules.scala 143:103:@19569.4]
  assign _T_72763 = $signed(_GEN_431) + $signed(_T_54353); // @[Modules.scala 143:103:@19569.4]
  assign _T_72764 = _T_72763[5:0]; // @[Modules.scala 143:103:@19570.4]
  assign _T_72765 = $signed(_T_72764); // @[Modules.scala 143:103:@19571.4]
  assign _T_72784 = $signed(_GEN_364) + $signed(_T_54381); // @[Modules.scala 143:103:@19587.4]
  assign _T_72785 = _T_72784[5:0]; // @[Modules.scala 143:103:@19588.4]
  assign _T_72786 = $signed(_T_72785); // @[Modules.scala 143:103:@19589.4]
  assign _T_72791 = $signed(_T_54383) + $signed(_T_54388); // @[Modules.scala 143:103:@19593.4]
  assign _T_72792 = _T_72791[5:0]; // @[Modules.scala 143:103:@19594.4]
  assign _T_72793 = $signed(_T_72792); // @[Modules.scala 143:103:@19595.4]
  assign _GEN_433 = {{1{_T_57416[4]}},_T_57416}; // @[Modules.scala 143:103:@19611.4]
  assign _T_72812 = $signed(_T_54409) + $signed(_GEN_433); // @[Modules.scala 143:103:@19611.4]
  assign _T_72813 = _T_72812[5:0]; // @[Modules.scala 143:103:@19612.4]
  assign _T_72814 = $signed(_T_72813); // @[Modules.scala 143:103:@19613.4]
  assign _GEN_434 = {{1{_T_57421[4]}},_T_57421}; // @[Modules.scala 143:103:@19617.4]
  assign _T_72819 = $signed(_GEN_434) + $signed(_T_54423); // @[Modules.scala 143:103:@19617.4]
  assign _T_72820 = _T_72819[5:0]; // @[Modules.scala 143:103:@19618.4]
  assign _T_72821 = $signed(_T_72820); // @[Modules.scala 143:103:@19619.4]
  assign _GEN_436 = {{1{_T_60474[4]}},_T_60474}; // @[Modules.scala 143:103:@19635.4]
  assign _T_72840 = $signed(_T_57442) + $signed(_GEN_436); // @[Modules.scala 143:103:@19635.4]
  assign _T_72841 = _T_72840[5:0]; // @[Modules.scala 143:103:@19636.4]
  assign _T_72842 = $signed(_T_72841); // @[Modules.scala 143:103:@19637.4]
  assign _T_72854 = $signed(_GEN_365) + $signed(_T_57456); // @[Modules.scala 143:103:@19647.4]
  assign _T_72855 = _T_72854[5:0]; // @[Modules.scala 143:103:@19648.4]
  assign _T_72856 = $signed(_T_72855); // @[Modules.scala 143:103:@19649.4]
  assign _T_72882 = $signed(_T_54481) + $signed(_T_54486); // @[Modules.scala 143:103:@19671.4]
  assign _T_72883 = _T_72882[5:0]; // @[Modules.scala 143:103:@19672.4]
  assign _T_72884 = $signed(_T_72883); // @[Modules.scala 143:103:@19673.4]
  assign _T_72917 = $signed(_GEN_86) + $signed(_T_57526); // @[Modules.scala 143:103:@19701.4]
  assign _T_72918 = _T_72917[5:0]; // @[Modules.scala 143:103:@19702.4]
  assign _T_72919 = $signed(_T_72918); // @[Modules.scala 143:103:@19703.4]
  assign _T_72924 = $signed(_T_54521) + $signed(_T_57533); // @[Modules.scala 143:103:@19707.4]
  assign _T_72925 = _T_72924[5:0]; // @[Modules.scala 143:103:@19708.4]
  assign _T_72926 = $signed(_T_72925); // @[Modules.scala 143:103:@19709.4]
  assign _T_72931 = $signed(_T_57535) + $signed(_T_57540); // @[Modules.scala 143:103:@19713.4]
  assign _T_72932 = _T_72931[5:0]; // @[Modules.scala 143:103:@19714.4]
  assign _T_72933 = $signed(_T_72932); // @[Modules.scala 143:103:@19715.4]
  assign _T_72959 = $signed(_T_63704) + $signed(_T_69826); // @[Modules.scala 143:103:@19737.4]
  assign _T_72960 = _T_72959[5:0]; // @[Modules.scala 143:103:@19738.4]
  assign _T_72961 = $signed(_T_72960); // @[Modules.scala 143:103:@19739.4]
  assign _T_72966 = $signed(_GEN_9) + $signed(_T_63723); // @[Modules.scala 143:103:@19743.4]
  assign _T_72967 = _T_72966[5:0]; // @[Modules.scala 143:103:@19744.4]
  assign _T_72968 = $signed(_T_72967); // @[Modules.scala 143:103:@19745.4]
  assign _T_73001 = $signed(_T_54586) + $signed(_T_54591); // @[Modules.scala 143:103:@19773.4]
  assign _T_73002 = _T_73001[5:0]; // @[Modules.scala 143:103:@19774.4]
  assign _T_73003 = $signed(_T_73002); // @[Modules.scala 143:103:@19775.4]
  assign _T_73008 = $signed(_T_54593) + $signed(_T_54598); // @[Modules.scala 143:103:@19779.4]
  assign _T_73009 = _T_73008[5:0]; // @[Modules.scala 143:103:@19780.4]
  assign _T_73010 = $signed(_T_73009); // @[Modules.scala 143:103:@19781.4]
  assign _T_73015 = $signed(_T_54600) + $signed(_T_54605); // @[Modules.scala 143:103:@19785.4]
  assign _T_73016 = _T_73015[5:0]; // @[Modules.scala 143:103:@19786.4]
  assign _T_73017 = $signed(_T_73016); // @[Modules.scala 143:103:@19787.4]
  assign _T_73021 = $signed(4'sh1) * $signed(io_in_178); // @[Modules.scala 144:80:@19790.4]
  assign _T_73022 = $signed(_T_69891) + $signed(_T_73021); // @[Modules.scala 143:103:@19791.4]
  assign _T_73023 = _T_73022[5:0]; // @[Modules.scala 143:103:@19792.4]
  assign _T_73024 = $signed(_T_73023); // @[Modules.scala 143:103:@19793.4]
  assign _T_73029 = $signed(_T_57626) + $signed(_T_57633); // @[Modules.scala 143:103:@19797.4]
  assign _T_73030 = _T_73029[5:0]; // @[Modules.scala 143:103:@19798.4]
  assign _T_73031 = $signed(_T_73030); // @[Modules.scala 143:103:@19799.4]
  assign _T_73036 = $signed(_T_57638) + $signed(_T_57645); // @[Modules.scala 143:103:@19803.4]
  assign _T_73037 = _T_73036[5:0]; // @[Modules.scala 143:103:@19804.4]
  assign _T_73038 = $signed(_T_73037); // @[Modules.scala 143:103:@19805.4]
  assign _GEN_443 = {{1{_T_54633[4]}},_T_54633}; // @[Modules.scala 143:103:@19809.4]
  assign _T_73043 = $signed(_T_66925) + $signed(_GEN_443); // @[Modules.scala 143:103:@19809.4]
  assign _T_73044 = _T_73043[5:0]; // @[Modules.scala 143:103:@19810.4]
  assign _T_73045 = $signed(_T_73044); // @[Modules.scala 143:103:@19811.4]
  assign _T_73049 = $signed(4'sh1) * $signed(io_in_189); // @[Modules.scala 144:80:@19814.4]
  assign _T_73050 = $signed(_T_69924) + $signed(_T_73049); // @[Modules.scala 143:103:@19815.4]
  assign _T_73051 = _T_73050[5:0]; // @[Modules.scala 143:103:@19816.4]
  assign _T_73052 = $signed(_T_73051); // @[Modules.scala 143:103:@19817.4]
  assign _T_73071 = $signed(_GEN_93) + $signed(_T_54654); // @[Modules.scala 143:103:@19833.4]
  assign _T_73072 = _T_73071[5:0]; // @[Modules.scala 143:103:@19834.4]
  assign _T_73073 = $signed(_T_73072); // @[Modules.scala 143:103:@19835.4]
  assign _T_73078 = $signed(_T_57675) + $signed(_T_54661); // @[Modules.scala 143:103:@19839.4]
  assign _T_73079 = _T_73078[5:0]; // @[Modules.scala 143:103:@19840.4]
  assign _T_73080 = $signed(_T_73079); // @[Modules.scala 143:103:@19841.4]
  assign _T_73092 = $signed(_T_54670) + $signed(_T_54675); // @[Modules.scala 143:103:@19851.4]
  assign _T_73093 = _T_73092[5:0]; // @[Modules.scala 143:103:@19852.4]
  assign _T_73094 = $signed(_T_73093); // @[Modules.scala 143:103:@19853.4]
  assign _T_73099 = $signed(_T_54677) + $signed(_T_54682); // @[Modules.scala 143:103:@19857.4]
  assign _T_73100 = _T_73099[5:0]; // @[Modules.scala 143:103:@19858.4]
  assign _T_73101 = $signed(_T_73100); // @[Modules.scala 143:103:@19859.4]
  assign _T_73106 = $signed(_T_69968) + $signed(_T_69973); // @[Modules.scala 143:103:@19863.4]
  assign _T_73107 = _T_73106[5:0]; // @[Modules.scala 143:103:@19864.4]
  assign _T_73108 = $signed(_T_73107); // @[Modules.scala 143:103:@19865.4]
  assign _T_73120 = $signed(_T_60754) + $signed(_T_60759); // @[Modules.scala 143:103:@19875.4]
  assign _T_73121 = _T_73120[4:0]; // @[Modules.scala 143:103:@19876.4]
  assign _T_73122 = $signed(_T_73121); // @[Modules.scala 143:103:@19877.4]
  assign _T_73127 = $signed(_GEN_17) + $signed(_T_63884); // @[Modules.scala 143:103:@19881.4]
  assign _T_73128 = _T_73127[5:0]; // @[Modules.scala 143:103:@19882.4]
  assign _T_73129 = $signed(_T_73128); // @[Modules.scala 143:103:@19883.4]
  assign _GEN_446 = {{1{_T_54710[4]}},_T_54710}; // @[Modules.scala 143:103:@19887.4]
  assign _T_73134 = $signed(_T_57736) + $signed(_GEN_446); // @[Modules.scala 143:103:@19887.4]
  assign _T_73135 = _T_73134[5:0]; // @[Modules.scala 143:103:@19888.4]
  assign _T_73136 = $signed(_T_73135); // @[Modules.scala 143:103:@19889.4]
  assign _T_73141 = $signed(_T_54712) + $signed(_T_54717); // @[Modules.scala 143:103:@19893.4]
  assign _T_73142 = _T_73141[4:0]; // @[Modules.scala 143:103:@19894.4]
  assign _T_73143 = $signed(_T_73142); // @[Modules.scala 143:103:@19895.4]
  assign _T_73148 = $signed(_T_54719) + $signed(_T_57757); // @[Modules.scala 143:103:@19899.4]
  assign _T_73149 = _T_73148[4:0]; // @[Modules.scala 143:103:@19900.4]
  assign _T_73150 = $signed(_T_73149); // @[Modules.scala 143:103:@19901.4]
  assign _T_73155 = $signed(_GEN_18) + $signed(_T_54731); // @[Modules.scala 143:103:@19905.4]
  assign _T_73156 = _T_73155[5:0]; // @[Modules.scala 143:103:@19906.4]
  assign _T_73157 = $signed(_T_73156); // @[Modules.scala 143:103:@19907.4]
  assign _T_73176 = $signed(_T_54747) + $signed(_T_54752); // @[Modules.scala 143:103:@19923.4]
  assign _T_73177 = _T_73176[5:0]; // @[Modules.scala 143:103:@19924.4]
  assign _T_73178 = $signed(_T_73177); // @[Modules.scala 143:103:@19925.4]
  assign _T_73183 = $signed(_T_54754) + $signed(_GEN_19); // @[Modules.scala 143:103:@19929.4]
  assign _T_73184 = _T_73183[5:0]; // @[Modules.scala 143:103:@19930.4]
  assign _T_73185 = $signed(_T_73184); // @[Modules.scala 143:103:@19931.4]
  assign _GEN_450 = {{1{_T_54794[4]}},_T_54794}; // @[Modules.scala 143:103:@19965.4]
  assign _T_73225 = $signed(_T_70099) + $signed(_GEN_450); // @[Modules.scala 143:103:@19965.4]
  assign _T_73226 = _T_73225[5:0]; // @[Modules.scala 143:103:@19966.4]
  assign _T_73227 = $signed(_T_73226); // @[Modules.scala 143:103:@19967.4]
  assign _GEN_451 = {{1{_T_54803[4]}},_T_54803}; // @[Modules.scala 143:103:@19977.4]
  assign _T_73239 = $signed(_GEN_451) + $signed(_T_54808); // @[Modules.scala 143:103:@19977.4]
  assign _T_73240 = _T_73239[5:0]; // @[Modules.scala 143:103:@19978.4]
  assign _T_73241 = $signed(_T_73240); // @[Modules.scala 143:103:@19979.4]
  assign _GEN_452 = {{1{_T_57869[4]}},_T_57869}; // @[Modules.scala 143:103:@20001.4]
  assign _T_73267 = $signed(_T_70143) + $signed(_GEN_452); // @[Modules.scala 143:103:@20001.4]
  assign _T_73268 = _T_73267[5:0]; // @[Modules.scala 143:103:@20002.4]
  assign _T_73269 = $signed(_T_73268); // @[Modules.scala 143:103:@20003.4]
  assign _T_73274 = $signed(_T_60920) + $signed(_T_54829); // @[Modules.scala 143:103:@20007.4]
  assign _T_73275 = _T_73274[4:0]; // @[Modules.scala 143:103:@20008.4]
  assign _T_73276 = $signed(_T_73275); // @[Modules.scala 143:103:@20009.4]
  assign _T_73281 = $signed(_T_54831) + $signed(_T_54836); // @[Modules.scala 143:103:@20013.4]
  assign _T_73282 = _T_73281[4:0]; // @[Modules.scala 143:103:@20014.4]
  assign _T_73283 = $signed(_T_73282); // @[Modules.scala 143:103:@20015.4]
  assign _GEN_453 = {{1{_T_54838[4]}},_T_54838}; // @[Modules.scala 143:103:@20019.4]
  assign _T_73288 = $signed(_GEN_453) + $signed(_T_54845); // @[Modules.scala 143:103:@20019.4]
  assign _T_73289 = _T_73288[5:0]; // @[Modules.scala 143:103:@20020.4]
  assign _T_73290 = $signed(_T_73289); // @[Modules.scala 143:103:@20021.4]
  assign _GEN_454 = {{1{_T_54878[4]}},_T_54878}; // @[Modules.scala 143:103:@20037.4]
  assign _T_73309 = $signed(_T_57899) + $signed(_GEN_454); // @[Modules.scala 143:103:@20037.4]
  assign _T_73310 = _T_73309[5:0]; // @[Modules.scala 143:103:@20038.4]
  assign _T_73311 = $signed(_T_73310); // @[Modules.scala 143:103:@20039.4]
  assign _T_73316 = $signed(_T_54880) + $signed(_T_54885); // @[Modules.scala 143:103:@20043.4]
  assign _T_73317 = _T_73316[4:0]; // @[Modules.scala 143:103:@20044.4]
  assign _T_73318 = $signed(_T_73317); // @[Modules.scala 143:103:@20045.4]
  assign _GEN_455 = {{1{_T_54887[4]}},_T_54887}; // @[Modules.scala 143:103:@20049.4]
  assign _T_73323 = $signed(_GEN_455) + $signed(_T_70213); // @[Modules.scala 143:103:@20049.4]
  assign _T_73324 = _T_73323[5:0]; // @[Modules.scala 143:103:@20050.4]
  assign _T_73325 = $signed(_T_73324); // @[Modules.scala 143:103:@20051.4]
  assign _T_73344 = $signed(_T_67200) + $signed(_T_64103); // @[Modules.scala 143:103:@20067.4]
  assign _T_73345 = _T_73344[5:0]; // @[Modules.scala 143:103:@20068.4]
  assign _T_73346 = $signed(_T_73345); // @[Modules.scala 143:103:@20069.4]
  assign _T_73386 = $signed(_T_57976) + $signed(_T_57981); // @[Modules.scala 143:103:@20103.4]
  assign _T_73387 = _T_73386[5:0]; // @[Modules.scala 143:103:@20104.4]
  assign _T_73388 = $signed(_T_73387); // @[Modules.scala 143:103:@20105.4]
  assign _GEN_457 = {{1{_T_54969[4]}},_T_54969}; // @[Modules.scala 143:103:@20109.4]
  assign _T_73393 = $signed(_T_57983) + $signed(_GEN_457); // @[Modules.scala 143:103:@20109.4]
  assign _T_73394 = _T_73393[5:0]; // @[Modules.scala 143:103:@20110.4]
  assign _T_73395 = $signed(_T_73394); // @[Modules.scala 143:103:@20111.4]
  assign _GEN_458 = {{1{_T_54978[4]}},_T_54978}; // @[Modules.scala 143:103:@20121.4]
  assign _T_73407 = $signed(_GEN_458) + $signed(_T_64171); // @[Modules.scala 143:103:@20121.4]
  assign _T_73408 = _T_73407[5:0]; // @[Modules.scala 143:103:@20122.4]
  assign _T_73409 = $signed(_T_73408); // @[Modules.scala 143:103:@20123.4]
  assign _GEN_459 = {{1{_T_55006[4]}},_T_55006}; // @[Modules.scala 143:103:@20145.4]
  assign _T_73435 = $signed(_T_64194) + $signed(_GEN_459); // @[Modules.scala 143:103:@20145.4]
  assign _T_73436 = _T_73435[5:0]; // @[Modules.scala 143:103:@20146.4]
  assign _T_73437 = $signed(_T_73436); // @[Modules.scala 143:103:@20147.4]
  assign _T_73463 = $signed(_GEN_28) + $signed(_T_58058); // @[Modules.scala 143:103:@20169.4]
  assign _T_73464 = _T_73463[5:0]; // @[Modules.scala 143:103:@20170.4]
  assign _T_73465 = $signed(_T_73464); // @[Modules.scala 143:103:@20171.4]
  assign _T_73505 = $signed(_T_58100) + $signed(_T_55076); // @[Modules.scala 143:103:@20205.4]
  assign _T_73506 = _T_73505[5:0]; // @[Modules.scala 143:103:@20206.4]
  assign _T_73507 = $signed(_T_73506); // @[Modules.scala 143:103:@20207.4]
  assign _GEN_461 = {{1{_T_55090[4]}},_T_55090}; // @[Modules.scala 143:103:@20217.4]
  assign _T_73519 = $signed(_T_58116) + $signed(_GEN_461); // @[Modules.scala 143:103:@20217.4]
  assign _T_73520 = _T_73519[5:0]; // @[Modules.scala 143:103:@20218.4]
  assign _T_73521 = $signed(_T_73520); // @[Modules.scala 143:103:@20219.4]
  assign _T_73554 = $signed(_GEN_172) + $signed(_T_55125); // @[Modules.scala 143:103:@20247.4]
  assign _T_73555 = _T_73554[5:0]; // @[Modules.scala 143:103:@20248.4]
  assign _T_73556 = $signed(_T_73555); // @[Modules.scala 143:103:@20249.4]
  assign _T_73561 = $signed(_T_58151) + $signed(_T_58156); // @[Modules.scala 143:103:@20253.4]
  assign _T_73562 = _T_73561[5:0]; // @[Modules.scala 143:103:@20254.4]
  assign _T_73563 = $signed(_T_73562); // @[Modules.scala 143:103:@20255.4]
  assign _T_73565 = $signed(-4'sh1) * $signed(io_in_354); // @[Modules.scala 143:74:@20257.4]
  assign _GEN_463 = {{1{_T_73565[4]}},_T_73565}; // @[Modules.scala 143:103:@20259.4]
  assign _T_73568 = $signed(_GEN_463) + $signed(_T_58163); // @[Modules.scala 143:103:@20259.4]
  assign _T_73569 = _T_73568[5:0]; // @[Modules.scala 143:103:@20260.4]
  assign _T_73570 = $signed(_T_73569); // @[Modules.scala 143:103:@20261.4]
  assign _T_73589 = $signed(_GEN_103) + $signed(_T_58177); // @[Modules.scala 143:103:@20277.4]
  assign _T_73590 = _T_73589[5:0]; // @[Modules.scala 143:103:@20278.4]
  assign _T_73591 = $signed(_T_73590); // @[Modules.scala 143:103:@20279.4]
  assign _T_73596 = $signed(_T_64355) + $signed(_T_55160); // @[Modules.scala 143:103:@20283.4]
  assign _T_73597 = _T_73596[5:0]; // @[Modules.scala 143:103:@20284.4]
  assign _T_73598 = $signed(_T_73597); // @[Modules.scala 143:103:@20285.4]
  assign _GEN_466 = {{1{_T_55181[4]}},_T_55181}; // @[Modules.scala 143:103:@20301.4]
  assign _T_73617 = $signed(_T_58200) + $signed(_GEN_466); // @[Modules.scala 143:103:@20301.4]
  assign _T_73618 = _T_73617[5:0]; // @[Modules.scala 143:103:@20302.4]
  assign _T_73619 = $signed(_T_73618); // @[Modules.scala 143:103:@20303.4]
  assign _T_73652 = $signed(_T_61284) + $signed(_T_70491); // @[Modules.scala 143:103:@20331.4]
  assign _T_73653 = _T_73652[4:0]; // @[Modules.scala 143:103:@20332.4]
  assign _T_73654 = $signed(_T_73653); // @[Modules.scala 143:103:@20333.4]
  assign _T_73663 = $signed(-4'sh1) * $signed(io_in_382); // @[Modules.scala 143:74:@20341.4]
  assign _T_73666 = $signed(_T_73663) + $signed(_T_55223); // @[Modules.scala 143:103:@20343.4]
  assign _T_73667 = _T_73666[4:0]; // @[Modules.scala 143:103:@20344.4]
  assign _T_73668 = $signed(_T_73667); // @[Modules.scala 143:103:@20345.4]
  assign _T_73764 = $signed(_T_58326) + $signed(_T_58331); // @[Modules.scala 143:103:@20427.4]
  assign _T_73765 = _T_73764[4:0]; // @[Modules.scala 143:103:@20428.4]
  assign _T_73766 = $signed(_T_73765); // @[Modules.scala 143:103:@20429.4]
  assign _GEN_469 = {{1{_T_58352[4]}},_T_58352}; // @[Modules.scala 143:103:@20451.4]
  assign _T_73792 = $signed(_GEN_469) + $signed(_T_61419); // @[Modules.scala 143:103:@20451.4]
  assign _T_73793 = _T_73792[5:0]; // @[Modules.scala 143:103:@20452.4]
  assign _T_73794 = $signed(_T_73793); // @[Modules.scala 143:103:@20453.4]
  assign _T_73806 = $signed(_T_58361) + $signed(_GEN_245); // @[Modules.scala 143:103:@20463.4]
  assign _T_73807 = _T_73806[5:0]; // @[Modules.scala 143:103:@20464.4]
  assign _T_73808 = $signed(_T_73807); // @[Modules.scala 143:103:@20465.4]
  assign _T_73834 = $signed(_T_61466) + $signed(_T_55384); // @[Modules.scala 143:103:@20487.4]
  assign _T_73835 = _T_73834[5:0]; // @[Modules.scala 143:103:@20488.4]
  assign _T_73836 = $signed(_T_73835); // @[Modules.scala 143:103:@20489.4]
  assign _T_73848 = $signed(_T_55398) + $signed(_T_55403); // @[Modules.scala 143:103:@20499.4]
  assign _T_73849 = _T_73848[4:0]; // @[Modules.scala 143:103:@20500.4]
  assign _T_73850 = $signed(_T_73849); // @[Modules.scala 143:103:@20501.4]
  assign _GEN_471 = {{1{_T_58410[4]}},_T_58410}; // @[Modules.scala 143:103:@20505.4]
  assign _T_73855 = $signed(_GEN_471) + $signed(_T_55405); // @[Modules.scala 143:103:@20505.4]
  assign _T_73856 = _T_73855[5:0]; // @[Modules.scala 143:103:@20506.4]
  assign _T_73857 = $signed(_T_73856); // @[Modules.scala 143:103:@20507.4]
  assign _T_73869 = $signed(_GEN_179) + $signed(_T_55424); // @[Modules.scala 143:103:@20517.4]
  assign _T_73870 = _T_73869[5:0]; // @[Modules.scala 143:103:@20518.4]
  assign _T_73871 = $signed(_T_73870); // @[Modules.scala 143:103:@20519.4]
  assign _T_73890 = $signed(_T_55438) + $signed(_T_64635); // @[Modules.scala 143:103:@20535.4]
  assign _T_73891 = _T_73890[5:0]; // @[Modules.scala 143:103:@20536.4]
  assign _T_73892 = $signed(_T_73891); // @[Modules.scala 143:103:@20537.4]
  assign _T_73904 = $signed(_T_64649) + $signed(_T_55452); // @[Modules.scala 143:103:@20547.4]
  assign _T_73905 = _T_73904[5:0]; // @[Modules.scala 143:103:@20548.4]
  assign _T_73906 = $signed(_T_73905); // @[Modules.scala 143:103:@20549.4]
  assign _T_73925 = $signed(_T_55468) + $signed(_T_61557); // @[Modules.scala 143:103:@20565.4]
  assign _T_73926 = _T_73925[5:0]; // @[Modules.scala 143:103:@20566.4]
  assign _T_73927 = $signed(_T_73926); // @[Modules.scala 143:103:@20567.4]
  assign _T_73932 = $signed(_T_55473) + $signed(_T_58485); // @[Modules.scala 143:103:@20571.4]
  assign _T_73933 = _T_73932[5:0]; // @[Modules.scala 143:103:@20572.4]
  assign _T_73934 = $signed(_T_73933); // @[Modules.scala 143:103:@20573.4]
  assign _T_73936 = $signed(4'sh1) * $signed(io_in_471); // @[Modules.scala 143:74:@20575.4]
  assign _T_73939 = $signed(_T_73936) + $signed(_T_70766); // @[Modules.scala 143:103:@20577.4]
  assign _T_73940 = _T_73939[5:0]; // @[Modules.scala 143:103:@20578.4]
  assign _T_73941 = $signed(_T_73940); // @[Modules.scala 143:103:@20579.4]
  assign _T_73953 = $signed(_T_58501) + $signed(_T_61580); // @[Modules.scala 143:103:@20589.4]
  assign _T_73954 = _T_73953[5:0]; // @[Modules.scala 143:103:@20590.4]
  assign _T_73955 = $signed(_T_73954); // @[Modules.scala 143:103:@20591.4]
  assign _T_73960 = $signed(_T_55489) + $signed(_T_55494); // @[Modules.scala 143:103:@20595.4]
  assign _T_73961 = _T_73960[5:0]; // @[Modules.scala 143:103:@20596.4]
  assign _T_73962 = $signed(_T_73961); // @[Modules.scala 143:103:@20597.4]
  assign _T_73967 = $signed(_T_55496) + $signed(_T_70799); // @[Modules.scala 143:103:@20601.4]
  assign _T_73968 = _T_73967[5:0]; // @[Modules.scala 143:103:@20602.4]
  assign _T_73969 = $signed(_T_73968); // @[Modules.scala 143:103:@20603.4]
  assign _T_73974 = $signed(_T_55501) + $signed(_T_61601); // @[Modules.scala 143:103:@20607.4]
  assign _T_73975 = _T_73974[5:0]; // @[Modules.scala 143:103:@20608.4]
  assign _T_73976 = $signed(_T_73975); // @[Modules.scala 143:103:@20609.4]
  assign _GEN_473 = {{1{_T_70815[4]}},_T_70815}; // @[Modules.scala 143:103:@20625.4]
  assign _T_73995 = $signed(_GEN_473) + $signed(_T_55522); // @[Modules.scala 143:103:@20625.4]
  assign _T_73996 = _T_73995[5:0]; // @[Modules.scala 143:103:@20626.4]
  assign _T_73997 = $signed(_T_73996); // @[Modules.scala 143:103:@20627.4]
  assign _T_74009 = $signed(_T_70829) + $signed(_T_58557); // @[Modules.scala 143:103:@20637.4]
  assign _T_74010 = _T_74009[5:0]; // @[Modules.scala 143:103:@20638.4]
  assign _T_74011 = $signed(_T_74010); // @[Modules.scala 143:103:@20639.4]
  assign _T_74023 = $signed(_T_55538) + $signed(_T_58569); // @[Modules.scala 143:103:@20649.4]
  assign _T_74024 = _T_74023[5:0]; // @[Modules.scala 143:103:@20650.4]
  assign _T_74025 = $signed(_T_74024); // @[Modules.scala 143:103:@20651.4]
  assign _GEN_475 = {{1{_T_58620[4]}},_T_58620}; // @[Modules.scala 143:103:@20703.4]
  assign _T_74086 = $signed(_GEN_475) + $signed(_T_55601); // @[Modules.scala 143:103:@20703.4]
  assign _T_74087 = _T_74086[5:0]; // @[Modules.scala 143:103:@20704.4]
  assign _T_74088 = $signed(_T_74087); // @[Modules.scala 143:103:@20705.4]
  assign _T_74093 = $signed(_T_55606) + $signed(_T_58632); // @[Modules.scala 143:103:@20709.4]
  assign _T_74094 = _T_74093[5:0]; // @[Modules.scala 143:103:@20710.4]
  assign _T_74095 = $signed(_T_74094); // @[Modules.scala 143:103:@20711.4]
  assign _T_74100 = $signed(_GEN_409) + $signed(_T_70918); // @[Modules.scala 143:103:@20715.4]
  assign _T_74101 = _T_74100[5:0]; // @[Modules.scala 143:103:@20716.4]
  assign _T_74102 = $signed(_T_74101); // @[Modules.scala 143:103:@20717.4]
  assign _GEN_478 = {{1{_T_58681[4]}},_T_58681}; // @[Modules.scala 143:103:@20757.4]
  assign _T_74149 = $signed(_T_70960) + $signed(_GEN_478); // @[Modules.scala 143:103:@20757.4]
  assign _T_74150 = _T_74149[5:0]; // @[Modules.scala 143:103:@20758.4]
  assign _T_74151 = $signed(_T_74150); // @[Modules.scala 143:103:@20759.4]
  assign _T_74170 = $signed(_T_55692) + $signed(_T_55697); // @[Modules.scala 143:103:@20775.4]
  assign _T_74171 = _T_74170[5:0]; // @[Modules.scala 143:103:@20776.4]
  assign _T_74172 = $signed(_T_74171); // @[Modules.scala 143:103:@20777.4]
  assign _T_74177 = $signed(_T_55699) + $signed(_T_55704); // @[Modules.scala 143:103:@20781.4]
  assign _T_74178 = _T_74177[5:0]; // @[Modules.scala 143:103:@20782.4]
  assign _T_74179 = $signed(_T_74178); // @[Modules.scala 143:103:@20783.4]
  assign _T_74184 = $signed(_T_70990) + $signed(_T_55706); // @[Modules.scala 143:103:@20787.4]
  assign _T_74185 = _T_74184[5:0]; // @[Modules.scala 143:103:@20788.4]
  assign _T_74186 = $signed(_T_74185); // @[Modules.scala 143:103:@20789.4]
  assign _T_74191 = $signed(_T_67928) + $signed(_T_58718); // @[Modules.scala 143:103:@20793.4]
  assign _T_74192 = _T_74191[4:0]; // @[Modules.scala 143:103:@20794.4]
  assign _T_74193 = $signed(_T_74192); // @[Modules.scala 143:103:@20795.4]
  assign _GEN_479 = {{1{_T_58723[4]}},_T_58723}; // @[Modules.scala 143:103:@20799.4]
  assign _T_74198 = $signed(_GEN_479) + $signed(_T_71009); // @[Modules.scala 143:103:@20799.4]
  assign _T_74199 = _T_74198[5:0]; // @[Modules.scala 143:103:@20800.4]
  assign _T_74200 = $signed(_T_74199); // @[Modules.scala 143:103:@20801.4]
  assign _T_74205 = $signed(_T_55713) + $signed(_T_55718); // @[Modules.scala 143:103:@20805.4]
  assign _T_74206 = _T_74205[5:0]; // @[Modules.scala 143:103:@20806.4]
  assign _T_74207 = $signed(_T_74206); // @[Modules.scala 143:103:@20807.4]
  assign _T_74212 = $signed(_T_55720) + $signed(_GEN_62); // @[Modules.scala 143:103:@20811.4]
  assign _T_74213 = _T_74212[5:0]; // @[Modules.scala 143:103:@20812.4]
  assign _T_74214 = $signed(_T_74213); // @[Modules.scala 143:103:@20813.4]
  assign _GEN_481 = {{1{_T_64948[4]}},_T_64948}; // @[Modules.scala 143:103:@20817.4]
  assign _T_74219 = $signed(_GEN_481) + $signed(_T_55727); // @[Modules.scala 143:103:@20817.4]
  assign _T_74220 = _T_74219[5:0]; // @[Modules.scala 143:103:@20818.4]
  assign _T_74221 = $signed(_T_74220); // @[Modules.scala 143:103:@20819.4]
  assign _GEN_482 = {{1{_T_61832[4]}},_T_61832}; // @[Modules.scala 143:103:@20835.4]
  assign _T_74240 = $signed(_T_55746) + $signed(_GEN_482); // @[Modules.scala 143:103:@20835.4]
  assign _T_74241 = _T_74240[5:0]; // @[Modules.scala 143:103:@20836.4]
  assign _T_74242 = $signed(_T_74241); // @[Modules.scala 143:103:@20837.4]
  assign _T_74260 = $signed(4'sh1) * $signed(io_in_577); // @[Modules.scala 144:80:@20852.4]
  assign _T_74261 = $signed(_T_61851) + $signed(_T_74260); // @[Modules.scala 143:103:@20853.4]
  assign _T_74262 = _T_74261[5:0]; // @[Modules.scala 143:103:@20854.4]
  assign _T_74263 = $signed(_T_74262); // @[Modules.scala 143:103:@20855.4]
  assign _T_74289 = $signed(_T_58809) + $signed(_GEN_342); // @[Modules.scala 143:103:@20877.4]
  assign _T_74290 = _T_74289[5:0]; // @[Modules.scala 143:103:@20878.4]
  assign _T_74291 = $signed(_T_74290); // @[Modules.scala 143:103:@20879.4]
  assign _T_74296 = $signed(_GEN_416) + $signed(_T_55797); // @[Modules.scala 143:103:@20883.4]
  assign _T_74297 = _T_74296[5:0]; // @[Modules.scala 143:103:@20884.4]
  assign _T_74298 = $signed(_T_74297); // @[Modules.scala 143:103:@20885.4]
  assign _T_74310 = $signed(_T_55809) + $signed(_T_61923); // @[Modules.scala 143:103:@20895.4]
  assign _T_74311 = _T_74310[5:0]; // @[Modules.scala 143:103:@20896.4]
  assign _T_74312 = $signed(_T_74311); // @[Modules.scala 143:103:@20897.4]
  assign _T_74317 = $signed(_T_58849) + $signed(_T_71163); // @[Modules.scala 143:103:@20901.4]
  assign _T_74318 = _T_74317[4:0]; // @[Modules.scala 143:103:@20902.4]
  assign _T_74319 = $signed(_T_74318); // @[Modules.scala 143:103:@20903.4]
  assign _T_74323 = $signed(4'sh1) * $signed(io_in_604); // @[Modules.scala 144:80:@20906.4]
  assign _GEN_485 = {{1{_T_68075[4]}},_T_68075}; // @[Modules.scala 143:103:@20907.4]
  assign _T_74324 = $signed(_GEN_485) + $signed(_T_74323); // @[Modules.scala 143:103:@20907.4]
  assign _T_74325 = _T_74324[5:0]; // @[Modules.scala 143:103:@20908.4]
  assign _T_74326 = $signed(_T_74325); // @[Modules.scala 143:103:@20909.4]
  assign _T_74330 = $signed(4'sh1) * $signed(io_in_606); // @[Modules.scala 144:80:@20912.4]
  assign _T_74331 = $signed(_T_61937) + $signed(_T_74330); // @[Modules.scala 143:103:@20913.4]
  assign _T_74332 = _T_74331[5:0]; // @[Modules.scala 143:103:@20914.4]
  assign _T_74333 = $signed(_T_74332); // @[Modules.scala 143:103:@20915.4]
  assign _T_74338 = $signed(_T_71179) + $signed(_T_55839); // @[Modules.scala 143:103:@20919.4]
  assign _T_74339 = _T_74338[5:0]; // @[Modules.scala 143:103:@20920.4]
  assign _T_74340 = $signed(_T_74339); // @[Modules.scala 143:103:@20921.4]
  assign _GEN_486 = {{1{_T_58870[4]}},_T_58870}; // @[Modules.scala 143:103:@20925.4]
  assign _T_74345 = $signed(_GEN_486) + $signed(_T_55851); // @[Modules.scala 143:103:@20925.4]
  assign _T_74346 = _T_74345[5:0]; // @[Modules.scala 143:103:@20926.4]
  assign _T_74347 = $signed(_T_74346); // @[Modules.scala 143:103:@20927.4]
  assign _T_74352 = $signed(_T_55853) + $signed(_T_55858); // @[Modules.scala 143:103:@20931.4]
  assign _T_74353 = _T_74352[5:0]; // @[Modules.scala 143:103:@20932.4]
  assign _T_74354 = $signed(_T_74353); // @[Modules.scala 143:103:@20933.4]
  assign _T_74359 = $signed(_T_58886) + $signed(_T_58891); // @[Modules.scala 143:103:@20937.4]
  assign _T_74360 = _T_74359[4:0]; // @[Modules.scala 143:103:@20938.4]
  assign _T_74361 = $signed(_T_74360); // @[Modules.scala 143:103:@20939.4]
  assign _T_74366 = $signed(_T_55867) + $signed(_T_55872); // @[Modules.scala 143:103:@20943.4]
  assign _T_74367 = _T_74366[5:0]; // @[Modules.scala 143:103:@20944.4]
  assign _T_74368 = $signed(_T_74367); // @[Modules.scala 143:103:@20945.4]
  assign _T_74373 = $signed(_T_55874) + $signed(_T_55879); // @[Modules.scala 143:103:@20949.4]
  assign _T_74374 = _T_74373[5:0]; // @[Modules.scala 143:103:@20950.4]
  assign _T_74375 = $signed(_T_74374); // @[Modules.scala 143:103:@20951.4]
  assign _T_74380 = $signed(_T_55881) + $signed(_GEN_66); // @[Modules.scala 143:103:@20955.4]
  assign _T_74381 = _T_74380[5:0]; // @[Modules.scala 143:103:@20956.4]
  assign _T_74382 = $signed(_T_74381); // @[Modules.scala 143:103:@20957.4]
  assign _T_74408 = $signed(_GEN_419) + $signed(_T_55921); // @[Modules.scala 143:103:@20979.4]
  assign _T_74409 = _T_74408[5:0]; // @[Modules.scala 143:103:@20980.4]
  assign _T_74410 = $signed(_T_74409); // @[Modules.scala 143:103:@20981.4]
  assign _T_74415 = $signed(_T_55923) + $signed(_T_55928); // @[Modules.scala 143:103:@20985.4]
  assign _T_74416 = _T_74415[5:0]; // @[Modules.scala 143:103:@20986.4]
  assign _T_74417 = $signed(_T_74416); // @[Modules.scala 143:103:@20987.4]
  assign _T_74422 = $signed(_T_55930) + $signed(_T_55935); // @[Modules.scala 143:103:@20991.4]
  assign _T_74423 = _T_74422[5:0]; // @[Modules.scala 143:103:@20992.4]
  assign _T_74424 = $signed(_T_74423); // @[Modules.scala 143:103:@20993.4]
  assign _T_74429 = $signed(_T_55937) + $signed(_T_55942); // @[Modules.scala 143:103:@20997.4]
  assign _T_74430 = _T_74429[5:0]; // @[Modules.scala 143:103:@20998.4]
  assign _T_74431 = $signed(_T_74430); // @[Modules.scala 143:103:@20999.4]
  assign _T_74450 = $signed(_T_55958) + $signed(_T_55963); // @[Modules.scala 143:103:@21015.4]
  assign _T_74451 = _T_74450[5:0]; // @[Modules.scala 143:103:@21016.4]
  assign _T_74452 = $signed(_T_74451); // @[Modules.scala 143:103:@21017.4]
  assign _GEN_490 = {{1{_T_55977[4]}},_T_55977}; // @[Modules.scala 143:103:@21021.4]
  assign _T_74457 = $signed(_T_55965) + $signed(_GEN_490); // @[Modules.scala 143:103:@21021.4]
  assign _T_74458 = _T_74457[5:0]; // @[Modules.scala 143:103:@21022.4]
  assign _T_74459 = $signed(_T_74458); // @[Modules.scala 143:103:@21023.4]
  assign _T_74464 = $signed(_T_55979) + $signed(_T_55984); // @[Modules.scala 143:103:@21027.4]
  assign _T_74465 = _T_74464[4:0]; // @[Modules.scala 143:103:@21028.4]
  assign _T_74466 = $signed(_T_74465); // @[Modules.scala 143:103:@21029.4]
  assign _T_74485 = $signed(_T_56000) + $signed(_T_56005); // @[Modules.scala 143:103:@21045.4]
  assign _T_74486 = _T_74485[4:0]; // @[Modules.scala 143:103:@21046.4]
  assign _T_74487 = $signed(_T_74486); // @[Modules.scala 143:103:@21047.4]
  assign _T_74492 = $signed(_T_56007) + $signed(_T_56014); // @[Modules.scala 143:103:@21051.4]
  assign _T_74493 = _T_74492[4:0]; // @[Modules.scala 143:103:@21052.4]
  assign _T_74494 = $signed(_T_74493); // @[Modules.scala 143:103:@21053.4]
  assign _T_74499 = $signed(_T_65221) + $signed(_T_56019); // @[Modules.scala 143:103:@21057.4]
  assign _T_74500 = _T_74499[5:0]; // @[Modules.scala 143:103:@21058.4]
  assign _T_74501 = $signed(_T_74500); // @[Modules.scala 143:103:@21059.4]
  assign _T_74506 = $signed(_T_68257) + $signed(_T_56021); // @[Modules.scala 143:103:@21063.4]
  assign _T_74507 = _T_74506[5:0]; // @[Modules.scala 143:103:@21064.4]
  assign _T_74508 = $signed(_T_74507); // @[Modules.scala 143:103:@21065.4]
  assign _T_74513 = $signed(_T_59033) + $signed(_T_56033); // @[Modules.scala 143:103:@21069.4]
  assign _T_74514 = _T_74513[5:0]; // @[Modules.scala 143:103:@21070.4]
  assign _T_74515 = $signed(_T_74514); // @[Modules.scala 143:103:@21071.4]
  assign _T_74520 = $signed(_T_56035) + $signed(_T_56040); // @[Modules.scala 143:103:@21075.4]
  assign _T_74521 = _T_74520[5:0]; // @[Modules.scala 143:103:@21076.4]
  assign _T_74522 = $signed(_T_74521); // @[Modules.scala 143:103:@21077.4]
  assign _T_74527 = $signed(_T_56042) + $signed(_T_56047); // @[Modules.scala 143:103:@21081.4]
  assign _T_74528 = _T_74527[5:0]; // @[Modules.scala 143:103:@21082.4]
  assign _T_74529 = $signed(_T_74528); // @[Modules.scala 143:103:@21083.4]
  assign _T_74555 = $signed(_T_56070) + $signed(_T_56075); // @[Modules.scala 143:103:@21105.4]
  assign _T_74556 = _T_74555[4:0]; // @[Modules.scala 143:103:@21106.4]
  assign _T_74557 = $signed(_T_74556); // @[Modules.scala 143:103:@21107.4]
  assign _T_74562 = $signed(_T_56077) + $signed(_T_56082); // @[Modules.scala 143:103:@21111.4]
  assign _T_74563 = _T_74562[4:0]; // @[Modules.scala 143:103:@21112.4]
  assign _T_74564 = $signed(_T_74563); // @[Modules.scala 143:103:@21113.4]
  assign _T_74569 = $signed(_T_56084) + $signed(_T_56089); // @[Modules.scala 143:103:@21117.4]
  assign _T_74570 = _T_74569[4:0]; // @[Modules.scala 143:103:@21118.4]
  assign _T_74571 = $signed(_T_74570); // @[Modules.scala 143:103:@21119.4]
  assign _T_74583 = $signed(_T_56098) + $signed(_T_56103); // @[Modules.scala 143:103:@21129.4]
  assign _T_74584 = _T_74583[5:0]; // @[Modules.scala 143:103:@21130.4]
  assign _T_74585 = $signed(_T_74584); // @[Modules.scala 143:103:@21131.4]
  assign _T_74590 = $signed(_T_56105) + $signed(_T_56110); // @[Modules.scala 143:103:@21135.4]
  assign _T_74591 = _T_74590[5:0]; // @[Modules.scala 143:103:@21136.4]
  assign _T_74592 = $signed(_T_74591); // @[Modules.scala 143:103:@21137.4]
  assign _T_74597 = $signed(_T_56112) + $signed(_T_56117); // @[Modules.scala 143:103:@21141.4]
  assign _T_74598 = _T_74597[5:0]; // @[Modules.scala 143:103:@21142.4]
  assign _T_74599 = $signed(_T_74598); // @[Modules.scala 143:103:@21143.4]
  assign _T_74604 = $signed(_T_59124) + $signed(_T_59129); // @[Modules.scala 143:103:@21147.4]
  assign _T_74605 = _T_74604[5:0]; // @[Modules.scala 143:103:@21148.4]
  assign _T_74606 = $signed(_T_74605); // @[Modules.scala 143:103:@21149.4]
  assign _T_74611 = $signed(_T_59131) + $signed(_T_56126); // @[Modules.scala 143:103:@21153.4]
  assign _T_74612 = _T_74611[5:0]; // @[Modules.scala 143:103:@21154.4]
  assign _T_74613 = $signed(_T_74612); // @[Modules.scala 143:103:@21155.4]
  assign _T_74632 = $signed(_T_59152) + $signed(_T_59157); // @[Modules.scala 143:103:@21171.4]
  assign _T_74633 = _T_74632[5:0]; // @[Modules.scala 143:103:@21172.4]
  assign _T_74634 = $signed(_T_74633); // @[Modules.scala 143:103:@21173.4]
  assign _T_74646 = $signed(_T_56161) + $signed(_T_56166); // @[Modules.scala 143:103:@21183.4]
  assign _T_74647 = _T_74646[4:0]; // @[Modules.scala 143:103:@21184.4]
  assign _T_74648 = $signed(_T_74647); // @[Modules.scala 143:103:@21185.4]
  assign _T_74653 = $signed(_T_56168) + $signed(_T_56173); // @[Modules.scala 143:103:@21189.4]
  assign _T_74654 = _T_74653[4:0]; // @[Modules.scala 143:103:@21190.4]
  assign _T_74655 = $signed(_T_74654); // @[Modules.scala 143:103:@21191.4]
  assign _T_74660 = $signed(_T_56175) + $signed(_T_56180); // @[Modules.scala 143:103:@21195.4]
  assign _T_74661 = _T_74660[4:0]; // @[Modules.scala 143:103:@21196.4]
  assign _T_74662 = $signed(_T_74661); // @[Modules.scala 143:103:@21197.4]
  assign _GEN_492 = {{1{_T_56182[4]}},_T_56182}; // @[Modules.scala 143:103:@21201.4]
  assign _T_74667 = $signed(_GEN_492) + $signed(_T_59185); // @[Modules.scala 143:103:@21201.4]
  assign _T_74668 = _T_74667[5:0]; // @[Modules.scala 143:103:@21202.4]
  assign _T_74669 = $signed(_T_74668); // @[Modules.scala 143:103:@21203.4]
  assign _T_74674 = $signed(_T_62273) + $signed(_GEN_72); // @[Modules.scala 143:103:@21207.4]
  assign _T_74675 = _T_74674[5:0]; // @[Modules.scala 143:103:@21208.4]
  assign _T_74676 = $signed(_T_74675); // @[Modules.scala 143:103:@21209.4]
  assign _GEN_494 = {{1{_T_59194[4]}},_T_59194}; // @[Modules.scala 143:103:@21213.4]
  assign _T_74681 = $signed(_GEN_494) + $signed(_T_62285); // @[Modules.scala 143:103:@21213.4]
  assign _T_74682 = _T_74681[5:0]; // @[Modules.scala 143:103:@21214.4]
  assign _T_74683 = $signed(_T_74682); // @[Modules.scala 143:103:@21215.4]
  assign _T_74730 = $signed(_T_59243) + $signed(_GEN_216); // @[Modules.scala 143:103:@21255.4]
  assign _T_74731 = _T_74730[5:0]; // @[Modules.scala 143:103:@21256.4]
  assign _T_74732 = $signed(_T_74731); // @[Modules.scala 143:103:@21257.4]
  assign _T_74737 = $signed(_T_56231) + $signed(_T_56236); // @[Modules.scala 143:103:@21261.4]
  assign _T_74738 = _T_74737[4:0]; // @[Modules.scala 143:103:@21262.4]
  assign _T_74739 = $signed(_T_74738); // @[Modules.scala 143:103:@21263.4]
  assign _GEN_497 = {{1{_T_56294[4]}},_T_56294}; // @[Modules.scala 143:103:@21327.4]
  assign _T_74814 = $signed(_GEN_497) + $signed(_T_56306); // @[Modules.scala 143:103:@21327.4]
  assign _T_74815 = _T_74814[5:0]; // @[Modules.scala 143:103:@21328.4]
  assign _T_74816 = $signed(_T_74815); // @[Modules.scala 143:103:@21329.4]
  assign buffer_6_2 = {{8{_T_72625[5]}},_T_72625}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_3 = {{9{_T_72632[4]}},_T_72632}; // @[Modules.scala 112:22:@8.4]
  assign _T_74820 = $signed(buffer_6_2) + $signed(buffer_6_3); // @[Modules.scala 160:64:@21335.4]
  assign _T_74821 = _T_74820[13:0]; // @[Modules.scala 160:64:@21336.4]
  assign buffer_6_317 = $signed(_T_74821); // @[Modules.scala 160:64:@21337.4]
  assign buffer_6_4 = {{9{_T_72639[4]}},_T_72639}; // @[Modules.scala 112:22:@8.4]
  assign _T_74823 = $signed(buffer_6_4) + $signed(buffer_4_3); // @[Modules.scala 160:64:@21339.4]
  assign _T_74824 = _T_74823[13:0]; // @[Modules.scala 160:64:@21340.4]
  assign buffer_6_318 = $signed(_T_74824); // @[Modules.scala 160:64:@21341.4]
  assign buffer_6_8 = {{8{_T_72667[5]}},_T_72667}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_9 = {{8{_T_72674[5]}},_T_72674}; // @[Modules.scala 112:22:@8.4]
  assign _T_74829 = $signed(buffer_6_8) + $signed(buffer_6_9); // @[Modules.scala 160:64:@21347.4]
  assign _T_74830 = _T_74829[13:0]; // @[Modules.scala 160:64:@21348.4]
  assign buffer_6_320 = $signed(_T_74830); // @[Modules.scala 160:64:@21349.4]
  assign buffer_6_10 = {{8{_T_72681[5]}},_T_72681}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_11 = {{8{_T_72688[5]}},_T_72688}; // @[Modules.scala 112:22:@8.4]
  assign _T_74832 = $signed(buffer_6_10) + $signed(buffer_6_11); // @[Modules.scala 160:64:@21351.4]
  assign _T_74833 = _T_74832[13:0]; // @[Modules.scala 160:64:@21352.4]
  assign buffer_6_321 = $signed(_T_74833); // @[Modules.scala 160:64:@21353.4]
  assign _T_74835 = $signed(buffer_5_12) + $signed(buffer_2_12); // @[Modules.scala 160:64:@21355.4]
  assign _T_74836 = _T_74835[13:0]; // @[Modules.scala 160:64:@21356.4]
  assign buffer_6_322 = $signed(_T_74836); // @[Modules.scala 160:64:@21357.4]
  assign buffer_6_20 = {{9{_T_72751[4]}},_T_72751}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_21 = {{9{_T_72758[4]}},_T_72758}; // @[Modules.scala 112:22:@8.4]
  assign _T_74847 = $signed(buffer_6_20) + $signed(buffer_6_21); // @[Modules.scala 160:64:@21371.4]
  assign _T_74848 = _T_74847[13:0]; // @[Modules.scala 160:64:@21372.4]
  assign buffer_6_326 = $signed(_T_74848); // @[Modules.scala 160:64:@21373.4]
  assign buffer_6_22 = {{8{_T_72765[5]}},_T_72765}; // @[Modules.scala 112:22:@8.4]
  assign _T_74850 = $signed(buffer_6_22) + $signed(buffer_3_22); // @[Modules.scala 160:64:@21375.4]
  assign _T_74851 = _T_74850[13:0]; // @[Modules.scala 160:64:@21376.4]
  assign buffer_6_327 = $signed(_T_74851); // @[Modules.scala 160:64:@21377.4]
  assign buffer_6_25 = {{8{_T_72786[5]}},_T_72786}; // @[Modules.scala 112:22:@8.4]
  assign _T_74853 = $signed(buffer_1_24) + $signed(buffer_6_25); // @[Modules.scala 160:64:@21379.4]
  assign _T_74854 = _T_74853[13:0]; // @[Modules.scala 160:64:@21380.4]
  assign buffer_6_328 = $signed(_T_74854); // @[Modules.scala 160:64:@21381.4]
  assign buffer_6_26 = {{8{_T_72793[5]}},_T_72793}; // @[Modules.scala 112:22:@8.4]
  assign _T_74856 = $signed(buffer_6_26) + $signed(buffer_0_28); // @[Modules.scala 160:64:@21383.4]
  assign _T_74857 = _T_74856[13:0]; // @[Modules.scala 160:64:@21384.4]
  assign buffer_6_329 = $signed(_T_74857); // @[Modules.scala 160:64:@21385.4]
  assign buffer_6_29 = {{8{_T_72814[5]}},_T_72814}; // @[Modules.scala 112:22:@8.4]
  assign _T_74859 = $signed(buffer_0_29) + $signed(buffer_6_29); // @[Modules.scala 160:64:@21387.4]
  assign _T_74860 = _T_74859[13:0]; // @[Modules.scala 160:64:@21388.4]
  assign buffer_6_330 = $signed(_T_74860); // @[Modules.scala 160:64:@21389.4]
  assign buffer_6_30 = {{8{_T_72821[5]}},_T_72821}; // @[Modules.scala 112:22:@8.4]
  assign _T_74862 = $signed(buffer_6_30) + $signed(buffer_1_31); // @[Modules.scala 160:64:@21391.4]
  assign _T_74863 = _T_74862[13:0]; // @[Modules.scala 160:64:@21392.4]
  assign buffer_6_331 = $signed(_T_74863); // @[Modules.scala 160:64:@21393.4]
  assign buffer_6_33 = {{8{_T_72842[5]}},_T_72842}; // @[Modules.scala 112:22:@8.4]
  assign _T_74865 = $signed(buffer_1_32) + $signed(buffer_6_33); // @[Modules.scala 160:64:@21395.4]
  assign _T_74866 = _T_74865[13:0]; // @[Modules.scala 160:64:@21396.4]
  assign buffer_6_332 = $signed(_T_74866); // @[Modules.scala 160:64:@21397.4]
  assign buffer_6_35 = {{8{_T_72856[5]}},_T_72856}; // @[Modules.scala 112:22:@8.4]
  assign _T_74868 = $signed(buffer_1_34) + $signed(buffer_6_35); // @[Modules.scala 160:64:@21399.4]
  assign _T_74869 = _T_74868[13:0]; // @[Modules.scala 160:64:@21400.4]
  assign buffer_6_333 = $signed(_T_74869); // @[Modules.scala 160:64:@21401.4]
  assign buffer_6_39 = {{8{_T_72884[5]}},_T_72884}; // @[Modules.scala 112:22:@8.4]
  assign _T_74874 = $signed(buffer_1_38) + $signed(buffer_6_39); // @[Modules.scala 160:64:@21407.4]
  assign _T_74875 = _T_74874[13:0]; // @[Modules.scala 160:64:@21408.4]
  assign buffer_6_335 = $signed(_T_74875); // @[Modules.scala 160:64:@21409.4]
  assign buffer_6_44 = {{8{_T_72919[5]}},_T_72919}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_45 = {{8{_T_72926[5]}},_T_72926}; // @[Modules.scala 112:22:@8.4]
  assign _T_74883 = $signed(buffer_6_44) + $signed(buffer_6_45); // @[Modules.scala 160:64:@21419.4]
  assign _T_74884 = _T_74883[13:0]; // @[Modules.scala 160:64:@21420.4]
  assign buffer_6_338 = $signed(_T_74884); // @[Modules.scala 160:64:@21421.4]
  assign buffer_6_46 = {{8{_T_72933[5]}},_T_72933}; // @[Modules.scala 112:22:@8.4]
  assign _T_74886 = $signed(buffer_6_46) + $signed(buffer_2_46); // @[Modules.scala 160:64:@21423.4]
  assign _T_74887 = _T_74886[13:0]; // @[Modules.scala 160:64:@21424.4]
  assign buffer_6_339 = $signed(_T_74887); // @[Modules.scala 160:64:@21425.4]
  assign buffer_6_50 = {{8{_T_72961[5]}},_T_72961}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_51 = {{8{_T_72968[5]}},_T_72968}; // @[Modules.scala 112:22:@8.4]
  assign _T_74892 = $signed(buffer_6_50) + $signed(buffer_6_51); // @[Modules.scala 160:64:@21431.4]
  assign _T_74893 = _T_74892[13:0]; // @[Modules.scala 160:64:@21432.4]
  assign buffer_6_341 = $signed(_T_74893); // @[Modules.scala 160:64:@21433.4]
  assign _T_74895 = $signed(buffer_0_51) + $signed(buffer_0_52); // @[Modules.scala 160:64:@21435.4]
  assign _T_74896 = _T_74895[13:0]; // @[Modules.scala 160:64:@21436.4]
  assign buffer_6_342 = $signed(_T_74896); // @[Modules.scala 160:64:@21437.4]
  assign _T_74898 = $signed(buffer_4_55) + $signed(buffer_3_58); // @[Modules.scala 160:64:@21439.4]
  assign _T_74899 = _T_74898[13:0]; // @[Modules.scala 160:64:@21440.4]
  assign buffer_6_343 = $signed(_T_74899); // @[Modules.scala 160:64:@21441.4]
  assign buffer_6_56 = {{8{_T_73003[5]}},_T_73003}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_57 = {{8{_T_73010[5]}},_T_73010}; // @[Modules.scala 112:22:@8.4]
  assign _T_74901 = $signed(buffer_6_56) + $signed(buffer_6_57); // @[Modules.scala 160:64:@21443.4]
  assign _T_74902 = _T_74901[13:0]; // @[Modules.scala 160:64:@21444.4]
  assign buffer_6_344 = $signed(_T_74902); // @[Modules.scala 160:64:@21445.4]
  assign buffer_6_58 = {{8{_T_73017[5]}},_T_73017}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_59 = {{8{_T_73024[5]}},_T_73024}; // @[Modules.scala 112:22:@8.4]
  assign _T_74904 = $signed(buffer_6_58) + $signed(buffer_6_59); // @[Modules.scala 160:64:@21447.4]
  assign _T_74905 = _T_74904[13:0]; // @[Modules.scala 160:64:@21448.4]
  assign buffer_6_345 = $signed(_T_74905); // @[Modules.scala 160:64:@21449.4]
  assign buffer_6_60 = {{8{_T_73031[5]}},_T_73031}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_61 = {{8{_T_73038[5]}},_T_73038}; // @[Modules.scala 112:22:@8.4]
  assign _T_74907 = $signed(buffer_6_60) + $signed(buffer_6_61); // @[Modules.scala 160:64:@21451.4]
  assign _T_74908 = _T_74907[13:0]; // @[Modules.scala 160:64:@21452.4]
  assign buffer_6_346 = $signed(_T_74908); // @[Modules.scala 160:64:@21453.4]
  assign buffer_6_62 = {{8{_T_73045[5]}},_T_73045}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_63 = {{8{_T_73052[5]}},_T_73052}; // @[Modules.scala 112:22:@8.4]
  assign _T_74910 = $signed(buffer_6_62) + $signed(buffer_6_63); // @[Modules.scala 160:64:@21455.4]
  assign _T_74911 = _T_74910[13:0]; // @[Modules.scala 160:64:@21456.4]
  assign buffer_6_347 = $signed(_T_74911); // @[Modules.scala 160:64:@21457.4]
  assign buffer_6_66 = {{8{_T_73073[5]}},_T_73073}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_67 = {{8{_T_73080[5]}},_T_73080}; // @[Modules.scala 112:22:@8.4]
  assign _T_74916 = $signed(buffer_6_66) + $signed(buffer_6_67); // @[Modules.scala 160:64:@21463.4]
  assign _T_74917 = _T_74916[13:0]; // @[Modules.scala 160:64:@21464.4]
  assign buffer_6_349 = $signed(_T_74917); // @[Modules.scala 160:64:@21465.4]
  assign buffer_6_69 = {{8{_T_73094[5]}},_T_73094}; // @[Modules.scala 112:22:@8.4]
  assign _T_74919 = $signed(buffer_5_69) + $signed(buffer_6_69); // @[Modules.scala 160:64:@21467.4]
  assign _T_74920 = _T_74919[13:0]; // @[Modules.scala 160:64:@21468.4]
  assign buffer_6_350 = $signed(_T_74920); // @[Modules.scala 160:64:@21469.4]
  assign buffer_6_70 = {{8{_T_73101[5]}},_T_73101}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_71 = {{8{_T_73108[5]}},_T_73108}; // @[Modules.scala 112:22:@8.4]
  assign _T_74922 = $signed(buffer_6_70) + $signed(buffer_6_71); // @[Modules.scala 160:64:@21471.4]
  assign _T_74923 = _T_74922[13:0]; // @[Modules.scala 160:64:@21472.4]
  assign buffer_6_351 = $signed(_T_74923); // @[Modules.scala 160:64:@21473.4]
  assign buffer_6_73 = {{9{_T_73122[4]}},_T_73122}; // @[Modules.scala 112:22:@8.4]
  assign _T_74925 = $signed(buffer_1_71) + $signed(buffer_6_73); // @[Modules.scala 160:64:@21475.4]
  assign _T_74926 = _T_74925[13:0]; // @[Modules.scala 160:64:@21476.4]
  assign buffer_6_352 = $signed(_T_74926); // @[Modules.scala 160:64:@21477.4]
  assign buffer_6_74 = {{8{_T_73129[5]}},_T_73129}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_75 = {{8{_T_73136[5]}},_T_73136}; // @[Modules.scala 112:22:@8.4]
  assign _T_74928 = $signed(buffer_6_74) + $signed(buffer_6_75); // @[Modules.scala 160:64:@21479.4]
  assign _T_74929 = _T_74928[13:0]; // @[Modules.scala 160:64:@21480.4]
  assign buffer_6_353 = $signed(_T_74929); // @[Modules.scala 160:64:@21481.4]
  assign buffer_6_76 = {{9{_T_73143[4]}},_T_73143}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_77 = {{9{_T_73150[4]}},_T_73150}; // @[Modules.scala 112:22:@8.4]
  assign _T_74931 = $signed(buffer_6_76) + $signed(buffer_6_77); // @[Modules.scala 160:64:@21483.4]
  assign _T_74932 = _T_74931[13:0]; // @[Modules.scala 160:64:@21484.4]
  assign buffer_6_354 = $signed(_T_74932); // @[Modules.scala 160:64:@21485.4]
  assign buffer_6_78 = {{8{_T_73157[5]}},_T_73157}; // @[Modules.scala 112:22:@8.4]
  assign _T_74934 = $signed(buffer_6_78) + $signed(buffer_1_80); // @[Modules.scala 160:64:@21487.4]
  assign _T_74935 = _T_74934[13:0]; // @[Modules.scala 160:64:@21488.4]
  assign buffer_6_355 = $signed(_T_74935); // @[Modules.scala 160:64:@21489.4]
  assign buffer_6_81 = {{8{_T_73178[5]}},_T_73178}; // @[Modules.scala 112:22:@8.4]
  assign _T_74937 = $signed(buffer_1_81) + $signed(buffer_6_81); // @[Modules.scala 160:64:@21491.4]
  assign _T_74938 = _T_74937[13:0]; // @[Modules.scala 160:64:@21492.4]
  assign buffer_6_356 = $signed(_T_74938); // @[Modules.scala 160:64:@21493.4]
  assign buffer_6_82 = {{8{_T_73185[5]}},_T_73185}; // @[Modules.scala 112:22:@8.4]
  assign _T_74940 = $signed(buffer_6_82) + $signed(buffer_4_82); // @[Modules.scala 160:64:@21495.4]
  assign _T_74941 = _T_74940[13:0]; // @[Modules.scala 160:64:@21496.4]
  assign buffer_6_357 = $signed(_T_74941); // @[Modules.scala 160:64:@21497.4]
  assign buffer_6_88 = {{8{_T_73227[5]}},_T_73227}; // @[Modules.scala 112:22:@8.4]
  assign _T_74949 = $signed(buffer_6_88) + $signed(buffer_2_90); // @[Modules.scala 160:64:@21507.4]
  assign _T_74950 = _T_74949[13:0]; // @[Modules.scala 160:64:@21508.4]
  assign buffer_6_360 = $signed(_T_74950); // @[Modules.scala 160:64:@21509.4]
  assign buffer_6_90 = {{8{_T_73241[5]}},_T_73241}; // @[Modules.scala 112:22:@8.4]
  assign _T_74952 = $signed(buffer_6_90) + $signed(buffer_4_90); // @[Modules.scala 160:64:@21511.4]
  assign _T_74953 = _T_74952[13:0]; // @[Modules.scala 160:64:@21512.4]
  assign buffer_6_361 = $signed(_T_74953); // @[Modules.scala 160:64:@21513.4]
  assign buffer_6_94 = {{8{_T_73269[5]}},_T_73269}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_95 = {{9{_T_73276[4]}},_T_73276}; // @[Modules.scala 112:22:@8.4]
  assign _T_74958 = $signed(buffer_6_94) + $signed(buffer_6_95); // @[Modules.scala 160:64:@21519.4]
  assign _T_74959 = _T_74958[13:0]; // @[Modules.scala 160:64:@21520.4]
  assign buffer_6_363 = $signed(_T_74959); // @[Modules.scala 160:64:@21521.4]
  assign buffer_6_96 = {{9{_T_73283[4]}},_T_73283}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_97 = {{8{_T_73290[5]}},_T_73290}; // @[Modules.scala 112:22:@8.4]
  assign _T_74961 = $signed(buffer_6_96) + $signed(buffer_6_97); // @[Modules.scala 160:64:@21523.4]
  assign _T_74962 = _T_74961[13:0]; // @[Modules.scala 160:64:@21524.4]
  assign buffer_6_364 = $signed(_T_74962); // @[Modules.scala 160:64:@21525.4]
  assign _T_74964 = $signed(buffer_4_95) + $signed(buffer_4_96); // @[Modules.scala 160:64:@21527.4]
  assign _T_74965 = _T_74964[13:0]; // @[Modules.scala 160:64:@21528.4]
  assign buffer_6_365 = $signed(_T_74965); // @[Modules.scala 160:64:@21529.4]
  assign buffer_6_100 = {{8{_T_73311[5]}},_T_73311}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_101 = {{9{_T_73318[4]}},_T_73318}; // @[Modules.scala 112:22:@8.4]
  assign _T_74967 = $signed(buffer_6_100) + $signed(buffer_6_101); // @[Modules.scala 160:64:@21531.4]
  assign _T_74968 = _T_74967[13:0]; // @[Modules.scala 160:64:@21532.4]
  assign buffer_6_366 = $signed(_T_74968); // @[Modules.scala 160:64:@21533.4]
  assign buffer_6_102 = {{8{_T_73325[5]}},_T_73325}; // @[Modules.scala 112:22:@8.4]
  assign _T_74970 = $signed(buffer_6_102) + $signed(buffer_0_100); // @[Modules.scala 160:64:@21535.4]
  assign _T_74971 = _T_74970[13:0]; // @[Modules.scala 160:64:@21536.4]
  assign buffer_6_367 = $signed(_T_74971); // @[Modules.scala 160:64:@21537.4]
  assign buffer_6_105 = {{8{_T_73346[5]}},_T_73346}; // @[Modules.scala 112:22:@8.4]
  assign _T_74973 = $signed(buffer_1_104) + $signed(buffer_6_105); // @[Modules.scala 160:64:@21539.4]
  assign _T_74974 = _T_74973[13:0]; // @[Modules.scala 160:64:@21540.4]
  assign buffer_6_368 = $signed(_T_74974); // @[Modules.scala 160:64:@21541.4]
  assign _T_74976 = $signed(buffer_0_103) + $signed(buffer_0_104); // @[Modules.scala 160:64:@21543.4]
  assign _T_74977 = _T_74976[13:0]; // @[Modules.scala 160:64:@21544.4]
  assign buffer_6_369 = $signed(_T_74977); // @[Modules.scala 160:64:@21545.4]
  assign _T_74979 = $signed(buffer_0_105) + $signed(buffer_0_106); // @[Modules.scala 160:64:@21547.4]
  assign _T_74980 = _T_74979[13:0]; // @[Modules.scala 160:64:@21548.4]
  assign buffer_6_370 = $signed(_T_74980); // @[Modules.scala 160:64:@21549.4]
  assign buffer_6_111 = {{8{_T_73388[5]}},_T_73388}; // @[Modules.scala 112:22:@8.4]
  assign _T_74982 = $signed(buffer_0_107) + $signed(buffer_6_111); // @[Modules.scala 160:64:@21551.4]
  assign _T_74983 = _T_74982[13:0]; // @[Modules.scala 160:64:@21552.4]
  assign buffer_6_371 = $signed(_T_74983); // @[Modules.scala 160:64:@21553.4]
  assign buffer_6_112 = {{8{_T_73395[5]}},_T_73395}; // @[Modules.scala 112:22:@8.4]
  assign _T_74985 = $signed(buffer_6_112) + $signed(buffer_1_112); // @[Modules.scala 160:64:@21555.4]
  assign _T_74986 = _T_74985[13:0]; // @[Modules.scala 160:64:@21556.4]
  assign buffer_6_372 = $signed(_T_74986); // @[Modules.scala 160:64:@21557.4]
  assign buffer_6_114 = {{8{_T_73409[5]}},_T_73409}; // @[Modules.scala 112:22:@8.4]
  assign _T_74988 = $signed(buffer_6_114) + $signed(buffer_1_114); // @[Modules.scala 160:64:@21559.4]
  assign _T_74989 = _T_74988[13:0]; // @[Modules.scala 160:64:@21560.4]
  assign buffer_6_373 = $signed(_T_74989); // @[Modules.scala 160:64:@21561.4]
  assign _T_74991 = $signed(buffer_1_115) + $signed(buffer_1_116); // @[Modules.scala 160:64:@21563.4]
  assign _T_74992 = _T_74991[13:0]; // @[Modules.scala 160:64:@21564.4]
  assign buffer_6_374 = $signed(_T_74992); // @[Modules.scala 160:64:@21565.4]
  assign buffer_6_118 = {{8{_T_73437[5]}},_T_73437}; // @[Modules.scala 112:22:@8.4]
  assign _T_74994 = $signed(buffer_6_118) + $signed(buffer_0_116); // @[Modules.scala 160:64:@21567.4]
  assign _T_74995 = _T_74994[13:0]; // @[Modules.scala 160:64:@21568.4]
  assign buffer_6_375 = $signed(_T_74995); // @[Modules.scala 160:64:@21569.4]
  assign _T_74997 = $signed(buffer_0_117) + $signed(buffer_0_118); // @[Modules.scala 160:64:@21571.4]
  assign _T_74998 = _T_74997[13:0]; // @[Modules.scala 160:64:@21572.4]
  assign buffer_6_376 = $signed(_T_74998); // @[Modules.scala 160:64:@21573.4]
  assign buffer_6_122 = {{8{_T_73465[5]}},_T_73465}; // @[Modules.scala 112:22:@8.4]
  assign _T_75000 = $signed(buffer_6_122) + $signed(buffer_4_118); // @[Modules.scala 160:64:@21575.4]
  assign _T_75001 = _T_75000[13:0]; // @[Modules.scala 160:64:@21576.4]
  assign buffer_6_377 = $signed(_T_75001); // @[Modules.scala 160:64:@21577.4]
  assign _T_75003 = $signed(buffer_2_124) + $signed(buffer_5_124); // @[Modules.scala 160:64:@21579.4]
  assign _T_75004 = _T_75003[13:0]; // @[Modules.scala 160:64:@21580.4]
  assign buffer_6_378 = $signed(_T_75004); // @[Modules.scala 160:64:@21581.4]
  assign _T_75006 = $signed(buffer_5_125) + $signed(buffer_1_125); // @[Modules.scala 160:64:@21583.4]
  assign _T_75007 = _T_75006[13:0]; // @[Modules.scala 160:64:@21584.4]
  assign buffer_6_379 = $signed(_T_75007); // @[Modules.scala 160:64:@21585.4]
  assign buffer_6_128 = {{8{_T_73507[5]}},_T_73507}; // @[Modules.scala 112:22:@8.4]
  assign _T_75009 = $signed(buffer_6_128) + $signed(buffer_0_126); // @[Modules.scala 160:64:@21587.4]
  assign _T_75010 = _T_75009[13:0]; // @[Modules.scala 160:64:@21588.4]
  assign buffer_6_380 = $signed(_T_75010); // @[Modules.scala 160:64:@21589.4]
  assign buffer_6_130 = {{8{_T_73521[5]}},_T_73521}; // @[Modules.scala 112:22:@8.4]
  assign _T_75012 = $signed(buffer_6_130) + $signed(buffer_0_128); // @[Modules.scala 160:64:@21591.4]
  assign _T_75013 = _T_75012[13:0]; // @[Modules.scala 160:64:@21592.4]
  assign buffer_6_381 = $signed(_T_75013); // @[Modules.scala 160:64:@21593.4]
  assign _T_75015 = $signed(buffer_0_129) + $signed(buffer_0_130); // @[Modules.scala 160:64:@21595.4]
  assign _T_75016 = _T_75015[13:0]; // @[Modules.scala 160:64:@21596.4]
  assign buffer_6_382 = $signed(_T_75016); // @[Modules.scala 160:64:@21597.4]
  assign buffer_6_135 = {{8{_T_73556[5]}},_T_73556}; // @[Modules.scala 112:22:@8.4]
  assign _T_75018 = $signed(buffer_0_131) + $signed(buffer_6_135); // @[Modules.scala 160:64:@21599.4]
  assign _T_75019 = _T_75018[13:0]; // @[Modules.scala 160:64:@21600.4]
  assign buffer_6_383 = $signed(_T_75019); // @[Modules.scala 160:64:@21601.4]
  assign buffer_6_136 = {{8{_T_73563[5]}},_T_73563}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_137 = {{8{_T_73570[5]}},_T_73570}; // @[Modules.scala 112:22:@8.4]
  assign _T_75021 = $signed(buffer_6_136) + $signed(buffer_6_137); // @[Modules.scala 160:64:@21603.4]
  assign _T_75022 = _T_75021[13:0]; // @[Modules.scala 160:64:@21604.4]
  assign buffer_6_384 = $signed(_T_75022); // @[Modules.scala 160:64:@21605.4]
  assign buffer_6_140 = {{8{_T_73591[5]}},_T_73591}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_141 = {{8{_T_73598[5]}},_T_73598}; // @[Modules.scala 112:22:@8.4]
  assign _T_75027 = $signed(buffer_6_140) + $signed(buffer_6_141); // @[Modules.scala 160:64:@21611.4]
  assign _T_75028 = _T_75027[13:0]; // @[Modules.scala 160:64:@21612.4]
  assign buffer_6_386 = $signed(_T_75028); // @[Modules.scala 160:64:@21613.4]
  assign buffer_6_144 = {{8{_T_73619[5]}},_T_73619}; // @[Modules.scala 112:22:@8.4]
  assign _T_75033 = $signed(buffer_6_144) + $signed(buffer_0_141); // @[Modules.scala 160:64:@21619.4]
  assign _T_75034 = _T_75033[13:0]; // @[Modules.scala 160:64:@21620.4]
  assign buffer_6_388 = $signed(_T_75034); // @[Modules.scala 160:64:@21621.4]
  assign buffer_6_149 = {{9{_T_73654[4]}},_T_73654}; // @[Modules.scala 112:22:@8.4]
  assign _T_75039 = $signed(buffer_0_144) + $signed(buffer_6_149); // @[Modules.scala 160:64:@21627.4]
  assign _T_75040 = _T_75039[13:0]; // @[Modules.scala 160:64:@21628.4]
  assign buffer_6_390 = $signed(_T_75040); // @[Modules.scala 160:64:@21629.4]
  assign buffer_6_151 = {{9{_T_73668[4]}},_T_73668}; // @[Modules.scala 112:22:@8.4]
  assign _T_75042 = $signed(buffer_2_149) + $signed(buffer_6_151); // @[Modules.scala 160:64:@21631.4]
  assign _T_75043 = _T_75042[13:0]; // @[Modules.scala 160:64:@21632.4]
  assign buffer_6_391 = $signed(_T_75043); // @[Modules.scala 160:64:@21633.4]
  assign _T_75045 = $signed(buffer_1_149) + $signed(buffer_1_150); // @[Modules.scala 160:64:@21635.4]
  assign _T_75046 = _T_75045[13:0]; // @[Modules.scala 160:64:@21636.4]
  assign buffer_6_392 = $signed(_T_75046); // @[Modules.scala 160:64:@21637.4]
  assign _T_75048 = $signed(buffer_1_151) + $signed(buffer_1_152); // @[Modules.scala 160:64:@21639.4]
  assign _T_75049 = _T_75048[13:0]; // @[Modules.scala 160:64:@21640.4]
  assign buffer_6_393 = $signed(_T_75049); // @[Modules.scala 160:64:@21641.4]
  assign _T_75051 = $signed(buffer_2_155) + $signed(buffer_2_156); // @[Modules.scala 160:64:@21643.4]
  assign _T_75052 = _T_75051[13:0]; // @[Modules.scala 160:64:@21644.4]
  assign buffer_6_394 = $signed(_T_75052); // @[Modules.scala 160:64:@21645.4]
  assign _T_75054 = $signed(buffer_5_153) + $signed(buffer_5_154); // @[Modules.scala 160:64:@21647.4]
  assign _T_75055 = _T_75054[13:0]; // @[Modules.scala 160:64:@21648.4]
  assign buffer_6_395 = $signed(_T_75055); // @[Modules.scala 160:64:@21649.4]
  assign _T_75057 = $signed(buffer_5_155) + $signed(buffer_1_156); // @[Modules.scala 160:64:@21651.4]
  assign _T_75058 = _T_75057[13:0]; // @[Modules.scala 160:64:@21652.4]
  assign buffer_6_396 = $signed(_T_75058); // @[Modules.scala 160:64:@21653.4]
  assign _T_75060 = $signed(buffer_5_157) + $signed(buffer_2_162); // @[Modules.scala 160:64:@21655.4]
  assign _T_75061 = _T_75060[13:0]; // @[Modules.scala 160:64:@21656.4]
  assign buffer_6_397 = $signed(_T_75061); // @[Modules.scala 160:64:@21657.4]
  assign buffer_6_165 = {{9{_T_73766[4]}},_T_73766}; // @[Modules.scala 112:22:@8.4]
  assign _T_75063 = $signed(buffer_4_155) + $signed(buffer_6_165); // @[Modules.scala 160:64:@21659.4]
  assign _T_75064 = _T_75063[13:0]; // @[Modules.scala 160:64:@21660.4]
  assign buffer_6_398 = $signed(_T_75064); // @[Modules.scala 160:64:@21661.4]
  assign _T_75066 = $signed(buffer_5_161) + $signed(buffer_5_162); // @[Modules.scala 160:64:@21663.4]
  assign _T_75067 = _T_75066[13:0]; // @[Modules.scala 160:64:@21664.4]
  assign buffer_6_399 = $signed(_T_75067); // @[Modules.scala 160:64:@21665.4]
  assign buffer_6_169 = {{8{_T_73794[5]}},_T_73794}; // @[Modules.scala 112:22:@8.4]
  assign _T_75069 = $signed(buffer_5_163) + $signed(buffer_6_169); // @[Modules.scala 160:64:@21667.4]
  assign _T_75070 = _T_75069[13:0]; // @[Modules.scala 160:64:@21668.4]
  assign buffer_6_400 = $signed(_T_75070); // @[Modules.scala 160:64:@21669.4]
  assign buffer_6_171 = {{8{_T_73808[5]}},_T_73808}; // @[Modules.scala 112:22:@8.4]
  assign _T_75072 = $signed(buffer_2_168) + $signed(buffer_6_171); // @[Modules.scala 160:64:@21671.4]
  assign _T_75073 = _T_75072[13:0]; // @[Modules.scala 160:64:@21672.4]
  assign buffer_6_401 = $signed(_T_75073); // @[Modules.scala 160:64:@21673.4]
  assign _T_75075 = $signed(buffer_5_167) + $signed(buffer_1_167); // @[Modules.scala 160:64:@21675.4]
  assign _T_75076 = _T_75075[13:0]; // @[Modules.scala 160:64:@21676.4]
  assign buffer_6_402 = $signed(_T_75076); // @[Modules.scala 160:64:@21677.4]
  assign buffer_6_175 = {{8{_T_73836[5]}},_T_73836}; // @[Modules.scala 112:22:@8.4]
  assign _T_75078 = $signed(buffer_2_173) + $signed(buffer_6_175); // @[Modules.scala 160:64:@21679.4]
  assign _T_75079 = _T_75078[13:0]; // @[Modules.scala 160:64:@21680.4]
  assign buffer_6_403 = $signed(_T_75079); // @[Modules.scala 160:64:@21681.4]
  assign buffer_6_177 = {{9{_T_73850[4]}},_T_73850}; // @[Modules.scala 112:22:@8.4]
  assign _T_75081 = $signed(buffer_0_170) + $signed(buffer_6_177); // @[Modules.scala 160:64:@21683.4]
  assign _T_75082 = _T_75081[13:0]; // @[Modules.scala 160:64:@21684.4]
  assign buffer_6_404 = $signed(_T_75082); // @[Modules.scala 160:64:@21685.4]
  assign buffer_6_178 = {{8{_T_73857[5]}},_T_73857}; // @[Modules.scala 112:22:@8.4]
  assign _T_75084 = $signed(buffer_6_178) + $signed(buffer_0_173); // @[Modules.scala 160:64:@21687.4]
  assign _T_75085 = _T_75084[13:0]; // @[Modules.scala 160:64:@21688.4]
  assign buffer_6_405 = $signed(_T_75085); // @[Modules.scala 160:64:@21689.4]
  assign buffer_6_180 = {{8{_T_73871[5]}},_T_73871}; // @[Modules.scala 112:22:@8.4]
  assign _T_75087 = $signed(buffer_6_180) + $signed(buffer_1_175); // @[Modules.scala 160:64:@21691.4]
  assign _T_75088 = _T_75087[13:0]; // @[Modules.scala 160:64:@21692.4]
  assign buffer_6_406 = $signed(_T_75088); // @[Modules.scala 160:64:@21693.4]
  assign buffer_6_183 = {{8{_T_73892[5]}},_T_73892}; // @[Modules.scala 112:22:@8.4]
  assign _T_75090 = $signed(buffer_1_176) + $signed(buffer_6_183); // @[Modules.scala 160:64:@21695.4]
  assign _T_75091 = _T_75090[13:0]; // @[Modules.scala 160:64:@21696.4]
  assign buffer_6_407 = $signed(_T_75091); // @[Modules.scala 160:64:@21697.4]
  assign buffer_6_185 = {{8{_T_73906[5]}},_T_73906}; // @[Modules.scala 112:22:@8.4]
  assign _T_75093 = $signed(buffer_4_172) + $signed(buffer_6_185); // @[Modules.scala 160:64:@21699.4]
  assign _T_75094 = _T_75093[13:0]; // @[Modules.scala 160:64:@21700.4]
  assign buffer_6_408 = $signed(_T_75094); // @[Modules.scala 160:64:@21701.4]
  assign _T_75096 = $signed(buffer_2_185) + $signed(buffer_1_181); // @[Modules.scala 160:64:@21703.4]
  assign _T_75097 = _T_75096[13:0]; // @[Modules.scala 160:64:@21704.4]
  assign buffer_6_409 = $signed(_T_75097); // @[Modules.scala 160:64:@21705.4]
  assign buffer_6_188 = {{8{_T_73927[5]}},_T_73927}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_189 = {{8{_T_73934[5]}},_T_73934}; // @[Modules.scala 112:22:@8.4]
  assign _T_75099 = $signed(buffer_6_188) + $signed(buffer_6_189); // @[Modules.scala 160:64:@21707.4]
  assign _T_75100 = _T_75099[13:0]; // @[Modules.scala 160:64:@21708.4]
  assign buffer_6_410 = $signed(_T_75100); // @[Modules.scala 160:64:@21709.4]
  assign buffer_6_190 = {{8{_T_73941[5]}},_T_73941}; // @[Modules.scala 112:22:@8.4]
  assign _T_75102 = $signed(buffer_6_190) + $signed(buffer_0_183); // @[Modules.scala 160:64:@21711.4]
  assign _T_75103 = _T_75102[13:0]; // @[Modules.scala 160:64:@21712.4]
  assign buffer_6_411 = $signed(_T_75103); // @[Modules.scala 160:64:@21713.4]
  assign buffer_6_192 = {{8{_T_73955[5]}},_T_73955}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_193 = {{8{_T_73962[5]}},_T_73962}; // @[Modules.scala 112:22:@8.4]
  assign _T_75105 = $signed(buffer_6_192) + $signed(buffer_6_193); // @[Modules.scala 160:64:@21715.4]
  assign _T_75106 = _T_75105[13:0]; // @[Modules.scala 160:64:@21716.4]
  assign buffer_6_412 = $signed(_T_75106); // @[Modules.scala 160:64:@21717.4]
  assign buffer_6_194 = {{8{_T_73969[5]}},_T_73969}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_195 = {{8{_T_73976[5]}},_T_73976}; // @[Modules.scala 112:22:@8.4]
  assign _T_75108 = $signed(buffer_6_194) + $signed(buffer_6_195); // @[Modules.scala 160:64:@21719.4]
  assign _T_75109 = _T_75108[13:0]; // @[Modules.scala 160:64:@21720.4]
  assign buffer_6_413 = $signed(_T_75109); // @[Modules.scala 160:64:@21721.4]
  assign _T_75111 = $signed(buffer_1_189) + $signed(buffer_1_190); // @[Modules.scala 160:64:@21723.4]
  assign _T_75112 = _T_75111[13:0]; // @[Modules.scala 160:64:@21724.4]
  assign buffer_6_414 = $signed(_T_75112); // @[Modules.scala 160:64:@21725.4]
  assign buffer_6_198 = {{8{_T_73997[5]}},_T_73997}; // @[Modules.scala 112:22:@8.4]
  assign _T_75114 = $signed(buffer_6_198) + $signed(buffer_2_196); // @[Modules.scala 160:64:@21727.4]
  assign _T_75115 = _T_75114[13:0]; // @[Modules.scala 160:64:@21728.4]
  assign buffer_6_415 = $signed(_T_75115); // @[Modules.scala 160:64:@21729.4]
  assign buffer_6_200 = {{8{_T_74011[5]}},_T_74011}; // @[Modules.scala 112:22:@8.4]
  assign _T_75117 = $signed(buffer_6_200) + $signed(buffer_4_184); // @[Modules.scala 160:64:@21731.4]
  assign _T_75118 = _T_75117[13:0]; // @[Modules.scala 160:64:@21732.4]
  assign buffer_6_416 = $signed(_T_75118); // @[Modules.scala 160:64:@21733.4]
  assign buffer_6_202 = {{8{_T_74025[5]}},_T_74025}; // @[Modules.scala 112:22:@8.4]
  assign _T_75120 = $signed(buffer_6_202) + $signed(buffer_0_192); // @[Modules.scala 160:64:@21735.4]
  assign _T_75121 = _T_75120[13:0]; // @[Modules.scala 160:64:@21736.4]
  assign buffer_6_417 = $signed(_T_75121); // @[Modules.scala 160:64:@21737.4]
  assign _T_75123 = $signed(buffer_0_193) + $signed(buffer_4_188); // @[Modules.scala 160:64:@21739.4]
  assign _T_75124 = _T_75123[13:0]; // @[Modules.scala 160:64:@21740.4]
  assign buffer_6_418 = $signed(_T_75124); // @[Modules.scala 160:64:@21741.4]
  assign _T_75126 = $signed(buffer_0_195) + $signed(buffer_0_196); // @[Modules.scala 160:64:@21743.4]
  assign _T_75127 = _T_75126[13:0]; // @[Modules.scala 160:64:@21744.4]
  assign buffer_6_419 = $signed(_T_75127); // @[Modules.scala 160:64:@21745.4]
  assign _T_75129 = $signed(buffer_0_197) + $signed(buffer_4_192); // @[Modules.scala 160:64:@21747.4]
  assign _T_75130 = _T_75129[13:0]; // @[Modules.scala 160:64:@21748.4]
  assign buffer_6_420 = $signed(_T_75130); // @[Modules.scala 160:64:@21749.4]
  assign buffer_6_211 = {{8{_T_74088[5]}},_T_74088}; // @[Modules.scala 112:22:@8.4]
  assign _T_75132 = $signed(buffer_4_193) + $signed(buffer_6_211); // @[Modules.scala 160:64:@21751.4]
  assign _T_75133 = _T_75132[13:0]; // @[Modules.scala 160:64:@21752.4]
  assign buffer_6_421 = $signed(_T_75133); // @[Modules.scala 160:64:@21753.4]
  assign buffer_6_212 = {{8{_T_74095[5]}},_T_74095}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_213 = {{8{_T_74102[5]}},_T_74102}; // @[Modules.scala 112:22:@8.4]
  assign _T_75135 = $signed(buffer_6_212) + $signed(buffer_6_213); // @[Modules.scala 160:64:@21755.4]
  assign _T_75136 = _T_75135[13:0]; // @[Modules.scala 160:64:@21756.4]
  assign buffer_6_422 = $signed(_T_75136); // @[Modules.scala 160:64:@21757.4]
  assign buffer_6_220 = {{8{_T_74151[5]}},_T_74151}; // @[Modules.scala 112:22:@8.4]
  assign _T_75147 = $signed(buffer_6_220) + $signed(buffer_4_203); // @[Modules.scala 160:64:@21771.4]
  assign _T_75148 = _T_75147[13:0]; // @[Modules.scala 160:64:@21772.4]
  assign buffer_6_426 = $signed(_T_75148); // @[Modules.scala 160:64:@21773.4]
  assign buffer_6_223 = {{8{_T_74172[5]}},_T_74172}; // @[Modules.scala 112:22:@8.4]
  assign _T_75150 = $signed(buffer_5_215) + $signed(buffer_6_223); // @[Modules.scala 160:64:@21775.4]
  assign _T_75151 = _T_75150[13:0]; // @[Modules.scala 160:64:@21776.4]
  assign buffer_6_427 = $signed(_T_75151); // @[Modules.scala 160:64:@21777.4]
  assign buffer_6_224 = {{8{_T_74179[5]}},_T_74179}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_225 = {{8{_T_74186[5]}},_T_74186}; // @[Modules.scala 112:22:@8.4]
  assign _T_75153 = $signed(buffer_6_224) + $signed(buffer_6_225); // @[Modules.scala 160:64:@21779.4]
  assign _T_75154 = _T_75153[13:0]; // @[Modules.scala 160:64:@21780.4]
  assign buffer_6_428 = $signed(_T_75154); // @[Modules.scala 160:64:@21781.4]
  assign buffer_6_226 = {{9{_T_74193[4]}},_T_74193}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_227 = {{8{_T_74200[5]}},_T_74200}; // @[Modules.scala 112:22:@8.4]
  assign _T_75156 = $signed(buffer_6_226) + $signed(buffer_6_227); // @[Modules.scala 160:64:@21783.4]
  assign _T_75157 = _T_75156[13:0]; // @[Modules.scala 160:64:@21784.4]
  assign buffer_6_429 = $signed(_T_75157); // @[Modules.scala 160:64:@21785.4]
  assign buffer_6_228 = {{8{_T_74207[5]}},_T_74207}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_229 = {{8{_T_74214[5]}},_T_74214}; // @[Modules.scala 112:22:@8.4]
  assign _T_75159 = $signed(buffer_6_228) + $signed(buffer_6_229); // @[Modules.scala 160:64:@21787.4]
  assign _T_75160 = _T_75159[13:0]; // @[Modules.scala 160:64:@21788.4]
  assign buffer_6_430 = $signed(_T_75160); // @[Modules.scala 160:64:@21789.4]
  assign buffer_6_230 = {{8{_T_74221[5]}},_T_74221}; // @[Modules.scala 112:22:@8.4]
  assign _T_75162 = $signed(buffer_6_230) + $signed(buffer_0_219); // @[Modules.scala 160:64:@21791.4]
  assign _T_75163 = _T_75162[13:0]; // @[Modules.scala 160:64:@21792.4]
  assign buffer_6_431 = $signed(_T_75163); // @[Modules.scala 160:64:@21793.4]
  assign buffer_6_233 = {{8{_T_74242[5]}},_T_74242}; // @[Modules.scala 112:22:@8.4]
  assign _T_75165 = $signed(buffer_0_220) + $signed(buffer_6_233); // @[Modules.scala 160:64:@21795.4]
  assign _T_75166 = _T_75165[13:0]; // @[Modules.scala 160:64:@21796.4]
  assign buffer_6_432 = $signed(_T_75166); // @[Modules.scala 160:64:@21797.4]
  assign _T_75168 = $signed(buffer_3_233) + $signed(buffer_3_234); // @[Modules.scala 160:64:@21799.4]
  assign _T_75169 = _T_75168[13:0]; // @[Modules.scala 160:64:@21800.4]
  assign buffer_6_433 = $signed(_T_75169); // @[Modules.scala 160:64:@21801.4]
  assign buffer_6_236 = {{8{_T_74263[5]}},_T_74263}; // @[Modules.scala 112:22:@8.4]
  assign _T_75171 = $signed(buffer_6_236) + $signed(buffer_5_230); // @[Modules.scala 160:64:@21803.4]
  assign _T_75172 = _T_75171[13:0]; // @[Modules.scala 160:64:@21804.4]
  assign buffer_6_434 = $signed(_T_75172); // @[Modules.scala 160:64:@21805.4]
  assign _T_75174 = $signed(buffer_1_226) + $signed(buffer_0_226); // @[Modules.scala 160:64:@21807.4]
  assign _T_75175 = _T_75174[13:0]; // @[Modules.scala 160:64:@21808.4]
  assign buffer_6_435 = $signed(_T_75175); // @[Modules.scala 160:64:@21809.4]
  assign buffer_6_240 = {{8{_T_74291[5]}},_T_74291}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_241 = {{8{_T_74298[5]}},_T_74298}; // @[Modules.scala 112:22:@8.4]
  assign _T_75177 = $signed(buffer_6_240) + $signed(buffer_6_241); // @[Modules.scala 160:64:@21811.4]
  assign _T_75178 = _T_75177[13:0]; // @[Modules.scala 160:64:@21812.4]
  assign buffer_6_436 = $signed(_T_75178); // @[Modules.scala 160:64:@21813.4]
  assign buffer_6_243 = {{8{_T_74312[5]}},_T_74312}; // @[Modules.scala 112:22:@8.4]
  assign _T_75180 = $signed(buffer_0_229) + $signed(buffer_6_243); // @[Modules.scala 160:64:@21815.4]
  assign _T_75181 = _T_75180[13:0]; // @[Modules.scala 160:64:@21816.4]
  assign buffer_6_437 = $signed(_T_75181); // @[Modules.scala 160:64:@21817.4]
  assign buffer_6_244 = {{9{_T_74319[4]}},_T_74319}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_245 = {{8{_T_74326[5]}},_T_74326}; // @[Modules.scala 112:22:@8.4]
  assign _T_75183 = $signed(buffer_6_244) + $signed(buffer_6_245); // @[Modules.scala 160:64:@21819.4]
  assign _T_75184 = _T_75183[13:0]; // @[Modules.scala 160:64:@21820.4]
  assign buffer_6_438 = $signed(_T_75184); // @[Modules.scala 160:64:@21821.4]
  assign buffer_6_246 = {{8{_T_74333[5]}},_T_74333}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_247 = {{8{_T_74340[5]}},_T_74340}; // @[Modules.scala 112:22:@8.4]
  assign _T_75186 = $signed(buffer_6_246) + $signed(buffer_6_247); // @[Modules.scala 160:64:@21823.4]
  assign _T_75187 = _T_75186[13:0]; // @[Modules.scala 160:64:@21824.4]
  assign buffer_6_439 = $signed(_T_75187); // @[Modules.scala 160:64:@21825.4]
  assign buffer_6_248 = {{8{_T_74347[5]}},_T_74347}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_249 = {{8{_T_74354[5]}},_T_74354}; // @[Modules.scala 112:22:@8.4]
  assign _T_75189 = $signed(buffer_6_248) + $signed(buffer_6_249); // @[Modules.scala 160:64:@21827.4]
  assign _T_75190 = _T_75189[13:0]; // @[Modules.scala 160:64:@21828.4]
  assign buffer_6_440 = $signed(_T_75190); // @[Modules.scala 160:64:@21829.4]
  assign buffer_6_250 = {{9{_T_74361[4]}},_T_74361}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_251 = {{8{_T_74368[5]}},_T_74368}; // @[Modules.scala 112:22:@8.4]
  assign _T_75192 = $signed(buffer_6_250) + $signed(buffer_6_251); // @[Modules.scala 160:64:@21831.4]
  assign _T_75193 = _T_75192[13:0]; // @[Modules.scala 160:64:@21832.4]
  assign buffer_6_441 = $signed(_T_75193); // @[Modules.scala 160:64:@21833.4]
  assign buffer_6_252 = {{8{_T_74375[5]}},_T_74375}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_253 = {{8{_T_74382[5]}},_T_74382}; // @[Modules.scala 112:22:@8.4]
  assign _T_75195 = $signed(buffer_6_252) + $signed(buffer_6_253); // @[Modules.scala 160:64:@21835.4]
  assign _T_75196 = _T_75195[13:0]; // @[Modules.scala 160:64:@21836.4]
  assign buffer_6_442 = $signed(_T_75196); // @[Modules.scala 160:64:@21837.4]
  assign _T_75198 = $signed(buffer_1_244) + $signed(buffer_0_243); // @[Modules.scala 160:64:@21839.4]
  assign _T_75199 = _T_75198[13:0]; // @[Modules.scala 160:64:@21840.4]
  assign buffer_6_443 = $signed(_T_75199); // @[Modules.scala 160:64:@21841.4]
  assign buffer_6_257 = {{8{_T_74410[5]}},_T_74410}; // @[Modules.scala 112:22:@8.4]
  assign _T_75201 = $signed(buffer_0_244) + $signed(buffer_6_257); // @[Modules.scala 160:64:@21843.4]
  assign _T_75202 = _T_75201[13:0]; // @[Modules.scala 160:64:@21844.4]
  assign buffer_6_444 = $signed(_T_75202); // @[Modules.scala 160:64:@21845.4]
  assign buffer_6_258 = {{8{_T_74417[5]}},_T_74417}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_259 = {{8{_T_74424[5]}},_T_74424}; // @[Modules.scala 112:22:@8.4]
  assign _T_75204 = $signed(buffer_6_258) + $signed(buffer_6_259); // @[Modules.scala 160:64:@21847.4]
  assign _T_75205 = _T_75204[13:0]; // @[Modules.scala 160:64:@21848.4]
  assign buffer_6_445 = $signed(_T_75205); // @[Modules.scala 160:64:@21849.4]
  assign buffer_6_260 = {{8{_T_74431[5]}},_T_74431}; // @[Modules.scala 112:22:@8.4]
  assign _T_75207 = $signed(buffer_6_260) + $signed(buffer_1_250); // @[Modules.scala 160:64:@21851.4]
  assign _T_75208 = _T_75207[13:0]; // @[Modules.scala 160:64:@21852.4]
  assign buffer_6_446 = $signed(_T_75208); // @[Modules.scala 160:64:@21853.4]
  assign buffer_6_263 = {{8{_T_74452[5]}},_T_74452}; // @[Modules.scala 112:22:@8.4]
  assign _T_75210 = $signed(buffer_5_259) + $signed(buffer_6_263); // @[Modules.scala 160:64:@21855.4]
  assign _T_75211 = _T_75210[13:0]; // @[Modules.scala 160:64:@21856.4]
  assign buffer_6_447 = $signed(_T_75211); // @[Modules.scala 160:64:@21857.4]
  assign buffer_6_264 = {{8{_T_74459[5]}},_T_74459}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_265 = {{9{_T_74466[4]}},_T_74466}; // @[Modules.scala 112:22:@8.4]
  assign _T_75213 = $signed(buffer_6_264) + $signed(buffer_6_265); // @[Modules.scala 160:64:@21859.4]
  assign _T_75214 = _T_75213[13:0]; // @[Modules.scala 160:64:@21860.4]
  assign buffer_6_448 = $signed(_T_75214); // @[Modules.scala 160:64:@21861.4]
  assign buffer_6_268 = {{9{_T_74487[4]}},_T_74487}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_269 = {{9{_T_74494[4]}},_T_74494}; // @[Modules.scala 112:22:@8.4]
  assign _T_75219 = $signed(buffer_6_268) + $signed(buffer_6_269); // @[Modules.scala 160:64:@21867.4]
  assign _T_75220 = _T_75219[13:0]; // @[Modules.scala 160:64:@21868.4]
  assign buffer_6_450 = $signed(_T_75220); // @[Modules.scala 160:64:@21869.4]
  assign buffer_6_270 = {{8{_T_74501[5]}},_T_74501}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_271 = {{8{_T_74508[5]}},_T_74508}; // @[Modules.scala 112:22:@8.4]
  assign _T_75222 = $signed(buffer_6_270) + $signed(buffer_6_271); // @[Modules.scala 160:64:@21871.4]
  assign _T_75223 = _T_75222[13:0]; // @[Modules.scala 160:64:@21872.4]
  assign buffer_6_451 = $signed(_T_75223); // @[Modules.scala 160:64:@21873.4]
  assign buffer_6_272 = {{8{_T_74515[5]}},_T_74515}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_273 = {{8{_T_74522[5]}},_T_74522}; // @[Modules.scala 112:22:@8.4]
  assign _T_75225 = $signed(buffer_6_272) + $signed(buffer_6_273); // @[Modules.scala 160:64:@21875.4]
  assign _T_75226 = _T_75225[13:0]; // @[Modules.scala 160:64:@21876.4]
  assign buffer_6_452 = $signed(_T_75226); // @[Modules.scala 160:64:@21877.4]
  assign buffer_6_274 = {{8{_T_74529[5]}},_T_74529}; // @[Modules.scala 112:22:@8.4]
  assign _T_75228 = $signed(buffer_6_274) + $signed(buffer_2_272); // @[Modules.scala 160:64:@21879.4]
  assign _T_75229 = _T_75228[13:0]; // @[Modules.scala 160:64:@21880.4]
  assign buffer_6_453 = $signed(_T_75229); // @[Modules.scala 160:64:@21881.4]
  assign _T_75231 = $signed(buffer_2_273) + $signed(buffer_3_276); // @[Modules.scala 160:64:@21883.4]
  assign _T_75232 = _T_75231[13:0]; // @[Modules.scala 160:64:@21884.4]
  assign buffer_6_454 = $signed(_T_75232); // @[Modules.scala 160:64:@21885.4]
  assign buffer_6_278 = {{9{_T_74557[4]}},_T_74557}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_279 = {{9{_T_74564[4]}},_T_74564}; // @[Modules.scala 112:22:@8.4]
  assign _T_75234 = $signed(buffer_6_278) + $signed(buffer_6_279); // @[Modules.scala 160:64:@21887.4]
  assign _T_75235 = _T_75234[13:0]; // @[Modules.scala 160:64:@21888.4]
  assign buffer_6_455 = $signed(_T_75235); // @[Modules.scala 160:64:@21889.4]
  assign buffer_6_280 = {{9{_T_74571[4]}},_T_74571}; // @[Modules.scala 112:22:@8.4]
  assign _T_75237 = $signed(buffer_6_280) + $signed(buffer_1_270); // @[Modules.scala 160:64:@21891.4]
  assign _T_75238 = _T_75237[13:0]; // @[Modules.scala 160:64:@21892.4]
  assign buffer_6_456 = $signed(_T_75238); // @[Modules.scala 160:64:@21893.4]
  assign buffer_6_282 = {{8{_T_74585[5]}},_T_74585}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_283 = {{8{_T_74592[5]}},_T_74592}; // @[Modules.scala 112:22:@8.4]
  assign _T_75240 = $signed(buffer_6_282) + $signed(buffer_6_283); // @[Modules.scala 160:64:@21895.4]
  assign _T_75241 = _T_75240[13:0]; // @[Modules.scala 160:64:@21896.4]
  assign buffer_6_457 = $signed(_T_75241); // @[Modules.scala 160:64:@21897.4]
  assign buffer_6_284 = {{8{_T_74599[5]}},_T_74599}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_285 = {{8{_T_74606[5]}},_T_74606}; // @[Modules.scala 112:22:@8.4]
  assign _T_75243 = $signed(buffer_6_284) + $signed(buffer_6_285); // @[Modules.scala 160:64:@21899.4]
  assign _T_75244 = _T_75243[13:0]; // @[Modules.scala 160:64:@21900.4]
  assign buffer_6_458 = $signed(_T_75244); // @[Modules.scala 160:64:@21901.4]
  assign buffer_6_286 = {{8{_T_74613[5]}},_T_74613}; // @[Modules.scala 112:22:@8.4]
  assign _T_75246 = $signed(buffer_6_286) + $signed(buffer_0_276); // @[Modules.scala 160:64:@21903.4]
  assign _T_75247 = _T_75246[13:0]; // @[Modules.scala 160:64:@21904.4]
  assign buffer_6_459 = $signed(_T_75247); // @[Modules.scala 160:64:@21905.4]
  assign buffer_6_289 = {{8{_T_74634[5]}},_T_74634}; // @[Modules.scala 112:22:@8.4]
  assign _T_75249 = $signed(buffer_0_277) + $signed(buffer_6_289); // @[Modules.scala 160:64:@21907.4]
  assign _T_75250 = _T_75249[13:0]; // @[Modules.scala 160:64:@21908.4]
  assign buffer_6_460 = $signed(_T_75250); // @[Modules.scala 160:64:@21909.4]
  assign buffer_6_291 = {{9{_T_74648[4]}},_T_74648}; // @[Modules.scala 112:22:@8.4]
  assign _T_75252 = $signed(buffer_0_279) + $signed(buffer_6_291); // @[Modules.scala 160:64:@21911.4]
  assign _T_75253 = _T_75252[13:0]; // @[Modules.scala 160:64:@21912.4]
  assign buffer_6_461 = $signed(_T_75253); // @[Modules.scala 160:64:@21913.4]
  assign buffer_6_292 = {{9{_T_74655[4]}},_T_74655}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_293 = {{9{_T_74662[4]}},_T_74662}; // @[Modules.scala 112:22:@8.4]
  assign _T_75255 = $signed(buffer_6_292) + $signed(buffer_6_293); // @[Modules.scala 160:64:@21915.4]
  assign _T_75256 = _T_75255[13:0]; // @[Modules.scala 160:64:@21916.4]
  assign buffer_6_462 = $signed(_T_75256); // @[Modules.scala 160:64:@21917.4]
  assign buffer_6_294 = {{8{_T_74669[5]}},_T_74669}; // @[Modules.scala 112:22:@8.4]
  assign buffer_6_295 = {{8{_T_74676[5]}},_T_74676}; // @[Modules.scala 112:22:@8.4]
  assign _T_75258 = $signed(buffer_6_294) + $signed(buffer_6_295); // @[Modules.scala 160:64:@21919.4]
  assign _T_75259 = _T_75258[13:0]; // @[Modules.scala 160:64:@21920.4]
  assign buffer_6_463 = $signed(_T_75259); // @[Modules.scala 160:64:@21921.4]
  assign buffer_6_296 = {{8{_T_74683[5]}},_T_74683}; // @[Modules.scala 112:22:@8.4]
  assign _T_75261 = $signed(buffer_6_296) + $signed(buffer_4_281); // @[Modules.scala 160:64:@21923.4]
  assign _T_75262 = _T_75261[13:0]; // @[Modules.scala 160:64:@21924.4]
  assign buffer_6_464 = $signed(_T_75262); // @[Modules.scala 160:64:@21925.4]
  assign buffer_6_303 = {{8{_T_74732[5]}},_T_74732}; // @[Modules.scala 112:22:@8.4]
  assign _T_75270 = $signed(buffer_4_286) + $signed(buffer_6_303); // @[Modules.scala 160:64:@21935.4]
  assign _T_75271 = _T_75270[13:0]; // @[Modules.scala 160:64:@21936.4]
  assign buffer_6_467 = $signed(_T_75271); // @[Modules.scala 160:64:@21937.4]
  assign buffer_6_304 = {{9{_T_74739[4]}},_T_74739}; // @[Modules.scala 112:22:@8.4]
  assign _T_75273 = $signed(buffer_6_304) + $signed(buffer_4_289); // @[Modules.scala 160:64:@21939.4]
  assign _T_75274 = _T_75273[13:0]; // @[Modules.scala 160:64:@21940.4]
  assign buffer_6_468 = $signed(_T_75274); // @[Modules.scala 160:64:@21941.4]
  assign _T_75276 = $signed(buffer_3_303) + $signed(buffer_0_293); // @[Modules.scala 160:64:@21943.4]
  assign _T_75277 = _T_75276[13:0]; // @[Modules.scala 160:64:@21944.4]
  assign buffer_6_469 = $signed(_T_75277); // @[Modules.scala 160:64:@21945.4]
  assign _T_75279 = $signed(buffer_4_292) + $signed(buffer_5_306); // @[Modules.scala 160:64:@21947.4]
  assign _T_75280 = _T_75279[13:0]; // @[Modules.scala 160:64:@21948.4]
  assign buffer_6_470 = $signed(_T_75280); // @[Modules.scala 160:64:@21949.4]
  assign _T_75282 = $signed(buffer_5_307) + $signed(buffer_5_308); // @[Modules.scala 160:64:@21951.4]
  assign _T_75283 = _T_75282[13:0]; // @[Modules.scala 160:64:@21952.4]
  assign buffer_6_471 = $signed(_T_75283); // @[Modules.scala 160:64:@21953.4]
  assign _T_75285 = $signed(buffer_0_297) + $signed(buffer_0_298); // @[Modules.scala 160:64:@21955.4]
  assign _T_75286 = _T_75285[13:0]; // @[Modules.scala 160:64:@21956.4]
  assign buffer_6_472 = $signed(_T_75286); // @[Modules.scala 160:64:@21957.4]
  assign buffer_6_315 = {{8{_T_74816[5]}},_T_74816}; // @[Modules.scala 112:22:@8.4]
  assign _T_75288 = $signed(buffer_5_311) + $signed(buffer_6_315); // @[Modules.scala 160:64:@21959.4]
  assign _T_75289 = _T_75288[13:0]; // @[Modules.scala 160:64:@21960.4]
  assign buffer_6_473 = $signed(_T_75289); // @[Modules.scala 160:64:@21961.4]
  assign _T_75291 = $signed(buffer_0_302) + $signed(buffer_6_317); // @[Modules.scala 160:64:@21963.4]
  assign _T_75292 = _T_75291[13:0]; // @[Modules.scala 160:64:@21964.4]
  assign buffer_6_474 = $signed(_T_75292); // @[Modules.scala 160:64:@21965.4]
  assign _T_75294 = $signed(buffer_6_318) + $signed(buffer_4_302); // @[Modules.scala 160:64:@21967.4]
  assign _T_75295 = _T_75294[13:0]; // @[Modules.scala 160:64:@21968.4]
  assign buffer_6_475 = $signed(_T_75295); // @[Modules.scala 160:64:@21969.4]
  assign _T_75297 = $signed(buffer_6_320) + $signed(buffer_6_321); // @[Modules.scala 160:64:@21971.4]
  assign _T_75298 = _T_75297[13:0]; // @[Modules.scala 160:64:@21972.4]
  assign buffer_6_476 = $signed(_T_75298); // @[Modules.scala 160:64:@21973.4]
  assign _T_75300 = $signed(buffer_6_322) + $signed(buffer_4_306); // @[Modules.scala 160:64:@21975.4]
  assign _T_75301 = _T_75300[13:0]; // @[Modules.scala 160:64:@21976.4]
  assign buffer_6_477 = $signed(_T_75301); // @[Modules.scala 160:64:@21977.4]
  assign _T_75306 = $signed(buffer_6_326) + $signed(buffer_6_327); // @[Modules.scala 160:64:@21983.4]
  assign _T_75307 = _T_75306[13:0]; // @[Modules.scala 160:64:@21984.4]
  assign buffer_6_479 = $signed(_T_75307); // @[Modules.scala 160:64:@21985.4]
  assign _T_75309 = $signed(buffer_6_328) + $signed(buffer_6_329); // @[Modules.scala 160:64:@21987.4]
  assign _T_75310 = _T_75309[13:0]; // @[Modules.scala 160:64:@21988.4]
  assign buffer_6_480 = $signed(_T_75310); // @[Modules.scala 160:64:@21989.4]
  assign _T_75312 = $signed(buffer_6_330) + $signed(buffer_6_331); // @[Modules.scala 160:64:@21991.4]
  assign _T_75313 = _T_75312[13:0]; // @[Modules.scala 160:64:@21992.4]
  assign buffer_6_481 = $signed(_T_75313); // @[Modules.scala 160:64:@21993.4]
  assign _T_75315 = $signed(buffer_6_332) + $signed(buffer_6_333); // @[Modules.scala 160:64:@21995.4]
  assign _T_75316 = _T_75315[13:0]; // @[Modules.scala 160:64:@21996.4]
  assign buffer_6_482 = $signed(_T_75316); // @[Modules.scala 160:64:@21997.4]
  assign _T_75318 = $signed(buffer_1_322) + $signed(buffer_6_335); // @[Modules.scala 160:64:@21999.4]
  assign _T_75319 = _T_75318[13:0]; // @[Modules.scala 160:64:@22000.4]
  assign buffer_6_483 = $signed(_T_75319); // @[Modules.scala 160:64:@22001.4]
  assign _T_75321 = $signed(buffer_1_324) + $signed(buffer_0_324); // @[Modules.scala 160:64:@22003.4]
  assign _T_75322 = _T_75321[13:0]; // @[Modules.scala 160:64:@22004.4]
  assign buffer_6_484 = $signed(_T_75322); // @[Modules.scala 160:64:@22005.4]
  assign _T_75324 = $signed(buffer_6_338) + $signed(buffer_6_339); // @[Modules.scala 160:64:@22007.4]
  assign _T_75325 = _T_75324[13:0]; // @[Modules.scala 160:64:@22008.4]
  assign buffer_6_485 = $signed(_T_75325); // @[Modules.scala 160:64:@22009.4]
  assign _T_75327 = $signed(buffer_1_328) + $signed(buffer_6_341); // @[Modules.scala 160:64:@22011.4]
  assign _T_75328 = _T_75327[13:0]; // @[Modules.scala 160:64:@22012.4]
  assign buffer_6_486 = $signed(_T_75328); // @[Modules.scala 160:64:@22013.4]
  assign _T_75330 = $signed(buffer_6_342) + $signed(buffer_6_343); // @[Modules.scala 160:64:@22015.4]
  assign _T_75331 = _T_75330[13:0]; // @[Modules.scala 160:64:@22016.4]
  assign buffer_6_487 = $signed(_T_75331); // @[Modules.scala 160:64:@22017.4]
  assign _T_75333 = $signed(buffer_6_344) + $signed(buffer_6_345); // @[Modules.scala 160:64:@22019.4]
  assign _T_75334 = _T_75333[13:0]; // @[Modules.scala 160:64:@22020.4]
  assign buffer_6_488 = $signed(_T_75334); // @[Modules.scala 160:64:@22021.4]
  assign _T_75336 = $signed(buffer_6_346) + $signed(buffer_6_347); // @[Modules.scala 160:64:@22023.4]
  assign _T_75337 = _T_75336[13:0]; // @[Modules.scala 160:64:@22024.4]
  assign buffer_6_489 = $signed(_T_75337); // @[Modules.scala 160:64:@22025.4]
  assign _T_75339 = $signed(buffer_1_336) + $signed(buffer_6_349); // @[Modules.scala 160:64:@22027.4]
  assign _T_75340 = _T_75339[13:0]; // @[Modules.scala 160:64:@22028.4]
  assign buffer_6_490 = $signed(_T_75340); // @[Modules.scala 160:64:@22029.4]
  assign _T_75342 = $signed(buffer_6_350) + $signed(buffer_6_351); // @[Modules.scala 160:64:@22031.4]
  assign _T_75343 = _T_75342[13:0]; // @[Modules.scala 160:64:@22032.4]
  assign buffer_6_491 = $signed(_T_75343); // @[Modules.scala 160:64:@22033.4]
  assign _T_75345 = $signed(buffer_6_352) + $signed(buffer_6_353); // @[Modules.scala 160:64:@22035.4]
  assign _T_75346 = _T_75345[13:0]; // @[Modules.scala 160:64:@22036.4]
  assign buffer_6_492 = $signed(_T_75346); // @[Modules.scala 160:64:@22037.4]
  assign _T_75348 = $signed(buffer_6_354) + $signed(buffer_6_355); // @[Modules.scala 160:64:@22039.4]
  assign _T_75349 = _T_75348[13:0]; // @[Modules.scala 160:64:@22040.4]
  assign buffer_6_493 = $signed(_T_75349); // @[Modules.scala 160:64:@22041.4]
  assign _T_75351 = $signed(buffer_6_356) + $signed(buffer_6_357); // @[Modules.scala 160:64:@22043.4]
  assign _T_75352 = _T_75351[13:0]; // @[Modules.scala 160:64:@22044.4]
  assign buffer_6_494 = $signed(_T_75352); // @[Modules.scala 160:64:@22045.4]
  assign _T_75354 = $signed(buffer_1_346) + $signed(buffer_3_358); // @[Modules.scala 160:64:@22047.4]
  assign _T_75355 = _T_75354[13:0]; // @[Modules.scala 160:64:@22048.4]
  assign buffer_6_495 = $signed(_T_75355); // @[Modules.scala 160:64:@22049.4]
  assign _T_75357 = $signed(buffer_6_360) + $signed(buffer_6_361); // @[Modules.scala 160:64:@22051.4]
  assign _T_75358 = _T_75357[13:0]; // @[Modules.scala 160:64:@22052.4]
  assign buffer_6_496 = $signed(_T_75358); // @[Modules.scala 160:64:@22053.4]
  assign _T_75360 = $signed(buffer_1_350) + $signed(buffer_6_363); // @[Modules.scala 160:64:@22055.4]
  assign _T_75361 = _T_75360[13:0]; // @[Modules.scala 160:64:@22056.4]
  assign buffer_6_497 = $signed(_T_75361); // @[Modules.scala 160:64:@22057.4]
  assign _T_75363 = $signed(buffer_6_364) + $signed(buffer_6_365); // @[Modules.scala 160:64:@22059.4]
  assign _T_75364 = _T_75363[13:0]; // @[Modules.scala 160:64:@22060.4]
  assign buffer_6_498 = $signed(_T_75364); // @[Modules.scala 160:64:@22061.4]
  assign _T_75366 = $signed(buffer_6_366) + $signed(buffer_6_367); // @[Modules.scala 160:64:@22063.4]
  assign _T_75367 = _T_75366[13:0]; // @[Modules.scala 160:64:@22064.4]
  assign buffer_6_499 = $signed(_T_75367); // @[Modules.scala 160:64:@22065.4]
  assign _T_75369 = $signed(buffer_6_368) + $signed(buffer_6_369); // @[Modules.scala 160:64:@22067.4]
  assign _T_75370 = _T_75369[13:0]; // @[Modules.scala 160:64:@22068.4]
  assign buffer_6_500 = $signed(_T_75370); // @[Modules.scala 160:64:@22069.4]
  assign _T_75372 = $signed(buffer_6_370) + $signed(buffer_6_371); // @[Modules.scala 160:64:@22071.4]
  assign _T_75373 = _T_75372[13:0]; // @[Modules.scala 160:64:@22072.4]
  assign buffer_6_501 = $signed(_T_75373); // @[Modules.scala 160:64:@22073.4]
  assign _T_75375 = $signed(buffer_6_372) + $signed(buffer_6_373); // @[Modules.scala 160:64:@22075.4]
  assign _T_75376 = _T_75375[13:0]; // @[Modules.scala 160:64:@22076.4]
  assign buffer_6_502 = $signed(_T_75376); // @[Modules.scala 160:64:@22077.4]
  assign _T_75378 = $signed(buffer_6_374) + $signed(buffer_6_375); // @[Modules.scala 160:64:@22079.4]
  assign _T_75379 = _T_75378[13:0]; // @[Modules.scala 160:64:@22080.4]
  assign buffer_6_503 = $signed(_T_75379); // @[Modules.scala 160:64:@22081.4]
  assign _T_75381 = $signed(buffer_6_376) + $signed(buffer_6_377); // @[Modules.scala 160:64:@22083.4]
  assign _T_75382 = _T_75381[13:0]; // @[Modules.scala 160:64:@22084.4]
  assign buffer_6_504 = $signed(_T_75382); // @[Modules.scala 160:64:@22085.4]
  assign _T_75384 = $signed(buffer_6_378) + $signed(buffer_6_379); // @[Modules.scala 160:64:@22087.4]
  assign _T_75385 = _T_75384[13:0]; // @[Modules.scala 160:64:@22088.4]
  assign buffer_6_505 = $signed(_T_75385); // @[Modules.scala 160:64:@22089.4]
  assign _T_75387 = $signed(buffer_6_380) + $signed(buffer_6_381); // @[Modules.scala 160:64:@22091.4]
  assign _T_75388 = _T_75387[13:0]; // @[Modules.scala 160:64:@22092.4]
  assign buffer_6_506 = $signed(_T_75388); // @[Modules.scala 160:64:@22093.4]
  assign _T_75390 = $signed(buffer_6_382) + $signed(buffer_6_383); // @[Modules.scala 160:64:@22095.4]
  assign _T_75391 = _T_75390[13:0]; // @[Modules.scala 160:64:@22096.4]
  assign buffer_6_507 = $signed(_T_75391); // @[Modules.scala 160:64:@22097.4]
  assign _T_75393 = $signed(buffer_6_384) + $signed(buffer_0_369); // @[Modules.scala 160:64:@22099.4]
  assign _T_75394 = _T_75393[13:0]; // @[Modules.scala 160:64:@22100.4]
  assign buffer_6_508 = $signed(_T_75394); // @[Modules.scala 160:64:@22101.4]
  assign _T_75396 = $signed(buffer_6_386) + $signed(buffer_0_371); // @[Modules.scala 160:64:@22103.4]
  assign _T_75397 = _T_75396[13:0]; // @[Modules.scala 160:64:@22104.4]
  assign buffer_6_509 = $signed(_T_75397); // @[Modules.scala 160:64:@22105.4]
  assign _T_75399 = $signed(buffer_6_388) + $signed(buffer_0_373); // @[Modules.scala 160:64:@22107.4]
  assign _T_75400 = _T_75399[13:0]; // @[Modules.scala 160:64:@22108.4]
  assign buffer_6_510 = $signed(_T_75400); // @[Modules.scala 160:64:@22109.4]
  assign _T_75402 = $signed(buffer_6_390) + $signed(buffer_6_391); // @[Modules.scala 160:64:@22111.4]
  assign _T_75403 = _T_75402[13:0]; // @[Modules.scala 160:64:@22112.4]
  assign buffer_6_511 = $signed(_T_75403); // @[Modules.scala 160:64:@22113.4]
  assign _T_75405 = $signed(buffer_6_392) + $signed(buffer_6_393); // @[Modules.scala 160:64:@22115.4]
  assign _T_75406 = _T_75405[13:0]; // @[Modules.scala 160:64:@22116.4]
  assign buffer_6_512 = $signed(_T_75406); // @[Modules.scala 160:64:@22117.4]
  assign _T_75408 = $signed(buffer_6_394) + $signed(buffer_6_395); // @[Modules.scala 160:64:@22119.4]
  assign _T_75409 = _T_75408[13:0]; // @[Modules.scala 160:64:@22120.4]
  assign buffer_6_513 = $signed(_T_75409); // @[Modules.scala 160:64:@22121.4]
  assign _T_75411 = $signed(buffer_6_396) + $signed(buffer_6_397); // @[Modules.scala 160:64:@22123.4]
  assign _T_75412 = _T_75411[13:0]; // @[Modules.scala 160:64:@22124.4]
  assign buffer_6_514 = $signed(_T_75412); // @[Modules.scala 160:64:@22125.4]
  assign _T_75414 = $signed(buffer_6_398) + $signed(buffer_6_399); // @[Modules.scala 160:64:@22127.4]
  assign _T_75415 = _T_75414[13:0]; // @[Modules.scala 160:64:@22128.4]
  assign buffer_6_515 = $signed(_T_75415); // @[Modules.scala 160:64:@22129.4]
  assign _T_75417 = $signed(buffer_6_400) + $signed(buffer_6_401); // @[Modules.scala 160:64:@22131.4]
  assign _T_75418 = _T_75417[13:0]; // @[Modules.scala 160:64:@22132.4]
  assign buffer_6_516 = $signed(_T_75418); // @[Modules.scala 160:64:@22133.4]
  assign _T_75420 = $signed(buffer_6_402) + $signed(buffer_6_403); // @[Modules.scala 160:64:@22135.4]
  assign _T_75421 = _T_75420[13:0]; // @[Modules.scala 160:64:@22136.4]
  assign buffer_6_517 = $signed(_T_75421); // @[Modules.scala 160:64:@22137.4]
  assign _T_75423 = $signed(buffer_6_404) + $signed(buffer_6_405); // @[Modules.scala 160:64:@22139.4]
  assign _T_75424 = _T_75423[13:0]; // @[Modules.scala 160:64:@22140.4]
  assign buffer_6_518 = $signed(_T_75424); // @[Modules.scala 160:64:@22141.4]
  assign _T_75426 = $signed(buffer_6_406) + $signed(buffer_6_407); // @[Modules.scala 160:64:@22143.4]
  assign _T_75427 = _T_75426[13:0]; // @[Modules.scala 160:64:@22144.4]
  assign buffer_6_519 = $signed(_T_75427); // @[Modules.scala 160:64:@22145.4]
  assign _T_75429 = $signed(buffer_6_408) + $signed(buffer_6_409); // @[Modules.scala 160:64:@22147.4]
  assign _T_75430 = _T_75429[13:0]; // @[Modules.scala 160:64:@22148.4]
  assign buffer_6_520 = $signed(_T_75430); // @[Modules.scala 160:64:@22149.4]
  assign _T_75432 = $signed(buffer_6_410) + $signed(buffer_6_411); // @[Modules.scala 160:64:@22151.4]
  assign _T_75433 = _T_75432[13:0]; // @[Modules.scala 160:64:@22152.4]
  assign buffer_6_521 = $signed(_T_75433); // @[Modules.scala 160:64:@22153.4]
  assign _T_75435 = $signed(buffer_6_412) + $signed(buffer_6_413); // @[Modules.scala 160:64:@22155.4]
  assign _T_75436 = _T_75435[13:0]; // @[Modules.scala 160:64:@22156.4]
  assign buffer_6_522 = $signed(_T_75436); // @[Modules.scala 160:64:@22157.4]
  assign _T_75438 = $signed(buffer_6_414) + $signed(buffer_6_415); // @[Modules.scala 160:64:@22159.4]
  assign _T_75439 = _T_75438[13:0]; // @[Modules.scala 160:64:@22160.4]
  assign buffer_6_523 = $signed(_T_75439); // @[Modules.scala 160:64:@22161.4]
  assign _T_75441 = $signed(buffer_6_416) + $signed(buffer_6_417); // @[Modules.scala 160:64:@22163.4]
  assign _T_75442 = _T_75441[13:0]; // @[Modules.scala 160:64:@22164.4]
  assign buffer_6_524 = $signed(_T_75442); // @[Modules.scala 160:64:@22165.4]
  assign _T_75444 = $signed(buffer_6_418) + $signed(buffer_6_419); // @[Modules.scala 160:64:@22167.4]
  assign _T_75445 = _T_75444[13:0]; // @[Modules.scala 160:64:@22168.4]
  assign buffer_6_525 = $signed(_T_75445); // @[Modules.scala 160:64:@22169.4]
  assign _T_75447 = $signed(buffer_6_420) + $signed(buffer_6_421); // @[Modules.scala 160:64:@22171.4]
  assign _T_75448 = _T_75447[13:0]; // @[Modules.scala 160:64:@22172.4]
  assign buffer_6_526 = $signed(_T_75448); // @[Modules.scala 160:64:@22173.4]
  assign _T_75450 = $signed(buffer_6_422) + $signed(buffer_0_404); // @[Modules.scala 160:64:@22175.4]
  assign _T_75451 = _T_75450[13:0]; // @[Modules.scala 160:64:@22176.4]
  assign buffer_6_527 = $signed(_T_75451); // @[Modules.scala 160:64:@22177.4]
  assign _T_75453 = $signed(buffer_0_405) + $signed(buffer_0_406); // @[Modules.scala 160:64:@22179.4]
  assign _T_75454 = _T_75453[13:0]; // @[Modules.scala 160:64:@22180.4]
  assign buffer_6_528 = $signed(_T_75454); // @[Modules.scala 160:64:@22181.4]
  assign _T_75456 = $signed(buffer_6_426) + $signed(buffer_6_427); // @[Modules.scala 160:64:@22183.4]
  assign _T_75457 = _T_75456[13:0]; // @[Modules.scala 160:64:@22184.4]
  assign buffer_6_529 = $signed(_T_75457); // @[Modules.scala 160:64:@22185.4]
  assign _T_75459 = $signed(buffer_6_428) + $signed(buffer_6_429); // @[Modules.scala 160:64:@22187.4]
  assign _T_75460 = _T_75459[13:0]; // @[Modules.scala 160:64:@22188.4]
  assign buffer_6_530 = $signed(_T_75460); // @[Modules.scala 160:64:@22189.4]
  assign _T_75462 = $signed(buffer_6_430) + $signed(buffer_6_431); // @[Modules.scala 160:64:@22191.4]
  assign _T_75463 = _T_75462[13:0]; // @[Modules.scala 160:64:@22192.4]
  assign buffer_6_531 = $signed(_T_75463); // @[Modules.scala 160:64:@22193.4]
  assign _T_75465 = $signed(buffer_6_432) + $signed(buffer_6_433); // @[Modules.scala 160:64:@22195.4]
  assign _T_75466 = _T_75465[13:0]; // @[Modules.scala 160:64:@22196.4]
  assign buffer_6_532 = $signed(_T_75466); // @[Modules.scala 160:64:@22197.4]
  assign _T_75468 = $signed(buffer_6_434) + $signed(buffer_6_435); // @[Modules.scala 160:64:@22199.4]
  assign _T_75469 = _T_75468[13:0]; // @[Modules.scala 160:64:@22200.4]
  assign buffer_6_533 = $signed(_T_75469); // @[Modules.scala 160:64:@22201.4]
  assign _T_75471 = $signed(buffer_6_436) + $signed(buffer_6_437); // @[Modules.scala 160:64:@22203.4]
  assign _T_75472 = _T_75471[13:0]; // @[Modules.scala 160:64:@22204.4]
  assign buffer_6_534 = $signed(_T_75472); // @[Modules.scala 160:64:@22205.4]
  assign _T_75474 = $signed(buffer_6_438) + $signed(buffer_6_439); // @[Modules.scala 160:64:@22207.4]
  assign _T_75475 = _T_75474[13:0]; // @[Modules.scala 160:64:@22208.4]
  assign buffer_6_535 = $signed(_T_75475); // @[Modules.scala 160:64:@22209.4]
  assign _T_75477 = $signed(buffer_6_440) + $signed(buffer_6_441); // @[Modules.scala 160:64:@22211.4]
  assign _T_75478 = _T_75477[13:0]; // @[Modules.scala 160:64:@22212.4]
  assign buffer_6_536 = $signed(_T_75478); // @[Modules.scala 160:64:@22213.4]
  assign _T_75480 = $signed(buffer_6_442) + $signed(buffer_6_443); // @[Modules.scala 160:64:@22215.4]
  assign _T_75481 = _T_75480[13:0]; // @[Modules.scala 160:64:@22216.4]
  assign buffer_6_537 = $signed(_T_75481); // @[Modules.scala 160:64:@22217.4]
  assign _T_75483 = $signed(buffer_6_444) + $signed(buffer_6_445); // @[Modules.scala 160:64:@22219.4]
  assign _T_75484 = _T_75483[13:0]; // @[Modules.scala 160:64:@22220.4]
  assign buffer_6_538 = $signed(_T_75484); // @[Modules.scala 160:64:@22221.4]
  assign _T_75486 = $signed(buffer_6_446) + $signed(buffer_6_447); // @[Modules.scala 160:64:@22223.4]
  assign _T_75487 = _T_75486[13:0]; // @[Modules.scala 160:64:@22224.4]
  assign buffer_6_539 = $signed(_T_75487); // @[Modules.scala 160:64:@22225.4]
  assign _T_75489 = $signed(buffer_6_448) + $signed(buffer_1_431); // @[Modules.scala 160:64:@22227.4]
  assign _T_75490 = _T_75489[13:0]; // @[Modules.scala 160:64:@22228.4]
  assign buffer_6_540 = $signed(_T_75490); // @[Modules.scala 160:64:@22229.4]
  assign _T_75492 = $signed(buffer_6_450) + $signed(buffer_6_451); // @[Modules.scala 160:64:@22231.4]
  assign _T_75493 = _T_75492[13:0]; // @[Modules.scala 160:64:@22232.4]
  assign buffer_6_541 = $signed(_T_75493); // @[Modules.scala 160:64:@22233.4]
  assign _T_75495 = $signed(buffer_6_452) + $signed(buffer_6_453); // @[Modules.scala 160:64:@22235.4]
  assign _T_75496 = _T_75495[13:0]; // @[Modules.scala 160:64:@22236.4]
  assign buffer_6_542 = $signed(_T_75496); // @[Modules.scala 160:64:@22237.4]
  assign _T_75498 = $signed(buffer_6_454) + $signed(buffer_6_455); // @[Modules.scala 160:64:@22239.4]
  assign _T_75499 = _T_75498[13:0]; // @[Modules.scala 160:64:@22240.4]
  assign buffer_6_543 = $signed(_T_75499); // @[Modules.scala 160:64:@22241.4]
  assign _T_75501 = $signed(buffer_6_456) + $signed(buffer_6_457); // @[Modules.scala 160:64:@22243.4]
  assign _T_75502 = _T_75501[13:0]; // @[Modules.scala 160:64:@22244.4]
  assign buffer_6_544 = $signed(_T_75502); // @[Modules.scala 160:64:@22245.4]
  assign _T_75504 = $signed(buffer_6_458) + $signed(buffer_6_459); // @[Modules.scala 160:64:@22247.4]
  assign _T_75505 = _T_75504[13:0]; // @[Modules.scala 160:64:@22248.4]
  assign buffer_6_545 = $signed(_T_75505); // @[Modules.scala 160:64:@22249.4]
  assign _T_75507 = $signed(buffer_6_460) + $signed(buffer_6_461); // @[Modules.scala 160:64:@22251.4]
  assign _T_75508 = _T_75507[13:0]; // @[Modules.scala 160:64:@22252.4]
  assign buffer_6_546 = $signed(_T_75508); // @[Modules.scala 160:64:@22253.4]
  assign _T_75510 = $signed(buffer_6_462) + $signed(buffer_6_463); // @[Modules.scala 160:64:@22255.4]
  assign _T_75511 = _T_75510[13:0]; // @[Modules.scala 160:64:@22256.4]
  assign buffer_6_547 = $signed(_T_75511); // @[Modules.scala 160:64:@22257.4]
  assign _T_75513 = $signed(buffer_6_464) + $signed(buffer_4_441); // @[Modules.scala 160:64:@22259.4]
  assign _T_75514 = _T_75513[13:0]; // @[Modules.scala 160:64:@22260.4]
  assign buffer_6_548 = $signed(_T_75514); // @[Modules.scala 160:64:@22261.4]
  assign _T_75516 = $signed(buffer_4_442) + $signed(buffer_6_467); // @[Modules.scala 160:64:@22263.4]
  assign _T_75517 = _T_75516[13:0]; // @[Modules.scala 160:64:@22264.4]
  assign buffer_6_549 = $signed(_T_75517); // @[Modules.scala 160:64:@22265.4]
  assign _T_75519 = $signed(buffer_6_468) + $signed(buffer_6_469); // @[Modules.scala 160:64:@22267.4]
  assign _T_75520 = _T_75519[13:0]; // @[Modules.scala 160:64:@22268.4]
  assign buffer_6_550 = $signed(_T_75520); // @[Modules.scala 160:64:@22269.4]
  assign _T_75522 = $signed(buffer_6_470) + $signed(buffer_6_471); // @[Modules.scala 160:64:@22271.4]
  assign _T_75523 = _T_75522[13:0]; // @[Modules.scala 160:64:@22272.4]
  assign buffer_6_551 = $signed(_T_75523); // @[Modules.scala 160:64:@22273.4]
  assign _T_75525 = $signed(buffer_6_472) + $signed(buffer_6_473); // @[Modules.scala 160:64:@22275.4]
  assign _T_75526 = _T_75525[13:0]; // @[Modules.scala 160:64:@22276.4]
  assign buffer_6_552 = $signed(_T_75526); // @[Modules.scala 160:64:@22277.4]
  assign _T_75528 = $signed(buffer_6_474) + $signed(buffer_6_475); // @[Modules.scala 166:64:@22279.4]
  assign _T_75529 = _T_75528[13:0]; // @[Modules.scala 166:64:@22280.4]
  assign buffer_6_553 = $signed(_T_75529); // @[Modules.scala 166:64:@22281.4]
  assign _T_75531 = $signed(buffer_6_476) + $signed(buffer_6_477); // @[Modules.scala 166:64:@22283.4]
  assign _T_75532 = _T_75531[13:0]; // @[Modules.scala 166:64:@22284.4]
  assign buffer_6_554 = $signed(_T_75532); // @[Modules.scala 166:64:@22285.4]
  assign _T_75534 = $signed(buffer_5_475) + $signed(buffer_6_479); // @[Modules.scala 166:64:@22287.4]
  assign _T_75535 = _T_75534[13:0]; // @[Modules.scala 166:64:@22288.4]
  assign buffer_6_555 = $signed(_T_75535); // @[Modules.scala 166:64:@22289.4]
  assign _T_75537 = $signed(buffer_6_480) + $signed(buffer_6_481); // @[Modules.scala 166:64:@22291.4]
  assign _T_75538 = _T_75537[13:0]; // @[Modules.scala 166:64:@22292.4]
  assign buffer_6_556 = $signed(_T_75538); // @[Modules.scala 166:64:@22293.4]
  assign _T_75540 = $signed(buffer_6_482) + $signed(buffer_6_483); // @[Modules.scala 166:64:@22295.4]
  assign _T_75541 = _T_75540[13:0]; // @[Modules.scala 166:64:@22296.4]
  assign buffer_6_557 = $signed(_T_75541); // @[Modules.scala 166:64:@22297.4]
  assign _T_75543 = $signed(buffer_6_484) + $signed(buffer_6_485); // @[Modules.scala 166:64:@22299.4]
  assign _T_75544 = _T_75543[13:0]; // @[Modules.scala 166:64:@22300.4]
  assign buffer_6_558 = $signed(_T_75544); // @[Modules.scala 166:64:@22301.4]
  assign _T_75546 = $signed(buffer_6_486) + $signed(buffer_6_487); // @[Modules.scala 166:64:@22303.4]
  assign _T_75547 = _T_75546[13:0]; // @[Modules.scala 166:64:@22304.4]
  assign buffer_6_559 = $signed(_T_75547); // @[Modules.scala 166:64:@22305.4]
  assign _T_75549 = $signed(buffer_6_488) + $signed(buffer_6_489); // @[Modules.scala 166:64:@22307.4]
  assign _T_75550 = _T_75549[13:0]; // @[Modules.scala 166:64:@22308.4]
  assign buffer_6_560 = $signed(_T_75550); // @[Modules.scala 166:64:@22309.4]
  assign _T_75552 = $signed(buffer_6_490) + $signed(buffer_6_491); // @[Modules.scala 166:64:@22311.4]
  assign _T_75553 = _T_75552[13:0]; // @[Modules.scala 166:64:@22312.4]
  assign buffer_6_561 = $signed(_T_75553); // @[Modules.scala 166:64:@22313.4]
  assign _T_75555 = $signed(buffer_6_492) + $signed(buffer_6_493); // @[Modules.scala 166:64:@22315.4]
  assign _T_75556 = _T_75555[13:0]; // @[Modules.scala 166:64:@22316.4]
  assign buffer_6_562 = $signed(_T_75556); // @[Modules.scala 166:64:@22317.4]
  assign _T_75558 = $signed(buffer_6_494) + $signed(buffer_6_495); // @[Modules.scala 166:64:@22319.4]
  assign _T_75559 = _T_75558[13:0]; // @[Modules.scala 166:64:@22320.4]
  assign buffer_6_563 = $signed(_T_75559); // @[Modules.scala 166:64:@22321.4]
  assign _T_75561 = $signed(buffer_6_496) + $signed(buffer_6_497); // @[Modules.scala 166:64:@22323.4]
  assign _T_75562 = _T_75561[13:0]; // @[Modules.scala 166:64:@22324.4]
  assign buffer_6_564 = $signed(_T_75562); // @[Modules.scala 166:64:@22325.4]
  assign _T_75564 = $signed(buffer_6_498) + $signed(buffer_6_499); // @[Modules.scala 166:64:@22327.4]
  assign _T_75565 = _T_75564[13:0]; // @[Modules.scala 166:64:@22328.4]
  assign buffer_6_565 = $signed(_T_75565); // @[Modules.scala 166:64:@22329.4]
  assign _T_75567 = $signed(buffer_6_500) + $signed(buffer_6_501); // @[Modules.scala 166:64:@22331.4]
  assign _T_75568 = _T_75567[13:0]; // @[Modules.scala 166:64:@22332.4]
  assign buffer_6_566 = $signed(_T_75568); // @[Modules.scala 166:64:@22333.4]
  assign _T_75570 = $signed(buffer_6_502) + $signed(buffer_6_503); // @[Modules.scala 166:64:@22335.4]
  assign _T_75571 = _T_75570[13:0]; // @[Modules.scala 166:64:@22336.4]
  assign buffer_6_567 = $signed(_T_75571); // @[Modules.scala 166:64:@22337.4]
  assign _T_75573 = $signed(buffer_6_504) + $signed(buffer_6_505); // @[Modules.scala 166:64:@22339.4]
  assign _T_75574 = _T_75573[13:0]; // @[Modules.scala 166:64:@22340.4]
  assign buffer_6_568 = $signed(_T_75574); // @[Modules.scala 166:64:@22341.4]
  assign _T_75576 = $signed(buffer_6_506) + $signed(buffer_6_507); // @[Modules.scala 166:64:@22343.4]
  assign _T_75577 = _T_75576[13:0]; // @[Modules.scala 166:64:@22344.4]
  assign buffer_6_569 = $signed(_T_75577); // @[Modules.scala 166:64:@22345.4]
  assign _T_75579 = $signed(buffer_6_508) + $signed(buffer_6_509); // @[Modules.scala 166:64:@22347.4]
  assign _T_75580 = _T_75579[13:0]; // @[Modules.scala 166:64:@22348.4]
  assign buffer_6_570 = $signed(_T_75580); // @[Modules.scala 166:64:@22349.4]
  assign _T_75582 = $signed(buffer_6_510) + $signed(buffer_6_511); // @[Modules.scala 166:64:@22351.4]
  assign _T_75583 = _T_75582[13:0]; // @[Modules.scala 166:64:@22352.4]
  assign buffer_6_571 = $signed(_T_75583); // @[Modules.scala 166:64:@22353.4]
  assign _T_75585 = $signed(buffer_6_512) + $signed(buffer_6_513); // @[Modules.scala 166:64:@22355.4]
  assign _T_75586 = _T_75585[13:0]; // @[Modules.scala 166:64:@22356.4]
  assign buffer_6_572 = $signed(_T_75586); // @[Modules.scala 166:64:@22357.4]
  assign _T_75588 = $signed(buffer_6_514) + $signed(buffer_6_515); // @[Modules.scala 166:64:@22359.4]
  assign _T_75589 = _T_75588[13:0]; // @[Modules.scala 166:64:@22360.4]
  assign buffer_6_573 = $signed(_T_75589); // @[Modules.scala 166:64:@22361.4]
  assign _T_75591 = $signed(buffer_6_516) + $signed(buffer_6_517); // @[Modules.scala 166:64:@22363.4]
  assign _T_75592 = _T_75591[13:0]; // @[Modules.scala 166:64:@22364.4]
  assign buffer_6_574 = $signed(_T_75592); // @[Modules.scala 166:64:@22365.4]
  assign _T_75594 = $signed(buffer_6_518) + $signed(buffer_6_519); // @[Modules.scala 166:64:@22367.4]
  assign _T_75595 = _T_75594[13:0]; // @[Modules.scala 166:64:@22368.4]
  assign buffer_6_575 = $signed(_T_75595); // @[Modules.scala 166:64:@22369.4]
  assign _T_75597 = $signed(buffer_6_520) + $signed(buffer_6_521); // @[Modules.scala 166:64:@22371.4]
  assign _T_75598 = _T_75597[13:0]; // @[Modules.scala 166:64:@22372.4]
  assign buffer_6_576 = $signed(_T_75598); // @[Modules.scala 166:64:@22373.4]
  assign _T_75600 = $signed(buffer_6_522) + $signed(buffer_6_523); // @[Modules.scala 166:64:@22375.4]
  assign _T_75601 = _T_75600[13:0]; // @[Modules.scala 166:64:@22376.4]
  assign buffer_6_577 = $signed(_T_75601); // @[Modules.scala 166:64:@22377.4]
  assign _T_75603 = $signed(buffer_6_524) + $signed(buffer_6_525); // @[Modules.scala 166:64:@22379.4]
  assign _T_75604 = _T_75603[13:0]; // @[Modules.scala 166:64:@22380.4]
  assign buffer_6_578 = $signed(_T_75604); // @[Modules.scala 166:64:@22381.4]
  assign _T_75606 = $signed(buffer_6_526) + $signed(buffer_6_527); // @[Modules.scala 166:64:@22383.4]
  assign _T_75607 = _T_75606[13:0]; // @[Modules.scala 166:64:@22384.4]
  assign buffer_6_579 = $signed(_T_75607); // @[Modules.scala 166:64:@22385.4]
  assign _T_75609 = $signed(buffer_6_528) + $signed(buffer_6_529); // @[Modules.scala 166:64:@22387.4]
  assign _T_75610 = _T_75609[13:0]; // @[Modules.scala 166:64:@22388.4]
  assign buffer_6_580 = $signed(_T_75610); // @[Modules.scala 166:64:@22389.4]
  assign _T_75612 = $signed(buffer_6_530) + $signed(buffer_6_531); // @[Modules.scala 166:64:@22391.4]
  assign _T_75613 = _T_75612[13:0]; // @[Modules.scala 166:64:@22392.4]
  assign buffer_6_581 = $signed(_T_75613); // @[Modules.scala 166:64:@22393.4]
  assign _T_75615 = $signed(buffer_6_532) + $signed(buffer_6_533); // @[Modules.scala 166:64:@22395.4]
  assign _T_75616 = _T_75615[13:0]; // @[Modules.scala 166:64:@22396.4]
  assign buffer_6_582 = $signed(_T_75616); // @[Modules.scala 166:64:@22397.4]
  assign _T_75618 = $signed(buffer_6_534) + $signed(buffer_6_535); // @[Modules.scala 166:64:@22399.4]
  assign _T_75619 = _T_75618[13:0]; // @[Modules.scala 166:64:@22400.4]
  assign buffer_6_583 = $signed(_T_75619); // @[Modules.scala 166:64:@22401.4]
  assign _T_75621 = $signed(buffer_6_536) + $signed(buffer_6_537); // @[Modules.scala 166:64:@22403.4]
  assign _T_75622 = _T_75621[13:0]; // @[Modules.scala 166:64:@22404.4]
  assign buffer_6_584 = $signed(_T_75622); // @[Modules.scala 166:64:@22405.4]
  assign _T_75624 = $signed(buffer_6_538) + $signed(buffer_6_539); // @[Modules.scala 166:64:@22407.4]
  assign _T_75625 = _T_75624[13:0]; // @[Modules.scala 166:64:@22408.4]
  assign buffer_6_585 = $signed(_T_75625); // @[Modules.scala 166:64:@22409.4]
  assign _T_75627 = $signed(buffer_6_540) + $signed(buffer_6_541); // @[Modules.scala 166:64:@22411.4]
  assign _T_75628 = _T_75627[13:0]; // @[Modules.scala 166:64:@22412.4]
  assign buffer_6_586 = $signed(_T_75628); // @[Modules.scala 166:64:@22413.4]
  assign _T_75630 = $signed(buffer_6_542) + $signed(buffer_6_543); // @[Modules.scala 166:64:@22415.4]
  assign _T_75631 = _T_75630[13:0]; // @[Modules.scala 166:64:@22416.4]
  assign buffer_6_587 = $signed(_T_75631); // @[Modules.scala 166:64:@22417.4]
  assign _T_75633 = $signed(buffer_6_544) + $signed(buffer_6_545); // @[Modules.scala 166:64:@22419.4]
  assign _T_75634 = _T_75633[13:0]; // @[Modules.scala 166:64:@22420.4]
  assign buffer_6_588 = $signed(_T_75634); // @[Modules.scala 166:64:@22421.4]
  assign _T_75636 = $signed(buffer_6_546) + $signed(buffer_6_547); // @[Modules.scala 166:64:@22423.4]
  assign _T_75637 = _T_75636[13:0]; // @[Modules.scala 166:64:@22424.4]
  assign buffer_6_589 = $signed(_T_75637); // @[Modules.scala 166:64:@22425.4]
  assign _T_75639 = $signed(buffer_6_548) + $signed(buffer_6_549); // @[Modules.scala 166:64:@22427.4]
  assign _T_75640 = _T_75639[13:0]; // @[Modules.scala 166:64:@22428.4]
  assign buffer_6_590 = $signed(_T_75640); // @[Modules.scala 166:64:@22429.4]
  assign _T_75642 = $signed(buffer_6_550) + $signed(buffer_6_551); // @[Modules.scala 166:64:@22431.4]
  assign _T_75643 = _T_75642[13:0]; // @[Modules.scala 166:64:@22432.4]
  assign buffer_6_591 = $signed(_T_75643); // @[Modules.scala 166:64:@22433.4]
  assign _T_75645 = $signed(buffer_6_553) + $signed(buffer_6_554); // @[Modules.scala 166:64:@22435.4]
  assign _T_75646 = _T_75645[13:0]; // @[Modules.scala 166:64:@22436.4]
  assign buffer_6_592 = $signed(_T_75646); // @[Modules.scala 166:64:@22437.4]
  assign _T_75648 = $signed(buffer_6_555) + $signed(buffer_6_556); // @[Modules.scala 166:64:@22439.4]
  assign _T_75649 = _T_75648[13:0]; // @[Modules.scala 166:64:@22440.4]
  assign buffer_6_593 = $signed(_T_75649); // @[Modules.scala 166:64:@22441.4]
  assign _T_75651 = $signed(buffer_6_557) + $signed(buffer_6_558); // @[Modules.scala 166:64:@22443.4]
  assign _T_75652 = _T_75651[13:0]; // @[Modules.scala 166:64:@22444.4]
  assign buffer_6_594 = $signed(_T_75652); // @[Modules.scala 166:64:@22445.4]
  assign _T_75654 = $signed(buffer_6_559) + $signed(buffer_6_560); // @[Modules.scala 166:64:@22447.4]
  assign _T_75655 = _T_75654[13:0]; // @[Modules.scala 166:64:@22448.4]
  assign buffer_6_595 = $signed(_T_75655); // @[Modules.scala 166:64:@22449.4]
  assign _T_75657 = $signed(buffer_6_561) + $signed(buffer_6_562); // @[Modules.scala 166:64:@22451.4]
  assign _T_75658 = _T_75657[13:0]; // @[Modules.scala 166:64:@22452.4]
  assign buffer_6_596 = $signed(_T_75658); // @[Modules.scala 166:64:@22453.4]
  assign _T_75660 = $signed(buffer_6_563) + $signed(buffer_6_564); // @[Modules.scala 166:64:@22455.4]
  assign _T_75661 = _T_75660[13:0]; // @[Modules.scala 166:64:@22456.4]
  assign buffer_6_597 = $signed(_T_75661); // @[Modules.scala 166:64:@22457.4]
  assign _T_75663 = $signed(buffer_6_565) + $signed(buffer_6_566); // @[Modules.scala 166:64:@22459.4]
  assign _T_75664 = _T_75663[13:0]; // @[Modules.scala 166:64:@22460.4]
  assign buffer_6_598 = $signed(_T_75664); // @[Modules.scala 166:64:@22461.4]
  assign _T_75666 = $signed(buffer_6_567) + $signed(buffer_6_568); // @[Modules.scala 166:64:@22463.4]
  assign _T_75667 = _T_75666[13:0]; // @[Modules.scala 166:64:@22464.4]
  assign buffer_6_599 = $signed(_T_75667); // @[Modules.scala 166:64:@22465.4]
  assign _T_75669 = $signed(buffer_6_569) + $signed(buffer_6_570); // @[Modules.scala 166:64:@22467.4]
  assign _T_75670 = _T_75669[13:0]; // @[Modules.scala 166:64:@22468.4]
  assign buffer_6_600 = $signed(_T_75670); // @[Modules.scala 166:64:@22469.4]
  assign _T_75672 = $signed(buffer_6_571) + $signed(buffer_6_572); // @[Modules.scala 166:64:@22471.4]
  assign _T_75673 = _T_75672[13:0]; // @[Modules.scala 166:64:@22472.4]
  assign buffer_6_601 = $signed(_T_75673); // @[Modules.scala 166:64:@22473.4]
  assign _T_75675 = $signed(buffer_6_573) + $signed(buffer_6_574); // @[Modules.scala 166:64:@22475.4]
  assign _T_75676 = _T_75675[13:0]; // @[Modules.scala 166:64:@22476.4]
  assign buffer_6_602 = $signed(_T_75676); // @[Modules.scala 166:64:@22477.4]
  assign _T_75678 = $signed(buffer_6_575) + $signed(buffer_6_576); // @[Modules.scala 166:64:@22479.4]
  assign _T_75679 = _T_75678[13:0]; // @[Modules.scala 166:64:@22480.4]
  assign buffer_6_603 = $signed(_T_75679); // @[Modules.scala 166:64:@22481.4]
  assign _T_75681 = $signed(buffer_6_577) + $signed(buffer_6_578); // @[Modules.scala 166:64:@22483.4]
  assign _T_75682 = _T_75681[13:0]; // @[Modules.scala 166:64:@22484.4]
  assign buffer_6_604 = $signed(_T_75682); // @[Modules.scala 166:64:@22485.4]
  assign _T_75684 = $signed(buffer_6_579) + $signed(buffer_6_580); // @[Modules.scala 166:64:@22487.4]
  assign _T_75685 = _T_75684[13:0]; // @[Modules.scala 166:64:@22488.4]
  assign buffer_6_605 = $signed(_T_75685); // @[Modules.scala 166:64:@22489.4]
  assign _T_75687 = $signed(buffer_6_581) + $signed(buffer_6_582); // @[Modules.scala 166:64:@22491.4]
  assign _T_75688 = _T_75687[13:0]; // @[Modules.scala 166:64:@22492.4]
  assign buffer_6_606 = $signed(_T_75688); // @[Modules.scala 166:64:@22493.4]
  assign _T_75690 = $signed(buffer_6_583) + $signed(buffer_6_584); // @[Modules.scala 166:64:@22495.4]
  assign _T_75691 = _T_75690[13:0]; // @[Modules.scala 166:64:@22496.4]
  assign buffer_6_607 = $signed(_T_75691); // @[Modules.scala 166:64:@22497.4]
  assign _T_75693 = $signed(buffer_6_585) + $signed(buffer_6_586); // @[Modules.scala 166:64:@22499.4]
  assign _T_75694 = _T_75693[13:0]; // @[Modules.scala 166:64:@22500.4]
  assign buffer_6_608 = $signed(_T_75694); // @[Modules.scala 166:64:@22501.4]
  assign _T_75696 = $signed(buffer_6_587) + $signed(buffer_6_588); // @[Modules.scala 166:64:@22503.4]
  assign _T_75697 = _T_75696[13:0]; // @[Modules.scala 166:64:@22504.4]
  assign buffer_6_609 = $signed(_T_75697); // @[Modules.scala 166:64:@22505.4]
  assign _T_75699 = $signed(buffer_6_589) + $signed(buffer_6_590); // @[Modules.scala 166:64:@22507.4]
  assign _T_75700 = _T_75699[13:0]; // @[Modules.scala 166:64:@22508.4]
  assign buffer_6_610 = $signed(_T_75700); // @[Modules.scala 166:64:@22509.4]
  assign _T_75702 = $signed(buffer_6_591) + $signed(buffer_6_552); // @[Modules.scala 172:66:@22511.4]
  assign _T_75703 = _T_75702[13:0]; // @[Modules.scala 172:66:@22512.4]
  assign buffer_6_611 = $signed(_T_75703); // @[Modules.scala 172:66:@22513.4]
  assign _T_75705 = $signed(buffer_6_592) + $signed(buffer_6_593); // @[Modules.scala 160:64:@22515.4]
  assign _T_75706 = _T_75705[13:0]; // @[Modules.scala 160:64:@22516.4]
  assign buffer_6_612 = $signed(_T_75706); // @[Modules.scala 160:64:@22517.4]
  assign _T_75708 = $signed(buffer_6_594) + $signed(buffer_6_595); // @[Modules.scala 160:64:@22519.4]
  assign _T_75709 = _T_75708[13:0]; // @[Modules.scala 160:64:@22520.4]
  assign buffer_6_613 = $signed(_T_75709); // @[Modules.scala 160:64:@22521.4]
  assign _T_75711 = $signed(buffer_6_596) + $signed(buffer_6_597); // @[Modules.scala 160:64:@22523.4]
  assign _T_75712 = _T_75711[13:0]; // @[Modules.scala 160:64:@22524.4]
  assign buffer_6_614 = $signed(_T_75712); // @[Modules.scala 160:64:@22525.4]
  assign _T_75714 = $signed(buffer_6_598) + $signed(buffer_6_599); // @[Modules.scala 160:64:@22527.4]
  assign _T_75715 = _T_75714[13:0]; // @[Modules.scala 160:64:@22528.4]
  assign buffer_6_615 = $signed(_T_75715); // @[Modules.scala 160:64:@22529.4]
  assign _T_75717 = $signed(buffer_6_600) + $signed(buffer_6_601); // @[Modules.scala 160:64:@22531.4]
  assign _T_75718 = _T_75717[13:0]; // @[Modules.scala 160:64:@22532.4]
  assign buffer_6_616 = $signed(_T_75718); // @[Modules.scala 160:64:@22533.4]
  assign _T_75720 = $signed(buffer_6_602) + $signed(buffer_6_603); // @[Modules.scala 160:64:@22535.4]
  assign _T_75721 = _T_75720[13:0]; // @[Modules.scala 160:64:@22536.4]
  assign buffer_6_617 = $signed(_T_75721); // @[Modules.scala 160:64:@22537.4]
  assign _T_75723 = $signed(buffer_6_604) + $signed(buffer_6_605); // @[Modules.scala 160:64:@22539.4]
  assign _T_75724 = _T_75723[13:0]; // @[Modules.scala 160:64:@22540.4]
  assign buffer_6_618 = $signed(_T_75724); // @[Modules.scala 160:64:@22541.4]
  assign _T_75726 = $signed(buffer_6_606) + $signed(buffer_6_607); // @[Modules.scala 160:64:@22543.4]
  assign _T_75727 = _T_75726[13:0]; // @[Modules.scala 160:64:@22544.4]
  assign buffer_6_619 = $signed(_T_75727); // @[Modules.scala 160:64:@22545.4]
  assign _T_75729 = $signed(buffer_6_608) + $signed(buffer_6_609); // @[Modules.scala 160:64:@22547.4]
  assign _T_75730 = _T_75729[13:0]; // @[Modules.scala 160:64:@22548.4]
  assign buffer_6_620 = $signed(_T_75730); // @[Modules.scala 160:64:@22549.4]
  assign _T_75732 = $signed(buffer_6_610) + $signed(buffer_6_611); // @[Modules.scala 160:64:@22551.4]
  assign _T_75733 = _T_75732[13:0]; // @[Modules.scala 160:64:@22552.4]
  assign buffer_6_621 = $signed(_T_75733); // @[Modules.scala 160:64:@22553.4]
  assign _T_75735 = $signed(buffer_6_612) + $signed(buffer_6_613); // @[Modules.scala 160:64:@22555.4]
  assign _T_75736 = _T_75735[13:0]; // @[Modules.scala 160:64:@22556.4]
  assign buffer_6_622 = $signed(_T_75736); // @[Modules.scala 160:64:@22557.4]
  assign _T_75738 = $signed(buffer_6_614) + $signed(buffer_6_615); // @[Modules.scala 160:64:@22559.4]
  assign _T_75739 = _T_75738[13:0]; // @[Modules.scala 160:64:@22560.4]
  assign buffer_6_623 = $signed(_T_75739); // @[Modules.scala 160:64:@22561.4]
  assign _T_75741 = $signed(buffer_6_616) + $signed(buffer_6_617); // @[Modules.scala 160:64:@22563.4]
  assign _T_75742 = _T_75741[13:0]; // @[Modules.scala 160:64:@22564.4]
  assign buffer_6_624 = $signed(_T_75742); // @[Modules.scala 160:64:@22565.4]
  assign _T_75744 = $signed(buffer_6_618) + $signed(buffer_6_619); // @[Modules.scala 160:64:@22567.4]
  assign _T_75745 = _T_75744[13:0]; // @[Modules.scala 160:64:@22568.4]
  assign buffer_6_625 = $signed(_T_75745); // @[Modules.scala 160:64:@22569.4]
  assign _T_75747 = $signed(buffer_6_620) + $signed(buffer_6_621); // @[Modules.scala 160:64:@22571.4]
  assign _T_75748 = _T_75747[13:0]; // @[Modules.scala 160:64:@22572.4]
  assign buffer_6_626 = $signed(_T_75748); // @[Modules.scala 160:64:@22573.4]
  assign _T_75750 = $signed(buffer_6_622) + $signed(buffer_6_623); // @[Modules.scala 166:64:@22575.4]
  assign _T_75751 = _T_75750[13:0]; // @[Modules.scala 166:64:@22576.4]
  assign buffer_6_627 = $signed(_T_75751); // @[Modules.scala 166:64:@22577.4]
  assign _T_75753 = $signed(buffer_6_624) + $signed(buffer_6_625); // @[Modules.scala 166:64:@22579.4]
  assign _T_75754 = _T_75753[13:0]; // @[Modules.scala 166:64:@22580.4]
  assign buffer_6_628 = $signed(_T_75754); // @[Modules.scala 166:64:@22581.4]
  assign _T_75756 = $signed(buffer_6_627) + $signed(buffer_6_628); // @[Modules.scala 160:64:@22583.4]
  assign _T_75757 = _T_75756[13:0]; // @[Modules.scala 160:64:@22584.4]
  assign buffer_6_629 = $signed(_T_75757); // @[Modules.scala 160:64:@22585.4]
  assign _T_75759 = $signed(buffer_6_629) + $signed(buffer_6_626); // @[Modules.scala 172:66:@22587.4]
  assign _T_75760 = _T_75759[13:0]; // @[Modules.scala 172:66:@22588.4]
  assign buffer_6_630 = $signed(_T_75760); // @[Modules.scala 172:66:@22589.4]
  assign _T_75763 = $signed(-4'sh1) * $signed(io_in_0); // @[Modules.scala 143:74:@22744.4]
  assign _T_75766 = $signed(_T_75763) + $signed(_T_69471); // @[Modules.scala 143:103:@22746.4]
  assign _T_75767 = _T_75766[4:0]; // @[Modules.scala 143:103:@22747.4]
  assign _T_75768 = $signed(_T_75767); // @[Modules.scala 143:103:@22748.4]
  assign _GEN_498 = {{1{_T_66500[4]}},_T_66500}; // @[Modules.scala 143:103:@22770.4]
  assign _T_75794 = $signed(_T_57232) + $signed(_GEN_498); // @[Modules.scala 143:103:@22770.4]
  assign _T_75795 = _T_75794[5:0]; // @[Modules.scala 143:103:@22771.4]
  assign _T_75796 = $signed(_T_75795); // @[Modules.scala 143:103:@22772.4]
  assign _T_75829 = $signed(_T_63403) + $signed(_T_63408); // @[Modules.scala 143:103:@22800.4]
  assign _T_75830 = _T_75829[4:0]; // @[Modules.scala 143:103:@22801.4]
  assign _T_75831 = $signed(_T_75830); // @[Modules.scala 143:103:@22802.4]
  assign _T_75857 = $signed(_T_54285) + $signed(_T_54290); // @[Modules.scala 143:103:@22824.4]
  assign _T_75858 = _T_75857[5:0]; // @[Modules.scala 143:103:@22825.4]
  assign _T_75859 = $signed(_T_75858); // @[Modules.scala 143:103:@22826.4]
  assign _T_75906 = $signed(_T_54339) + $signed(_GEN_282); // @[Modules.scala 143:103:@22866.4]
  assign _T_75907 = _T_75906[5:0]; // @[Modules.scala 143:103:@22867.4]
  assign _T_75908 = $signed(_T_75907); // @[Modules.scala 143:103:@22868.4]
  assign _T_75920 = $signed(_T_66624) + $signed(_T_54360); // @[Modules.scala 143:103:@22878.4]
  assign _T_75921 = _T_75920[5:0]; // @[Modules.scala 143:103:@22879.4]
  assign _T_75922 = $signed(_T_75921); // @[Modules.scala 143:103:@22880.4]
  assign _GEN_502 = {{1{_T_57381[4]}},_T_57381}; // @[Modules.scala 143:103:@22890.4]
  assign _T_75934 = $signed(_T_54369) + $signed(_GEN_502); // @[Modules.scala 143:103:@22890.4]
  assign _T_75935 = _T_75934[5:0]; // @[Modules.scala 143:103:@22891.4]
  assign _T_75936 = $signed(_T_75935); // @[Modules.scala 143:103:@22892.4]
  assign _GEN_503 = {{1{_T_63571[4]}},_T_63571}; // @[Modules.scala 143:103:@22944.4]
  assign _T_75997 = $signed(_T_54432) + $signed(_GEN_503); // @[Modules.scala 143:103:@22944.4]
  assign _T_75998 = _T_75997[5:0]; // @[Modules.scala 143:103:@22945.4]
  assign _T_75999 = $signed(_T_75998); // @[Modules.scala 143:103:@22946.4]
  assign _GEN_505 = {{1{_T_63585[4]}},_T_63585}; // @[Modules.scala 143:103:@22956.4]
  assign _T_76011 = $signed(_T_57449) + $signed(_GEN_505); // @[Modules.scala 143:103:@22956.4]
  assign _T_76012 = _T_76011[5:0]; // @[Modules.scala 143:103:@22957.4]
  assign _T_76013 = $signed(_T_76012); // @[Modules.scala 143:103:@22958.4]
  assign _GEN_506 = {{1{_T_63604[4]}},_T_63604}; // @[Modules.scala 143:103:@22974.4]
  assign _T_76032 = $signed(_GEN_506) + $signed(_T_54467); // @[Modules.scala 143:103:@22974.4]
  assign _T_76033 = _T_76032[5:0]; // @[Modules.scala 143:103:@22975.4]
  assign _T_76034 = $signed(_T_76033); // @[Modules.scala 143:103:@22976.4]
  assign _T_76046 = $signed(_T_60509) + $signed(_T_57486); // @[Modules.scala 143:103:@22986.4]
  assign _T_76047 = _T_76046[4:0]; // @[Modules.scala 143:103:@22987.4]
  assign _T_76048 = $signed(_T_76047); // @[Modules.scala 143:103:@22988.4]
  assign _T_76052 = $signed(-4'sh1) * $signed(io_in_130); // @[Modules.scala 144:80:@22991.4]
  assign _T_76053 = $signed(_T_66750) + $signed(_T_76052); // @[Modules.scala 143:103:@22992.4]
  assign _T_76054 = _T_76053[4:0]; // @[Modules.scala 143:103:@22993.4]
  assign _T_76055 = $signed(_T_76054); // @[Modules.scala 143:103:@22994.4]
  assign _T_76057 = $signed(-4'sh1) * $signed(io_in_131); // @[Modules.scala 143:74:@22996.4]
  assign _T_76060 = $signed(_T_76057) + $signed(_T_69765); // @[Modules.scala 143:103:@22998.4]
  assign _T_76061 = _T_76060[4:0]; // @[Modules.scala 143:103:@22999.4]
  assign _T_76062 = $signed(_T_76061); // @[Modules.scala 143:103:@23000.4]
  assign _GEN_507 = {{1{_T_69770[4]}},_T_69770}; // @[Modules.scala 143:103:@23004.4]
  assign _T_76067 = $signed(_GEN_507) + $signed(_T_57507); // @[Modules.scala 143:103:@23004.4]
  assign _T_76068 = _T_76067[5:0]; // @[Modules.scala 143:103:@23005.4]
  assign _T_76069 = $signed(_T_76068); // @[Modules.scala 143:103:@23006.4]
  assign _T_76081 = $signed(_T_54516) + $signed(_T_57526); // @[Modules.scala 143:103:@23016.4]
  assign _T_76082 = _T_76081[5:0]; // @[Modules.scala 143:103:@23017.4]
  assign _T_76083 = $signed(_T_76082); // @[Modules.scala 143:103:@23018.4]
  assign _GEN_509 = {{1{_T_60584[4]}},_T_60584}; // @[Modules.scala 143:103:@23040.4]
  assign _T_76109 = $signed(_T_54535) + $signed(_GEN_509); // @[Modules.scala 143:103:@23040.4]
  assign _T_76110 = _T_76109[5:0]; // @[Modules.scala 143:103:@23041.4]
  assign _T_76111 = $signed(_T_76110); // @[Modules.scala 143:103:@23042.4]
  assign _T_76122 = $signed(4'sh1) * $signed(io_in_158); // @[Modules.scala 144:80:@23051.4]
  assign _T_76123 = $signed(_T_69833) + $signed(_T_76122); // @[Modules.scala 143:103:@23052.4]
  assign _T_76124 = _T_76123[5:0]; // @[Modules.scala 143:103:@23053.4]
  assign _T_76125 = $signed(_T_76124); // @[Modules.scala 143:103:@23054.4]
  assign _T_76130 = $signed(_T_54556) + $signed(_T_63730); // @[Modules.scala 143:103:@23058.4]
  assign _T_76131 = _T_76130[5:0]; // @[Modules.scala 143:103:@23059.4]
  assign _T_76132 = $signed(_T_76131); // @[Modules.scala 143:103:@23060.4]
  assign _T_76137 = $signed(_T_60614) + $signed(_T_60619); // @[Modules.scala 143:103:@23064.4]
  assign _T_76138 = _T_76137[5:0]; // @[Modules.scala 143:103:@23065.4]
  assign _T_76139 = $signed(_T_76138); // @[Modules.scala 143:103:@23066.4]
  assign _T_76144 = $signed(_T_63739) + $signed(_T_54572); // @[Modules.scala 143:103:@23070.4]
  assign _T_76145 = _T_76144[5:0]; // @[Modules.scala 143:103:@23071.4]
  assign _T_76146 = $signed(_T_76145); // @[Modules.scala 143:103:@23072.4]
  assign _T_76150 = $signed(4'sh1) * $signed(io_in_168); // @[Modules.scala 144:80:@23075.4]
  assign _T_76151 = $signed(_GEN_225) + $signed(_T_76150); // @[Modules.scala 143:103:@23076.4]
  assign _T_76152 = _T_76151[5:0]; // @[Modules.scala 143:103:@23077.4]
  assign _T_76153 = $signed(_T_76152); // @[Modules.scala 143:103:@23078.4]
  assign _T_76165 = $signed(_GEN_159) + $signed(_T_54598); // @[Modules.scala 143:103:@23088.4]
  assign _T_76166 = _T_76165[5:0]; // @[Modules.scala 143:103:@23089.4]
  assign _T_76167 = $signed(_T_76166); // @[Modules.scala 143:103:@23090.4]
  assign _T_76186 = $signed(_T_60656) + $signed(_T_54614); // @[Modules.scala 143:103:@23106.4]
  assign _T_76187 = _T_76186[4:0]; // @[Modules.scala 143:103:@23107.4]
  assign _T_76188 = $signed(_T_76187); // @[Modules.scala 143:103:@23108.4]
  assign _GEN_513 = {{1{_T_54628[4]}},_T_54628}; // @[Modules.scala 143:103:@23124.4]
  assign _T_76207 = $signed(_GEN_513) + $signed(_T_73049); // @[Modules.scala 143:103:@23124.4]
  assign _T_76208 = _T_76207[5:0]; // @[Modules.scala 143:103:@23125.4]
  assign _T_76209 = $signed(_T_76208); // @[Modules.scala 143:103:@23126.4]
  assign _T_76228 = $signed(_T_69938) + $signed(_T_54654); // @[Modules.scala 143:103:@23142.4]
  assign _T_76229 = _T_76228[5:0]; // @[Modules.scala 143:103:@23143.4]
  assign _T_76230 = $signed(_T_76229); // @[Modules.scala 143:103:@23144.4]
  assign _T_76242 = $signed(_T_54668) + $signed(_T_54675); // @[Modules.scala 143:103:@23154.4]
  assign _T_76243 = _T_76242[5:0]; // @[Modules.scala 143:103:@23155.4]
  assign _T_76244 = $signed(_T_76243); // @[Modules.scala 143:103:@23156.4]
  assign _T_76284 = $signed(_GEN_230) + $signed(_T_70010); // @[Modules.scala 143:103:@23190.4]
  assign _T_76285 = _T_76284[5:0]; // @[Modules.scala 143:103:@23191.4]
  assign _T_76286 = $signed(_T_76285); // @[Modules.scala 143:103:@23192.4]
  assign _T_76291 = $signed(_T_63893) + $signed(_T_63898); // @[Modules.scala 143:103:@23196.4]
  assign _T_76292 = _T_76291[5:0]; // @[Modules.scala 143:103:@23197.4]
  assign _T_76293 = $signed(_T_76292); // @[Modules.scala 143:103:@23198.4]
  assign _T_76298 = $signed(_T_63900) + $signed(_T_63905); // @[Modules.scala 143:103:@23202.4]
  assign _T_76299 = _T_76298[5:0]; // @[Modules.scala 143:103:@23203.4]
  assign _T_76300 = $signed(_T_76299); // @[Modules.scala 143:103:@23204.4]
  assign _T_76305 = $signed(_T_63907) + $signed(_T_54724); // @[Modules.scala 143:103:@23208.4]
  assign _T_76306 = _T_76305[5:0]; // @[Modules.scala 143:103:@23209.4]
  assign _T_76307 = $signed(_T_76306); // @[Modules.scala 143:103:@23210.4]
  assign _T_76340 = $signed(_T_54754) + $signed(_T_70057); // @[Modules.scala 143:103:@23238.4]
  assign _T_76341 = _T_76340[5:0]; // @[Modules.scala 143:103:@23239.4]
  assign _T_76342 = $signed(_T_76341); // @[Modules.scala 143:103:@23240.4]
  assign _T_76347 = $signed(_T_70059) + $signed(_T_54761); // @[Modules.scala 143:103:@23244.4]
  assign _T_76348 = _T_76347[5:0]; // @[Modules.scala 143:103:@23245.4]
  assign _T_76349 = $signed(_T_76348); // @[Modules.scala 143:103:@23246.4]
  assign _GEN_516 = {{1{_T_60845[4]}},_T_60845}; // @[Modules.scala 143:103:@23250.4]
  assign _T_76354 = $signed(_T_67053) + $signed(_GEN_516); // @[Modules.scala 143:103:@23250.4]
  assign _T_76355 = _T_76354[5:0]; // @[Modules.scala 143:103:@23251.4]
  assign _T_76356 = $signed(_T_76355); // @[Modules.scala 143:103:@23252.4]
  assign _T_76368 = $signed(_T_57813) + $signed(_T_63970); // @[Modules.scala 143:103:@23262.4]
  assign _T_76369 = _T_76368[5:0]; // @[Modules.scala 143:103:@23263.4]
  assign _T_76370 = $signed(_T_76369); // @[Modules.scala 143:103:@23264.4]
  assign _T_76466 = $signed(_T_70192) + $signed(_T_64061); // @[Modules.scala 143:103:@23346.4]
  assign _T_76467 = _T_76466[5:0]; // @[Modules.scala 143:103:@23347.4]
  assign _T_76468 = $signed(_T_76467); // @[Modules.scala 143:103:@23348.4]
  assign _GEN_518 = {{1{_T_54955[4]}},_T_54955}; // @[Modules.scala 143:103:@23418.4]
  assign _T_76550 = $signed(_T_57976) + $signed(_GEN_518); // @[Modules.scala 143:103:@23418.4]
  assign _T_76551 = _T_76550[5:0]; // @[Modules.scala 143:103:@23419.4]
  assign _T_76552 = $signed(_T_76551); // @[Modules.scala 143:103:@23420.4]
  assign _GEN_519 = {{1{_T_54985[4]}},_T_54985}; // @[Modules.scala 143:103:@23436.4]
  assign _T_76571 = $signed(_GEN_519) + $signed(_T_58018); // @[Modules.scala 143:103:@23436.4]
  assign _T_76572 = _T_76571[5:0]; // @[Modules.scala 143:103:@23437.4]
  assign _T_76573 = $signed(_T_76572); // @[Modules.scala 143:103:@23438.4]
  assign _T_76606 = $signed(_T_61097) + $signed(_GEN_28); // @[Modules.scala 143:103:@23466.4]
  assign _T_76607 = _T_76606[5:0]; // @[Modules.scala 143:103:@23467.4]
  assign _T_76608 = $signed(_T_76607); // @[Modules.scala 143:103:@23468.4]
  assign _GEN_521 = {{1{_T_55067[4]}},_T_55067}; // @[Modules.scala 143:103:@23496.4]
  assign _T_76641 = $signed(_GEN_521) + $signed(_T_64262); // @[Modules.scala 143:103:@23496.4]
  assign _T_76642 = _T_76641[5:0]; // @[Modules.scala 143:103:@23497.4]
  assign _T_76643 = $signed(_T_76642); // @[Modules.scala 143:103:@23498.4]
  assign _T_76648 = $signed(_T_64264) + $signed(_T_58100); // @[Modules.scala 143:103:@23502.4]
  assign _T_76649 = _T_76648[5:0]; // @[Modules.scala 143:103:@23503.4]
  assign _T_76650 = $signed(_T_76649); // @[Modules.scala 143:103:@23504.4]
  assign _GEN_523 = {{1{_T_55104[4]}},_T_55104}; // @[Modules.scala 143:103:@23520.4]
  assign _T_76669 = $signed(_T_58116) + $signed(_GEN_523); // @[Modules.scala 143:103:@23520.4]
  assign _T_76670 = _T_76669[5:0]; // @[Modules.scala 143:103:@23521.4]
  assign _T_76671 = $signed(_T_76670); // @[Modules.scala 143:103:@23522.4]
  assign _T_76696 = $signed(-4'sh1) * $signed(io_in_355); // @[Modules.scala 144:80:@23543.4]
  assign _T_76697 = $signed(_T_55132) + $signed(_T_76696); // @[Modules.scala 143:103:@23544.4]
  assign _T_76698 = _T_76697[4:0]; // @[Modules.scala 143:103:@23545.4]
  assign _T_76699 = $signed(_T_76698); // @[Modules.scala 143:103:@23546.4]
  assign _T_76778 = $signed(-4'sh1) * $signed(io_in_380); // @[Modules.scala 143:74:@23614.4]
  assign _T_76781 = $signed(_T_76778) + $signed(_T_55216); // @[Modules.scala 143:103:@23616.4]
  assign _T_76782 = _T_76781[4:0]; // @[Modules.scala 143:103:@23617.4]
  assign _T_76783 = $signed(_T_76782); // @[Modules.scala 143:103:@23618.4]
  assign _T_76787 = $signed(-4'sh1) * $signed(io_in_383); // @[Modules.scala 144:80:@23621.4]
  assign _T_76788 = $signed(_T_73663) + $signed(_T_76787); // @[Modules.scala 143:103:@23622.4]
  assign _T_76789 = _T_76788[4:0]; // @[Modules.scala 143:103:@23623.4]
  assign _T_76790 = $signed(_T_76789); // @[Modules.scala 143:103:@23624.4]
  assign _T_76809 = $signed(_GEN_36) + $signed(_T_58270); // @[Modules.scala 143:103:@23640.4]
  assign _T_76810 = _T_76809[5:0]; // @[Modules.scala 143:103:@23641.4]
  assign _T_76811 = $signed(_T_76810); // @[Modules.scala 143:103:@23642.4]
  assign _T_76816 = $signed(_T_55244) + $signed(_T_55249); // @[Modules.scala 143:103:@23646.4]
  assign _T_76817 = _T_76816[5:0]; // @[Modules.scala 143:103:@23647.4]
  assign _T_76818 = $signed(_T_76817); // @[Modules.scala 143:103:@23648.4]
  assign _T_76823 = $signed(_GEN_38) + $signed(_T_55256); // @[Modules.scala 143:103:@23652.4]
  assign _T_76824 = _T_76823[5:0]; // @[Modules.scala 143:103:@23653.4]
  assign _T_76825 = $signed(_T_76824); // @[Modules.scala 143:103:@23654.4]
  assign _GEN_528 = {{1{_T_55263[4]}},_T_55263}; // @[Modules.scala 143:103:@23658.4]
  assign _T_76830 = $signed(_T_55258) + $signed(_GEN_528); // @[Modules.scala 143:103:@23658.4]
  assign _T_76831 = _T_76830[5:0]; // @[Modules.scala 143:103:@23659.4]
  assign _T_76832 = $signed(_T_76831); // @[Modules.scala 143:103:@23660.4]
  assign _GEN_529 = {{1{_T_67550[4]}},_T_67550}; // @[Modules.scala 143:103:@23688.4]
  assign _T_76865 = $signed(_GEN_529) + $signed(_T_55293); // @[Modules.scala 143:103:@23688.4]
  assign _T_76866 = _T_76865[5:0]; // @[Modules.scala 143:103:@23689.4]
  assign _T_76867 = $signed(_T_76866); // @[Modules.scala 143:103:@23690.4]
  assign _T_76872 = $signed(_T_55300) + $signed(_T_55305); // @[Modules.scala 143:103:@23694.4]
  assign _T_76873 = _T_76872[4:0]; // @[Modules.scala 143:103:@23695.4]
  assign _T_76874 = $signed(_T_76873); // @[Modules.scala 143:103:@23696.4]
  assign _T_76879 = $signed(_T_70584) + $signed(_T_70589); // @[Modules.scala 143:103:@23700.4]
  assign _T_76880 = _T_76879[4:0]; // @[Modules.scala 143:103:@23701.4]
  assign _T_76881 = $signed(_T_76880); // @[Modules.scala 143:103:@23702.4]
  assign _T_76900 = $signed(_T_58340) + $signed(_T_55321); // @[Modules.scala 143:103:@23718.4]
  assign _T_76901 = _T_76900[4:0]; // @[Modules.scala 143:103:@23719.4]
  assign _T_76902 = $signed(_T_76901); // @[Modules.scala 143:103:@23720.4]
  assign _T_76914 = $signed(_T_55333) + $signed(_T_67597); // @[Modules.scala 143:103:@23730.4]
  assign _T_76915 = _T_76914[4:0]; // @[Modules.scala 143:103:@23731.4]
  assign _T_76916 = $signed(_T_76915); // @[Modules.scala 143:103:@23732.4]
  assign _T_76921 = $signed(_T_70626) + $signed(_T_55342); // @[Modules.scala 143:103:@23736.4]
  assign _T_76922 = _T_76921[4:0]; // @[Modules.scala 143:103:@23737.4]
  assign _T_76923 = $signed(_T_76922); // @[Modules.scala 143:103:@23738.4]
  assign _T_76942 = $signed(_T_55356) + $signed(_T_55361); // @[Modules.scala 143:103:@23754.4]
  assign _T_76943 = _T_76942[4:0]; // @[Modules.scala 143:103:@23755.4]
  assign _T_76944 = $signed(_T_76943); // @[Modules.scala 143:103:@23756.4]
  assign _T_76963 = $signed(_T_70666) + $signed(_T_55377); // @[Modules.scala 143:103:@23772.4]
  assign _T_76964 = _T_76963[4:0]; // @[Modules.scala 143:103:@23773.4]
  assign _T_76965 = $signed(_T_76964); // @[Modules.scala 143:103:@23774.4]
  assign _T_76998 = $signed(_T_55405) + $signed(_T_55410); // @[Modules.scala 143:103:@23802.4]
  assign _T_76999 = _T_76998[5:0]; // @[Modules.scala 143:103:@23803.4]
  assign _T_77000 = $signed(_T_76999); // @[Modules.scala 143:103:@23804.4]
  assign _T_77005 = $signed(_T_55412) + $signed(_GEN_179); // @[Modules.scala 143:103:@23808.4]
  assign _T_77006 = _T_77005[5:0]; // @[Modules.scala 143:103:@23809.4]
  assign _T_77007 = $signed(_T_77006); // @[Modules.scala 143:103:@23810.4]
  assign _GEN_533 = {{1{_T_58492[4]}},_T_58492}; // @[Modules.scala 143:103:@23880.4]
  assign _T_77089 = $signed(_GEN_533) + $signed(_T_55480); // @[Modules.scala 143:103:@23880.4]
  assign _T_77090 = _T_77089[5:0]; // @[Modules.scala 143:103:@23881.4]
  assign _T_77091 = $signed(_T_77090); // @[Modules.scala 143:103:@23882.4]
  assign _T_77103 = $signed(_T_55487) + $signed(_T_61585); // @[Modules.scala 143:103:@23892.4]
  assign _T_77104 = _T_77103[4:0]; // @[Modules.scala 143:103:@23893.4]
  assign _T_77105 = $signed(_T_77104); // @[Modules.scala 143:103:@23894.4]
  assign _T_77152 = $signed(_T_55531) + $signed(_T_55536); // @[Modules.scala 143:103:@23934.4]
  assign _T_77153 = _T_77152[4:0]; // @[Modules.scala 143:103:@23935.4]
  assign _T_77154 = $signed(_T_77153); // @[Modules.scala 143:103:@23936.4]
  assign _T_77166 = $signed(_T_64754) + $signed(_T_61629); // @[Modules.scala 143:103:@23946.4]
  assign _T_77167 = _T_77166[4:0]; // @[Modules.scala 143:103:@23947.4]
  assign _T_77168 = $signed(_T_77167); // @[Modules.scala 143:103:@23948.4]
  assign _T_77187 = $signed(_T_55557) + $signed(_GEN_406); // @[Modules.scala 143:103:@23964.4]
  assign _T_77188 = _T_77187[5:0]; // @[Modules.scala 143:103:@23965.4]
  assign _T_77189 = $signed(_T_77188); // @[Modules.scala 143:103:@23966.4]
  assign _T_77194 = $signed(_T_64782) + $signed(_T_61657); // @[Modules.scala 143:103:@23970.4]
  assign _T_77195 = _T_77194[4:0]; // @[Modules.scala 143:103:@23971.4]
  assign _T_77196 = $signed(_T_77195); // @[Modules.scala 143:103:@23972.4]
  assign _T_77215 = $signed(_T_55587) + $signed(_T_55592); // @[Modules.scala 143:103:@23988.4]
  assign _T_77216 = _T_77215[5:0]; // @[Modules.scala 143:103:@23989.4]
  assign _T_77217 = $signed(_T_77216); // @[Modules.scala 143:103:@23990.4]
  assign _T_77222 = $signed(_T_55594) + $signed(_T_55599); // @[Modules.scala 143:103:@23994.4]
  assign _T_77223 = _T_77222[5:0]; // @[Modules.scala 143:103:@23995.4]
  assign _T_77224 = $signed(_T_77223); // @[Modules.scala 143:103:@23996.4]
  assign _T_77229 = $signed(_T_55601) + $signed(_T_55606); // @[Modules.scala 143:103:@24000.4]
  assign _T_77230 = _T_77229[5:0]; // @[Modules.scala 143:103:@24001.4]
  assign _T_77231 = $signed(_T_77230); // @[Modules.scala 143:103:@24002.4]
  assign _T_77243 = $signed(_T_61699) + $signed(_T_64829); // @[Modules.scala 143:103:@24012.4]
  assign _T_77244 = _T_77243[4:0]; // @[Modules.scala 143:103:@24013.4]
  assign _T_77245 = $signed(_T_77244); // @[Modules.scala 143:103:@24014.4]
  assign _T_77250 = $signed(_GEN_409) + $signed(_T_55622); // @[Modules.scala 143:103:@24018.4]
  assign _T_77251 = _T_77250[5:0]; // @[Modules.scala 143:103:@24019.4]
  assign _T_77252 = $signed(_T_77251); // @[Modules.scala 143:103:@24020.4]
  assign _T_77257 = $signed(_T_64838) + $signed(_T_61706); // @[Modules.scala 143:103:@24024.4]
  assign _T_77258 = _T_77257[4:0]; // @[Modules.scala 143:103:@24025.4]
  assign _T_77259 = $signed(_T_77258); // @[Modules.scala 143:103:@24026.4]
  assign _GEN_537 = {{1{_T_58639[4]}},_T_58639}; // @[Modules.scala 143:103:@24030.4]
  assign _T_77264 = $signed(_GEN_537) + $signed(_T_55634); // @[Modules.scala 143:103:@24030.4]
  assign _T_77265 = _T_77264[5:0]; // @[Modules.scala 143:103:@24031.4]
  assign _T_77266 = $signed(_T_77265); // @[Modules.scala 143:103:@24032.4]
  assign _T_77278 = $signed(_T_55643) + $signed(_GEN_61); // @[Modules.scala 143:103:@24042.4]
  assign _T_77279 = _T_77278[5:0]; // @[Modules.scala 143:103:@24043.4]
  assign _T_77280 = $signed(_T_77279); // @[Modules.scala 143:103:@24044.4]
  assign _T_77327 = $signed(_T_55697) + $signed(_GEN_120); // @[Modules.scala 143:103:@24084.4]
  assign _T_77328 = _T_77327[5:0]; // @[Modules.scala 143:103:@24085.4]
  assign _T_77329 = $signed(_T_77328); // @[Modules.scala 143:103:@24086.4]
  assign _T_77334 = $signed(_T_64920) + $signed(_T_58718); // @[Modules.scala 143:103:@24090.4]
  assign _T_77335 = _T_77334[4:0]; // @[Modules.scala 143:103:@24091.4]
  assign _T_77336 = $signed(_T_77335); // @[Modules.scala 143:103:@24092.4]
  assign _T_77355 = $signed(_T_55720) + $signed(_T_64943); // @[Modules.scala 143:103:@24108.4]
  assign _T_77356 = _T_77355[5:0]; // @[Modules.scala 143:103:@24109.4]
  assign _T_77357 = $signed(_T_77356); // @[Modules.scala 143:103:@24110.4]
  assign _T_77382 = $signed(4'sh1) * $signed(io_in_569); // @[Modules.scala 144:80:@24131.4]
  assign _T_77383 = $signed(_T_64969) + $signed(_T_77382); // @[Modules.scala 143:103:@24132.4]
  assign _T_77384 = _T_77383[5:0]; // @[Modules.scala 143:103:@24133.4]
  assign _T_77385 = $signed(_T_77384); // @[Modules.scala 143:103:@24134.4]
  assign _T_77390 = $signed(_T_55748) + $signed(_T_55753); // @[Modules.scala 143:103:@24138.4]
  assign _T_77391 = _T_77390[5:0]; // @[Modules.scala 143:103:@24139.4]
  assign _T_77392 = $signed(_T_77391); // @[Modules.scala 143:103:@24140.4]
  assign _T_77397 = $signed(_T_55755) + $signed(_T_55760); // @[Modules.scala 143:103:@24144.4]
  assign _T_77398 = _T_77397[5:0]; // @[Modules.scala 143:103:@24145.4]
  assign _T_77399 = $signed(_T_77398); // @[Modules.scala 143:103:@24146.4]
  assign _T_77404 = $signed(_T_55762) + $signed(_T_74260); // @[Modules.scala 143:103:@24150.4]
  assign _T_77405 = _T_77404[5:0]; // @[Modules.scala 143:103:@24151.4]
  assign _T_77406 = $signed(_T_77405); // @[Modules.scala 143:103:@24152.4]
  assign _GEN_540 = {{1{_T_61858[4]}},_T_61858}; // @[Modules.scala 143:103:@24156.4]
  assign _T_77411 = $signed(_T_55767) + $signed(_GEN_540); // @[Modules.scala 143:103:@24156.4]
  assign _T_77412 = _T_77411[5:0]; // @[Modules.scala 143:103:@24157.4]
  assign _T_77413 = $signed(_T_77412); // @[Modules.scala 143:103:@24158.4]
  assign _T_77418 = $signed(_T_55769) + $signed(_T_58793); // @[Modules.scala 143:103:@24162.4]
  assign _T_77419 = _T_77418[4:0]; // @[Modules.scala 143:103:@24163.4]
  assign _T_77420 = $signed(_T_77419); // @[Modules.scala 143:103:@24164.4]
  assign _T_77425 = $signed(_GEN_64) + $signed(_T_55781); // @[Modules.scala 143:103:@24168.4]
  assign _T_77426 = _T_77425[5:0]; // @[Modules.scala 143:103:@24169.4]
  assign _T_77427 = $signed(_T_77426); // @[Modules.scala 143:103:@24170.4]
  assign _T_77432 = $signed(_T_55783) + $signed(_T_58809); // @[Modules.scala 143:103:@24174.4]
  assign _T_77433 = _T_77432[5:0]; // @[Modules.scala 143:103:@24175.4]
  assign _T_77434 = $signed(_T_77433); // @[Modules.scala 143:103:@24176.4]
  assign _T_77446 = $signed(_T_71116) + $signed(_T_68038); // @[Modules.scala 143:103:@24186.4]
  assign _T_77447 = _T_77446[4:0]; // @[Modules.scala 143:103:@24187.4]
  assign _T_77448 = $signed(_T_77447); // @[Modules.scala 143:103:@24188.4]
  assign _GEN_542 = {{1{_T_61902[4]}},_T_61902}; // @[Modules.scala 143:103:@24198.4]
  assign _T_77460 = $signed(_GEN_542) + $signed(_T_55811); // @[Modules.scala 143:103:@24198.4]
  assign _T_77461 = _T_77460[5:0]; // @[Modules.scala 143:103:@24199.4]
  assign _T_77462 = $signed(_T_77461); // @[Modules.scala 143:103:@24200.4]
  assign _T_77464 = $signed(4'sh1) * $signed(io_in_597); // @[Modules.scala 143:74:@24202.4]
  assign _T_77467 = $signed(_T_77464) + $signed(_GEN_126); // @[Modules.scala 143:103:@24204.4]
  assign _T_77468 = _T_77467[5:0]; // @[Modules.scala 143:103:@24205.4]
  assign _T_77469 = $signed(_T_77468); // @[Modules.scala 143:103:@24206.4]
  assign _T_77481 = $signed(_GEN_485) + $signed(_T_74330); // @[Modules.scala 143:103:@24216.4]
  assign _T_77482 = _T_77481[5:0]; // @[Modules.scala 143:103:@24217.4]
  assign _T_77483 = $signed(_T_77482); // @[Modules.scala 143:103:@24218.4]
  assign _GEN_545 = {{1{_T_61944[4]}},_T_61944}; // @[Modules.scala 143:103:@24222.4]
  assign _T_77488 = $signed(_GEN_545) + $signed(_T_71179); // @[Modules.scala 143:103:@24222.4]
  assign _T_77489 = _T_77488[5:0]; // @[Modules.scala 143:103:@24223.4]
  assign _T_77490 = $signed(_T_77489); // @[Modules.scala 143:103:@24224.4]
  assign _T_77495 = $signed(_GEN_486) + $signed(_T_55846); // @[Modules.scala 143:103:@24228.4]
  assign _T_77496 = _T_77495[5:0]; // @[Modules.scala 143:103:@24229.4]
  assign _T_77497 = $signed(_T_77496); // @[Modules.scala 143:103:@24230.4]
  assign _T_77516 = $signed(_T_65083) + $signed(_T_61979); // @[Modules.scala 143:103:@24246.4]
  assign _T_77517 = _T_77516[4:0]; // @[Modules.scala 143:103:@24247.4]
  assign _T_77518 = $signed(_T_77517); // @[Modules.scala 143:103:@24248.4]
  assign _GEN_547 = {{1{_T_61984[4]}},_T_61984}; // @[Modules.scala 143:103:@24252.4]
  assign _T_77523 = $signed(_GEN_547) + $signed(_T_55879); // @[Modules.scala 143:103:@24252.4]
  assign _T_77524 = _T_77523[5:0]; // @[Modules.scala 143:103:@24253.4]
  assign _T_77525 = $signed(_T_77524); // @[Modules.scala 143:103:@24254.4]
  assign _T_77544 = $signed(_T_55895) + $signed(_T_55907); // @[Modules.scala 143:103:@24270.4]
  assign _T_77545 = _T_77544[4:0]; // @[Modules.scala 143:103:@24271.4]
  assign _T_77546 = $signed(_T_77545); // @[Modules.scala 143:103:@24272.4]
  assign _GEN_549 = {{1{_T_55909[4]}},_T_55909}; // @[Modules.scala 143:103:@24276.4]
  assign _T_77551 = $signed(_GEN_549) + $signed(_T_62026); // @[Modules.scala 143:103:@24276.4]
  assign _T_77552 = _T_77551[5:0]; // @[Modules.scala 143:103:@24277.4]
  assign _T_77553 = $signed(_T_77552); // @[Modules.scala 143:103:@24278.4]
  assign _T_77558 = $signed(_T_55928) + $signed(_T_55935); // @[Modules.scala 143:103:@24282.4]
  assign _T_77559 = _T_77558[5:0]; // @[Modules.scala 143:103:@24283.4]
  assign _T_77560 = $signed(_T_77559); // @[Modules.scala 143:103:@24284.4]
  assign _GEN_551 = {{1{_T_62056[4]}},_T_62056}; // @[Modules.scala 143:103:@24306.4]
  assign _T_77586 = $signed(_GEN_551) + $signed(_T_55963); // @[Modules.scala 143:103:@24306.4]
  assign _T_77587 = _T_77586[5:0]; // @[Modules.scala 143:103:@24307.4]
  assign _T_77588 = $signed(_T_77587); // @[Modules.scala 143:103:@24308.4]
  assign _T_77600 = $signed(_T_55972) + $signed(_T_55977); // @[Modules.scala 143:103:@24318.4]
  assign _T_77601 = _T_77600[4:0]; // @[Modules.scala 143:103:@24319.4]
  assign _T_77602 = $signed(_T_77601); // @[Modules.scala 143:103:@24320.4]
  assign _T_77607 = $signed(_GEN_347) + $signed(_T_65188); // @[Modules.scala 143:103:@24324.4]
  assign _T_77608 = _T_77607[5:0]; // @[Modules.scala 143:103:@24325.4]
  assign _T_77609 = $signed(_T_77608); // @[Modules.scala 143:103:@24326.4]
  assign _T_77642 = $signed(_T_56021) + $signed(_T_56026); // @[Modules.scala 143:103:@24354.4]
  assign _T_77643 = _T_77642[5:0]; // @[Modules.scala 143:103:@24355.4]
  assign _T_77644 = $signed(_T_77643); // @[Modules.scala 143:103:@24356.4]
  assign _T_77649 = $signed(_T_56028) + $signed(_T_62138); // @[Modules.scala 143:103:@24360.4]
  assign _T_77650 = _T_77649[4:0]; // @[Modules.scala 143:103:@24361.4]
  assign _T_77651 = $signed(_T_77650); // @[Modules.scala 143:103:@24362.4]
  assign _T_77670 = $signed(_GEN_68) + $signed(_T_59061); // @[Modules.scala 143:103:@24378.4]
  assign _T_77671 = _T_77670[5:0]; // @[Modules.scala 143:103:@24379.4]
  assign _T_77672 = $signed(_T_77671); // @[Modules.scala 143:103:@24380.4]
  assign _T_77677 = $signed(_T_71389) + $signed(_T_59075); // @[Modules.scala 143:103:@24384.4]
  assign _T_77678 = _T_77677[5:0]; // @[Modules.scala 143:103:@24385.4]
  assign _T_77679 = $signed(_T_77678); // @[Modules.scala 143:103:@24386.4]
  assign _T_77712 = $signed(_GEN_136) + $signed(_T_56103); // @[Modules.scala 143:103:@24414.4]
  assign _T_77713 = _T_77712[5:0]; // @[Modules.scala 143:103:@24415.4]
  assign _T_77714 = $signed(_T_77713); // @[Modules.scala 143:103:@24416.4]
  assign _T_77726 = $signed(_T_56112) + $signed(_GEN_354); // @[Modules.scala 143:103:@24426.4]
  assign _T_77727 = _T_77726[5:0]; // @[Modules.scala 143:103:@24427.4]
  assign _T_77728 = $signed(_T_77727); // @[Modules.scala 143:103:@24428.4]
  assign _T_77733 = $signed(_T_62215) + $signed(_T_56119); // @[Modules.scala 143:103:@24432.4]
  assign _T_77734 = _T_77733[4:0]; // @[Modules.scala 143:103:@24433.4]
  assign _T_77735 = $signed(_T_77734); // @[Modules.scala 143:103:@24434.4]
  assign _T_77740 = $signed(_T_56126) + $signed(_T_56133); // @[Modules.scala 143:103:@24438.4]
  assign _T_77741 = _T_77740[5:0]; // @[Modules.scala 143:103:@24439.4]
  assign _T_77742 = $signed(_T_77741); // @[Modules.scala 143:103:@24440.4]
  assign _GEN_558 = {{1{_T_65354[4]}},_T_65354}; // @[Modules.scala 143:103:@24444.4]
  assign _T_77747 = $signed(_T_56138) + $signed(_GEN_558); // @[Modules.scala 143:103:@24444.4]
  assign _T_77748 = _T_77747[5:0]; // @[Modules.scala 143:103:@24445.4]
  assign _T_77749 = $signed(_T_77748); // @[Modules.scala 143:103:@24446.4]
  assign _T_77789 = $signed(_T_59185) + $signed(_T_62273); // @[Modules.scala 143:103:@24480.4]
  assign _T_77790 = _T_77789[5:0]; // @[Modules.scala 143:103:@24481.4]
  assign _T_77791 = $signed(_T_77790); // @[Modules.scala 143:103:@24482.4]
  assign _T_77802 = $signed(-4'sh1) * $signed(io_in_734); // @[Modules.scala 144:80:@24491.4]
  assign _T_77803 = $signed(_T_59199) + $signed(_T_77802); // @[Modules.scala 143:103:@24492.4]
  assign _T_77804 = _T_77803[4:0]; // @[Modules.scala 143:103:@24493.4]
  assign _T_77805 = $signed(_T_77804); // @[Modules.scala 143:103:@24494.4]
  assign _GEN_559 = {{1{_T_62299[4]}},_T_62299}; // @[Modules.scala 143:103:@24504.4]
  assign _T_77817 = $signed(_GEN_559) + $signed(_T_56203); // @[Modules.scala 143:103:@24504.4]
  assign _T_77818 = _T_77817[5:0]; // @[Modules.scala 143:103:@24505.4]
  assign _T_77819 = $signed(_T_77818); // @[Modules.scala 143:103:@24506.4]
  assign _T_77838 = $signed(_T_59234) + $signed(_GEN_74); // @[Modules.scala 143:103:@24522.4]
  assign _T_77839 = _T_77838[5:0]; // @[Modules.scala 143:103:@24523.4]
  assign _T_77840 = $signed(_T_77839); // @[Modules.scala 143:103:@24524.4]
  assign _GEN_561 = {{1{_T_56236[4]}},_T_56236}; // @[Modules.scala 143:103:@24534.4]
  assign _T_77852 = $signed(_GEN_561) + $signed(_T_68500); // @[Modules.scala 143:103:@24534.4]
  assign _T_77853 = _T_77852[5:0]; // @[Modules.scala 143:103:@24535.4]
  assign _T_77854 = $signed(_T_77853); // @[Modules.scala 143:103:@24536.4]
  assign _GEN_562 = {{1{_T_62348[4]}},_T_62348}; // @[Modules.scala 143:103:@24540.4]
  assign _T_77859 = $signed(_T_68502) + $signed(_GEN_562); // @[Modules.scala 143:103:@24540.4]
  assign _T_77860 = _T_77859[5:0]; // @[Modules.scala 143:103:@24541.4]
  assign _T_77861 = $signed(_T_77860); // @[Modules.scala 143:103:@24542.4]
  assign _T_77866 = $signed(_GEN_278) + $signed(_T_56250); // @[Modules.scala 143:103:@24546.4]
  assign _T_77867 = _T_77866[5:0]; // @[Modules.scala 143:103:@24547.4]
  assign _T_77868 = $signed(_T_77867); // @[Modules.scala 143:103:@24548.4]
  assign _GEN_564 = {{1{_T_56257[4]}},_T_56257}; // @[Modules.scala 143:103:@24552.4]
  assign _T_77873 = $signed(_T_56252) + $signed(_GEN_564); // @[Modules.scala 143:103:@24552.4]
  assign _T_77874 = _T_77873[5:0]; // @[Modules.scala 143:103:@24553.4]
  assign _T_77875 = $signed(_T_77874); // @[Modules.scala 143:103:@24554.4]
  assign _T_77887 = $signed(_T_56271) + $signed(_T_71625); // @[Modules.scala 143:103:@24564.4]
  assign _T_77888 = _T_77887[5:0]; // @[Modules.scala 143:103:@24565.4]
  assign _T_77889 = $signed(_T_77888); // @[Modules.scala 143:103:@24566.4]
  assign _T_77915 = $signed(_T_59318) + $signed(_GEN_497); // @[Modules.scala 143:103:@24588.4]
  assign _T_77916 = _T_77915[5:0]; // @[Modules.scala 143:103:@24589.4]
  assign _T_77917 = $signed(_T_77916); // @[Modules.scala 143:103:@24590.4]
  assign _T_77922 = $signed(_T_56301) + $signed(_T_56306); // @[Modules.scala 143:103:@24594.4]
  assign _T_77923 = _T_77922[5:0]; // @[Modules.scala 143:103:@24595.4]
  assign _T_77924 = $signed(_T_77923); // @[Modules.scala 143:103:@24596.4]
  assign buffer_7_0 = {{9{_T_75768[4]}},_T_75768}; // @[Modules.scala 112:22:@8.4]
  assign _T_77925 = $signed(buffer_7_0) + $signed(buffer_0_0); // @[Modules.scala 166:64:@24598.4]
  assign _T_77926 = _T_77925[13:0]; // @[Modules.scala 166:64:@24599.4]
  assign buffer_7_309 = $signed(_T_77926); // @[Modules.scala 166:64:@24600.4]
  assign _T_77928 = $signed(buffer_0_1) + $signed(buffer_3_2); // @[Modules.scala 166:64:@24602.4]
  assign _T_77929 = _T_77928[13:0]; // @[Modules.scala 166:64:@24603.4]
  assign buffer_7_310 = $signed(_T_77929); // @[Modules.scala 166:64:@24604.4]
  assign buffer_7_4 = {{8{_T_75796[5]}},_T_75796}; // @[Modules.scala 112:22:@8.4]
  assign _T_77931 = $signed(buffer_7_4) + $signed(buffer_4_4); // @[Modules.scala 166:64:@24606.4]
  assign _T_77932 = _T_77931[13:0]; // @[Modules.scala 166:64:@24607.4]
  assign buffer_7_311 = $signed(_T_77932); // @[Modules.scala 166:64:@24608.4]
  assign _T_77934 = $signed(buffer_1_6) + $signed(buffer_6_8); // @[Modules.scala 166:64:@24610.4]
  assign _T_77935 = _T_77934[13:0]; // @[Modules.scala 166:64:@24611.4]
  assign buffer_7_312 = $signed(_T_77935); // @[Modules.scala 166:64:@24612.4]
  assign buffer_7_9 = {{9{_T_75831[4]}},_T_75831}; // @[Modules.scala 112:22:@8.4]
  assign _T_77937 = $signed(buffer_6_9) + $signed(buffer_7_9); // @[Modules.scala 166:64:@24614.4]
  assign _T_77938 = _T_77937[13:0]; // @[Modules.scala 166:64:@24615.4]
  assign buffer_7_313 = $signed(_T_77938); // @[Modules.scala 166:64:@24616.4]
  assign buffer_7_13 = {{8{_T_75859[5]}},_T_75859}; // @[Modules.scala 112:22:@8.4]
  assign _T_77943 = $signed(buffer_3_12) + $signed(buffer_7_13); // @[Modules.scala 166:64:@24622.4]
  assign _T_77944 = _T_77943[13:0]; // @[Modules.scala 166:64:@24623.4]
  assign buffer_7_315 = $signed(_T_77944); // @[Modules.scala 166:64:@24624.4]
  assign _T_77946 = $signed(buffer_4_13) + $signed(buffer_2_14); // @[Modules.scala 166:64:@24626.4]
  assign _T_77947 = _T_77946[13:0]; // @[Modules.scala 166:64:@24627.4]
  assign buffer_7_316 = $signed(_T_77947); // @[Modules.scala 166:64:@24628.4]
  assign _T_77949 = $signed(buffer_2_15) + $signed(buffer_2_16); // @[Modules.scala 166:64:@24630.4]
  assign _T_77950 = _T_77949[13:0]; // @[Modules.scala 166:64:@24631.4]
  assign buffer_7_317 = $signed(_T_77950); // @[Modules.scala 166:64:@24632.4]
  assign _T_77952 = $signed(buffer_3_17) + $signed(buffer_6_20); // @[Modules.scala 166:64:@24634.4]
  assign _T_77953 = _T_77952[13:0]; // @[Modules.scala 166:64:@24635.4]
  assign buffer_7_318 = $signed(_T_77953); // @[Modules.scala 166:64:@24636.4]
  assign buffer_7_20 = {{8{_T_75908[5]}},_T_75908}; // @[Modules.scala 112:22:@8.4]
  assign _T_77955 = $signed(buffer_7_20) + $signed(buffer_1_21); // @[Modules.scala 166:64:@24638.4]
  assign _T_77956 = _T_77955[13:0]; // @[Modules.scala 166:64:@24639.4]
  assign buffer_7_319 = $signed(_T_77956); // @[Modules.scala 166:64:@24640.4]
  assign buffer_7_22 = {{8{_T_75922[5]}},_T_75922}; // @[Modules.scala 112:22:@8.4]
  assign _T_77958 = $signed(buffer_7_22) + $signed(buffer_1_23); // @[Modules.scala 166:64:@24642.4]
  assign _T_77959 = _T_77958[13:0]; // @[Modules.scala 166:64:@24643.4]
  assign buffer_7_320 = $signed(_T_77959); // @[Modules.scala 166:64:@24644.4]
  assign buffer_7_24 = {{8{_T_75936[5]}},_T_75936}; // @[Modules.scala 112:22:@8.4]
  assign _T_77961 = $signed(buffer_7_24) + $signed(buffer_1_25); // @[Modules.scala 166:64:@24646.4]
  assign _T_77962 = _T_77961[13:0]; // @[Modules.scala 166:64:@24647.4]
  assign buffer_7_321 = $signed(_T_77962); // @[Modules.scala 166:64:@24648.4]
  assign _T_77967 = $signed(buffer_5_27) + $signed(buffer_5_28); // @[Modules.scala 166:64:@24654.4]
  assign _T_77968 = _T_77967[13:0]; // @[Modules.scala 166:64:@24655.4]
  assign buffer_7_323 = $signed(_T_77968); // @[Modules.scala 166:64:@24656.4]
  assign _T_77970 = $signed(buffer_1_29) + $signed(buffer_1_30); // @[Modules.scala 166:64:@24658.4]
  assign _T_77971 = _T_77970[13:0]; // @[Modules.scala 166:64:@24659.4]
  assign buffer_7_324 = $signed(_T_77971); // @[Modules.scala 166:64:@24660.4]
  assign buffer_7_33 = {{8{_T_75999[5]}},_T_75999}; // @[Modules.scala 112:22:@8.4]
  assign _T_77973 = $signed(buffer_1_31) + $signed(buffer_7_33); // @[Modules.scala 166:64:@24662.4]
  assign _T_77974 = _T_77973[13:0]; // @[Modules.scala 166:64:@24663.4]
  assign buffer_7_325 = $signed(_T_77974); // @[Modules.scala 166:64:@24664.4]
  assign buffer_7_35 = {{8{_T_76013[5]}},_T_76013}; // @[Modules.scala 112:22:@8.4]
  assign _T_77976 = $signed(buffer_6_33) + $signed(buffer_7_35); // @[Modules.scala 166:64:@24666.4]
  assign _T_77977 = _T_77976[13:0]; // @[Modules.scala 166:64:@24667.4]
  assign buffer_7_326 = $signed(_T_77977); // @[Modules.scala 166:64:@24668.4]
  assign _T_77979 = $signed(buffer_3_35) + $signed(buffer_3_36); // @[Modules.scala 166:64:@24670.4]
  assign _T_77980 = _T_77979[13:0]; // @[Modules.scala 166:64:@24671.4]
  assign buffer_7_327 = $signed(_T_77980); // @[Modules.scala 166:64:@24672.4]
  assign buffer_7_38 = {{8{_T_76034[5]}},_T_76034}; // @[Modules.scala 112:22:@8.4]
  assign _T_77982 = $signed(buffer_7_38) + $signed(buffer_0_39); // @[Modules.scala 166:64:@24674.4]
  assign _T_77983 = _T_77982[13:0]; // @[Modules.scala 166:64:@24675.4]
  assign buffer_7_328 = $signed(_T_77983); // @[Modules.scala 166:64:@24676.4]
  assign buffer_7_40 = {{9{_T_76048[4]}},_T_76048}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_41 = {{9{_T_76055[4]}},_T_76055}; // @[Modules.scala 112:22:@8.4]
  assign _T_77985 = $signed(buffer_7_40) + $signed(buffer_7_41); // @[Modules.scala 166:64:@24678.4]
  assign _T_77986 = _T_77985[13:0]; // @[Modules.scala 166:64:@24679.4]
  assign buffer_7_329 = $signed(_T_77986); // @[Modules.scala 166:64:@24680.4]
  assign buffer_7_42 = {{9{_T_76062[4]}},_T_76062}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_43 = {{8{_T_76069[5]}},_T_76069}; // @[Modules.scala 112:22:@8.4]
  assign _T_77988 = $signed(buffer_7_42) + $signed(buffer_7_43); // @[Modules.scala 166:64:@24682.4]
  assign _T_77989 = _T_77988[13:0]; // @[Modules.scala 166:64:@24683.4]
  assign buffer_7_330 = $signed(_T_77989); // @[Modules.scala 166:64:@24684.4]
  assign buffer_7_45 = {{8{_T_76083[5]}},_T_76083}; // @[Modules.scala 112:22:@8.4]
  assign _T_77991 = $signed(buffer_1_43) + $signed(buffer_7_45); // @[Modules.scala 166:64:@24686.4]
  assign _T_77992 = _T_77991[13:0]; // @[Modules.scala 166:64:@24687.4]
  assign buffer_7_331 = $signed(_T_77992); // @[Modules.scala 166:64:@24688.4]
  assign buffer_7_49 = {{8{_T_76111[5]}},_T_76111}; // @[Modules.scala 112:22:@8.4]
  assign _T_77997 = $signed(buffer_0_47) + $signed(buffer_7_49); // @[Modules.scala 166:64:@24694.4]
  assign _T_77998 = _T_77997[13:0]; // @[Modules.scala 166:64:@24695.4]
  assign buffer_7_333 = $signed(_T_77998); // @[Modules.scala 166:64:@24696.4]
  assign buffer_7_51 = {{8{_T_76125[5]}},_T_76125}; // @[Modules.scala 112:22:@8.4]
  assign _T_78000 = $signed(buffer_5_50) + $signed(buffer_7_51); // @[Modules.scala 166:64:@24698.4]
  assign _T_78001 = _T_78000[13:0]; // @[Modules.scala 166:64:@24699.4]
  assign buffer_7_334 = $signed(_T_78001); // @[Modules.scala 166:64:@24700.4]
  assign buffer_7_52 = {{8{_T_76132[5]}},_T_76132}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_53 = {{8{_T_76139[5]}},_T_76139}; // @[Modules.scala 112:22:@8.4]
  assign _T_78003 = $signed(buffer_7_52) + $signed(buffer_7_53); // @[Modules.scala 166:64:@24702.4]
  assign _T_78004 = _T_78003[13:0]; // @[Modules.scala 166:64:@24703.4]
  assign buffer_7_335 = $signed(_T_78004); // @[Modules.scala 166:64:@24704.4]
  assign buffer_7_54 = {{8{_T_76146[5]}},_T_76146}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_55 = {{8{_T_76153[5]}},_T_76153}; // @[Modules.scala 112:22:@8.4]
  assign _T_78006 = $signed(buffer_7_54) + $signed(buffer_7_55); // @[Modules.scala 166:64:@24706.4]
  assign _T_78007 = _T_78006[13:0]; // @[Modules.scala 166:64:@24707.4]
  assign buffer_7_336 = $signed(_T_78007); // @[Modules.scala 166:64:@24708.4]
  assign buffer_7_57 = {{8{_T_76167[5]}},_T_76167}; // @[Modules.scala 112:22:@8.4]
  assign _T_78009 = $signed(buffer_3_58) + $signed(buffer_7_57); // @[Modules.scala 166:64:@24710.4]
  assign _T_78010 = _T_78009[13:0]; // @[Modules.scala 166:64:@24711.4]
  assign buffer_7_337 = $signed(_T_78010); // @[Modules.scala 166:64:@24712.4]
  assign _T_78012 = $signed(buffer_6_58) + $signed(buffer_3_62); // @[Modules.scala 166:64:@24714.4]
  assign _T_78013 = _T_78012[13:0]; // @[Modules.scala 166:64:@24715.4]
  assign buffer_7_338 = $signed(_T_78013); // @[Modules.scala 166:64:@24716.4]
  assign buffer_7_60 = {{9{_T_76188[4]}},_T_76188}; // @[Modules.scala 112:22:@8.4]
  assign _T_78015 = $signed(buffer_7_60) + $signed(buffer_2_60); // @[Modules.scala 166:64:@24718.4]
  assign _T_78016 = _T_78015[13:0]; // @[Modules.scala 166:64:@24719.4]
  assign buffer_7_339 = $signed(_T_78016); // @[Modules.scala 166:64:@24720.4]
  assign buffer_7_63 = {{8{_T_76209[5]}},_T_76209}; // @[Modules.scala 112:22:@8.4]
  assign _T_78018 = $signed(buffer_2_61) + $signed(buffer_7_63); // @[Modules.scala 166:64:@24722.4]
  assign _T_78019 = _T_78018[13:0]; // @[Modules.scala 166:64:@24723.4]
  assign buffer_7_340 = $signed(_T_78019); // @[Modules.scala 166:64:@24724.4]
  assign _T_78021 = $signed(buffer_3_67) + $signed(buffer_3_68); // @[Modules.scala 166:64:@24726.4]
  assign _T_78022 = _T_78021[13:0]; // @[Modules.scala 166:64:@24727.4]
  assign buffer_7_341 = $signed(_T_78022); // @[Modules.scala 166:64:@24728.4]
  assign buffer_7_66 = {{8{_T_76230[5]}},_T_76230}; // @[Modules.scala 112:22:@8.4]
  assign _T_78024 = $signed(buffer_7_66) + $signed(buffer_6_67); // @[Modules.scala 166:64:@24730.4]
  assign _T_78025 = _T_78024[13:0]; // @[Modules.scala 166:64:@24731.4]
  assign buffer_7_342 = $signed(_T_78025); // @[Modules.scala 166:64:@24732.4]
  assign buffer_7_68 = {{8{_T_76244[5]}},_T_76244}; // @[Modules.scala 112:22:@8.4]
  assign _T_78027 = $signed(buffer_7_68) + $signed(buffer_6_70); // @[Modules.scala 166:64:@24734.4]
  assign _T_78028 = _T_78027[13:0]; // @[Modules.scala 166:64:@24735.4]
  assign buffer_7_343 = $signed(_T_78028); // @[Modules.scala 166:64:@24736.4]
  assign _T_78030 = $signed(buffer_5_72) + $signed(buffer_2_72); // @[Modules.scala 166:64:@24738.4]
  assign _T_78031 = _T_78030[13:0]; // @[Modules.scala 166:64:@24739.4]
  assign buffer_7_344 = $signed(_T_78031); // @[Modules.scala 166:64:@24740.4]
  assign _T_78033 = $signed(buffer_2_73) + $signed(buffer_0_71); // @[Modules.scala 166:64:@24742.4]
  assign _T_78034 = _T_78033[13:0]; // @[Modules.scala 166:64:@24743.4]
  assign buffer_7_345 = $signed(_T_78034); // @[Modules.scala 166:64:@24744.4]
  assign buffer_7_74 = {{8{_T_76286[5]}},_T_76286}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_75 = {{8{_T_76293[5]}},_T_76293}; // @[Modules.scala 112:22:@8.4]
  assign _T_78036 = $signed(buffer_7_74) + $signed(buffer_7_75); // @[Modules.scala 166:64:@24746.4]
  assign _T_78037 = _T_78036[13:0]; // @[Modules.scala 166:64:@24747.4]
  assign buffer_7_346 = $signed(_T_78037); // @[Modules.scala 166:64:@24748.4]
  assign buffer_7_76 = {{8{_T_76300[5]}},_T_76300}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_77 = {{8{_T_76307[5]}},_T_76307}; // @[Modules.scala 112:22:@8.4]
  assign _T_78039 = $signed(buffer_7_76) + $signed(buffer_7_77); // @[Modules.scala 166:64:@24750.4]
  assign _T_78040 = _T_78039[13:0]; // @[Modules.scala 166:64:@24751.4]
  assign buffer_7_347 = $signed(_T_78040); // @[Modules.scala 166:64:@24752.4]
  assign buffer_7_82 = {{8{_T_76342[5]}},_T_76342}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_83 = {{8{_T_76349[5]}},_T_76349}; // @[Modules.scala 112:22:@8.4]
  assign _T_78048 = $signed(buffer_7_82) + $signed(buffer_7_83); // @[Modules.scala 166:64:@24762.4]
  assign _T_78049 = _T_78048[13:0]; // @[Modules.scala 166:64:@24763.4]
  assign buffer_7_350 = $signed(_T_78049); // @[Modules.scala 166:64:@24764.4]
  assign buffer_7_84 = {{8{_T_76356[5]}},_T_76356}; // @[Modules.scala 112:22:@8.4]
  assign _T_78051 = $signed(buffer_7_84) + $signed(buffer_2_86); // @[Modules.scala 166:64:@24766.4]
  assign _T_78052 = _T_78051[13:0]; // @[Modules.scala 166:64:@24767.4]
  assign buffer_7_351 = $signed(_T_78052); // @[Modules.scala 166:64:@24768.4]
  assign buffer_7_86 = {{8{_T_76370[5]}},_T_76370}; // @[Modules.scala 112:22:@8.4]
  assign _T_78054 = $signed(buffer_7_86) + $signed(buffer_5_90); // @[Modules.scala 166:64:@24770.4]
  assign _T_78055 = _T_78054[13:0]; // @[Modules.scala 166:64:@24771.4]
  assign buffer_7_352 = $signed(_T_78055); // @[Modules.scala 166:64:@24772.4]
  assign _T_78057 = $signed(buffer_5_91) + $signed(buffer_5_92); // @[Modules.scala 166:64:@24774.4]
  assign _T_78058 = _T_78057[13:0]; // @[Modules.scala 166:64:@24775.4]
  assign buffer_7_353 = $signed(_T_78058); // @[Modules.scala 166:64:@24776.4]
  assign _T_78060 = $signed(buffer_5_93) + $signed(buffer_0_88); // @[Modules.scala 166:64:@24778.4]
  assign _T_78061 = _T_78060[13:0]; // @[Modules.scala 166:64:@24779.4]
  assign buffer_7_354 = $signed(_T_78061); // @[Modules.scala 166:64:@24780.4]
  assign _T_78063 = $signed(buffer_5_95) + $signed(buffer_5_96); // @[Modules.scala 166:64:@24782.4]
  assign _T_78064 = _T_78063[13:0]; // @[Modules.scala 166:64:@24783.4]
  assign buffer_7_355 = $signed(_T_78064); // @[Modules.scala 166:64:@24784.4]
  assign _T_78066 = $signed(buffer_5_97) + $signed(buffer_5_98); // @[Modules.scala 166:64:@24786.4]
  assign _T_78067 = _T_78066[13:0]; // @[Modules.scala 166:64:@24787.4]
  assign buffer_7_356 = $signed(_T_78067); // @[Modules.scala 166:64:@24788.4]
  assign _T_78069 = $signed(buffer_4_93) + $signed(buffer_4_94); // @[Modules.scala 166:64:@24790.4]
  assign _T_78070 = _T_78069[13:0]; // @[Modules.scala 166:64:@24791.4]
  assign buffer_7_357 = $signed(_T_78070); // @[Modules.scala 166:64:@24792.4]
  assign buffer_7_100 = {{8{_T_76468[5]}},_T_76468}; // @[Modules.scala 112:22:@8.4]
  assign _T_78075 = $signed(buffer_7_100) + $signed(buffer_3_103); // @[Modules.scala 166:64:@24798.4]
  assign _T_78076 = _T_78075[13:0]; // @[Modules.scala 166:64:@24799.4]
  assign buffer_7_359 = $signed(_T_78076); // @[Modules.scala 166:64:@24800.4]
  assign _T_78078 = $signed(buffer_3_104) + $signed(buffer_1_102); // @[Modules.scala 166:64:@24802.4]
  assign _T_78079 = _T_78078[13:0]; // @[Modules.scala 166:64:@24803.4]
  assign buffer_7_360 = $signed(_T_78079); // @[Modules.scala 166:64:@24804.4]
  assign _T_78081 = $signed(buffer_0_100) + $signed(buffer_1_104); // @[Modules.scala 166:64:@24806.4]
  assign _T_78082 = _T_78081[13:0]; // @[Modules.scala 166:64:@24807.4]
  assign buffer_7_361 = $signed(_T_78082); // @[Modules.scala 166:64:@24808.4]
  assign _T_78084 = $signed(buffer_6_105) + $signed(buffer_3_109); // @[Modules.scala 166:64:@24810.4]
  assign _T_78085 = _T_78084[13:0]; // @[Modules.scala 166:64:@24811.4]
  assign buffer_7_362 = $signed(_T_78085); // @[Modules.scala 166:64:@24812.4]
  assign buffer_7_112 = {{8{_T_76552[5]}},_T_76552}; // @[Modules.scala 112:22:@8.4]
  assign _T_78093 = $signed(buffer_7_112) + $signed(buffer_1_112); // @[Modules.scala 166:64:@24822.4]
  assign _T_78094 = _T_78093[13:0]; // @[Modules.scala 166:64:@24823.4]
  assign buffer_7_365 = $signed(_T_78094); // @[Modules.scala 166:64:@24824.4]
  assign buffer_7_115 = {{8{_T_76573[5]}},_T_76573}; // @[Modules.scala 112:22:@8.4]
  assign _T_78096 = $signed(buffer_5_117) + $signed(buffer_7_115); // @[Modules.scala 166:64:@24826.4]
  assign _T_78097 = _T_78096[13:0]; // @[Modules.scala 166:64:@24827.4]
  assign buffer_7_366 = $signed(_T_78097); // @[Modules.scala 166:64:@24828.4]
  assign _T_78099 = $signed(buffer_1_116) + $signed(buffer_4_115); // @[Modules.scala 166:64:@24830.4]
  assign _T_78100 = _T_78099[13:0]; // @[Modules.scala 166:64:@24831.4]
  assign buffer_7_367 = $signed(_T_78100); // @[Modules.scala 166:64:@24832.4]
  assign _T_78102 = $signed(buffer_2_119) + $signed(buffer_1_119); // @[Modules.scala 166:64:@24834.4]
  assign _T_78103 = _T_78102[13:0]; // @[Modules.scala 166:64:@24835.4]
  assign buffer_7_368 = $signed(_T_78103); // @[Modules.scala 166:64:@24836.4]
  assign buffer_7_120 = {{8{_T_76608[5]}},_T_76608}; // @[Modules.scala 112:22:@8.4]
  assign _T_78105 = $signed(buffer_7_120) + $signed(buffer_1_121); // @[Modules.scala 166:64:@24838.4]
  assign _T_78106 = _T_78105[13:0]; // @[Modules.scala 166:64:@24839.4]
  assign buffer_7_369 = $signed(_T_78106); // @[Modules.scala 166:64:@24840.4]
  assign _T_78108 = $signed(buffer_0_120) + $signed(buffer_0_122); // @[Modules.scala 166:64:@24842.4]
  assign _T_78109 = _T_78108[13:0]; // @[Modules.scala 166:64:@24843.4]
  assign buffer_7_370 = $signed(_T_78109); // @[Modules.scala 166:64:@24844.4]
  assign buffer_7_125 = {{8{_T_76643[5]}},_T_76643}; // @[Modules.scala 112:22:@8.4]
  assign _T_78111 = $signed(buffer_0_123) + $signed(buffer_7_125); // @[Modules.scala 166:64:@24846.4]
  assign _T_78112 = _T_78111[13:0]; // @[Modules.scala 166:64:@24847.4]
  assign buffer_7_371 = $signed(_T_78112); // @[Modules.scala 166:64:@24848.4]
  assign buffer_7_126 = {{8{_T_76650[5]}},_T_76650}; // @[Modules.scala 112:22:@8.4]
  assign _T_78114 = $signed(buffer_7_126) + $signed(buffer_0_125); // @[Modules.scala 166:64:@24850.4]
  assign _T_78115 = _T_78114[13:0]; // @[Modules.scala 166:64:@24851.4]
  assign buffer_7_372 = $signed(_T_78115); // @[Modules.scala 166:64:@24852.4]
  assign buffer_7_129 = {{8{_T_76671[5]}},_T_76671}; // @[Modules.scala 112:22:@8.4]
  assign _T_78117 = $signed(buffer_0_126) + $signed(buffer_7_129); // @[Modules.scala 166:64:@24854.4]
  assign _T_78118 = _T_78117[13:0]; // @[Modules.scala 166:64:@24855.4]
  assign buffer_7_373 = $signed(_T_78118); // @[Modules.scala 166:64:@24856.4]
  assign buffer_7_133 = {{9{_T_76699[4]}},_T_76699}; // @[Modules.scala 112:22:@8.4]
  assign _T_78123 = $signed(buffer_5_135) + $signed(buffer_7_133); // @[Modules.scala 166:64:@24862.4]
  assign _T_78124 = _T_78123[13:0]; // @[Modules.scala 166:64:@24863.4]
  assign buffer_7_375 = $signed(_T_78124); // @[Modules.scala 166:64:@24864.4]
  assign _T_78126 = $signed(buffer_0_135) + $signed(buffer_6_140); // @[Modules.scala 166:64:@24866.4]
  assign _T_78127 = _T_78126[13:0]; // @[Modules.scala 166:64:@24867.4]
  assign buffer_7_376 = $signed(_T_78127); // @[Modules.scala 166:64:@24868.4]
  assign _T_78129 = $signed(buffer_6_141) + $signed(buffer_0_138); // @[Modules.scala 166:64:@24870.4]
  assign _T_78130 = _T_78129[13:0]; // @[Modules.scala 166:64:@24871.4]
  assign buffer_7_377 = $signed(_T_78130); // @[Modules.scala 166:64:@24872.4]
  assign _T_78132 = $signed(buffer_0_139) + $signed(buffer_6_144); // @[Modules.scala 166:64:@24874.4]
  assign _T_78133 = _T_78132[13:0]; // @[Modules.scala 166:64:@24875.4]
  assign buffer_7_378 = $signed(_T_78133); // @[Modules.scala 166:64:@24876.4]
  assign _T_78135 = $signed(buffer_0_141) + $signed(buffer_0_142); // @[Modules.scala 166:64:@24878.4]
  assign _T_78136 = _T_78135[13:0]; // @[Modules.scala 166:64:@24879.4]
  assign buffer_7_379 = $signed(_T_78136); // @[Modules.scala 166:64:@24880.4]
  assign _T_78138 = $signed(buffer_0_143) + $signed(buffer_0_144); // @[Modules.scala 166:64:@24882.4]
  assign _T_78139 = _T_78138[13:0]; // @[Modules.scala 166:64:@24883.4]
  assign buffer_7_380 = $signed(_T_78139); // @[Modules.scala 166:64:@24884.4]
  assign buffer_7_145 = {{9{_T_76783[4]}},_T_76783}; // @[Modules.scala 112:22:@8.4]
  assign _T_78141 = $signed(buffer_6_149) + $signed(buffer_7_145); // @[Modules.scala 166:64:@24886.4]
  assign _T_78142 = _T_78141[13:0]; // @[Modules.scala 166:64:@24887.4]
  assign buffer_7_381 = $signed(_T_78142); // @[Modules.scala 166:64:@24888.4]
  assign buffer_7_146 = {{9{_T_76790[4]}},_T_76790}; // @[Modules.scala 112:22:@8.4]
  assign _T_78144 = $signed(buffer_7_146) + $signed(buffer_1_149); // @[Modules.scala 166:64:@24890.4]
  assign _T_78145 = _T_78144[13:0]; // @[Modules.scala 166:64:@24891.4]
  assign buffer_7_382 = $signed(_T_78145); // @[Modules.scala 166:64:@24892.4]
  assign buffer_7_149 = {{8{_T_76811[5]}},_T_76811}; // @[Modules.scala 112:22:@8.4]
  assign _T_78147 = $signed(buffer_1_150) + $signed(buffer_7_149); // @[Modules.scala 166:64:@24894.4]
  assign _T_78148 = _T_78147[13:0]; // @[Modules.scala 166:64:@24895.4]
  assign buffer_7_383 = $signed(_T_78148); // @[Modules.scala 166:64:@24896.4]
  assign buffer_7_150 = {{8{_T_76818[5]}},_T_76818}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_151 = {{8{_T_76825[5]}},_T_76825}; // @[Modules.scala 112:22:@8.4]
  assign _T_78150 = $signed(buffer_7_150) + $signed(buffer_7_151); // @[Modules.scala 166:64:@24898.4]
  assign _T_78151 = _T_78150[13:0]; // @[Modules.scala 166:64:@24899.4]
  assign buffer_7_384 = $signed(_T_78151); // @[Modules.scala 166:64:@24900.4]
  assign buffer_7_152 = {{8{_T_76832[5]}},_T_76832}; // @[Modules.scala 112:22:@8.4]
  assign _T_78153 = $signed(buffer_7_152) + $signed(buffer_5_153); // @[Modules.scala 166:64:@24902.4]
  assign _T_78154 = _T_78153[13:0]; // @[Modules.scala 166:64:@24903.4]
  assign buffer_7_385 = $signed(_T_78154); // @[Modules.scala 166:64:@24904.4]
  assign buffer_7_157 = {{8{_T_76867[5]}},_T_76867}; // @[Modules.scala 112:22:@8.4]
  assign _T_78159 = $signed(buffer_1_156) + $signed(buffer_7_157); // @[Modules.scala 166:64:@24910.4]
  assign _T_78160 = _T_78159[13:0]; // @[Modules.scala 166:64:@24911.4]
  assign buffer_7_387 = $signed(_T_78160); // @[Modules.scala 166:64:@24912.4]
  assign buffer_7_158 = {{9{_T_76874[4]}},_T_76874}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_159 = {{9{_T_76881[4]}},_T_76881}; // @[Modules.scala 112:22:@8.4]
  assign _T_78162 = $signed(buffer_7_158) + $signed(buffer_7_159); // @[Modules.scala 166:64:@24914.4]
  assign _T_78163 = _T_78162[13:0]; // @[Modules.scala 166:64:@24915.4]
  assign buffer_7_388 = $signed(_T_78163); // @[Modules.scala 166:64:@24916.4]
  assign _T_78165 = $signed(buffer_6_165) + $signed(buffer_5_161); // @[Modules.scala 166:64:@24918.4]
  assign _T_78166 = _T_78165[13:0]; // @[Modules.scala 166:64:@24919.4]
  assign buffer_7_389 = $signed(_T_78166); // @[Modules.scala 166:64:@24920.4]
  assign buffer_7_162 = {{9{_T_76902[4]}},_T_76902}; // @[Modules.scala 112:22:@8.4]
  assign _T_78168 = $signed(buffer_7_162) + $signed(buffer_5_163); // @[Modules.scala 166:64:@24922.4]
  assign _T_78169 = _T_78168[13:0]; // @[Modules.scala 166:64:@24923.4]
  assign buffer_7_390 = $signed(_T_78169); // @[Modules.scala 166:64:@24924.4]
  assign buffer_7_164 = {{9{_T_76916[4]}},_T_76916}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_165 = {{9{_T_76923[4]}},_T_76923}; // @[Modules.scala 112:22:@8.4]
  assign _T_78171 = $signed(buffer_7_164) + $signed(buffer_7_165); // @[Modules.scala 166:64:@24926.4]
  assign _T_78172 = _T_78171[13:0]; // @[Modules.scala 166:64:@24927.4]
  assign buffer_7_391 = $signed(_T_78172); // @[Modules.scala 166:64:@24928.4]
  assign _T_78174 = $signed(buffer_0_164) + $signed(buffer_1_166); // @[Modules.scala 166:64:@24930.4]
  assign _T_78175 = _T_78174[13:0]; // @[Modules.scala 166:64:@24931.4]
  assign buffer_7_392 = $signed(_T_78175); // @[Modules.scala 166:64:@24932.4]
  assign buffer_7_168 = {{9{_T_76944[4]}},_T_76944}; // @[Modules.scala 112:22:@8.4]
  assign _T_78177 = $signed(buffer_7_168) + $signed(buffer_4_163); // @[Modules.scala 166:64:@24934.4]
  assign _T_78178 = _T_78177[13:0]; // @[Modules.scala 166:64:@24935.4]
  assign buffer_7_393 = $signed(_T_78178); // @[Modules.scala 166:64:@24936.4]
  assign buffer_7_171 = {{9{_T_76965[4]}},_T_76965}; // @[Modules.scala 112:22:@8.4]
  assign _T_78180 = $signed(buffer_0_167) + $signed(buffer_7_171); // @[Modules.scala 166:64:@24938.4]
  assign _T_78181 = _T_78180[13:0]; // @[Modules.scala 166:64:@24939.4]
  assign buffer_7_394 = $signed(_T_78181); // @[Modules.scala 166:64:@24940.4]
  assign _T_78183 = $signed(buffer_3_175) + $signed(buffer_3_176); // @[Modules.scala 166:64:@24942.4]
  assign _T_78184 = _T_78183[13:0]; // @[Modules.scala 166:64:@24943.4]
  assign buffer_7_395 = $signed(_T_78184); // @[Modules.scala 166:64:@24944.4]
  assign _T_78186 = $signed(buffer_3_177) + $signed(buffer_1_171); // @[Modules.scala 166:64:@24946.4]
  assign _T_78187 = _T_78186[13:0]; // @[Modules.scala 166:64:@24947.4]
  assign buffer_7_396 = $signed(_T_78187); // @[Modules.scala 166:64:@24948.4]
  assign buffer_7_176 = {{8{_T_77000[5]}},_T_77000}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_177 = {{8{_T_77007[5]}},_T_77007}; // @[Modules.scala 112:22:@8.4]
  assign _T_78189 = $signed(buffer_7_176) + $signed(buffer_7_177); // @[Modules.scala 166:64:@24950.4]
  assign _T_78190 = _T_78189[13:0]; // @[Modules.scala 166:64:@24951.4]
  assign buffer_7_397 = $signed(_T_78190); // @[Modules.scala 166:64:@24952.4]
  assign _T_78192 = $signed(buffer_3_181) + $signed(buffer_3_182); // @[Modules.scala 166:64:@24954.4]
  assign _T_78193 = _T_78192[13:0]; // @[Modules.scala 166:64:@24955.4]
  assign buffer_7_398 = $signed(_T_78193); // @[Modules.scala 166:64:@24956.4]
  assign _T_78198 = $signed(buffer_1_178) + $signed(buffer_5_180); // @[Modules.scala 166:64:@24962.4]
  assign _T_78199 = _T_78198[13:0]; // @[Modules.scala 166:64:@24963.4]
  assign buffer_7_400 = $signed(_T_78199); // @[Modules.scala 166:64:@24964.4]
  assign _T_78201 = $signed(buffer_0_179) + $signed(buffer_0_180); // @[Modules.scala 166:64:@24966.4]
  assign _T_78202 = _T_78201[13:0]; // @[Modules.scala 166:64:@24967.4]
  assign buffer_7_401 = $signed(_T_78202); // @[Modules.scala 166:64:@24968.4]
  assign _T_78204 = $signed(buffer_3_189) + $signed(buffer_3_190); // @[Modules.scala 166:64:@24970.4]
  assign _T_78205 = _T_78204[13:0]; // @[Modules.scala 166:64:@24971.4]
  assign buffer_7_402 = $signed(_T_78205); // @[Modules.scala 166:64:@24972.4]
  assign buffer_7_189 = {{8{_T_77091[5]}},_T_77091}; // @[Modules.scala 112:22:@8.4]
  assign _T_78207 = $signed(buffer_2_188) + $signed(buffer_7_189); // @[Modules.scala 166:64:@24974.4]
  assign _T_78208 = _T_78207[13:0]; // @[Modules.scala 166:64:@24975.4]
  assign buffer_7_403 = $signed(_T_78208); // @[Modules.scala 166:64:@24976.4]
  assign buffer_7_191 = {{9{_T_77105[4]}},_T_77105}; // @[Modules.scala 112:22:@8.4]
  assign _T_78210 = $signed(buffer_1_184) + $signed(buffer_7_191); // @[Modules.scala 166:64:@24978.4]
  assign _T_78211 = _T_78210[13:0]; // @[Modules.scala 166:64:@24979.4]
  assign buffer_7_404 = $signed(_T_78211); // @[Modules.scala 166:64:@24980.4]
  assign _T_78213 = $signed(buffer_3_195) + $signed(buffer_1_187); // @[Modules.scala 166:64:@24982.4]
  assign _T_78214 = _T_78213[13:0]; // @[Modules.scala 166:64:@24983.4]
  assign buffer_7_405 = $signed(_T_78214); // @[Modules.scala 166:64:@24984.4]
  assign _T_78216 = $signed(buffer_1_188) + $signed(buffer_0_187); // @[Modules.scala 166:64:@24986.4]
  assign _T_78217 = _T_78216[13:0]; // @[Modules.scala 166:64:@24987.4]
  assign buffer_7_406 = $signed(_T_78217); // @[Modules.scala 166:64:@24988.4]
  assign buffer_7_198 = {{9{_T_77154[4]}},_T_77154}; // @[Modules.scala 112:22:@8.4]
  assign _T_78222 = $signed(buffer_7_198) + $signed(buffer_1_193); // @[Modules.scala 166:64:@24994.4]
  assign _T_78223 = _T_78222[13:0]; // @[Modules.scala 166:64:@24995.4]
  assign buffer_7_408 = $signed(_T_78223); // @[Modules.scala 166:64:@24996.4]
  assign buffer_7_200 = {{9{_T_77168[4]}},_T_77168}; // @[Modules.scala 112:22:@8.4]
  assign _T_78225 = $signed(buffer_7_200) + $signed(buffer_2_198); // @[Modules.scala 166:64:@24998.4]
  assign _T_78226 = _T_78225[13:0]; // @[Modules.scala 166:64:@24999.4]
  assign buffer_7_409 = $signed(_T_78226); // @[Modules.scala 166:64:@25000.4]
  assign buffer_7_203 = {{8{_T_77189[5]}},_T_77189}; // @[Modules.scala 112:22:@8.4]
  assign _T_78228 = $signed(buffer_0_193) + $signed(buffer_7_203); // @[Modules.scala 166:64:@25002.4]
  assign _T_78229 = _T_78228[13:0]; // @[Modules.scala 166:64:@25003.4]
  assign buffer_7_410 = $signed(_T_78229); // @[Modules.scala 166:64:@25004.4]
  assign buffer_7_204 = {{9{_T_77196[4]}},_T_77196}; // @[Modules.scala 112:22:@8.4]
  assign _T_78231 = $signed(buffer_7_204) + $signed(buffer_2_202); // @[Modules.scala 166:64:@25006.4]
  assign _T_78232 = _T_78231[13:0]; // @[Modules.scala 166:64:@25007.4]
  assign buffer_7_411 = $signed(_T_78232); // @[Modules.scala 166:64:@25008.4]
  assign buffer_7_207 = {{8{_T_77217[5]}},_T_77217}; // @[Modules.scala 112:22:@8.4]
  assign _T_78234 = $signed(buffer_1_199) + $signed(buffer_7_207); // @[Modules.scala 166:64:@25010.4]
  assign _T_78235 = _T_78234[13:0]; // @[Modules.scala 166:64:@25011.4]
  assign buffer_7_412 = $signed(_T_78235); // @[Modules.scala 166:64:@25012.4]
  assign buffer_7_208 = {{8{_T_77224[5]}},_T_77224}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_209 = {{8{_T_77231[5]}},_T_77231}; // @[Modules.scala 112:22:@8.4]
  assign _T_78237 = $signed(buffer_7_208) + $signed(buffer_7_209); // @[Modules.scala 166:64:@25014.4]
  assign _T_78238 = _T_78237[13:0]; // @[Modules.scala 166:64:@25015.4]
  assign buffer_7_413 = $signed(_T_78238); // @[Modules.scala 166:64:@25016.4]
  assign buffer_7_211 = {{9{_T_77245[4]}},_T_77245}; // @[Modules.scala 112:22:@8.4]
  assign _T_78240 = $signed(buffer_1_203) + $signed(buffer_7_211); // @[Modules.scala 166:64:@25018.4]
  assign _T_78241 = _T_78240[13:0]; // @[Modules.scala 166:64:@25019.4]
  assign buffer_7_414 = $signed(_T_78241); // @[Modules.scala 166:64:@25020.4]
  assign buffer_7_212 = {{8{_T_77252[5]}},_T_77252}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_213 = {{9{_T_77259[4]}},_T_77259}; // @[Modules.scala 112:22:@8.4]
  assign _T_78243 = $signed(buffer_7_212) + $signed(buffer_7_213); // @[Modules.scala 166:64:@25022.4]
  assign _T_78244 = _T_78243[13:0]; // @[Modules.scala 166:64:@25023.4]
  assign buffer_7_415 = $signed(_T_78244); // @[Modules.scala 166:64:@25024.4]
  assign buffer_7_214 = {{8{_T_77266[5]}},_T_77266}; // @[Modules.scala 112:22:@8.4]
  assign _T_78246 = $signed(buffer_7_214) + $signed(buffer_5_209); // @[Modules.scala 166:64:@25026.4]
  assign _T_78247 = _T_78246[13:0]; // @[Modules.scala 166:64:@25027.4]
  assign buffer_7_416 = $signed(_T_78247); // @[Modules.scala 166:64:@25028.4]
  assign buffer_7_216 = {{8{_T_77280[5]}},_T_77280}; // @[Modules.scala 112:22:@8.4]
  assign _T_78249 = $signed(buffer_7_216) + $signed(buffer_3_218); // @[Modules.scala 166:64:@25030.4]
  assign _T_78250 = _T_78249[13:0]; // @[Modules.scala 166:64:@25031.4]
  assign buffer_7_417 = $signed(_T_78250); // @[Modules.scala 166:64:@25032.4]
  assign _T_78252 = $signed(buffer_3_219) + $signed(buffer_0_210); // @[Modules.scala 166:64:@25034.4]
  assign _T_78253 = _T_78252[13:0]; // @[Modules.scala 166:64:@25035.4]
  assign buffer_7_418 = $signed(_T_78253); // @[Modules.scala 166:64:@25036.4]
  assign _T_78255 = $signed(buffer_0_211) + $signed(buffer_0_212); // @[Modules.scala 166:64:@25038.4]
  assign _T_78256 = _T_78255[13:0]; // @[Modules.scala 166:64:@25039.4]
  assign buffer_7_419 = $signed(_T_78256); // @[Modules.scala 166:64:@25040.4]
  assign buffer_7_223 = {{8{_T_77329[5]}},_T_77329}; // @[Modules.scala 112:22:@8.4]
  assign _T_78258 = $signed(buffer_0_213) + $signed(buffer_7_223); // @[Modules.scala 166:64:@25042.4]
  assign _T_78259 = _T_78258[13:0]; // @[Modules.scala 166:64:@25043.4]
  assign buffer_7_420 = $signed(_T_78259); // @[Modules.scala 166:64:@25044.4]
  assign buffer_7_224 = {{9{_T_77336[4]}},_T_77336}; // @[Modules.scala 112:22:@8.4]
  assign _T_78261 = $signed(buffer_7_224) + $signed(buffer_1_216); // @[Modules.scala 166:64:@25046.4]
  assign _T_78262 = _T_78261[13:0]; // @[Modules.scala 166:64:@25047.4]
  assign buffer_7_421 = $signed(_T_78262); // @[Modules.scala 166:64:@25048.4]
  assign buffer_7_227 = {{8{_T_77357[5]}},_T_77357}; // @[Modules.scala 112:22:@8.4]
  assign _T_78264 = $signed(buffer_6_228) + $signed(buffer_7_227); // @[Modules.scala 166:64:@25050.4]
  assign _T_78265 = _T_78264[13:0]; // @[Modules.scala 166:64:@25051.4]
  assign buffer_7_422 = $signed(_T_78265); // @[Modules.scala 166:64:@25052.4]
  assign _T_78267 = $signed(buffer_3_229) + $signed(buffer_2_224); // @[Modules.scala 166:64:@25054.4]
  assign _T_78268 = _T_78267[13:0]; // @[Modules.scala 166:64:@25055.4]
  assign buffer_7_423 = $signed(_T_78268); // @[Modules.scala 166:64:@25056.4]
  assign buffer_7_231 = {{8{_T_77385[5]}},_T_77385}; // @[Modules.scala 112:22:@8.4]
  assign _T_78270 = $signed(buffer_5_225) + $signed(buffer_7_231); // @[Modules.scala 166:64:@25058.4]
  assign _T_78271 = _T_78270[13:0]; // @[Modules.scala 166:64:@25059.4]
  assign buffer_7_424 = $signed(_T_78271); // @[Modules.scala 166:64:@25060.4]
  assign buffer_7_232 = {{8{_T_77392[5]}},_T_77392}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_233 = {{8{_T_77399[5]}},_T_77399}; // @[Modules.scala 112:22:@8.4]
  assign _T_78273 = $signed(buffer_7_232) + $signed(buffer_7_233); // @[Modules.scala 166:64:@25062.4]
  assign _T_78274 = _T_78273[13:0]; // @[Modules.scala 166:64:@25063.4]
  assign buffer_7_425 = $signed(_T_78274); // @[Modules.scala 166:64:@25064.4]
  assign buffer_7_234 = {{8{_T_77406[5]}},_T_77406}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_235 = {{8{_T_77413[5]}},_T_77413}; // @[Modules.scala 112:22:@8.4]
  assign _T_78276 = $signed(buffer_7_234) + $signed(buffer_7_235); // @[Modules.scala 166:64:@25066.4]
  assign _T_78277 = _T_78276[13:0]; // @[Modules.scala 166:64:@25067.4]
  assign buffer_7_426 = $signed(_T_78277); // @[Modules.scala 166:64:@25068.4]
  assign buffer_7_236 = {{9{_T_77420[4]}},_T_77420}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_237 = {{8{_T_77427[5]}},_T_77427}; // @[Modules.scala 112:22:@8.4]
  assign _T_78279 = $signed(buffer_7_236) + $signed(buffer_7_237); // @[Modules.scala 166:64:@25070.4]
  assign _T_78280 = _T_78279[13:0]; // @[Modules.scala 166:64:@25071.4]
  assign buffer_7_427 = $signed(_T_78280); // @[Modules.scala 166:64:@25072.4]
  assign buffer_7_238 = {{8{_T_77434[5]}},_T_77434}; // @[Modules.scala 112:22:@8.4]
  assign _T_78282 = $signed(buffer_7_238) + $signed(buffer_1_229); // @[Modules.scala 166:64:@25074.4]
  assign _T_78283 = _T_78282[13:0]; // @[Modules.scala 166:64:@25075.4]
  assign buffer_7_428 = $signed(_T_78283); // @[Modules.scala 166:64:@25076.4]
  assign buffer_7_240 = {{9{_T_77448[4]}},_T_77448}; // @[Modules.scala 112:22:@8.4]
  assign _T_78285 = $signed(buffer_7_240) + $signed(buffer_3_240); // @[Modules.scala 166:64:@25078.4]
  assign _T_78286 = _T_78285[13:0]; // @[Modules.scala 166:64:@25079.4]
  assign buffer_7_429 = $signed(_T_78286); // @[Modules.scala 166:64:@25080.4]
  assign buffer_7_242 = {{8{_T_77462[5]}},_T_77462}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_243 = {{8{_T_77469[5]}},_T_77469}; // @[Modules.scala 112:22:@8.4]
  assign _T_78288 = $signed(buffer_7_242) + $signed(buffer_7_243); // @[Modules.scala 166:64:@25082.4]
  assign _T_78289 = _T_78288[13:0]; // @[Modules.scala 166:64:@25083.4]
  assign buffer_7_430 = $signed(_T_78289); // @[Modules.scala 166:64:@25084.4]
  assign buffer_7_245 = {{8{_T_77483[5]}},_T_77483}; // @[Modules.scala 112:22:@8.4]
  assign _T_78291 = $signed(buffer_6_244) + $signed(buffer_7_245); // @[Modules.scala 166:64:@25086.4]
  assign _T_78292 = _T_78291[13:0]; // @[Modules.scala 166:64:@25087.4]
  assign buffer_7_431 = $signed(_T_78292); // @[Modules.scala 166:64:@25088.4]
  assign buffer_7_246 = {{8{_T_77490[5]}},_T_77490}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_247 = {{8{_T_77497[5]}},_T_77497}; // @[Modules.scala 112:22:@8.4]
  assign _T_78294 = $signed(buffer_7_246) + $signed(buffer_7_247); // @[Modules.scala 166:64:@25090.4]
  assign _T_78295 = _T_78294[13:0]; // @[Modules.scala 166:64:@25091.4]
  assign buffer_7_432 = $signed(_T_78295); // @[Modules.scala 166:64:@25092.4]
  assign buffer_7_250 = {{9{_T_77518[4]}},_T_77518}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_251 = {{8{_T_77525[5]}},_T_77525}; // @[Modules.scala 112:22:@8.4]
  assign _T_78300 = $signed(buffer_7_250) + $signed(buffer_7_251); // @[Modules.scala 166:64:@25098.4]
  assign _T_78301 = _T_78300[13:0]; // @[Modules.scala 166:64:@25099.4]
  assign buffer_7_434 = $signed(_T_78301); // @[Modules.scala 166:64:@25100.4]
  assign _T_78303 = $signed(buffer_6_253) + $signed(buffer_3_252); // @[Modules.scala 166:64:@25102.4]
  assign _T_78304 = _T_78303[13:0]; // @[Modules.scala 166:64:@25103.4]
  assign buffer_7_435 = $signed(_T_78304); // @[Modules.scala 166:64:@25104.4]
  assign buffer_7_254 = {{9{_T_77546[4]}},_T_77546}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_255 = {{8{_T_77553[5]}},_T_77553}; // @[Modules.scala 112:22:@8.4]
  assign _T_78306 = $signed(buffer_7_254) + $signed(buffer_7_255); // @[Modules.scala 166:64:@25106.4]
  assign _T_78307 = _T_78306[13:0]; // @[Modules.scala 166:64:@25107.4]
  assign buffer_7_436 = $signed(_T_78307); // @[Modules.scala 166:64:@25108.4]
  assign buffer_7_256 = {{8{_T_77560[5]}},_T_77560}; // @[Modules.scala 112:22:@8.4]
  assign _T_78309 = $signed(buffer_7_256) + $signed(buffer_6_260); // @[Modules.scala 166:64:@25110.4]
  assign _T_78310 = _T_78309[13:0]; // @[Modules.scala 166:64:@25111.4]
  assign buffer_7_437 = $signed(_T_78310); // @[Modules.scala 166:64:@25112.4]
  assign _T_78312 = $signed(buffer_4_245) + $signed(buffer_4_246); // @[Modules.scala 166:64:@25114.4]
  assign _T_78313 = _T_78312[13:0]; // @[Modules.scala 166:64:@25115.4]
  assign buffer_7_438 = $signed(_T_78313); // @[Modules.scala 166:64:@25116.4]
  assign buffer_7_260 = {{8{_T_77588[5]}},_T_77588}; // @[Modules.scala 112:22:@8.4]
  assign _T_78315 = $signed(buffer_7_260) + $signed(buffer_5_261); // @[Modules.scala 166:64:@25118.4]
  assign _T_78316 = _T_78315[13:0]; // @[Modules.scala 166:64:@25119.4]
  assign buffer_7_439 = $signed(_T_78316); // @[Modules.scala 166:64:@25120.4]
  assign buffer_7_262 = {{9{_T_77602[4]}},_T_77602}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_263 = {{8{_T_77609[5]}},_T_77609}; // @[Modules.scala 112:22:@8.4]
  assign _T_78318 = $signed(buffer_7_262) + $signed(buffer_7_263); // @[Modules.scala 166:64:@25122.4]
  assign _T_78319 = _T_78318[13:0]; // @[Modules.scala 166:64:@25123.4]
  assign buffer_7_440 = $signed(_T_78319); // @[Modules.scala 166:64:@25124.4]
  assign _T_78324 = $signed(buffer_2_266) + $signed(buffer_3_268); // @[Modules.scala 166:64:@25130.4]
  assign _T_78325 = _T_78324[13:0]; // @[Modules.scala 166:64:@25131.4]
  assign buffer_7_442 = $signed(_T_78325); // @[Modules.scala 166:64:@25132.4]
  assign buffer_7_268 = {{8{_T_77644[5]}},_T_77644}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_269 = {{9{_T_77651[4]}},_T_77651}; // @[Modules.scala 112:22:@8.4]
  assign _T_78327 = $signed(buffer_7_268) + $signed(buffer_7_269); // @[Modules.scala 166:64:@25134.4]
  assign _T_78328 = _T_78327[13:0]; // @[Modules.scala 166:64:@25135.4]
  assign buffer_7_443 = $signed(_T_78328); // @[Modules.scala 166:64:@25136.4]
  assign _T_78330 = $signed(buffer_3_271) + $signed(buffer_3_272); // @[Modules.scala 166:64:@25138.4]
  assign _T_78331 = _T_78330[13:0]; // @[Modules.scala 166:64:@25139.4]
  assign buffer_7_444 = $signed(_T_78331); // @[Modules.scala 166:64:@25140.4]
  assign buffer_7_272 = {{8{_T_77672[5]}},_T_77672}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_273 = {{8{_T_77679[5]}},_T_77679}; // @[Modules.scala 112:22:@8.4]
  assign _T_78333 = $signed(buffer_7_272) + $signed(buffer_7_273); // @[Modules.scala 166:64:@25142.4]
  assign _T_78334 = _T_78333[13:0]; // @[Modules.scala 166:64:@25143.4]
  assign buffer_7_445 = $signed(_T_78334); // @[Modules.scala 166:64:@25144.4]
  assign buffer_7_278 = {{8{_T_77714[5]}},_T_77714}; // @[Modules.scala 112:22:@8.4]
  assign _T_78342 = $signed(buffer_7_278) + $signed(buffer_2_279); // @[Modules.scala 166:64:@25154.4]
  assign _T_78343 = _T_78342[13:0]; // @[Modules.scala 166:64:@25155.4]
  assign buffer_7_448 = $signed(_T_78343); // @[Modules.scala 166:64:@25156.4]
  assign buffer_7_280 = {{8{_T_77728[5]}},_T_77728}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_281 = {{9{_T_77735[4]}},_T_77735}; // @[Modules.scala 112:22:@8.4]
  assign _T_78345 = $signed(buffer_7_280) + $signed(buffer_7_281); // @[Modules.scala 166:64:@25158.4]
  assign _T_78346 = _T_78345[13:0]; // @[Modules.scala 166:64:@25159.4]
  assign buffer_7_449 = $signed(_T_78346); // @[Modules.scala 166:64:@25160.4]
  assign buffer_7_282 = {{8{_T_77742[5]}},_T_77742}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_283 = {{8{_T_77749[5]}},_T_77749}; // @[Modules.scala 112:22:@8.4]
  assign _T_78348 = $signed(buffer_7_282) + $signed(buffer_7_283); // @[Modules.scala 166:64:@25162.4]
  assign _T_78349 = _T_78348[13:0]; // @[Modules.scala 166:64:@25163.4]
  assign buffer_7_450 = $signed(_T_78349); // @[Modules.scala 166:64:@25164.4]
  assign _T_78351 = $signed(buffer_0_278) + $signed(buffer_0_280); // @[Modules.scala 166:64:@25166.4]
  assign _T_78352 = _T_78351[13:0]; // @[Modules.scala 166:64:@25167.4]
  assign buffer_7_451 = $signed(_T_78352); // @[Modules.scala 166:64:@25168.4]
  assign _T_78354 = $signed(buffer_0_281) + $signed(buffer_0_282); // @[Modules.scala 166:64:@25170.4]
  assign _T_78355 = _T_78354[13:0]; // @[Modules.scala 166:64:@25171.4]
  assign buffer_7_452 = $signed(_T_78355); // @[Modules.scala 166:64:@25172.4]
  assign buffer_7_289 = {{8{_T_77791[5]}},_T_77791}; // @[Modules.scala 112:22:@8.4]
  assign _T_78357 = $signed(buffer_0_283) + $signed(buffer_7_289); // @[Modules.scala 166:64:@25174.4]
  assign _T_78358 = _T_78357[13:0]; // @[Modules.scala 166:64:@25175.4]
  assign buffer_7_453 = $signed(_T_78358); // @[Modules.scala 166:64:@25176.4]
  assign buffer_7_291 = {{9{_T_77805[4]}},_T_77805}; // @[Modules.scala 112:22:@8.4]
  assign _T_78360 = $signed(buffer_1_283) + $signed(buffer_7_291); // @[Modules.scala 166:64:@25178.4]
  assign _T_78361 = _T_78360[13:0]; // @[Modules.scala 166:64:@25179.4]
  assign buffer_7_454 = $signed(_T_78361); // @[Modules.scala 166:64:@25180.4]
  assign buffer_7_293 = {{8{_T_77819[5]}},_T_77819}; // @[Modules.scala 112:22:@8.4]
  assign _T_78363 = $signed(buffer_3_295) + $signed(buffer_7_293); // @[Modules.scala 166:64:@25182.4]
  assign _T_78364 = _T_78363[13:0]; // @[Modules.scala 166:64:@25183.4]
  assign buffer_7_455 = $signed(_T_78364); // @[Modules.scala 166:64:@25184.4]
  assign _T_78366 = $signed(buffer_0_287) + $signed(buffer_1_288); // @[Modules.scala 166:64:@25186.4]
  assign _T_78367 = _T_78366[13:0]; // @[Modules.scala 166:64:@25187.4]
  assign buffer_7_456 = $signed(_T_78367); // @[Modules.scala 166:64:@25188.4]
  assign buffer_7_296 = {{8{_T_77840[5]}},_T_77840}; // @[Modules.scala 112:22:@8.4]
  assign _T_78369 = $signed(buffer_7_296) + $signed(buffer_0_290); // @[Modules.scala 166:64:@25190.4]
  assign _T_78370 = _T_78369[13:0]; // @[Modules.scala 166:64:@25191.4]
  assign buffer_7_457 = $signed(_T_78370); // @[Modules.scala 166:64:@25192.4]
  assign buffer_7_298 = {{8{_T_77854[5]}},_T_77854}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_299 = {{8{_T_77861[5]}},_T_77861}; // @[Modules.scala 112:22:@8.4]
  assign _T_78372 = $signed(buffer_7_298) + $signed(buffer_7_299); // @[Modules.scala 166:64:@25194.4]
  assign _T_78373 = _T_78372[13:0]; // @[Modules.scala 166:64:@25195.4]
  assign buffer_7_458 = $signed(_T_78373); // @[Modules.scala 166:64:@25196.4]
  assign buffer_7_300 = {{8{_T_77868[5]}},_T_77868}; // @[Modules.scala 112:22:@8.4]
  assign buffer_7_301 = {{8{_T_77875[5]}},_T_77875}; // @[Modules.scala 112:22:@8.4]
  assign _T_78375 = $signed(buffer_7_300) + $signed(buffer_7_301); // @[Modules.scala 166:64:@25198.4]
  assign _T_78376 = _T_78375[13:0]; // @[Modules.scala 166:64:@25199.4]
  assign buffer_7_459 = $signed(_T_78376); // @[Modules.scala 166:64:@25200.4]
  assign buffer_7_303 = {{8{_T_77889[5]}},_T_77889}; // @[Modules.scala 112:22:@8.4]
  assign _T_78378 = $signed(buffer_0_295) + $signed(buffer_7_303); // @[Modules.scala 166:64:@25202.4]
  assign _T_78379 = _T_78378[13:0]; // @[Modules.scala 166:64:@25203.4]
  assign buffer_7_460 = $signed(_T_78379); // @[Modules.scala 166:64:@25204.4]
  assign buffer_7_307 = {{8{_T_77917[5]}},_T_77917}; // @[Modules.scala 112:22:@8.4]
  assign _T_78384 = $signed(buffer_1_300) + $signed(buffer_7_307); // @[Modules.scala 166:64:@25210.4]
  assign _T_78385 = _T_78384[13:0]; // @[Modules.scala 166:64:@25211.4]
  assign buffer_7_462 = $signed(_T_78385); // @[Modules.scala 166:64:@25212.4]
  assign _T_78387 = $signed(buffer_7_309) + $signed(buffer_7_310); // @[Modules.scala 160:64:@25214.4]
  assign _T_78388 = _T_78387[13:0]; // @[Modules.scala 160:64:@25215.4]
  assign buffer_7_463 = $signed(_T_78388); // @[Modules.scala 160:64:@25216.4]
  assign _T_78390 = $signed(buffer_7_311) + $signed(buffer_7_312); // @[Modules.scala 160:64:@25218.4]
  assign _T_78391 = _T_78390[13:0]; // @[Modules.scala 160:64:@25219.4]
  assign buffer_7_464 = $signed(_T_78391); // @[Modules.scala 160:64:@25220.4]
  assign _T_78393 = $signed(buffer_7_313) + $signed(buffer_0_307); // @[Modules.scala 160:64:@25222.4]
  assign _T_78394 = _T_78393[13:0]; // @[Modules.scala 160:64:@25223.4]
  assign buffer_7_465 = $signed(_T_78394); // @[Modules.scala 160:64:@25224.4]
  assign _T_78396 = $signed(buffer_7_315) + $signed(buffer_7_316); // @[Modules.scala 160:64:@25226.4]
  assign _T_78397 = _T_78396[13:0]; // @[Modules.scala 160:64:@25227.4]
  assign buffer_7_466 = $signed(_T_78397); // @[Modules.scala 160:64:@25228.4]
  assign _T_78399 = $signed(buffer_7_317) + $signed(buffer_7_318); // @[Modules.scala 160:64:@25230.4]
  assign _T_78400 = _T_78399[13:0]; // @[Modules.scala 160:64:@25231.4]
  assign buffer_7_467 = $signed(_T_78400); // @[Modules.scala 160:64:@25232.4]
  assign _T_78402 = $signed(buffer_7_319) + $signed(buffer_7_320); // @[Modules.scala 160:64:@25234.4]
  assign _T_78403 = _T_78402[13:0]; // @[Modules.scala 160:64:@25235.4]
  assign buffer_7_468 = $signed(_T_78403); // @[Modules.scala 160:64:@25236.4]
  assign _T_78405 = $signed(buffer_7_321) + $signed(buffer_1_317); // @[Modules.scala 160:64:@25238.4]
  assign _T_78406 = _T_78405[13:0]; // @[Modules.scala 160:64:@25239.4]
  assign buffer_7_469 = $signed(_T_78406); // @[Modules.scala 160:64:@25240.4]
  assign _T_78408 = $signed(buffer_7_323) + $signed(buffer_7_324); // @[Modules.scala 160:64:@25242.4]
  assign _T_78409 = _T_78408[13:0]; // @[Modules.scala 160:64:@25243.4]
  assign buffer_7_470 = $signed(_T_78409); // @[Modules.scala 160:64:@25244.4]
  assign _T_78411 = $signed(buffer_7_325) + $signed(buffer_7_326); // @[Modules.scala 160:64:@25246.4]
  assign _T_78412 = _T_78411[13:0]; // @[Modules.scala 160:64:@25247.4]
  assign buffer_7_471 = $signed(_T_78412); // @[Modules.scala 160:64:@25248.4]
  assign _T_78414 = $signed(buffer_7_327) + $signed(buffer_7_328); // @[Modules.scala 160:64:@25250.4]
  assign _T_78415 = _T_78414[13:0]; // @[Modules.scala 160:64:@25251.4]
  assign buffer_7_472 = $signed(_T_78415); // @[Modules.scala 160:64:@25252.4]
  assign _T_78417 = $signed(buffer_7_329) + $signed(buffer_7_330); // @[Modules.scala 160:64:@25254.4]
  assign _T_78418 = _T_78417[13:0]; // @[Modules.scala 160:64:@25255.4]
  assign buffer_7_473 = $signed(_T_78418); // @[Modules.scala 160:64:@25256.4]
  assign _T_78420 = $signed(buffer_7_331) + $signed(buffer_3_337); // @[Modules.scala 160:64:@25258.4]
  assign _T_78421 = _T_78420[13:0]; // @[Modules.scala 160:64:@25259.4]
  assign buffer_7_474 = $signed(_T_78421); // @[Modules.scala 160:64:@25260.4]
  assign _T_78423 = $signed(buffer_7_333) + $signed(buffer_7_334); // @[Modules.scala 160:64:@25262.4]
  assign _T_78424 = _T_78423[13:0]; // @[Modules.scala 160:64:@25263.4]
  assign buffer_7_475 = $signed(_T_78424); // @[Modules.scala 160:64:@25264.4]
  assign _T_78426 = $signed(buffer_7_335) + $signed(buffer_7_336); // @[Modules.scala 160:64:@25266.4]
  assign _T_78427 = _T_78426[13:0]; // @[Modules.scala 160:64:@25267.4]
  assign buffer_7_476 = $signed(_T_78427); // @[Modules.scala 160:64:@25268.4]
  assign _T_78429 = $signed(buffer_7_337) + $signed(buffer_7_338); // @[Modules.scala 160:64:@25270.4]
  assign _T_78430 = _T_78429[13:0]; // @[Modules.scala 160:64:@25271.4]
  assign buffer_7_477 = $signed(_T_78430); // @[Modules.scala 160:64:@25272.4]
  assign _T_78432 = $signed(buffer_7_339) + $signed(buffer_7_340); // @[Modules.scala 160:64:@25274.4]
  assign _T_78433 = _T_78432[13:0]; // @[Modules.scala 160:64:@25275.4]
  assign buffer_7_478 = $signed(_T_78433); // @[Modules.scala 160:64:@25276.4]
  assign _T_78435 = $signed(buffer_7_341) + $signed(buffer_7_342); // @[Modules.scala 160:64:@25278.4]
  assign _T_78436 = _T_78435[13:0]; // @[Modules.scala 160:64:@25279.4]
  assign buffer_7_479 = $signed(_T_78436); // @[Modules.scala 160:64:@25280.4]
  assign _T_78438 = $signed(buffer_7_343) + $signed(buffer_7_344); // @[Modules.scala 160:64:@25282.4]
  assign _T_78439 = _T_78438[13:0]; // @[Modules.scala 160:64:@25283.4]
  assign buffer_7_480 = $signed(_T_78439); // @[Modules.scala 160:64:@25284.4]
  assign _T_78441 = $signed(buffer_7_345) + $signed(buffer_7_346); // @[Modules.scala 160:64:@25286.4]
  assign _T_78442 = _T_78441[13:0]; // @[Modules.scala 160:64:@25287.4]
  assign buffer_7_481 = $signed(_T_78442); // @[Modules.scala 160:64:@25288.4]
  assign _T_78444 = $signed(buffer_7_347) + $signed(buffer_6_355); // @[Modules.scala 160:64:@25290.4]
  assign _T_78445 = _T_78444[13:0]; // @[Modules.scala 160:64:@25291.4]
  assign buffer_7_482 = $signed(_T_78445); // @[Modules.scala 160:64:@25292.4]
  assign _T_78447 = $signed(buffer_6_356) + $signed(buffer_7_350); // @[Modules.scala 160:64:@25294.4]
  assign _T_78448 = _T_78447[13:0]; // @[Modules.scala 160:64:@25295.4]
  assign buffer_7_483 = $signed(_T_78448); // @[Modules.scala 160:64:@25296.4]
  assign _T_78450 = $signed(buffer_7_351) + $signed(buffer_7_352); // @[Modules.scala 160:64:@25298.4]
  assign _T_78451 = _T_78450[13:0]; // @[Modules.scala 160:64:@25299.4]
  assign buffer_7_484 = $signed(_T_78451); // @[Modules.scala 160:64:@25300.4]
  assign _T_78453 = $signed(buffer_7_353) + $signed(buffer_7_354); // @[Modules.scala 160:64:@25302.4]
  assign _T_78454 = _T_78453[13:0]; // @[Modules.scala 160:64:@25303.4]
  assign buffer_7_485 = $signed(_T_78454); // @[Modules.scala 160:64:@25304.4]
  assign _T_78456 = $signed(buffer_7_355) + $signed(buffer_7_356); // @[Modules.scala 160:64:@25306.4]
  assign _T_78457 = _T_78456[13:0]; // @[Modules.scala 160:64:@25307.4]
  assign buffer_7_486 = $signed(_T_78457); // @[Modules.scala 160:64:@25308.4]
  assign _T_78459 = $signed(buffer_7_357) + $signed(buffer_6_365); // @[Modules.scala 160:64:@25310.4]
  assign _T_78460 = _T_78459[13:0]; // @[Modules.scala 160:64:@25311.4]
  assign buffer_7_487 = $signed(_T_78460); // @[Modules.scala 160:64:@25312.4]
  assign _T_78462 = $signed(buffer_7_359) + $signed(buffer_7_360); // @[Modules.scala 160:64:@25314.4]
  assign _T_78463 = _T_78462[13:0]; // @[Modules.scala 160:64:@25315.4]
  assign buffer_7_488 = $signed(_T_78463); // @[Modules.scala 160:64:@25316.4]
  assign _T_78465 = $signed(buffer_7_361) + $signed(buffer_7_362); // @[Modules.scala 160:64:@25318.4]
  assign _T_78466 = _T_78465[13:0]; // @[Modules.scala 160:64:@25319.4]
  assign buffer_7_489 = $signed(_T_78466); // @[Modules.scala 160:64:@25320.4]
  assign _T_78468 = $signed(buffer_3_369) + $signed(buffer_4_353); // @[Modules.scala 160:64:@25322.4]
  assign _T_78469 = _T_78468[13:0]; // @[Modules.scala 160:64:@25323.4]
  assign buffer_7_490 = $signed(_T_78469); // @[Modules.scala 160:64:@25324.4]
  assign _T_78471 = $signed(buffer_7_365) + $signed(buffer_7_366); // @[Modules.scala 160:64:@25326.4]
  assign _T_78472 = _T_78471[13:0]; // @[Modules.scala 160:64:@25327.4]
  assign buffer_7_491 = $signed(_T_78472); // @[Modules.scala 160:64:@25328.4]
  assign _T_78474 = $signed(buffer_7_367) + $signed(buffer_7_368); // @[Modules.scala 160:64:@25330.4]
  assign _T_78475 = _T_78474[13:0]; // @[Modules.scala 160:64:@25331.4]
  assign buffer_7_492 = $signed(_T_78475); // @[Modules.scala 160:64:@25332.4]
  assign _T_78477 = $signed(buffer_7_369) + $signed(buffer_7_370); // @[Modules.scala 160:64:@25334.4]
  assign _T_78478 = _T_78477[13:0]; // @[Modules.scala 160:64:@25335.4]
  assign buffer_7_493 = $signed(_T_78478); // @[Modules.scala 160:64:@25336.4]
  assign _T_78480 = $signed(buffer_7_371) + $signed(buffer_7_372); // @[Modules.scala 160:64:@25338.4]
  assign _T_78481 = _T_78480[13:0]; // @[Modules.scala 160:64:@25339.4]
  assign buffer_7_494 = $signed(_T_78481); // @[Modules.scala 160:64:@25340.4]
  assign _T_78483 = $signed(buffer_7_373) + $signed(buffer_0_367); // @[Modules.scala 160:64:@25342.4]
  assign _T_78484 = _T_78483[13:0]; // @[Modules.scala 160:64:@25343.4]
  assign buffer_7_495 = $signed(_T_78484); // @[Modules.scala 160:64:@25344.4]
  assign _T_78486 = $signed(buffer_7_375) + $signed(buffer_7_376); // @[Modules.scala 160:64:@25346.4]
  assign _T_78487 = _T_78486[13:0]; // @[Modules.scala 160:64:@25347.4]
  assign buffer_7_496 = $signed(_T_78487); // @[Modules.scala 160:64:@25348.4]
  assign _T_78489 = $signed(buffer_7_377) + $signed(buffer_7_378); // @[Modules.scala 160:64:@25350.4]
  assign _T_78490 = _T_78489[13:0]; // @[Modules.scala 160:64:@25351.4]
  assign buffer_7_497 = $signed(_T_78490); // @[Modules.scala 160:64:@25352.4]
  assign _T_78492 = $signed(buffer_7_379) + $signed(buffer_7_380); // @[Modules.scala 160:64:@25354.4]
  assign _T_78493 = _T_78492[13:0]; // @[Modules.scala 160:64:@25355.4]
  assign buffer_7_498 = $signed(_T_78493); // @[Modules.scala 160:64:@25356.4]
  assign _T_78495 = $signed(buffer_7_381) + $signed(buffer_7_382); // @[Modules.scala 160:64:@25358.4]
  assign _T_78496 = _T_78495[13:0]; // @[Modules.scala 160:64:@25359.4]
  assign buffer_7_499 = $signed(_T_78496); // @[Modules.scala 160:64:@25360.4]
  assign _T_78498 = $signed(buffer_7_383) + $signed(buffer_7_384); // @[Modules.scala 160:64:@25362.4]
  assign _T_78499 = _T_78498[13:0]; // @[Modules.scala 160:64:@25363.4]
  assign buffer_7_500 = $signed(_T_78499); // @[Modules.scala 160:64:@25364.4]
  assign _T_78501 = $signed(buffer_7_385) + $signed(buffer_5_391); // @[Modules.scala 160:64:@25366.4]
  assign _T_78502 = _T_78501[13:0]; // @[Modules.scala 160:64:@25367.4]
  assign buffer_7_501 = $signed(_T_78502); // @[Modules.scala 160:64:@25368.4]
  assign _T_78504 = $signed(buffer_7_387) + $signed(buffer_7_388); // @[Modules.scala 160:64:@25370.4]
  assign _T_78505 = _T_78504[13:0]; // @[Modules.scala 160:64:@25371.4]
  assign buffer_7_502 = $signed(_T_78505); // @[Modules.scala 160:64:@25372.4]
  assign _T_78507 = $signed(buffer_7_389) + $signed(buffer_7_390); // @[Modules.scala 160:64:@25374.4]
  assign _T_78508 = _T_78507[13:0]; // @[Modules.scala 160:64:@25375.4]
  assign buffer_7_503 = $signed(_T_78508); // @[Modules.scala 160:64:@25376.4]
  assign _T_78510 = $signed(buffer_7_391) + $signed(buffer_7_392); // @[Modules.scala 160:64:@25378.4]
  assign _T_78511 = _T_78510[13:0]; // @[Modules.scala 160:64:@25379.4]
  assign buffer_7_504 = $signed(_T_78511); // @[Modules.scala 160:64:@25380.4]
  assign _T_78513 = $signed(buffer_7_393) + $signed(buffer_7_394); // @[Modules.scala 160:64:@25382.4]
  assign _T_78514 = _T_78513[13:0]; // @[Modules.scala 160:64:@25383.4]
  assign buffer_7_505 = $signed(_T_78514); // @[Modules.scala 160:64:@25384.4]
  assign _T_78516 = $signed(buffer_7_395) + $signed(buffer_7_396); // @[Modules.scala 160:64:@25386.4]
  assign _T_78517 = _T_78516[13:0]; // @[Modules.scala 160:64:@25387.4]
  assign buffer_7_506 = $signed(_T_78517); // @[Modules.scala 160:64:@25388.4]
  assign _T_78519 = $signed(buffer_7_397) + $signed(buffer_7_398); // @[Modules.scala 160:64:@25390.4]
  assign _T_78520 = _T_78519[13:0]; // @[Modules.scala 160:64:@25391.4]
  assign buffer_7_507 = $signed(_T_78520); // @[Modules.scala 160:64:@25392.4]
  assign _T_78522 = $signed(buffer_1_392) + $signed(buffer_7_400); // @[Modules.scala 160:64:@25394.4]
  assign _T_78523 = _T_78522[13:0]; // @[Modules.scala 160:64:@25395.4]
  assign buffer_7_508 = $signed(_T_78523); // @[Modules.scala 160:64:@25396.4]
  assign _T_78525 = $signed(buffer_7_401) + $signed(buffer_7_402); // @[Modules.scala 160:64:@25398.4]
  assign _T_78526 = _T_78525[13:0]; // @[Modules.scala 160:64:@25399.4]
  assign buffer_7_509 = $signed(_T_78526); // @[Modules.scala 160:64:@25400.4]
  assign _T_78528 = $signed(buffer_7_403) + $signed(buffer_7_404); // @[Modules.scala 160:64:@25402.4]
  assign _T_78529 = _T_78528[13:0]; // @[Modules.scala 160:64:@25403.4]
  assign buffer_7_510 = $signed(_T_78529); // @[Modules.scala 160:64:@25404.4]
  assign _T_78531 = $signed(buffer_7_405) + $signed(buffer_7_406); // @[Modules.scala 160:64:@25406.4]
  assign _T_78532 = _T_78531[13:0]; // @[Modules.scala 160:64:@25407.4]
  assign buffer_7_511 = $signed(_T_78532); // @[Modules.scala 160:64:@25408.4]
  assign _T_78534 = $signed(buffer_0_396) + $signed(buffer_7_408); // @[Modules.scala 160:64:@25410.4]
  assign _T_78535 = _T_78534[13:0]; // @[Modules.scala 160:64:@25411.4]
  assign buffer_7_512 = $signed(_T_78535); // @[Modules.scala 160:64:@25412.4]
  assign _T_78537 = $signed(buffer_7_409) + $signed(buffer_7_410); // @[Modules.scala 160:64:@25414.4]
  assign _T_78538 = _T_78537[13:0]; // @[Modules.scala 160:64:@25415.4]
  assign buffer_7_513 = $signed(_T_78538); // @[Modules.scala 160:64:@25416.4]
  assign _T_78540 = $signed(buffer_7_411) + $signed(buffer_7_412); // @[Modules.scala 160:64:@25418.4]
  assign _T_78541 = _T_78540[13:0]; // @[Modules.scala 160:64:@25419.4]
  assign buffer_7_514 = $signed(_T_78541); // @[Modules.scala 160:64:@25420.4]
  assign _T_78543 = $signed(buffer_7_413) + $signed(buffer_7_414); // @[Modules.scala 160:64:@25422.4]
  assign _T_78544 = _T_78543[13:0]; // @[Modules.scala 160:64:@25423.4]
  assign buffer_7_515 = $signed(_T_78544); // @[Modules.scala 160:64:@25424.4]
  assign _T_78546 = $signed(buffer_7_415) + $signed(buffer_7_416); // @[Modules.scala 160:64:@25426.4]
  assign _T_78547 = _T_78546[13:0]; // @[Modules.scala 160:64:@25427.4]
  assign buffer_7_516 = $signed(_T_78547); // @[Modules.scala 160:64:@25428.4]
  assign _T_78549 = $signed(buffer_7_417) + $signed(buffer_7_418); // @[Modules.scala 160:64:@25430.4]
  assign _T_78550 = _T_78549[13:0]; // @[Modules.scala 160:64:@25431.4]
  assign buffer_7_517 = $signed(_T_78550); // @[Modules.scala 160:64:@25432.4]
  assign _T_78552 = $signed(buffer_7_419) + $signed(buffer_7_420); // @[Modules.scala 160:64:@25434.4]
  assign _T_78553 = _T_78552[13:0]; // @[Modules.scala 160:64:@25435.4]
  assign buffer_7_518 = $signed(_T_78553); // @[Modules.scala 160:64:@25436.4]
  assign _T_78555 = $signed(buffer_7_421) + $signed(buffer_7_422); // @[Modules.scala 160:64:@25438.4]
  assign _T_78556 = _T_78555[13:0]; // @[Modules.scala 160:64:@25439.4]
  assign buffer_7_519 = $signed(_T_78556); // @[Modules.scala 160:64:@25440.4]
  assign _T_78558 = $signed(buffer_7_423) + $signed(buffer_7_424); // @[Modules.scala 160:64:@25442.4]
  assign _T_78559 = _T_78558[13:0]; // @[Modules.scala 160:64:@25443.4]
  assign buffer_7_520 = $signed(_T_78559); // @[Modules.scala 160:64:@25444.4]
  assign _T_78561 = $signed(buffer_7_425) + $signed(buffer_7_426); // @[Modules.scala 160:64:@25446.4]
  assign _T_78562 = _T_78561[13:0]; // @[Modules.scala 160:64:@25447.4]
  assign buffer_7_521 = $signed(_T_78562); // @[Modules.scala 160:64:@25448.4]
  assign _T_78564 = $signed(buffer_7_427) + $signed(buffer_7_428); // @[Modules.scala 160:64:@25450.4]
  assign _T_78565 = _T_78564[13:0]; // @[Modules.scala 160:64:@25451.4]
  assign buffer_7_522 = $signed(_T_78565); // @[Modules.scala 160:64:@25452.4]
  assign _T_78567 = $signed(buffer_7_429) + $signed(buffer_7_430); // @[Modules.scala 160:64:@25454.4]
  assign _T_78568 = _T_78567[13:0]; // @[Modules.scala 160:64:@25455.4]
  assign buffer_7_523 = $signed(_T_78568); // @[Modules.scala 160:64:@25456.4]
  assign _T_78570 = $signed(buffer_7_431) + $signed(buffer_7_432); // @[Modules.scala 160:64:@25458.4]
  assign _T_78571 = _T_78570[13:0]; // @[Modules.scala 160:64:@25459.4]
  assign buffer_7_524 = $signed(_T_78571); // @[Modules.scala 160:64:@25460.4]
  assign _T_78573 = $signed(buffer_4_416) + $signed(buffer_7_434); // @[Modules.scala 160:64:@25462.4]
  assign _T_78574 = _T_78573[13:0]; // @[Modules.scala 160:64:@25463.4]
  assign buffer_7_525 = $signed(_T_78574); // @[Modules.scala 160:64:@25464.4]
  assign _T_78576 = $signed(buffer_7_435) + $signed(buffer_7_436); // @[Modules.scala 160:64:@25466.4]
  assign _T_78577 = _T_78576[13:0]; // @[Modules.scala 160:64:@25467.4]
  assign buffer_7_526 = $signed(_T_78577); // @[Modules.scala 160:64:@25468.4]
  assign _T_78579 = $signed(buffer_7_437) + $signed(buffer_7_438); // @[Modules.scala 160:64:@25470.4]
  assign _T_78580 = _T_78579[13:0]; // @[Modules.scala 160:64:@25471.4]
  assign buffer_7_527 = $signed(_T_78580); // @[Modules.scala 160:64:@25472.4]
  assign _T_78582 = $signed(buffer_7_439) + $signed(buffer_7_440); // @[Modules.scala 160:64:@25474.4]
  assign _T_78583 = _T_78582[13:0]; // @[Modules.scala 160:64:@25475.4]
  assign buffer_7_528 = $signed(_T_78583); // @[Modules.scala 160:64:@25476.4]
  assign _T_78585 = $signed(buffer_5_446) + $signed(buffer_7_442); // @[Modules.scala 160:64:@25478.4]
  assign _T_78586 = _T_78585[13:0]; // @[Modules.scala 160:64:@25479.4]
  assign buffer_7_529 = $signed(_T_78586); // @[Modules.scala 160:64:@25480.4]
  assign _T_78588 = $signed(buffer_7_443) + $signed(buffer_7_444); // @[Modules.scala 160:64:@25482.4]
  assign _T_78589 = _T_78588[13:0]; // @[Modules.scala 160:64:@25483.4]
  assign buffer_7_530 = $signed(_T_78589); // @[Modules.scala 160:64:@25484.4]
  assign _T_78591 = $signed(buffer_7_445) + $signed(buffer_6_455); // @[Modules.scala 160:64:@25486.4]
  assign _T_78592 = _T_78591[13:0]; // @[Modules.scala 160:64:@25487.4]
  assign buffer_7_531 = $signed(_T_78592); // @[Modules.scala 160:64:@25488.4]
  assign _T_78594 = $signed(buffer_6_456) + $signed(buffer_7_448); // @[Modules.scala 160:64:@25490.4]
  assign _T_78595 = _T_78594[13:0]; // @[Modules.scala 160:64:@25491.4]
  assign buffer_7_532 = $signed(_T_78595); // @[Modules.scala 160:64:@25492.4]
  assign _T_78597 = $signed(buffer_7_449) + $signed(buffer_7_450); // @[Modules.scala 160:64:@25494.4]
  assign _T_78598 = _T_78597[13:0]; // @[Modules.scala 160:64:@25495.4]
  assign buffer_7_533 = $signed(_T_78598); // @[Modules.scala 160:64:@25496.4]
  assign _T_78600 = $signed(buffer_7_451) + $signed(buffer_7_452); // @[Modules.scala 160:64:@25498.4]
  assign _T_78601 = _T_78600[13:0]; // @[Modules.scala 160:64:@25499.4]
  assign buffer_7_534 = $signed(_T_78601); // @[Modules.scala 160:64:@25500.4]
  assign _T_78603 = $signed(buffer_7_453) + $signed(buffer_7_454); // @[Modules.scala 160:64:@25502.4]
  assign _T_78604 = _T_78603[13:0]; // @[Modules.scala 160:64:@25503.4]
  assign buffer_7_535 = $signed(_T_78604); // @[Modules.scala 160:64:@25504.4]
  assign _T_78606 = $signed(buffer_7_455) + $signed(buffer_7_456); // @[Modules.scala 160:64:@25506.4]
  assign _T_78607 = _T_78606[13:0]; // @[Modules.scala 160:64:@25507.4]
  assign buffer_7_536 = $signed(_T_78607); // @[Modules.scala 160:64:@25508.4]
  assign _T_78609 = $signed(buffer_7_457) + $signed(buffer_7_458); // @[Modules.scala 160:64:@25510.4]
  assign _T_78610 = _T_78609[13:0]; // @[Modules.scala 160:64:@25511.4]
  assign buffer_7_537 = $signed(_T_78610); // @[Modules.scala 160:64:@25512.4]
  assign _T_78612 = $signed(buffer_7_459) + $signed(buffer_7_460); // @[Modules.scala 160:64:@25514.4]
  assign _T_78613 = _T_78612[13:0]; // @[Modules.scala 160:64:@25515.4]
  assign buffer_7_538 = $signed(_T_78613); // @[Modules.scala 160:64:@25516.4]
  assign _T_78615 = $signed(buffer_1_453) + $signed(buffer_7_462); // @[Modules.scala 160:64:@25518.4]
  assign _T_78616 = _T_78615[13:0]; // @[Modules.scala 160:64:@25519.4]
  assign buffer_7_539 = $signed(_T_78616); // @[Modules.scala 160:64:@25520.4]
  assign _T_78618 = $signed(buffer_7_463) + $signed(buffer_7_464); // @[Modules.scala 166:64:@25522.4]
  assign _T_78619 = _T_78618[13:0]; // @[Modules.scala 166:64:@25523.4]
  assign buffer_7_540 = $signed(_T_78619); // @[Modules.scala 166:64:@25524.4]
  assign _T_78621 = $signed(buffer_7_465) + $signed(buffer_7_466); // @[Modules.scala 166:64:@25526.4]
  assign _T_78622 = _T_78621[13:0]; // @[Modules.scala 166:64:@25527.4]
  assign buffer_7_541 = $signed(_T_78622); // @[Modules.scala 166:64:@25528.4]
  assign _T_78624 = $signed(buffer_7_467) + $signed(buffer_7_468); // @[Modules.scala 166:64:@25530.4]
  assign _T_78625 = _T_78624[13:0]; // @[Modules.scala 166:64:@25531.4]
  assign buffer_7_542 = $signed(_T_78625); // @[Modules.scala 166:64:@25532.4]
  assign _T_78627 = $signed(buffer_7_469) + $signed(buffer_7_470); // @[Modules.scala 166:64:@25534.4]
  assign _T_78628 = _T_78627[13:0]; // @[Modules.scala 166:64:@25535.4]
  assign buffer_7_543 = $signed(_T_78628); // @[Modules.scala 166:64:@25536.4]
  assign _T_78630 = $signed(buffer_7_471) + $signed(buffer_7_472); // @[Modules.scala 166:64:@25538.4]
  assign _T_78631 = _T_78630[13:0]; // @[Modules.scala 166:64:@25539.4]
  assign buffer_7_544 = $signed(_T_78631); // @[Modules.scala 166:64:@25540.4]
  assign _T_78633 = $signed(buffer_7_473) + $signed(buffer_7_474); // @[Modules.scala 166:64:@25542.4]
  assign _T_78634 = _T_78633[13:0]; // @[Modules.scala 166:64:@25543.4]
  assign buffer_7_545 = $signed(_T_78634); // @[Modules.scala 166:64:@25544.4]
  assign _T_78636 = $signed(buffer_7_475) + $signed(buffer_7_476); // @[Modules.scala 166:64:@25546.4]
  assign _T_78637 = _T_78636[13:0]; // @[Modules.scala 166:64:@25547.4]
  assign buffer_7_546 = $signed(_T_78637); // @[Modules.scala 166:64:@25548.4]
  assign _T_78639 = $signed(buffer_7_477) + $signed(buffer_7_478); // @[Modules.scala 166:64:@25550.4]
  assign _T_78640 = _T_78639[13:0]; // @[Modules.scala 166:64:@25551.4]
  assign buffer_7_547 = $signed(_T_78640); // @[Modules.scala 166:64:@25552.4]
  assign _T_78642 = $signed(buffer_7_479) + $signed(buffer_7_480); // @[Modules.scala 166:64:@25554.4]
  assign _T_78643 = _T_78642[13:0]; // @[Modules.scala 166:64:@25555.4]
  assign buffer_7_548 = $signed(_T_78643); // @[Modules.scala 166:64:@25556.4]
  assign _T_78645 = $signed(buffer_7_481) + $signed(buffer_7_482); // @[Modules.scala 166:64:@25558.4]
  assign _T_78646 = _T_78645[13:0]; // @[Modules.scala 166:64:@25559.4]
  assign buffer_7_549 = $signed(_T_78646); // @[Modules.scala 166:64:@25560.4]
  assign _T_78648 = $signed(buffer_7_483) + $signed(buffer_7_484); // @[Modules.scala 166:64:@25562.4]
  assign _T_78649 = _T_78648[13:0]; // @[Modules.scala 166:64:@25563.4]
  assign buffer_7_550 = $signed(_T_78649); // @[Modules.scala 166:64:@25564.4]
  assign _T_78651 = $signed(buffer_7_485) + $signed(buffer_7_486); // @[Modules.scala 166:64:@25566.4]
  assign _T_78652 = _T_78651[13:0]; // @[Modules.scala 166:64:@25567.4]
  assign buffer_7_551 = $signed(_T_78652); // @[Modules.scala 166:64:@25568.4]
  assign _T_78654 = $signed(buffer_7_487) + $signed(buffer_7_488); // @[Modules.scala 166:64:@25570.4]
  assign _T_78655 = _T_78654[13:0]; // @[Modules.scala 166:64:@25571.4]
  assign buffer_7_552 = $signed(_T_78655); // @[Modules.scala 166:64:@25572.4]
  assign _T_78657 = $signed(buffer_7_489) + $signed(buffer_7_490); // @[Modules.scala 166:64:@25574.4]
  assign _T_78658 = _T_78657[13:0]; // @[Modules.scala 166:64:@25575.4]
  assign buffer_7_553 = $signed(_T_78658); // @[Modules.scala 166:64:@25576.4]
  assign _T_78660 = $signed(buffer_7_491) + $signed(buffer_7_492); // @[Modules.scala 166:64:@25578.4]
  assign _T_78661 = _T_78660[13:0]; // @[Modules.scala 166:64:@25579.4]
  assign buffer_7_554 = $signed(_T_78661); // @[Modules.scala 166:64:@25580.4]
  assign _T_78663 = $signed(buffer_7_493) + $signed(buffer_7_494); // @[Modules.scala 166:64:@25582.4]
  assign _T_78664 = _T_78663[13:0]; // @[Modules.scala 166:64:@25583.4]
  assign buffer_7_555 = $signed(_T_78664); // @[Modules.scala 166:64:@25584.4]
  assign _T_78666 = $signed(buffer_7_495) + $signed(buffer_7_496); // @[Modules.scala 166:64:@25586.4]
  assign _T_78667 = _T_78666[13:0]; // @[Modules.scala 166:64:@25587.4]
  assign buffer_7_556 = $signed(_T_78667); // @[Modules.scala 166:64:@25588.4]
  assign _T_78669 = $signed(buffer_7_497) + $signed(buffer_7_498); // @[Modules.scala 166:64:@25590.4]
  assign _T_78670 = _T_78669[13:0]; // @[Modules.scala 166:64:@25591.4]
  assign buffer_7_557 = $signed(_T_78670); // @[Modules.scala 166:64:@25592.4]
  assign _T_78672 = $signed(buffer_7_499) + $signed(buffer_7_500); // @[Modules.scala 166:64:@25594.4]
  assign _T_78673 = _T_78672[13:0]; // @[Modules.scala 166:64:@25595.4]
  assign buffer_7_558 = $signed(_T_78673); // @[Modules.scala 166:64:@25596.4]
  assign _T_78675 = $signed(buffer_7_501) + $signed(buffer_7_502); // @[Modules.scala 166:64:@25598.4]
  assign _T_78676 = _T_78675[13:0]; // @[Modules.scala 166:64:@25599.4]
  assign buffer_7_559 = $signed(_T_78676); // @[Modules.scala 166:64:@25600.4]
  assign _T_78678 = $signed(buffer_7_503) + $signed(buffer_7_504); // @[Modules.scala 166:64:@25602.4]
  assign _T_78679 = _T_78678[13:0]; // @[Modules.scala 166:64:@25603.4]
  assign buffer_7_560 = $signed(_T_78679); // @[Modules.scala 166:64:@25604.4]
  assign _T_78681 = $signed(buffer_7_505) + $signed(buffer_7_506); // @[Modules.scala 166:64:@25606.4]
  assign _T_78682 = _T_78681[13:0]; // @[Modules.scala 166:64:@25607.4]
  assign buffer_7_561 = $signed(_T_78682); // @[Modules.scala 166:64:@25608.4]
  assign _T_78684 = $signed(buffer_7_507) + $signed(buffer_7_508); // @[Modules.scala 166:64:@25610.4]
  assign _T_78685 = _T_78684[13:0]; // @[Modules.scala 166:64:@25611.4]
  assign buffer_7_562 = $signed(_T_78685); // @[Modules.scala 166:64:@25612.4]
  assign _T_78687 = $signed(buffer_7_509) + $signed(buffer_7_510); // @[Modules.scala 166:64:@25614.4]
  assign _T_78688 = _T_78687[13:0]; // @[Modules.scala 166:64:@25615.4]
  assign buffer_7_563 = $signed(_T_78688); // @[Modules.scala 166:64:@25616.4]
  assign _T_78690 = $signed(buffer_7_511) + $signed(buffer_7_512); // @[Modules.scala 166:64:@25618.4]
  assign _T_78691 = _T_78690[13:0]; // @[Modules.scala 166:64:@25619.4]
  assign buffer_7_564 = $signed(_T_78691); // @[Modules.scala 166:64:@25620.4]
  assign _T_78693 = $signed(buffer_7_513) + $signed(buffer_7_514); // @[Modules.scala 166:64:@25622.4]
  assign _T_78694 = _T_78693[13:0]; // @[Modules.scala 166:64:@25623.4]
  assign buffer_7_565 = $signed(_T_78694); // @[Modules.scala 166:64:@25624.4]
  assign _T_78696 = $signed(buffer_7_515) + $signed(buffer_7_516); // @[Modules.scala 166:64:@25626.4]
  assign _T_78697 = _T_78696[13:0]; // @[Modules.scala 166:64:@25627.4]
  assign buffer_7_566 = $signed(_T_78697); // @[Modules.scala 166:64:@25628.4]
  assign _T_78699 = $signed(buffer_7_517) + $signed(buffer_7_518); // @[Modules.scala 166:64:@25630.4]
  assign _T_78700 = _T_78699[13:0]; // @[Modules.scala 166:64:@25631.4]
  assign buffer_7_567 = $signed(_T_78700); // @[Modules.scala 166:64:@25632.4]
  assign _T_78702 = $signed(buffer_7_519) + $signed(buffer_7_520); // @[Modules.scala 166:64:@25634.4]
  assign _T_78703 = _T_78702[13:0]; // @[Modules.scala 166:64:@25635.4]
  assign buffer_7_568 = $signed(_T_78703); // @[Modules.scala 166:64:@25636.4]
  assign _T_78705 = $signed(buffer_7_521) + $signed(buffer_7_522); // @[Modules.scala 166:64:@25638.4]
  assign _T_78706 = _T_78705[13:0]; // @[Modules.scala 166:64:@25639.4]
  assign buffer_7_569 = $signed(_T_78706); // @[Modules.scala 166:64:@25640.4]
  assign _T_78708 = $signed(buffer_7_523) + $signed(buffer_7_524); // @[Modules.scala 166:64:@25642.4]
  assign _T_78709 = _T_78708[13:0]; // @[Modules.scala 166:64:@25643.4]
  assign buffer_7_570 = $signed(_T_78709); // @[Modules.scala 166:64:@25644.4]
  assign _T_78711 = $signed(buffer_7_525) + $signed(buffer_7_526); // @[Modules.scala 166:64:@25646.4]
  assign _T_78712 = _T_78711[13:0]; // @[Modules.scala 166:64:@25647.4]
  assign buffer_7_571 = $signed(_T_78712); // @[Modules.scala 166:64:@25648.4]
  assign _T_78714 = $signed(buffer_7_527) + $signed(buffer_7_528); // @[Modules.scala 166:64:@25650.4]
  assign _T_78715 = _T_78714[13:0]; // @[Modules.scala 166:64:@25651.4]
  assign buffer_7_572 = $signed(_T_78715); // @[Modules.scala 166:64:@25652.4]
  assign _T_78717 = $signed(buffer_7_529) + $signed(buffer_7_530); // @[Modules.scala 166:64:@25654.4]
  assign _T_78718 = _T_78717[13:0]; // @[Modules.scala 166:64:@25655.4]
  assign buffer_7_573 = $signed(_T_78718); // @[Modules.scala 166:64:@25656.4]
  assign _T_78720 = $signed(buffer_7_531) + $signed(buffer_7_532); // @[Modules.scala 166:64:@25658.4]
  assign _T_78721 = _T_78720[13:0]; // @[Modules.scala 166:64:@25659.4]
  assign buffer_7_574 = $signed(_T_78721); // @[Modules.scala 166:64:@25660.4]
  assign _T_78723 = $signed(buffer_7_533) + $signed(buffer_7_534); // @[Modules.scala 166:64:@25662.4]
  assign _T_78724 = _T_78723[13:0]; // @[Modules.scala 166:64:@25663.4]
  assign buffer_7_575 = $signed(_T_78724); // @[Modules.scala 166:64:@25664.4]
  assign _T_78726 = $signed(buffer_7_535) + $signed(buffer_7_536); // @[Modules.scala 166:64:@25666.4]
  assign _T_78727 = _T_78726[13:0]; // @[Modules.scala 166:64:@25667.4]
  assign buffer_7_576 = $signed(_T_78727); // @[Modules.scala 166:64:@25668.4]
  assign _T_78729 = $signed(buffer_7_537) + $signed(buffer_7_538); // @[Modules.scala 166:64:@25670.4]
  assign _T_78730 = _T_78729[13:0]; // @[Modules.scala 166:64:@25671.4]
  assign buffer_7_577 = $signed(_T_78730); // @[Modules.scala 166:64:@25672.4]
  assign buffer_7_308 = {{8{_T_77924[5]}},_T_77924}; // @[Modules.scala 112:22:@8.4]
  assign _T_78732 = $signed(buffer_7_539) + $signed(buffer_7_308); // @[Modules.scala 172:66:@25674.4]
  assign _T_78733 = _T_78732[13:0]; // @[Modules.scala 172:66:@25675.4]
  assign buffer_7_578 = $signed(_T_78733); // @[Modules.scala 172:66:@25676.4]
  assign _T_78735 = $signed(buffer_7_540) + $signed(buffer_7_541); // @[Modules.scala 166:64:@25678.4]
  assign _T_78736 = _T_78735[13:0]; // @[Modules.scala 166:64:@25679.4]
  assign buffer_7_579 = $signed(_T_78736); // @[Modules.scala 166:64:@25680.4]
  assign _T_78738 = $signed(buffer_7_542) + $signed(buffer_7_543); // @[Modules.scala 166:64:@25682.4]
  assign _T_78739 = _T_78738[13:0]; // @[Modules.scala 166:64:@25683.4]
  assign buffer_7_580 = $signed(_T_78739); // @[Modules.scala 166:64:@25684.4]
  assign _T_78741 = $signed(buffer_7_544) + $signed(buffer_7_545); // @[Modules.scala 166:64:@25686.4]
  assign _T_78742 = _T_78741[13:0]; // @[Modules.scala 166:64:@25687.4]
  assign buffer_7_581 = $signed(_T_78742); // @[Modules.scala 166:64:@25688.4]
  assign _T_78744 = $signed(buffer_7_546) + $signed(buffer_7_547); // @[Modules.scala 166:64:@25690.4]
  assign _T_78745 = _T_78744[13:0]; // @[Modules.scala 166:64:@25691.4]
  assign buffer_7_582 = $signed(_T_78745); // @[Modules.scala 166:64:@25692.4]
  assign _T_78747 = $signed(buffer_7_548) + $signed(buffer_7_549); // @[Modules.scala 166:64:@25694.4]
  assign _T_78748 = _T_78747[13:0]; // @[Modules.scala 166:64:@25695.4]
  assign buffer_7_583 = $signed(_T_78748); // @[Modules.scala 166:64:@25696.4]
  assign _T_78750 = $signed(buffer_7_550) + $signed(buffer_7_551); // @[Modules.scala 166:64:@25698.4]
  assign _T_78751 = _T_78750[13:0]; // @[Modules.scala 166:64:@25699.4]
  assign buffer_7_584 = $signed(_T_78751); // @[Modules.scala 166:64:@25700.4]
  assign _T_78753 = $signed(buffer_7_552) + $signed(buffer_7_553); // @[Modules.scala 166:64:@25702.4]
  assign _T_78754 = _T_78753[13:0]; // @[Modules.scala 166:64:@25703.4]
  assign buffer_7_585 = $signed(_T_78754); // @[Modules.scala 166:64:@25704.4]
  assign _T_78756 = $signed(buffer_7_554) + $signed(buffer_7_555); // @[Modules.scala 166:64:@25706.4]
  assign _T_78757 = _T_78756[13:0]; // @[Modules.scala 166:64:@25707.4]
  assign buffer_7_586 = $signed(_T_78757); // @[Modules.scala 166:64:@25708.4]
  assign _T_78759 = $signed(buffer_7_556) + $signed(buffer_7_557); // @[Modules.scala 166:64:@25710.4]
  assign _T_78760 = _T_78759[13:0]; // @[Modules.scala 166:64:@25711.4]
  assign buffer_7_587 = $signed(_T_78760); // @[Modules.scala 166:64:@25712.4]
  assign _T_78762 = $signed(buffer_7_558) + $signed(buffer_7_559); // @[Modules.scala 166:64:@25714.4]
  assign _T_78763 = _T_78762[13:0]; // @[Modules.scala 166:64:@25715.4]
  assign buffer_7_588 = $signed(_T_78763); // @[Modules.scala 166:64:@25716.4]
  assign _T_78765 = $signed(buffer_7_560) + $signed(buffer_7_561); // @[Modules.scala 166:64:@25718.4]
  assign _T_78766 = _T_78765[13:0]; // @[Modules.scala 166:64:@25719.4]
  assign buffer_7_589 = $signed(_T_78766); // @[Modules.scala 166:64:@25720.4]
  assign _T_78768 = $signed(buffer_7_562) + $signed(buffer_7_563); // @[Modules.scala 166:64:@25722.4]
  assign _T_78769 = _T_78768[13:0]; // @[Modules.scala 166:64:@25723.4]
  assign buffer_7_590 = $signed(_T_78769); // @[Modules.scala 166:64:@25724.4]
  assign _T_78771 = $signed(buffer_7_564) + $signed(buffer_7_565); // @[Modules.scala 166:64:@25726.4]
  assign _T_78772 = _T_78771[13:0]; // @[Modules.scala 166:64:@25727.4]
  assign buffer_7_591 = $signed(_T_78772); // @[Modules.scala 166:64:@25728.4]
  assign _T_78774 = $signed(buffer_7_566) + $signed(buffer_7_567); // @[Modules.scala 166:64:@25730.4]
  assign _T_78775 = _T_78774[13:0]; // @[Modules.scala 166:64:@25731.4]
  assign buffer_7_592 = $signed(_T_78775); // @[Modules.scala 166:64:@25732.4]
  assign _T_78777 = $signed(buffer_7_568) + $signed(buffer_7_569); // @[Modules.scala 166:64:@25734.4]
  assign _T_78778 = _T_78777[13:0]; // @[Modules.scala 166:64:@25735.4]
  assign buffer_7_593 = $signed(_T_78778); // @[Modules.scala 166:64:@25736.4]
  assign _T_78780 = $signed(buffer_7_570) + $signed(buffer_7_571); // @[Modules.scala 166:64:@25738.4]
  assign _T_78781 = _T_78780[13:0]; // @[Modules.scala 166:64:@25739.4]
  assign buffer_7_594 = $signed(_T_78781); // @[Modules.scala 166:64:@25740.4]
  assign _T_78783 = $signed(buffer_7_572) + $signed(buffer_7_573); // @[Modules.scala 166:64:@25742.4]
  assign _T_78784 = _T_78783[13:0]; // @[Modules.scala 166:64:@25743.4]
  assign buffer_7_595 = $signed(_T_78784); // @[Modules.scala 166:64:@25744.4]
  assign _T_78786 = $signed(buffer_7_574) + $signed(buffer_7_575); // @[Modules.scala 166:64:@25746.4]
  assign _T_78787 = _T_78786[13:0]; // @[Modules.scala 166:64:@25747.4]
  assign buffer_7_596 = $signed(_T_78787); // @[Modules.scala 166:64:@25748.4]
  assign _T_78789 = $signed(buffer_7_576) + $signed(buffer_7_577); // @[Modules.scala 166:64:@25750.4]
  assign _T_78790 = _T_78789[13:0]; // @[Modules.scala 166:64:@25751.4]
  assign buffer_7_597 = $signed(_T_78790); // @[Modules.scala 166:64:@25752.4]
  assign _T_78792 = $signed(buffer_7_579) + $signed(buffer_7_580); // @[Modules.scala 166:64:@25754.4]
  assign _T_78793 = _T_78792[13:0]; // @[Modules.scala 166:64:@25755.4]
  assign buffer_7_598 = $signed(_T_78793); // @[Modules.scala 166:64:@25756.4]
  assign _T_78795 = $signed(buffer_7_581) + $signed(buffer_7_582); // @[Modules.scala 166:64:@25758.4]
  assign _T_78796 = _T_78795[13:0]; // @[Modules.scala 166:64:@25759.4]
  assign buffer_7_599 = $signed(_T_78796); // @[Modules.scala 166:64:@25760.4]
  assign _T_78798 = $signed(buffer_7_583) + $signed(buffer_7_584); // @[Modules.scala 166:64:@25762.4]
  assign _T_78799 = _T_78798[13:0]; // @[Modules.scala 166:64:@25763.4]
  assign buffer_7_600 = $signed(_T_78799); // @[Modules.scala 166:64:@25764.4]
  assign _T_78801 = $signed(buffer_7_585) + $signed(buffer_7_586); // @[Modules.scala 166:64:@25766.4]
  assign _T_78802 = _T_78801[13:0]; // @[Modules.scala 166:64:@25767.4]
  assign buffer_7_601 = $signed(_T_78802); // @[Modules.scala 166:64:@25768.4]
  assign _T_78804 = $signed(buffer_7_587) + $signed(buffer_7_588); // @[Modules.scala 166:64:@25770.4]
  assign _T_78805 = _T_78804[13:0]; // @[Modules.scala 166:64:@25771.4]
  assign buffer_7_602 = $signed(_T_78805); // @[Modules.scala 166:64:@25772.4]
  assign _T_78807 = $signed(buffer_7_589) + $signed(buffer_7_590); // @[Modules.scala 166:64:@25774.4]
  assign _T_78808 = _T_78807[13:0]; // @[Modules.scala 166:64:@25775.4]
  assign buffer_7_603 = $signed(_T_78808); // @[Modules.scala 166:64:@25776.4]
  assign _T_78810 = $signed(buffer_7_591) + $signed(buffer_7_592); // @[Modules.scala 166:64:@25778.4]
  assign _T_78811 = _T_78810[13:0]; // @[Modules.scala 166:64:@25779.4]
  assign buffer_7_604 = $signed(_T_78811); // @[Modules.scala 166:64:@25780.4]
  assign _T_78813 = $signed(buffer_7_593) + $signed(buffer_7_594); // @[Modules.scala 166:64:@25782.4]
  assign _T_78814 = _T_78813[13:0]; // @[Modules.scala 166:64:@25783.4]
  assign buffer_7_605 = $signed(_T_78814); // @[Modules.scala 166:64:@25784.4]
  assign _T_78816 = $signed(buffer_7_595) + $signed(buffer_7_596); // @[Modules.scala 166:64:@25786.4]
  assign _T_78817 = _T_78816[13:0]; // @[Modules.scala 166:64:@25787.4]
  assign buffer_7_606 = $signed(_T_78817); // @[Modules.scala 166:64:@25788.4]
  assign _T_78819 = $signed(buffer_7_597) + $signed(buffer_7_578); // @[Modules.scala 172:66:@25790.4]
  assign _T_78820 = _T_78819[13:0]; // @[Modules.scala 172:66:@25791.4]
  assign buffer_7_607 = $signed(_T_78820); // @[Modules.scala 172:66:@25792.4]
  assign _T_78822 = $signed(buffer_7_598) + $signed(buffer_7_599); // @[Modules.scala 160:64:@25794.4]
  assign _T_78823 = _T_78822[13:0]; // @[Modules.scala 160:64:@25795.4]
  assign buffer_7_608 = $signed(_T_78823); // @[Modules.scala 160:64:@25796.4]
  assign _T_78825 = $signed(buffer_7_600) + $signed(buffer_7_601); // @[Modules.scala 160:64:@25798.4]
  assign _T_78826 = _T_78825[13:0]; // @[Modules.scala 160:64:@25799.4]
  assign buffer_7_609 = $signed(_T_78826); // @[Modules.scala 160:64:@25800.4]
  assign _T_78828 = $signed(buffer_7_602) + $signed(buffer_7_603); // @[Modules.scala 160:64:@25802.4]
  assign _T_78829 = _T_78828[13:0]; // @[Modules.scala 160:64:@25803.4]
  assign buffer_7_610 = $signed(_T_78829); // @[Modules.scala 160:64:@25804.4]
  assign _T_78831 = $signed(buffer_7_604) + $signed(buffer_7_605); // @[Modules.scala 160:64:@25806.4]
  assign _T_78832 = _T_78831[13:0]; // @[Modules.scala 160:64:@25807.4]
  assign buffer_7_611 = $signed(_T_78832); // @[Modules.scala 160:64:@25808.4]
  assign _T_78834 = $signed(buffer_7_606) + $signed(buffer_7_607); // @[Modules.scala 160:64:@25810.4]
  assign _T_78835 = _T_78834[13:0]; // @[Modules.scala 160:64:@25811.4]
  assign buffer_7_612 = $signed(_T_78835); // @[Modules.scala 160:64:@25812.4]
  assign _T_78837 = $signed(buffer_7_608) + $signed(buffer_7_609); // @[Modules.scala 166:64:@25814.4]
  assign _T_78838 = _T_78837[13:0]; // @[Modules.scala 166:64:@25815.4]
  assign buffer_7_613 = $signed(_T_78838); // @[Modules.scala 166:64:@25816.4]
  assign _T_78840 = $signed(buffer_7_610) + $signed(buffer_7_611); // @[Modules.scala 166:64:@25818.4]
  assign _T_78841 = _T_78840[13:0]; // @[Modules.scala 166:64:@25819.4]
  assign buffer_7_614 = $signed(_T_78841); // @[Modules.scala 166:64:@25820.4]
  assign _T_78843 = $signed(buffer_7_613) + $signed(buffer_7_614); // @[Modules.scala 160:64:@25822.4]
  assign _T_78844 = _T_78843[13:0]; // @[Modules.scala 160:64:@25823.4]
  assign buffer_7_615 = $signed(_T_78844); // @[Modules.scala 160:64:@25824.4]
  assign _T_78846 = $signed(buffer_7_615) + $signed(buffer_7_612); // @[Modules.scala 172:66:@25826.4]
  assign _T_78847 = _T_78846[13:0]; // @[Modules.scala 172:66:@25827.4]
  assign buffer_7_616 = $signed(_T_78847); // @[Modules.scala 172:66:@25828.4]
  assign _T_78864 = $signed(4'sh1) * $signed(io_in_25); // @[Modules.scala 143:74:@26009.4]
  assign _T_78866 = $signed(4'sh1) * $signed(io_in_29); // @[Modules.scala 144:80:@26010.4]
  assign _T_78867 = $signed(_T_78864) + $signed(_T_78866); // @[Modules.scala 143:103:@26011.4]
  assign _T_78868 = _T_78867[5:0]; // @[Modules.scala 143:103:@26012.4]
  assign _T_78869 = $signed(_T_78868); // @[Modules.scala 143:103:@26013.4]
  assign _GEN_566 = {{1{_T_57241[4]}},_T_57241}; // @[Modules.scala 143:103:@26029.4]
  assign _T_78888 = $signed(_T_54222) + $signed(_GEN_566); // @[Modules.scala 143:103:@26029.4]
  assign _T_78889 = _T_78888[5:0]; // @[Modules.scala 143:103:@26030.4]
  assign _T_78890 = $signed(_T_78889); // @[Modules.scala 143:103:@26031.4]
  assign _T_78909 = $signed(_T_57255) + $signed(_T_57260); // @[Modules.scala 143:103:@26047.4]
  assign _T_78910 = _T_78909[4:0]; // @[Modules.scala 143:103:@26048.4]
  assign _T_78911 = $signed(_T_78910); // @[Modules.scala 143:103:@26049.4]
  assign _GEN_568 = {{1{_T_57276[4]}},_T_57276}; // @[Modules.scala 143:103:@26071.4]
  assign _T_78937 = $signed(_GEN_568) + $signed(_T_54276); // @[Modules.scala 143:103:@26071.4]
  assign _T_78938 = _T_78937[5:0]; // @[Modules.scala 143:103:@26072.4]
  assign _T_78939 = $signed(_T_78938); // @[Modules.scala 143:103:@26073.4]
  assign _GEN_570 = {{1{_T_66605[4]}},_T_66605}; // @[Modules.scala 143:103:@26131.4]
  assign _T_79007 = $signed(_GEN_570) + $signed(_T_54341); // @[Modules.scala 143:103:@26131.4]
  assign _T_79008 = _T_79007[5:0]; // @[Modules.scala 143:103:@26132.4]
  assign _T_79009 = $signed(_T_79008); // @[Modules.scala 143:103:@26133.4]
  assign _GEN_571 = {{1{_T_63492[4]}},_T_63492}; // @[Modules.scala 143:103:@26143.4]
  assign _T_79021 = $signed(_GEN_571) + $signed(_T_66624); // @[Modules.scala 143:103:@26143.4]
  assign _T_79022 = _T_79021[5:0]; // @[Modules.scala 143:103:@26144.4]
  assign _T_79023 = $signed(_T_79022); // @[Modules.scala 143:103:@26145.4]
  assign _T_79091 = $signed(_T_57430) + $signed(_T_57435); // @[Modules.scala 143:103:@26203.4]
  assign _T_79092 = _T_79091[4:0]; // @[Modules.scala 143:103:@26204.4]
  assign _T_79093 = $signed(_T_79092); // @[Modules.scala 143:103:@26205.4]
  assign _T_79098 = $signed(_GEN_503) + $signed(_T_57442); // @[Modules.scala 143:103:@26209.4]
  assign _T_79099 = _T_79098[5:0]; // @[Modules.scala 143:103:@26210.4]
  assign _T_79100 = $signed(_T_79099); // @[Modules.scala 143:103:@26211.4]
  assign _T_79105 = $signed(_GEN_436) + $signed(_T_57449); // @[Modules.scala 143:103:@26215.4]
  assign _T_79106 = _T_79105[5:0]; // @[Modules.scala 143:103:@26216.4]
  assign _T_79107 = $signed(_T_79106); // @[Modules.scala 143:103:@26217.4]
  assign _GEN_575 = {{1{_T_60507[4]}},_T_60507}; // @[Modules.scala 143:103:@26239.4]
  assign _T_79133 = $signed(_T_54472) + $signed(_GEN_575); // @[Modules.scala 143:103:@26239.4]
  assign _T_79134 = _T_79133[5:0]; // @[Modules.scala 143:103:@26240.4]
  assign _T_79135 = $signed(_T_79134); // @[Modules.scala 143:103:@26241.4]
  assign _T_79140 = $signed(_GEN_85) + $signed(_T_54488); // @[Modules.scala 143:103:@26245.4]
  assign _T_79141 = _T_79140[5:0]; // @[Modules.scala 143:103:@26246.4]
  assign _T_79142 = $signed(_T_79141); // @[Modules.scala 143:103:@26247.4]
  assign _GEN_578 = {{1{_T_63683[4]}},_T_63683}; // @[Modules.scala 143:103:@26275.4]
  assign _T_79175 = $signed(_T_57535) + $signed(_GEN_578); // @[Modules.scala 143:103:@26275.4]
  assign _T_79176 = _T_79175[5:0]; // @[Modules.scala 143:103:@26276.4]
  assign _T_79177 = $signed(_T_79176); // @[Modules.scala 143:103:@26277.4]
  assign _GEN_579 = {{1{_T_60577[4]}},_T_60577}; // @[Modules.scala 143:103:@26281.4]
  assign _T_79182 = $signed(_T_54535) + $signed(_GEN_579); // @[Modules.scala 143:103:@26281.4]
  assign _T_79183 = _T_79182[5:0]; // @[Modules.scala 143:103:@26282.4]
  assign _T_79184 = $signed(_T_79183); // @[Modules.scala 143:103:@26283.4]
  assign _T_79189 = $signed(_T_57556) + $signed(_GEN_224); // @[Modules.scala 143:103:@26287.4]
  assign _T_79190 = _T_79189[5:0]; // @[Modules.scala 143:103:@26288.4]
  assign _T_79191 = $signed(_T_79190); // @[Modules.scala 143:103:@26289.4]
  assign _T_79196 = $signed(_GEN_9) + $signed(_T_76122); // @[Modules.scala 143:103:@26293.4]
  assign _T_79197 = _T_79196[5:0]; // @[Modules.scala 143:103:@26294.4]
  assign _T_79198 = $signed(_T_79197); // @[Modules.scala 143:103:@26295.4]
  assign _T_79238 = $signed(_T_60647) + $signed(_T_63772); // @[Modules.scala 143:103:@26329.4]
  assign _T_79239 = _T_79238[4:0]; // @[Modules.scala 143:103:@26330.4]
  assign _T_79240 = $signed(_T_79239); // @[Modules.scala 143:103:@26331.4]
  assign _T_79245 = $signed(_T_54605) + $signed(_T_57626); // @[Modules.scala 143:103:@26335.4]
  assign _T_79246 = _T_79245[5:0]; // @[Modules.scala 143:103:@26336.4]
  assign _T_79247 = $signed(_T_79246); // @[Modules.scala 143:103:@26337.4]
  assign _T_79266 = $signed(_GEN_513) + $signed(_T_69924); // @[Modules.scala 143:103:@26353.4]
  assign _T_79267 = _T_79266[5:0]; // @[Modules.scala 143:103:@26354.4]
  assign _T_79268 = $signed(_T_79267); // @[Modules.scala 143:103:@26355.4]
  assign _T_79273 = $signed(_GEN_293) + $signed(_T_63814); // @[Modules.scala 143:103:@26359.4]
  assign _T_79274 = _T_79273[5:0]; // @[Modules.scala 143:103:@26360.4]
  assign _T_79275 = $signed(_T_79274); // @[Modules.scala 143:103:@26361.4]
  assign _T_79280 = $signed(_T_60698) + $signed(_T_63821); // @[Modules.scala 143:103:@26365.4]
  assign _T_79281 = _T_79280[5:0]; // @[Modules.scala 143:103:@26366.4]
  assign _T_79282 = $signed(_T_79281); // @[Modules.scala 143:103:@26367.4]
  assign _T_79287 = $signed(_T_63823) + $signed(_T_69938); // @[Modules.scala 143:103:@26371.4]
  assign _T_79288 = _T_79287[5:0]; // @[Modules.scala 143:103:@26372.4]
  assign _T_79289 = $signed(_T_79288); // @[Modules.scala 143:103:@26373.4]
  assign _T_79294 = $signed(_GEN_15) + $signed(_T_54661); // @[Modules.scala 143:103:@26377.4]
  assign _T_79295 = _T_79294[5:0]; // @[Modules.scala 143:103:@26378.4]
  assign _T_79296 = $signed(_T_79295); // @[Modules.scala 143:103:@26379.4]
  assign _T_79301 = $signed(_T_54668) + $signed(_GEN_377); // @[Modules.scala 143:103:@26383.4]
  assign _T_79302 = _T_79301[5:0]; // @[Modules.scala 143:103:@26384.4]
  assign _T_79303 = $signed(_T_79302); // @[Modules.scala 143:103:@26385.4]
  assign _GEN_587 = {{1{_T_57701[4]}},_T_57701}; // @[Modules.scala 143:103:@26395.4]
  assign _T_79315 = $signed(_GEN_587) + $signed(_T_69968); // @[Modules.scala 143:103:@26395.4]
  assign _T_79316 = _T_79315[5:0]; // @[Modules.scala 143:103:@26396.4]
  assign _T_79317 = $signed(_T_79316); // @[Modules.scala 143:103:@26397.4]
  assign _GEN_588 = {{1{_T_60747[4]}},_T_60747}; // @[Modules.scala 143:103:@26401.4]
  assign _T_79322 = $signed(_T_69973) + $signed(_GEN_588); // @[Modules.scala 143:103:@26401.4]
  assign _T_79323 = _T_79322[5:0]; // @[Modules.scala 143:103:@26402.4]
  assign _T_79324 = $signed(_T_79323); // @[Modules.scala 143:103:@26403.4]
  assign _GEN_589 = {{1{_T_54696[4]}},_T_54696}; // @[Modules.scala 143:103:@26413.4]
  assign _T_79336 = $signed(_T_57724) + $signed(_GEN_589); // @[Modules.scala 143:103:@26413.4]
  assign _T_79337 = _T_79336[5:0]; // @[Modules.scala 143:103:@26414.4]
  assign _T_79338 = $signed(_T_79337); // @[Modules.scala 143:103:@26415.4]
  assign _T_79343 = $signed(_T_63884) + $signed(_T_57738); // @[Modules.scala 143:103:@26419.4]
  assign _T_79344 = _T_79343[5:0]; // @[Modules.scala 143:103:@26420.4]
  assign _T_79345 = $signed(_T_79344); // @[Modules.scala 143:103:@26421.4]
  assign _T_79350 = $signed(_T_70010) + $signed(_T_63893); // @[Modules.scala 143:103:@26425.4]
  assign _T_79351 = _T_79350[5:0]; // @[Modules.scala 143:103:@26426.4]
  assign _T_79352 = $signed(_T_79351); // @[Modules.scala 143:103:@26427.4]
  assign _T_79371 = $signed(_T_54726) + $signed(_T_70036); // @[Modules.scala 143:103:@26443.4]
  assign _T_79372 = _T_79371[4:0]; // @[Modules.scala 143:103:@26444.4]
  assign _T_79373 = $signed(_T_79372); // @[Modules.scala 143:103:@26445.4]
  assign _GEN_590 = {{1{_T_60817[4]}},_T_60817}; // @[Modules.scala 143:103:@26455.4]
  assign _T_79385 = $signed(_T_54740) + $signed(_GEN_590); // @[Modules.scala 143:103:@26455.4]
  assign _T_79386 = _T_79385[5:0]; // @[Modules.scala 143:103:@26456.4]
  assign _T_79387 = $signed(_T_79386); // @[Modules.scala 143:103:@26457.4]
  assign _T_79392 = $signed(_GEN_95) + $signed(_T_54754); // @[Modules.scala 143:103:@26461.4]
  assign _T_79393 = _T_79392[5:0]; // @[Modules.scala 143:103:@26462.4]
  assign _T_79394 = $signed(_T_79393); // @[Modules.scala 143:103:@26463.4]
  assign _T_79399 = $signed(_T_70057) + $signed(_T_54761); // @[Modules.scala 143:103:@26467.4]
  assign _T_79400 = _T_79399[5:0]; // @[Modules.scala 143:103:@26468.4]
  assign _T_79401 = $signed(_T_79400); // @[Modules.scala 143:103:@26469.4]
  assign _T_79406 = $signed(_T_67053) + $signed(_T_57799); // @[Modules.scala 143:103:@26473.4]
  assign _T_79407 = _T_79406[5:0]; // @[Modules.scala 143:103:@26474.4]
  assign _T_79408 = $signed(_T_79407); // @[Modules.scala 143:103:@26475.4]
  assign _T_79413 = $signed(_T_60845) + $signed(_T_60850); // @[Modules.scala 143:103:@26479.4]
  assign _T_79414 = _T_79413[4:0]; // @[Modules.scala 143:103:@26480.4]
  assign _T_79415 = $signed(_T_79414); // @[Modules.scala 143:103:@26481.4]
  assign _T_79420 = $signed(_T_57808) + $signed(_T_57815); // @[Modules.scala 143:103:@26485.4]
  assign _T_79421 = _T_79420[5:0]; // @[Modules.scala 143:103:@26486.4]
  assign _T_79422 = $signed(_T_79421); // @[Modules.scala 143:103:@26487.4]
  assign _GEN_592 = {{1{_T_54782[4]}},_T_54782}; // @[Modules.scala 143:103:@26491.4]
  assign _T_79427 = $signed(_T_63968) + $signed(_GEN_592); // @[Modules.scala 143:103:@26491.4]
  assign _T_79428 = _T_79427[5:0]; // @[Modules.scala 143:103:@26492.4]
  assign _T_79429 = $signed(_T_79428); // @[Modules.scala 143:103:@26493.4]
  assign _T_79448 = $signed(_T_63989) + $signed(_T_54808); // @[Modules.scala 143:103:@26509.4]
  assign _T_79449 = _T_79448[5:0]; // @[Modules.scala 143:103:@26510.4]
  assign _T_79450 = $signed(_T_79449); // @[Modules.scala 143:103:@26511.4]
  assign _T_79455 = $signed(_T_54810) + $signed(_T_63996); // @[Modules.scala 143:103:@26515.4]
  assign _T_79456 = _T_79455[4:0]; // @[Modules.scala 143:103:@26516.4]
  assign _T_79457 = $signed(_T_79456); // @[Modules.scala 143:103:@26517.4]
  assign _GEN_593 = {{1{_T_60899[4]}},_T_60899}; // @[Modules.scala 143:103:@26521.4]
  assign _T_79462 = $signed(_GEN_593) + $signed(_T_57857); // @[Modules.scala 143:103:@26521.4]
  assign _T_79463 = _T_79462[5:0]; // @[Modules.scala 143:103:@26522.4]
  assign _T_79464 = $signed(_T_79463); // @[Modules.scala 143:103:@26523.4]
  assign _T_79476 = $signed(_T_70143) + $signed(_T_70148); // @[Modules.scala 143:103:@26533.4]
  assign _T_79477 = _T_79476[5:0]; // @[Modules.scala 143:103:@26534.4]
  assign _T_79478 = $signed(_T_79477); // @[Modules.scala 143:103:@26535.4]
  assign _T_79497 = $signed(_T_67130) + $signed(_GEN_22); // @[Modules.scala 143:103:@26551.4]
  assign _T_79498 = _T_79497[5:0]; // @[Modules.scala 143:103:@26552.4]
  assign _T_79499 = $signed(_T_79498); // @[Modules.scala 143:103:@26553.4]
  assign _GEN_595 = {{1{_T_54857[4]}},_T_54857}; // @[Modules.scala 143:103:@26563.4]
  assign _T_79511 = $signed(_T_57890) + $signed(_GEN_595); // @[Modules.scala 143:103:@26563.4]
  assign _T_79512 = _T_79511[5:0]; // @[Modules.scala 143:103:@26564.4]
  assign _T_79513 = $signed(_T_79512); // @[Modules.scala 143:103:@26565.4]
  assign _T_79518 = $signed(_T_57897) + $signed(_T_70192); // @[Modules.scala 143:103:@26569.4]
  assign _T_79519 = _T_79518[5:0]; // @[Modules.scala 143:103:@26570.4]
  assign _T_79520 = $signed(_T_79519); // @[Modules.scala 143:103:@26571.4]
  assign _GEN_596 = {{1{_T_60985[4]}},_T_60985}; // @[Modules.scala 143:103:@26599.4]
  assign _T_79553 = $signed(_T_54901) + $signed(_GEN_596); // @[Modules.scala 143:103:@26599.4]
  assign _T_79554 = _T_79553[5:0]; // @[Modules.scala 143:103:@26600.4]
  assign _T_79555 = $signed(_T_79554); // @[Modules.scala 143:103:@26601.4]
  assign _T_79560 = $signed(_T_57941) + $signed(_T_64103); // @[Modules.scala 143:103:@26605.4]
  assign _T_79561 = _T_79560[5:0]; // @[Modules.scala 143:103:@26606.4]
  assign _T_79562 = $signed(_T_79561); // @[Modules.scala 143:103:@26607.4]
  assign _T_79602 = $signed(_GEN_518) + $signed(_T_57988); // @[Modules.scala 143:103:@26641.4]
  assign _T_79603 = _T_79602[5:0]; // @[Modules.scala 143:103:@26642.4]
  assign _T_79604 = $signed(_T_79603); // @[Modules.scala 143:103:@26643.4]
  assign _T_79609 = $signed(_T_54964) + $signed(_T_54971); // @[Modules.scala 143:103:@26647.4]
  assign _T_79610 = _T_79609[4:0]; // @[Modules.scala 143:103:@26648.4]
  assign _T_79611 = $signed(_T_79610); // @[Modules.scala 143:103:@26649.4]
  assign _T_79623 = $signed(_T_64171) + $signed(_T_58009); // @[Modules.scala 143:103:@26659.4]
  assign _T_79624 = _T_79623[5:0]; // @[Modules.scala 143:103:@26660.4]
  assign _T_79625 = $signed(_T_79624); // @[Modules.scala 143:103:@26661.4]
  assign _T_79630 = $signed(_T_58011) + $signed(_T_58018); // @[Modules.scala 143:103:@26665.4]
  assign _T_79631 = _T_79630[5:0]; // @[Modules.scala 143:103:@26666.4]
  assign _T_79632 = $signed(_T_79631); // @[Modules.scala 143:103:@26667.4]
  assign _GEN_598 = {{1{_T_61069[4]}},_T_61069}; // @[Modules.scala 143:103:@26671.4]
  assign _T_79637 = $signed(_GEN_598) + $signed(_T_58025); // @[Modules.scala 143:103:@26671.4]
  assign _T_79638 = _T_79637[5:0]; // @[Modules.scala 143:103:@26672.4]
  assign _T_79639 = $signed(_T_79638); // @[Modules.scala 143:103:@26673.4]
  assign _T_79721 = $signed(_T_55076) + $signed(_T_55081); // @[Modules.scala 143:103:@26743.4]
  assign _T_79722 = _T_79721[5:0]; // @[Modules.scala 143:103:@26744.4]
  assign _T_79723 = $signed(_T_79722); // @[Modules.scala 143:103:@26745.4]
  assign _T_79784 = $signed(_T_76696) + $signed(_T_55139); // @[Modules.scala 143:103:@26797.4]
  assign _T_79785 = _T_79784[4:0]; // @[Modules.scala 143:103:@26798.4]
  assign _T_79786 = $signed(_T_79785); // @[Modules.scala 143:103:@26799.4]
  assign _T_79896 = $signed(_T_58270) + $signed(_GEN_106); // @[Modules.scala 143:103:@26893.4]
  assign _T_79897 = _T_79896[5:0]; // @[Modules.scala 143:103:@26894.4]
  assign _T_79898 = $signed(_T_79897); // @[Modules.scala 143:103:@26895.4]
  assign _T_79903 = $signed(_T_58282) + $signed(_GEN_242); // @[Modules.scala 143:103:@26899.4]
  assign _T_79904 = _T_79903[5:0]; // @[Modules.scala 143:103:@26900.4]
  assign _T_79905 = $signed(_T_79904); // @[Modules.scala 143:103:@26901.4]
  assign _T_79924 = $signed(_GEN_107) + $signed(_T_61370); // @[Modules.scala 143:103:@26917.4]
  assign _T_79925 = _T_79924[5:0]; // @[Modules.scala 143:103:@26918.4]
  assign _T_79926 = $signed(_T_79925); // @[Modules.scala 143:103:@26919.4]
  assign _T_79938 = $signed(_T_55298) + $signed(_T_61382); // @[Modules.scala 143:103:@26929.4]
  assign _T_79939 = _T_79938[5:0]; // @[Modules.scala 143:103:@26930.4]
  assign _T_79940 = $signed(_T_79939); // @[Modules.scala 143:103:@26931.4]
  assign _T_79945 = $signed(_T_61384) + $signed(_T_55307); // @[Modules.scala 143:103:@26935.4]
  assign _T_79946 = _T_79945[5:0]; // @[Modules.scala 143:103:@26936.4]
  assign _T_79947 = $signed(_T_79946); // @[Modules.scala 143:103:@26937.4]
  assign _T_79952 = $signed(_T_55312) + $signed(_GEN_243); // @[Modules.scala 143:103:@26941.4]
  assign _T_79953 = _T_79952[5:0]; // @[Modules.scala 143:103:@26942.4]
  assign _T_79954 = $signed(_T_79953); // @[Modules.scala 143:103:@26943.4]
  assign _T_79966 = $signed(_T_55321) + $signed(_T_61412); // @[Modules.scala 143:103:@26953.4]
  assign _T_79967 = _T_79966[4:0]; // @[Modules.scala 143:103:@26954.4]
  assign _T_79968 = $signed(_T_79967); // @[Modules.scala 143:103:@26955.4]
  assign _T_79973 = $signed(_GEN_469) + $signed(_T_55335); // @[Modules.scala 143:103:@26959.4]
  assign _T_79974 = _T_79973[5:0]; // @[Modules.scala 143:103:@26960.4]
  assign _T_79975 = $signed(_T_79974); // @[Modules.scala 143:103:@26961.4]
  assign _GEN_607 = {{1{_T_58382[4]}},_T_58382}; // @[Modules.scala 143:103:@26989.4]
  assign _T_80008 = $signed(_GEN_607) + $signed(_T_55363); // @[Modules.scala 143:103:@26989.4]
  assign _T_80009 = _T_80008[5:0]; // @[Modules.scala 143:103:@26990.4]
  assign _T_80010 = $signed(_T_80009); // @[Modules.scala 143:103:@26991.4]
  assign _T_80022 = $signed(_T_55375) + $signed(_T_61466); // @[Modules.scala 143:103:@27001.4]
  assign _T_80023 = _T_80022[5:0]; // @[Modules.scala 143:103:@27002.4]
  assign _T_80024 = $signed(_T_80023); // @[Modules.scala 143:103:@27003.4]
  assign _T_80050 = $signed(_T_58410) + $signed(_T_58415); // @[Modules.scala 143:103:@27025.4]
  assign _T_80051 = _T_80050[4:0]; // @[Modules.scala 143:103:@27026.4]
  assign _T_80052 = $signed(_T_80051); // @[Modules.scala 143:103:@27027.4]
  assign _T_80064 = $signed(_T_58424) + $signed(_T_61503); // @[Modules.scala 143:103:@27037.4]
  assign _T_80065 = _T_80064[5:0]; // @[Modules.scala 143:103:@27038.4]
  assign _T_80066 = $signed(_T_80065); // @[Modules.scala 143:103:@27039.4]
  assign _T_80085 = $signed(_T_58445) + $signed(_T_58450); // @[Modules.scala 143:103:@27055.4]
  assign _T_80086 = _T_80085[4:0]; // @[Modules.scala 143:103:@27056.4]
  assign _T_80087 = $signed(_T_80086); // @[Modules.scala 143:103:@27057.4]
  assign _T_80092 = $signed(_T_58452) + $signed(_T_58457); // @[Modules.scala 143:103:@27061.4]
  assign _T_80093 = _T_80092[4:0]; // @[Modules.scala 143:103:@27062.4]
  assign _T_80094 = $signed(_T_80093); // @[Modules.scala 143:103:@27063.4]
  assign _T_80113 = $signed(_T_55454) + $signed(_T_55459); // @[Modules.scala 143:103:@27079.4]
  assign _T_80114 = _T_80113[5:0]; // @[Modules.scala 143:103:@27080.4]
  assign _T_80115 = $signed(_T_80114); // @[Modules.scala 143:103:@27081.4]
  assign _T_80120 = $signed(_T_61545) + $signed(_GEN_183); // @[Modules.scala 143:103:@27085.4]
  assign _T_80121 = _T_80120[5:0]; // @[Modules.scala 143:103:@27086.4]
  assign _T_80122 = $signed(_T_80121); // @[Modules.scala 143:103:@27087.4]
  assign _T_80169 = $signed(_T_58522) + $signed(_T_58527); // @[Modules.scala 143:103:@27127.4]
  assign _T_80170 = _T_80169[4:0]; // @[Modules.scala 143:103:@27128.4]
  assign _T_80171 = $signed(_T_80170); // @[Modules.scala 143:103:@27129.4]
  assign _T_80176 = $signed(_T_58529) + $signed(_T_55503); // @[Modules.scala 143:103:@27133.4]
  assign _T_80177 = _T_80176[4:0]; // @[Modules.scala 143:103:@27134.4]
  assign _T_80178 = $signed(_T_80177); // @[Modules.scala 143:103:@27135.4]
  assign _T_80183 = $signed(_T_58536) + $signed(_T_58541); // @[Modules.scala 143:103:@27139.4]
  assign _T_80184 = _T_80183[4:0]; // @[Modules.scala 143:103:@27140.4]
  assign _T_80185 = $signed(_T_80184); // @[Modules.scala 143:103:@27141.4]
  assign _GEN_610 = {{1{_T_58543[4]}},_T_58543}; // @[Modules.scala 143:103:@27145.4]
  assign _T_80190 = $signed(_GEN_610) + $signed(_T_55517); // @[Modules.scala 143:103:@27145.4]
  assign _T_80191 = _T_80190[5:0]; // @[Modules.scala 143:103:@27146.4]
  assign _T_80192 = $signed(_T_80191); // @[Modules.scala 143:103:@27147.4]
  assign _T_80232 = $signed(_T_64768) + $signed(_T_61643); // @[Modules.scala 143:103:@27181.4]
  assign _T_80233 = _T_80232[4:0]; // @[Modules.scala 143:103:@27182.4]
  assign _T_80234 = $signed(_T_80233); // @[Modules.scala 143:103:@27183.4]
  assign _T_80239 = $signed(_T_58590) + $signed(_T_55564); // @[Modules.scala 143:103:@27187.4]
  assign _T_80240 = _T_80239[5:0]; // @[Modules.scala 143:103:@27188.4]
  assign _T_80241 = $signed(_T_80240); // @[Modules.scala 143:103:@27189.4]
  assign _T_80246 = $signed(_T_55566) + $signed(_T_55571); // @[Modules.scala 143:103:@27193.4]
  assign _T_80247 = _T_80246[5:0]; // @[Modules.scala 143:103:@27194.4]
  assign _T_80248 = $signed(_T_80247); // @[Modules.scala 143:103:@27195.4]
  assign _T_80274 = $signed(_T_58620) + $signed(_T_58625); // @[Modules.scala 143:103:@27217.4]
  assign _T_80275 = _T_80274[4:0]; // @[Modules.scala 143:103:@27218.4]
  assign _T_80276 = $signed(_T_80275); // @[Modules.scala 143:103:@27219.4]
  assign _T_80281 = $signed(_T_58627) + $signed(_T_70897); // @[Modules.scala 143:103:@27223.4]
  assign _T_80282 = _T_80281[4:0]; // @[Modules.scala 143:103:@27224.4]
  assign _T_80283 = $signed(_T_80282); // @[Modules.scala 143:103:@27225.4]
  assign _T_80288 = $signed(_T_55608) + $signed(_T_55613); // @[Modules.scala 143:103:@27229.4]
  assign _T_80289 = _T_80288[4:0]; // @[Modules.scala 143:103:@27230.4]
  assign _T_80290 = $signed(_T_80289); // @[Modules.scala 143:103:@27231.4]
  assign _T_80301 = $signed(-4'sh1) * $signed(io_in_524); // @[Modules.scala 144:80:@27240.4]
  assign _T_80302 = $signed(_T_64831) + $signed(_T_80301); // @[Modules.scala 143:103:@27241.4]
  assign _T_80303 = _T_80302[4:0]; // @[Modules.scala 143:103:@27242.4]
  assign _T_80304 = $signed(_T_80303); // @[Modules.scala 143:103:@27243.4]
  assign _T_80309 = $signed(_T_64838) + $signed(_T_58639); // @[Modules.scala 143:103:@27247.4]
  assign _T_80310 = _T_80309[4:0]; // @[Modules.scala 143:103:@27248.4]
  assign _T_80311 = $signed(_T_80310); // @[Modules.scala 143:103:@27249.4]
  assign _T_80323 = $signed(_T_58648) + $signed(_T_61725); // @[Modules.scala 143:103:@27259.4]
  assign _T_80324 = _T_80323[4:0]; // @[Modules.scala 143:103:@27260.4]
  assign _T_80325 = $signed(_T_80324); // @[Modules.scala 143:103:@27261.4]
  assign _T_80330 = $signed(_T_58655) + $signed(_T_55650); // @[Modules.scala 143:103:@27265.4]
  assign _T_80331 = _T_80330[5:0]; // @[Modules.scala 143:103:@27266.4]
  assign _T_80332 = $signed(_T_80331); // @[Modules.scala 143:103:@27267.4]
  assign _GEN_612 = {{1{_T_58676[4]}},_T_58676}; // @[Modules.scala 143:103:@27277.4]
  assign _T_80344 = $signed(_T_55662) + $signed(_GEN_612); // @[Modules.scala 143:103:@27277.4]
  assign _T_80345 = _T_80344[5:0]; // @[Modules.scala 143:103:@27278.4]
  assign _T_80346 = $signed(_T_80345); // @[Modules.scala 143:103:@27279.4]
  assign _T_80372 = $signed(_T_61774) + $signed(_T_64906); // @[Modules.scala 143:103:@27301.4]
  assign _T_80373 = _T_80372[4:0]; // @[Modules.scala 143:103:@27302.4]
  assign _T_80374 = $signed(_T_80373); // @[Modules.scala 143:103:@27303.4]
  assign _T_80379 = $signed(_T_58704) + $signed(_T_58709); // @[Modules.scala 143:103:@27307.4]
  assign _T_80380 = _T_80379[4:0]; // @[Modules.scala 143:103:@27308.4]
  assign _T_80381 = $signed(_T_80380); // @[Modules.scala 143:103:@27309.4]
  assign _T_80386 = $signed(_T_58711) + $signed(_T_64920); // @[Modules.scala 143:103:@27313.4]
  assign _T_80387 = _T_80386[4:0]; // @[Modules.scala 143:103:@27314.4]
  assign _T_80388 = $signed(_T_80387); // @[Modules.scala 143:103:@27315.4]
  assign _T_80407 = $signed(_T_58732) + $signed(_T_58737); // @[Modules.scala 143:103:@27331.4]
  assign _T_80408 = _T_80407[4:0]; // @[Modules.scala 143:103:@27332.4]
  assign _T_80409 = $signed(_T_80408); // @[Modules.scala 143:103:@27333.4]
  assign _T_80414 = $signed(_GEN_62) + $signed(_T_61809); // @[Modules.scala 143:103:@27337.4]
  assign _T_80415 = _T_80414[5:0]; // @[Modules.scala 143:103:@27338.4]
  assign _T_80416 = $signed(_T_80415); // @[Modules.scala 143:103:@27339.4]
  assign _T_80435 = $signed(_T_55746) + $signed(_T_64969); // @[Modules.scala 143:103:@27355.4]
  assign _T_80436 = _T_80435[5:0]; // @[Modules.scala 143:103:@27356.4]
  assign _T_80437 = $signed(_T_80436); // @[Modules.scala 143:103:@27357.4]
  assign _T_80442 = $signed(_T_77382) + $signed(_GEN_262); // @[Modules.scala 143:103:@27361.4]
  assign _T_80443 = _T_80442[5:0]; // @[Modules.scala 143:103:@27362.4]
  assign _T_80444 = $signed(_T_80443); // @[Modules.scala 143:103:@27363.4]
  assign _T_80470 = $signed(_T_58781) + $signed(_T_61858); // @[Modules.scala 143:103:@27385.4]
  assign _T_80471 = _T_80470[4:0]; // @[Modules.scala 143:103:@27386.4]
  assign _T_80472 = $signed(_T_80471); // @[Modules.scala 143:103:@27387.4]
  assign _T_80491 = $signed(_T_58802) + $signed(_T_58807); // @[Modules.scala 143:103:@27403.4]
  assign _T_80492 = _T_80491[4:0]; // @[Modules.scala 143:103:@27404.4]
  assign _T_80493 = $signed(_T_80492); // @[Modules.scala 143:103:@27405.4]
  assign _T_80498 = $signed(_T_61879) + $signed(_T_58814); // @[Modules.scala 143:103:@27409.4]
  assign _T_80499 = _T_80498[4:0]; // @[Modules.scala 143:103:@27410.4]
  assign _T_80500 = $signed(_T_80499); // @[Modules.scala 143:103:@27411.4]
  assign _T_80505 = $signed(_GEN_342) + $signed(_T_55797); // @[Modules.scala 143:103:@27415.4]
  assign _T_80506 = _T_80505[5:0]; // @[Modules.scala 143:103:@27416.4]
  assign _T_80507 = $signed(_T_80506); // @[Modules.scala 143:103:@27417.4]
  assign _GEN_616 = {{1{_T_71151[4]}},_T_71151}; // @[Modules.scala 143:103:@27433.4]
  assign _T_80526 = $signed(_T_55816) + $signed(_GEN_616); // @[Modules.scala 143:103:@27433.4]
  assign _T_80527 = _T_80526[5:0]; // @[Modules.scala 143:103:@27434.4]
  assign _T_80528 = $signed(_T_80527); // @[Modules.scala 143:103:@27435.4]
  assign _T_80596 = $signed(_T_55874) + $signed(_T_55881); // @[Modules.scala 143:103:@27493.4]
  assign _T_80597 = _T_80596[5:0]; // @[Modules.scala 143:103:@27494.4]
  assign _T_80598 = $signed(_T_80597); // @[Modules.scala 143:103:@27495.4]
  assign _GEN_617 = {{1{_T_61998[4]}},_T_61998}; // @[Modules.scala 143:103:@27499.4]
  assign _T_80603 = $signed(_T_71221) + $signed(_GEN_617); // @[Modules.scala 143:103:@27499.4]
  assign _T_80604 = _T_80603[5:0]; // @[Modules.scala 143:103:@27500.4]
  assign _T_80605 = $signed(_T_80604); // @[Modules.scala 143:103:@27501.4]
  assign _T_80617 = $signed(_GEN_130) + $signed(_T_71247); // @[Modules.scala 143:103:@27511.4]
  assign _T_80618 = _T_80617[5:0]; // @[Modules.scala 143:103:@27512.4]
  assign _T_80619 = $signed(_T_80618); // @[Modules.scala 143:103:@27513.4]
  assign _T_80624 = $signed(_T_65125) + $signed(_GEN_549); // @[Modules.scala 143:103:@27517.4]
  assign _T_80625 = _T_80624[5:0]; // @[Modules.scala 143:103:@27518.4]
  assign _T_80626 = $signed(_T_80625); // @[Modules.scala 143:103:@27519.4]
  assign _T_80652 = $signed(_T_58949) + $signed(_T_65165); // @[Modules.scala 143:103:@27541.4]
  assign _T_80653 = _T_80652[4:0]; // @[Modules.scala 143:103:@27542.4]
  assign _T_80654 = $signed(_T_80653); // @[Modules.scala 143:103:@27543.4]
  assign _T_80659 = $signed(_T_55949) + $signed(_GEN_551); // @[Modules.scala 143:103:@27547.4]
  assign _T_80660 = _T_80659[5:0]; // @[Modules.scala 143:103:@27548.4]
  assign _T_80661 = $signed(_T_80660); // @[Modules.scala 143:103:@27549.4]
  assign _T_80673 = $signed(_T_58982) + $signed(_GEN_490); // @[Modules.scala 143:103:@27559.4]
  assign _T_80674 = _T_80673[5:0]; // @[Modules.scala 143:103:@27560.4]
  assign _T_80675 = $signed(_T_80674); // @[Modules.scala 143:103:@27561.4]
  assign _T_80680 = $signed(_T_58984) + $signed(_T_71317); // @[Modules.scala 143:103:@27565.4]
  assign _T_80681 = _T_80680[5:0]; // @[Modules.scala 143:103:@27566.4]
  assign _T_80682 = $signed(_T_80681); // @[Modules.scala 143:103:@27567.4]
  assign _T_80708 = $signed(_GEN_349) + $signed(_T_65221); // @[Modules.scala 143:103:@27589.4]
  assign _T_80709 = _T_80708[5:0]; // @[Modules.scala 143:103:@27590.4]
  assign _T_80710 = $signed(_T_80709); // @[Modules.scala 143:103:@27591.4]
  assign _T_80715 = $signed(_T_56019) + $signed(_T_68257); // @[Modules.scala 143:103:@27595.4]
  assign _T_80716 = _T_80715[5:0]; // @[Modules.scala 143:103:@27596.4]
  assign _T_80717 = $signed(_T_80716); // @[Modules.scala 143:103:@27597.4]
  assign _T_80799 = $signed(_GEN_208) + $signed(_T_56112); // @[Modules.scala 143:103:@27667.4]
  assign _T_80800 = _T_80799[5:0]; // @[Modules.scala 143:103:@27668.4]
  assign _T_80801 = $signed(_T_80800); // @[Modules.scala 143:103:@27669.4]
  assign _T_80883 = $signed(_T_62278) + $signed(_GEN_140); // @[Modules.scala 143:103:@27739.4]
  assign _T_80884 = _T_80883[5:0]; // @[Modules.scala 143:103:@27740.4]
  assign _T_80885 = $signed(_T_80884); // @[Modules.scala 143:103:@27741.4]
  assign _GEN_627 = {{1{_T_77802[4]}},_T_77802}; // @[Modules.scala 143:103:@27745.4]
  assign _T_80890 = $signed(_GEN_627) + $signed(_T_59206); // @[Modules.scala 143:103:@27745.4]
  assign _T_80891 = _T_80890[5:0]; // @[Modules.scala 143:103:@27746.4]
  assign _T_80892 = $signed(_T_80891); // @[Modules.scala 143:103:@27747.4]
  assign _T_80943 = $signed(4'sh1) * $signed(io_in_756); // @[Modules.scala 143:74:@27791.4]
  assign _T_80945 = $signed(4'sh1) * $signed(io_in_758); // @[Modules.scala 144:80:@27792.4]
  assign _T_80946 = $signed(_T_80943) + $signed(_T_80945); // @[Modules.scala 143:103:@27793.4]
  assign _T_80947 = _T_80946[5:0]; // @[Modules.scala 143:103:@27794.4]
  assign _T_80948 = $signed(_T_80947); // @[Modules.scala 143:103:@27795.4]
  assign _T_80953 = $signed(_GEN_142) + $signed(_T_59276); // @[Modules.scala 143:103:@27799.4]
  assign _T_80954 = _T_80953[5:0]; // @[Modules.scala 143:103:@27800.4]
  assign _T_80955 = $signed(_T_80954); // @[Modules.scala 143:103:@27801.4]
  assign _GEN_630 = {{1{_T_62392[4]}},_T_62392}; // @[Modules.scala 143:103:@27823.4]
  assign _T_80981 = $signed(_T_56278) + $signed(_GEN_630); // @[Modules.scala 143:103:@27823.4]
  assign _T_80982 = _T_80981[5:0]; // @[Modules.scala 143:103:@27824.4]
  assign _T_80983 = $signed(_T_80982); // @[Modules.scala 143:103:@27825.4]
  assign _GEN_631 = {{1{_T_56292[4]}},_T_56292}; // @[Modules.scala 143:103:@27835.4]
  assign _T_80995 = $signed(_T_59313) + $signed(_GEN_631); // @[Modules.scala 143:103:@27835.4]
  assign _T_80996 = _T_80995[5:0]; // @[Modules.scala 143:103:@27836.4]
  assign _T_80997 = $signed(_T_80996); // @[Modules.scala 143:103:@27837.4]
  assign buffer_8_2 = {{8{_T_78869[5]}},_T_78869}; // @[Modules.scala 112:22:@8.4]
  assign _T_81015 = $signed(buffer_8_2) + $signed(buffer_2_2); // @[Modules.scala 166:64:@27855.4]
  assign _T_81016 = _T_81015[13:0]; // @[Modules.scala 166:64:@27856.4]
  assign buffer_8_310 = $signed(_T_81016); // @[Modules.scala 166:64:@27857.4]
  assign buffer_8_5 = {{8{_T_78890[5]}},_T_78890}; // @[Modules.scala 112:22:@8.4]
  assign _T_81018 = $signed(buffer_2_3) + $signed(buffer_8_5); // @[Modules.scala 166:64:@27859.4]
  assign _T_81019 = _T_81018[13:0]; // @[Modules.scala 166:64:@27860.4]
  assign buffer_8_311 = $signed(_T_81019); // @[Modules.scala 166:64:@27861.4]
  assign _T_81021 = $signed(buffer_5_6) + $signed(buffer_2_6); // @[Modules.scala 166:64:@27863.4]
  assign _T_81022 = _T_81021[13:0]; // @[Modules.scala 166:64:@27864.4]
  assign buffer_8_312 = $signed(_T_81022); // @[Modules.scala 166:64:@27865.4]
  assign buffer_8_8 = {{9{_T_78911[4]}},_T_78911}; // @[Modules.scala 112:22:@8.4]
  assign _T_81024 = $signed(buffer_8_8) + $signed(buffer_3_7); // @[Modules.scala 166:64:@27867.4]
  assign _T_81025 = _T_81024[13:0]; // @[Modules.scala 166:64:@27868.4]
  assign buffer_8_313 = $signed(_T_81025); // @[Modules.scala 166:64:@27869.4]
  assign _T_81027 = $signed(buffer_5_9) + $signed(buffer_3_9); // @[Modules.scala 166:64:@27871.4]
  assign _T_81028 = _T_81027[13:0]; // @[Modules.scala 166:64:@27872.4]
  assign buffer_8_314 = $signed(_T_81028); // @[Modules.scala 166:64:@27873.4]
  assign buffer_8_12 = {{8{_T_78939[5]}},_T_78939}; // @[Modules.scala 112:22:@8.4]
  assign _T_81030 = $signed(buffer_8_12) + $signed(buffer_5_12); // @[Modules.scala 166:64:@27875.4]
  assign _T_81031 = _T_81030[13:0]; // @[Modules.scala 166:64:@27876.4]
  assign buffer_8_315 = $signed(_T_81031); // @[Modules.scala 166:64:@27877.4]
  assign _T_81033 = $signed(buffer_2_12) + $signed(buffer_4_12); // @[Modules.scala 166:64:@27879.4]
  assign _T_81034 = _T_81033[13:0]; // @[Modules.scala 166:64:@27880.4]
  assign buffer_8_316 = $signed(_T_81034); // @[Modules.scala 166:64:@27881.4]
  assign buffer_8_22 = {{8{_T_79009[5]}},_T_79009}; // @[Modules.scala 112:22:@8.4]
  assign _T_81045 = $signed(buffer_8_22) + $signed(buffer_3_20); // @[Modules.scala 166:64:@27895.4]
  assign _T_81046 = _T_81045[13:0]; // @[Modules.scala 166:64:@27896.4]
  assign buffer_8_320 = $signed(_T_81046); // @[Modules.scala 166:64:@27897.4]
  assign buffer_8_24 = {{8{_T_79023[5]}},_T_79023}; // @[Modules.scala 112:22:@8.4]
  assign _T_81048 = $signed(buffer_8_24) + $signed(buffer_0_23); // @[Modules.scala 166:64:@27899.4]
  assign _T_81049 = _T_81048[13:0]; // @[Modules.scala 166:64:@27900.4]
  assign buffer_8_321 = $signed(_T_81049); // @[Modules.scala 166:64:@27901.4]
  assign buffer_8_34 = {{9{_T_79093[4]}},_T_79093}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_35 = {{8{_T_79100[5]}},_T_79100}; // @[Modules.scala 112:22:@8.4]
  assign _T_81063 = $signed(buffer_8_34) + $signed(buffer_8_35); // @[Modules.scala 166:64:@27919.4]
  assign _T_81064 = _T_81063[13:0]; // @[Modules.scala 166:64:@27920.4]
  assign buffer_8_326 = $signed(_T_81064); // @[Modules.scala 166:64:@27921.4]
  assign buffer_8_36 = {{8{_T_79107[5]}},_T_79107}; // @[Modules.scala 112:22:@8.4]
  assign _T_81066 = $signed(buffer_8_36) + $signed(buffer_4_34); // @[Modules.scala 166:64:@27923.4]
  assign _T_81067 = _T_81066[13:0]; // @[Modules.scala 166:64:@27924.4]
  assign buffer_8_327 = $signed(_T_81067); // @[Modules.scala 166:64:@27925.4]
  assign _T_81069 = $signed(buffer_1_35) + $signed(buffer_7_38); // @[Modules.scala 166:64:@27927.4]
  assign _T_81070 = _T_81069[13:0]; // @[Modules.scala 166:64:@27928.4]
  assign buffer_8_328 = $signed(_T_81070); // @[Modules.scala 166:64:@27929.4]
  assign buffer_8_40 = {{8{_T_79135[5]}},_T_79135}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_41 = {{8{_T_79142[5]}},_T_79142}; // @[Modules.scala 112:22:@8.4]
  assign _T_81072 = $signed(buffer_8_40) + $signed(buffer_8_41); // @[Modules.scala 166:64:@27931.4]
  assign _T_81073 = _T_81072[13:0]; // @[Modules.scala 166:64:@27932.4]
  assign buffer_8_329 = $signed(_T_81073); // @[Modules.scala 166:64:@27933.4]
  assign _T_81075 = $signed(buffer_0_42) + $signed(buffer_3_44); // @[Modules.scala 166:64:@27935.4]
  assign _T_81076 = _T_81075[13:0]; // @[Modules.scala 166:64:@27936.4]
  assign buffer_8_330 = $signed(_T_81076); // @[Modules.scala 166:64:@27937.4]
  assign buffer_8_46 = {{8{_T_79177[5]}},_T_79177}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_47 = {{8{_T_79184[5]}},_T_79184}; // @[Modules.scala 112:22:@8.4]
  assign _T_81081 = $signed(buffer_8_46) + $signed(buffer_8_47); // @[Modules.scala 166:64:@27943.4]
  assign _T_81082 = _T_81081[13:0]; // @[Modules.scala 166:64:@27944.4]
  assign buffer_8_332 = $signed(_T_81082); // @[Modules.scala 166:64:@27945.4]
  assign buffer_8_48 = {{8{_T_79191[5]}},_T_79191}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_49 = {{8{_T_79198[5]}},_T_79198}; // @[Modules.scala 112:22:@8.4]
  assign _T_81084 = $signed(buffer_8_48) + $signed(buffer_8_49); // @[Modules.scala 166:64:@27947.4]
  assign _T_81085 = _T_81084[13:0]; // @[Modules.scala 166:64:@27948.4]
  assign buffer_8_333 = $signed(_T_81085); // @[Modules.scala 166:64:@27949.4]
  assign _T_81087 = $signed(buffer_5_53) + $signed(buffer_7_53); // @[Modules.scala 166:64:@27951.4]
  assign _T_81088 = _T_81087[13:0]; // @[Modules.scala 166:64:@27952.4]
  assign buffer_8_334 = $signed(_T_81088); // @[Modules.scala 166:64:@27953.4]
  assign _T_81090 = $signed(buffer_7_54) + $signed(buffer_0_55); // @[Modules.scala 166:64:@27955.4]
  assign _T_81091 = _T_81090[13:0]; // @[Modules.scala 166:64:@27956.4]
  assign buffer_8_335 = $signed(_T_81091); // @[Modules.scala 166:64:@27957.4]
  assign buffer_8_55 = {{9{_T_79240[4]}},_T_79240}; // @[Modules.scala 112:22:@8.4]
  assign _T_81093 = $signed(buffer_5_58) + $signed(buffer_8_55); // @[Modules.scala 166:64:@27959.4]
  assign _T_81094 = _T_81093[13:0]; // @[Modules.scala 166:64:@27960.4]
  assign buffer_8_336 = $signed(_T_81094); // @[Modules.scala 166:64:@27961.4]
  assign buffer_8_56 = {{8{_T_79247[5]}},_T_79247}; // @[Modules.scala 112:22:@8.4]
  assign _T_81096 = $signed(buffer_8_56) + $signed(buffer_0_59); // @[Modules.scala 166:64:@27963.4]
  assign _T_81097 = _T_81096[13:0]; // @[Modules.scala 166:64:@27964.4]
  assign buffer_8_337 = $signed(_T_81097); // @[Modules.scala 166:64:@27965.4]
  assign buffer_8_59 = {{8{_T_79268[5]}},_T_79268}; // @[Modules.scala 112:22:@8.4]
  assign _T_81099 = $signed(buffer_2_61) + $signed(buffer_8_59); // @[Modules.scala 166:64:@27967.4]
  assign _T_81100 = _T_81099[13:0]; // @[Modules.scala 166:64:@27968.4]
  assign buffer_8_338 = $signed(_T_81100); // @[Modules.scala 166:64:@27969.4]
  assign buffer_8_60 = {{8{_T_79275[5]}},_T_79275}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_61 = {{8{_T_79282[5]}},_T_79282}; // @[Modules.scala 112:22:@8.4]
  assign _T_81102 = $signed(buffer_8_60) + $signed(buffer_8_61); // @[Modules.scala 166:64:@27971.4]
  assign _T_81103 = _T_81102[13:0]; // @[Modules.scala 166:64:@27972.4]
  assign buffer_8_339 = $signed(_T_81103); // @[Modules.scala 166:64:@27973.4]
  assign buffer_8_62 = {{8{_T_79289[5]}},_T_79289}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_63 = {{8{_T_79296[5]}},_T_79296}; // @[Modules.scala 112:22:@8.4]
  assign _T_81105 = $signed(buffer_8_62) + $signed(buffer_8_63); // @[Modules.scala 166:64:@27975.4]
  assign _T_81106 = _T_81105[13:0]; // @[Modules.scala 166:64:@27976.4]
  assign buffer_8_340 = $signed(_T_81106); // @[Modules.scala 166:64:@27977.4]
  assign buffer_8_64 = {{8{_T_79303[5]}},_T_79303}; // @[Modules.scala 112:22:@8.4]
  assign _T_81108 = $signed(buffer_8_64) + $signed(buffer_2_68); // @[Modules.scala 166:64:@27979.4]
  assign _T_81109 = _T_81108[13:0]; // @[Modules.scala 166:64:@27980.4]
  assign buffer_8_341 = $signed(_T_81109); // @[Modules.scala 166:64:@27981.4]
  assign buffer_8_66 = {{8{_T_79317[5]}},_T_79317}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_67 = {{8{_T_79324[5]}},_T_79324}; // @[Modules.scala 112:22:@8.4]
  assign _T_81111 = $signed(buffer_8_66) + $signed(buffer_8_67); // @[Modules.scala 166:64:@27983.4]
  assign _T_81112 = _T_81111[13:0]; // @[Modules.scala 166:64:@27984.4]
  assign buffer_8_342 = $signed(_T_81112); // @[Modules.scala 166:64:@27985.4]
  assign buffer_8_69 = {{8{_T_79338[5]}},_T_79338}; // @[Modules.scala 112:22:@8.4]
  assign _T_81114 = $signed(buffer_2_72) + $signed(buffer_8_69); // @[Modules.scala 166:64:@27987.4]
  assign _T_81115 = _T_81114[13:0]; // @[Modules.scala 166:64:@27988.4]
  assign buffer_8_343 = $signed(_T_81115); // @[Modules.scala 166:64:@27989.4]
  assign buffer_8_70 = {{8{_T_79345[5]}},_T_79345}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_71 = {{8{_T_79352[5]}},_T_79352}; // @[Modules.scala 112:22:@8.4]
  assign _T_81117 = $signed(buffer_8_70) + $signed(buffer_8_71); // @[Modules.scala 166:64:@27991.4]
  assign _T_81118 = _T_81117[13:0]; // @[Modules.scala 166:64:@27992.4]
  assign buffer_8_344 = $signed(_T_81118); // @[Modules.scala 166:64:@27993.4]
  assign buffer_8_74 = {{9{_T_79373[4]}},_T_79373}; // @[Modules.scala 112:22:@8.4]
  assign _T_81123 = $signed(buffer_8_74) + $signed(buffer_1_80); // @[Modules.scala 166:64:@27999.4]
  assign _T_81124 = _T_81123[13:0]; // @[Modules.scala 166:64:@28000.4]
  assign buffer_8_346 = $signed(_T_81124); // @[Modules.scala 166:64:@28001.4]
  assign buffer_8_76 = {{8{_T_79387[5]}},_T_79387}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_77 = {{8{_T_79394[5]}},_T_79394}; // @[Modules.scala 112:22:@8.4]
  assign _T_81126 = $signed(buffer_8_76) + $signed(buffer_8_77); // @[Modules.scala 166:64:@28003.4]
  assign _T_81127 = _T_81126[13:0]; // @[Modules.scala 166:64:@28004.4]
  assign buffer_8_347 = $signed(_T_81127); // @[Modules.scala 166:64:@28005.4]
  assign buffer_8_78 = {{8{_T_79401[5]}},_T_79401}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_79 = {{8{_T_79408[5]}},_T_79408}; // @[Modules.scala 112:22:@8.4]
  assign _T_81129 = $signed(buffer_8_78) + $signed(buffer_8_79); // @[Modules.scala 166:64:@28007.4]
  assign _T_81130 = _T_81129[13:0]; // @[Modules.scala 166:64:@28008.4]
  assign buffer_8_348 = $signed(_T_81130); // @[Modules.scala 166:64:@28009.4]
  assign buffer_8_80 = {{9{_T_79415[4]}},_T_79415}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_81 = {{8{_T_79422[5]}},_T_79422}; // @[Modules.scala 112:22:@8.4]
  assign _T_81132 = $signed(buffer_8_80) + $signed(buffer_8_81); // @[Modules.scala 166:64:@28011.4]
  assign _T_81133 = _T_81132[13:0]; // @[Modules.scala 166:64:@28012.4]
  assign buffer_8_349 = $signed(_T_81133); // @[Modules.scala 166:64:@28013.4]
  assign buffer_8_82 = {{8{_T_79429[5]}},_T_79429}; // @[Modules.scala 112:22:@8.4]
  assign _T_81135 = $signed(buffer_8_82) + $signed(buffer_3_90); // @[Modules.scala 166:64:@28015.4]
  assign _T_81136 = _T_81135[13:0]; // @[Modules.scala 166:64:@28016.4]
  assign buffer_8_350 = $signed(_T_81136); // @[Modules.scala 166:64:@28017.4]
  assign buffer_8_85 = {{8{_T_79450[5]}},_T_79450}; // @[Modules.scala 112:22:@8.4]
  assign _T_81138 = $signed(buffer_3_91) + $signed(buffer_8_85); // @[Modules.scala 166:64:@28019.4]
  assign _T_81139 = _T_81138[13:0]; // @[Modules.scala 166:64:@28020.4]
  assign buffer_8_351 = $signed(_T_81139); // @[Modules.scala 166:64:@28021.4]
  assign buffer_8_86 = {{9{_T_79457[4]}},_T_79457}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_87 = {{8{_T_79464[5]}},_T_79464}; // @[Modules.scala 112:22:@8.4]
  assign _T_81141 = $signed(buffer_8_86) + $signed(buffer_8_87); // @[Modules.scala 166:64:@28023.4]
  assign _T_81142 = _T_81141[13:0]; // @[Modules.scala 166:64:@28024.4]
  assign buffer_8_352 = $signed(_T_81142); // @[Modules.scala 166:64:@28025.4]
  assign buffer_8_89 = {{8{_T_79478[5]}},_T_79478}; // @[Modules.scala 112:22:@8.4]
  assign _T_81144 = $signed(buffer_1_93) + $signed(buffer_8_89); // @[Modules.scala 166:64:@28027.4]
  assign _T_81145 = _T_81144[13:0]; // @[Modules.scala 166:64:@28028.4]
  assign buffer_8_353 = $signed(_T_81145); // @[Modules.scala 166:64:@28029.4]
  assign buffer_8_92 = {{8{_T_79499[5]}},_T_79499}; // @[Modules.scala 112:22:@8.4]
  assign _T_81150 = $signed(buffer_8_92) + $signed(buffer_2_98); // @[Modules.scala 166:64:@28035.4]
  assign _T_81151 = _T_81150[13:0]; // @[Modules.scala 166:64:@28036.4]
  assign buffer_8_355 = $signed(_T_81151); // @[Modules.scala 166:64:@28037.4]
  assign buffer_8_94 = {{8{_T_79513[5]}},_T_79513}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_95 = {{8{_T_79520[5]}},_T_79520}; // @[Modules.scala 112:22:@8.4]
  assign _T_81153 = $signed(buffer_8_94) + $signed(buffer_8_95); // @[Modules.scala 166:64:@28039.4]
  assign _T_81154 = _T_81153[13:0]; // @[Modules.scala 166:64:@28040.4]
  assign buffer_8_356 = $signed(_T_81154); // @[Modules.scala 166:64:@28041.4]
  assign _T_81159 = $signed(buffer_5_106) + $signed(buffer_4_101); // @[Modules.scala 166:64:@28047.4]
  assign _T_81160 = _T_81159[13:0]; // @[Modules.scala 166:64:@28048.4]
  assign buffer_8_358 = $signed(_T_81160); // @[Modules.scala 166:64:@28049.4]
  assign buffer_8_100 = {{8{_T_79555[5]}},_T_79555}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_101 = {{8{_T_79562[5]}},_T_79562}; // @[Modules.scala 112:22:@8.4]
  assign _T_81162 = $signed(buffer_8_100) + $signed(buffer_8_101); // @[Modules.scala 166:64:@28051.4]
  assign _T_81163 = _T_81162[13:0]; // @[Modules.scala 166:64:@28052.4]
  assign buffer_8_359 = $signed(_T_81163); // @[Modules.scala 166:64:@28053.4]
  assign _T_81165 = $signed(buffer_3_109) + $signed(buffer_3_110); // @[Modules.scala 166:64:@28055.4]
  assign _T_81166 = _T_81165[13:0]; // @[Modules.scala 166:64:@28056.4]
  assign buffer_8_360 = $signed(_T_81166); // @[Modules.scala 166:64:@28057.4]
  assign _T_81168 = $signed(buffer_3_111) + $signed(buffer_4_106); // @[Modules.scala 166:64:@28059.4]
  assign _T_81169 = _T_81168[13:0]; // @[Modules.scala 166:64:@28060.4]
  assign buffer_8_361 = $signed(_T_81169); // @[Modules.scala 166:64:@28061.4]
  assign buffer_8_107 = {{8{_T_79604[5]}},_T_79604}; // @[Modules.scala 112:22:@8.4]
  assign _T_81171 = $signed(buffer_0_107) + $signed(buffer_8_107); // @[Modules.scala 166:64:@28063.4]
  assign _T_81172 = _T_81171[13:0]; // @[Modules.scala 166:64:@28064.4]
  assign buffer_8_362 = $signed(_T_81172); // @[Modules.scala 166:64:@28065.4]
  assign buffer_8_108 = {{9{_T_79611[4]}},_T_79611}; // @[Modules.scala 112:22:@8.4]
  assign _T_81174 = $signed(buffer_8_108) + $signed(buffer_3_117); // @[Modules.scala 166:64:@28067.4]
  assign _T_81175 = _T_81174[13:0]; // @[Modules.scala 166:64:@28068.4]
  assign buffer_8_363 = $signed(_T_81175); // @[Modules.scala 166:64:@28069.4]
  assign buffer_8_110 = {{8{_T_79625[5]}},_T_79625}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_111 = {{8{_T_79632[5]}},_T_79632}; // @[Modules.scala 112:22:@8.4]
  assign _T_81177 = $signed(buffer_8_110) + $signed(buffer_8_111); // @[Modules.scala 166:64:@28071.4]
  assign _T_81178 = _T_81177[13:0]; // @[Modules.scala 166:64:@28072.4]
  assign buffer_8_364 = $signed(_T_81178); // @[Modules.scala 166:64:@28073.4]
  assign buffer_8_112 = {{8{_T_79639[5]}},_T_79639}; // @[Modules.scala 112:22:@8.4]
  assign _T_81180 = $signed(buffer_8_112) + $signed(buffer_3_122); // @[Modules.scala 166:64:@28075.4]
  assign _T_81181 = _T_81180[13:0]; // @[Modules.scala 166:64:@28076.4]
  assign buffer_8_365 = $signed(_T_81181); // @[Modules.scala 166:64:@28077.4]
  assign _T_81183 = $signed(buffer_3_123) + $signed(buffer_3_124); // @[Modules.scala 166:64:@28079.4]
  assign _T_81184 = _T_81183[13:0]; // @[Modules.scala 166:64:@28080.4]
  assign buffer_8_366 = $signed(_T_81184); // @[Modules.scala 166:64:@28081.4]
  assign _T_81186 = $signed(buffer_3_125) + $signed(buffer_1_121); // @[Modules.scala 166:64:@28083.4]
  assign _T_81187 = _T_81186[13:0]; // @[Modules.scala 166:64:@28084.4]
  assign buffer_8_367 = $signed(_T_81187); // @[Modules.scala 166:64:@28085.4]
  assign _T_81189 = $signed(buffer_1_122) + $signed(buffer_0_121); // @[Modules.scala 166:64:@28087.4]
  assign _T_81190 = _T_81189[13:0]; // @[Modules.scala 166:64:@28088.4]
  assign buffer_8_368 = $signed(_T_81190); // @[Modules.scala 166:64:@28089.4]
  assign _T_81195 = $signed(buffer_3_131) + $signed(buffer_1_127); // @[Modules.scala 166:64:@28095.4]
  assign _T_81196 = _T_81195[13:0]; // @[Modules.scala 166:64:@28096.4]
  assign buffer_8_370 = $signed(_T_81196); // @[Modules.scala 166:64:@28097.4]
  assign buffer_8_124 = {{8{_T_79723[5]}},_T_79723}; // @[Modules.scala 112:22:@8.4]
  assign _T_81198 = $signed(buffer_8_124) + $signed(buffer_1_129); // @[Modules.scala 166:64:@28099.4]
  assign _T_81199 = _T_81198[13:0]; // @[Modules.scala 166:64:@28100.4]
  assign buffer_8_371 = $signed(_T_81199); // @[Modules.scala 166:64:@28101.4]
  assign _T_81201 = $signed(buffer_3_135) + $signed(buffer_2_131); // @[Modules.scala 166:64:@28103.4]
  assign _T_81202 = _T_81201[13:0]; // @[Modules.scala 166:64:@28104.4]
  assign buffer_8_372 = $signed(_T_81202); // @[Modules.scala 166:64:@28105.4]
  assign _T_81207 = $signed(buffer_1_133) + $signed(buffer_1_134); // @[Modules.scala 166:64:@28111.4]
  assign _T_81208 = _T_81207[13:0]; // @[Modules.scala 166:64:@28112.4]
  assign buffer_8_374 = $signed(_T_81208); // @[Modules.scala 166:64:@28113.4]
  assign buffer_8_133 = {{9{_T_79786[4]}},_T_79786}; // @[Modules.scala 112:22:@8.4]
  assign _T_81210 = $signed(buffer_1_135) + $signed(buffer_8_133); // @[Modules.scala 166:64:@28115.4]
  assign _T_81211 = _T_81210[13:0]; // @[Modules.scala 166:64:@28116.4]
  assign buffer_8_375 = $signed(_T_81211); // @[Modules.scala 166:64:@28117.4]
  assign _T_81219 = $signed(buffer_0_139) + $signed(buffer_2_144); // @[Modules.scala 166:64:@28127.4]
  assign _T_81220 = _T_81219[13:0]; // @[Modules.scala 166:64:@28128.4]
  assign buffer_8_378 = $signed(_T_81220); // @[Modules.scala 166:64:@28129.4]
  assign _T_81222 = $signed(buffer_2_145) + $signed(buffer_2_146); // @[Modules.scala 166:64:@28131.4]
  assign _T_81223 = _T_81222[13:0]; // @[Modules.scala 166:64:@28132.4]
  assign buffer_8_379 = $signed(_T_81223); // @[Modules.scala 166:64:@28133.4]
  assign _T_81225 = $signed(buffer_2_147) + $signed(buffer_3_152); // @[Modules.scala 166:64:@28135.4]
  assign _T_81226 = _T_81225[13:0]; // @[Modules.scala 166:64:@28136.4]
  assign buffer_8_380 = $signed(_T_81226); // @[Modules.scala 166:64:@28137.4]
  assign _T_81228 = $signed(buffer_2_149) + $signed(buffer_2_150); // @[Modules.scala 166:64:@28139.4]
  assign _T_81229 = _T_81228[13:0]; // @[Modules.scala 166:64:@28140.4]
  assign buffer_8_381 = $signed(_T_81229); // @[Modules.scala 166:64:@28141.4]
  assign _T_81231 = $signed(buffer_5_147) + $signed(buffer_3_156); // @[Modules.scala 166:64:@28143.4]
  assign _T_81232 = _T_81231[13:0]; // @[Modules.scala 166:64:@28144.4]
  assign buffer_8_382 = $signed(_T_81232); // @[Modules.scala 166:64:@28145.4]
  assign buffer_8_149 = {{8{_T_79898[5]}},_T_79898}; // @[Modules.scala 112:22:@8.4]
  assign _T_81234 = $signed(buffer_3_157) + $signed(buffer_8_149); // @[Modules.scala 166:64:@28147.4]
  assign _T_81235 = _T_81234[13:0]; // @[Modules.scala 166:64:@28148.4]
  assign buffer_8_383 = $signed(_T_81235); // @[Modules.scala 166:64:@28149.4]
  assign buffer_8_150 = {{8{_T_79905[5]}},_T_79905}; // @[Modules.scala 112:22:@8.4]
  assign _T_81237 = $signed(buffer_8_150) + $signed(buffer_7_152); // @[Modules.scala 166:64:@28151.4]
  assign _T_81238 = _T_81237[13:0]; // @[Modules.scala 166:64:@28152.4]
  assign buffer_8_384 = $signed(_T_81238); // @[Modules.scala 166:64:@28153.4]
  assign buffer_8_153 = {{8{_T_79926[5]}},_T_79926}; // @[Modules.scala 112:22:@8.4]
  assign _T_81240 = $signed(buffer_5_153) + $signed(buffer_8_153); // @[Modules.scala 166:64:@28155.4]
  assign _T_81241 = _T_81240[13:0]; // @[Modules.scala 166:64:@28156.4]
  assign buffer_8_385 = $signed(_T_81241); // @[Modules.scala 166:64:@28157.4]
  assign buffer_8_155 = {{8{_T_79940[5]}},_T_79940}; // @[Modules.scala 112:22:@8.4]
  assign _T_81243 = $signed(buffer_1_157) + $signed(buffer_8_155); // @[Modules.scala 166:64:@28159.4]
  assign _T_81244 = _T_81243[13:0]; // @[Modules.scala 166:64:@28160.4]
  assign buffer_8_386 = $signed(_T_81244); // @[Modules.scala 166:64:@28161.4]
  assign buffer_8_156 = {{8{_T_79947[5]}},_T_79947}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_157 = {{8{_T_79954[5]}},_T_79954}; // @[Modules.scala 112:22:@8.4]
  assign _T_81246 = $signed(buffer_8_156) + $signed(buffer_8_157); // @[Modules.scala 166:64:@28163.4]
  assign _T_81247 = _T_81246[13:0]; // @[Modules.scala 166:64:@28164.4]
  assign buffer_8_387 = $signed(_T_81247); // @[Modules.scala 166:64:@28165.4]
  assign buffer_8_159 = {{9{_T_79968[4]}},_T_79968}; // @[Modules.scala 112:22:@8.4]
  assign _T_81249 = $signed(buffer_1_161) + $signed(buffer_8_159); // @[Modules.scala 166:64:@28167.4]
  assign _T_81250 = _T_81249[13:0]; // @[Modules.scala 166:64:@28168.4]
  assign buffer_8_388 = $signed(_T_81250); // @[Modules.scala 166:64:@28169.4]
  assign buffer_8_160 = {{8{_T_79975[5]}},_T_79975}; // @[Modules.scala 112:22:@8.4]
  assign _T_81252 = $signed(buffer_8_160) + $signed(buffer_7_165); // @[Modules.scala 166:64:@28171.4]
  assign _T_81253 = _T_81252[13:0]; // @[Modules.scala 166:64:@28172.4]
  assign buffer_8_389 = $signed(_T_81253); // @[Modules.scala 166:64:@28173.4]
  assign buffer_8_165 = {{8{_T_80010[5]}},_T_80010}; // @[Modules.scala 112:22:@8.4]
  assign _T_81258 = $signed(buffer_7_168) + $signed(buffer_8_165); // @[Modules.scala 166:64:@28179.4]
  assign _T_81259 = _T_81258[13:0]; // @[Modules.scala 166:64:@28180.4]
  assign buffer_8_391 = $signed(_T_81259); // @[Modules.scala 166:64:@28181.4]
  assign buffer_8_167 = {{8{_T_80024[5]}},_T_80024}; // @[Modules.scala 112:22:@8.4]
  assign _T_81261 = $signed(buffer_0_167) + $signed(buffer_8_167); // @[Modules.scala 166:64:@28183.4]
  assign _T_81262 = _T_81261[13:0]; // @[Modules.scala 166:64:@28184.4]
  assign buffer_8_392 = $signed(_T_81262); // @[Modules.scala 166:64:@28185.4]
  assign _T_81264 = $signed(buffer_4_165) + $signed(buffer_4_166); // @[Modules.scala 166:64:@28187.4]
  assign _T_81265 = _T_81264[13:0]; // @[Modules.scala 166:64:@28188.4]
  assign buffer_8_393 = $signed(_T_81265); // @[Modules.scala 166:64:@28189.4]
  assign buffer_8_171 = {{9{_T_80052[4]}},_T_80052}; // @[Modules.scala 112:22:@8.4]
  assign _T_81267 = $signed(buffer_6_177) + $signed(buffer_8_171); // @[Modules.scala 166:64:@28191.4]
  assign _T_81268 = _T_81267[13:0]; // @[Modules.scala 166:64:@28192.4]
  assign buffer_8_394 = $signed(_T_81268); // @[Modules.scala 166:64:@28193.4]
  assign buffer_8_173 = {{8{_T_80066[5]}},_T_80066}; // @[Modules.scala 112:22:@8.4]
  assign _T_81270 = $signed(buffer_2_178) + $signed(buffer_8_173); // @[Modules.scala 166:64:@28195.4]
  assign _T_81271 = _T_81270[13:0]; // @[Modules.scala 166:64:@28196.4]
  assign buffer_8_395 = $signed(_T_81271); // @[Modules.scala 166:64:@28197.4]
  assign _T_81273 = $signed(buffer_0_175) + $signed(buffer_0_176); // @[Modules.scala 166:64:@28199.4]
  assign _T_81274 = _T_81273[13:0]; // @[Modules.scala 166:64:@28200.4]
  assign buffer_8_396 = $signed(_T_81274); // @[Modules.scala 166:64:@28201.4]
  assign buffer_8_176 = {{9{_T_80087[4]}},_T_80087}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_177 = {{9{_T_80094[4]}},_T_80094}; // @[Modules.scala 112:22:@8.4]
  assign _T_81276 = $signed(buffer_8_176) + $signed(buffer_8_177); // @[Modules.scala 166:64:@28203.4]
  assign _T_81277 = _T_81276[13:0]; // @[Modules.scala 166:64:@28204.4]
  assign buffer_8_397 = $signed(_T_81277); // @[Modules.scala 166:64:@28205.4]
  assign buffer_8_180 = {{8{_T_80115[5]}},_T_80115}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_181 = {{8{_T_80122[5]}},_T_80122}; // @[Modules.scala 112:22:@8.4]
  assign _T_81282 = $signed(buffer_8_180) + $signed(buffer_8_181); // @[Modules.scala 166:64:@28211.4]
  assign _T_81283 = _T_81282[13:0]; // @[Modules.scala 166:64:@28212.4]
  assign buffer_8_399 = $signed(_T_81283); // @[Modules.scala 166:64:@28213.4]
  assign _T_81291 = $signed(buffer_6_193) + $signed(buffer_2_192); // @[Modules.scala 166:64:@28223.4]
  assign _T_81292 = _T_81291[13:0]; // @[Modules.scala 166:64:@28224.4]
  assign buffer_8_402 = $signed(_T_81292); // @[Modules.scala 166:64:@28225.4]
  assign buffer_8_188 = {{9{_T_80171[4]}},_T_80171}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_189 = {{9{_T_80178[4]}},_T_80178}; // @[Modules.scala 112:22:@8.4]
  assign _T_81294 = $signed(buffer_8_188) + $signed(buffer_8_189); // @[Modules.scala 166:64:@28227.4]
  assign _T_81295 = _T_81294[13:0]; // @[Modules.scala 166:64:@28228.4]
  assign buffer_8_403 = $signed(_T_81295); // @[Modules.scala 166:64:@28229.4]
  assign buffer_8_190 = {{9{_T_80185[4]}},_T_80185}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_191 = {{8{_T_80192[5]}},_T_80192}; // @[Modules.scala 112:22:@8.4]
  assign _T_81297 = $signed(buffer_8_190) + $signed(buffer_8_191); // @[Modules.scala 166:64:@28231.4]
  assign _T_81298 = _T_81297[13:0]; // @[Modules.scala 166:64:@28232.4]
  assign buffer_8_404 = $signed(_T_81298); // @[Modules.scala 166:64:@28233.4]
  assign _T_81300 = $signed(buffer_3_200) + $signed(buffer_7_198); // @[Modules.scala 166:64:@28235.4]
  assign _T_81301 = _T_81300[13:0]; // @[Modules.scala 166:64:@28236.4]
  assign buffer_8_405 = $signed(_T_81301); // @[Modules.scala 166:64:@28237.4]
  assign _T_81303 = $signed(buffer_1_193) + $signed(buffer_7_200); // @[Modules.scala 166:64:@28239.4]
  assign _T_81304 = _T_81303[13:0]; // @[Modules.scala 166:64:@28240.4]
  assign buffer_8_406 = $signed(_T_81304); // @[Modules.scala 166:64:@28241.4]
  assign buffer_8_197 = {{9{_T_80234[4]}},_T_80234}; // @[Modules.scala 112:22:@8.4]
  assign _T_81306 = $signed(buffer_1_195) + $signed(buffer_8_197); // @[Modules.scala 166:64:@28243.4]
  assign _T_81307 = _T_81306[13:0]; // @[Modules.scala 166:64:@28244.4]
  assign buffer_8_407 = $signed(_T_81307); // @[Modules.scala 166:64:@28245.4]
  assign buffer_8_198 = {{8{_T_80241[5]}},_T_80241}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_199 = {{8{_T_80248[5]}},_T_80248}; // @[Modules.scala 112:22:@8.4]
  assign _T_81309 = $signed(buffer_8_198) + $signed(buffer_8_199); // @[Modules.scala 166:64:@28247.4]
  assign _T_81310 = _T_81309[13:0]; // @[Modules.scala 166:64:@28248.4]
  assign buffer_8_408 = $signed(_T_81310); // @[Modules.scala 166:64:@28249.4]
  assign _T_81312 = $signed(buffer_2_202) + $signed(buffer_4_192); // @[Modules.scala 166:64:@28251.4]
  assign _T_81313 = _T_81312[13:0]; // @[Modules.scala 166:64:@28252.4]
  assign buffer_8_409 = $signed(_T_81313); // @[Modules.scala 166:64:@28253.4]
  assign buffer_8_203 = {{9{_T_80276[4]}},_T_80276}; // @[Modules.scala 112:22:@8.4]
  assign _T_81315 = $signed(buffer_4_193) + $signed(buffer_8_203); // @[Modules.scala 166:64:@28255.4]
  assign _T_81316 = _T_81315[13:0]; // @[Modules.scala 166:64:@28256.4]
  assign buffer_8_410 = $signed(_T_81316); // @[Modules.scala 166:64:@28257.4]
  assign buffer_8_204 = {{9{_T_80283[4]}},_T_80283}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_205 = {{9{_T_80290[4]}},_T_80290}; // @[Modules.scala 112:22:@8.4]
  assign _T_81318 = $signed(buffer_8_204) + $signed(buffer_8_205); // @[Modules.scala 166:64:@28259.4]
  assign _T_81319 = _T_81318[13:0]; // @[Modules.scala 166:64:@28260.4]
  assign buffer_8_411 = $signed(_T_81319); // @[Modules.scala 166:64:@28261.4]
  assign buffer_8_207 = {{9{_T_80304[4]}},_T_80304}; // @[Modules.scala 112:22:@8.4]
  assign _T_81321 = $signed(buffer_7_211) + $signed(buffer_8_207); // @[Modules.scala 166:64:@28263.4]
  assign _T_81322 = _T_81321[13:0]; // @[Modules.scala 166:64:@28264.4]
  assign buffer_8_412 = $signed(_T_81322); // @[Modules.scala 166:64:@28265.4]
  assign buffer_8_208 = {{9{_T_80311[4]}},_T_80311}; // @[Modules.scala 112:22:@8.4]
  assign _T_81324 = $signed(buffer_8_208) + $signed(buffer_3_215); // @[Modules.scala 166:64:@28267.4]
  assign _T_81325 = _T_81324[13:0]; // @[Modules.scala 166:64:@28268.4]
  assign buffer_8_413 = $signed(_T_81325); // @[Modules.scala 166:64:@28269.4]
  assign buffer_8_210 = {{9{_T_80325[4]}},_T_80325}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_211 = {{8{_T_80332[5]}},_T_80332}; // @[Modules.scala 112:22:@8.4]
  assign _T_81327 = $signed(buffer_8_210) + $signed(buffer_8_211); // @[Modules.scala 166:64:@28271.4]
  assign _T_81328 = _T_81327[13:0]; // @[Modules.scala 166:64:@28272.4]
  assign buffer_8_414 = $signed(_T_81328); // @[Modules.scala 166:64:@28273.4]
  assign buffer_8_213 = {{8{_T_80346[5]}},_T_80346}; // @[Modules.scala 112:22:@8.4]
  assign _T_81330 = $signed(buffer_0_208) + $signed(buffer_8_213); // @[Modules.scala 166:64:@28275.4]
  assign _T_81331 = _T_81330[13:0]; // @[Modules.scala 166:64:@28276.4]
  assign buffer_8_415 = $signed(_T_81331); // @[Modules.scala 166:64:@28277.4]
  assign buffer_8_217 = {{9{_T_80374[4]}},_T_80374}; // @[Modules.scala 112:22:@8.4]
  assign _T_81336 = $signed(buffer_1_212) + $signed(buffer_8_217); // @[Modules.scala 166:64:@28283.4]
  assign _T_81337 = _T_81336[13:0]; // @[Modules.scala 166:64:@28284.4]
  assign buffer_8_417 = $signed(_T_81337); // @[Modules.scala 166:64:@28285.4]
  assign buffer_8_218 = {{9{_T_80381[4]}},_T_80381}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_219 = {{9{_T_80388[4]}},_T_80388}; // @[Modules.scala 112:22:@8.4]
  assign _T_81339 = $signed(buffer_8_218) + $signed(buffer_8_219); // @[Modules.scala 166:64:@28287.4]
  assign _T_81340 = _T_81339[13:0]; // @[Modules.scala 166:64:@28288.4]
  assign buffer_8_418 = $signed(_T_81340); // @[Modules.scala 166:64:@28289.4]
  assign buffer_8_222 = {{9{_T_80409[4]}},_T_80409}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_223 = {{8{_T_80416[5]}},_T_80416}; // @[Modules.scala 112:22:@8.4]
  assign _T_81345 = $signed(buffer_8_222) + $signed(buffer_8_223); // @[Modules.scala 166:64:@28295.4]
  assign _T_81346 = _T_81345[13:0]; // @[Modules.scala 166:64:@28296.4]
  assign buffer_8_420 = $signed(_T_81346); // @[Modules.scala 166:64:@28297.4]
  assign _T_81348 = $signed(buffer_1_219) + $signed(buffer_5_224); // @[Modules.scala 166:64:@28299.4]
  assign _T_81349 = _T_81348[13:0]; // @[Modules.scala 166:64:@28300.4]
  assign buffer_8_421 = $signed(_T_81349); // @[Modules.scala 166:64:@28301.4]
  assign buffer_8_226 = {{8{_T_80437[5]}},_T_80437}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_227 = {{8{_T_80444[5]}},_T_80444}; // @[Modules.scala 112:22:@8.4]
  assign _T_81351 = $signed(buffer_8_226) + $signed(buffer_8_227); // @[Modules.scala 166:64:@28303.4]
  assign _T_81352 = _T_81351[13:0]; // @[Modules.scala 166:64:@28304.4]
  assign buffer_8_422 = $signed(_T_81352); // @[Modules.scala 166:64:@28305.4]
  assign _T_81354 = $signed(buffer_3_233) + $signed(buffer_5_228); // @[Modules.scala 166:64:@28307.4]
  assign _T_81355 = _T_81354[13:0]; // @[Modules.scala 166:64:@28308.4]
  assign buffer_8_423 = $signed(_T_81355); // @[Modules.scala 166:64:@28309.4]
  assign buffer_8_231 = {{9{_T_80472[4]}},_T_80472}; // @[Modules.scala 112:22:@8.4]
  assign _T_81357 = $signed(buffer_5_229) + $signed(buffer_8_231); // @[Modules.scala 166:64:@28311.4]
  assign _T_81358 = _T_81357[13:0]; // @[Modules.scala 166:64:@28312.4]
  assign buffer_8_424 = $signed(_T_81358); // @[Modules.scala 166:64:@28313.4]
  assign _T_81360 = $signed(buffer_7_236) + $signed(buffer_2_231); // @[Modules.scala 166:64:@28315.4]
  assign _T_81361 = _T_81360[13:0]; // @[Modules.scala 166:64:@28316.4]
  assign buffer_8_425 = $signed(_T_81361); // @[Modules.scala 166:64:@28317.4]
  assign buffer_8_234 = {{9{_T_80493[4]}},_T_80493}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_235 = {{9{_T_80500[4]}},_T_80500}; // @[Modules.scala 112:22:@8.4]
  assign _T_81363 = $signed(buffer_8_234) + $signed(buffer_8_235); // @[Modules.scala 166:64:@28319.4]
  assign _T_81364 = _T_81363[13:0]; // @[Modules.scala 166:64:@28320.4]
  assign buffer_8_426 = $signed(_T_81364); // @[Modules.scala 166:64:@28321.4]
  assign buffer_8_236 = {{8{_T_80507[5]}},_T_80507}; // @[Modules.scala 112:22:@8.4]
  assign _T_81366 = $signed(buffer_8_236) + $signed(buffer_0_229); // @[Modules.scala 166:64:@28323.4]
  assign _T_81367 = _T_81366[13:0]; // @[Modules.scala 166:64:@28324.4]
  assign buffer_8_427 = $signed(_T_81367); // @[Modules.scala 166:64:@28325.4]
  assign buffer_8_239 = {{8{_T_80528[5]}},_T_80528}; // @[Modules.scala 112:22:@8.4]
  assign _T_81369 = $signed(buffer_5_238) + $signed(buffer_8_239); // @[Modules.scala 166:64:@28327.4]
  assign _T_81370 = _T_81369[13:0]; // @[Modules.scala 166:64:@28328.4]
  assign buffer_8_428 = $signed(_T_81370); // @[Modules.scala 166:64:@28329.4]
  assign _T_81372 = $signed(buffer_5_241) + $signed(buffer_5_242); // @[Modules.scala 166:64:@28331.4]
  assign _T_81373 = _T_81372[13:0]; // @[Modules.scala 166:64:@28332.4]
  assign buffer_8_429 = $signed(_T_81373); // @[Modules.scala 166:64:@28333.4]
  assign _T_81375 = $signed(buffer_5_243) + $signed(buffer_2_242); // @[Modules.scala 166:64:@28335.4]
  assign _T_81376 = _T_81375[13:0]; // @[Modules.scala 166:64:@28336.4]
  assign buffer_8_430 = $signed(_T_81376); // @[Modules.scala 166:64:@28337.4]
  assign _T_81381 = $signed(buffer_1_238) + $signed(buffer_4_233); // @[Modules.scala 166:64:@28343.4]
  assign _T_81382 = _T_81381[13:0]; // @[Modules.scala 166:64:@28344.4]
  assign buffer_8_432 = $signed(_T_81382); // @[Modules.scala 166:64:@28345.4]
  assign buffer_8_249 = {{8{_T_80598[5]}},_T_80598}; // @[Modules.scala 112:22:@8.4]
  assign _T_81384 = $signed(buffer_6_251) + $signed(buffer_8_249); // @[Modules.scala 166:64:@28347.4]
  assign _T_81385 = _T_81384[13:0]; // @[Modules.scala 166:64:@28348.4]
  assign buffer_8_433 = $signed(_T_81385); // @[Modules.scala 166:64:@28349.4]
  assign buffer_8_250 = {{8{_T_80605[5]}},_T_80605}; // @[Modules.scala 112:22:@8.4]
  assign _T_81387 = $signed(buffer_8_250) + $signed(buffer_2_251); // @[Modules.scala 166:64:@28351.4]
  assign _T_81388 = _T_81387[13:0]; // @[Modules.scala 166:64:@28352.4]
  assign buffer_8_434 = $signed(_T_81388); // @[Modules.scala 166:64:@28353.4]
  assign buffer_8_252 = {{8{_T_80619[5]}},_T_80619}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_253 = {{8{_T_80626[5]}},_T_80626}; // @[Modules.scala 112:22:@8.4]
  assign _T_81390 = $signed(buffer_8_252) + $signed(buffer_8_253); // @[Modules.scala 166:64:@28355.4]
  assign _T_81391 = _T_81390[13:0]; // @[Modules.scala 166:64:@28356.4]
  assign buffer_8_435 = $signed(_T_81391); // @[Modules.scala 166:64:@28357.4]
  assign _T_81393 = $signed(buffer_0_245) + $signed(buffer_4_242); // @[Modules.scala 166:64:@28359.4]
  assign _T_81394 = _T_81393[13:0]; // @[Modules.scala 166:64:@28360.4]
  assign buffer_8_436 = $signed(_T_81394); // @[Modules.scala 166:64:@28361.4]
  assign buffer_8_257 = {{9{_T_80654[4]}},_T_80654}; // @[Modules.scala 112:22:@8.4]
  assign _T_81396 = $signed(buffer_4_243) + $signed(buffer_8_257); // @[Modules.scala 166:64:@28363.4]
  assign _T_81397 = _T_81396[13:0]; // @[Modules.scala 166:64:@28364.4]
  assign buffer_8_437 = $signed(_T_81397); // @[Modules.scala 166:64:@28365.4]
  assign buffer_8_258 = {{8{_T_80661[5]}},_T_80661}; // @[Modules.scala 112:22:@8.4]
  assign _T_81399 = $signed(buffer_8_258) + $signed(buffer_2_259); // @[Modules.scala 166:64:@28367.4]
  assign _T_81400 = _T_81399[13:0]; // @[Modules.scala 166:64:@28368.4]
  assign buffer_8_438 = $signed(_T_81400); // @[Modules.scala 166:64:@28369.4]
  assign buffer_8_260 = {{8{_T_80675[5]}},_T_80675}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_261 = {{8{_T_80682[5]}},_T_80682}; // @[Modules.scala 112:22:@8.4]
  assign _T_81402 = $signed(buffer_8_260) + $signed(buffer_8_261); // @[Modules.scala 166:64:@28371.4]
  assign _T_81403 = _T_81402[13:0]; // @[Modules.scala 166:64:@28372.4]
  assign buffer_8_439 = $signed(_T_81403); // @[Modules.scala 166:64:@28373.4]
  assign _T_81405 = $signed(buffer_3_264) + $signed(buffer_4_252); // @[Modules.scala 166:64:@28375.4]
  assign _T_81406 = _T_81405[13:0]; // @[Modules.scala 166:64:@28376.4]
  assign buffer_8_440 = $signed(_T_81406); // @[Modules.scala 166:64:@28377.4]
  assign buffer_8_265 = {{8{_T_80710[5]}},_T_80710}; // @[Modules.scala 112:22:@8.4]
  assign _T_81408 = $signed(buffer_4_253) + $signed(buffer_8_265); // @[Modules.scala 166:64:@28379.4]
  assign _T_81409 = _T_81408[13:0]; // @[Modules.scala 166:64:@28380.4]
  assign buffer_8_441 = $signed(_T_81409); // @[Modules.scala 166:64:@28381.4]
  assign buffer_8_266 = {{8{_T_80717[5]}},_T_80717}; // @[Modules.scala 112:22:@8.4]
  assign _T_81411 = $signed(buffer_8_266) + $signed(buffer_3_269); // @[Modules.scala 166:64:@28383.4]
  assign _T_81412 = _T_81411[13:0]; // @[Modules.scala 166:64:@28384.4]
  assign buffer_8_442 = $signed(_T_81412); // @[Modules.scala 166:64:@28385.4]
  assign _T_81414 = $signed(buffer_7_269) + $signed(buffer_0_263); // @[Modules.scala 166:64:@28387.4]
  assign _T_81415 = _T_81414[13:0]; // @[Modules.scala 166:64:@28388.4]
  assign buffer_8_443 = $signed(_T_81415); // @[Modules.scala 166:64:@28389.4]
  assign _T_81417 = $signed(buffer_1_263) + $signed(buffer_1_264); // @[Modules.scala 166:64:@28391.4]
  assign _T_81418 = _T_81417[13:0]; // @[Modules.scala 166:64:@28392.4]
  assign buffer_8_444 = $signed(_T_81418); // @[Modules.scala 166:64:@28393.4]
  assign _T_81426 = $signed(buffer_4_265) + $signed(buffer_0_272); // @[Modules.scala 166:64:@28403.4]
  assign _T_81427 = _T_81426[13:0]; // @[Modules.scala 166:64:@28404.4]
  assign buffer_8_447 = $signed(_T_81427); // @[Modules.scala 166:64:@28405.4]
  assign buffer_8_278 = {{8{_T_80801[5]}},_T_80801}; // @[Modules.scala 112:22:@8.4]
  assign _T_81429 = $signed(buffer_8_278) + $signed(buffer_3_283); // @[Modules.scala 166:64:@28407.4]
  assign _T_81430 = _T_81429[13:0]; // @[Modules.scala 166:64:@28408.4]
  assign buffer_8_448 = $signed(_T_81430); // @[Modules.scala 166:64:@28409.4]
  assign _T_81444 = $signed(buffer_3_291) + $signed(buffer_7_289); // @[Modules.scala 166:64:@28427.4]
  assign _T_81445 = _T_81444[13:0]; // @[Modules.scala 166:64:@28428.4]
  assign buffer_8_453 = $signed(_T_81445); // @[Modules.scala 166:64:@28429.4]
  assign buffer_8_290 = {{8{_T_80885[5]}},_T_80885}; // @[Modules.scala 112:22:@8.4]
  assign buffer_8_291 = {{8{_T_80892[5]}},_T_80892}; // @[Modules.scala 112:22:@8.4]
  assign _T_81447 = $signed(buffer_8_290) + $signed(buffer_8_291); // @[Modules.scala 166:64:@28431.4]
  assign _T_81448 = _T_81447[13:0]; // @[Modules.scala 166:64:@28432.4]
  assign buffer_8_454 = $signed(_T_81448); // @[Modules.scala 166:64:@28433.4]
  assign _T_81453 = $signed(buffer_1_289) + $signed(buffer_1_290); // @[Modules.scala 166:64:@28439.4]
  assign _T_81454 = _T_81453[13:0]; // @[Modules.scala 166:64:@28440.4]
  assign buffer_8_456 = $signed(_T_81454); // @[Modules.scala 166:64:@28441.4]
  assign _T_81456 = $signed(buffer_1_291) + $signed(buffer_5_302); // @[Modules.scala 166:64:@28443.4]
  assign _T_81457 = _T_81456[13:0]; // @[Modules.scala 166:64:@28444.4]
  assign buffer_8_457 = $signed(_T_81457); // @[Modules.scala 166:64:@28445.4]
  assign buffer_8_299 = {{8{_T_80948[5]}},_T_80948}; // @[Modules.scala 112:22:@8.4]
  assign _T_81459 = $signed(buffer_7_299) + $signed(buffer_8_299); // @[Modules.scala 166:64:@28447.4]
  assign _T_81460 = _T_81459[13:0]; // @[Modules.scala 166:64:@28448.4]
  assign buffer_8_458 = $signed(_T_81460); // @[Modules.scala 166:64:@28449.4]
  assign buffer_8_300 = {{8{_T_80955[5]}},_T_80955}; // @[Modules.scala 112:22:@8.4]
  assign _T_81462 = $signed(buffer_8_300) + $signed(buffer_0_294); // @[Modules.scala 166:64:@28451.4]
  assign _T_81463 = _T_81462[13:0]; // @[Modules.scala 166:64:@28452.4]
  assign buffer_8_459 = $signed(_T_81463); // @[Modules.scala 166:64:@28453.4]
  assign buffer_8_304 = {{8{_T_80983[5]}},_T_80983}; // @[Modules.scala 112:22:@8.4]
  assign _T_81468 = $signed(buffer_8_304) + $signed(buffer_0_298); // @[Modules.scala 166:64:@28459.4]
  assign _T_81469 = _T_81468[13:0]; // @[Modules.scala 166:64:@28460.4]
  assign buffer_8_461 = $signed(_T_81469); // @[Modules.scala 166:64:@28461.4]
  assign buffer_8_306 = {{8{_T_80997[5]}},_T_80997}; // @[Modules.scala 112:22:@8.4]
  assign _T_81471 = $signed(buffer_8_306) + $signed(buffer_2_309); // @[Modules.scala 166:64:@28463.4]
  assign _T_81472 = _T_81471[13:0]; // @[Modules.scala 166:64:@28464.4]
  assign buffer_8_462 = $signed(_T_81472); // @[Modules.scala 166:64:@28465.4]
  assign _T_81474 = $signed(buffer_2_310) + $signed(buffer_8_310); // @[Modules.scala 160:64:@28467.4]
  assign _T_81475 = _T_81474[13:0]; // @[Modules.scala 160:64:@28468.4]
  assign buffer_8_463 = $signed(_T_81475); // @[Modules.scala 160:64:@28469.4]
  assign _T_81477 = $signed(buffer_8_311) + $signed(buffer_8_312); // @[Modules.scala 160:64:@28471.4]
  assign _T_81478 = _T_81477[13:0]; // @[Modules.scala 160:64:@28472.4]
  assign buffer_8_464 = $signed(_T_81478); // @[Modules.scala 160:64:@28473.4]
  assign _T_81480 = $signed(buffer_8_313) + $signed(buffer_8_314); // @[Modules.scala 160:64:@28475.4]
  assign _T_81481 = _T_81480[13:0]; // @[Modules.scala 160:64:@28476.4]
  assign buffer_8_465 = $signed(_T_81481); // @[Modules.scala 160:64:@28477.4]
  assign _T_81483 = $signed(buffer_8_315) + $signed(buffer_8_316); // @[Modules.scala 160:64:@28479.4]
  assign _T_81484 = _T_81483[13:0]; // @[Modules.scala 160:64:@28480.4]
  assign buffer_8_466 = $signed(_T_81484); // @[Modules.scala 160:64:@28481.4]
  assign _T_81486 = $signed(buffer_7_316) + $signed(buffer_7_317); // @[Modules.scala 160:64:@28483.4]
  assign _T_81487 = _T_81486[13:0]; // @[Modules.scala 160:64:@28484.4]
  assign buffer_8_467 = $signed(_T_81487); // @[Modules.scala 160:64:@28485.4]
  assign _T_81489 = $signed(buffer_7_318) + $signed(buffer_8_320); // @[Modules.scala 160:64:@28487.4]
  assign _T_81490 = _T_81489[13:0]; // @[Modules.scala 160:64:@28488.4]
  assign buffer_8_468 = $signed(_T_81490); // @[Modules.scala 160:64:@28489.4]
  assign _T_81492 = $signed(buffer_8_321) + $signed(buffer_1_316); // @[Modules.scala 160:64:@28491.4]
  assign _T_81493 = _T_81492[13:0]; // @[Modules.scala 160:64:@28492.4]
  assign buffer_8_469 = $signed(_T_81493); // @[Modules.scala 160:64:@28493.4]
  assign _T_81495 = $signed(buffer_1_317) + $signed(buffer_7_323); // @[Modules.scala 160:64:@28495.4]
  assign _T_81496 = _T_81495[13:0]; // @[Modules.scala 160:64:@28496.4]
  assign buffer_8_470 = $signed(_T_81496); // @[Modules.scala 160:64:@28497.4]
  assign _T_81498 = $signed(buffer_7_324) + $signed(buffer_8_326); // @[Modules.scala 160:64:@28499.4]
  assign _T_81499 = _T_81498[13:0]; // @[Modules.scala 160:64:@28500.4]
  assign buffer_8_471 = $signed(_T_81499); // @[Modules.scala 160:64:@28501.4]
  assign _T_81501 = $signed(buffer_8_327) + $signed(buffer_8_328); // @[Modules.scala 160:64:@28503.4]
  assign _T_81502 = _T_81501[13:0]; // @[Modules.scala 160:64:@28504.4]
  assign buffer_8_472 = $signed(_T_81502); // @[Modules.scala 160:64:@28505.4]
  assign _T_81504 = $signed(buffer_8_329) + $signed(buffer_8_330); // @[Modules.scala 160:64:@28507.4]
  assign _T_81505 = _T_81504[13:0]; // @[Modules.scala 160:64:@28508.4]
  assign buffer_8_473 = $signed(_T_81505); // @[Modules.scala 160:64:@28509.4]
  assign _T_81507 = $signed(buffer_6_338) + $signed(buffer_8_332); // @[Modules.scala 160:64:@28511.4]
  assign _T_81508 = _T_81507[13:0]; // @[Modules.scala 160:64:@28512.4]
  assign buffer_8_474 = $signed(_T_81508); // @[Modules.scala 160:64:@28513.4]
  assign _T_81510 = $signed(buffer_8_333) + $signed(buffer_8_334); // @[Modules.scala 160:64:@28515.4]
  assign _T_81511 = _T_81510[13:0]; // @[Modules.scala 160:64:@28516.4]
  assign buffer_8_475 = $signed(_T_81511); // @[Modules.scala 160:64:@28517.4]
  assign _T_81513 = $signed(buffer_8_335) + $signed(buffer_8_336); // @[Modules.scala 160:64:@28519.4]
  assign _T_81514 = _T_81513[13:0]; // @[Modules.scala 160:64:@28520.4]
  assign buffer_8_476 = $signed(_T_81514); // @[Modules.scala 160:64:@28521.4]
  assign _T_81516 = $signed(buffer_8_337) + $signed(buffer_8_338); // @[Modules.scala 160:64:@28523.4]
  assign _T_81517 = _T_81516[13:0]; // @[Modules.scala 160:64:@28524.4]
  assign buffer_8_477 = $signed(_T_81517); // @[Modules.scala 160:64:@28525.4]
  assign _T_81519 = $signed(buffer_8_339) + $signed(buffer_8_340); // @[Modules.scala 160:64:@28527.4]
  assign _T_81520 = _T_81519[13:0]; // @[Modules.scala 160:64:@28528.4]
  assign buffer_8_478 = $signed(_T_81520); // @[Modules.scala 160:64:@28529.4]
  assign _T_81522 = $signed(buffer_8_341) + $signed(buffer_8_342); // @[Modules.scala 160:64:@28531.4]
  assign _T_81523 = _T_81522[13:0]; // @[Modules.scala 160:64:@28532.4]
  assign buffer_8_479 = $signed(_T_81523); // @[Modules.scala 160:64:@28533.4]
  assign _T_81525 = $signed(buffer_8_343) + $signed(buffer_8_344); // @[Modules.scala 160:64:@28535.4]
  assign _T_81526 = _T_81525[13:0]; // @[Modules.scala 160:64:@28536.4]
  assign buffer_8_480 = $signed(_T_81526); // @[Modules.scala 160:64:@28537.4]
  assign _T_81528 = $signed(buffer_5_353) + $signed(buffer_8_346); // @[Modules.scala 160:64:@28539.4]
  assign _T_81529 = _T_81528[13:0]; // @[Modules.scala 160:64:@28540.4]
  assign buffer_8_481 = $signed(_T_81529); // @[Modules.scala 160:64:@28541.4]
  assign _T_81531 = $signed(buffer_8_347) + $signed(buffer_8_348); // @[Modules.scala 160:64:@28543.4]
  assign _T_81532 = _T_81531[13:0]; // @[Modules.scala 160:64:@28544.4]
  assign buffer_8_482 = $signed(_T_81532); // @[Modules.scala 160:64:@28545.4]
  assign _T_81534 = $signed(buffer_8_349) + $signed(buffer_8_350); // @[Modules.scala 160:64:@28547.4]
  assign _T_81535 = _T_81534[13:0]; // @[Modules.scala 160:64:@28548.4]
  assign buffer_8_483 = $signed(_T_81535); // @[Modules.scala 160:64:@28549.4]
  assign _T_81537 = $signed(buffer_8_351) + $signed(buffer_8_352); // @[Modules.scala 160:64:@28551.4]
  assign _T_81538 = _T_81537[13:0]; // @[Modules.scala 160:64:@28552.4]
  assign buffer_8_484 = $signed(_T_81538); // @[Modules.scala 160:64:@28553.4]
  assign _T_81540 = $signed(buffer_8_353) + $signed(buffer_3_362); // @[Modules.scala 160:64:@28555.4]
  assign _T_81541 = _T_81540[13:0]; // @[Modules.scala 160:64:@28556.4]
  assign buffer_8_485 = $signed(_T_81541); // @[Modules.scala 160:64:@28557.4]
  assign _T_81543 = $signed(buffer_8_355) + $signed(buffer_8_356); // @[Modules.scala 160:64:@28559.4]
  assign _T_81544 = _T_81543[13:0]; // @[Modules.scala 160:64:@28560.4]
  assign buffer_8_486 = $signed(_T_81544); // @[Modules.scala 160:64:@28561.4]
  assign _T_81546 = $signed(buffer_5_366) + $signed(buffer_8_358); // @[Modules.scala 160:64:@28563.4]
  assign _T_81547 = _T_81546[13:0]; // @[Modules.scala 160:64:@28564.4]
  assign buffer_8_487 = $signed(_T_81547); // @[Modules.scala 160:64:@28565.4]
  assign _T_81549 = $signed(buffer_8_359) + $signed(buffer_8_360); // @[Modules.scala 160:64:@28567.4]
  assign _T_81550 = _T_81549[13:0]; // @[Modules.scala 160:64:@28568.4]
  assign buffer_8_488 = $signed(_T_81550); // @[Modules.scala 160:64:@28569.4]
  assign _T_81552 = $signed(buffer_8_361) + $signed(buffer_8_362); // @[Modules.scala 160:64:@28571.4]
  assign _T_81553 = _T_81552[13:0]; // @[Modules.scala 160:64:@28572.4]
  assign buffer_8_489 = $signed(_T_81553); // @[Modules.scala 160:64:@28573.4]
  assign _T_81555 = $signed(buffer_8_363) + $signed(buffer_8_364); // @[Modules.scala 160:64:@28575.4]
  assign _T_81556 = _T_81555[13:0]; // @[Modules.scala 160:64:@28576.4]
  assign buffer_8_490 = $signed(_T_81556); // @[Modules.scala 160:64:@28577.4]
  assign _T_81558 = $signed(buffer_8_365) + $signed(buffer_8_366); // @[Modules.scala 160:64:@28579.4]
  assign _T_81559 = _T_81558[13:0]; // @[Modules.scala 160:64:@28580.4]
  assign buffer_8_491 = $signed(_T_81559); // @[Modules.scala 160:64:@28581.4]
  assign _T_81561 = $signed(buffer_8_367) + $signed(buffer_8_368); // @[Modules.scala 160:64:@28583.4]
  assign _T_81562 = _T_81561[13:0]; // @[Modules.scala 160:64:@28584.4]
  assign buffer_8_492 = $signed(_T_81562); // @[Modules.scala 160:64:@28585.4]
  assign _T_81564 = $signed(buffer_0_363) + $signed(buffer_8_370); // @[Modules.scala 160:64:@28587.4]
  assign _T_81565 = _T_81564[13:0]; // @[Modules.scala 160:64:@28588.4]
  assign buffer_8_493 = $signed(_T_81565); // @[Modules.scala 160:64:@28589.4]
  assign _T_81567 = $signed(buffer_8_371) + $signed(buffer_8_372); // @[Modules.scala 160:64:@28591.4]
  assign _T_81568 = _T_81567[13:0]; // @[Modules.scala 160:64:@28592.4]
  assign buffer_8_494 = $signed(_T_81568); // @[Modules.scala 160:64:@28593.4]
  assign _T_81570 = $signed(buffer_2_376) + $signed(buffer_8_374); // @[Modules.scala 160:64:@28595.4]
  assign _T_81571 = _T_81570[13:0]; // @[Modules.scala 160:64:@28596.4]
  assign buffer_8_495 = $signed(_T_81571); // @[Modules.scala 160:64:@28597.4]
  assign _T_81573 = $signed(buffer_8_375) + $signed(buffer_7_376); // @[Modules.scala 160:64:@28599.4]
  assign _T_81574 = _T_81573[13:0]; // @[Modules.scala 160:64:@28600.4]
  assign buffer_8_496 = $signed(_T_81574); // @[Modules.scala 160:64:@28601.4]
  assign _T_81576 = $signed(buffer_7_377) + $signed(buffer_8_378); // @[Modules.scala 160:64:@28603.4]
  assign _T_81577 = _T_81576[13:0]; // @[Modules.scala 160:64:@28604.4]
  assign buffer_8_497 = $signed(_T_81577); // @[Modules.scala 160:64:@28605.4]
  assign _T_81579 = $signed(buffer_8_379) + $signed(buffer_8_380); // @[Modules.scala 160:64:@28607.4]
  assign _T_81580 = _T_81579[13:0]; // @[Modules.scala 160:64:@28608.4]
  assign buffer_8_498 = $signed(_T_81580); // @[Modules.scala 160:64:@28609.4]
  assign _T_81582 = $signed(buffer_8_381) + $signed(buffer_8_382); // @[Modules.scala 160:64:@28611.4]
  assign _T_81583 = _T_81582[13:0]; // @[Modules.scala 160:64:@28612.4]
  assign buffer_8_499 = $signed(_T_81583); // @[Modules.scala 160:64:@28613.4]
  assign _T_81585 = $signed(buffer_8_383) + $signed(buffer_8_384); // @[Modules.scala 160:64:@28615.4]
  assign _T_81586 = _T_81585[13:0]; // @[Modules.scala 160:64:@28616.4]
  assign buffer_8_500 = $signed(_T_81586); // @[Modules.scala 160:64:@28617.4]
  assign _T_81588 = $signed(buffer_8_385) + $signed(buffer_8_386); // @[Modules.scala 160:64:@28619.4]
  assign _T_81589 = _T_81588[13:0]; // @[Modules.scala 160:64:@28620.4]
  assign buffer_8_501 = $signed(_T_81589); // @[Modules.scala 160:64:@28621.4]
  assign _T_81591 = $signed(buffer_8_387) + $signed(buffer_8_388); // @[Modules.scala 160:64:@28623.4]
  assign _T_81592 = _T_81591[13:0]; // @[Modules.scala 160:64:@28624.4]
  assign buffer_8_502 = $signed(_T_81592); // @[Modules.scala 160:64:@28625.4]
  assign _T_81594 = $signed(buffer_8_389) + $signed(buffer_7_392); // @[Modules.scala 160:64:@28627.4]
  assign _T_81595 = _T_81594[13:0]; // @[Modules.scala 160:64:@28628.4]
  assign buffer_8_503 = $signed(_T_81595); // @[Modules.scala 160:64:@28629.4]
  assign _T_81597 = $signed(buffer_8_391) + $signed(buffer_8_392); // @[Modules.scala 160:64:@28631.4]
  assign _T_81598 = _T_81597[13:0]; // @[Modules.scala 160:64:@28632.4]
  assign buffer_8_504 = $signed(_T_81598); // @[Modules.scala 160:64:@28633.4]
  assign _T_81600 = $signed(buffer_8_393) + $signed(buffer_8_394); // @[Modules.scala 160:64:@28635.4]
  assign _T_81601 = _T_81600[13:0]; // @[Modules.scala 160:64:@28636.4]
  assign buffer_8_505 = $signed(_T_81601); // @[Modules.scala 160:64:@28637.4]
  assign _T_81603 = $signed(buffer_8_395) + $signed(buffer_8_396); // @[Modules.scala 160:64:@28639.4]
  assign _T_81604 = _T_81603[13:0]; // @[Modules.scala 160:64:@28640.4]
  assign buffer_8_506 = $signed(_T_81604); // @[Modules.scala 160:64:@28641.4]
  assign _T_81606 = $signed(buffer_8_397) + $signed(buffer_6_408); // @[Modules.scala 160:64:@28643.4]
  assign _T_81607 = _T_81606[13:0]; // @[Modules.scala 160:64:@28644.4]
  assign buffer_8_507 = $signed(_T_81607); // @[Modules.scala 160:64:@28645.4]
  assign _T_81609 = $signed(buffer_8_399) + $signed(buffer_3_409); // @[Modules.scala 160:64:@28647.4]
  assign _T_81610 = _T_81609[13:0]; // @[Modules.scala 160:64:@28648.4]
  assign buffer_8_508 = $signed(_T_81610); // @[Modules.scala 160:64:@28649.4]
  assign _T_81612 = $signed(buffer_3_410) + $signed(buffer_8_402); // @[Modules.scala 160:64:@28651.4]
  assign _T_81613 = _T_81612[13:0]; // @[Modules.scala 160:64:@28652.4]
  assign buffer_8_509 = $signed(_T_81613); // @[Modules.scala 160:64:@28653.4]
  assign _T_81615 = $signed(buffer_8_403) + $signed(buffer_8_404); // @[Modules.scala 160:64:@28655.4]
  assign _T_81616 = _T_81615[13:0]; // @[Modules.scala 160:64:@28656.4]
  assign buffer_8_510 = $signed(_T_81616); // @[Modules.scala 160:64:@28657.4]
  assign _T_81618 = $signed(buffer_8_405) + $signed(buffer_8_406); // @[Modules.scala 160:64:@28659.4]
  assign _T_81619 = _T_81618[13:0]; // @[Modules.scala 160:64:@28660.4]
  assign buffer_8_511 = $signed(_T_81619); // @[Modules.scala 160:64:@28661.4]
  assign _T_81621 = $signed(buffer_8_407) + $signed(buffer_8_408); // @[Modules.scala 160:64:@28663.4]
  assign _T_81622 = _T_81621[13:0]; // @[Modules.scala 160:64:@28664.4]
  assign buffer_8_512 = $signed(_T_81622); // @[Modules.scala 160:64:@28665.4]
  assign _T_81624 = $signed(buffer_8_409) + $signed(buffer_8_410); // @[Modules.scala 160:64:@28667.4]
  assign _T_81625 = _T_81624[13:0]; // @[Modules.scala 160:64:@28668.4]
  assign buffer_8_513 = $signed(_T_81625); // @[Modules.scala 160:64:@28669.4]
  assign _T_81627 = $signed(buffer_8_411) + $signed(buffer_8_412); // @[Modules.scala 160:64:@28671.4]
  assign _T_81628 = _T_81627[13:0]; // @[Modules.scala 160:64:@28672.4]
  assign buffer_8_514 = $signed(_T_81628); // @[Modules.scala 160:64:@28673.4]
  assign _T_81630 = $signed(buffer_8_413) + $signed(buffer_8_414); // @[Modules.scala 160:64:@28675.4]
  assign _T_81631 = _T_81630[13:0]; // @[Modules.scala 160:64:@28676.4]
  assign buffer_8_515 = $signed(_T_81631); // @[Modules.scala 160:64:@28677.4]
  assign _T_81633 = $signed(buffer_8_415) + $signed(buffer_1_409); // @[Modules.scala 160:64:@28679.4]
  assign _T_81634 = _T_81633[13:0]; // @[Modules.scala 160:64:@28680.4]
  assign buffer_8_516 = $signed(_T_81634); // @[Modules.scala 160:64:@28681.4]
  assign _T_81636 = $signed(buffer_8_417) + $signed(buffer_8_418); // @[Modules.scala 160:64:@28683.4]
  assign _T_81637 = _T_81636[13:0]; // @[Modules.scala 160:64:@28684.4]
  assign buffer_8_517 = $signed(_T_81637); // @[Modules.scala 160:64:@28685.4]
  assign _T_81639 = $signed(buffer_4_404) + $signed(buffer_8_420); // @[Modules.scala 160:64:@28687.4]
  assign _T_81640 = _T_81639[13:0]; // @[Modules.scala 160:64:@28688.4]
  assign buffer_8_518 = $signed(_T_81640); // @[Modules.scala 160:64:@28689.4]
  assign _T_81642 = $signed(buffer_8_421) + $signed(buffer_8_422); // @[Modules.scala 160:64:@28691.4]
  assign _T_81643 = _T_81642[13:0]; // @[Modules.scala 160:64:@28692.4]
  assign buffer_8_519 = $signed(_T_81643); // @[Modules.scala 160:64:@28693.4]
  assign _T_81645 = $signed(buffer_8_423) + $signed(buffer_8_424); // @[Modules.scala 160:64:@28695.4]
  assign _T_81646 = _T_81645[13:0]; // @[Modules.scala 160:64:@28696.4]
  assign buffer_8_520 = $signed(_T_81646); // @[Modules.scala 160:64:@28697.4]
  assign _T_81648 = $signed(buffer_8_425) + $signed(buffer_8_426); // @[Modules.scala 160:64:@28699.4]
  assign _T_81649 = _T_81648[13:0]; // @[Modules.scala 160:64:@28700.4]
  assign buffer_8_521 = $signed(_T_81649); // @[Modules.scala 160:64:@28701.4]
  assign _T_81651 = $signed(buffer_8_427) + $signed(buffer_8_428); // @[Modules.scala 160:64:@28703.4]
  assign _T_81652 = _T_81651[13:0]; // @[Modules.scala 160:64:@28704.4]
  assign buffer_8_522 = $signed(_T_81652); // @[Modules.scala 160:64:@28705.4]
  assign _T_81654 = $signed(buffer_8_429) + $signed(buffer_8_430); // @[Modules.scala 160:64:@28707.4]
  assign _T_81655 = _T_81654[13:0]; // @[Modules.scala 160:64:@28708.4]
  assign buffer_8_523 = $signed(_T_81655); // @[Modules.scala 160:64:@28709.4]
  assign _T_81657 = $signed(buffer_1_422) + $signed(buffer_8_432); // @[Modules.scala 160:64:@28711.4]
  assign _T_81658 = _T_81657[13:0]; // @[Modules.scala 160:64:@28712.4]
  assign buffer_8_524 = $signed(_T_81658); // @[Modules.scala 160:64:@28713.4]
  assign _T_81660 = $signed(buffer_8_433) + $signed(buffer_8_434); // @[Modules.scala 160:64:@28715.4]
  assign _T_81661 = _T_81660[13:0]; // @[Modules.scala 160:64:@28716.4]
  assign buffer_8_525 = $signed(_T_81661); // @[Modules.scala 160:64:@28717.4]
  assign _T_81663 = $signed(buffer_8_435) + $signed(buffer_8_436); // @[Modules.scala 160:64:@28719.4]
  assign _T_81664 = _T_81663[13:0]; // @[Modules.scala 160:64:@28720.4]
  assign buffer_8_526 = $signed(_T_81664); // @[Modules.scala 160:64:@28721.4]
  assign _T_81666 = $signed(buffer_8_437) + $signed(buffer_8_438); // @[Modules.scala 160:64:@28723.4]
  assign _T_81667 = _T_81666[13:0]; // @[Modules.scala 160:64:@28724.4]
  assign buffer_8_527 = $signed(_T_81667); // @[Modules.scala 160:64:@28725.4]
  assign _T_81669 = $signed(buffer_8_439) + $signed(buffer_8_440); // @[Modules.scala 160:64:@28727.4]
  assign _T_81670 = _T_81669[13:0]; // @[Modules.scala 160:64:@28728.4]
  assign buffer_8_528 = $signed(_T_81670); // @[Modules.scala 160:64:@28729.4]
  assign _T_81672 = $signed(buffer_8_441) + $signed(buffer_8_442); // @[Modules.scala 160:64:@28731.4]
  assign _T_81673 = _T_81672[13:0]; // @[Modules.scala 160:64:@28732.4]
  assign buffer_8_529 = $signed(_T_81673); // @[Modules.scala 160:64:@28733.4]
  assign _T_81675 = $signed(buffer_8_443) + $signed(buffer_8_444); // @[Modules.scala 160:64:@28735.4]
  assign _T_81676 = _T_81675[13:0]; // @[Modules.scala 160:64:@28736.4]
  assign buffer_8_530 = $signed(_T_81676); // @[Modules.scala 160:64:@28737.4]
  assign _T_81681 = $signed(buffer_8_447) + $signed(buffer_8_448); // @[Modules.scala 160:64:@28743.4]
  assign _T_81682 = _T_81681[13:0]; // @[Modules.scala 160:64:@28744.4]
  assign buffer_8_532 = $signed(_T_81682); // @[Modules.scala 160:64:@28745.4]
  assign _T_81684 = $signed(buffer_1_441) + $signed(buffer_1_442); // @[Modules.scala 160:64:@28747.4]
  assign _T_81685 = _T_81684[13:0]; // @[Modules.scala 160:64:@28748.4]
  assign buffer_8_533 = $signed(_T_81685); // @[Modules.scala 160:64:@28749.4]
  assign _T_81687 = $signed(buffer_1_443) + $signed(buffer_1_444); // @[Modules.scala 160:64:@28751.4]
  assign _T_81688 = _T_81687[13:0]; // @[Modules.scala 160:64:@28752.4]
  assign buffer_8_534 = $signed(_T_81688); // @[Modules.scala 160:64:@28753.4]
  assign _T_81690 = $signed(buffer_8_453) + $signed(buffer_8_454); // @[Modules.scala 160:64:@28755.4]
  assign _T_81691 = _T_81690[13:0]; // @[Modules.scala 160:64:@28756.4]
  assign buffer_8_535 = $signed(_T_81691); // @[Modules.scala 160:64:@28757.4]
  assign _T_81693 = $signed(buffer_7_456) + $signed(buffer_8_456); // @[Modules.scala 160:64:@28759.4]
  assign _T_81694 = _T_81693[13:0]; // @[Modules.scala 160:64:@28760.4]
  assign buffer_8_536 = $signed(_T_81694); // @[Modules.scala 160:64:@28761.4]
  assign _T_81696 = $signed(buffer_8_457) + $signed(buffer_8_458); // @[Modules.scala 160:64:@28763.4]
  assign _T_81697 = _T_81696[13:0]; // @[Modules.scala 160:64:@28764.4]
  assign buffer_8_537 = $signed(_T_81697); // @[Modules.scala 160:64:@28765.4]
  assign _T_81699 = $signed(buffer_8_459) + $signed(buffer_2_462); // @[Modules.scala 160:64:@28767.4]
  assign _T_81700 = _T_81699[13:0]; // @[Modules.scala 160:64:@28768.4]
  assign buffer_8_538 = $signed(_T_81700); // @[Modules.scala 160:64:@28769.4]
  assign _T_81702 = $signed(buffer_8_461) + $signed(buffer_8_462); // @[Modules.scala 160:64:@28771.4]
  assign _T_81703 = _T_81702[13:0]; // @[Modules.scala 160:64:@28772.4]
  assign buffer_8_539 = $signed(_T_81703); // @[Modules.scala 160:64:@28773.4]
  assign _T_81705 = $signed(buffer_8_463) + $signed(buffer_8_464); // @[Modules.scala 166:64:@28775.4]
  assign _T_81706 = _T_81705[13:0]; // @[Modules.scala 166:64:@28776.4]
  assign buffer_8_540 = $signed(_T_81706); // @[Modules.scala 166:64:@28777.4]
  assign _T_81708 = $signed(buffer_8_465) + $signed(buffer_8_466); // @[Modules.scala 166:64:@28779.4]
  assign _T_81709 = _T_81708[13:0]; // @[Modules.scala 166:64:@28780.4]
  assign buffer_8_541 = $signed(_T_81709); // @[Modules.scala 166:64:@28781.4]
  assign _T_81711 = $signed(buffer_8_467) + $signed(buffer_8_468); // @[Modules.scala 166:64:@28783.4]
  assign _T_81712 = _T_81711[13:0]; // @[Modules.scala 166:64:@28784.4]
  assign buffer_8_542 = $signed(_T_81712); // @[Modules.scala 166:64:@28785.4]
  assign _T_81714 = $signed(buffer_8_469) + $signed(buffer_8_470); // @[Modules.scala 166:64:@28787.4]
  assign _T_81715 = _T_81714[13:0]; // @[Modules.scala 166:64:@28788.4]
  assign buffer_8_543 = $signed(_T_81715); // @[Modules.scala 166:64:@28789.4]
  assign _T_81717 = $signed(buffer_8_471) + $signed(buffer_8_472); // @[Modules.scala 166:64:@28791.4]
  assign _T_81718 = _T_81717[13:0]; // @[Modules.scala 166:64:@28792.4]
  assign buffer_8_544 = $signed(_T_81718); // @[Modules.scala 166:64:@28793.4]
  assign _T_81720 = $signed(buffer_8_473) + $signed(buffer_8_474); // @[Modules.scala 166:64:@28795.4]
  assign _T_81721 = _T_81720[13:0]; // @[Modules.scala 166:64:@28796.4]
  assign buffer_8_545 = $signed(_T_81721); // @[Modules.scala 166:64:@28797.4]
  assign _T_81723 = $signed(buffer_8_475) + $signed(buffer_8_476); // @[Modules.scala 166:64:@28799.4]
  assign _T_81724 = _T_81723[13:0]; // @[Modules.scala 166:64:@28800.4]
  assign buffer_8_546 = $signed(_T_81724); // @[Modules.scala 166:64:@28801.4]
  assign _T_81726 = $signed(buffer_8_477) + $signed(buffer_8_478); // @[Modules.scala 166:64:@28803.4]
  assign _T_81727 = _T_81726[13:0]; // @[Modules.scala 166:64:@28804.4]
  assign buffer_8_547 = $signed(_T_81727); // @[Modules.scala 166:64:@28805.4]
  assign _T_81729 = $signed(buffer_8_479) + $signed(buffer_8_480); // @[Modules.scala 166:64:@28807.4]
  assign _T_81730 = _T_81729[13:0]; // @[Modules.scala 166:64:@28808.4]
  assign buffer_8_548 = $signed(_T_81730); // @[Modules.scala 166:64:@28809.4]
  assign _T_81732 = $signed(buffer_8_481) + $signed(buffer_8_482); // @[Modules.scala 166:64:@28811.4]
  assign _T_81733 = _T_81732[13:0]; // @[Modules.scala 166:64:@28812.4]
  assign buffer_8_549 = $signed(_T_81733); // @[Modules.scala 166:64:@28813.4]
  assign _T_81735 = $signed(buffer_8_483) + $signed(buffer_8_484); // @[Modules.scala 166:64:@28815.4]
  assign _T_81736 = _T_81735[13:0]; // @[Modules.scala 166:64:@28816.4]
  assign buffer_8_550 = $signed(_T_81736); // @[Modules.scala 166:64:@28817.4]
  assign _T_81738 = $signed(buffer_8_485) + $signed(buffer_8_486); // @[Modules.scala 166:64:@28819.4]
  assign _T_81739 = _T_81738[13:0]; // @[Modules.scala 166:64:@28820.4]
  assign buffer_8_551 = $signed(_T_81739); // @[Modules.scala 166:64:@28821.4]
  assign _T_81741 = $signed(buffer_8_487) + $signed(buffer_8_488); // @[Modules.scala 166:64:@28823.4]
  assign _T_81742 = _T_81741[13:0]; // @[Modules.scala 166:64:@28824.4]
  assign buffer_8_552 = $signed(_T_81742); // @[Modules.scala 166:64:@28825.4]
  assign _T_81744 = $signed(buffer_8_489) + $signed(buffer_8_490); // @[Modules.scala 166:64:@28827.4]
  assign _T_81745 = _T_81744[13:0]; // @[Modules.scala 166:64:@28828.4]
  assign buffer_8_553 = $signed(_T_81745); // @[Modules.scala 166:64:@28829.4]
  assign _T_81747 = $signed(buffer_8_491) + $signed(buffer_8_492); // @[Modules.scala 166:64:@28831.4]
  assign _T_81748 = _T_81747[13:0]; // @[Modules.scala 166:64:@28832.4]
  assign buffer_8_554 = $signed(_T_81748); // @[Modules.scala 166:64:@28833.4]
  assign _T_81750 = $signed(buffer_8_493) + $signed(buffer_8_494); // @[Modules.scala 166:64:@28835.4]
  assign _T_81751 = _T_81750[13:0]; // @[Modules.scala 166:64:@28836.4]
  assign buffer_8_555 = $signed(_T_81751); // @[Modules.scala 166:64:@28837.4]
  assign _T_81753 = $signed(buffer_8_495) + $signed(buffer_8_496); // @[Modules.scala 166:64:@28839.4]
  assign _T_81754 = _T_81753[13:0]; // @[Modules.scala 166:64:@28840.4]
  assign buffer_8_556 = $signed(_T_81754); // @[Modules.scala 166:64:@28841.4]
  assign _T_81756 = $signed(buffer_8_497) + $signed(buffer_8_498); // @[Modules.scala 166:64:@28843.4]
  assign _T_81757 = _T_81756[13:0]; // @[Modules.scala 166:64:@28844.4]
  assign buffer_8_557 = $signed(_T_81757); // @[Modules.scala 166:64:@28845.4]
  assign _T_81759 = $signed(buffer_8_499) + $signed(buffer_8_500); // @[Modules.scala 166:64:@28847.4]
  assign _T_81760 = _T_81759[13:0]; // @[Modules.scala 166:64:@28848.4]
  assign buffer_8_558 = $signed(_T_81760); // @[Modules.scala 166:64:@28849.4]
  assign _T_81762 = $signed(buffer_8_501) + $signed(buffer_8_502); // @[Modules.scala 166:64:@28851.4]
  assign _T_81763 = _T_81762[13:0]; // @[Modules.scala 166:64:@28852.4]
  assign buffer_8_559 = $signed(_T_81763); // @[Modules.scala 166:64:@28853.4]
  assign _T_81765 = $signed(buffer_8_503) + $signed(buffer_8_504); // @[Modules.scala 166:64:@28855.4]
  assign _T_81766 = _T_81765[13:0]; // @[Modules.scala 166:64:@28856.4]
  assign buffer_8_560 = $signed(_T_81766); // @[Modules.scala 166:64:@28857.4]
  assign _T_81768 = $signed(buffer_8_505) + $signed(buffer_8_506); // @[Modules.scala 166:64:@28859.4]
  assign _T_81769 = _T_81768[13:0]; // @[Modules.scala 166:64:@28860.4]
  assign buffer_8_561 = $signed(_T_81769); // @[Modules.scala 166:64:@28861.4]
  assign _T_81771 = $signed(buffer_8_507) + $signed(buffer_8_508); // @[Modules.scala 166:64:@28863.4]
  assign _T_81772 = _T_81771[13:0]; // @[Modules.scala 166:64:@28864.4]
  assign buffer_8_562 = $signed(_T_81772); // @[Modules.scala 166:64:@28865.4]
  assign _T_81774 = $signed(buffer_8_509) + $signed(buffer_8_510); // @[Modules.scala 166:64:@28867.4]
  assign _T_81775 = _T_81774[13:0]; // @[Modules.scala 166:64:@28868.4]
  assign buffer_8_563 = $signed(_T_81775); // @[Modules.scala 166:64:@28869.4]
  assign _T_81777 = $signed(buffer_8_511) + $signed(buffer_8_512); // @[Modules.scala 166:64:@28871.4]
  assign _T_81778 = _T_81777[13:0]; // @[Modules.scala 166:64:@28872.4]
  assign buffer_8_564 = $signed(_T_81778); // @[Modules.scala 166:64:@28873.4]
  assign _T_81780 = $signed(buffer_8_513) + $signed(buffer_8_514); // @[Modules.scala 166:64:@28875.4]
  assign _T_81781 = _T_81780[13:0]; // @[Modules.scala 166:64:@28876.4]
  assign buffer_8_565 = $signed(_T_81781); // @[Modules.scala 166:64:@28877.4]
  assign _T_81783 = $signed(buffer_8_515) + $signed(buffer_8_516); // @[Modules.scala 166:64:@28879.4]
  assign _T_81784 = _T_81783[13:0]; // @[Modules.scala 166:64:@28880.4]
  assign buffer_8_566 = $signed(_T_81784); // @[Modules.scala 166:64:@28881.4]
  assign _T_81786 = $signed(buffer_8_517) + $signed(buffer_8_518); // @[Modules.scala 166:64:@28883.4]
  assign _T_81787 = _T_81786[13:0]; // @[Modules.scala 166:64:@28884.4]
  assign buffer_8_567 = $signed(_T_81787); // @[Modules.scala 166:64:@28885.4]
  assign _T_81789 = $signed(buffer_8_519) + $signed(buffer_8_520); // @[Modules.scala 166:64:@28887.4]
  assign _T_81790 = _T_81789[13:0]; // @[Modules.scala 166:64:@28888.4]
  assign buffer_8_568 = $signed(_T_81790); // @[Modules.scala 166:64:@28889.4]
  assign _T_81792 = $signed(buffer_8_521) + $signed(buffer_8_522); // @[Modules.scala 166:64:@28891.4]
  assign _T_81793 = _T_81792[13:0]; // @[Modules.scala 166:64:@28892.4]
  assign buffer_8_569 = $signed(_T_81793); // @[Modules.scala 166:64:@28893.4]
  assign _T_81795 = $signed(buffer_8_523) + $signed(buffer_8_524); // @[Modules.scala 166:64:@28895.4]
  assign _T_81796 = _T_81795[13:0]; // @[Modules.scala 166:64:@28896.4]
  assign buffer_8_570 = $signed(_T_81796); // @[Modules.scala 166:64:@28897.4]
  assign _T_81798 = $signed(buffer_8_525) + $signed(buffer_8_526); // @[Modules.scala 166:64:@28899.4]
  assign _T_81799 = _T_81798[13:0]; // @[Modules.scala 166:64:@28900.4]
  assign buffer_8_571 = $signed(_T_81799); // @[Modules.scala 166:64:@28901.4]
  assign _T_81801 = $signed(buffer_8_527) + $signed(buffer_8_528); // @[Modules.scala 166:64:@28903.4]
  assign _T_81802 = _T_81801[13:0]; // @[Modules.scala 166:64:@28904.4]
  assign buffer_8_572 = $signed(_T_81802); // @[Modules.scala 166:64:@28905.4]
  assign _T_81804 = $signed(buffer_8_529) + $signed(buffer_8_530); // @[Modules.scala 166:64:@28907.4]
  assign _T_81805 = _T_81804[13:0]; // @[Modules.scala 166:64:@28908.4]
  assign buffer_8_573 = $signed(_T_81805); // @[Modules.scala 166:64:@28909.4]
  assign _T_81807 = $signed(buffer_5_540) + $signed(buffer_8_532); // @[Modules.scala 166:64:@28911.4]
  assign _T_81808 = _T_81807[13:0]; // @[Modules.scala 166:64:@28912.4]
  assign buffer_8_574 = $signed(_T_81808); // @[Modules.scala 166:64:@28913.4]
  assign _T_81810 = $signed(buffer_8_533) + $signed(buffer_8_534); // @[Modules.scala 166:64:@28915.4]
  assign _T_81811 = _T_81810[13:0]; // @[Modules.scala 166:64:@28916.4]
  assign buffer_8_575 = $signed(_T_81811); // @[Modules.scala 166:64:@28917.4]
  assign _T_81813 = $signed(buffer_8_535) + $signed(buffer_8_536); // @[Modules.scala 166:64:@28919.4]
  assign _T_81814 = _T_81813[13:0]; // @[Modules.scala 166:64:@28920.4]
  assign buffer_8_576 = $signed(_T_81814); // @[Modules.scala 166:64:@28921.4]
  assign _T_81816 = $signed(buffer_8_537) + $signed(buffer_8_538); // @[Modules.scala 166:64:@28923.4]
  assign _T_81817 = _T_81816[13:0]; // @[Modules.scala 166:64:@28924.4]
  assign buffer_8_577 = $signed(_T_81817); // @[Modules.scala 166:64:@28925.4]
  assign _T_81819 = $signed(buffer_8_539) + $signed(buffer_5_313); // @[Modules.scala 172:66:@28927.4]
  assign _T_81820 = _T_81819[13:0]; // @[Modules.scala 172:66:@28928.4]
  assign buffer_8_578 = $signed(_T_81820); // @[Modules.scala 172:66:@28929.4]
  assign _T_81822 = $signed(buffer_8_540) + $signed(buffer_8_541); // @[Modules.scala 166:64:@28931.4]
  assign _T_81823 = _T_81822[13:0]; // @[Modules.scala 166:64:@28932.4]
  assign buffer_8_579 = $signed(_T_81823); // @[Modules.scala 166:64:@28933.4]
  assign _T_81825 = $signed(buffer_8_542) + $signed(buffer_8_543); // @[Modules.scala 166:64:@28935.4]
  assign _T_81826 = _T_81825[13:0]; // @[Modules.scala 166:64:@28936.4]
  assign buffer_8_580 = $signed(_T_81826); // @[Modules.scala 166:64:@28937.4]
  assign _T_81828 = $signed(buffer_8_544) + $signed(buffer_8_545); // @[Modules.scala 166:64:@28939.4]
  assign _T_81829 = _T_81828[13:0]; // @[Modules.scala 166:64:@28940.4]
  assign buffer_8_581 = $signed(_T_81829); // @[Modules.scala 166:64:@28941.4]
  assign _T_81831 = $signed(buffer_8_546) + $signed(buffer_8_547); // @[Modules.scala 166:64:@28943.4]
  assign _T_81832 = _T_81831[13:0]; // @[Modules.scala 166:64:@28944.4]
  assign buffer_8_582 = $signed(_T_81832); // @[Modules.scala 166:64:@28945.4]
  assign _T_81834 = $signed(buffer_8_548) + $signed(buffer_8_549); // @[Modules.scala 166:64:@28947.4]
  assign _T_81835 = _T_81834[13:0]; // @[Modules.scala 166:64:@28948.4]
  assign buffer_8_583 = $signed(_T_81835); // @[Modules.scala 166:64:@28949.4]
  assign _T_81837 = $signed(buffer_8_550) + $signed(buffer_8_551); // @[Modules.scala 166:64:@28951.4]
  assign _T_81838 = _T_81837[13:0]; // @[Modules.scala 166:64:@28952.4]
  assign buffer_8_584 = $signed(_T_81838); // @[Modules.scala 166:64:@28953.4]
  assign _T_81840 = $signed(buffer_8_552) + $signed(buffer_8_553); // @[Modules.scala 166:64:@28955.4]
  assign _T_81841 = _T_81840[13:0]; // @[Modules.scala 166:64:@28956.4]
  assign buffer_8_585 = $signed(_T_81841); // @[Modules.scala 166:64:@28957.4]
  assign _T_81843 = $signed(buffer_8_554) + $signed(buffer_8_555); // @[Modules.scala 166:64:@28959.4]
  assign _T_81844 = _T_81843[13:0]; // @[Modules.scala 166:64:@28960.4]
  assign buffer_8_586 = $signed(_T_81844); // @[Modules.scala 166:64:@28961.4]
  assign _T_81846 = $signed(buffer_8_556) + $signed(buffer_8_557); // @[Modules.scala 166:64:@28963.4]
  assign _T_81847 = _T_81846[13:0]; // @[Modules.scala 166:64:@28964.4]
  assign buffer_8_587 = $signed(_T_81847); // @[Modules.scala 166:64:@28965.4]
  assign _T_81849 = $signed(buffer_8_558) + $signed(buffer_8_559); // @[Modules.scala 166:64:@28967.4]
  assign _T_81850 = _T_81849[13:0]; // @[Modules.scala 166:64:@28968.4]
  assign buffer_8_588 = $signed(_T_81850); // @[Modules.scala 166:64:@28969.4]
  assign _T_81852 = $signed(buffer_8_560) + $signed(buffer_8_561); // @[Modules.scala 166:64:@28971.4]
  assign _T_81853 = _T_81852[13:0]; // @[Modules.scala 166:64:@28972.4]
  assign buffer_8_589 = $signed(_T_81853); // @[Modules.scala 166:64:@28973.4]
  assign _T_81855 = $signed(buffer_8_562) + $signed(buffer_8_563); // @[Modules.scala 166:64:@28975.4]
  assign _T_81856 = _T_81855[13:0]; // @[Modules.scala 166:64:@28976.4]
  assign buffer_8_590 = $signed(_T_81856); // @[Modules.scala 166:64:@28977.4]
  assign _T_81858 = $signed(buffer_8_564) + $signed(buffer_8_565); // @[Modules.scala 166:64:@28979.4]
  assign _T_81859 = _T_81858[13:0]; // @[Modules.scala 166:64:@28980.4]
  assign buffer_8_591 = $signed(_T_81859); // @[Modules.scala 166:64:@28981.4]
  assign _T_81861 = $signed(buffer_8_566) + $signed(buffer_8_567); // @[Modules.scala 166:64:@28983.4]
  assign _T_81862 = _T_81861[13:0]; // @[Modules.scala 166:64:@28984.4]
  assign buffer_8_592 = $signed(_T_81862); // @[Modules.scala 166:64:@28985.4]
  assign _T_81864 = $signed(buffer_8_568) + $signed(buffer_8_569); // @[Modules.scala 166:64:@28987.4]
  assign _T_81865 = _T_81864[13:0]; // @[Modules.scala 166:64:@28988.4]
  assign buffer_8_593 = $signed(_T_81865); // @[Modules.scala 166:64:@28989.4]
  assign _T_81867 = $signed(buffer_8_570) + $signed(buffer_8_571); // @[Modules.scala 166:64:@28991.4]
  assign _T_81868 = _T_81867[13:0]; // @[Modules.scala 166:64:@28992.4]
  assign buffer_8_594 = $signed(_T_81868); // @[Modules.scala 166:64:@28993.4]
  assign _T_81870 = $signed(buffer_8_572) + $signed(buffer_8_573); // @[Modules.scala 166:64:@28995.4]
  assign _T_81871 = _T_81870[13:0]; // @[Modules.scala 166:64:@28996.4]
  assign buffer_8_595 = $signed(_T_81871); // @[Modules.scala 166:64:@28997.4]
  assign _T_81873 = $signed(buffer_8_574) + $signed(buffer_8_575); // @[Modules.scala 166:64:@28999.4]
  assign _T_81874 = _T_81873[13:0]; // @[Modules.scala 166:64:@29000.4]
  assign buffer_8_596 = $signed(_T_81874); // @[Modules.scala 166:64:@29001.4]
  assign _T_81876 = $signed(buffer_8_576) + $signed(buffer_8_577); // @[Modules.scala 166:64:@29003.4]
  assign _T_81877 = _T_81876[13:0]; // @[Modules.scala 166:64:@29004.4]
  assign buffer_8_597 = $signed(_T_81877); // @[Modules.scala 166:64:@29005.4]
  assign _T_81879 = $signed(buffer_8_579) + $signed(buffer_8_580); // @[Modules.scala 166:64:@29007.4]
  assign _T_81880 = _T_81879[13:0]; // @[Modules.scala 166:64:@29008.4]
  assign buffer_8_598 = $signed(_T_81880); // @[Modules.scala 166:64:@29009.4]
  assign _T_81882 = $signed(buffer_8_581) + $signed(buffer_8_582); // @[Modules.scala 166:64:@29011.4]
  assign _T_81883 = _T_81882[13:0]; // @[Modules.scala 166:64:@29012.4]
  assign buffer_8_599 = $signed(_T_81883); // @[Modules.scala 166:64:@29013.4]
  assign _T_81885 = $signed(buffer_8_583) + $signed(buffer_8_584); // @[Modules.scala 166:64:@29015.4]
  assign _T_81886 = _T_81885[13:0]; // @[Modules.scala 166:64:@29016.4]
  assign buffer_8_600 = $signed(_T_81886); // @[Modules.scala 166:64:@29017.4]
  assign _T_81888 = $signed(buffer_8_585) + $signed(buffer_8_586); // @[Modules.scala 166:64:@29019.4]
  assign _T_81889 = _T_81888[13:0]; // @[Modules.scala 166:64:@29020.4]
  assign buffer_8_601 = $signed(_T_81889); // @[Modules.scala 166:64:@29021.4]
  assign _T_81891 = $signed(buffer_8_587) + $signed(buffer_8_588); // @[Modules.scala 166:64:@29023.4]
  assign _T_81892 = _T_81891[13:0]; // @[Modules.scala 166:64:@29024.4]
  assign buffer_8_602 = $signed(_T_81892); // @[Modules.scala 166:64:@29025.4]
  assign _T_81894 = $signed(buffer_8_589) + $signed(buffer_8_590); // @[Modules.scala 166:64:@29027.4]
  assign _T_81895 = _T_81894[13:0]; // @[Modules.scala 166:64:@29028.4]
  assign buffer_8_603 = $signed(_T_81895); // @[Modules.scala 166:64:@29029.4]
  assign _T_81897 = $signed(buffer_8_591) + $signed(buffer_8_592); // @[Modules.scala 166:64:@29031.4]
  assign _T_81898 = _T_81897[13:0]; // @[Modules.scala 166:64:@29032.4]
  assign buffer_8_604 = $signed(_T_81898); // @[Modules.scala 166:64:@29033.4]
  assign _T_81900 = $signed(buffer_8_593) + $signed(buffer_8_594); // @[Modules.scala 166:64:@29035.4]
  assign _T_81901 = _T_81900[13:0]; // @[Modules.scala 166:64:@29036.4]
  assign buffer_8_605 = $signed(_T_81901); // @[Modules.scala 166:64:@29037.4]
  assign _T_81903 = $signed(buffer_8_595) + $signed(buffer_8_596); // @[Modules.scala 166:64:@29039.4]
  assign _T_81904 = _T_81903[13:0]; // @[Modules.scala 166:64:@29040.4]
  assign buffer_8_606 = $signed(_T_81904); // @[Modules.scala 166:64:@29041.4]
  assign _T_81906 = $signed(buffer_8_597) + $signed(buffer_8_578); // @[Modules.scala 172:66:@29043.4]
  assign _T_81907 = _T_81906[13:0]; // @[Modules.scala 172:66:@29044.4]
  assign buffer_8_607 = $signed(_T_81907); // @[Modules.scala 172:66:@29045.4]
  assign _T_81909 = $signed(buffer_8_598) + $signed(buffer_8_599); // @[Modules.scala 160:64:@29047.4]
  assign _T_81910 = _T_81909[13:0]; // @[Modules.scala 160:64:@29048.4]
  assign buffer_8_608 = $signed(_T_81910); // @[Modules.scala 160:64:@29049.4]
  assign _T_81912 = $signed(buffer_8_600) + $signed(buffer_8_601); // @[Modules.scala 160:64:@29051.4]
  assign _T_81913 = _T_81912[13:0]; // @[Modules.scala 160:64:@29052.4]
  assign buffer_8_609 = $signed(_T_81913); // @[Modules.scala 160:64:@29053.4]
  assign _T_81915 = $signed(buffer_8_602) + $signed(buffer_8_603); // @[Modules.scala 160:64:@29055.4]
  assign _T_81916 = _T_81915[13:0]; // @[Modules.scala 160:64:@29056.4]
  assign buffer_8_610 = $signed(_T_81916); // @[Modules.scala 160:64:@29057.4]
  assign _T_81918 = $signed(buffer_8_604) + $signed(buffer_8_605); // @[Modules.scala 160:64:@29059.4]
  assign _T_81919 = _T_81918[13:0]; // @[Modules.scala 160:64:@29060.4]
  assign buffer_8_611 = $signed(_T_81919); // @[Modules.scala 160:64:@29061.4]
  assign _T_81921 = $signed(buffer_8_606) + $signed(buffer_8_607); // @[Modules.scala 160:64:@29063.4]
  assign _T_81922 = _T_81921[13:0]; // @[Modules.scala 160:64:@29064.4]
  assign buffer_8_612 = $signed(_T_81922); // @[Modules.scala 160:64:@29065.4]
  assign _T_81924 = $signed(buffer_8_608) + $signed(buffer_8_609); // @[Modules.scala 166:64:@29067.4]
  assign _T_81925 = _T_81924[13:0]; // @[Modules.scala 166:64:@29068.4]
  assign buffer_8_613 = $signed(_T_81925); // @[Modules.scala 166:64:@29069.4]
  assign _T_81927 = $signed(buffer_8_610) + $signed(buffer_8_611); // @[Modules.scala 166:64:@29071.4]
  assign _T_81928 = _T_81927[13:0]; // @[Modules.scala 166:64:@29072.4]
  assign buffer_8_614 = $signed(_T_81928); // @[Modules.scala 166:64:@29073.4]
  assign _T_81930 = $signed(buffer_8_613) + $signed(buffer_8_614); // @[Modules.scala 160:64:@29075.4]
  assign _T_81931 = _T_81930[13:0]; // @[Modules.scala 160:64:@29076.4]
  assign buffer_8_615 = $signed(_T_81931); // @[Modules.scala 160:64:@29077.4]
  assign _T_81933 = $signed(buffer_8_615) + $signed(buffer_8_612); // @[Modules.scala 172:66:@29079.4]
  assign _T_81934 = _T_81933[13:0]; // @[Modules.scala 172:66:@29080.4]
  assign buffer_8_616 = $signed(_T_81934); // @[Modules.scala 172:66:@29081.4]
  assign _GEN_633 = {{1{_T_60269[4]}},_T_60269}; // @[Modules.scala 143:103:@29270.4]
  assign _T_81961 = $signed(_GEN_633) + $signed(_T_57234); // @[Modules.scala 143:103:@29270.4]
  assign _T_81962 = _T_81961[5:0]; // @[Modules.scala 143:103:@29271.4]
  assign _T_81963 = $signed(_T_81962); // @[Modules.scala 143:103:@29272.4]
  assign _T_81982 = $signed(_T_54236) + $signed(_T_54241); // @[Modules.scala 143:103:@29288.4]
  assign _T_81983 = _T_81982[5:0]; // @[Modules.scala 143:103:@29289.4]
  assign _T_81984 = $signed(_T_81983); // @[Modules.scala 143:103:@29290.4]
  assign _T_81989 = $signed(_T_54243) + $signed(_T_54248); // @[Modules.scala 143:103:@29294.4]
  assign _T_81990 = _T_81989[5:0]; // @[Modules.scala 143:103:@29295.4]
  assign _T_81991 = $signed(_T_81990); // @[Modules.scala 143:103:@29296.4]
  assign _T_81996 = $signed(_T_54250) + $signed(_T_54255); // @[Modules.scala 143:103:@29300.4]
  assign _T_81997 = _T_81996[5:0]; // @[Modules.scala 143:103:@29301.4]
  assign _T_81998 = $signed(_T_81997); // @[Modules.scala 143:103:@29302.4]
  assign _T_82010 = $signed(_T_54264) + $signed(_T_54269); // @[Modules.scala 143:103:@29312.4]
  assign _T_82011 = _T_82010[5:0]; // @[Modules.scala 143:103:@29313.4]
  assign _T_82012 = $signed(_T_82011); // @[Modules.scala 143:103:@29314.4]
  assign _T_82038 = $signed(_GEN_81) + $signed(_T_54292); // @[Modules.scala 143:103:@29336.4]
  assign _T_82039 = _T_82038[5:0]; // @[Modules.scala 143:103:@29337.4]
  assign _T_82040 = $signed(_T_82039); // @[Modules.scala 143:103:@29338.4]
  assign _T_82094 = $signed(_T_54346) + $signed(_GEN_431); // @[Modules.scala 143:103:@29384.4]
  assign _T_82095 = _T_82094[5:0]; // @[Modules.scala 143:103:@29385.4]
  assign _T_82096 = $signed(_T_82095); // @[Modules.scala 143:103:@29386.4]
  assign _T_82143 = $signed(_T_54397) + $signed(_T_54402); // @[Modules.scala 143:103:@29426.4]
  assign _T_82144 = _T_82143[5:0]; // @[Modules.scala 143:103:@29427.4]
  assign _T_82145 = $signed(_T_82144); // @[Modules.scala 143:103:@29428.4]
  assign _T_82199 = $signed(_T_54451) + $signed(_T_60488); // @[Modules.scala 143:103:@29474.4]
  assign _T_82200 = _T_82199[5:0]; // @[Modules.scala 143:103:@29475.4]
  assign _T_82201 = $signed(_T_82200); // @[Modules.scala 143:103:@29476.4]
  assign _GEN_637 = {{1{_T_63606[4]}},_T_63606}; // @[Modules.scala 143:103:@29480.4]
  assign _T_82206 = $signed(_T_54460) + $signed(_GEN_637); // @[Modules.scala 143:103:@29480.4]
  assign _T_82207 = _T_82206[5:0]; // @[Modules.scala 143:103:@29481.4]
  assign _T_82208 = $signed(_T_82207); // @[Modules.scala 143:103:@29482.4]
  assign _T_82227 = $signed(_T_60509) + $signed(_T_60514); // @[Modules.scala 143:103:@29498.4]
  assign _T_82228 = _T_82227[4:0]; // @[Modules.scala 143:103:@29499.4]
  assign _T_82229 = $signed(_T_82228); // @[Modules.scala 143:103:@29500.4]
  assign _T_82234 = $signed(_GEN_85) + $signed(_T_54493); // @[Modules.scala 143:103:@29504.4]
  assign _T_82235 = _T_82234[5:0]; // @[Modules.scala 143:103:@29505.4]
  assign _T_82236 = $signed(_T_82235); // @[Modules.scala 143:103:@29506.4]
  assign _GEN_639 = {{1{_T_69763[4]}},_T_69763}; // @[Modules.scala 143:103:@29510.4]
  assign _T_82241 = $signed(_T_54495) + $signed(_GEN_639); // @[Modules.scala 143:103:@29510.4]
  assign _T_82242 = _T_82241[5:0]; // @[Modules.scala 143:103:@29511.4]
  assign _T_82243 = $signed(_T_82242); // @[Modules.scala 143:103:@29512.4]
  assign _T_82262 = $signed(_T_57514) + $signed(_GEN_152); // @[Modules.scala 143:103:@29528.4]
  assign _T_82263 = _T_82262[5:0]; // @[Modules.scala 143:103:@29529.4]
  assign _T_82264 = $signed(_T_82263); // @[Modules.scala 143:103:@29530.4]
  assign _GEN_642 = {{1{_T_60579[4]}},_T_60579}; // @[Modules.scala 143:103:@29558.4]
  assign _T_82297 = $signed(_T_54535) + $signed(_GEN_642); // @[Modules.scala 143:103:@29558.4]
  assign _T_82298 = _T_82297[5:0]; // @[Modules.scala 143:103:@29559.4]
  assign _T_82299 = $signed(_T_82298); // @[Modules.scala 143:103:@29560.4]
  assign _T_82325 = $signed(_GEN_87) + $signed(_T_60605); // @[Modules.scala 143:103:@29582.4]
  assign _T_82326 = _T_82325[5:0]; // @[Modules.scala 143:103:@29583.4]
  assign _T_82327 = $signed(_T_82326); // @[Modules.scala 143:103:@29584.4]
  assign _T_82353 = $signed(_T_54572) + $signed(_GEN_12); // @[Modules.scala 143:103:@29606.4]
  assign _T_82354 = _T_82353[5:0]; // @[Modules.scala 143:103:@29607.4]
  assign _T_82355 = $signed(_T_82354); // @[Modules.scala 143:103:@29608.4]
  assign _T_82360 = $signed(_T_60633) + $signed(_T_54586); // @[Modules.scala 143:103:@29612.4]
  assign _T_82361 = _T_82360[5:0]; // @[Modules.scala 143:103:@29613.4]
  assign _T_82362 = $signed(_T_82361); // @[Modules.scala 143:103:@29614.4]
  assign _T_82381 = $signed(_T_54605) + $signed(_T_73021); // @[Modules.scala 143:103:@29630.4]
  assign _T_82382 = _T_82381[5:0]; // @[Modules.scala 143:103:@29631.4]
  assign _T_82383 = $signed(_T_82382); // @[Modules.scala 143:103:@29632.4]
  assign _GEN_646 = {{1{_T_63835[4]}},_T_63835}; // @[Modules.scala 143:103:@29678.4]
  assign _T_82437 = $signed(_T_57675) + $signed(_GEN_646); // @[Modules.scala 143:103:@29678.4]
  assign _T_82438 = _T_82437[5:0]; // @[Modules.scala 143:103:@29679.4]
  assign _T_82439 = $signed(_T_82438); // @[Modules.scala 143:103:@29680.4]
  assign _T_82451 = $signed(_T_54675) + $signed(_GEN_164); // @[Modules.scala 143:103:@29690.4]
  assign _T_82452 = _T_82451[5:0]; // @[Modules.scala 143:103:@29691.4]
  assign _T_82453 = $signed(_T_82452); // @[Modules.scala 143:103:@29692.4]
  assign _T_82458 = $signed(_GEN_16) + $signed(_T_57708); // @[Modules.scala 143:103:@29696.4]
  assign _T_82459 = _T_82458[5:0]; // @[Modules.scala 143:103:@29697.4]
  assign _T_82460 = $signed(_T_82459); // @[Modules.scala 143:103:@29698.4]
  assign _T_82465 = $signed(_T_57710) + $signed(_GEN_229); // @[Modules.scala 143:103:@29702.4]
  assign _T_82466 = _T_82465[5:0]; // @[Modules.scala 143:103:@29703.4]
  assign _T_82467 = $signed(_T_82466); // @[Modules.scala 143:103:@29704.4]
  assign _T_82479 = $signed(_T_54691) + $signed(_T_54696); // @[Modules.scala 143:103:@29714.4]
  assign _T_82480 = _T_82479[4:0]; // @[Modules.scala 143:103:@29715.4]
  assign _T_82481 = $signed(_T_82480); // @[Modules.scala 143:103:@29716.4]
  assign _T_82486 = $signed(_T_63884) + $signed(_GEN_446); // @[Modules.scala 143:103:@29720.4]
  assign _T_82487 = _T_82486[5:0]; // @[Modules.scala 143:103:@29721.4]
  assign _T_82488 = $signed(_T_82487); // @[Modules.scala 143:103:@29722.4]
  assign _T_82528 = $signed(_T_57787) + $signed(_T_60829); // @[Modules.scala 143:103:@29756.4]
  assign _T_82529 = _T_82528[4:0]; // @[Modules.scala 143:103:@29757.4]
  assign _T_82530 = $signed(_T_82529); // @[Modules.scala 143:103:@29758.4]
  assign _T_82535 = $signed(_T_54759) + $signed(_T_60831); // @[Modules.scala 143:103:@29762.4]
  assign _T_82536 = _T_82535[4:0]; // @[Modules.scala 143:103:@29763.4]
  assign _T_82537 = $signed(_T_82536); // @[Modules.scala 143:103:@29764.4]
  assign _T_82542 = $signed(_T_57794) + $signed(_T_60838); // @[Modules.scala 143:103:@29768.4]
  assign _T_82543 = _T_82542[4:0]; // @[Modules.scala 143:103:@29769.4]
  assign _T_82544 = $signed(_T_82543); // @[Modules.scala 143:103:@29770.4]
  assign _T_82570 = $signed(_GEN_299) + $signed(_T_63970); // @[Modules.scala 143:103:@29792.4]
  assign _T_82571 = _T_82570[5:0]; // @[Modules.scala 143:103:@29793.4]
  assign _T_82572 = $signed(_T_82571); // @[Modules.scala 143:103:@29794.4]
  assign _GEN_652 = {{1{_T_54789[4]}},_T_54789}; // @[Modules.scala 143:103:@29798.4]
  assign _T_82577 = $signed(_GEN_652) + $signed(_T_63977); // @[Modules.scala 143:103:@29798.4]
  assign _T_82578 = _T_82577[5:0]; // @[Modules.scala 143:103:@29799.4]
  assign _T_82579 = $signed(_T_82578); // @[Modules.scala 143:103:@29800.4]
  assign _T_82619 = $signed(_T_57869) + $signed(_T_54829); // @[Modules.scala 143:103:@29834.4]
  assign _T_82620 = _T_82619[4:0]; // @[Modules.scala 143:103:@29835.4]
  assign _T_82621 = $signed(_T_82620); // @[Modules.scala 143:103:@29836.4]
  assign _T_82654 = $signed(_T_54859) + $signed(_T_54864); // @[Modules.scala 143:103:@29864.4]
  assign _T_82655 = _T_82654[4:0]; // @[Modules.scala 143:103:@29865.4]
  assign _T_82656 = $signed(_T_82655); // @[Modules.scala 143:103:@29866.4]
  assign _T_82661 = $signed(_T_54866) + $signed(_T_54871); // @[Modules.scala 143:103:@29870.4]
  assign _T_82662 = _T_82661[4:0]; // @[Modules.scala 143:103:@29871.4]
  assign _T_82663 = $signed(_T_82662); // @[Modules.scala 143:103:@29872.4]
  assign _T_82668 = $signed(_T_54873) + $signed(_T_54878); // @[Modules.scala 143:103:@29876.4]
  assign _T_82669 = _T_82668[4:0]; // @[Modules.scala 143:103:@29877.4]
  assign _T_82670 = $signed(_T_82669); // @[Modules.scala 143:103:@29878.4]
  assign _GEN_654 = {{1{_T_54894[4]}},_T_54894}; // @[Modules.scala 143:103:@29894.4]
  assign _T_82689 = $signed(_GEN_654) + $signed(_T_54899); // @[Modules.scala 143:103:@29894.4]
  assign _T_82690 = _T_82689[5:0]; // @[Modules.scala 143:103:@29895.4]
  assign _T_82691 = $signed(_T_82690); // @[Modules.scala 143:103:@29896.4]
  assign _T_82731 = $signed(_T_54936) + $signed(_T_54941); // @[Modules.scala 143:103:@29930.4]
  assign _T_82732 = _T_82731[4:0]; // @[Modules.scala 143:103:@29931.4]
  assign _T_82733 = $signed(_T_82732); // @[Modules.scala 143:103:@29932.4]
  assign _GEN_655 = {{1{_T_61025[4]}},_T_61025}; // @[Modules.scala 143:103:@29936.4]
  assign _T_82738 = $signed(_T_54948) + $signed(_GEN_655); // @[Modules.scala 143:103:@29936.4]
  assign _T_82739 = _T_82738[5:0]; // @[Modules.scala 143:103:@29937.4]
  assign _T_82740 = $signed(_T_82739); // @[Modules.scala 143:103:@29938.4]
  assign _T_82780 = $signed(_GEN_519) + $signed(_T_54990); // @[Modules.scala 143:103:@29972.4]
  assign _T_82781 = _T_82780[5:0]; // @[Modules.scala 143:103:@29973.4]
  assign _T_82782 = $signed(_T_82781); // @[Modules.scala 143:103:@29974.4]
  assign _T_82787 = $signed(_T_54992) + $signed(_T_54999); // @[Modules.scala 143:103:@29978.4]
  assign _T_82788 = _T_82787[4:0]; // @[Modules.scala 143:103:@29979.4]
  assign _T_82789 = $signed(_T_82788); // @[Modules.scala 143:103:@29980.4]
  assign _GEN_657 = {{1{_T_55011[4]}},_T_55011}; // @[Modules.scala 143:103:@29990.4]
  assign _T_82801 = $signed(_GEN_657) + $signed(_T_61088); // @[Modules.scala 143:103:@29990.4]
  assign _T_82802 = _T_82801[5:0]; // @[Modules.scala 143:103:@29991.4]
  assign _T_82803 = $signed(_T_82802); // @[Modules.scala 143:103:@29992.4]
  assign _GEN_658 = {{1{_T_55020[4]}},_T_55020}; // @[Modules.scala 143:103:@29996.4]
  assign _T_82808 = $signed(_GEN_658) + $signed(_T_61097); // @[Modules.scala 143:103:@29996.4]
  assign _T_82809 = _T_82808[5:0]; // @[Modules.scala 143:103:@29997.4]
  assign _T_82810 = $signed(_T_82809); // @[Modules.scala 143:103:@29998.4]
  assign _T_82815 = $signed(_T_58053) + $signed(_T_58058); // @[Modules.scala 143:103:@30002.4]
  assign _T_82816 = _T_82815[5:0]; // @[Modules.scala 143:103:@30003.4]
  assign _T_82817 = $signed(_T_82816); // @[Modules.scala 143:103:@30004.4]
  assign _T_82829 = $signed(_T_55041) + $signed(_T_55046); // @[Modules.scala 143:103:@30014.4]
  assign _T_82830 = _T_82829[4:0]; // @[Modules.scala 143:103:@30015.4]
  assign _T_82831 = $signed(_T_82830); // @[Modules.scala 143:103:@30016.4]
  assign _T_82836 = $signed(_T_55048) + $signed(_T_55053); // @[Modules.scala 143:103:@30020.4]
  assign _T_82837 = _T_82836[4:0]; // @[Modules.scala 143:103:@30021.4]
  assign _T_82838 = $signed(_T_82837); // @[Modules.scala 143:103:@30022.4]
  assign _T_82878 = $signed(_T_61153) + $signed(_T_55088); // @[Modules.scala 143:103:@30056.4]
  assign _T_82879 = _T_82878[4:0]; // @[Modules.scala 143:103:@30057.4]
  assign _T_82880 = $signed(_T_82879); // @[Modules.scala 143:103:@30058.4]
  assign _T_82885 = $signed(_GEN_461) + $signed(_T_61160); // @[Modules.scala 143:103:@30062.4]
  assign _T_82886 = _T_82885[5:0]; // @[Modules.scala 143:103:@30063.4]
  assign _T_82887 = $signed(_T_82886); // @[Modules.scala 143:103:@30064.4]
  assign _T_82920 = $signed(_T_55125) + $signed(_GEN_312); // @[Modules.scala 143:103:@30092.4]
  assign _T_82921 = _T_82920[5:0]; // @[Modules.scala 143:103:@30093.4]
  assign _T_82922 = $signed(_T_82921); // @[Modules.scala 143:103:@30094.4]
  assign _T_82927 = $signed(_T_73565) + $signed(_T_76696); // @[Modules.scala 143:103:@30098.4]
  assign _T_82928 = _T_82927[4:0]; // @[Modules.scala 143:103:@30099.4]
  assign _T_82929 = $signed(_T_82928); // @[Modules.scala 143:103:@30100.4]
  assign _T_82934 = $signed(_T_64334) + $signed(_T_55139); // @[Modules.scala 143:103:@30104.4]
  assign _T_82935 = _T_82934[4:0]; // @[Modules.scala 143:103:@30105.4]
  assign _T_82936 = $signed(_T_82935); // @[Modules.scala 143:103:@30106.4]
  assign _T_82962 = $signed(_T_61235) + $signed(_T_58191); // @[Modules.scala 143:103:@30128.4]
  assign _T_82963 = _T_82962[4:0]; // @[Modules.scala 143:103:@30129.4]
  assign _T_82964 = $signed(_T_82963); // @[Modules.scala 143:103:@30130.4]
  assign _T_83011 = $signed(_T_55214) + $signed(_T_58240); // @[Modules.scala 143:103:@30170.4]
  assign _T_83012 = _T_83011[5:0]; // @[Modules.scala 143:103:@30171.4]
  assign _T_83013 = $signed(_T_83012); // @[Modules.scala 143:103:@30172.4]
  assign _T_83018 = $signed(_T_76787) + $signed(_T_55223); // @[Modules.scala 143:103:@30176.4]
  assign _T_83019 = _T_83018[4:0]; // @[Modules.scala 143:103:@30177.4]
  assign _T_83020 = $signed(_T_83019); // @[Modules.scala 143:103:@30178.4]
  assign _T_83039 = $signed(_T_61326) + $signed(_T_58277); // @[Modules.scala 143:103:@30194.4]
  assign _T_83040 = _T_83039[4:0]; // @[Modules.scala 143:103:@30195.4]
  assign _T_83041 = $signed(_T_83040); // @[Modules.scala 143:103:@30196.4]
  assign _T_83088 = $signed(_GEN_390) + $signed(_T_61384); // @[Modules.scala 143:103:@30236.4]
  assign _T_83089 = _T_83088[5:0]; // @[Modules.scala 143:103:@30237.4]
  assign _T_83090 = $signed(_T_83089); // @[Modules.scala 143:103:@30238.4]
  assign _T_83095 = $signed(_T_61391) + $signed(_T_55314); // @[Modules.scala 143:103:@30242.4]
  assign _T_83096 = _T_83095[5:0]; // @[Modules.scala 143:103:@30243.4]
  assign _T_83097 = $signed(_T_83096); // @[Modules.scala 143:103:@30244.4]
  assign _T_83102 = $signed(_T_61398) + $signed(_T_61403); // @[Modules.scala 143:103:@30248.4]
  assign _T_83103 = _T_83102[5:0]; // @[Modules.scala 143:103:@30249.4]
  assign _T_83104 = $signed(_T_83103); // @[Modules.scala 143:103:@30250.4]
  assign _T_83116 = $signed(_T_61412) + $signed(_T_58352); // @[Modules.scala 143:103:@30260.4]
  assign _T_83117 = _T_83116[4:0]; // @[Modules.scala 143:103:@30261.4]
  assign _T_83118 = $signed(_T_83117); // @[Modules.scala 143:103:@30262.4]
  assign _T_83123 = $signed(_T_61419) + $signed(_T_55335); // @[Modules.scala 143:103:@30266.4]
  assign _T_83124 = _T_83123[5:0]; // @[Modules.scala 143:103:@30267.4]
  assign _T_83125 = $signed(_T_83124); // @[Modules.scala 143:103:@30268.4]
  assign _T_83144 = $signed(_T_61438) + $signed(_T_64549); // @[Modules.scala 143:103:@30284.4]
  assign _T_83145 = _T_83144[5:0]; // @[Modules.scala 143:103:@30285.4]
  assign _T_83146 = $signed(_T_83145); // @[Modules.scala 143:103:@30286.4]
  assign _T_83151 = $signed(_T_61440) + $signed(_T_61447); // @[Modules.scala 143:103:@30290.4]
  assign _T_83152 = _T_83151[5:0]; // @[Modules.scala 143:103:@30291.4]
  assign _T_83153 = $signed(_T_83152); // @[Modules.scala 143:103:@30292.4]
  assign _T_83165 = $signed(_T_55375) + $signed(_T_61468); // @[Modules.scala 143:103:@30302.4]
  assign _T_83166 = _T_83165[5:0]; // @[Modules.scala 143:103:@30303.4]
  assign _T_83167 = $signed(_T_83166); // @[Modules.scala 143:103:@30304.4]
  assign _T_83179 = $signed(_T_55396) + $signed(_T_58403); // @[Modules.scala 143:103:@30314.4]
  assign _T_83180 = _T_83179[5:0]; // @[Modules.scala 143:103:@30315.4]
  assign _T_83181 = $signed(_T_83180); // @[Modules.scala 143:103:@30316.4]
  assign _T_83183 = $signed(4'sh1) * $signed(io_in_443); // @[Modules.scala 143:74:@30318.4]
  assign _T_83186 = $signed(_T_83183) + $signed(_T_61489); // @[Modules.scala 143:103:@30320.4]
  assign _T_83187 = _T_83186[5:0]; // @[Modules.scala 143:103:@30321.4]
  assign _T_83188 = $signed(_T_83187); // @[Modules.scala 143:103:@30322.4]
  assign _GEN_664 = {{1{_T_58417[4]}},_T_58417}; // @[Modules.scala 143:103:@30326.4]
  assign _T_83193 = $signed(_T_55405) + $signed(_GEN_664); // @[Modules.scala 143:103:@30326.4]
  assign _T_83194 = _T_83193[5:0]; // @[Modules.scala 143:103:@30327.4]
  assign _T_83195 = $signed(_T_83194); // @[Modules.scala 143:103:@30328.4]
  assign _T_83207 = $signed(_T_61503) + $signed(_T_55424); // @[Modules.scala 143:103:@30338.4]
  assign _T_83208 = _T_83207[5:0]; // @[Modules.scala 143:103:@30339.4]
  assign _T_83209 = $signed(_T_83208); // @[Modules.scala 143:103:@30340.4]
  assign _GEN_665 = {{1{_T_55431[4]}},_T_55431}; // @[Modules.scala 143:103:@30344.4]
  assign _T_83214 = $signed(_T_55426) + $signed(_GEN_665); // @[Modules.scala 143:103:@30344.4]
  assign _T_83215 = _T_83214[5:0]; // @[Modules.scala 143:103:@30345.4]
  assign _T_83216 = $signed(_T_83215); // @[Modules.scala 143:103:@30346.4]
  assign _T_83256 = $signed(_T_55459) + $signed(_T_58480); // @[Modules.scala 143:103:@30380.4]
  assign _T_83257 = _T_83256[5:0]; // @[Modules.scala 143:103:@30381.4]
  assign _T_83258 = $signed(_T_83257); // @[Modules.scala 143:103:@30382.4]
  assign _T_83284 = $signed(_T_58494) + $signed(_T_61573); // @[Modules.scala 143:103:@30404.4]
  assign _T_83285 = _T_83284[4:0]; // @[Modules.scala 143:103:@30405.4]
  assign _T_83286 = $signed(_T_83285); // @[Modules.scala 143:103:@30406.4]
  assign _T_83340 = $signed(_T_55522) + $signed(_T_70829); // @[Modules.scala 143:103:@30452.4]
  assign _T_83341 = _T_83340[5:0]; // @[Modules.scala 143:103:@30453.4]
  assign _T_83342 = $signed(_T_83341); // @[Modules.scala 143:103:@30454.4]
  assign _T_83347 = $signed(_T_58557) + $signed(_T_67765); // @[Modules.scala 143:103:@30458.4]
  assign _T_83348 = _T_83347[5:0]; // @[Modules.scala 143:103:@30459.4]
  assign _T_83349 = $signed(_T_83348); // @[Modules.scala 143:103:@30460.4]
  assign _T_83354 = $signed(_T_67767) + $signed(_T_58569); // @[Modules.scala 143:103:@30464.4]
  assign _T_83355 = _T_83354[5:0]; // @[Modules.scala 143:103:@30465.4]
  assign _T_83356 = $signed(_T_83355); // @[Modules.scala 143:103:@30466.4]
  assign _GEN_668 = {{1{_T_58576[4]}},_T_58576}; // @[Modules.scala 143:103:@30470.4]
  assign _T_83361 = $signed(_T_55543) + $signed(_GEN_668); // @[Modules.scala 143:103:@30470.4]
  assign _T_83362 = _T_83361[5:0]; // @[Modules.scala 143:103:@30471.4]
  assign _T_83363 = $signed(_T_83362); // @[Modules.scala 143:103:@30472.4]
  assign _T_83375 = $signed(_T_61643) + $signed(_T_55559); // @[Modules.scala 143:103:@30482.4]
  assign _T_83376 = _T_83375[4:0]; // @[Modules.scala 143:103:@30483.4]
  assign _T_83377 = $signed(_T_83376); // @[Modules.scala 143:103:@30484.4]
  assign _GEN_669 = {{1{_T_61662[4]}},_T_61662}; // @[Modules.scala 143:103:@30494.4]
  assign _T_83389 = $signed(_T_55571) + $signed(_GEN_669); // @[Modules.scala 143:103:@30494.4]
  assign _T_83390 = _T_83389[5:0]; // @[Modules.scala 143:103:@30495.4]
  assign _T_83391 = $signed(_T_83390); // @[Modules.scala 143:103:@30496.4]
  assign _T_83438 = $signed(_T_55620) + $signed(_T_55627); // @[Modules.scala 143:103:@30536.4]
  assign _T_83439 = _T_83438[5:0]; // @[Modules.scala 143:103:@30537.4]
  assign _T_83440 = $signed(_T_83439); // @[Modules.scala 143:103:@30538.4]
  assign _GEN_672 = {{1{_T_58641[4]}},_T_58641}; // @[Modules.scala 143:103:@30542.4]
  assign _T_83445 = $signed(_T_55629) + $signed(_GEN_672); // @[Modules.scala 143:103:@30542.4]
  assign _T_83446 = _T_83445[5:0]; // @[Modules.scala 143:103:@30543.4]
  assign _T_83447 = $signed(_T_83446); // @[Modules.scala 143:103:@30544.4]
  assign _GEN_673 = {{1{_T_58674[4]}},_T_58674}; // @[Modules.scala 143:103:@30566.4]
  assign _T_83473 = $signed(_T_55657) + $signed(_GEN_673); // @[Modules.scala 143:103:@30566.4]
  assign _T_83474 = _T_83473[5:0]; // @[Modules.scala 143:103:@30567.4]
  assign _T_83475 = $signed(_T_83474); // @[Modules.scala 143:103:@30568.4]
  assign _T_83501 = $signed(_T_55690) + $signed(_GEN_194); // @[Modules.scala 143:103:@30590.4]
  assign _T_83502 = _T_83501[5:0]; // @[Modules.scala 143:103:@30591.4]
  assign _T_83503 = $signed(_T_83502); // @[Modules.scala 143:103:@30592.4]
  assign _T_83508 = $signed(_T_55706) + $signed(_T_55711); // @[Modules.scala 143:103:@30596.4]
  assign _T_83509 = _T_83508[5:0]; // @[Modules.scala 143:103:@30597.4]
  assign _T_83510 = $signed(_T_83509); // @[Modules.scala 143:103:@30598.4]
  assign _T_83515 = $signed(_T_71002) + $signed(_GEN_479); // @[Modules.scala 143:103:@30602.4]
  assign _T_83516 = _T_83515[5:0]; // @[Modules.scala 143:103:@30603.4]
  assign _T_83517 = $signed(_T_83516); // @[Modules.scala 143:103:@30604.4]
  assign _T_83543 = $signed(_T_61818) + $signed(_T_58753); // @[Modules.scala 143:103:@30626.4]
  assign _T_83544 = _T_83543[4:0]; // @[Modules.scala 143:103:@30627.4]
  assign _T_83545 = $signed(_T_83544); // @[Modules.scala 143:103:@30628.4]
  assign _T_83550 = $signed(_T_55746) + $signed(_T_77382); // @[Modules.scala 143:103:@30632.4]
  assign _T_83551 = _T_83550[5:0]; // @[Modules.scala 143:103:@30633.4]
  assign _T_83552 = $signed(_T_83551); // @[Modules.scala 143:103:@30634.4]
  assign _GEN_676 = {{1{_T_58765[4]}},_T_58765}; // @[Modules.scala 143:103:@30638.4]
  assign _T_83557 = $signed(_T_55748) + $signed(_GEN_676); // @[Modules.scala 143:103:@30638.4]
  assign _T_83558 = _T_83557[5:0]; // @[Modules.scala 143:103:@30639.4]
  assign _T_83559 = $signed(_T_83558); // @[Modules.scala 143:103:@30640.4]
  assign _T_83585 = $signed(_T_58788) + $signed(_GEN_64); // @[Modules.scala 143:103:@30662.4]
  assign _T_83586 = _T_83585[5:0]; // @[Modules.scala 143:103:@30663.4]
  assign _T_83587 = $signed(_T_83586); // @[Modules.scala 143:103:@30664.4]
  assign _T_83599 = $signed(_T_58807) + $signed(_T_61879); // @[Modules.scala 143:103:@30674.4]
  assign _T_83600 = _T_83599[4:0]; // @[Modules.scala 143:103:@30675.4]
  assign _T_83601 = $signed(_T_83600); // @[Modules.scala 143:103:@30676.4]
  assign _T_83606 = $signed(_T_55788) + $signed(_GEN_342); // @[Modules.scala 143:103:@30680.4]
  assign _T_83607 = _T_83606[5:0]; // @[Modules.scala 143:103:@30681.4]
  assign _T_83608 = $signed(_T_83607); // @[Modules.scala 143:103:@30682.4]
  assign _GEN_679 = {{1{_T_61907[4]}},_T_61907}; // @[Modules.scala 143:103:@30698.4]
  assign _T_83627 = $signed(_GEN_679) + $signed(_T_55816); // @[Modules.scala 143:103:@30698.4]
  assign _T_83628 = _T_83627[5:0]; // @[Modules.scala 143:103:@30699.4]
  assign _T_83629 = $signed(_T_83628); // @[Modules.scala 143:103:@30700.4]
  assign _T_83634 = $signed(_T_77464) + $signed(_GEN_616); // @[Modules.scala 143:103:@30704.4]
  assign _T_83635 = _T_83634[5:0]; // @[Modules.scala 143:103:@30705.4]
  assign _T_83636 = $signed(_T_83635); // @[Modules.scala 143:103:@30706.4]
  assign _T_83641 = $signed(_GEN_126) + $signed(_T_55825); // @[Modules.scala 143:103:@30710.4]
  assign _T_83642 = _T_83641[5:0]; // @[Modules.scala 143:103:@30711.4]
  assign _T_83643 = $signed(_T_83642); // @[Modules.scala 143:103:@30712.4]
  assign _T_83655 = $signed(_T_74323) + $signed(_T_61937); // @[Modules.scala 143:103:@30722.4]
  assign _T_83656 = _T_83655[5:0]; // @[Modules.scala 143:103:@30723.4]
  assign _T_83657 = $signed(_T_83656); // @[Modules.scala 143:103:@30724.4]
  assign _T_83662 = $signed(_T_74330) + $signed(_T_71179); // @[Modules.scala 143:103:@30728.4]
  assign _T_83663 = _T_83662[5:0]; // @[Modules.scala 143:103:@30729.4]
  assign _T_83664 = $signed(_T_83663); // @[Modules.scala 143:103:@30730.4]
  assign _T_83669 = $signed(_T_55839) + $signed(_GEN_486); // @[Modules.scala 143:103:@30734.4]
  assign _T_83670 = _T_83669[5:0]; // @[Modules.scala 143:103:@30735.4]
  assign _T_83671 = $signed(_T_83670); // @[Modules.scala 143:103:@30736.4]
  assign _T_83676 = $signed(_T_58872) + $signed(_T_58877); // @[Modules.scala 143:103:@30740.4]
  assign _T_83677 = _T_83676[4:0]; // @[Modules.scala 143:103:@30741.4]
  assign _T_83678 = $signed(_T_83677); // @[Modules.scala 143:103:@30742.4]
  assign _T_83697 = $signed(_T_55867) + $signed(_GEN_418); // @[Modules.scala 143:103:@30758.4]
  assign _T_83698 = _T_83697[5:0]; // @[Modules.scala 143:103:@30759.4]
  assign _T_83699 = $signed(_T_83698); // @[Modules.scala 143:103:@30760.4]
  assign _T_83753 = $signed(_T_58949) + $signed(_T_58954); // @[Modules.scala 143:103:@30806.4]
  assign _T_83754 = _T_83753[4:0]; // @[Modules.scala 143:103:@30807.4]
  assign _T_83755 = $signed(_T_83754); // @[Modules.scala 143:103:@30808.4]
  assign _T_83760 = $signed(_GEN_344) + $signed(_T_55949); // @[Modules.scala 143:103:@30812.4]
  assign _T_83761 = _T_83760[5:0]; // @[Modules.scala 143:103:@30813.4]
  assign _T_83762 = $signed(_T_83761); // @[Modules.scala 143:103:@30814.4]
  assign _T_83781 = $signed(_T_55965) + $signed(_T_58982); // @[Modules.scala 143:103:@30830.4]
  assign _T_83782 = _T_83781[5:0]; // @[Modules.scala 143:103:@30831.4]
  assign _T_83783 = $signed(_T_83782); // @[Modules.scala 143:103:@30832.4]
  assign _GEN_686 = {{1{_T_56000[4]}},_T_56000}; // @[Modules.scala 143:103:@30854.4]
  assign _T_83809 = $signed(_GEN_686) + $signed(_T_59005); // @[Modules.scala 143:103:@30854.4]
  assign _T_83810 = _T_83809[5:0]; // @[Modules.scala 143:103:@30855.4]
  assign _T_83811 = $signed(_T_83810); // @[Modules.scala 143:103:@30856.4]
  assign _T_83816 = $signed(_T_62110) + $signed(_GEN_349); // @[Modules.scala 143:103:@30860.4]
  assign _T_83817 = _T_83816[5:0]; // @[Modules.scala 143:103:@30861.4]
  assign _T_83818 = $signed(_T_83817); // @[Modules.scala 143:103:@30862.4]
  assign _T_83837 = $signed(_T_56026) + $signed(_T_56033); // @[Modules.scala 143:103:@30878.4]
  assign _T_83838 = _T_83837[5:0]; // @[Modules.scala 143:103:@30879.4]
  assign _T_83839 = $signed(_T_83838); // @[Modules.scala 143:103:@30880.4]
  assign _T_83858 = $signed(_T_59054) + $signed(_T_59061); // @[Modules.scala 143:103:@30896.4]
  assign _T_83859 = _T_83858[5:0]; // @[Modules.scala 143:103:@30897.4]
  assign _T_83860 = $signed(_T_83859); // @[Modules.scala 143:103:@30898.4]
  assign _T_83865 = $signed(_GEN_206) + $signed(_T_71394); // @[Modules.scala 143:103:@30902.4]
  assign _T_83866 = _T_83865[5:0]; // @[Modules.scala 143:103:@30903.4]
  assign _T_83867 = $signed(_T_83866); // @[Modules.scala 143:103:@30904.4]
  assign _GEN_689 = {{1{_T_56068[4]}},_T_56068}; // @[Modules.scala 143:103:@30908.4]
  assign _T_83872 = $signed(_T_71396) + $signed(_GEN_689); // @[Modules.scala 143:103:@30908.4]
  assign _T_83873 = _T_83872[5:0]; // @[Modules.scala 143:103:@30909.4]
  assign _T_83874 = $signed(_T_83873); // @[Modules.scala 143:103:@30910.4]
  assign _GEN_690 = {{1{_T_56077[4]}},_T_56077}; // @[Modules.scala 143:103:@30920.4]
  assign _T_83886 = $signed(_GEN_690) + $signed(_T_59089); // @[Modules.scala 143:103:@30920.4]
  assign _T_83887 = _T_83886[5:0]; // @[Modules.scala 143:103:@30921.4]
  assign _T_83888 = $signed(_T_83887); // @[Modules.scala 143:103:@30922.4]
  assign _T_83900 = $signed(_T_56091) + $signed(_T_59108); // @[Modules.scala 143:103:@30932.4]
  assign _T_83901 = _T_83900[4:0]; // @[Modules.scala 143:103:@30933.4]
  assign _T_83902 = $signed(_T_83901); // @[Modules.scala 143:103:@30934.4]
  assign _T_83907 = $signed(_GEN_275) + $signed(_T_56105); // @[Modules.scala 143:103:@30938.4]
  assign _T_83908 = _T_83907[5:0]; // @[Modules.scala 143:103:@30939.4]
  assign _T_83909 = $signed(_T_83908); // @[Modules.scala 143:103:@30940.4]
  assign _T_83984 = $signed(_T_65384) + $signed(_T_68423); // @[Modules.scala 143:103:@31004.4]
  assign _T_83985 = _T_83984[5:0]; // @[Modules.scala 143:103:@31005.4]
  assign _T_83986 = $signed(_T_83985); // @[Modules.scala 143:103:@31006.4]
  assign _T_84012 = $signed(_T_62294) + $signed(_T_62299); // @[Modules.scala 143:103:@31028.4]
  assign _T_84013 = _T_84012[4:0]; // @[Modules.scala 143:103:@31029.4]
  assign _T_84014 = $signed(_T_84013); // @[Modules.scala 143:103:@31030.4]
  assign _T_84019 = $signed(_T_62301) + $signed(_T_62306); // @[Modules.scala 143:103:@31034.4]
  assign _T_84020 = _T_84019[4:0]; // @[Modules.scala 143:103:@31035.4]
  assign _T_84021 = $signed(_T_84020); // @[Modules.scala 143:103:@31036.4]
  assign _T_84026 = $signed(_T_62308) + $signed(_T_62313); // @[Modules.scala 143:103:@31040.4]
  assign _T_84027 = _T_84026[4:0]; // @[Modules.scala 143:103:@31041.4]
  assign _T_84028 = $signed(_T_84027); // @[Modules.scala 143:103:@31042.4]
  assign _T_84033 = $signed(_T_56215) + $signed(_T_62320); // @[Modules.scala 143:103:@31046.4]
  assign _T_84034 = _T_84033[4:0]; // @[Modules.scala 143:103:@31047.4]
  assign _T_84035 = $signed(_T_84034); // @[Modules.scala 143:103:@31048.4]
  assign _T_84040 = $signed(_T_62322) + $signed(_T_62327); // @[Modules.scala 143:103:@31052.4]
  assign _T_84041 = _T_84040[4:0]; // @[Modules.scala 143:103:@31053.4]
  assign _T_84042 = $signed(_T_84041); // @[Modules.scala 143:103:@31054.4]
  assign _T_84047 = $signed(_T_56224) + $signed(_T_56229); // @[Modules.scala 143:103:@31058.4]
  assign _T_84048 = _T_84047[4:0]; // @[Modules.scala 143:103:@31059.4]
  assign _T_84049 = $signed(_T_84048); // @[Modules.scala 143:103:@31060.4]
  assign _T_84075 = $signed(_T_59269) + $signed(_T_62362); // @[Modules.scala 143:103:@31082.4]
  assign _T_84076 = _T_84075[4:0]; // @[Modules.scala 143:103:@31083.4]
  assign _T_84077 = $signed(_T_84076); // @[Modules.scala 143:103:@31084.4]
  assign _T_84089 = $signed(_T_62371) + $signed(_T_62376); // @[Modules.scala 143:103:@31094.4]
  assign _T_84090 = _T_84089[4:0]; // @[Modules.scala 143:103:@31095.4]
  assign _T_84091 = $signed(_T_84090); // @[Modules.scala 143:103:@31096.4]
  assign _T_84103 = $signed(_T_62385) + $signed(_T_62390); // @[Modules.scala 143:103:@31106.4]
  assign _T_84104 = _T_84103[4:0]; // @[Modules.scala 143:103:@31107.4]
  assign _T_84105 = $signed(_T_84104); // @[Modules.scala 143:103:@31108.4]
  assign _T_84110 = $signed(_T_62392) + $signed(_T_62397); // @[Modules.scala 143:103:@31112.4]
  assign _T_84111 = _T_84110[4:0]; // @[Modules.scala 143:103:@31113.4]
  assign _T_84112 = $signed(_T_84111); // @[Modules.scala 143:103:@31114.4]
  assign _T_84117 = $signed(_T_62399) + $signed(_T_62404); // @[Modules.scala 143:103:@31118.4]
  assign _T_84118 = _T_84117[4:0]; // @[Modules.scala 143:103:@31119.4]
  assign _T_84119 = $signed(_T_84118); // @[Modules.scala 143:103:@31120.4]
  assign _GEN_693 = {{1{_T_65529[4]}},_T_65529}; // @[Modules.scala 143:103:@31124.4]
  assign _T_84124 = $signed(_T_59318) + $signed(_GEN_693); // @[Modules.scala 143:103:@31124.4]
  assign _T_84125 = _T_84124[5:0]; // @[Modules.scala 143:103:@31125.4]
  assign _T_84126 = $signed(_T_84125); // @[Modules.scala 143:103:@31126.4]
  assign _T_84131 = $signed(_T_59327) + $signed(_T_59332); // @[Modules.scala 143:103:@31130.4]
  assign _T_84132 = _T_84131[4:0]; // @[Modules.scala 143:103:@31131.4]
  assign _T_84133 = $signed(_T_84132); // @[Modules.scala 143:103:@31132.4]
  assign buffer_9_3 = {{8{_T_81963[5]}},_T_81963}; // @[Modules.scala 112:22:@8.4]
  assign _T_84137 = $signed(buffer_2_2) + $signed(buffer_9_3); // @[Modules.scala 160:64:@31138.4]
  assign _T_84138 = _T_84137[13:0]; // @[Modules.scala 160:64:@31139.4]
  assign buffer_9_315 = $signed(_T_84138); // @[Modules.scala 160:64:@31140.4]
  assign buffer_9_6 = {{8{_T_81984[5]}},_T_81984}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_7 = {{8{_T_81991[5]}},_T_81991}; // @[Modules.scala 112:22:@8.4]
  assign _T_84143 = $signed(buffer_9_6) + $signed(buffer_9_7); // @[Modules.scala 160:64:@31146.4]
  assign _T_84144 = _T_84143[13:0]; // @[Modules.scala 160:64:@31147.4]
  assign buffer_9_317 = $signed(_T_84144); // @[Modules.scala 160:64:@31148.4]
  assign buffer_9_8 = {{8{_T_81998[5]}},_T_81998}; // @[Modules.scala 112:22:@8.4]
  assign _T_84146 = $signed(buffer_9_8) + $signed(buffer_4_7); // @[Modules.scala 160:64:@31150.4]
  assign _T_84147 = _T_84146[13:0]; // @[Modules.scala 160:64:@31151.4]
  assign buffer_9_318 = $signed(_T_84147); // @[Modules.scala 160:64:@31152.4]
  assign buffer_9_10 = {{8{_T_82012[5]}},_T_82012}; // @[Modules.scala 112:22:@8.4]
  assign _T_84149 = $signed(buffer_9_10) + $signed(buffer_6_11); // @[Modules.scala 160:64:@31154.4]
  assign _T_84150 = _T_84149[13:0]; // @[Modules.scala 160:64:@31155.4]
  assign buffer_9_319 = $signed(_T_84150); // @[Modules.scala 160:64:@31156.4]
  assign _T_84152 = $signed(buffer_4_10) + $signed(buffer_2_12); // @[Modules.scala 160:64:@31158.4]
  assign _T_84153 = _T_84152[13:0]; // @[Modules.scala 160:64:@31159.4]
  assign buffer_9_320 = $signed(_T_84153); // @[Modules.scala 160:64:@31160.4]
  assign buffer_9_14 = {{8{_T_82040[5]}},_T_82040}; // @[Modules.scala 112:22:@8.4]
  assign _T_84155 = $signed(buffer_9_14) + $signed(buffer_0_14); // @[Modules.scala 160:64:@31162.4]
  assign _T_84156 = _T_84155[13:0]; // @[Modules.scala 160:64:@31163.4]
  assign buffer_9_321 = $signed(_T_84156); // @[Modules.scala 160:64:@31164.4]
  assign _T_84158 = $signed(buffer_0_15) + $signed(buffer_0_16); // @[Modules.scala 160:64:@31166.4]
  assign _T_84159 = _T_84158[13:0]; // @[Modules.scala 160:64:@31167.4]
  assign buffer_9_322 = $signed(_T_84159); // @[Modules.scala 160:64:@31168.4]
  assign _T_84161 = $signed(buffer_0_17) + $signed(buffer_0_18); // @[Modules.scala 160:64:@31170.4]
  assign _T_84162 = _T_84161[13:0]; // @[Modules.scala 160:64:@31171.4]
  assign buffer_9_323 = $signed(_T_84162); // @[Modules.scala 160:64:@31172.4]
  assign _T_84164 = $signed(buffer_0_19) + $signed(buffer_0_20); // @[Modules.scala 160:64:@31174.4]
  assign _T_84165 = _T_84164[13:0]; // @[Modules.scala 160:64:@31175.4]
  assign buffer_9_324 = $signed(_T_84165); // @[Modules.scala 160:64:@31176.4]
  assign buffer_9_22 = {{8{_T_82096[5]}},_T_82096}; // @[Modules.scala 112:22:@8.4]
  assign _T_84167 = $signed(buffer_9_22) + $signed(buffer_3_21); // @[Modules.scala 160:64:@31178.4]
  assign _T_84168 = _T_84167[13:0]; // @[Modules.scala 160:64:@31179.4]
  assign buffer_9_325 = $signed(_T_84168); // @[Modules.scala 160:64:@31180.4]
  assign _T_84170 = $signed(buffer_0_23) + $signed(buffer_0_24); // @[Modules.scala 160:64:@31182.4]
  assign _T_84171 = _T_84170[13:0]; // @[Modules.scala 160:64:@31183.4]
  assign buffer_9_326 = $signed(_T_84171); // @[Modules.scala 160:64:@31184.4]
  assign _T_84173 = $signed(buffer_0_25) + $signed(buffer_1_26); // @[Modules.scala 160:64:@31186.4]
  assign _T_84174 = _T_84173[13:0]; // @[Modules.scala 160:64:@31187.4]
  assign buffer_9_327 = $signed(_T_84174); // @[Modules.scala 160:64:@31188.4]
  assign buffer_9_29 = {{8{_T_82145[5]}},_T_82145}; // @[Modules.scala 112:22:@8.4]
  assign _T_84176 = $signed(buffer_1_27) + $signed(buffer_9_29); // @[Modules.scala 160:64:@31190.4]
  assign _T_84177 = _T_84176[13:0]; // @[Modules.scala 160:64:@31191.4]
  assign buffer_9_328 = $signed(_T_84177); // @[Modules.scala 160:64:@31192.4]
  assign _T_84179 = $signed(buffer_2_27) + $signed(buffer_2_28); // @[Modules.scala 160:64:@31194.4]
  assign _T_84180 = _T_84179[13:0]; // @[Modules.scala 160:64:@31195.4]
  assign buffer_9_329 = $signed(_T_84180); // @[Modules.scala 160:64:@31196.4]
  assign _T_84182 = $signed(buffer_2_29) + $signed(buffer_2_30); // @[Modules.scala 160:64:@31198.4]
  assign _T_84183 = _T_84182[13:0]; // @[Modules.scala 160:64:@31199.4]
  assign buffer_9_330 = $signed(_T_84183); // @[Modules.scala 160:64:@31200.4]
  assign _T_84185 = $signed(buffer_3_32) + $signed(buffer_2_32); // @[Modules.scala 160:64:@31202.4]
  assign _T_84186 = _T_84185[13:0]; // @[Modules.scala 160:64:@31203.4]
  assign buffer_9_331 = $signed(_T_84186); // @[Modules.scala 160:64:@31204.4]
  assign buffer_9_37 = {{8{_T_82201[5]}},_T_82201}; // @[Modules.scala 112:22:@8.4]
  assign _T_84188 = $signed(buffer_1_34) + $signed(buffer_9_37); // @[Modules.scala 160:64:@31206.4]
  assign _T_84189 = _T_84188[13:0]; // @[Modules.scala 160:64:@31207.4]
  assign buffer_9_332 = $signed(_T_84189); // @[Modules.scala 160:64:@31208.4]
  assign buffer_9_38 = {{8{_T_82208[5]}},_T_82208}; // @[Modules.scala 112:22:@8.4]
  assign _T_84191 = $signed(buffer_9_38) + $signed(buffer_3_38); // @[Modules.scala 160:64:@31210.4]
  assign _T_84192 = _T_84191[13:0]; // @[Modules.scala 160:64:@31211.4]
  assign buffer_9_333 = $signed(_T_84192); // @[Modules.scala 160:64:@31212.4]
  assign buffer_9_41 = {{9{_T_82229[4]}},_T_82229}; // @[Modules.scala 112:22:@8.4]
  assign _T_84194 = $signed(buffer_3_39) + $signed(buffer_9_41); // @[Modules.scala 160:64:@31214.4]
  assign _T_84195 = _T_84194[13:0]; // @[Modules.scala 160:64:@31215.4]
  assign buffer_9_334 = $signed(_T_84195); // @[Modules.scala 160:64:@31216.4]
  assign buffer_9_42 = {{8{_T_82236[5]}},_T_82236}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_43 = {{8{_T_82243[5]}},_T_82243}; // @[Modules.scala 112:22:@8.4]
  assign _T_84197 = $signed(buffer_9_42) + $signed(buffer_9_43); // @[Modules.scala 160:64:@31218.4]
  assign _T_84198 = _T_84197[13:0]; // @[Modules.scala 160:64:@31219.4]
  assign buffer_9_335 = $signed(_T_84198); // @[Modules.scala 160:64:@31220.4]
  assign buffer_9_46 = {{8{_T_82264[5]}},_T_82264}; // @[Modules.scala 112:22:@8.4]
  assign _T_84203 = $signed(buffer_9_46) + $signed(buffer_2_43); // @[Modules.scala 160:64:@31226.4]
  assign _T_84204 = _T_84203[13:0]; // @[Modules.scala 160:64:@31227.4]
  assign buffer_9_337 = $signed(_T_84204); // @[Modules.scala 160:64:@31228.4]
  assign _T_84206 = $signed(buffer_6_45) + $signed(buffer_6_46); // @[Modules.scala 160:64:@31230.4]
  assign _T_84207 = _T_84206[13:0]; // @[Modules.scala 160:64:@31231.4]
  assign buffer_9_338 = $signed(_T_84207); // @[Modules.scala 160:64:@31232.4]
  assign buffer_9_51 = {{8{_T_82299[5]}},_T_82299}; // @[Modules.scala 112:22:@8.4]
  assign _T_84209 = $signed(buffer_2_46) + $signed(buffer_9_51); // @[Modules.scala 160:64:@31234.4]
  assign _T_84210 = _T_84209[13:0]; // @[Modules.scala 160:64:@31235.4]
  assign buffer_9_339 = $signed(_T_84210); // @[Modules.scala 160:64:@31236.4]
  assign buffer_9_55 = {{8{_T_82327[5]}},_T_82327}; // @[Modules.scala 112:22:@8.4]
  assign _T_84215 = $signed(buffer_1_51) + $signed(buffer_9_55); // @[Modules.scala 160:64:@31242.4]
  assign _T_84216 = _T_84215[13:0]; // @[Modules.scala 160:64:@31243.4]
  assign buffer_9_341 = $signed(_T_84216); // @[Modules.scala 160:64:@31244.4]
  assign buffer_9_59 = {{8{_T_82355[5]}},_T_82355}; // @[Modules.scala 112:22:@8.4]
  assign _T_84221 = $signed(buffer_3_56) + $signed(buffer_9_59); // @[Modules.scala 160:64:@31250.4]
  assign _T_84222 = _T_84221[13:0]; // @[Modules.scala 160:64:@31251.4]
  assign buffer_9_343 = $signed(_T_84222); // @[Modules.scala 160:64:@31252.4]
  assign buffer_9_60 = {{8{_T_82362[5]}},_T_82362}; // @[Modules.scala 112:22:@8.4]
  assign _T_84224 = $signed(buffer_9_60) + $signed(buffer_0_56); // @[Modules.scala 160:64:@31254.4]
  assign _T_84225 = _T_84224[13:0]; // @[Modules.scala 160:64:@31255.4]
  assign buffer_9_344 = $signed(_T_84225); // @[Modules.scala 160:64:@31256.4]
  assign buffer_9_63 = {{8{_T_82383[5]}},_T_82383}; // @[Modules.scala 112:22:@8.4]
  assign _T_84227 = $signed(buffer_0_57) + $signed(buffer_9_63); // @[Modules.scala 160:64:@31258.4]
  assign _T_84228 = _T_84227[13:0]; // @[Modules.scala 160:64:@31259.4]
  assign buffer_9_345 = $signed(_T_84228); // @[Modules.scala 160:64:@31260.4]
  assign buffer_9_71 = {{8{_T_82439[5]}},_T_82439}; // @[Modules.scala 112:22:@8.4]
  assign _T_84239 = $signed(buffer_7_66) + $signed(buffer_9_71); // @[Modules.scala 160:64:@31274.4]
  assign _T_84240 = _T_84239[13:0]; // @[Modules.scala 160:64:@31275.4]
  assign buffer_9_349 = $signed(_T_84240); // @[Modules.scala 160:64:@31276.4]
  assign buffer_9_73 = {{8{_T_82453[5]}},_T_82453}; // @[Modules.scala 112:22:@8.4]
  assign _T_84242 = $signed(buffer_0_67) + $signed(buffer_9_73); // @[Modules.scala 160:64:@31278.4]
  assign _T_84243 = _T_84242[13:0]; // @[Modules.scala 160:64:@31279.4]
  assign buffer_9_350 = $signed(_T_84243); // @[Modules.scala 160:64:@31280.4]
  assign buffer_9_74 = {{8{_T_82460[5]}},_T_82460}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_75 = {{8{_T_82467[5]}},_T_82467}; // @[Modules.scala 112:22:@8.4]
  assign _T_84245 = $signed(buffer_9_74) + $signed(buffer_9_75); // @[Modules.scala 160:64:@31282.4]
  assign _T_84246 = _T_84245[13:0]; // @[Modules.scala 160:64:@31283.4]
  assign buffer_9_351 = $signed(_T_84246); // @[Modules.scala 160:64:@31284.4]
  assign buffer_9_77 = {{9{_T_82481[4]}},_T_82481}; // @[Modules.scala 112:22:@8.4]
  assign _T_84248 = $signed(buffer_6_73) + $signed(buffer_9_77); // @[Modules.scala 160:64:@31286.4]
  assign _T_84249 = _T_84248[13:0]; // @[Modules.scala 160:64:@31287.4]
  assign buffer_9_352 = $signed(_T_84249); // @[Modules.scala 160:64:@31288.4]
  assign buffer_9_78 = {{8{_T_82488[5]}},_T_82488}; // @[Modules.scala 112:22:@8.4]
  assign _T_84251 = $signed(buffer_9_78) + $signed(buffer_3_79); // @[Modules.scala 160:64:@31290.4]
  assign _T_84252 = _T_84251[13:0]; // @[Modules.scala 160:64:@31291.4]
  assign buffer_9_353 = $signed(_T_84252); // @[Modules.scala 160:64:@31292.4]
  assign _T_84254 = $signed(buffer_3_80) + $signed(buffer_1_79); // @[Modules.scala 160:64:@31294.4]
  assign _T_84255 = _T_84254[13:0]; // @[Modules.scala 160:64:@31295.4]
  assign buffer_9_354 = $signed(_T_84255); // @[Modules.scala 160:64:@31296.4]
  assign buffer_9_84 = {{9{_T_82530[4]}},_T_82530}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_85 = {{9{_T_82537[4]}},_T_82537}; // @[Modules.scala 112:22:@8.4]
  assign _T_84260 = $signed(buffer_9_84) + $signed(buffer_9_85); // @[Modules.scala 160:64:@31302.4]
  assign _T_84261 = _T_84260[13:0]; // @[Modules.scala 160:64:@31303.4]
  assign buffer_9_356 = $signed(_T_84261); // @[Modules.scala 160:64:@31304.4]
  assign buffer_9_86 = {{9{_T_82544[4]}},_T_82544}; // @[Modules.scala 112:22:@8.4]
  assign _T_84263 = $signed(buffer_9_86) + $signed(buffer_2_85); // @[Modules.scala 160:64:@31306.4]
  assign _T_84264 = _T_84263[13:0]; // @[Modules.scala 160:64:@31307.4]
  assign buffer_9_357 = $signed(_T_84264); // @[Modules.scala 160:64:@31308.4]
  assign _T_84266 = $signed(buffer_2_86) + $signed(buffer_0_82); // @[Modules.scala 160:64:@31310.4]
  assign _T_84267 = _T_84266[13:0]; // @[Modules.scala 160:64:@31311.4]
  assign buffer_9_358 = $signed(_T_84267); // @[Modules.scala 160:64:@31312.4]
  assign buffer_9_90 = {{8{_T_82572[5]}},_T_82572}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_91 = {{8{_T_82579[5]}},_T_82579}; // @[Modules.scala 112:22:@8.4]
  assign _T_84269 = $signed(buffer_9_90) + $signed(buffer_9_91); // @[Modules.scala 160:64:@31314.4]
  assign _T_84270 = _T_84269[13:0]; // @[Modules.scala 160:64:@31315.4]
  assign buffer_9_359 = $signed(_T_84270); // @[Modules.scala 160:64:@31316.4]
  assign buffer_9_97 = {{9{_T_82621[4]}},_T_82621}; // @[Modules.scala 112:22:@8.4]
  assign _T_84278 = $signed(buffer_2_94) + $signed(buffer_9_97); // @[Modules.scala 160:64:@31326.4]
  assign _T_84279 = _T_84278[13:0]; // @[Modules.scala 160:64:@31327.4]
  assign buffer_9_362 = $signed(_T_84279); // @[Modules.scala 160:64:@31328.4]
  assign _T_84281 = $signed(buffer_6_96) + $signed(buffer_2_97); // @[Modules.scala 160:64:@31330.4]
  assign _T_84282 = _T_84281[13:0]; // @[Modules.scala 160:64:@31331.4]
  assign buffer_9_363 = $signed(_T_84282); // @[Modules.scala 160:64:@31332.4]
  assign buffer_9_102 = {{9{_T_82656[4]}},_T_82656}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_103 = {{9{_T_82663[4]}},_T_82663}; // @[Modules.scala 112:22:@8.4]
  assign _T_84287 = $signed(buffer_9_102) + $signed(buffer_9_103); // @[Modules.scala 160:64:@31338.4]
  assign _T_84288 = _T_84287[13:0]; // @[Modules.scala 160:64:@31339.4]
  assign buffer_9_365 = $signed(_T_84288); // @[Modules.scala 160:64:@31340.4]
  assign buffer_9_104 = {{9{_T_82670[4]}},_T_82670}; // @[Modules.scala 112:22:@8.4]
  assign _T_84290 = $signed(buffer_9_104) + $signed(buffer_5_105); // @[Modules.scala 160:64:@31342.4]
  assign _T_84291 = _T_84290[13:0]; // @[Modules.scala 160:64:@31343.4]
  assign buffer_9_366 = $signed(_T_84291); // @[Modules.scala 160:64:@31344.4]
  assign buffer_9_107 = {{8{_T_82691[5]}},_T_82691}; // @[Modules.scala 112:22:@8.4]
  assign _T_84293 = $signed(buffer_5_106) + $signed(buffer_9_107); // @[Modules.scala 160:64:@31346.4]
  assign _T_84294 = _T_84293[13:0]; // @[Modules.scala 160:64:@31347.4]
  assign buffer_9_367 = $signed(_T_84294); // @[Modules.scala 160:64:@31348.4]
  assign _T_84296 = $signed(buffer_2_105) + $signed(buffer_2_106); // @[Modules.scala 160:64:@31350.4]
  assign _T_84297 = _T_84296[13:0]; // @[Modules.scala 160:64:@31351.4]
  assign buffer_9_368 = $signed(_T_84297); // @[Modules.scala 160:64:@31352.4]
  assign _T_84299 = $signed(buffer_2_107) + $signed(buffer_1_105); // @[Modules.scala 160:64:@31354.4]
  assign _T_84300 = _T_84299[13:0]; // @[Modules.scala 160:64:@31355.4]
  assign buffer_9_369 = $signed(_T_84300); // @[Modules.scala 160:64:@31356.4]
  assign buffer_9_113 = {{9{_T_82733[4]}},_T_82733}; // @[Modules.scala 112:22:@8.4]
  assign _T_84302 = $signed(buffer_1_106) + $signed(buffer_9_113); // @[Modules.scala 160:64:@31358.4]
  assign _T_84303 = _T_84302[13:0]; // @[Modules.scala 160:64:@31359.4]
  assign buffer_9_370 = $signed(_T_84303); // @[Modules.scala 160:64:@31360.4]
  assign buffer_9_114 = {{8{_T_82740[5]}},_T_82740}; // @[Modules.scala 112:22:@8.4]
  assign _T_84305 = $signed(buffer_9_114) + $signed(buffer_0_108); // @[Modules.scala 160:64:@31362.4]
  assign _T_84306 = _T_84305[13:0]; // @[Modules.scala 160:64:@31363.4]
  assign buffer_9_371 = $signed(_T_84306); // @[Modules.scala 160:64:@31364.4]
  assign _T_84308 = $signed(buffer_0_109) + $signed(buffer_0_110); // @[Modules.scala 160:64:@31366.4]
  assign _T_84309 = _T_84308[13:0]; // @[Modules.scala 160:64:@31367.4]
  assign buffer_9_372 = $signed(_T_84309); // @[Modules.scala 160:64:@31368.4]
  assign _T_84311 = $signed(buffer_3_117) + $signed(buffer_8_110); // @[Modules.scala 160:64:@31370.4]
  assign _T_84312 = _T_84311[13:0]; // @[Modules.scala 160:64:@31371.4]
  assign buffer_9_373 = $signed(_T_84312); // @[Modules.scala 160:64:@31372.4]
  assign buffer_9_120 = {{8{_T_82782[5]}},_T_82782}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_121 = {{9{_T_82789[4]}},_T_82789}; // @[Modules.scala 112:22:@8.4]
  assign _T_84314 = $signed(buffer_9_120) + $signed(buffer_9_121); // @[Modules.scala 160:64:@31374.4]
  assign _T_84315 = _T_84314[13:0]; // @[Modules.scala 160:64:@31375.4]
  assign buffer_9_374 = $signed(_T_84315); // @[Modules.scala 160:64:@31376.4]
  assign buffer_9_123 = {{8{_T_82803[5]}},_T_82803}; // @[Modules.scala 112:22:@8.4]
  assign _T_84317 = $signed(buffer_0_115) + $signed(buffer_9_123); // @[Modules.scala 160:64:@31378.4]
  assign _T_84318 = _T_84317[13:0]; // @[Modules.scala 160:64:@31379.4]
  assign buffer_9_375 = $signed(_T_84318); // @[Modules.scala 160:64:@31380.4]
  assign buffer_9_124 = {{8{_T_82810[5]}},_T_82810}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_125 = {{8{_T_82817[5]}},_T_82817}; // @[Modules.scala 112:22:@8.4]
  assign _T_84320 = $signed(buffer_9_124) + $signed(buffer_9_125); // @[Modules.scala 160:64:@31382.4]
  assign _T_84321 = _T_84320[13:0]; // @[Modules.scala 160:64:@31383.4]
  assign buffer_9_376 = $signed(_T_84321); // @[Modules.scala 160:64:@31384.4]
  assign buffer_9_127 = {{9{_T_82831[4]}},_T_82831}; // @[Modules.scala 112:22:@8.4]
  assign _T_84323 = $signed(buffer_4_118) + $signed(buffer_9_127); // @[Modules.scala 160:64:@31386.4]
  assign _T_84324 = _T_84323[13:0]; // @[Modules.scala 160:64:@31387.4]
  assign buffer_9_377 = $signed(_T_84324); // @[Modules.scala 160:64:@31388.4]
  assign buffer_9_128 = {{9{_T_82838[4]}},_T_82838}; // @[Modules.scala 112:22:@8.4]
  assign _T_84326 = $signed(buffer_9_128) + $signed(buffer_5_125); // @[Modules.scala 160:64:@31390.4]
  assign _T_84327 = _T_84326[13:0]; // @[Modules.scala 160:64:@31391.4]
  assign buffer_9_378 = $signed(_T_84327); // @[Modules.scala 160:64:@31392.4]
  assign _T_84329 = $signed(buffer_1_125) + $signed(buffer_3_131); // @[Modules.scala 160:64:@31394.4]
  assign _T_84330 = _T_84329[13:0]; // @[Modules.scala 160:64:@31395.4]
  assign buffer_9_379 = $signed(_T_84330); // @[Modules.scala 160:64:@31396.4]
  assign _T_84332 = $signed(buffer_1_127) + $signed(buffer_1_128); // @[Modules.scala 160:64:@31398.4]
  assign _T_84333 = _T_84332[13:0]; // @[Modules.scala 160:64:@31399.4]
  assign buffer_9_380 = $signed(_T_84333); // @[Modules.scala 160:64:@31400.4]
  assign buffer_9_134 = {{9{_T_82880[4]}},_T_82880}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_135 = {{8{_T_82887[5]}},_T_82887}; // @[Modules.scala 112:22:@8.4]
  assign _T_84335 = $signed(buffer_9_134) + $signed(buffer_9_135); // @[Modules.scala 160:64:@31402.4]
  assign _T_84336 = _T_84335[13:0]; // @[Modules.scala 160:64:@31403.4]
  assign buffer_9_381 = $signed(_T_84336); // @[Modules.scala 160:64:@31404.4]
  assign buffer_9_140 = {{8{_T_82922[5]}},_T_82922}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_141 = {{9{_T_82929[4]}},_T_82929}; // @[Modules.scala 112:22:@8.4]
  assign _T_84344 = $signed(buffer_9_140) + $signed(buffer_9_141); // @[Modules.scala 160:64:@31414.4]
  assign _T_84345 = _T_84344[13:0]; // @[Modules.scala 160:64:@31415.4]
  assign buffer_9_384 = $signed(_T_84345); // @[Modules.scala 160:64:@31416.4]
  assign buffer_9_142 = {{9{_T_82936[4]}},_T_82936}; // @[Modules.scala 112:22:@8.4]
  assign _T_84347 = $signed(buffer_9_142) + $signed(buffer_0_135); // @[Modules.scala 160:64:@31418.4]
  assign _T_84348 = _T_84347[13:0]; // @[Modules.scala 160:64:@31419.4]
  assign buffer_9_385 = $signed(_T_84348); // @[Modules.scala 160:64:@31420.4]
  assign _T_84350 = $signed(buffer_2_139) + $signed(buffer_2_140); // @[Modules.scala 160:64:@31422.4]
  assign _T_84351 = _T_84350[13:0]; // @[Modules.scala 160:64:@31423.4]
  assign buffer_9_386 = $signed(_T_84351); // @[Modules.scala 160:64:@31424.4]
  assign buffer_9_146 = {{9{_T_82964[4]}},_T_82964}; // @[Modules.scala 112:22:@8.4]
  assign _T_84353 = $signed(buffer_9_146) + $signed(buffer_2_142); // @[Modules.scala 160:64:@31426.4]
  assign _T_84354 = _T_84353[13:0]; // @[Modules.scala 160:64:@31427.4]
  assign buffer_9_387 = $signed(_T_84354); // @[Modules.scala 160:64:@31428.4]
  assign _T_84356 = $signed(buffer_2_143) + $signed(buffer_2_144); // @[Modules.scala 160:64:@31430.4]
  assign _T_84357 = _T_84356[13:0]; // @[Modules.scala 160:64:@31431.4]
  assign buffer_9_388 = $signed(_T_84357); // @[Modules.scala 160:64:@31432.4]
  assign buffer_9_153 = {{8{_T_83013[5]}},_T_83013}; // @[Modules.scala 112:22:@8.4]
  assign _T_84362 = $signed(buffer_2_147) + $signed(buffer_9_153); // @[Modules.scala 160:64:@31438.4]
  assign _T_84363 = _T_84362[13:0]; // @[Modules.scala 160:64:@31439.4]
  assign buffer_9_390 = $signed(_T_84363); // @[Modules.scala 160:64:@31440.4]
  assign buffer_9_154 = {{9{_T_83020[4]}},_T_83020}; // @[Modules.scala 112:22:@8.4]
  assign _T_84365 = $signed(buffer_9_154) + $signed(buffer_3_156); // @[Modules.scala 160:64:@31442.4]
  assign _T_84366 = _T_84365[13:0]; // @[Modules.scala 160:64:@31443.4]
  assign buffer_9_391 = $signed(_T_84366); // @[Modules.scala 160:64:@31444.4]
  assign buffer_9_157 = {{9{_T_83041[4]}},_T_83041}; // @[Modules.scala 112:22:@8.4]
  assign _T_84368 = $signed(buffer_2_153) + $signed(buffer_9_157); // @[Modules.scala 160:64:@31446.4]
  assign _T_84369 = _T_84368[13:0]; // @[Modules.scala 160:64:@31447.4]
  assign buffer_9_392 = $signed(_T_84369); // @[Modules.scala 160:64:@31448.4]
  assign _T_84371 = $signed(buffer_8_150) + $signed(buffer_2_156); // @[Modules.scala 160:64:@31450.4]
  assign _T_84372 = _T_84371[13:0]; // @[Modules.scala 160:64:@31451.4]
  assign buffer_9_393 = $signed(_T_84372); // @[Modules.scala 160:64:@31452.4]
  assign buffer_9_164 = {{8{_T_83090[5]}},_T_83090}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_165 = {{8{_T_83097[5]}},_T_83097}; // @[Modules.scala 112:22:@8.4]
  assign _T_84380 = $signed(buffer_9_164) + $signed(buffer_9_165); // @[Modules.scala 160:64:@31462.4]
  assign _T_84381 = _T_84380[13:0]; // @[Modules.scala 160:64:@31463.4]
  assign buffer_9_396 = $signed(_T_84381); // @[Modules.scala 160:64:@31464.4]
  assign buffer_9_166 = {{8{_T_83104[5]}},_T_83104}; // @[Modules.scala 112:22:@8.4]
  assign _T_84383 = $signed(buffer_9_166) + $signed(buffer_1_162); // @[Modules.scala 160:64:@31466.4]
  assign _T_84384 = _T_84383[13:0]; // @[Modules.scala 160:64:@31467.4]
  assign buffer_9_397 = $signed(_T_84384); // @[Modules.scala 160:64:@31468.4]
  assign buffer_9_168 = {{9{_T_83118[4]}},_T_83118}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_169 = {{8{_T_83125[5]}},_T_83125}; // @[Modules.scala 112:22:@8.4]
  assign _T_84386 = $signed(buffer_9_168) + $signed(buffer_9_169); // @[Modules.scala 160:64:@31470.4]
  assign _T_84387 = _T_84386[13:0]; // @[Modules.scala 160:64:@31471.4]
  assign buffer_9_398 = $signed(_T_84387); // @[Modules.scala 160:64:@31472.4]
  assign _T_84389 = $signed(buffer_1_164) + $signed(buffer_2_169); // @[Modules.scala 160:64:@31474.4]
  assign _T_84390 = _T_84389[13:0]; // @[Modules.scala 160:64:@31475.4]
  assign buffer_9_399 = $signed(_T_84390); // @[Modules.scala 160:64:@31476.4]
  assign buffer_9_172 = {{8{_T_83146[5]}},_T_83146}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_173 = {{8{_T_83153[5]}},_T_83153}; // @[Modules.scala 112:22:@8.4]
  assign _T_84392 = $signed(buffer_9_172) + $signed(buffer_9_173); // @[Modules.scala 160:64:@31478.4]
  assign _T_84393 = _T_84392[13:0]; // @[Modules.scala 160:64:@31479.4]
  assign buffer_9_400 = $signed(_T_84393); // @[Modules.scala 160:64:@31480.4]
  assign buffer_9_175 = {{8{_T_83167[5]}},_T_83167}; // @[Modules.scala 112:22:@8.4]
  assign _T_84395 = $signed(buffer_0_167) + $signed(buffer_9_175); // @[Modules.scala 160:64:@31482.4]
  assign _T_84396 = _T_84395[13:0]; // @[Modules.scala 160:64:@31483.4]
  assign buffer_9_401 = $signed(_T_84396); // @[Modules.scala 160:64:@31484.4]
  assign buffer_9_177 = {{8{_T_83181[5]}},_T_83181}; // @[Modules.scala 112:22:@8.4]
  assign _T_84398 = $signed(buffer_0_170) + $signed(buffer_9_177); // @[Modules.scala 160:64:@31486.4]
  assign _T_84399 = _T_84398[13:0]; // @[Modules.scala 160:64:@31487.4]
  assign buffer_9_402 = $signed(_T_84399); // @[Modules.scala 160:64:@31488.4]
  assign buffer_9_178 = {{8{_T_83188[5]}},_T_83188}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_179 = {{8{_T_83195[5]}},_T_83195}; // @[Modules.scala 112:22:@8.4]
  assign _T_84401 = $signed(buffer_9_178) + $signed(buffer_9_179); // @[Modules.scala 160:64:@31490.4]
  assign _T_84402 = _T_84401[13:0]; // @[Modules.scala 160:64:@31491.4]
  assign buffer_9_403 = $signed(_T_84402); // @[Modules.scala 160:64:@31492.4]
  assign buffer_9_181 = {{8{_T_83209[5]}},_T_83209}; // @[Modules.scala 112:22:@8.4]
  assign _T_84404 = $signed(buffer_3_180) + $signed(buffer_9_181); // @[Modules.scala 160:64:@31494.4]
  assign _T_84405 = _T_84404[13:0]; // @[Modules.scala 160:64:@31495.4]
  assign buffer_9_404 = $signed(_T_84405); // @[Modules.scala 160:64:@31496.4]
  assign buffer_9_182 = {{8{_T_83216[5]}},_T_83216}; // @[Modules.scala 112:22:@8.4]
  assign _T_84407 = $signed(buffer_9_182) + $signed(buffer_1_176); // @[Modules.scala 160:64:@31498.4]
  assign _T_84408 = _T_84407[13:0]; // @[Modules.scala 160:64:@31499.4]
  assign buffer_9_405 = $signed(_T_84408); // @[Modules.scala 160:64:@31500.4]
  assign _T_84410 = $signed(buffer_1_177) + $signed(buffer_1_178); // @[Modules.scala 160:64:@31502.4]
  assign _T_84411 = _T_84410[13:0]; // @[Modules.scala 160:64:@31503.4]
  assign buffer_9_406 = $signed(_T_84411); // @[Modules.scala 160:64:@31504.4]
  assign _T_84413 = $signed(buffer_1_179) + $signed(buffer_0_179); // @[Modules.scala 160:64:@31506.4]
  assign _T_84414 = _T_84413[13:0]; // @[Modules.scala 160:64:@31507.4]
  assign buffer_9_407 = $signed(_T_84414); // @[Modules.scala 160:64:@31508.4]
  assign buffer_9_188 = {{8{_T_83258[5]}},_T_83258}; // @[Modules.scala 112:22:@8.4]
  assign _T_84416 = $signed(buffer_9_188) + $signed(buffer_6_188); // @[Modules.scala 160:64:@31510.4]
  assign _T_84417 = _T_84416[13:0]; // @[Modules.scala 160:64:@31511.4]
  assign buffer_9_408 = $signed(_T_84417); // @[Modules.scala 160:64:@31512.4]
  assign _T_84419 = $signed(buffer_6_189) + $signed(buffer_6_190); // @[Modules.scala 160:64:@31514.4]
  assign _T_84420 = _T_84419[13:0]; // @[Modules.scala 160:64:@31515.4]
  assign buffer_9_409 = $signed(_T_84420); // @[Modules.scala 160:64:@31516.4]
  assign buffer_9_192 = {{9{_T_83286[4]}},_T_83286}; // @[Modules.scala 112:22:@8.4]
  assign _T_84422 = $signed(buffer_9_192) + $signed(buffer_2_190); // @[Modules.scala 160:64:@31518.4]
  assign _T_84423 = _T_84422[13:0]; // @[Modules.scala 160:64:@31519.4]
  assign buffer_9_410 = $signed(_T_84423); // @[Modules.scala 160:64:@31520.4]
  assign buffer_9_200 = {{8{_T_83342[5]}},_T_83342}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_201 = {{8{_T_83349[5]}},_T_83349}; // @[Modules.scala 112:22:@8.4]
  assign _T_84434 = $signed(buffer_9_200) + $signed(buffer_9_201); // @[Modules.scala 160:64:@31534.4]
  assign _T_84435 = _T_84434[13:0]; // @[Modules.scala 160:64:@31535.4]
  assign buffer_9_414 = $signed(_T_84435); // @[Modules.scala 160:64:@31536.4]
  assign buffer_9_202 = {{8{_T_83356[5]}},_T_83356}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_203 = {{8{_T_83363[5]}},_T_83363}; // @[Modules.scala 112:22:@8.4]
  assign _T_84437 = $signed(buffer_9_202) + $signed(buffer_9_203); // @[Modules.scala 160:64:@31538.4]
  assign _T_84438 = _T_84437[13:0]; // @[Modules.scala 160:64:@31539.4]
  assign buffer_9_415 = $signed(_T_84438); // @[Modules.scala 160:64:@31540.4]
  assign buffer_9_205 = {{9{_T_83377[4]}},_T_83377}; // @[Modules.scala 112:22:@8.4]
  assign _T_84440 = $signed(buffer_3_203) + $signed(buffer_9_205); // @[Modules.scala 160:64:@31542.4]
  assign _T_84441 = _T_84440[13:0]; // @[Modules.scala 160:64:@31543.4]
  assign buffer_9_416 = $signed(_T_84441); // @[Modules.scala 160:64:@31544.4]
  assign buffer_9_207 = {{8{_T_83391[5]}},_T_83391}; // @[Modules.scala 112:22:@8.4]
  assign _T_84443 = $signed(buffer_0_195) + $signed(buffer_9_207); // @[Modules.scala 160:64:@31546.4]
  assign _T_84444 = _T_84443[13:0]; // @[Modules.scala 160:64:@31547.4]
  assign buffer_9_417 = $signed(_T_84444); // @[Modules.scala 160:64:@31548.4]
  assign _T_84446 = $signed(buffer_4_191) + $signed(buffer_4_192); // @[Modules.scala 160:64:@31550.4]
  assign _T_84447 = _T_84446[13:0]; // @[Modules.scala 160:64:@31551.4]
  assign buffer_9_418 = $signed(_T_84447); // @[Modules.scala 160:64:@31552.4]
  assign _T_84452 = $signed(buffer_0_201) + $signed(buffer_0_202); // @[Modules.scala 160:64:@31558.4]
  assign _T_84453 = _T_84452[13:0]; // @[Modules.scala 160:64:@31559.4]
  assign buffer_9_420 = $signed(_T_84453); // @[Modules.scala 160:64:@31560.4]
  assign buffer_9_214 = {{8{_T_83440[5]}},_T_83440}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_215 = {{8{_T_83447[5]}},_T_83447}; // @[Modules.scala 112:22:@8.4]
  assign _T_84455 = $signed(buffer_9_214) + $signed(buffer_9_215); // @[Modules.scala 160:64:@31562.4]
  assign _T_84456 = _T_84455[13:0]; // @[Modules.scala 160:64:@31563.4]
  assign buffer_9_421 = $signed(_T_84456); // @[Modules.scala 160:64:@31564.4]
  assign _T_84458 = $signed(buffer_1_205) + $signed(buffer_1_206); // @[Modules.scala 160:64:@31566.4]
  assign _T_84459 = _T_84458[13:0]; // @[Modules.scala 160:64:@31567.4]
  assign buffer_9_422 = $signed(_T_84459); // @[Modules.scala 160:64:@31568.4]
  assign buffer_9_219 = {{8{_T_83475[5]}},_T_83475}; // @[Modules.scala 112:22:@8.4]
  assign _T_84461 = $signed(buffer_2_212) + $signed(buffer_9_219); // @[Modules.scala 160:64:@31570.4]
  assign _T_84462 = _T_84461[13:0]; // @[Modules.scala 160:64:@31571.4]
  assign buffer_9_423 = $signed(_T_84462); // @[Modules.scala 160:64:@31572.4]
  assign buffer_9_223 = {{8{_T_83503[5]}},_T_83503}; // @[Modules.scala 112:22:@8.4]
  assign _T_84467 = $signed(buffer_5_215) + $signed(buffer_9_223); // @[Modules.scala 160:64:@31578.4]
  assign _T_84468 = _T_84467[13:0]; // @[Modules.scala 160:64:@31579.4]
  assign buffer_9_425 = $signed(_T_84468); // @[Modules.scala 160:64:@31580.4]
  assign buffer_9_224 = {{8{_T_83510[5]}},_T_83510}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_225 = {{8{_T_83517[5]}},_T_83517}; // @[Modules.scala 112:22:@8.4]
  assign _T_84470 = $signed(buffer_9_224) + $signed(buffer_9_225); // @[Modules.scala 160:64:@31582.4]
  assign _T_84471 = _T_84470[13:0]; // @[Modules.scala 160:64:@31583.4]
  assign buffer_9_426 = $signed(_T_84471); // @[Modules.scala 160:64:@31584.4]
  assign _T_84473 = $signed(buffer_4_209) + $signed(buffer_8_222); // @[Modules.scala 160:64:@31586.4]
  assign _T_84474 = _T_84473[13:0]; // @[Modules.scala 160:64:@31587.4]
  assign buffer_9_427 = $signed(_T_84474); // @[Modules.scala 160:64:@31588.4]
  assign buffer_9_229 = {{9{_T_83545[4]}},_T_83545}; // @[Modules.scala 112:22:@8.4]
  assign _T_84476 = $signed(buffer_1_219) + $signed(buffer_9_229); // @[Modules.scala 160:64:@31590.4]
  assign _T_84477 = _T_84476[13:0]; // @[Modules.scala 160:64:@31591.4]
  assign buffer_9_428 = $signed(_T_84477); // @[Modules.scala 160:64:@31592.4]
  assign buffer_9_230 = {{8{_T_83552[5]}},_T_83552}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_231 = {{8{_T_83559[5]}},_T_83559}; // @[Modules.scala 112:22:@8.4]
  assign _T_84479 = $signed(buffer_9_230) + $signed(buffer_9_231); // @[Modules.scala 160:64:@31594.4]
  assign _T_84480 = _T_84479[13:0]; // @[Modules.scala 160:64:@31595.4]
  assign buffer_9_429 = $signed(_T_84480); // @[Modules.scala 160:64:@31596.4]
  assign _T_84482 = $signed(buffer_0_223) + $signed(buffer_6_236); // @[Modules.scala 160:64:@31598.4]
  assign _T_84483 = _T_84482[13:0]; // @[Modules.scala 160:64:@31599.4]
  assign buffer_9_430 = $signed(_T_84483); // @[Modules.scala 160:64:@31600.4]
  assign buffer_9_235 = {{8{_T_83587[5]}},_T_83587}; // @[Modules.scala 112:22:@8.4]
  assign _T_84485 = $signed(buffer_5_230) + $signed(buffer_9_235); // @[Modules.scala 160:64:@31602.4]
  assign _T_84486 = _T_84485[13:0]; // @[Modules.scala 160:64:@31603.4]
  assign buffer_9_431 = $signed(_T_84486); // @[Modules.scala 160:64:@31604.4]
  assign buffer_9_237 = {{9{_T_83601[4]}},_T_83601}; // @[Modules.scala 112:22:@8.4]
  assign _T_84488 = $signed(buffer_1_227) + $signed(buffer_9_237); // @[Modules.scala 160:64:@31606.4]
  assign _T_84489 = _T_84488[13:0]; // @[Modules.scala 160:64:@31607.4]
  assign buffer_9_432 = $signed(_T_84489); // @[Modules.scala 160:64:@31608.4]
  assign buffer_9_238 = {{8{_T_83608[5]}},_T_83608}; // @[Modules.scala 112:22:@8.4]
  assign _T_84491 = $signed(buffer_9_238) + $signed(buffer_5_236); // @[Modules.scala 160:64:@31610.4]
  assign _T_84492 = _T_84491[13:0]; // @[Modules.scala 160:64:@31611.4]
  assign buffer_9_433 = $signed(_T_84492); // @[Modules.scala 160:64:@31612.4]
  assign buffer_9_241 = {{8{_T_83629[5]}},_T_83629}; // @[Modules.scala 112:22:@8.4]
  assign _T_84494 = $signed(buffer_2_236) + $signed(buffer_9_241); // @[Modules.scala 160:64:@31614.4]
  assign _T_84495 = _T_84494[13:0]; // @[Modules.scala 160:64:@31615.4]
  assign buffer_9_434 = $signed(_T_84495); // @[Modules.scala 160:64:@31616.4]
  assign buffer_9_242 = {{8{_T_83636[5]}},_T_83636}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_243 = {{8{_T_83643[5]}},_T_83643}; // @[Modules.scala 112:22:@8.4]
  assign _T_84497 = $signed(buffer_9_242) + $signed(buffer_9_243); // @[Modules.scala 160:64:@31618.4]
  assign _T_84498 = _T_84497[13:0]; // @[Modules.scala 160:64:@31619.4]
  assign buffer_9_435 = $signed(_T_84498); // @[Modules.scala 160:64:@31620.4]
  assign buffer_9_245 = {{8{_T_83657[5]}},_T_83657}; // @[Modules.scala 112:22:@8.4]
  assign _T_84500 = $signed(buffer_0_233) + $signed(buffer_9_245); // @[Modules.scala 160:64:@31622.4]
  assign _T_84501 = _T_84500[13:0]; // @[Modules.scala 160:64:@31623.4]
  assign buffer_9_436 = $signed(_T_84501); // @[Modules.scala 160:64:@31624.4]
  assign buffer_9_246 = {{8{_T_83664[5]}},_T_83664}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_247 = {{8{_T_83671[5]}},_T_83671}; // @[Modules.scala 112:22:@8.4]
  assign _T_84503 = $signed(buffer_9_246) + $signed(buffer_9_247); // @[Modules.scala 160:64:@31626.4]
  assign _T_84504 = _T_84503[13:0]; // @[Modules.scala 160:64:@31627.4]
  assign buffer_9_437 = $signed(_T_84504); // @[Modules.scala 160:64:@31628.4]
  assign buffer_9_248 = {{9{_T_83678[4]}},_T_83678}; // @[Modules.scala 112:22:@8.4]
  assign _T_84506 = $signed(buffer_9_248) + $signed(buffer_5_247); // @[Modules.scala 160:64:@31630.4]
  assign _T_84507 = _T_84506[13:0]; // @[Modules.scala 160:64:@31631.4]
  assign buffer_9_438 = $signed(_T_84507); // @[Modules.scala 160:64:@31632.4]
  assign buffer_9_251 = {{8{_T_83699[5]}},_T_83699}; // @[Modules.scala 112:22:@8.4]
  assign _T_84509 = $signed(buffer_6_250) + $signed(buffer_9_251); // @[Modules.scala 160:64:@31634.4]
  assign _T_84510 = _T_84509[13:0]; // @[Modules.scala 160:64:@31635.4]
  assign buffer_9_439 = $signed(_T_84510); // @[Modules.scala 160:64:@31636.4]
  assign _T_84512 = $signed(buffer_2_249) + $signed(buffer_3_252); // @[Modules.scala 160:64:@31638.4]
  assign _T_84513 = _T_84512[13:0]; // @[Modules.scala 160:64:@31639.4]
  assign buffer_9_440 = $signed(_T_84513); // @[Modules.scala 160:64:@31640.4]
  assign _T_84518 = $signed(buffer_3_255) + $signed(buffer_3_256); // @[Modules.scala 160:64:@31646.4]
  assign _T_84519 = _T_84518[13:0]; // @[Modules.scala 160:64:@31647.4]
  assign buffer_9_442 = $signed(_T_84519); // @[Modules.scala 160:64:@31648.4]
  assign buffer_9_259 = {{9{_T_83755[4]}},_T_83755}; // @[Modules.scala 112:22:@8.4]
  assign _T_84521 = $signed(buffer_6_258) + $signed(buffer_9_259); // @[Modules.scala 160:64:@31650.4]
  assign _T_84522 = _T_84521[13:0]; // @[Modules.scala 160:64:@31651.4]
  assign buffer_9_443 = $signed(_T_84522); // @[Modules.scala 160:64:@31652.4]
  assign buffer_9_260 = {{8{_T_83762[5]}},_T_83762}; // @[Modules.scala 112:22:@8.4]
  assign _T_84524 = $signed(buffer_9_260) + $signed(buffer_5_259); // @[Modules.scala 160:64:@31654.4]
  assign _T_84525 = _T_84524[13:0]; // @[Modules.scala 160:64:@31655.4]
  assign buffer_9_444 = $signed(_T_84525); // @[Modules.scala 160:64:@31656.4]
  assign buffer_9_263 = {{8{_T_83783[5]}},_T_83783}; // @[Modules.scala 112:22:@8.4]
  assign _T_84527 = $signed(buffer_6_263) + $signed(buffer_9_263); // @[Modules.scala 160:64:@31658.4]
  assign _T_84528 = _T_84527[13:0]; // @[Modules.scala 160:64:@31659.4]
  assign buffer_9_445 = $signed(_T_84528); // @[Modules.scala 160:64:@31660.4]
  assign _T_84530 = $signed(buffer_4_249) + $signed(buffer_0_255); // @[Modules.scala 160:64:@31662.4]
  assign _T_84531 = _T_84530[13:0]; // @[Modules.scala 160:64:@31663.4]
  assign buffer_9_446 = $signed(_T_84531); // @[Modules.scala 160:64:@31664.4]
  assign buffer_9_267 = {{8{_T_83811[5]}},_T_83811}; // @[Modules.scala 112:22:@8.4]
  assign _T_84533 = $signed(buffer_0_256) + $signed(buffer_9_267); // @[Modules.scala 160:64:@31666.4]
  assign _T_84534 = _T_84533[13:0]; // @[Modules.scala 160:64:@31667.4]
  assign buffer_9_447 = $signed(_T_84534); // @[Modules.scala 160:64:@31668.4]
  assign buffer_9_268 = {{8{_T_83818[5]}},_T_83818}; // @[Modules.scala 112:22:@8.4]
  assign _T_84536 = $signed(buffer_9_268) + $signed(buffer_1_258); // @[Modules.scala 160:64:@31670.4]
  assign _T_84537 = _T_84536[13:0]; // @[Modules.scala 160:64:@31671.4]
  assign buffer_9_448 = $signed(_T_84537); // @[Modules.scala 160:64:@31672.4]
  assign buffer_9_271 = {{8{_T_83839[5]}},_T_83839}; // @[Modules.scala 112:22:@8.4]
  assign _T_84539 = $signed(buffer_2_268) + $signed(buffer_9_271); // @[Modules.scala 160:64:@31674.4]
  assign _T_84540 = _T_84539[13:0]; // @[Modules.scala 160:64:@31675.4]
  assign buffer_9_449 = $signed(_T_84540); // @[Modules.scala 160:64:@31676.4]
  assign _T_84542 = $signed(buffer_6_273) + $signed(buffer_6_274); // @[Modules.scala 160:64:@31678.4]
  assign _T_84543 = _T_84542[13:0]; // @[Modules.scala 160:64:@31679.4]
  assign buffer_9_450 = $signed(_T_84543); // @[Modules.scala 160:64:@31680.4]
  assign buffer_9_274 = {{8{_T_83860[5]}},_T_83860}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_275 = {{8{_T_83867[5]}},_T_83867}; // @[Modules.scala 112:22:@8.4]
  assign _T_84545 = $signed(buffer_9_274) + $signed(buffer_9_275); // @[Modules.scala 160:64:@31682.4]
  assign _T_84546 = _T_84545[13:0]; // @[Modules.scala 160:64:@31683.4]
  assign buffer_9_451 = $signed(_T_84546); // @[Modules.scala 160:64:@31684.4]
  assign buffer_9_276 = {{8{_T_83874[5]}},_T_83874}; // @[Modules.scala 112:22:@8.4]
  assign _T_84548 = $signed(buffer_9_276) + $signed(buffer_6_278); // @[Modules.scala 160:64:@31686.4]
  assign _T_84549 = _T_84548[13:0]; // @[Modules.scala 160:64:@31687.4]
  assign buffer_9_452 = $signed(_T_84549); // @[Modules.scala 160:64:@31688.4]
  assign buffer_9_278 = {{8{_T_83888[5]}},_T_83888}; // @[Modules.scala 112:22:@8.4]
  assign _T_84551 = $signed(buffer_9_278) + $signed(buffer_6_280); // @[Modules.scala 160:64:@31690.4]
  assign _T_84552 = _T_84551[13:0]; // @[Modules.scala 160:64:@31691.4]
  assign buffer_9_453 = $signed(_T_84552); // @[Modules.scala 160:64:@31692.4]
  assign buffer_9_280 = {{9{_T_83902[4]}},_T_83902}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_281 = {{8{_T_83909[5]}},_T_83909}; // @[Modules.scala 112:22:@8.4]
  assign _T_84554 = $signed(buffer_9_280) + $signed(buffer_9_281); // @[Modules.scala 160:64:@31694.4]
  assign _T_84555 = _T_84554[13:0]; // @[Modules.scala 160:64:@31695.4]
  assign buffer_9_454 = $signed(_T_84555); // @[Modules.scala 160:64:@31696.4]
  assign _T_84569 = $signed(buffer_6_291) + $signed(buffer_6_292); // @[Modules.scala 160:64:@31714.4]
  assign _T_84570 = _T_84569[13:0]; // @[Modules.scala 160:64:@31715.4]
  assign buffer_9_459 = $signed(_T_84570); // @[Modules.scala 160:64:@31716.4]
  assign buffer_9_292 = {{8{_T_83986[5]}},_T_83986}; // @[Modules.scala 112:22:@8.4]
  assign _T_84572 = $signed(buffer_9_292) + $signed(buffer_0_284); // @[Modules.scala 160:64:@31718.4]
  assign _T_84573 = _T_84572[13:0]; // @[Modules.scala 160:64:@31719.4]
  assign buffer_9_460 = $signed(_T_84573); // @[Modules.scala 160:64:@31720.4]
  assign buffer_9_296 = {{9{_T_84014[4]}},_T_84014}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_297 = {{9{_T_84021[4]}},_T_84021}; // @[Modules.scala 112:22:@8.4]
  assign _T_84578 = $signed(buffer_9_296) + $signed(buffer_9_297); // @[Modules.scala 160:64:@31726.4]
  assign _T_84579 = _T_84578[13:0]; // @[Modules.scala 160:64:@31727.4]
  assign buffer_9_462 = $signed(_T_84579); // @[Modules.scala 160:64:@31728.4]
  assign buffer_9_298 = {{9{_T_84028[4]}},_T_84028}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_299 = {{9{_T_84035[4]}},_T_84035}; // @[Modules.scala 112:22:@8.4]
  assign _T_84581 = $signed(buffer_9_298) + $signed(buffer_9_299); // @[Modules.scala 160:64:@31730.4]
  assign _T_84582 = _T_84581[13:0]; // @[Modules.scala 160:64:@31731.4]
  assign buffer_9_463 = $signed(_T_84582); // @[Modules.scala 160:64:@31732.4]
  assign buffer_9_300 = {{9{_T_84042[4]}},_T_84042}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_301 = {{9{_T_84049[4]}},_T_84049}; // @[Modules.scala 112:22:@8.4]
  assign _T_84584 = $signed(buffer_9_300) + $signed(buffer_9_301); // @[Modules.scala 160:64:@31734.4]
  assign _T_84585 = _T_84584[13:0]; // @[Modules.scala 160:64:@31735.4]
  assign buffer_9_464 = $signed(_T_84585); // @[Modules.scala 160:64:@31736.4]
  assign _T_84587 = $signed(buffer_6_304) + $signed(buffer_2_299); // @[Modules.scala 160:64:@31738.4]
  assign _T_84588 = _T_84587[13:0]; // @[Modules.scala 160:64:@31739.4]
  assign buffer_9_465 = $signed(_T_84588); // @[Modules.scala 160:64:@31740.4]
  assign buffer_9_305 = {{9{_T_84077[4]}},_T_84077}; // @[Modules.scala 112:22:@8.4]
  assign _T_84590 = $signed(buffer_2_300) + $signed(buffer_9_305); // @[Modules.scala 160:64:@31742.4]
  assign _T_84591 = _T_84590[13:0]; // @[Modules.scala 160:64:@31743.4]
  assign buffer_9_466 = $signed(_T_84591); // @[Modules.scala 160:64:@31744.4]
  assign buffer_9_307 = {{9{_T_84091[4]}},_T_84091}; // @[Modules.scala 112:22:@8.4]
  assign _T_84593 = $signed(buffer_0_294) + $signed(buffer_9_307); // @[Modules.scala 160:64:@31746.4]
  assign _T_84594 = _T_84593[13:0]; // @[Modules.scala 160:64:@31747.4]
  assign buffer_9_467 = $signed(_T_84594); // @[Modules.scala 160:64:@31748.4]
  assign buffer_9_309 = {{9{_T_84105[4]}},_T_84105}; // @[Modules.scala 112:22:@8.4]
  assign _T_84596 = $signed(buffer_1_297) + $signed(buffer_9_309); // @[Modules.scala 160:64:@31750.4]
  assign _T_84597 = _T_84596[13:0]; // @[Modules.scala 160:64:@31751.4]
  assign buffer_9_468 = $signed(_T_84597); // @[Modules.scala 160:64:@31752.4]
  assign buffer_9_310 = {{9{_T_84112[4]}},_T_84112}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_311 = {{9{_T_84119[4]}},_T_84119}; // @[Modules.scala 112:22:@8.4]
  assign _T_84599 = $signed(buffer_9_310) + $signed(buffer_9_311); // @[Modules.scala 160:64:@31754.4]
  assign _T_84600 = _T_84599[13:0]; // @[Modules.scala 160:64:@31755.4]
  assign buffer_9_469 = $signed(_T_84600); // @[Modules.scala 160:64:@31756.4]
  assign buffer_9_312 = {{8{_T_84126[5]}},_T_84126}; // @[Modules.scala 112:22:@8.4]
  assign buffer_9_313 = {{9{_T_84133[4]}},_T_84133}; // @[Modules.scala 112:22:@8.4]
  assign _T_84602 = $signed(buffer_9_312) + $signed(buffer_9_313); // @[Modules.scala 160:64:@31758.4]
  assign _T_84603 = _T_84602[13:0]; // @[Modules.scala 160:64:@31759.4]
  assign buffer_9_470 = $signed(_T_84603); // @[Modules.scala 160:64:@31760.4]
  assign _T_84605 = $signed(buffer_2_310) + $signed(buffer_9_315); // @[Modules.scala 166:64:@31762.4]
  assign _T_84606 = _T_84605[13:0]; // @[Modules.scala 166:64:@31763.4]
  assign buffer_9_471 = $signed(_T_84606); // @[Modules.scala 166:64:@31764.4]
  assign _T_84608 = $signed(buffer_2_312) + $signed(buffer_9_317); // @[Modules.scala 166:64:@31766.4]
  assign _T_84609 = _T_84608[13:0]; // @[Modules.scala 166:64:@31767.4]
  assign buffer_9_472 = $signed(_T_84609); // @[Modules.scala 166:64:@31768.4]
  assign _T_84611 = $signed(buffer_9_318) + $signed(buffer_9_319); // @[Modules.scala 166:64:@31770.4]
  assign _T_84612 = _T_84611[13:0]; // @[Modules.scala 166:64:@31771.4]
  assign buffer_9_473 = $signed(_T_84612); // @[Modules.scala 166:64:@31772.4]
  assign _T_84614 = $signed(buffer_9_320) + $signed(buffer_9_321); // @[Modules.scala 166:64:@31774.4]
  assign _T_84615 = _T_84614[13:0]; // @[Modules.scala 166:64:@31775.4]
  assign buffer_9_474 = $signed(_T_84615); // @[Modules.scala 166:64:@31776.4]
  assign _T_84617 = $signed(buffer_9_322) + $signed(buffer_9_323); // @[Modules.scala 166:64:@31778.4]
  assign _T_84618 = _T_84617[13:0]; // @[Modules.scala 166:64:@31779.4]
  assign buffer_9_475 = $signed(_T_84618); // @[Modules.scala 166:64:@31780.4]
  assign _T_84620 = $signed(buffer_9_324) + $signed(buffer_9_325); // @[Modules.scala 166:64:@31782.4]
  assign _T_84621 = _T_84620[13:0]; // @[Modules.scala 166:64:@31783.4]
  assign buffer_9_476 = $signed(_T_84621); // @[Modules.scala 166:64:@31784.4]
  assign _T_84623 = $signed(buffer_9_326) + $signed(buffer_9_327); // @[Modules.scala 166:64:@31786.4]
  assign _T_84624 = _T_84623[13:0]; // @[Modules.scala 166:64:@31787.4]
  assign buffer_9_477 = $signed(_T_84624); // @[Modules.scala 166:64:@31788.4]
  assign _T_84626 = $signed(buffer_9_328) + $signed(buffer_9_329); // @[Modules.scala 166:64:@31790.4]
  assign _T_84627 = _T_84626[13:0]; // @[Modules.scala 166:64:@31791.4]
  assign buffer_9_478 = $signed(_T_84627); // @[Modules.scala 166:64:@31792.4]
  assign _T_84629 = $signed(buffer_9_330) + $signed(buffer_9_331); // @[Modules.scala 166:64:@31794.4]
  assign _T_84630 = _T_84629[13:0]; // @[Modules.scala 166:64:@31795.4]
  assign buffer_9_479 = $signed(_T_84630); // @[Modules.scala 166:64:@31796.4]
  assign _T_84632 = $signed(buffer_9_332) + $signed(buffer_9_333); // @[Modules.scala 166:64:@31798.4]
  assign _T_84633 = _T_84632[13:0]; // @[Modules.scala 166:64:@31799.4]
  assign buffer_9_480 = $signed(_T_84633); // @[Modules.scala 166:64:@31800.4]
  assign _T_84635 = $signed(buffer_9_334) + $signed(buffer_9_335); // @[Modules.scala 166:64:@31802.4]
  assign _T_84636 = _T_84635[13:0]; // @[Modules.scala 166:64:@31803.4]
  assign buffer_9_481 = $signed(_T_84636); // @[Modules.scala 166:64:@31804.4]
  assign _T_84638 = $signed(buffer_3_335) + $signed(buffer_9_337); // @[Modules.scala 166:64:@31806.4]
  assign _T_84639 = _T_84638[13:0]; // @[Modules.scala 166:64:@31807.4]
  assign buffer_9_482 = $signed(_T_84639); // @[Modules.scala 166:64:@31808.4]
  assign _T_84641 = $signed(buffer_9_338) + $signed(buffer_9_339); // @[Modules.scala 166:64:@31810.4]
  assign _T_84642 = _T_84641[13:0]; // @[Modules.scala 166:64:@31811.4]
  assign buffer_9_483 = $signed(_T_84642); // @[Modules.scala 166:64:@31812.4]
  assign _T_84644 = $signed(buffer_2_334) + $signed(buffer_9_341); // @[Modules.scala 166:64:@31814.4]
  assign _T_84645 = _T_84644[13:0]; // @[Modules.scala 166:64:@31815.4]
  assign buffer_9_484 = $signed(_T_84645); // @[Modules.scala 166:64:@31816.4]
  assign _T_84647 = $signed(buffer_3_341) + $signed(buffer_9_343); // @[Modules.scala 166:64:@31818.4]
  assign _T_84648 = _T_84647[13:0]; // @[Modules.scala 166:64:@31819.4]
  assign buffer_9_485 = $signed(_T_84648); // @[Modules.scala 166:64:@31820.4]
  assign _T_84650 = $signed(buffer_9_344) + $signed(buffer_9_345); // @[Modules.scala 166:64:@31822.4]
  assign _T_84651 = _T_84650[13:0]; // @[Modules.scala 166:64:@31823.4]
  assign buffer_9_486 = $signed(_T_84651); // @[Modules.scala 166:64:@31824.4]
  assign _T_84656 = $signed(buffer_7_341) + $signed(buffer_9_349); // @[Modules.scala 166:64:@31830.4]
  assign _T_84657 = _T_84656[13:0]; // @[Modules.scala 166:64:@31831.4]
  assign buffer_9_488 = $signed(_T_84657); // @[Modules.scala 166:64:@31832.4]
  assign _T_84659 = $signed(buffer_9_350) + $signed(buffer_9_351); // @[Modules.scala 166:64:@31834.4]
  assign _T_84660 = _T_84659[13:0]; // @[Modules.scala 166:64:@31835.4]
  assign buffer_9_489 = $signed(_T_84660); // @[Modules.scala 166:64:@31836.4]
  assign _T_84662 = $signed(buffer_9_352) + $signed(buffer_9_353); // @[Modules.scala 166:64:@31838.4]
  assign _T_84663 = _T_84662[13:0]; // @[Modules.scala 166:64:@31839.4]
  assign buffer_9_490 = $signed(_T_84663); // @[Modules.scala 166:64:@31840.4]
  assign _T_84665 = $signed(buffer_9_354) + $signed(buffer_2_350); // @[Modules.scala 166:64:@31842.4]
  assign _T_84666 = _T_84665[13:0]; // @[Modules.scala 166:64:@31843.4]
  assign buffer_9_491 = $signed(_T_84666); // @[Modules.scala 166:64:@31844.4]
  assign _T_84668 = $signed(buffer_9_356) + $signed(buffer_9_357); // @[Modules.scala 166:64:@31846.4]
  assign _T_84669 = _T_84668[13:0]; // @[Modules.scala 166:64:@31847.4]
  assign buffer_9_492 = $signed(_T_84669); // @[Modules.scala 166:64:@31848.4]
  assign _T_84671 = $signed(buffer_9_358) + $signed(buffer_9_359); // @[Modules.scala 166:64:@31850.4]
  assign _T_84672 = _T_84671[13:0]; // @[Modules.scala 166:64:@31851.4]
  assign buffer_9_493 = $signed(_T_84672); // @[Modules.scala 166:64:@31852.4]
  assign _T_84674 = $signed(buffer_8_351) + $signed(buffer_2_356); // @[Modules.scala 166:64:@31854.4]
  assign _T_84675 = _T_84674[13:0]; // @[Modules.scala 166:64:@31855.4]
  assign buffer_9_494 = $signed(_T_84675); // @[Modules.scala 166:64:@31856.4]
  assign _T_84677 = $signed(buffer_9_362) + $signed(buffer_9_363); // @[Modules.scala 166:64:@31858.4]
  assign _T_84678 = _T_84677[13:0]; // @[Modules.scala 166:64:@31859.4]
  assign buffer_9_495 = $signed(_T_84678); // @[Modules.scala 166:64:@31860.4]
  assign _T_84680 = $signed(buffer_2_359) + $signed(buffer_9_365); // @[Modules.scala 166:64:@31862.4]
  assign _T_84681 = _T_84680[13:0]; // @[Modules.scala 166:64:@31863.4]
  assign buffer_9_496 = $signed(_T_84681); // @[Modules.scala 166:64:@31864.4]
  assign _T_84683 = $signed(buffer_9_366) + $signed(buffer_9_367); // @[Modules.scala 166:64:@31866.4]
  assign _T_84684 = _T_84683[13:0]; // @[Modules.scala 166:64:@31867.4]
  assign buffer_9_497 = $signed(_T_84684); // @[Modules.scala 166:64:@31868.4]
  assign _T_84686 = $signed(buffer_9_368) + $signed(buffer_9_369); // @[Modules.scala 166:64:@31870.4]
  assign _T_84687 = _T_84686[13:0]; // @[Modules.scala 166:64:@31871.4]
  assign buffer_9_498 = $signed(_T_84687); // @[Modules.scala 166:64:@31872.4]
  assign _T_84689 = $signed(buffer_9_370) + $signed(buffer_9_371); // @[Modules.scala 166:64:@31874.4]
  assign _T_84690 = _T_84689[13:0]; // @[Modules.scala 166:64:@31875.4]
  assign buffer_9_499 = $signed(_T_84690); // @[Modules.scala 166:64:@31876.4]
  assign _T_84692 = $signed(buffer_9_372) + $signed(buffer_9_373); // @[Modules.scala 166:64:@31878.4]
  assign _T_84693 = _T_84692[13:0]; // @[Modules.scala 166:64:@31879.4]
  assign buffer_9_500 = $signed(_T_84693); // @[Modules.scala 166:64:@31880.4]
  assign _T_84695 = $signed(buffer_9_374) + $signed(buffer_9_375); // @[Modules.scala 166:64:@31882.4]
  assign _T_84696 = _T_84695[13:0]; // @[Modules.scala 166:64:@31883.4]
  assign buffer_9_501 = $signed(_T_84696); // @[Modules.scala 166:64:@31884.4]
  assign _T_84698 = $signed(buffer_9_376) + $signed(buffer_9_377); // @[Modules.scala 166:64:@31886.4]
  assign _T_84699 = _T_84698[13:0]; // @[Modules.scala 166:64:@31887.4]
  assign buffer_9_502 = $signed(_T_84699); // @[Modules.scala 166:64:@31888.4]
  assign _T_84701 = $signed(buffer_9_378) + $signed(buffer_9_379); // @[Modules.scala 166:64:@31890.4]
  assign _T_84702 = _T_84701[13:0]; // @[Modules.scala 166:64:@31891.4]
  assign buffer_9_503 = $signed(_T_84702); // @[Modules.scala 166:64:@31892.4]
  assign _T_84704 = $signed(buffer_9_380) + $signed(buffer_9_381); // @[Modules.scala 166:64:@31894.4]
  assign _T_84705 = _T_84704[13:0]; // @[Modules.scala 166:64:@31895.4]
  assign buffer_9_504 = $signed(_T_84705); // @[Modules.scala 166:64:@31896.4]
  assign _T_84710 = $signed(buffer_9_384) + $signed(buffer_9_385); // @[Modules.scala 166:64:@31902.4]
  assign _T_84711 = _T_84710[13:0]; // @[Modules.scala 166:64:@31903.4]
  assign buffer_9_506 = $signed(_T_84711); // @[Modules.scala 166:64:@31904.4]
  assign _T_84713 = $signed(buffer_9_386) + $signed(buffer_9_387); // @[Modules.scala 166:64:@31906.4]
  assign _T_84714 = _T_84713[13:0]; // @[Modules.scala 166:64:@31907.4]
  assign buffer_9_507 = $signed(_T_84714); // @[Modules.scala 166:64:@31908.4]
  assign _T_84716 = $signed(buffer_9_388) + $signed(buffer_8_379); // @[Modules.scala 166:64:@31910.4]
  assign _T_84717 = _T_84716[13:0]; // @[Modules.scala 166:64:@31911.4]
  assign buffer_9_508 = $signed(_T_84717); // @[Modules.scala 166:64:@31912.4]
  assign _T_84719 = $signed(buffer_9_390) + $signed(buffer_9_391); // @[Modules.scala 166:64:@31914.4]
  assign _T_84720 = _T_84719[13:0]; // @[Modules.scala 166:64:@31915.4]
  assign buffer_9_509 = $signed(_T_84720); // @[Modules.scala 166:64:@31916.4]
  assign _T_84722 = $signed(buffer_9_392) + $signed(buffer_9_393); // @[Modules.scala 166:64:@31918.4]
  assign _T_84723 = _T_84722[13:0]; // @[Modules.scala 166:64:@31919.4]
  assign buffer_9_510 = $signed(_T_84723); // @[Modules.scala 166:64:@31920.4]
  assign _T_84728 = $signed(buffer_9_396) + $signed(buffer_9_397); // @[Modules.scala 166:64:@31926.4]
  assign _T_84729 = _T_84728[13:0]; // @[Modules.scala 166:64:@31927.4]
  assign buffer_9_512 = $signed(_T_84729); // @[Modules.scala 166:64:@31928.4]
  assign _T_84731 = $signed(buffer_9_398) + $signed(buffer_9_399); // @[Modules.scala 166:64:@31930.4]
  assign _T_84732 = _T_84731[13:0]; // @[Modules.scala 166:64:@31931.4]
  assign buffer_9_513 = $signed(_T_84732); // @[Modules.scala 166:64:@31932.4]
  assign _T_84734 = $signed(buffer_9_400) + $signed(buffer_9_401); // @[Modules.scala 166:64:@31934.4]
  assign _T_84735 = _T_84734[13:0]; // @[Modules.scala 166:64:@31935.4]
  assign buffer_9_514 = $signed(_T_84735); // @[Modules.scala 166:64:@31936.4]
  assign _T_84737 = $signed(buffer_9_402) + $signed(buffer_9_403); // @[Modules.scala 166:64:@31938.4]
  assign _T_84738 = _T_84737[13:0]; // @[Modules.scala 166:64:@31939.4]
  assign buffer_9_515 = $signed(_T_84738); // @[Modules.scala 166:64:@31940.4]
  assign _T_84740 = $signed(buffer_9_404) + $signed(buffer_9_405); // @[Modules.scala 166:64:@31942.4]
  assign _T_84741 = _T_84740[13:0]; // @[Modules.scala 166:64:@31943.4]
  assign buffer_9_516 = $signed(_T_84741); // @[Modules.scala 166:64:@31944.4]
  assign _T_84743 = $signed(buffer_9_406) + $signed(buffer_9_407); // @[Modules.scala 166:64:@31946.4]
  assign _T_84744 = _T_84743[13:0]; // @[Modules.scala 166:64:@31947.4]
  assign buffer_9_517 = $signed(_T_84744); // @[Modules.scala 166:64:@31948.4]
  assign _T_84746 = $signed(buffer_9_408) + $signed(buffer_9_409); // @[Modules.scala 166:64:@31950.4]
  assign _T_84747 = _T_84746[13:0]; // @[Modules.scala 166:64:@31951.4]
  assign buffer_9_518 = $signed(_T_84747); // @[Modules.scala 166:64:@31952.4]
  assign _T_84749 = $signed(buffer_9_410) + $signed(buffer_8_402); // @[Modules.scala 166:64:@31954.4]
  assign _T_84750 = _T_84749[13:0]; // @[Modules.scala 166:64:@31955.4]
  assign buffer_9_519 = $signed(_T_84750); // @[Modules.scala 166:64:@31956.4]
  assign _T_84755 = $signed(buffer_9_414) + $signed(buffer_9_415); // @[Modules.scala 166:64:@31962.4]
  assign _T_84756 = _T_84755[13:0]; // @[Modules.scala 166:64:@31963.4]
  assign buffer_9_521 = $signed(_T_84756); // @[Modules.scala 166:64:@31964.4]
  assign _T_84758 = $signed(buffer_9_416) + $signed(buffer_9_417); // @[Modules.scala 166:64:@31966.4]
  assign _T_84759 = _T_84758[13:0]; // @[Modules.scala 166:64:@31967.4]
  assign buffer_9_522 = $signed(_T_84759); // @[Modules.scala 166:64:@31968.4]
  assign _T_84761 = $signed(buffer_9_418) + $signed(buffer_8_410); // @[Modules.scala 166:64:@31970.4]
  assign _T_84762 = _T_84761[13:0]; // @[Modules.scala 166:64:@31971.4]
  assign buffer_9_523 = $signed(_T_84762); // @[Modules.scala 166:64:@31972.4]
  assign _T_84764 = $signed(buffer_9_420) + $signed(buffer_9_421); // @[Modules.scala 166:64:@31974.4]
  assign _T_84765 = _T_84764[13:0]; // @[Modules.scala 166:64:@31975.4]
  assign buffer_9_524 = $signed(_T_84765); // @[Modules.scala 166:64:@31976.4]
  assign _T_84767 = $signed(buffer_9_422) + $signed(buffer_9_423); // @[Modules.scala 166:64:@31978.4]
  assign _T_84768 = _T_84767[13:0]; // @[Modules.scala 166:64:@31979.4]
  assign buffer_9_525 = $signed(_T_84768); // @[Modules.scala 166:64:@31980.4]
  assign _T_84770 = $signed(buffer_4_401) + $signed(buffer_9_425); // @[Modules.scala 166:64:@31982.4]
  assign _T_84771 = _T_84770[13:0]; // @[Modules.scala 166:64:@31983.4]
  assign buffer_9_526 = $signed(_T_84771); // @[Modules.scala 166:64:@31984.4]
  assign _T_84773 = $signed(buffer_9_426) + $signed(buffer_9_427); // @[Modules.scala 166:64:@31986.4]
  assign _T_84774 = _T_84773[13:0]; // @[Modules.scala 166:64:@31987.4]
  assign buffer_9_527 = $signed(_T_84774); // @[Modules.scala 166:64:@31988.4]
  assign _T_84776 = $signed(buffer_9_428) + $signed(buffer_9_429); // @[Modules.scala 166:64:@31990.4]
  assign _T_84777 = _T_84776[13:0]; // @[Modules.scala 166:64:@31991.4]
  assign buffer_9_528 = $signed(_T_84777); // @[Modules.scala 166:64:@31992.4]
  assign _T_84779 = $signed(buffer_9_430) + $signed(buffer_9_431); // @[Modules.scala 166:64:@31994.4]
  assign _T_84780 = _T_84779[13:0]; // @[Modules.scala 166:64:@31995.4]
  assign buffer_9_529 = $signed(_T_84780); // @[Modules.scala 166:64:@31996.4]
  assign _T_84782 = $signed(buffer_9_432) + $signed(buffer_9_433); // @[Modules.scala 166:64:@31998.4]
  assign _T_84783 = _T_84782[13:0]; // @[Modules.scala 166:64:@31999.4]
  assign buffer_9_530 = $signed(_T_84783); // @[Modules.scala 166:64:@32000.4]
  assign _T_84785 = $signed(buffer_9_434) + $signed(buffer_9_435); // @[Modules.scala 166:64:@32002.4]
  assign _T_84786 = _T_84785[13:0]; // @[Modules.scala 166:64:@32003.4]
  assign buffer_9_531 = $signed(_T_84786); // @[Modules.scala 166:64:@32004.4]
  assign _T_84788 = $signed(buffer_9_436) + $signed(buffer_9_437); // @[Modules.scala 166:64:@32006.4]
  assign _T_84789 = _T_84788[13:0]; // @[Modules.scala 166:64:@32007.4]
  assign buffer_9_532 = $signed(_T_84789); // @[Modules.scala 166:64:@32008.4]
  assign _T_84791 = $signed(buffer_9_438) + $signed(buffer_9_439); // @[Modules.scala 166:64:@32010.4]
  assign _T_84792 = _T_84791[13:0]; // @[Modules.scala 166:64:@32011.4]
  assign buffer_9_533 = $signed(_T_84792); // @[Modules.scala 166:64:@32012.4]
  assign _T_84794 = $signed(buffer_9_440) + $signed(buffer_0_423); // @[Modules.scala 166:64:@32014.4]
  assign _T_84795 = _T_84794[13:0]; // @[Modules.scala 166:64:@32015.4]
  assign buffer_9_534 = $signed(_T_84795); // @[Modules.scala 166:64:@32016.4]
  assign _T_84797 = $signed(buffer_9_442) + $signed(buffer_9_443); // @[Modules.scala 166:64:@32018.4]
  assign _T_84798 = _T_84797[13:0]; // @[Modules.scala 166:64:@32019.4]
  assign buffer_9_535 = $signed(_T_84798); // @[Modules.scala 166:64:@32020.4]
  assign _T_84800 = $signed(buffer_9_444) + $signed(buffer_9_445); // @[Modules.scala 166:64:@32022.4]
  assign _T_84801 = _T_84800[13:0]; // @[Modules.scala 166:64:@32023.4]
  assign buffer_9_536 = $signed(_T_84801); // @[Modules.scala 166:64:@32024.4]
  assign _T_84803 = $signed(buffer_9_446) + $signed(buffer_9_447); // @[Modules.scala 166:64:@32026.4]
  assign _T_84804 = _T_84803[13:0]; // @[Modules.scala 166:64:@32027.4]
  assign buffer_9_537 = $signed(_T_84804); // @[Modules.scala 166:64:@32028.4]
  assign _T_84806 = $signed(buffer_9_448) + $signed(buffer_9_449); // @[Modules.scala 166:64:@32030.4]
  assign _T_84807 = _T_84806[13:0]; // @[Modules.scala 166:64:@32031.4]
  assign buffer_9_538 = $signed(_T_84807); // @[Modules.scala 166:64:@32032.4]
  assign _T_84809 = $signed(buffer_9_450) + $signed(buffer_9_451); // @[Modules.scala 166:64:@32034.4]
  assign _T_84810 = _T_84809[13:0]; // @[Modules.scala 166:64:@32035.4]
  assign buffer_9_539 = $signed(_T_84810); // @[Modules.scala 166:64:@32036.4]
  assign _T_84812 = $signed(buffer_9_452) + $signed(buffer_9_453); // @[Modules.scala 166:64:@32038.4]
  assign _T_84813 = _T_84812[13:0]; // @[Modules.scala 166:64:@32039.4]
  assign buffer_9_540 = $signed(_T_84813); // @[Modules.scala 166:64:@32040.4]
  assign _T_84815 = $signed(buffer_9_454) + $signed(buffer_3_455); // @[Modules.scala 166:64:@32042.4]
  assign _T_84816 = _T_84815[13:0]; // @[Modules.scala 166:64:@32043.4]
  assign buffer_9_541 = $signed(_T_84816); // @[Modules.scala 166:64:@32044.4]
  assign _T_84821 = $signed(buffer_2_452) + $signed(buffer_9_459); // @[Modules.scala 166:64:@32050.4]
  assign _T_84822 = _T_84821[13:0]; // @[Modules.scala 166:64:@32051.4]
  assign buffer_9_543 = $signed(_T_84822); // @[Modules.scala 166:64:@32052.4]
  assign _T_84824 = $signed(buffer_9_460) + $signed(buffer_7_454); // @[Modules.scala 166:64:@32054.4]
  assign _T_84825 = _T_84824[13:0]; // @[Modules.scala 166:64:@32055.4]
  assign buffer_9_544 = $signed(_T_84825); // @[Modules.scala 166:64:@32056.4]
  assign _T_84827 = $signed(buffer_9_462) + $signed(buffer_9_463); // @[Modules.scala 166:64:@32058.4]
  assign _T_84828 = _T_84827[13:0]; // @[Modules.scala 166:64:@32059.4]
  assign buffer_9_545 = $signed(_T_84828); // @[Modules.scala 166:64:@32060.4]
  assign _T_84830 = $signed(buffer_9_464) + $signed(buffer_9_465); // @[Modules.scala 166:64:@32062.4]
  assign _T_84831 = _T_84830[13:0]; // @[Modules.scala 166:64:@32063.4]
  assign buffer_9_546 = $signed(_T_84831); // @[Modules.scala 166:64:@32064.4]
  assign _T_84833 = $signed(buffer_9_466) + $signed(buffer_9_467); // @[Modules.scala 166:64:@32066.4]
  assign _T_84834 = _T_84833[13:0]; // @[Modules.scala 166:64:@32067.4]
  assign buffer_9_547 = $signed(_T_84834); // @[Modules.scala 166:64:@32068.4]
  assign _T_84836 = $signed(buffer_9_468) + $signed(buffer_9_469); // @[Modules.scala 166:64:@32070.4]
  assign _T_84837 = _T_84836[13:0]; // @[Modules.scala 166:64:@32071.4]
  assign buffer_9_548 = $signed(_T_84837); // @[Modules.scala 166:64:@32072.4]
  assign _T_84839 = $signed(buffer_9_471) + $signed(buffer_9_472); // @[Modules.scala 160:64:@32074.4]
  assign _T_84840 = _T_84839[13:0]; // @[Modules.scala 160:64:@32075.4]
  assign buffer_9_549 = $signed(_T_84840); // @[Modules.scala 160:64:@32076.4]
  assign _T_84842 = $signed(buffer_9_473) + $signed(buffer_9_474); // @[Modules.scala 160:64:@32078.4]
  assign _T_84843 = _T_84842[13:0]; // @[Modules.scala 160:64:@32079.4]
  assign buffer_9_550 = $signed(_T_84843); // @[Modules.scala 160:64:@32080.4]
  assign _T_84845 = $signed(buffer_9_475) + $signed(buffer_9_476); // @[Modules.scala 160:64:@32082.4]
  assign _T_84846 = _T_84845[13:0]; // @[Modules.scala 160:64:@32083.4]
  assign buffer_9_551 = $signed(_T_84846); // @[Modules.scala 160:64:@32084.4]
  assign _T_84848 = $signed(buffer_9_477) + $signed(buffer_9_478); // @[Modules.scala 160:64:@32086.4]
  assign _T_84849 = _T_84848[13:0]; // @[Modules.scala 160:64:@32087.4]
  assign buffer_9_552 = $signed(_T_84849); // @[Modules.scala 160:64:@32088.4]
  assign _T_84851 = $signed(buffer_9_479) + $signed(buffer_9_480); // @[Modules.scala 160:64:@32090.4]
  assign _T_84852 = _T_84851[13:0]; // @[Modules.scala 160:64:@32091.4]
  assign buffer_9_553 = $signed(_T_84852); // @[Modules.scala 160:64:@32092.4]
  assign _T_84854 = $signed(buffer_9_481) + $signed(buffer_9_482); // @[Modules.scala 160:64:@32094.4]
  assign _T_84855 = _T_84854[13:0]; // @[Modules.scala 160:64:@32095.4]
  assign buffer_9_554 = $signed(_T_84855); // @[Modules.scala 160:64:@32096.4]
  assign _T_84857 = $signed(buffer_9_483) + $signed(buffer_9_484); // @[Modules.scala 160:64:@32098.4]
  assign _T_84858 = _T_84857[13:0]; // @[Modules.scala 160:64:@32099.4]
  assign buffer_9_555 = $signed(_T_84858); // @[Modules.scala 160:64:@32100.4]
  assign _T_84860 = $signed(buffer_9_485) + $signed(buffer_9_486); // @[Modules.scala 160:64:@32102.4]
  assign _T_84861 = _T_84860[13:0]; // @[Modules.scala 160:64:@32103.4]
  assign buffer_9_556 = $signed(_T_84861); // @[Modules.scala 160:64:@32104.4]
  assign _T_84863 = $signed(buffer_7_478) + $signed(buffer_9_488); // @[Modules.scala 160:64:@32106.4]
  assign _T_84864 = _T_84863[13:0]; // @[Modules.scala 160:64:@32107.4]
  assign buffer_9_557 = $signed(_T_84864); // @[Modules.scala 160:64:@32108.4]
  assign _T_84866 = $signed(buffer_9_489) + $signed(buffer_9_490); // @[Modules.scala 160:64:@32110.4]
  assign _T_84867 = _T_84866[13:0]; // @[Modules.scala 160:64:@32111.4]
  assign buffer_9_558 = $signed(_T_84867); // @[Modules.scala 160:64:@32112.4]
  assign _T_84869 = $signed(buffer_9_491) + $signed(buffer_9_492); // @[Modules.scala 160:64:@32114.4]
  assign _T_84870 = _T_84869[13:0]; // @[Modules.scala 160:64:@32115.4]
  assign buffer_9_559 = $signed(_T_84870); // @[Modules.scala 160:64:@32116.4]
  assign _T_84872 = $signed(buffer_9_493) + $signed(buffer_9_494); // @[Modules.scala 160:64:@32118.4]
  assign _T_84873 = _T_84872[13:0]; // @[Modules.scala 160:64:@32119.4]
  assign buffer_9_560 = $signed(_T_84873); // @[Modules.scala 160:64:@32120.4]
  assign _T_84875 = $signed(buffer_9_495) + $signed(buffer_9_496); // @[Modules.scala 160:64:@32122.4]
  assign _T_84876 = _T_84875[13:0]; // @[Modules.scala 160:64:@32123.4]
  assign buffer_9_561 = $signed(_T_84876); // @[Modules.scala 160:64:@32124.4]
  assign _T_84878 = $signed(buffer_9_497) + $signed(buffer_9_498); // @[Modules.scala 160:64:@32126.4]
  assign _T_84879 = _T_84878[13:0]; // @[Modules.scala 160:64:@32127.4]
  assign buffer_9_562 = $signed(_T_84879); // @[Modules.scala 160:64:@32128.4]
  assign _T_84881 = $signed(buffer_9_499) + $signed(buffer_9_500); // @[Modules.scala 160:64:@32130.4]
  assign _T_84882 = _T_84881[13:0]; // @[Modules.scala 160:64:@32131.4]
  assign buffer_9_563 = $signed(_T_84882); // @[Modules.scala 160:64:@32132.4]
  assign _T_84884 = $signed(buffer_9_501) + $signed(buffer_9_502); // @[Modules.scala 160:64:@32134.4]
  assign _T_84885 = _T_84884[13:0]; // @[Modules.scala 160:64:@32135.4]
  assign buffer_9_564 = $signed(_T_84885); // @[Modules.scala 160:64:@32136.4]
  assign _T_84887 = $signed(buffer_9_503) + $signed(buffer_9_504); // @[Modules.scala 160:64:@32138.4]
  assign _T_84888 = _T_84887[13:0]; // @[Modules.scala 160:64:@32139.4]
  assign buffer_9_565 = $signed(_T_84888); // @[Modules.scala 160:64:@32140.4]
  assign _T_84890 = $signed(buffer_3_505) + $signed(buffer_9_506); // @[Modules.scala 160:64:@32142.4]
  assign _T_84891 = _T_84890[13:0]; // @[Modules.scala 160:64:@32143.4]
  assign buffer_9_566 = $signed(_T_84891); // @[Modules.scala 160:64:@32144.4]
  assign _T_84893 = $signed(buffer_9_507) + $signed(buffer_9_508); // @[Modules.scala 160:64:@32146.4]
  assign _T_84894 = _T_84893[13:0]; // @[Modules.scala 160:64:@32147.4]
  assign buffer_9_567 = $signed(_T_84894); // @[Modules.scala 160:64:@32148.4]
  assign _T_84896 = $signed(buffer_9_509) + $signed(buffer_9_510); // @[Modules.scala 160:64:@32150.4]
  assign _T_84897 = _T_84896[13:0]; // @[Modules.scala 160:64:@32151.4]
  assign buffer_9_568 = $signed(_T_84897); // @[Modules.scala 160:64:@32152.4]
  assign _T_84899 = $signed(buffer_3_511) + $signed(buffer_9_512); // @[Modules.scala 160:64:@32154.4]
  assign _T_84900 = _T_84899[13:0]; // @[Modules.scala 160:64:@32155.4]
  assign buffer_9_569 = $signed(_T_84900); // @[Modules.scala 160:64:@32156.4]
  assign _T_84902 = $signed(buffer_9_513) + $signed(buffer_9_514); // @[Modules.scala 160:64:@32158.4]
  assign _T_84903 = _T_84902[13:0]; // @[Modules.scala 160:64:@32159.4]
  assign buffer_9_570 = $signed(_T_84903); // @[Modules.scala 160:64:@32160.4]
  assign _T_84905 = $signed(buffer_9_515) + $signed(buffer_9_516); // @[Modules.scala 160:64:@32162.4]
  assign _T_84906 = _T_84905[13:0]; // @[Modules.scala 160:64:@32163.4]
  assign buffer_9_571 = $signed(_T_84906); // @[Modules.scala 160:64:@32164.4]
  assign _T_84908 = $signed(buffer_9_517) + $signed(buffer_9_518); // @[Modules.scala 160:64:@32166.4]
  assign _T_84909 = _T_84908[13:0]; // @[Modules.scala 160:64:@32167.4]
  assign buffer_9_572 = $signed(_T_84909); // @[Modules.scala 160:64:@32168.4]
  assign _T_84911 = $signed(buffer_9_519) + $signed(buffer_8_510); // @[Modules.scala 160:64:@32170.4]
  assign _T_84912 = _T_84911[13:0]; // @[Modules.scala 160:64:@32171.4]
  assign buffer_9_573 = $signed(_T_84912); // @[Modules.scala 160:64:@32172.4]
  assign _T_84914 = $signed(buffer_9_521) + $signed(buffer_9_522); // @[Modules.scala 160:64:@32174.4]
  assign _T_84915 = _T_84914[13:0]; // @[Modules.scala 160:64:@32175.4]
  assign buffer_9_574 = $signed(_T_84915); // @[Modules.scala 160:64:@32176.4]
  assign _T_84917 = $signed(buffer_9_523) + $signed(buffer_9_524); // @[Modules.scala 160:64:@32178.4]
  assign _T_84918 = _T_84917[13:0]; // @[Modules.scala 160:64:@32179.4]
  assign buffer_9_575 = $signed(_T_84918); // @[Modules.scala 160:64:@32180.4]
  assign _T_84920 = $signed(buffer_9_525) + $signed(buffer_9_526); // @[Modules.scala 160:64:@32182.4]
  assign _T_84921 = _T_84920[13:0]; // @[Modules.scala 160:64:@32183.4]
  assign buffer_9_576 = $signed(_T_84921); // @[Modules.scala 160:64:@32184.4]
  assign _T_84923 = $signed(buffer_9_527) + $signed(buffer_9_528); // @[Modules.scala 160:64:@32186.4]
  assign _T_84924 = _T_84923[13:0]; // @[Modules.scala 160:64:@32187.4]
  assign buffer_9_577 = $signed(_T_84924); // @[Modules.scala 160:64:@32188.4]
  assign _T_84926 = $signed(buffer_9_529) + $signed(buffer_9_530); // @[Modules.scala 160:64:@32190.4]
  assign _T_84927 = _T_84926[13:0]; // @[Modules.scala 160:64:@32191.4]
  assign buffer_9_578 = $signed(_T_84927); // @[Modules.scala 160:64:@32192.4]
  assign _T_84929 = $signed(buffer_9_531) + $signed(buffer_9_532); // @[Modules.scala 160:64:@32194.4]
  assign _T_84930 = _T_84929[13:0]; // @[Modules.scala 160:64:@32195.4]
  assign buffer_9_579 = $signed(_T_84930); // @[Modules.scala 160:64:@32196.4]
  assign _T_84932 = $signed(buffer_9_533) + $signed(buffer_9_534); // @[Modules.scala 160:64:@32198.4]
  assign _T_84933 = _T_84932[13:0]; // @[Modules.scala 160:64:@32199.4]
  assign buffer_9_580 = $signed(_T_84933); // @[Modules.scala 160:64:@32200.4]
  assign _T_84935 = $signed(buffer_9_535) + $signed(buffer_9_536); // @[Modules.scala 160:64:@32202.4]
  assign _T_84936 = _T_84935[13:0]; // @[Modules.scala 160:64:@32203.4]
  assign buffer_9_581 = $signed(_T_84936); // @[Modules.scala 160:64:@32204.4]
  assign _T_84938 = $signed(buffer_9_537) + $signed(buffer_9_538); // @[Modules.scala 160:64:@32206.4]
  assign _T_84939 = _T_84938[13:0]; // @[Modules.scala 160:64:@32207.4]
  assign buffer_9_582 = $signed(_T_84939); // @[Modules.scala 160:64:@32208.4]
  assign _T_84941 = $signed(buffer_9_539) + $signed(buffer_9_540); // @[Modules.scala 160:64:@32210.4]
  assign _T_84942 = _T_84941[13:0]; // @[Modules.scala 160:64:@32211.4]
  assign buffer_9_583 = $signed(_T_84942); // @[Modules.scala 160:64:@32212.4]
  assign _T_84944 = $signed(buffer_9_541) + $signed(buffer_3_542); // @[Modules.scala 160:64:@32214.4]
  assign _T_84945 = _T_84944[13:0]; // @[Modules.scala 160:64:@32215.4]
  assign buffer_9_584 = $signed(_T_84945); // @[Modules.scala 160:64:@32216.4]
  assign _T_84947 = $signed(buffer_9_543) + $signed(buffer_9_544); // @[Modules.scala 160:64:@32218.4]
  assign _T_84948 = _T_84947[13:0]; // @[Modules.scala 160:64:@32219.4]
  assign buffer_9_585 = $signed(_T_84948); // @[Modules.scala 160:64:@32220.4]
  assign _T_84950 = $signed(buffer_9_545) + $signed(buffer_9_546); // @[Modules.scala 160:64:@32222.4]
  assign _T_84951 = _T_84950[13:0]; // @[Modules.scala 160:64:@32223.4]
  assign buffer_9_586 = $signed(_T_84951); // @[Modules.scala 160:64:@32224.4]
  assign _T_84953 = $signed(buffer_9_547) + $signed(buffer_9_548); // @[Modules.scala 160:64:@32226.4]
  assign _T_84954 = _T_84953[13:0]; // @[Modules.scala 160:64:@32227.4]
  assign buffer_9_587 = $signed(_T_84954); // @[Modules.scala 160:64:@32228.4]
  assign _T_84956 = $signed(buffer_9_549) + $signed(buffer_9_550); // @[Modules.scala 166:64:@32230.4]
  assign _T_84957 = _T_84956[13:0]; // @[Modules.scala 166:64:@32231.4]
  assign buffer_9_588 = $signed(_T_84957); // @[Modules.scala 166:64:@32232.4]
  assign _T_84959 = $signed(buffer_9_551) + $signed(buffer_9_552); // @[Modules.scala 166:64:@32234.4]
  assign _T_84960 = _T_84959[13:0]; // @[Modules.scala 166:64:@32235.4]
  assign buffer_9_589 = $signed(_T_84960); // @[Modules.scala 166:64:@32236.4]
  assign _T_84962 = $signed(buffer_9_553) + $signed(buffer_9_554); // @[Modules.scala 166:64:@32238.4]
  assign _T_84963 = _T_84962[13:0]; // @[Modules.scala 166:64:@32239.4]
  assign buffer_9_590 = $signed(_T_84963); // @[Modules.scala 166:64:@32240.4]
  assign _T_84965 = $signed(buffer_9_555) + $signed(buffer_9_556); // @[Modules.scala 166:64:@32242.4]
  assign _T_84966 = _T_84965[13:0]; // @[Modules.scala 166:64:@32243.4]
  assign buffer_9_591 = $signed(_T_84966); // @[Modules.scala 166:64:@32244.4]
  assign _T_84968 = $signed(buffer_9_557) + $signed(buffer_9_558); // @[Modules.scala 166:64:@32246.4]
  assign _T_84969 = _T_84968[13:0]; // @[Modules.scala 166:64:@32247.4]
  assign buffer_9_592 = $signed(_T_84969); // @[Modules.scala 166:64:@32248.4]
  assign _T_84971 = $signed(buffer_9_559) + $signed(buffer_9_560); // @[Modules.scala 166:64:@32250.4]
  assign _T_84972 = _T_84971[13:0]; // @[Modules.scala 166:64:@32251.4]
  assign buffer_9_593 = $signed(_T_84972); // @[Modules.scala 166:64:@32252.4]
  assign _T_84974 = $signed(buffer_9_561) + $signed(buffer_9_562); // @[Modules.scala 166:64:@32254.4]
  assign _T_84975 = _T_84974[13:0]; // @[Modules.scala 166:64:@32255.4]
  assign buffer_9_594 = $signed(_T_84975); // @[Modules.scala 166:64:@32256.4]
  assign _T_84977 = $signed(buffer_9_563) + $signed(buffer_9_564); // @[Modules.scala 166:64:@32258.4]
  assign _T_84978 = _T_84977[13:0]; // @[Modules.scala 166:64:@32259.4]
  assign buffer_9_595 = $signed(_T_84978); // @[Modules.scala 166:64:@32260.4]
  assign _T_84980 = $signed(buffer_9_565) + $signed(buffer_9_566); // @[Modules.scala 166:64:@32262.4]
  assign _T_84981 = _T_84980[13:0]; // @[Modules.scala 166:64:@32263.4]
  assign buffer_9_596 = $signed(_T_84981); // @[Modules.scala 166:64:@32264.4]
  assign _T_84983 = $signed(buffer_9_567) + $signed(buffer_9_568); // @[Modules.scala 166:64:@32266.4]
  assign _T_84984 = _T_84983[13:0]; // @[Modules.scala 166:64:@32267.4]
  assign buffer_9_597 = $signed(_T_84984); // @[Modules.scala 166:64:@32268.4]
  assign _T_84986 = $signed(buffer_9_569) + $signed(buffer_9_570); // @[Modules.scala 166:64:@32270.4]
  assign _T_84987 = _T_84986[13:0]; // @[Modules.scala 166:64:@32271.4]
  assign buffer_9_598 = $signed(_T_84987); // @[Modules.scala 166:64:@32272.4]
  assign _T_84989 = $signed(buffer_9_571) + $signed(buffer_9_572); // @[Modules.scala 166:64:@32274.4]
  assign _T_84990 = _T_84989[13:0]; // @[Modules.scala 166:64:@32275.4]
  assign buffer_9_599 = $signed(_T_84990); // @[Modules.scala 166:64:@32276.4]
  assign _T_84992 = $signed(buffer_9_573) + $signed(buffer_9_574); // @[Modules.scala 166:64:@32278.4]
  assign _T_84993 = _T_84992[13:0]; // @[Modules.scala 166:64:@32279.4]
  assign buffer_9_600 = $signed(_T_84993); // @[Modules.scala 166:64:@32280.4]
  assign _T_84995 = $signed(buffer_9_575) + $signed(buffer_9_576); // @[Modules.scala 166:64:@32282.4]
  assign _T_84996 = _T_84995[13:0]; // @[Modules.scala 166:64:@32283.4]
  assign buffer_9_601 = $signed(_T_84996); // @[Modules.scala 166:64:@32284.4]
  assign _T_84998 = $signed(buffer_9_577) + $signed(buffer_9_578); // @[Modules.scala 166:64:@32286.4]
  assign _T_84999 = _T_84998[13:0]; // @[Modules.scala 166:64:@32287.4]
  assign buffer_9_602 = $signed(_T_84999); // @[Modules.scala 166:64:@32288.4]
  assign _T_85001 = $signed(buffer_9_579) + $signed(buffer_9_580); // @[Modules.scala 166:64:@32290.4]
  assign _T_85002 = _T_85001[13:0]; // @[Modules.scala 166:64:@32291.4]
  assign buffer_9_603 = $signed(_T_85002); // @[Modules.scala 166:64:@32292.4]
  assign _T_85004 = $signed(buffer_9_581) + $signed(buffer_9_582); // @[Modules.scala 166:64:@32294.4]
  assign _T_85005 = _T_85004[13:0]; // @[Modules.scala 166:64:@32295.4]
  assign buffer_9_604 = $signed(_T_85005); // @[Modules.scala 166:64:@32296.4]
  assign _T_85007 = $signed(buffer_9_583) + $signed(buffer_9_584); // @[Modules.scala 166:64:@32298.4]
  assign _T_85008 = _T_85007[13:0]; // @[Modules.scala 166:64:@32299.4]
  assign buffer_9_605 = $signed(_T_85008); // @[Modules.scala 166:64:@32300.4]
  assign _T_85010 = $signed(buffer_9_585) + $signed(buffer_9_586); // @[Modules.scala 166:64:@32302.4]
  assign _T_85011 = _T_85010[13:0]; // @[Modules.scala 166:64:@32303.4]
  assign buffer_9_606 = $signed(_T_85011); // @[Modules.scala 166:64:@32304.4]
  assign _T_85013 = $signed(buffer_9_587) + $signed(buffer_9_470); // @[Modules.scala 172:66:@32306.4]
  assign _T_85014 = _T_85013[13:0]; // @[Modules.scala 172:66:@32307.4]
  assign buffer_9_607 = $signed(_T_85014); // @[Modules.scala 172:66:@32308.4]
  assign _T_85016 = $signed(buffer_9_588) + $signed(buffer_9_589); // @[Modules.scala 160:64:@32310.4]
  assign _T_85017 = _T_85016[13:0]; // @[Modules.scala 160:64:@32311.4]
  assign buffer_9_608 = $signed(_T_85017); // @[Modules.scala 160:64:@32312.4]
  assign _T_85019 = $signed(buffer_9_590) + $signed(buffer_9_591); // @[Modules.scala 160:64:@32314.4]
  assign _T_85020 = _T_85019[13:0]; // @[Modules.scala 160:64:@32315.4]
  assign buffer_9_609 = $signed(_T_85020); // @[Modules.scala 160:64:@32316.4]
  assign _T_85022 = $signed(buffer_9_592) + $signed(buffer_9_593); // @[Modules.scala 160:64:@32318.4]
  assign _T_85023 = _T_85022[13:0]; // @[Modules.scala 160:64:@32319.4]
  assign buffer_9_610 = $signed(_T_85023); // @[Modules.scala 160:64:@32320.4]
  assign _T_85025 = $signed(buffer_9_594) + $signed(buffer_9_595); // @[Modules.scala 160:64:@32322.4]
  assign _T_85026 = _T_85025[13:0]; // @[Modules.scala 160:64:@32323.4]
  assign buffer_9_611 = $signed(_T_85026); // @[Modules.scala 160:64:@32324.4]
  assign _T_85028 = $signed(buffer_9_596) + $signed(buffer_9_597); // @[Modules.scala 160:64:@32326.4]
  assign _T_85029 = _T_85028[13:0]; // @[Modules.scala 160:64:@32327.4]
  assign buffer_9_612 = $signed(_T_85029); // @[Modules.scala 160:64:@32328.4]
  assign _T_85031 = $signed(buffer_9_598) + $signed(buffer_9_599); // @[Modules.scala 160:64:@32330.4]
  assign _T_85032 = _T_85031[13:0]; // @[Modules.scala 160:64:@32331.4]
  assign buffer_9_613 = $signed(_T_85032); // @[Modules.scala 160:64:@32332.4]
  assign _T_85034 = $signed(buffer_9_600) + $signed(buffer_9_601); // @[Modules.scala 160:64:@32334.4]
  assign _T_85035 = _T_85034[13:0]; // @[Modules.scala 160:64:@32335.4]
  assign buffer_9_614 = $signed(_T_85035); // @[Modules.scala 160:64:@32336.4]
  assign _T_85037 = $signed(buffer_9_602) + $signed(buffer_9_603); // @[Modules.scala 160:64:@32338.4]
  assign _T_85038 = _T_85037[13:0]; // @[Modules.scala 160:64:@32339.4]
  assign buffer_9_615 = $signed(_T_85038); // @[Modules.scala 160:64:@32340.4]
  assign _T_85040 = $signed(buffer_9_604) + $signed(buffer_9_605); // @[Modules.scala 160:64:@32342.4]
  assign _T_85041 = _T_85040[13:0]; // @[Modules.scala 160:64:@32343.4]
  assign buffer_9_616 = $signed(_T_85041); // @[Modules.scala 160:64:@32344.4]
  assign _T_85043 = $signed(buffer_9_606) + $signed(buffer_9_607); // @[Modules.scala 160:64:@32346.4]
  assign _T_85044 = _T_85043[13:0]; // @[Modules.scala 160:64:@32347.4]
  assign buffer_9_617 = $signed(_T_85044); // @[Modules.scala 160:64:@32348.4]
  assign _T_85046 = $signed(buffer_9_608) + $signed(buffer_9_609); // @[Modules.scala 160:64:@32350.4]
  assign _T_85047 = _T_85046[13:0]; // @[Modules.scala 160:64:@32351.4]
  assign buffer_9_618 = $signed(_T_85047); // @[Modules.scala 160:64:@32352.4]
  assign _T_85049 = $signed(buffer_9_610) + $signed(buffer_9_611); // @[Modules.scala 160:64:@32354.4]
  assign _T_85050 = _T_85049[13:0]; // @[Modules.scala 160:64:@32355.4]
  assign buffer_9_619 = $signed(_T_85050); // @[Modules.scala 160:64:@32356.4]
  assign _T_85052 = $signed(buffer_9_612) + $signed(buffer_9_613); // @[Modules.scala 160:64:@32358.4]
  assign _T_85053 = _T_85052[13:0]; // @[Modules.scala 160:64:@32359.4]
  assign buffer_9_620 = $signed(_T_85053); // @[Modules.scala 160:64:@32360.4]
  assign _T_85055 = $signed(buffer_9_614) + $signed(buffer_9_615); // @[Modules.scala 160:64:@32362.4]
  assign _T_85056 = _T_85055[13:0]; // @[Modules.scala 160:64:@32363.4]
  assign buffer_9_621 = $signed(_T_85056); // @[Modules.scala 160:64:@32364.4]
  assign _T_85058 = $signed(buffer_9_616) + $signed(buffer_9_617); // @[Modules.scala 160:64:@32366.4]
  assign _T_85059 = _T_85058[13:0]; // @[Modules.scala 160:64:@32367.4]
  assign buffer_9_622 = $signed(_T_85059); // @[Modules.scala 160:64:@32368.4]
  assign _T_85061 = $signed(buffer_9_618) + $signed(buffer_9_619); // @[Modules.scala 166:64:@32370.4]
  assign _T_85062 = _T_85061[13:0]; // @[Modules.scala 166:64:@32371.4]
  assign buffer_9_623 = $signed(_T_85062); // @[Modules.scala 166:64:@32372.4]
  assign _T_85064 = $signed(buffer_9_620) + $signed(buffer_9_621); // @[Modules.scala 166:64:@32374.4]
  assign _T_85065 = _T_85064[13:0]; // @[Modules.scala 166:64:@32375.4]
  assign buffer_9_624 = $signed(_T_85065); // @[Modules.scala 166:64:@32376.4]
  assign _T_85067 = $signed(buffer_9_623) + $signed(buffer_9_624); // @[Modules.scala 160:64:@32378.4]
  assign _T_85068 = _T_85067[13:0]; // @[Modules.scala 160:64:@32379.4]
  assign buffer_9_625 = $signed(_T_85068); // @[Modules.scala 160:64:@32380.4]
  assign _T_85070 = $signed(buffer_9_625) + $signed(buffer_9_622); // @[Modules.scala 172:66:@32382.4]
  assign _T_85071 = _T_85070[13:0]; // @[Modules.scala 172:66:@32383.4]
  assign buffer_9_626 = $signed(_T_85071); // @[Modules.scala 172:66:@32384.4]
  assign _GEN_694 = {{1{_T_60255[4]}},_T_60255}; // @[Modules.scala 150:103:@32545.4]
  assign _T_85077 = $signed(_T_54199) + $signed(_GEN_694); // @[Modules.scala 150:103:@32545.4]
  assign _T_85078 = _T_85077[5:0]; // @[Modules.scala 150:103:@32546.4]
  assign _T_85079 = $signed(_T_85078); // @[Modules.scala 150:103:@32547.4]
  assign _T_85084 = $signed(_T_60257) + $signed(_T_57227); // @[Modules.scala 150:103:@32551.4]
  assign _T_85085 = _T_85084[4:0]; // @[Modules.scala 150:103:@32552.4]
  assign _T_85086 = $signed(_T_85085); // @[Modules.scala 150:103:@32553.4]
  assign _GEN_695 = {{1{_T_60264[4]}},_T_60264}; // @[Modules.scala 150:103:@32557.4]
  assign _T_85091 = $signed(_GEN_695) + $signed(_T_57232); // @[Modules.scala 150:103:@32557.4]
  assign _T_85092 = _T_85091[5:0]; // @[Modules.scala 150:103:@32558.4]
  assign _T_85093 = $signed(_T_85092); // @[Modules.scala 150:103:@32559.4]
  assign _T_85098 = $signed(_T_57234) + $signed(_T_54222); // @[Modules.scala 150:103:@32563.4]
  assign _T_85099 = _T_85098[5:0]; // @[Modules.scala 150:103:@32564.4]
  assign _T_85100 = $signed(_T_85099); // @[Modules.scala 150:103:@32565.4]
  assign _GEN_696 = {{1{_T_57274[4]}},_T_57274}; // @[Modules.scala 150:103:@32599.4]
  assign _T_85140 = $signed(_T_54264) + $signed(_GEN_696); // @[Modules.scala 150:103:@32599.4]
  assign _T_85141 = _T_85140[5:0]; // @[Modules.scala 150:103:@32600.4]
  assign _T_85142 = $signed(_T_85141); // @[Modules.scala 150:103:@32601.4]
  assign _T_85154 = $signed(_T_60327) + $signed(_T_57288); // @[Modules.scala 150:103:@32611.4]
  assign _T_85155 = _T_85154[4:0]; // @[Modules.scala 150:103:@32612.4]
  assign _T_85156 = $signed(_T_85155); // @[Modules.scala 150:103:@32613.4]
  assign _T_85231 = $signed(_T_54355) + $signed(_T_63499); // @[Modules.scala 150:103:@32677.4]
  assign _T_85232 = _T_85231[4:0]; // @[Modules.scala 150:103:@32678.4]
  assign _T_85233 = $signed(_T_85232); // @[Modules.scala 150:103:@32679.4]
  assign _T_85252 = $signed(_T_54376) + $signed(_T_54381); // @[Modules.scala 150:103:@32695.4]
  assign _T_85253 = _T_85252[5:0]; // @[Modules.scala 150:103:@32696.4]
  assign _T_85254 = $signed(_T_85253); // @[Modules.scala 150:103:@32697.4]
  assign _T_85266 = $signed(_T_54390) + $signed(_T_54395); // @[Modules.scala 150:103:@32707.4]
  assign _T_85267 = _T_85266[5:0]; // @[Modules.scala 150:103:@32708.4]
  assign _T_85268 = $signed(_T_85267); // @[Modules.scala 150:103:@32709.4]
  assign _T_85322 = $signed(_T_63585) + $signed(_T_63590); // @[Modules.scala 150:103:@32755.4]
  assign _T_85323 = _T_85322[4:0]; // @[Modules.scala 150:103:@32756.4]
  assign _T_85324 = $signed(_T_85323); // @[Modules.scala 150:103:@32757.4]
  assign _T_85329 = $signed(_GEN_4) + $signed(_T_60488); // @[Modules.scala 150:103:@32761.4]
  assign _T_85330 = _T_85329[5:0]; // @[Modules.scala 150:103:@32762.4]
  assign _T_85331 = $signed(_T_85330); // @[Modules.scala 150:103:@32763.4]
  assign _T_85357 = $signed(_T_54481) + $signed(_T_69749); // @[Modules.scala 150:103:@32785.4]
  assign _T_85358 = _T_85357[5:0]; // @[Modules.scala 150:103:@32786.4]
  assign _T_85359 = $signed(_T_85358); // @[Modules.scala 150:103:@32787.4]
  assign _T_85371 = $signed(_T_76057) + $signed(_T_69763); // @[Modules.scala 150:103:@32797.4]
  assign _T_85372 = _T_85371[4:0]; // @[Modules.scala 150:103:@32798.4]
  assign _T_85373 = $signed(_T_85372); // @[Modules.scala 150:103:@32799.4]
  assign _T_85378 = $signed(_T_69765) + $signed(_T_69770); // @[Modules.scala 150:103:@32803.4]
  assign _T_85379 = _T_85378[4:0]; // @[Modules.scala 150:103:@32804.4]
  assign _T_85380 = $signed(_T_85379); // @[Modules.scala 150:103:@32805.4]
  assign _T_85399 = $signed(_T_57526) + $signed(_GEN_154); // @[Modules.scala 150:103:@32821.4]
  assign _T_85400 = _T_85399[5:0]; // @[Modules.scala 150:103:@32822.4]
  assign _T_85401 = $signed(_T_85400); // @[Modules.scala 150:103:@32823.4]
  assign _T_85406 = $signed(_T_63669) + $signed(_T_60563); // @[Modules.scala 150:103:@32827.4]
  assign _T_85407 = _T_85406[4:0]; // @[Modules.scala 150:103:@32828.4]
  assign _T_85408 = $signed(_T_85407); // @[Modules.scala 150:103:@32829.4]
  assign _T_85413 = $signed(_T_54523) + $signed(_T_54528); // @[Modules.scala 150:103:@32833.4]
  assign _T_85414 = _T_85413[4:0]; // @[Modules.scala 150:103:@32834.4]
  assign _T_85415 = $signed(_T_85414); // @[Modules.scala 150:103:@32835.4]
  assign _GEN_701 = {{1{_T_63688[4]}},_T_63688}; // @[Modules.scala 150:103:@32839.4]
  assign _T_85420 = $signed(_T_54530) + $signed(_GEN_701); // @[Modules.scala 150:103:@32839.4]
  assign _T_85421 = _T_85420[5:0]; // @[Modules.scala 150:103:@32840.4]
  assign _T_85422 = $signed(_T_85421); // @[Modules.scala 150:103:@32841.4]
  assign _T_85434 = $signed(_T_63704) + $signed(_T_76122); // @[Modules.scala 150:103:@32851.4]
  assign _T_85435 = _T_85434[5:0]; // @[Modules.scala 150:103:@32852.4]
  assign _T_85436 = $signed(_T_85435); // @[Modules.scala 150:103:@32853.4]
  assign _T_85469 = $signed(_T_60628) + $signed(_T_60633); // @[Modules.scala 150:103:@32881.4]
  assign _T_85470 = _T_85469[5:0]; // @[Modules.scala 150:103:@32882.4]
  assign _T_85471 = $signed(_T_85470); // @[Modules.scala 150:103:@32883.4]
  assign _T_85476 = $signed(_T_54586) + $signed(_GEN_160); // @[Modules.scala 150:103:@32887.4]
  assign _T_85477 = _T_85476[5:0]; // @[Modules.scala 150:103:@32888.4]
  assign _T_85478 = $signed(_T_85477); // @[Modules.scala 150:103:@32889.4]
  assign _T_85490 = $signed(_T_63774) + $signed(_T_57619); // @[Modules.scala 150:103:@32899.4]
  assign _T_85491 = _T_85490[4:0]; // @[Modules.scala 150:103:@32900.4]
  assign _T_85492 = $signed(_T_85491); // @[Modules.scala 150:103:@32901.4]
  assign _GEN_703 = {{1{_T_60689[4]}},_T_60689}; // @[Modules.scala 150:103:@32923.4]
  assign _T_85518 = $signed(_T_66920) + $signed(_GEN_703); // @[Modules.scala 150:103:@32923.4]
  assign _T_85519 = _T_85518[5:0]; // @[Modules.scala 150:103:@32924.4]
  assign _T_85520 = $signed(_T_85519); // @[Modules.scala 150:103:@32925.4]
  assign _T_85525 = $signed(_T_60691) + $signed(_T_54635); // @[Modules.scala 150:103:@32929.4]
  assign _T_85526 = _T_85525[4:0]; // @[Modules.scala 150:103:@32930.4]
  assign _T_85527 = $signed(_T_85526); // @[Modules.scala 150:103:@32931.4]
  assign _T_85539 = $signed(_T_54649) + $signed(_T_63828); // @[Modules.scala 150:103:@32941.4]
  assign _T_85540 = _T_85539[4:0]; // @[Modules.scala 150:103:@32942.4]
  assign _T_85541 = $signed(_T_85540); // @[Modules.scala 150:103:@32943.4]
  assign _GEN_704 = {{1{_T_69947[4]}},_T_69947}; // @[Modules.scala 150:103:@32947.4]
  assign _T_85546 = $signed(_T_57675) + $signed(_GEN_704); // @[Modules.scala 150:103:@32947.4]
  assign _T_85547 = _T_85546[5:0]; // @[Modules.scala 150:103:@32948.4]
  assign _T_85548 = $signed(_T_85547); // @[Modules.scala 150:103:@32949.4]
  assign _GEN_705 = {{1{_T_60724[4]}},_T_60724}; // @[Modules.scala 150:103:@32953.4]
  assign _T_85553 = $signed(_T_54668) + $signed(_GEN_705); // @[Modules.scala 150:103:@32953.4]
  assign _T_85554 = _T_85553[5:0]; // @[Modules.scala 150:103:@32954.4]
  assign _T_85555 = $signed(_T_85554); // @[Modules.scala 150:103:@32955.4]
  assign _T_85588 = $signed(_T_54698) + $signed(_T_54705); // @[Modules.scala 150:103:@32983.4]
  assign _T_85589 = _T_85588[4:0]; // @[Modules.scala 150:103:@32984.4]
  assign _T_85590 = $signed(_T_85589); // @[Modules.scala 150:103:@32985.4]
  assign _T_85609 = $signed(_GEN_296) + $signed(_T_57764); // @[Modules.scala 150:103:@33001.4]
  assign _T_85610 = _T_85609[5:0]; // @[Modules.scala 150:103:@33002.4]
  assign _T_85611 = $signed(_T_85610); // @[Modules.scala 150:103:@33003.4]
  assign _T_85616 = $signed(_T_70036) + $signed(_T_60808); // @[Modules.scala 150:103:@33007.4]
  assign _T_85617 = _T_85616[4:0]; // @[Modules.scala 150:103:@33008.4]
  assign _T_85618 = $signed(_T_85617); // @[Modules.scala 150:103:@33009.4]
  assign _T_85637 = $signed(_T_60829) + $signed(_T_54759); // @[Modules.scala 150:103:@33025.4]
  assign _T_85638 = _T_85637[4:0]; // @[Modules.scala 150:103:@33026.4]
  assign _T_85639 = $signed(_T_85638); // @[Modules.scala 150:103:@33027.4]
  assign _GEN_707 = {{1{_T_54787[4]}},_T_54787}; // @[Modules.scala 150:103:@33049.4]
  assign _T_85665 = $signed(_T_63970) + $signed(_GEN_707); // @[Modules.scala 150:103:@33049.4]
  assign _T_85666 = _T_85665[5:0]; // @[Modules.scala 150:103:@33050.4]
  assign _T_85667 = $signed(_T_85666); // @[Modules.scala 150:103:@33051.4]
  assign _GEN_709 = {{1{_T_63996[4]}},_T_63996}; // @[Modules.scala 150:103:@33073.4]
  assign _T_85693 = $signed(_T_57850) + $signed(_GEN_709); // @[Modules.scala 150:103:@33073.4]
  assign _T_85694 = _T_85693[5:0]; // @[Modules.scala 150:103:@33074.4]
  assign _T_85695 = $signed(_T_85694); // @[Modules.scala 150:103:@33075.4]
  assign _T_85707 = $signed(_T_60906) + $signed(_T_57869); // @[Modules.scala 150:103:@33085.4]
  assign _T_85708 = _T_85707[4:0]; // @[Modules.scala 150:103:@33086.4]
  assign _T_85709 = $signed(_T_85708); // @[Modules.scala 150:103:@33087.4]
  assign _T_85714 = $signed(_GEN_167) + $signed(_T_64019); // @[Modules.scala 150:103:@33091.4]
  assign _T_85715 = _T_85714[5:0]; // @[Modules.scala 150:103:@33092.4]
  assign _T_85716 = $signed(_T_85715); // @[Modules.scala 150:103:@33093.4]
  assign _T_85728 = $signed(_GEN_453) + $signed(_T_67135); // @[Modules.scala 150:103:@33103.4]
  assign _T_85729 = _T_85728[5:0]; // @[Modules.scala 150:103:@33104.4]
  assign _T_85730 = $signed(_T_85729); // @[Modules.scala 150:103:@33105.4]
  assign _T_85777 = $signed(_T_54887) + $signed(_T_54892); // @[Modules.scala 150:103:@33145.4]
  assign _T_85778 = _T_85777[4:0]; // @[Modules.scala 150:103:@33146.4]
  assign _T_85779 = $signed(_T_85778); // @[Modules.scala 150:103:@33147.4]
  assign _T_85805 = $signed(_T_64103) + $signed(_T_64108); // @[Modules.scala 150:103:@33169.4]
  assign _T_85806 = _T_85805[5:0]; // @[Modules.scala 150:103:@33170.4]
  assign _T_85807 = $signed(_T_85806); // @[Modules.scala 150:103:@33171.4]
  assign _T_85819 = $signed(_T_61006) + $signed(_GEN_99); // @[Modules.scala 150:103:@33181.4]
  assign _T_85820 = _T_85819[5:0]; // @[Modules.scala 150:103:@33182.4]
  assign _T_85821 = $signed(_T_85820); // @[Modules.scala 150:103:@33183.4]
  assign _T_85840 = $signed(_T_61025) + $signed(_T_54957); // @[Modules.scala 150:103:@33199.4]
  assign _T_85841 = _T_85840[4:0]; // @[Modules.scala 150:103:@33200.4]
  assign _T_85842 = $signed(_T_85841); // @[Modules.scala 150:103:@33201.4]
  assign _T_85868 = $signed(_T_64173) + $signed(_T_54985); // @[Modules.scala 150:103:@33223.4]
  assign _T_85869 = _T_85868[4:0]; // @[Modules.scala 150:103:@33224.4]
  assign _T_85870 = $signed(_T_85869); // @[Modules.scala 150:103:@33225.4]
  assign _T_85875 = $signed(_T_61062) + $signed(_T_54992); // @[Modules.scala 150:103:@33229.4]
  assign _T_85876 = _T_85875[4:0]; // @[Modules.scala 150:103:@33230.4]
  assign _T_85877 = $signed(_T_85876); // @[Modules.scala 150:103:@33231.4]
  assign _T_85882 = $signed(_T_61069) + $signed(_T_54999); // @[Modules.scala 150:103:@33235.4]
  assign _T_85883 = _T_85882[4:0]; // @[Modules.scala 150:103:@33236.4]
  assign _T_85884 = $signed(_T_85883); // @[Modules.scala 150:103:@33237.4]
  assign _T_85924 = $signed(_GEN_306) + $signed(_T_58072); // @[Modules.scala 150:103:@33271.4]
  assign _T_85925 = _T_85924[5:0]; // @[Modules.scala 150:103:@33272.4]
  assign _T_85926 = $signed(_T_85925); // @[Modules.scala 150:103:@33273.4]
  assign _T_85938 = $signed(_T_58081) + $signed(_T_67324); // @[Modules.scala 150:103:@33283.4]
  assign _T_85939 = _T_85938[5:0]; // @[Modules.scala 150:103:@33284.4]
  assign _T_85940 = $signed(_T_85939); // @[Modules.scala 150:103:@33285.4]
  assign _T_85987 = $signed(_T_61165) + $signed(_GEN_102); // @[Modules.scala 150:103:@33325.4]
  assign _T_85988 = _T_85987[5:0]; // @[Modules.scala 150:103:@33326.4]
  assign _T_85989 = $signed(_T_85988); // @[Modules.scala 150:103:@33327.4]
  assign _GEN_719 = {{1{_T_55116[4]}},_T_55116}; // @[Modules.scala 150:103:@33337.4]
  assign _T_86001 = $signed(_GEN_719) + $signed(_T_58142); // @[Modules.scala 150:103:@33337.4]
  assign _T_86002 = _T_86001[5:0]; // @[Modules.scala 150:103:@33338.4]
  assign _T_86003 = $signed(_T_86002); // @[Modules.scala 150:103:@33339.4]
  assign _T_86015 = $signed(_T_58151) + $signed(_T_58158); // @[Modules.scala 150:103:@33349.4]
  assign _T_86016 = _T_86015[5:0]; // @[Modules.scala 150:103:@33350.4]
  assign _T_86017 = $signed(_T_86016); // @[Modules.scala 150:103:@33351.4]
  assign _T_86036 = $signed(_T_61216) + $signed(_T_55151); // @[Modules.scala 150:103:@33367.4]
  assign _T_86037 = _T_86036[5:0]; // @[Modules.scala 150:103:@33368.4]
  assign _T_86038 = $signed(_T_86037); // @[Modules.scala 150:103:@33369.4]
  assign _T_86106 = $signed(_T_58235) + $signed(_GEN_33); // @[Modules.scala 150:103:@33427.4]
  assign _T_86107 = _T_86106[5:0]; // @[Modules.scala 150:103:@33428.4]
  assign _T_86108 = $signed(_T_86107); // @[Modules.scala 150:103:@33429.4]
  assign _T_86127 = $signed(_T_61307) + $signed(_GEN_317); // @[Modules.scala 150:103:@33445.4]
  assign _T_86128 = _T_86127[5:0]; // @[Modules.scala 150:103:@33446.4]
  assign _T_86129 = $signed(_T_86128); // @[Modules.scala 150:103:@33447.4]
  assign _T_86134 = $signed(_T_55235) + $signed(_T_58268); // @[Modules.scala 150:103:@33451.4]
  assign _T_86135 = _T_86134[5:0]; // @[Modules.scala 150:103:@33452.4]
  assign _T_86136 = $signed(_T_86135); // @[Modules.scala 150:103:@33453.4]
  assign _T_86155 = $signed(_T_64458) + $signed(_T_70533); // @[Modules.scala 150:103:@33469.4]
  assign _T_86156 = _T_86155[4:0]; // @[Modules.scala 150:103:@33470.4]
  assign _T_86157 = $signed(_T_86156); // @[Modules.scala 150:103:@33471.4]
  assign _T_86204 = $signed(_T_55305) + $signed(_T_70589); // @[Modules.scala 150:103:@33511.4]
  assign _T_86205 = _T_86204[4:0]; // @[Modules.scala 150:103:@33512.4]
  assign _T_86206 = $signed(_T_86205); // @[Modules.scala 150:103:@33513.4]
  assign _T_86225 = $signed(_T_55319) + $signed(_T_70605); // @[Modules.scala 150:103:@33529.4]
  assign _T_86226 = _T_86225[5:0]; // @[Modules.scala 150:103:@33530.4]
  assign _T_86227 = $signed(_T_86226); // @[Modules.scala 150:103:@33531.4]
  assign _GEN_726 = {{1{_T_55356[4]}},_T_55356}; // @[Modules.scala 150:103:@33565.4]
  assign _T_86267 = $signed(_GEN_726) + $signed(_T_61447); // @[Modules.scala 150:103:@33565.4]
  assign _T_86268 = _T_86267[5:0]; // @[Modules.scala 150:103:@33566.4]
  assign _T_86269 = $signed(_T_86268); // @[Modules.scala 150:103:@33567.4]
  assign _T_86274 = $signed(_T_55363) + $signed(_T_55368); // @[Modules.scala 150:103:@33571.4]
  assign _T_86275 = _T_86274[5:0]; // @[Modules.scala 150:103:@33572.4]
  assign _T_86276 = $signed(_T_86275); // @[Modules.scala 150:103:@33573.4]
  assign _GEN_729 = {{1{_T_64614[4]}},_T_64614}; // @[Modules.scala 150:103:@33619.4]
  assign _T_86330 = $signed(_T_61503) + $signed(_GEN_729); // @[Modules.scala 150:103:@33619.4]
  assign _T_86331 = _T_86330[5:0]; // @[Modules.scala 150:103:@33620.4]
  assign _T_86332 = $signed(_T_86331); // @[Modules.scala 150:103:@33621.4]
  assign _T_86344 = $signed(_GEN_325) + $signed(_T_55438); // @[Modules.scala 150:103:@33631.4]
  assign _T_86345 = _T_86344[5:0]; // @[Modules.scala 150:103:@33632.4]
  assign _T_86346 = $signed(_T_86345); // @[Modules.scala 150:103:@33633.4]
  assign _GEN_731 = {{1{_T_58452[4]}},_T_58452}; // @[Modules.scala 150:103:@33637.4]
  assign _T_86351 = $signed(_GEN_731) + $signed(_T_55440); // @[Modules.scala 150:103:@33637.4]
  assign _T_86352 = _T_86351[5:0]; // @[Modules.scala 150:103:@33638.4]
  assign _T_86353 = $signed(_T_86352); // @[Modules.scala 150:103:@33639.4]
  assign _GEN_732 = {{1{_T_58473[4]}},_T_58473}; // @[Modules.scala 150:103:@33655.4]
  assign _T_86372 = $signed(_T_55454) + $signed(_GEN_732); // @[Modules.scala 150:103:@33655.4]
  assign _T_86373 = _T_86372[5:0]; // @[Modules.scala 150:103:@33656.4]
  assign _T_86374 = $signed(_T_86373); // @[Modules.scala 150:103:@33657.4]
  assign _T_86379 = $signed(_T_55461) + $signed(_T_55466); // @[Modules.scala 150:103:@33661.4]
  assign _T_86380 = _T_86379[4:0]; // @[Modules.scala 150:103:@33662.4]
  assign _T_86381 = $signed(_T_86380); // @[Modules.scala 150:103:@33663.4]
  assign _T_86386 = $signed(_T_61552) + $signed(_T_64675); // @[Modules.scala 150:103:@33667.4]
  assign _T_86387 = _T_86386[4:0]; // @[Modules.scala 150:103:@33668.4]
  assign _T_86388 = $signed(_T_86387); // @[Modules.scala 150:103:@33669.4]
  assign _T_86393 = $signed(_T_64677) + $signed(_T_61564); // @[Modules.scala 150:103:@33673.4]
  assign _T_86394 = _T_86393[4:0]; // @[Modules.scala 150:103:@33674.4]
  assign _T_86395 = $signed(_T_86394); // @[Modules.scala 150:103:@33675.4]
  assign _T_86414 = $signed(_T_58501) + $signed(_GEN_53); // @[Modules.scala 150:103:@33691.4]
  assign _T_86415 = _T_86414[5:0]; // @[Modules.scala 150:103:@33692.4]
  assign _T_86416 = $signed(_T_86415); // @[Modules.scala 150:103:@33693.4]
  assign _T_86456 = $signed(_T_55522) + $signed(_GEN_331); // @[Modules.scala 150:103:@33727.4]
  assign _T_86457 = _T_86456[5:0]; // @[Modules.scala 150:103:@33728.4]
  assign _T_86458 = $signed(_T_86457); // @[Modules.scala 150:103:@33729.4]
  assign _T_86463 = $signed(_T_55536) + $signed(_T_58562); // @[Modules.scala 150:103:@33733.4]
  assign _T_86464 = _T_86463[4:0]; // @[Modules.scala 150:103:@33734.4]
  assign _T_86465 = $signed(_T_86464); // @[Modules.scala 150:103:@33735.4]
  assign _T_86470 = $signed(_T_58564) + $signed(_T_64754); // @[Modules.scala 150:103:@33739.4]
  assign _T_86471 = _T_86470[4:0]; // @[Modules.scala 150:103:@33740.4]
  assign _T_86472 = $signed(_T_86471); // @[Modules.scala 150:103:@33741.4]
  assign _T_86484 = $signed(_T_55552) + $signed(_GEN_251); // @[Modules.scala 150:103:@33751.4]
  assign _T_86485 = _T_86484[5:0]; // @[Modules.scala 150:103:@33752.4]
  assign _T_86486 = $signed(_T_86485); // @[Modules.scala 150:103:@33753.4]
  assign _T_86491 = $signed(_T_55559) + $signed(_T_70855); // @[Modules.scala 150:103:@33757.4]
  assign _T_86492 = _T_86491[4:0]; // @[Modules.scala 150:103:@33758.4]
  assign _T_86493 = $signed(_T_86492); // @[Modules.scala 150:103:@33759.4]
  assign _T_86568 = $signed(_T_58660) + $signed(_T_64871); // @[Modules.scala 150:103:@33823.4]
  assign _T_86569 = _T_86568[4:0]; // @[Modules.scala 150:103:@33824.4]
  assign _T_86570 = $signed(_T_86569); // @[Modules.scala 150:103:@33825.4]
  assign _GEN_738 = {{1{_T_64906[4]}},_T_64906}; // @[Modules.scala 150:103:@33859.4]
  assign _T_86610 = $signed(_T_55690) + $signed(_GEN_738); // @[Modules.scala 150:103:@33859.4]
  assign _T_86611 = _T_86610[5:0]; // @[Modules.scala 150:103:@33860.4]
  assign _T_86612 = $signed(_T_86611); // @[Modules.scala 150:103:@33861.4]
  assign _GEN_739 = {{1{_T_67928[4]}},_T_67928}; // @[Modules.scala 150:103:@33871.4]
  assign _T_86624 = $signed(_GEN_739) + $signed(_T_71004); // @[Modules.scala 150:103:@33871.4]
  assign _T_86625 = _T_86624[5:0]; // @[Modules.scala 150:103:@33872.4]
  assign _T_86626 = $signed(_T_86625); // @[Modules.scala 150:103:@33873.4]
  assign _T_86659 = $signed(_GEN_122) + $signed(_T_55746); // @[Modules.scala 150:103:@33901.4]
  assign _T_86660 = _T_86659[5:0]; // @[Modules.scala 150:103:@33902.4]
  assign _T_86661 = $signed(_T_86660); // @[Modules.scala 150:103:@33903.4]
  assign _GEN_742 = {{1{_T_58767[4]}},_T_58767}; // @[Modules.scala 150:103:@33919.4]
  assign _T_86680 = $signed(_GEN_742) + $signed(_T_61846); // @[Modules.scala 150:103:@33919.4]
  assign _T_86681 = _T_86680[5:0]; // @[Modules.scala 150:103:@33920.4]
  assign _T_86682 = $signed(_T_86681); // @[Modules.scala 150:103:@33921.4]
  assign _T_86687 = $signed(_T_58779) + $signed(_T_55769); // @[Modules.scala 150:103:@33925.4]
  assign _T_86688 = _T_86687[4:0]; // @[Modules.scala 150:103:@33926.4]
  assign _T_86689 = $signed(_T_86688); // @[Modules.scala 150:103:@33927.4]
  assign _T_86694 = $signed(_T_71088) + $signed(_T_65004); // @[Modules.scala 150:103:@33931.4]
  assign _T_86695 = _T_86694[5:0]; // @[Modules.scala 150:103:@33932.4]
  assign _T_86696 = $signed(_T_86695); // @[Modules.scala 150:103:@33933.4]
  assign _T_86708 = $signed(_T_58809) + $signed(_T_55788); // @[Modules.scala 150:103:@33943.4]
  assign _T_86709 = _T_86708[5:0]; // @[Modules.scala 150:103:@33944.4]
  assign _T_86710 = $signed(_T_86709); // @[Modules.scala 150:103:@33945.4]
  assign _T_86736 = $signed(_GEN_679) + $signed(_T_71137); // @[Modules.scala 150:103:@33967.4]
  assign _T_86737 = _T_86736[5:0]; // @[Modules.scala 150:103:@33968.4]
  assign _T_86738 = $signed(_T_86737); // @[Modules.scala 150:103:@33969.4]
  assign _T_86757 = $signed(_T_68075) + $signed(_T_65048); // @[Modules.scala 150:103:@33985.4]
  assign _T_86758 = _T_86757[4:0]; // @[Modules.scala 150:103:@33986.4]
  assign _T_86759 = $signed(_T_86758); // @[Modules.scala 150:103:@33987.4]
  assign _T_86764 = $signed(_T_71179) + $signed(_T_55844); // @[Modules.scala 150:103:@33991.4]
  assign _T_86765 = _T_86764[5:0]; // @[Modules.scala 150:103:@33992.4]
  assign _T_86766 = $signed(_T_86765); // @[Modules.scala 150:103:@33993.4]
  assign _T_86785 = $signed(_T_55860) + $signed(_GEN_129); // @[Modules.scala 150:103:@34009.4]
  assign _T_86786 = _T_86785[5:0]; // @[Modules.scala 150:103:@34010.4]
  assign _T_86787 = $signed(_T_86786); // @[Modules.scala 150:103:@34011.4]
  assign _T_86834 = $signed(_GEN_549) + $signed(_T_58933); // @[Modules.scala 150:103:@34051.4]
  assign _T_86835 = _T_86834[5:0]; // @[Modules.scala 150:103:@34052.4]
  assign _T_86836 = $signed(_T_86835); // @[Modules.scala 150:103:@34053.4]
  assign _T_86841 = $signed(_T_55916) + $signed(_T_68171); // @[Modules.scala 150:103:@34057.4]
  assign _T_86842 = _T_86841[4:0]; // @[Modules.scala 150:103:@34058.4]
  assign _T_86843 = $signed(_T_86842); // @[Modules.scala 150:103:@34059.4]
  assign _T_86862 = $signed(_T_55937) + $signed(_T_55944); // @[Modules.scala 150:103:@34075.4]
  assign _T_86863 = _T_86862[5:0]; // @[Modules.scala 150:103:@34076.4]
  assign _T_86864 = $signed(_T_86863); // @[Modules.scala 150:103:@34077.4]
  assign _T_86869 = $signed(_T_68194) + $signed(_T_62049); // @[Modules.scala 150:103:@34081.4]
  assign _T_86870 = _T_86869[4:0]; // @[Modules.scala 150:103:@34082.4]
  assign _T_86871 = $signed(_T_86870); // @[Modules.scala 150:103:@34083.4]
  assign _T_86883 = $signed(_T_62063) + $signed(_T_55972); // @[Modules.scala 150:103:@34093.4]
  assign _T_86884 = _T_86883[4:0]; // @[Modules.scala 150:103:@34094.4]
  assign _T_86885 = $signed(_T_86884); // @[Modules.scala 150:103:@34095.4]
  assign _GEN_749 = {{1{_T_56007[4]}},_T_56007}; // @[Modules.scala 150:103:@34117.4]
  assign _T_86911 = $signed(_GEN_749) + $signed(_T_62110); // @[Modules.scala 150:103:@34117.4]
  assign _T_86912 = _T_86911[5:0]; // @[Modules.scala 150:103:@34118.4]
  assign _T_86913 = $signed(_T_86912); // @[Modules.scala 150:103:@34119.4]
  assign _T_86918 = $signed(_T_62112) + $signed(_T_65221); // @[Modules.scala 150:103:@34123.4]
  assign _T_86919 = _T_86918[5:0]; // @[Modules.scala 150:103:@34124.4]
  assign _T_86920 = $signed(_T_86919); // @[Modules.scala 150:103:@34125.4]
  assign _T_86974 = $signed(_T_71389) + $signed(_T_71394); // @[Modules.scala 150:103:@34171.4]
  assign _T_86975 = _T_86974[5:0]; // @[Modules.scala 150:103:@34172.4]
  assign _T_86976 = $signed(_T_86975); // @[Modules.scala 150:103:@34173.4]
  assign _T_86981 = $signed(_T_71396) + $signed(_T_59080); // @[Modules.scala 150:103:@34177.4]
  assign _T_86982 = _T_86981[5:0]; // @[Modules.scala 150:103:@34178.4]
  assign _T_86983 = $signed(_T_86982); // @[Modules.scala 150:103:@34179.4]
  assign _T_87009 = $signed(_T_56103) + $signed(_GEN_423); // @[Modules.scala 150:103:@34201.4]
  assign _T_87010 = _T_87009[5:0]; // @[Modules.scala 150:103:@34202.4]
  assign _T_87011 = $signed(_T_87010); // @[Modules.scala 150:103:@34203.4]
  assign _T_87016 = $signed(_T_56110) + $signed(_GEN_138); // @[Modules.scala 150:103:@34207.4]
  assign _T_87017 = _T_87016[5:0]; // @[Modules.scala 150:103:@34208.4]
  assign _T_87018 = $signed(_T_87017); // @[Modules.scala 150:103:@34209.4]
  assign _T_87023 = $signed(_T_62210) + $signed(_T_62215); // @[Modules.scala 150:103:@34213.4]
  assign _T_87024 = _T_87023[4:0]; // @[Modules.scala 150:103:@34214.4]
  assign _T_87025 = $signed(_T_87024); // @[Modules.scala 150:103:@34215.4]
  assign _GEN_753 = {{1{_T_56180[4]}},_T_56180}; // @[Modules.scala 150:103:@34267.4]
  assign _T_87086 = $signed(_T_65382) + $signed(_GEN_753); // @[Modules.scala 150:103:@34267.4]
  assign _T_87087 = _T_87086[5:0]; // @[Modules.scala 150:103:@34268.4]
  assign _T_87088 = $signed(_T_87087); // @[Modules.scala 150:103:@34269.4]
  assign _GEN_756 = {{1{_T_65410[4]}},_T_65410}; // @[Modules.scala 150:103:@34291.4]
  assign _T_87114 = $signed(_GEN_756) + $signed(_T_56196); // @[Modules.scala 150:103:@34291.4]
  assign _T_87115 = _T_87114[5:0]; // @[Modules.scala 150:103:@34292.4]
  assign _T_87116 = $signed(_T_87115); // @[Modules.scala 150:103:@34293.4]
  assign _GEN_757 = {{1{_T_62306[4]}},_T_62306}; // @[Modules.scala 150:103:@34297.4]
  assign _T_87121 = $signed(_T_56201) + $signed(_GEN_757); // @[Modules.scala 150:103:@34297.4]
  assign _T_87122 = _T_87121[5:0]; // @[Modules.scala 150:103:@34298.4]
  assign _T_87123 = $signed(_T_87122); // @[Modules.scala 150:103:@34299.4]
  assign _T_87163 = $signed(_T_56243) + $signed(_T_62348); // @[Modules.scala 150:103:@34333.4]
  assign _T_87164 = _T_87163[4:0]; // @[Modules.scala 150:103:@34334.4]
  assign _T_87165 = $signed(_T_87164); // @[Modules.scala 150:103:@34335.4]
  assign _T_87170 = $signed(_T_59264) + $signed(_GEN_142); // @[Modules.scala 150:103:@34339.4]
  assign _T_87171 = _T_87170[5:0]; // @[Modules.scala 150:103:@34340.4]
  assign _T_87172 = $signed(_T_87171); // @[Modules.scala 150:103:@34341.4]
  assign _GEN_759 = {{1{_T_65475[4]}},_T_65475}; // @[Modules.scala 150:103:@34345.4]
  assign _T_87177 = $signed(_GEN_759) + $signed(_T_56264); // @[Modules.scala 150:103:@34345.4]
  assign _T_87178 = _T_87177[5:0]; // @[Modules.scala 150:103:@34346.4]
  assign _T_87179 = $signed(_T_87178); // @[Modules.scala 150:103:@34347.4]
  assign buffer_10_0 = {{8{_T_85079[5]}},_T_85079}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_1 = {{9{_T_85086[4]}},_T_85086}; // @[Modules.scala 112:22:@8.4]
  assign _T_87224 = $signed(buffer_10_0) + $signed(buffer_10_1); // @[Modules.scala 160:64:@34387.4]
  assign _T_87225 = _T_87224[13:0]; // @[Modules.scala 160:64:@34388.4]
  assign buffer_10_308 = $signed(_T_87225); // @[Modules.scala 160:64:@34389.4]
  assign buffer_10_2 = {{8{_T_85093[5]}},_T_85093}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_3 = {{8{_T_85100[5]}},_T_85100}; // @[Modules.scala 112:22:@8.4]
  assign _T_87227 = $signed(buffer_10_2) + $signed(buffer_10_3); // @[Modules.scala 160:64:@34391.4]
  assign _T_87228 = _T_87227[13:0]; // @[Modules.scala 160:64:@34392.4]
  assign buffer_10_309 = $signed(_T_87228); // @[Modules.scala 160:64:@34393.4]
  assign _T_87233 = $signed(buffer_0_6) + $signed(buffer_3_7); // @[Modules.scala 160:64:@34399.4]
  assign _T_87234 = _T_87233[13:0]; // @[Modules.scala 160:64:@34400.4]
  assign buffer_10_311 = $signed(_T_87234); // @[Modules.scala 160:64:@34401.4]
  assign buffer_10_9 = {{8{_T_85142[5]}},_T_85142}; // @[Modules.scala 112:22:@8.4]
  assign _T_87236 = $signed(buffer_4_7) + $signed(buffer_10_9); // @[Modules.scala 160:64:@34403.4]
  assign _T_87237 = _T_87236[13:0]; // @[Modules.scala 160:64:@34404.4]
  assign buffer_10_312 = $signed(_T_87237); // @[Modules.scala 160:64:@34405.4]
  assign buffer_10_11 = {{9{_T_85156[4]}},_T_85156}; // @[Modules.scala 112:22:@8.4]
  assign _T_87239 = $signed(buffer_4_9) + $signed(buffer_10_11); // @[Modules.scala 160:64:@34407.4]
  assign _T_87240 = _T_87239[13:0]; // @[Modules.scala 160:64:@34408.4]
  assign buffer_10_313 = $signed(_T_87240); // @[Modules.scala 160:64:@34409.4]
  assign _T_87254 = $signed(buffer_0_20) + $signed(buffer_1_21); // @[Modules.scala 160:64:@34427.4]
  assign _T_87255 = _T_87254[13:0]; // @[Modules.scala 160:64:@34428.4]
  assign buffer_10_318 = $signed(_T_87255); // @[Modules.scala 160:64:@34429.4]
  assign buffer_10_22 = {{9{_T_85233[4]}},_T_85233}; // @[Modules.scala 112:22:@8.4]
  assign _T_87257 = $signed(buffer_10_22) + $signed(buffer_2_22); // @[Modules.scala 160:64:@34431.4]
  assign _T_87258 = _T_87257[13:0]; // @[Modules.scala 160:64:@34432.4]
  assign buffer_10_319 = $signed(_T_87258); // @[Modules.scala 160:64:@34433.4]
  assign buffer_10_25 = {{8{_T_85254[5]}},_T_85254}; // @[Modules.scala 112:22:@8.4]
  assign _T_87260 = $signed(buffer_2_23) + $signed(buffer_10_25); // @[Modules.scala 160:64:@34435.4]
  assign _T_87261 = _T_87260[13:0]; // @[Modules.scala 160:64:@34436.4]
  assign buffer_10_320 = $signed(_T_87261); // @[Modules.scala 160:64:@34437.4]
  assign buffer_10_27 = {{8{_T_85268[5]}},_T_85268}; // @[Modules.scala 112:22:@8.4]
  assign _T_87263 = $signed(buffer_6_26) + $signed(buffer_10_27); // @[Modules.scala 160:64:@34439.4]
  assign _T_87264 = _T_87263[13:0]; // @[Modules.scala 160:64:@34440.4]
  assign buffer_10_321 = $signed(_T_87264); // @[Modules.scala 160:64:@34441.4]
  assign _T_87266 = $signed(buffer_9_29) + $signed(buffer_2_27); // @[Modules.scala 160:64:@34443.4]
  assign _T_87267 = _T_87266[13:0]; // @[Modules.scala 160:64:@34444.4]
  assign buffer_10_322 = $signed(_T_87267); // @[Modules.scala 160:64:@34445.4]
  assign _T_87272 = $signed(buffer_8_34) + $signed(buffer_5_32); // @[Modules.scala 160:64:@34451.4]
  assign _T_87273 = _T_87272[13:0]; // @[Modules.scala 160:64:@34452.4]
  assign buffer_10_324 = $signed(_T_87273); // @[Modules.scala 160:64:@34453.4]
  assign buffer_10_35 = {{9{_T_85324[4]}},_T_85324}; // @[Modules.scala 112:22:@8.4]
  assign _T_87275 = $signed(buffer_0_35) + $signed(buffer_10_35); // @[Modules.scala 160:64:@34455.4]
  assign _T_87276 = _T_87275[13:0]; // @[Modules.scala 160:64:@34456.4]
  assign buffer_10_325 = $signed(_T_87276); // @[Modules.scala 160:64:@34457.4]
  assign buffer_10_36 = {{8{_T_85331[5]}},_T_85331}; // @[Modules.scala 112:22:@8.4]
  assign _T_87278 = $signed(buffer_10_36) + $signed(buffer_1_36); // @[Modules.scala 160:64:@34459.4]
  assign _T_87279 = _T_87278[13:0]; // @[Modules.scala 160:64:@34460.4]
  assign buffer_10_326 = $signed(_T_87279); // @[Modules.scala 160:64:@34461.4]
  assign _T_87281 = $signed(buffer_1_37) + $signed(buffer_1_38); // @[Modules.scala 160:64:@34463.4]
  assign _T_87282 = _T_87281[13:0]; // @[Modules.scala 160:64:@34464.4]
  assign buffer_10_327 = $signed(_T_87282); // @[Modules.scala 160:64:@34465.4]
  assign buffer_10_40 = {{8{_T_85359[5]}},_T_85359}; // @[Modules.scala 112:22:@8.4]
  assign _T_87284 = $signed(buffer_10_40) + $signed(buffer_0_41); // @[Modules.scala 160:64:@34467.4]
  assign _T_87285 = _T_87284[13:0]; // @[Modules.scala 160:64:@34468.4]
  assign buffer_10_328 = $signed(_T_87285); // @[Modules.scala 160:64:@34469.4]
  assign buffer_10_42 = {{9{_T_85373[4]}},_T_85373}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_43 = {{9{_T_85380[4]}},_T_85380}; // @[Modules.scala 112:22:@8.4]
  assign _T_87287 = $signed(buffer_10_42) + $signed(buffer_10_43); // @[Modules.scala 160:64:@34471.4]
  assign _T_87288 = _T_87287[13:0]; // @[Modules.scala 160:64:@34472.4]
  assign buffer_10_329 = $signed(_T_87288); // @[Modules.scala 160:64:@34473.4]
  assign buffer_10_46 = {{8{_T_85401[5]}},_T_85401}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_47 = {{9{_T_85408[4]}},_T_85408}; // @[Modules.scala 112:22:@8.4]
  assign _T_87293 = $signed(buffer_10_46) + $signed(buffer_10_47); // @[Modules.scala 160:64:@34479.4]
  assign _T_87294 = _T_87293[13:0]; // @[Modules.scala 160:64:@34480.4]
  assign buffer_10_331 = $signed(_T_87294); // @[Modules.scala 160:64:@34481.4]
  assign buffer_10_48 = {{9{_T_85415[4]}},_T_85415}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_49 = {{8{_T_85422[5]}},_T_85422}; // @[Modules.scala 112:22:@8.4]
  assign _T_87296 = $signed(buffer_10_48) + $signed(buffer_10_49); // @[Modules.scala 160:64:@34483.4]
  assign _T_87297 = _T_87296[13:0]; // @[Modules.scala 160:64:@34484.4]
  assign buffer_10_332 = $signed(_T_87297); // @[Modules.scala 160:64:@34485.4]
  assign buffer_10_51 = {{8{_T_85436[5]}},_T_85436}; // @[Modules.scala 112:22:@8.4]
  assign _T_87299 = $signed(buffer_1_49) + $signed(buffer_10_51); // @[Modules.scala 160:64:@34487.4]
  assign _T_87300 = _T_87299[13:0]; // @[Modules.scala 160:64:@34488.4]
  assign buffer_10_333 = $signed(_T_87300); // @[Modules.scala 160:64:@34489.4]
  assign buffer_10_56 = {{8{_T_85471[5]}},_T_85471}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_57 = {{8{_T_85478[5]}},_T_85478}; // @[Modules.scala 112:22:@8.4]
  assign _T_87308 = $signed(buffer_10_56) + $signed(buffer_10_57); // @[Modules.scala 160:64:@34499.4]
  assign _T_87309 = _T_87308[13:0]; // @[Modules.scala 160:64:@34500.4]
  assign buffer_10_336 = $signed(_T_87309); // @[Modules.scala 160:64:@34501.4]
  assign buffer_10_59 = {{9{_T_85492[4]}},_T_85492}; // @[Modules.scala 112:22:@8.4]
  assign _T_87311 = $signed(buffer_8_55) + $signed(buffer_10_59); // @[Modules.scala 160:64:@34503.4]
  assign _T_87312 = _T_87311[13:0]; // @[Modules.scala 160:64:@34504.4]
  assign buffer_10_337 = $signed(_T_87312); // @[Modules.scala 160:64:@34505.4]
  assign _T_87314 = $signed(buffer_5_61) + $signed(buffer_4_62); // @[Modules.scala 160:64:@34507.4]
  assign _T_87315 = _T_87314[13:0]; // @[Modules.scala 160:64:@34508.4]
  assign buffer_10_338 = $signed(_T_87315); // @[Modules.scala 160:64:@34509.4]
  assign buffer_10_63 = {{8{_T_85520[5]}},_T_85520}; // @[Modules.scala 112:22:@8.4]
  assign _T_87317 = $signed(buffer_5_63) + $signed(buffer_10_63); // @[Modules.scala 160:64:@34511.4]
  assign _T_87318 = _T_87317[13:0]; // @[Modules.scala 160:64:@34512.4]
  assign buffer_10_339 = $signed(_T_87318); // @[Modules.scala 160:64:@34513.4]
  assign buffer_10_64 = {{9{_T_85527[4]}},_T_85527}; // @[Modules.scala 112:22:@8.4]
  assign _T_87320 = $signed(buffer_10_64) + $signed(buffer_1_65); // @[Modules.scala 160:64:@34515.4]
  assign _T_87321 = _T_87320[13:0]; // @[Modules.scala 160:64:@34516.4]
  assign buffer_10_340 = $signed(_T_87321); // @[Modules.scala 160:64:@34517.4]
  assign buffer_10_66 = {{9{_T_85541[4]}},_T_85541}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_67 = {{8{_T_85548[5]}},_T_85548}; // @[Modules.scala 112:22:@8.4]
  assign _T_87323 = $signed(buffer_10_66) + $signed(buffer_10_67); // @[Modules.scala 160:64:@34519.4]
  assign _T_87324 = _T_87323[13:0]; // @[Modules.scala 160:64:@34520.4]
  assign buffer_10_341 = $signed(_T_87324); // @[Modules.scala 160:64:@34521.4]
  assign buffer_10_68 = {{8{_T_85555[5]}},_T_85555}; // @[Modules.scala 112:22:@8.4]
  assign _T_87326 = $signed(buffer_10_68) + $signed(buffer_3_72); // @[Modules.scala 160:64:@34523.4]
  assign _T_87327 = _T_87326[13:0]; // @[Modules.scala 160:64:@34524.4]
  assign buffer_10_342 = $signed(_T_87327); // @[Modules.scala 160:64:@34525.4]
  assign _T_87329 = $signed(buffer_3_73) + $signed(buffer_1_72); // @[Modules.scala 160:64:@34527.4]
  assign _T_87330 = _T_87329[13:0]; // @[Modules.scala 160:64:@34528.4]
  assign buffer_10_343 = $signed(_T_87330); // @[Modules.scala 160:64:@34529.4]
  assign buffer_10_73 = {{9{_T_85590[4]}},_T_85590}; // @[Modules.scala 112:22:@8.4]
  assign _T_87332 = $signed(buffer_1_73) + $signed(buffer_10_73); // @[Modules.scala 160:64:@34531.4]
  assign _T_87333 = _T_87332[13:0]; // @[Modules.scala 160:64:@34532.4]
  assign buffer_10_344 = $signed(_T_87333); // @[Modules.scala 160:64:@34533.4]
  assign buffer_10_76 = {{8{_T_85611[5]}},_T_85611}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_77 = {{9{_T_85618[4]}},_T_85618}; // @[Modules.scala 112:22:@8.4]
  assign _T_87338 = $signed(buffer_10_76) + $signed(buffer_10_77); // @[Modules.scala 160:64:@34539.4]
  assign _T_87339 = _T_87338[13:0]; // @[Modules.scala 160:64:@34540.4]
  assign buffer_10_346 = $signed(_T_87339); // @[Modules.scala 160:64:@34541.4]
  assign _T_87341 = $signed(buffer_2_81) + $signed(buffer_2_82); // @[Modules.scala 160:64:@34543.4]
  assign _T_87342 = _T_87341[13:0]; // @[Modules.scala 160:64:@34544.4]
  assign buffer_10_347 = $signed(_T_87342); // @[Modules.scala 160:64:@34545.4]
  assign buffer_10_80 = {{9{_T_85639[4]}},_T_85639}; // @[Modules.scala 112:22:@8.4]
  assign _T_87344 = $signed(buffer_10_80) + $signed(buffer_5_85); // @[Modules.scala 160:64:@34547.4]
  assign _T_87345 = _T_87344[13:0]; // @[Modules.scala 160:64:@34548.4]
  assign buffer_10_348 = $signed(_T_87345); // @[Modules.scala 160:64:@34549.4]
  assign buffer_10_84 = {{8{_T_85667[5]}},_T_85667}; // @[Modules.scala 112:22:@8.4]
  assign _T_87350 = $signed(buffer_10_84) + $signed(buffer_2_89); // @[Modules.scala 160:64:@34555.4]
  assign _T_87351 = _T_87350[13:0]; // @[Modules.scala 160:64:@34556.4]
  assign buffer_10_350 = $signed(_T_87351); // @[Modules.scala 160:64:@34557.4]
  assign _T_87353 = $signed(buffer_2_90) + $signed(buffer_6_90); // @[Modules.scala 160:64:@34559.4]
  assign _T_87354 = _T_87353[13:0]; // @[Modules.scala 160:64:@34560.4]
  assign buffer_10_351 = $signed(_T_87354); // @[Modules.scala 160:64:@34561.4]
  assign buffer_10_88 = {{8{_T_85695[5]}},_T_85695}; // @[Modules.scala 112:22:@8.4]
  assign _T_87356 = $signed(buffer_10_88) + $signed(buffer_2_93); // @[Modules.scala 160:64:@34563.4]
  assign _T_87357 = _T_87356[13:0]; // @[Modules.scala 160:64:@34564.4]
  assign buffer_10_352 = $signed(_T_87357); // @[Modules.scala 160:64:@34565.4]
  assign buffer_10_90 = {{9{_T_85709[4]}},_T_85709}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_91 = {{8{_T_85716[5]}},_T_85716}; // @[Modules.scala 112:22:@8.4]
  assign _T_87359 = $signed(buffer_10_90) + $signed(buffer_10_91); // @[Modules.scala 160:64:@34567.4]
  assign _T_87360 = _T_87359[13:0]; // @[Modules.scala 160:64:@34568.4]
  assign buffer_10_353 = $signed(_T_87360); // @[Modules.scala 160:64:@34569.4]
  assign buffer_10_93 = {{8{_T_85730[5]}},_T_85730}; // @[Modules.scala 112:22:@8.4]
  assign _T_87362 = $signed(buffer_6_96) + $signed(buffer_10_93); // @[Modules.scala 160:64:@34571.4]
  assign _T_87363 = _T_87362[13:0]; // @[Modules.scala 160:64:@34572.4]
  assign buffer_10_354 = $signed(_T_87363); // @[Modules.scala 160:64:@34573.4]
  assign _T_87365 = $signed(buffer_1_96) + $signed(buffer_2_99); // @[Modules.scala 160:64:@34575.4]
  assign _T_87366 = _T_87365[13:0]; // @[Modules.scala 160:64:@34576.4]
  assign buffer_10_355 = $signed(_T_87366); // @[Modules.scala 160:64:@34577.4]
  assign _T_87371 = $signed(buffer_9_104) + $signed(buffer_6_101); // @[Modules.scala 160:64:@34583.4]
  assign _T_87372 = _T_87371[13:0]; // @[Modules.scala 160:64:@34584.4]
  assign buffer_10_357 = $signed(_T_87372); // @[Modules.scala 160:64:@34585.4]
  assign buffer_10_100 = {{9{_T_85779[4]}},_T_85779}; // @[Modules.scala 112:22:@8.4]
  assign _T_87374 = $signed(buffer_10_100) + $signed(buffer_5_107); // @[Modules.scala 160:64:@34587.4]
  assign _T_87375 = _T_87374[13:0]; // @[Modules.scala 160:64:@34588.4]
  assign buffer_10_358 = $signed(_T_87375); // @[Modules.scala 160:64:@34589.4]
  assign buffer_10_104 = {{8{_T_85807[5]}},_T_85807}; // @[Modules.scala 112:22:@8.4]
  assign _T_87380 = $signed(buffer_10_104) + $signed(buffer_5_110); // @[Modules.scala 160:64:@34595.4]
  assign _T_87381 = _T_87380[13:0]; // @[Modules.scala 160:64:@34596.4]
  assign buffer_10_360 = $signed(_T_87381); // @[Modules.scala 160:64:@34597.4]
  assign buffer_10_106 = {{8{_T_85821[5]}},_T_85821}; // @[Modules.scala 112:22:@8.4]
  assign _T_87383 = $signed(buffer_10_106) + $signed(buffer_2_109); // @[Modules.scala 160:64:@34599.4]
  assign _T_87384 = _T_87383[13:0]; // @[Modules.scala 160:64:@34600.4]
  assign buffer_10_361 = $signed(_T_87384); // @[Modules.scala 160:64:@34601.4]
  assign buffer_10_109 = {{9{_T_85842[4]}},_T_85842}; // @[Modules.scala 112:22:@8.4]
  assign _T_87386 = $signed(buffer_2_110) + $signed(buffer_10_109); // @[Modules.scala 160:64:@34603.4]
  assign _T_87387 = _T_87386[13:0]; // @[Modules.scala 160:64:@34604.4]
  assign buffer_10_362 = $signed(_T_87387); // @[Modules.scala 160:64:@34605.4]
  assign _T_87389 = $signed(buffer_5_115) + $signed(buffer_1_112); // @[Modules.scala 160:64:@34607.4]
  assign _T_87390 = _T_87389[13:0]; // @[Modules.scala 160:64:@34608.4]
  assign buffer_10_363 = $signed(_T_87390); // @[Modules.scala 160:64:@34609.4]
  assign buffer_10_113 = {{9{_T_85870[4]}},_T_85870}; // @[Modules.scala 112:22:@8.4]
  assign _T_87392 = $signed(buffer_1_113) + $signed(buffer_10_113); // @[Modules.scala 160:64:@34611.4]
  assign _T_87393 = _T_87392[13:0]; // @[Modules.scala 160:64:@34612.4]
  assign buffer_10_364 = $signed(_T_87393); // @[Modules.scala 160:64:@34613.4]
  assign buffer_10_114 = {{9{_T_85877[4]}},_T_85877}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_115 = {{9{_T_85884[4]}},_T_85884}; // @[Modules.scala 112:22:@8.4]
  assign _T_87395 = $signed(buffer_10_114) + $signed(buffer_10_115); // @[Modules.scala 160:64:@34615.4]
  assign _T_87396 = _T_87395[13:0]; // @[Modules.scala 160:64:@34616.4]
  assign buffer_10_365 = $signed(_T_87396); // @[Modules.scala 160:64:@34617.4]
  assign _T_87398 = $signed(buffer_4_115) + $signed(buffer_2_119); // @[Modules.scala 160:64:@34619.4]
  assign _T_87399 = _T_87398[13:0]; // @[Modules.scala 160:64:@34620.4]
  assign buffer_10_366 = $signed(_T_87399); // @[Modules.scala 160:64:@34621.4]
  assign _T_87401 = $signed(buffer_2_120) + $signed(buffer_0_118); // @[Modules.scala 160:64:@34623.4]
  assign _T_87402 = _T_87401[13:0]; // @[Modules.scala 160:64:@34624.4]
  assign buffer_10_367 = $signed(_T_87402); // @[Modules.scala 160:64:@34625.4]
  assign buffer_10_121 = {{8{_T_85926[5]}},_T_85926}; // @[Modules.scala 112:22:@8.4]
  assign _T_87404 = $signed(buffer_0_119) + $signed(buffer_10_121); // @[Modules.scala 160:64:@34627.4]
  assign _T_87405 = _T_87404[13:0]; // @[Modules.scala 160:64:@34628.4]
  assign buffer_10_368 = $signed(_T_87405); // @[Modules.scala 160:64:@34629.4]
  assign buffer_10_123 = {{8{_T_85940[5]}},_T_85940}; // @[Modules.scala 112:22:@8.4]
  assign _T_87407 = $signed(buffer_5_124) + $signed(buffer_10_123); // @[Modules.scala 160:64:@34631.4]
  assign _T_87408 = _T_87407[13:0]; // @[Modules.scala 160:64:@34632.4]
  assign buffer_10_369 = $signed(_T_87408); // @[Modules.scala 160:64:@34633.4]
  assign _T_87410 = $signed(buffer_5_126) + $signed(buffer_1_126); // @[Modules.scala 160:64:@34635.4]
  assign _T_87411 = _T_87410[13:0]; // @[Modules.scala 160:64:@34636.4]
  assign buffer_10_370 = $signed(_T_87411); // @[Modules.scala 160:64:@34637.4]
  assign _T_87413 = $signed(buffer_5_128) + $signed(buffer_1_128); // @[Modules.scala 160:64:@34639.4]
  assign _T_87414 = _T_87413[13:0]; // @[Modules.scala 160:64:@34640.4]
  assign buffer_10_371 = $signed(_T_87414); // @[Modules.scala 160:64:@34641.4]
  assign buffer_10_130 = {{8{_T_85989[5]}},_T_85989}; // @[Modules.scala 112:22:@8.4]
  assign _T_87419 = $signed(buffer_10_130) + $signed(buffer_0_130); // @[Modules.scala 160:64:@34647.4]
  assign _T_87420 = _T_87419[13:0]; // @[Modules.scala 160:64:@34648.4]
  assign buffer_10_373 = $signed(_T_87420); // @[Modules.scala 160:64:@34649.4]
  assign buffer_10_132 = {{8{_T_86003[5]}},_T_86003}; // @[Modules.scala 112:22:@8.4]
  assign _T_87422 = $signed(buffer_10_132) + $signed(buffer_0_132); // @[Modules.scala 160:64:@34651.4]
  assign _T_87423 = _T_87422[13:0]; // @[Modules.scala 160:64:@34652.4]
  assign buffer_10_374 = $signed(_T_87423); // @[Modules.scala 160:64:@34653.4]
  assign buffer_10_134 = {{8{_T_86017[5]}},_T_86017}; // @[Modules.scala 112:22:@8.4]
  assign _T_87425 = $signed(buffer_10_134) + $signed(buffer_1_136); // @[Modules.scala 160:64:@34655.4]
  assign _T_87426 = _T_87425[13:0]; // @[Modules.scala 160:64:@34656.4]
  assign buffer_10_375 = $signed(_T_87426); // @[Modules.scala 160:64:@34657.4]
  assign buffer_10_137 = {{8{_T_86038[5]}},_T_86038}; // @[Modules.scala 112:22:@8.4]
  assign _T_87428 = $signed(buffer_4_133) + $signed(buffer_10_137); // @[Modules.scala 160:64:@34659.4]
  assign _T_87429 = _T_87428[13:0]; // @[Modules.scala 160:64:@34660.4]
  assign buffer_10_376 = $signed(_T_87429); // @[Modules.scala 160:64:@34661.4]
  assign _T_87434 = $signed(buffer_1_140) + $signed(buffer_6_144); // @[Modules.scala 160:64:@34667.4]
  assign _T_87435 = _T_87434[13:0]; // @[Modules.scala 160:64:@34668.4]
  assign buffer_10_378 = $signed(_T_87435); // @[Modules.scala 160:64:@34669.4]
  assign _T_87440 = $signed(buffer_0_143) + $signed(buffer_2_147); // @[Modules.scala 160:64:@34675.4]
  assign _T_87441 = _T_87440[13:0]; // @[Modules.scala 160:64:@34676.4]
  assign buffer_10_380 = $signed(_T_87441); // @[Modules.scala 160:64:@34677.4]
  assign buffer_10_147 = {{8{_T_86108[5]}},_T_86108}; // @[Modules.scala 112:22:@8.4]
  assign _T_87443 = $signed(buffer_3_152) + $signed(buffer_10_147); // @[Modules.scala 160:64:@34679.4]
  assign _T_87444 = _T_87443[13:0]; // @[Modules.scala 160:64:@34680.4]
  assign buffer_10_381 = $signed(_T_87444); // @[Modules.scala 160:64:@34681.4]
  assign buffer_10_150 = {{8{_T_86129[5]}},_T_86129}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_151 = {{8{_T_86136[5]}},_T_86136}; // @[Modules.scala 112:22:@8.4]
  assign _T_87449 = $signed(buffer_10_150) + $signed(buffer_10_151); // @[Modules.scala 160:64:@34687.4]
  assign _T_87450 = _T_87449[13:0]; // @[Modules.scala 160:64:@34688.4]
  assign buffer_10_383 = $signed(_T_87450); // @[Modules.scala 160:64:@34689.4]
  assign buffer_10_154 = {{9{_T_86157[4]}},_T_86157}; // @[Modules.scala 112:22:@8.4]
  assign _T_87455 = $signed(buffer_10_154) + $signed(buffer_0_152); // @[Modules.scala 160:64:@34695.4]
  assign _T_87456 = _T_87455[13:0]; // @[Modules.scala 160:64:@34696.4]
  assign buffer_10_385 = $signed(_T_87456); // @[Modules.scala 160:64:@34697.4]
  assign _T_87461 = $signed(buffer_8_153) + $signed(buffer_1_157); // @[Modules.scala 160:64:@34703.4]
  assign _T_87462 = _T_87461[13:0]; // @[Modules.scala 160:64:@34704.4]
  assign buffer_10_387 = $signed(_T_87462); // @[Modules.scala 160:64:@34705.4]
  assign buffer_10_161 = {{9{_T_86206[4]}},_T_86206}; // @[Modules.scala 112:22:@8.4]
  assign _T_87464 = $signed(buffer_8_155) + $signed(buffer_10_161); // @[Modules.scala 160:64:@34707.4]
  assign _T_87465 = _T_87464[13:0]; // @[Modules.scala 160:64:@34708.4]
  assign buffer_10_388 = $signed(_T_87465); // @[Modules.scala 160:64:@34709.4]
  assign buffer_10_164 = {{8{_T_86227[5]}},_T_86227}; // @[Modules.scala 112:22:@8.4]
  assign _T_87470 = $signed(buffer_10_164) + $signed(buffer_5_163); // @[Modules.scala 160:64:@34715.4]
  assign _T_87471 = _T_87470[13:0]; // @[Modules.scala 160:64:@34716.4]
  assign buffer_10_390 = $signed(_T_87471); // @[Modules.scala 160:64:@34717.4]
  assign _T_87473 = $signed(buffer_6_169) + $signed(buffer_5_165); // @[Modules.scala 160:64:@34719.4]
  assign _T_87474 = _T_87473[13:0]; // @[Modules.scala 160:64:@34720.4]
  assign buffer_10_391 = $signed(_T_87474); // @[Modules.scala 160:64:@34721.4]
  assign _T_87476 = $signed(buffer_5_166) + $signed(buffer_1_166); // @[Modules.scala 160:64:@34723.4]
  assign _T_87477 = _T_87476[13:0]; // @[Modules.scala 160:64:@34724.4]
  assign buffer_10_392 = $signed(_T_87477); // @[Modules.scala 160:64:@34725.4]
  assign buffer_10_170 = {{8{_T_86269[5]}},_T_86269}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_171 = {{8{_T_86276[5]}},_T_86276}; // @[Modules.scala 112:22:@8.4]
  assign _T_87479 = $signed(buffer_10_170) + $signed(buffer_10_171); // @[Modules.scala 160:64:@34727.4]
  assign _T_87480 = _T_87479[13:0]; // @[Modules.scala 160:64:@34728.4]
  assign buffer_10_393 = $signed(_T_87480); // @[Modules.scala 160:64:@34729.4]
  assign _T_87482 = $signed(buffer_2_173) + $signed(buffer_3_175); // @[Modules.scala 160:64:@34731.4]
  assign _T_87483 = _T_87482[13:0]; // @[Modules.scala 160:64:@34732.4]
  assign buffer_10_394 = $signed(_T_87483); // @[Modules.scala 160:64:@34733.4]
  assign _T_87488 = $signed(buffer_2_177) + $signed(buffer_7_176); // @[Modules.scala 160:64:@34739.4]
  assign _T_87489 = _T_87488[13:0]; // @[Modules.scala 160:64:@34740.4]
  assign buffer_10_396 = $signed(_T_87489); // @[Modules.scala 160:64:@34741.4]
  assign buffer_10_179 = {{8{_T_86332[5]}},_T_86332}; // @[Modules.scala 112:22:@8.4]
  assign _T_87491 = $signed(buffer_7_177) + $signed(buffer_10_179); // @[Modules.scala 160:64:@34743.4]
  assign _T_87492 = _T_87491[13:0]; // @[Modules.scala 160:64:@34744.4]
  assign buffer_10_397 = $signed(_T_87492); // @[Modules.scala 160:64:@34745.4]
  assign buffer_10_181 = {{8{_T_86346[5]}},_T_86346}; // @[Modules.scala 112:22:@8.4]
  assign _T_87494 = $signed(buffer_3_182) + $signed(buffer_10_181); // @[Modules.scala 160:64:@34747.4]
  assign _T_87495 = _T_87494[13:0]; // @[Modules.scala 160:64:@34748.4]
  assign buffer_10_398 = $signed(_T_87495); // @[Modules.scala 160:64:@34749.4]
  assign buffer_10_182 = {{8{_T_86353[5]}},_T_86353}; // @[Modules.scala 112:22:@8.4]
  assign _T_87497 = $signed(buffer_10_182) + $signed(buffer_0_178); // @[Modules.scala 160:64:@34751.4]
  assign _T_87498 = _T_87497[13:0]; // @[Modules.scala 160:64:@34752.4]
  assign buffer_10_399 = $signed(_T_87498); // @[Modules.scala 160:64:@34753.4]
  assign buffer_10_185 = {{8{_T_86374[5]}},_T_86374}; // @[Modules.scala 112:22:@8.4]
  assign _T_87500 = $signed(buffer_6_185) + $signed(buffer_10_185); // @[Modules.scala 160:64:@34755.4]
  assign _T_87501 = _T_87500[13:0]; // @[Modules.scala 160:64:@34756.4]
  assign buffer_10_400 = $signed(_T_87501); // @[Modules.scala 160:64:@34757.4]
  assign buffer_10_186 = {{9{_T_86381[4]}},_T_86381}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_187 = {{9{_T_86388[4]}},_T_86388}; // @[Modules.scala 112:22:@8.4]
  assign _T_87503 = $signed(buffer_10_186) + $signed(buffer_10_187); // @[Modules.scala 160:64:@34759.4]
  assign _T_87504 = _T_87503[13:0]; // @[Modules.scala 160:64:@34760.4]
  assign buffer_10_401 = $signed(_T_87504); // @[Modules.scala 160:64:@34761.4]
  assign buffer_10_188 = {{9{_T_86395[4]}},_T_86395}; // @[Modules.scala 112:22:@8.4]
  assign _T_87506 = $signed(buffer_10_188) + $signed(buffer_6_190); // @[Modules.scala 160:64:@34763.4]
  assign _T_87507 = _T_87506[13:0]; // @[Modules.scala 160:64:@34764.4]
  assign buffer_10_402 = $signed(_T_87507); // @[Modules.scala 160:64:@34765.4]
  assign buffer_10_191 = {{8{_T_86416[5]}},_T_86416}; // @[Modules.scala 112:22:@8.4]
  assign _T_87509 = $signed(buffer_0_183) + $signed(buffer_10_191); // @[Modules.scala 160:64:@34767.4]
  assign _T_87510 = _T_87509[13:0]; // @[Modules.scala 160:64:@34768.4]
  assign buffer_10_403 = $signed(_T_87510); // @[Modules.scala 160:64:@34769.4]
  assign _T_87512 = $signed(buffer_2_191) + $signed(buffer_1_187); // @[Modules.scala 160:64:@34771.4]
  assign _T_87513 = _T_87512[13:0]; // @[Modules.scala 160:64:@34772.4]
  assign buffer_10_404 = $signed(_T_87513); // @[Modules.scala 160:64:@34773.4]
  assign _T_87515 = $signed(buffer_3_197) + $signed(buffer_0_187); // @[Modules.scala 160:64:@34775.4]
  assign _T_87516 = _T_87515[13:0]; // @[Modules.scala 160:64:@34776.4]
  assign buffer_10_405 = $signed(_T_87516); // @[Modules.scala 160:64:@34777.4]
  assign buffer_10_197 = {{8{_T_86458[5]}},_T_86458}; // @[Modules.scala 112:22:@8.4]
  assign _T_87518 = $signed(buffer_0_188) + $signed(buffer_10_197); // @[Modules.scala 160:64:@34779.4]
  assign _T_87519 = _T_87518[13:0]; // @[Modules.scala 160:64:@34780.4]
  assign buffer_10_406 = $signed(_T_87519); // @[Modules.scala 160:64:@34781.4]
  assign buffer_10_198 = {{9{_T_86465[4]}},_T_86465}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_199 = {{9{_T_86472[4]}},_T_86472}; // @[Modules.scala 112:22:@8.4]
  assign _T_87521 = $signed(buffer_10_198) + $signed(buffer_10_199); // @[Modules.scala 160:64:@34783.4]
  assign _T_87522 = _T_87521[13:0]; // @[Modules.scala 160:64:@34784.4]
  assign buffer_10_407 = $signed(_T_87522); // @[Modules.scala 160:64:@34785.4]
  assign buffer_10_201 = {{8{_T_86486[5]}},_T_86486}; // @[Modules.scala 112:22:@8.4]
  assign _T_87524 = $signed(buffer_5_196) + $signed(buffer_10_201); // @[Modules.scala 160:64:@34787.4]
  assign _T_87525 = _T_87524[13:0]; // @[Modules.scala 160:64:@34788.4]
  assign buffer_10_408 = $signed(_T_87525); // @[Modules.scala 160:64:@34789.4]
  assign buffer_10_202 = {{9{_T_86493[4]}},_T_86493}; // @[Modules.scala 112:22:@8.4]
  assign _T_87527 = $signed(buffer_10_202) + $signed(buffer_7_204); // @[Modules.scala 160:64:@34791.4]
  assign _T_87528 = _T_87527[13:0]; // @[Modules.scala 160:64:@34792.4]
  assign buffer_10_409 = $signed(_T_87528); // @[Modules.scala 160:64:@34793.4]
  assign _T_87530 = $signed(buffer_4_191) + $signed(buffer_2_204); // @[Modules.scala 160:64:@34795.4]
  assign _T_87531 = _T_87530[13:0]; // @[Modules.scala 160:64:@34796.4]
  assign buffer_10_410 = $signed(_T_87531); // @[Modules.scala 160:64:@34797.4]
  assign _T_87533 = $signed(buffer_0_199) + $signed(buffer_0_200); // @[Modules.scala 160:64:@34799.4]
  assign _T_87534 = _T_87533[13:0]; // @[Modules.scala 160:64:@34800.4]
  assign buffer_10_411 = $signed(_T_87534); // @[Modules.scala 160:64:@34801.4]
  assign _T_87536 = $signed(buffer_0_201) + $signed(buffer_9_214); // @[Modules.scala 160:64:@34803.4]
  assign _T_87537 = _T_87536[13:0]; // @[Modules.scala 160:64:@34804.4]
  assign buffer_10_412 = $signed(_T_87537); // @[Modules.scala 160:64:@34805.4]
  assign buffer_10_213 = {{9{_T_86570[4]}},_T_86570}; // @[Modules.scala 112:22:@8.4]
  assign _T_87542 = $signed(buffer_2_211) + $signed(buffer_10_213); // @[Modules.scala 160:64:@34811.4]
  assign _T_87543 = _T_87542[13:0]; // @[Modules.scala 160:64:@34812.4]
  assign buffer_10_414 = $signed(_T_87543); // @[Modules.scala 160:64:@34813.4]
  assign buffer_10_219 = {{8{_T_86612[5]}},_T_86612}; // @[Modules.scala 112:22:@8.4]
  assign _T_87551 = $signed(buffer_0_212) + $signed(buffer_10_219); // @[Modules.scala 160:64:@34823.4]
  assign _T_87552 = _T_87551[13:0]; // @[Modules.scala 160:64:@34824.4]
  assign buffer_10_417 = $signed(_T_87552); // @[Modules.scala 160:64:@34825.4]
  assign buffer_10_221 = {{8{_T_86626[5]}},_T_86626}; // @[Modules.scala 112:22:@8.4]
  assign _T_87554 = $signed(buffer_6_224) + $signed(buffer_10_221); // @[Modules.scala 160:64:@34827.4]
  assign _T_87555 = _T_87554[13:0]; // @[Modules.scala 160:64:@34828.4]
  assign buffer_10_418 = $signed(_T_87555); // @[Modules.scala 160:64:@34829.4]
  assign buffer_10_226 = {{8{_T_86661[5]}},_T_86661}; // @[Modules.scala 112:22:@8.4]
  assign _T_87563 = $signed(buffer_10_226) + $signed(buffer_7_231); // @[Modules.scala 160:64:@34839.4]
  assign _T_87564 = _T_87563[13:0]; // @[Modules.scala 160:64:@34840.4]
  assign buffer_10_421 = $signed(_T_87564); // @[Modules.scala 160:64:@34841.4]
  assign buffer_10_229 = {{8{_T_86682[5]}},_T_86682}; // @[Modules.scala 112:22:@8.4]
  assign _T_87566 = $signed(buffer_7_232) + $signed(buffer_10_229); // @[Modules.scala 160:64:@34843.4]
  assign _T_87567 = _T_87566[13:0]; // @[Modules.scala 160:64:@34844.4]
  assign buffer_10_422 = $signed(_T_87567); // @[Modules.scala 160:64:@34845.4]
  assign buffer_10_230 = {{9{_T_86689[4]}},_T_86689}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_231 = {{8{_T_86696[5]}},_T_86696}; // @[Modules.scala 112:22:@8.4]
  assign _T_87569 = $signed(buffer_10_230) + $signed(buffer_10_231); // @[Modules.scala 160:64:@34847.4]
  assign _T_87570 = _T_87569[13:0]; // @[Modules.scala 160:64:@34848.4]
  assign buffer_10_423 = $signed(_T_87570); // @[Modules.scala 160:64:@34849.4]
  assign buffer_10_233 = {{8{_T_86710[5]}},_T_86710}; // @[Modules.scala 112:22:@8.4]
  assign _T_87572 = $signed(buffer_0_226) + $signed(buffer_10_233); // @[Modules.scala 160:64:@34851.4]
  assign _T_87573 = _T_87572[13:0]; // @[Modules.scala 160:64:@34852.4]
  assign buffer_10_424 = $signed(_T_87573); // @[Modules.scala 160:64:@34853.4]
  assign _T_87575 = $signed(buffer_5_235) + $signed(buffer_4_223); // @[Modules.scala 160:64:@34855.4]
  assign _T_87576 = _T_87575[13:0]; // @[Modules.scala 160:64:@34856.4]
  assign buffer_10_425 = $signed(_T_87576); // @[Modules.scala 160:64:@34857.4]
  assign buffer_10_237 = {{8{_T_86738[5]}},_T_86738}; // @[Modules.scala 112:22:@8.4]
  assign _T_87578 = $signed(buffer_2_236) + $signed(buffer_10_237); // @[Modules.scala 160:64:@34859.4]
  assign _T_87579 = _T_87578[13:0]; // @[Modules.scala 160:64:@34860.4]
  assign buffer_10_426 = $signed(_T_87579); // @[Modules.scala 160:64:@34861.4]
  assign _T_87581 = $signed(buffer_1_233) + $signed(buffer_6_244); // @[Modules.scala 160:64:@34863.4]
  assign _T_87582 = _T_87581[13:0]; // @[Modules.scala 160:64:@34864.4]
  assign buffer_10_427 = $signed(_T_87582); // @[Modules.scala 160:64:@34865.4]
  assign buffer_10_240 = {{9{_T_86759[4]}},_T_86759}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_241 = {{8{_T_86766[5]}},_T_86766}; // @[Modules.scala 112:22:@8.4]
  assign _T_87584 = $signed(buffer_10_240) + $signed(buffer_10_241); // @[Modules.scala 160:64:@34867.4]
  assign _T_87585 = _T_87584[13:0]; // @[Modules.scala 160:64:@34868.4]
  assign buffer_10_428 = $signed(_T_87585); // @[Modules.scala 160:64:@34869.4]
  assign _T_87587 = $signed(buffer_5_246) + $signed(buffer_6_249); // @[Modules.scala 160:64:@34871.4]
  assign _T_87588 = _T_87587[13:0]; // @[Modules.scala 160:64:@34872.4]
  assign buffer_10_429 = $signed(_T_87588); // @[Modules.scala 160:64:@34873.4]
  assign buffer_10_244 = {{8{_T_86787[5]}},_T_86787}; // @[Modules.scala 112:22:@8.4]
  assign _T_87590 = $signed(buffer_10_244) + $signed(buffer_7_250); // @[Modules.scala 160:64:@34875.4]
  assign _T_87591 = _T_87590[13:0]; // @[Modules.scala 160:64:@34876.4]
  assign buffer_10_430 = $signed(_T_87591); // @[Modules.scala 160:64:@34877.4]
  assign _T_87593 = $signed(buffer_2_248) + $signed(buffer_3_251); // @[Modules.scala 160:64:@34879.4]
  assign _T_87594 = _T_87593[13:0]; // @[Modules.scala 160:64:@34880.4]
  assign buffer_10_431 = $signed(_T_87594); // @[Modules.scala 160:64:@34881.4]
  assign buffer_10_251 = {{8{_T_86836[5]}},_T_86836}; // @[Modules.scala 112:22:@8.4]
  assign _T_87599 = $signed(buffer_0_243) + $signed(buffer_10_251); // @[Modules.scala 160:64:@34887.4]
  assign _T_87600 = _T_87599[13:0]; // @[Modules.scala 160:64:@34888.4]
  assign buffer_10_433 = $signed(_T_87600); // @[Modules.scala 160:64:@34889.4]
  assign buffer_10_252 = {{9{_T_86843[4]}},_T_86843}; // @[Modules.scala 112:22:@8.4]
  assign _T_87602 = $signed(buffer_10_252) + $signed(buffer_3_257); // @[Modules.scala 160:64:@34891.4]
  assign _T_87603 = _T_87602[13:0]; // @[Modules.scala 160:64:@34892.4]
  assign buffer_10_434 = $signed(_T_87603); // @[Modules.scala 160:64:@34893.4]
  assign buffer_10_255 = {{8{_T_86864[5]}},_T_86864}; // @[Modules.scala 112:22:@8.4]
  assign _T_87605 = $signed(buffer_6_259) + $signed(buffer_10_255); // @[Modules.scala 160:64:@34895.4]
  assign _T_87606 = _T_87605[13:0]; // @[Modules.scala 160:64:@34896.4]
  assign buffer_10_435 = $signed(_T_87606); // @[Modules.scala 160:64:@34897.4]
  assign buffer_10_256 = {{9{_T_86871[4]}},_T_86871}; // @[Modules.scala 112:22:@8.4]
  assign _T_87608 = $signed(buffer_10_256) + $signed(buffer_2_258); // @[Modules.scala 160:64:@34899.4]
  assign _T_87609 = _T_87608[13:0]; // @[Modules.scala 160:64:@34900.4]
  assign buffer_10_436 = $signed(_T_87609); // @[Modules.scala 160:64:@34901.4]
  assign buffer_10_258 = {{9{_T_86885[4]}},_T_86885}; // @[Modules.scala 112:22:@8.4]
  assign _T_87611 = $signed(buffer_10_258) + $signed(buffer_0_254); // @[Modules.scala 160:64:@34903.4]
  assign _T_87612 = _T_87611[13:0]; // @[Modules.scala 160:64:@34904.4]
  assign buffer_10_437 = $signed(_T_87612); // @[Modules.scala 160:64:@34905.4]
  assign buffer_10_262 = {{8{_T_86913[5]}},_T_86913}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_263 = {{8{_T_86920[5]}},_T_86920}; // @[Modules.scala 112:22:@8.4]
  assign _T_87617 = $signed(buffer_10_262) + $signed(buffer_10_263); // @[Modules.scala 160:64:@34911.4]
  assign _T_87618 = _T_87617[13:0]; // @[Modules.scala 160:64:@34912.4]
  assign buffer_10_439 = $signed(_T_87618); // @[Modules.scala 160:64:@34913.4]
  assign _T_87620 = $signed(buffer_8_266) + $signed(buffer_7_268); // @[Modules.scala 160:64:@34915.4]
  assign _T_87621 = _T_87620[13:0]; // @[Modules.scala 160:64:@34916.4]
  assign buffer_10_440 = $signed(_T_87621); // @[Modules.scala 160:64:@34917.4]
  assign buffer_10_271 = {{8{_T_86976[5]}},_T_86976}; // @[Modules.scala 112:22:@8.4]
  assign _T_87629 = $signed(buffer_3_274) + $signed(buffer_10_271); // @[Modules.scala 160:64:@34927.4]
  assign _T_87630 = _T_87629[13:0]; // @[Modules.scala 160:64:@34928.4]
  assign buffer_10_443 = $signed(_T_87630); // @[Modules.scala 160:64:@34929.4]
  assign buffer_10_272 = {{8{_T_86983[5]}},_T_86983}; // @[Modules.scala 112:22:@8.4]
  assign _T_87632 = $signed(buffer_10_272) + $signed(buffer_1_268); // @[Modules.scala 160:64:@34931.4]
  assign _T_87633 = _T_87632[13:0]; // @[Modules.scala 160:64:@34932.4]
  assign buffer_10_444 = $signed(_T_87633); // @[Modules.scala 160:64:@34933.4]
  assign _T_87635 = $signed(buffer_3_279) + $signed(buffer_3_280); // @[Modules.scala 160:64:@34935.4]
  assign _T_87636 = _T_87635[13:0]; // @[Modules.scala 160:64:@34936.4]
  assign buffer_10_445 = $signed(_T_87636); // @[Modules.scala 160:64:@34937.4]
  assign buffer_10_276 = {{8{_T_87011[5]}},_T_87011}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_277 = {{8{_T_87018[5]}},_T_87018}; // @[Modules.scala 112:22:@8.4]
  assign _T_87638 = $signed(buffer_10_276) + $signed(buffer_10_277); // @[Modules.scala 160:64:@34939.4]
  assign _T_87639 = _T_87638[13:0]; // @[Modules.scala 160:64:@34940.4]
  assign buffer_10_446 = $signed(_T_87639); // @[Modules.scala 160:64:@34941.4]
  assign buffer_10_278 = {{9{_T_87025[4]}},_T_87025}; // @[Modules.scala 112:22:@8.4]
  assign _T_87641 = $signed(buffer_10_278) + $signed(buffer_3_284); // @[Modules.scala 160:64:@34943.4]
  assign _T_87642 = _T_87641[13:0]; // @[Modules.scala 160:64:@34944.4]
  assign buffer_10_447 = $signed(_T_87642); // @[Modules.scala 160:64:@34945.4]
  assign _T_87644 = $signed(buffer_3_285) + $signed(buffer_3_286); // @[Modules.scala 160:64:@34947.4]
  assign _T_87645 = _T_87644[13:0]; // @[Modules.scala 160:64:@34948.4]
  assign buffer_10_448 = $signed(_T_87645); // @[Modules.scala 160:64:@34949.4]
  assign buffer_10_287 = {{8{_T_87088[5]}},_T_87088}; // @[Modules.scala 112:22:@8.4]
  assign _T_87653 = $signed(buffer_1_281) + $signed(buffer_10_287); // @[Modules.scala 160:64:@34959.4]
  assign _T_87654 = _T_87653[13:0]; // @[Modules.scala 160:64:@34960.4]
  assign buffer_10_451 = $signed(_T_87654); // @[Modules.scala 160:64:@34961.4]
  assign _T_87656 = $signed(buffer_6_294) + $signed(buffer_4_279); // @[Modules.scala 160:64:@34963.4]
  assign _T_87657 = _T_87656[13:0]; // @[Modules.scala 160:64:@34964.4]
  assign buffer_10_452 = $signed(_T_87657); // @[Modules.scala 160:64:@34965.4]
  assign buffer_10_291 = {{8{_T_87116[5]}},_T_87116}; // @[Modules.scala 112:22:@8.4]
  assign _T_87659 = $signed(buffer_3_294) + $signed(buffer_10_291); // @[Modules.scala 160:64:@34967.4]
  assign _T_87660 = _T_87659[13:0]; // @[Modules.scala 160:64:@34968.4]
  assign buffer_10_453 = $signed(_T_87660); // @[Modules.scala 160:64:@34969.4]
  assign buffer_10_292 = {{8{_T_87123[5]}},_T_87123}; // @[Modules.scala 112:22:@8.4]
  assign _T_87662 = $signed(buffer_10_292) + $signed(buffer_4_284); // @[Modules.scala 160:64:@34971.4]
  assign _T_87663 = _T_87662[13:0]; // @[Modules.scala 160:64:@34972.4]
  assign buffer_10_454 = $signed(_T_87663); // @[Modules.scala 160:64:@34973.4]
  assign _T_87665 = $signed(buffer_4_285) + $signed(buffer_4_286); // @[Modules.scala 160:64:@34975.4]
  assign _T_87666 = _T_87665[13:0]; // @[Modules.scala 160:64:@34976.4]
  assign buffer_10_455 = $signed(_T_87666); // @[Modules.scala 160:64:@34977.4]
  assign _T_87668 = $signed(buffer_4_287) + $signed(buffer_4_288); // @[Modules.scala 160:64:@34979.4]
  assign _T_87669 = _T_87668[13:0]; // @[Modules.scala 160:64:@34980.4]
  assign buffer_10_456 = $signed(_T_87669); // @[Modules.scala 160:64:@34981.4]
  assign buffer_10_298 = {{9{_T_87165[4]}},_T_87165}; // @[Modules.scala 112:22:@8.4]
  assign buffer_10_299 = {{8{_T_87172[5]}},_T_87172}; // @[Modules.scala 112:22:@8.4]
  assign _T_87671 = $signed(buffer_10_298) + $signed(buffer_10_299); // @[Modules.scala 160:64:@34983.4]
  assign _T_87672 = _T_87671[13:0]; // @[Modules.scala 160:64:@34984.4]
  assign buffer_10_457 = $signed(_T_87672); // @[Modules.scala 160:64:@34985.4]
  assign buffer_10_300 = {{8{_T_87179[5]}},_T_87179}; // @[Modules.scala 112:22:@8.4]
  assign _T_87674 = $signed(buffer_10_300) + $signed(buffer_2_304); // @[Modules.scala 160:64:@34987.4]
  assign _T_87675 = _T_87674[13:0]; // @[Modules.scala 160:64:@34988.4]
  assign buffer_10_458 = $signed(_T_87675); // @[Modules.scala 160:64:@34989.4]
  assign _T_87677 = $signed(buffer_2_305) + $signed(buffer_9_310); // @[Modules.scala 160:64:@34991.4]
  assign _T_87678 = _T_87677[13:0]; // @[Modules.scala 160:64:@34992.4]
  assign buffer_10_459 = $signed(_T_87678); // @[Modules.scala 160:64:@34993.4]
  assign _T_87686 = $signed(buffer_10_308) + $signed(buffer_10_309); // @[Modules.scala 160:64:@35003.4]
  assign _T_87687 = _T_87686[13:0]; // @[Modules.scala 160:64:@35004.4]
  assign buffer_10_462 = $signed(_T_87687); // @[Modules.scala 160:64:@35005.4]
  assign _T_87689 = $signed(buffer_0_304) + $signed(buffer_10_311); // @[Modules.scala 160:64:@35007.4]
  assign _T_87690 = _T_87689[13:0]; // @[Modules.scala 160:64:@35008.4]
  assign buffer_10_463 = $signed(_T_87690); // @[Modules.scala 160:64:@35009.4]
  assign _T_87692 = $signed(buffer_10_312) + $signed(buffer_10_313); // @[Modules.scala 160:64:@35011.4]
  assign _T_87693 = _T_87692[13:0]; // @[Modules.scala 160:64:@35012.4]
  assign buffer_10_464 = $signed(_T_87693); // @[Modules.scala 160:64:@35013.4]
  assign _T_87701 = $signed(buffer_10_318) + $signed(buffer_10_319); // @[Modules.scala 160:64:@35023.4]
  assign _T_87702 = _T_87701[13:0]; // @[Modules.scala 160:64:@35024.4]
  assign buffer_10_467 = $signed(_T_87702); // @[Modules.scala 160:64:@35025.4]
  assign _T_87704 = $signed(buffer_10_320) + $signed(buffer_10_321); // @[Modules.scala 160:64:@35027.4]
  assign _T_87705 = _T_87704[13:0]; // @[Modules.scala 160:64:@35028.4]
  assign buffer_10_468 = $signed(_T_87705); // @[Modules.scala 160:64:@35029.4]
  assign _T_87707 = $signed(buffer_10_322) + $signed(buffer_2_324); // @[Modules.scala 160:64:@35031.4]
  assign _T_87708 = _T_87707[13:0]; // @[Modules.scala 160:64:@35032.4]
  assign buffer_10_469 = $signed(_T_87708); // @[Modules.scala 160:64:@35033.4]
  assign _T_87710 = $signed(buffer_10_324) + $signed(buffer_10_325); // @[Modules.scala 160:64:@35035.4]
  assign _T_87711 = _T_87710[13:0]; // @[Modules.scala 160:64:@35036.4]
  assign buffer_10_470 = $signed(_T_87711); // @[Modules.scala 160:64:@35037.4]
  assign _T_87713 = $signed(buffer_10_326) + $signed(buffer_10_327); // @[Modules.scala 160:64:@35039.4]
  assign _T_87714 = _T_87713[13:0]; // @[Modules.scala 160:64:@35040.4]
  assign buffer_10_471 = $signed(_T_87714); // @[Modules.scala 160:64:@35041.4]
  assign _T_87716 = $signed(buffer_10_328) + $signed(buffer_10_329); // @[Modules.scala 160:64:@35043.4]
  assign _T_87717 = _T_87716[13:0]; // @[Modules.scala 160:64:@35044.4]
  assign buffer_10_472 = $signed(_T_87717); // @[Modules.scala 160:64:@35045.4]
  assign _T_87719 = $signed(buffer_0_324) + $signed(buffer_10_331); // @[Modules.scala 160:64:@35047.4]
  assign _T_87720 = _T_87719[13:0]; // @[Modules.scala 160:64:@35048.4]
  assign buffer_10_473 = $signed(_T_87720); // @[Modules.scala 160:64:@35049.4]
  assign _T_87722 = $signed(buffer_10_332) + $signed(buffer_10_333); // @[Modules.scala 160:64:@35051.4]
  assign _T_87723 = _T_87722[13:0]; // @[Modules.scala 160:64:@35052.4]
  assign buffer_10_474 = $signed(_T_87723); // @[Modules.scala 160:64:@35053.4]
  assign _T_87728 = $signed(buffer_10_336) + $signed(buffer_10_337); // @[Modules.scala 160:64:@35059.4]
  assign _T_87729 = _T_87728[13:0]; // @[Modules.scala 160:64:@35060.4]
  assign buffer_10_476 = $signed(_T_87729); // @[Modules.scala 160:64:@35061.4]
  assign _T_87731 = $signed(buffer_10_338) + $signed(buffer_10_339); // @[Modules.scala 160:64:@35063.4]
  assign _T_87732 = _T_87731[13:0]; // @[Modules.scala 160:64:@35064.4]
  assign buffer_10_477 = $signed(_T_87732); // @[Modules.scala 160:64:@35065.4]
  assign _T_87734 = $signed(buffer_10_340) + $signed(buffer_10_341); // @[Modules.scala 160:64:@35067.4]
  assign _T_87735 = _T_87734[13:0]; // @[Modules.scala 160:64:@35068.4]
  assign buffer_10_478 = $signed(_T_87735); // @[Modules.scala 160:64:@35069.4]
  assign _T_87737 = $signed(buffer_10_342) + $signed(buffer_10_343); // @[Modules.scala 160:64:@35071.4]
  assign _T_87738 = _T_87737[13:0]; // @[Modules.scala 160:64:@35072.4]
  assign buffer_10_479 = $signed(_T_87738); // @[Modules.scala 160:64:@35073.4]
  assign _T_87740 = $signed(buffer_10_344) + $signed(buffer_1_342); // @[Modules.scala 160:64:@35075.4]
  assign _T_87741 = _T_87740[13:0]; // @[Modules.scala 160:64:@35076.4]
  assign buffer_10_480 = $signed(_T_87741); // @[Modules.scala 160:64:@35077.4]
  assign _T_87743 = $signed(buffer_10_346) + $signed(buffer_10_347); // @[Modules.scala 160:64:@35079.4]
  assign _T_87744 = _T_87743[13:0]; // @[Modules.scala 160:64:@35080.4]
  assign buffer_10_481 = $signed(_T_87744); // @[Modules.scala 160:64:@35081.4]
  assign _T_87746 = $signed(buffer_10_348) + $signed(buffer_1_346); // @[Modules.scala 160:64:@35083.4]
  assign _T_87747 = _T_87746[13:0]; // @[Modules.scala 160:64:@35084.4]
  assign buffer_10_482 = $signed(_T_87747); // @[Modules.scala 160:64:@35085.4]
  assign _T_87749 = $signed(buffer_10_350) + $signed(buffer_10_351); // @[Modules.scala 160:64:@35087.4]
  assign _T_87750 = _T_87749[13:0]; // @[Modules.scala 160:64:@35088.4]
  assign buffer_10_483 = $signed(_T_87750); // @[Modules.scala 160:64:@35089.4]
  assign _T_87752 = $signed(buffer_10_352) + $signed(buffer_10_353); // @[Modules.scala 160:64:@35091.4]
  assign _T_87753 = _T_87752[13:0]; // @[Modules.scala 160:64:@35092.4]
  assign buffer_10_484 = $signed(_T_87753); // @[Modules.scala 160:64:@35093.4]
  assign _T_87755 = $signed(buffer_10_354) + $signed(buffer_10_355); // @[Modules.scala 160:64:@35095.4]
  assign _T_87756 = _T_87755[13:0]; // @[Modules.scala 160:64:@35096.4]
  assign buffer_10_485 = $signed(_T_87756); // @[Modules.scala 160:64:@35097.4]
  assign _T_87758 = $signed(buffer_9_365) + $signed(buffer_10_357); // @[Modules.scala 160:64:@35099.4]
  assign _T_87759 = _T_87758[13:0]; // @[Modules.scala 160:64:@35100.4]
  assign buffer_10_486 = $signed(_T_87759); // @[Modules.scala 160:64:@35101.4]
  assign _T_87761 = $signed(buffer_10_358) + $signed(buffer_4_351); // @[Modules.scala 160:64:@35103.4]
  assign _T_87762 = _T_87761[13:0]; // @[Modules.scala 160:64:@35104.4]
  assign buffer_10_487 = $signed(_T_87762); // @[Modules.scala 160:64:@35105.4]
  assign _T_87764 = $signed(buffer_10_360) + $signed(buffer_10_361); // @[Modules.scala 160:64:@35107.4]
  assign _T_87765 = _T_87764[13:0]; // @[Modules.scala 160:64:@35108.4]
  assign buffer_10_488 = $signed(_T_87765); // @[Modules.scala 160:64:@35109.4]
  assign _T_87767 = $signed(buffer_10_362) + $signed(buffer_10_363); // @[Modules.scala 160:64:@35111.4]
  assign _T_87768 = _T_87767[13:0]; // @[Modules.scala 160:64:@35112.4]
  assign buffer_10_489 = $signed(_T_87768); // @[Modules.scala 160:64:@35113.4]
  assign _T_87770 = $signed(buffer_10_364) + $signed(buffer_10_365); // @[Modules.scala 160:64:@35115.4]
  assign _T_87771 = _T_87770[13:0]; // @[Modules.scala 160:64:@35116.4]
  assign buffer_10_490 = $signed(_T_87771); // @[Modules.scala 160:64:@35117.4]
  assign _T_87773 = $signed(buffer_10_366) + $signed(buffer_10_367); // @[Modules.scala 160:64:@35119.4]
  assign _T_87774 = _T_87773[13:0]; // @[Modules.scala 160:64:@35120.4]
  assign buffer_10_491 = $signed(_T_87774); // @[Modules.scala 160:64:@35121.4]
  assign _T_87776 = $signed(buffer_10_368) + $signed(buffer_10_369); // @[Modules.scala 160:64:@35123.4]
  assign _T_87777 = _T_87776[13:0]; // @[Modules.scala 160:64:@35124.4]
  assign buffer_10_492 = $signed(_T_87777); // @[Modules.scala 160:64:@35125.4]
  assign _T_87779 = $signed(buffer_10_370) + $signed(buffer_10_371); // @[Modules.scala 160:64:@35127.4]
  assign _T_87780 = _T_87779[13:0]; // @[Modules.scala 160:64:@35128.4]
  assign buffer_10_493 = $signed(_T_87780); // @[Modules.scala 160:64:@35129.4]
  assign _T_87782 = $signed(buffer_3_381) + $signed(buffer_10_373); // @[Modules.scala 160:64:@35131.4]
  assign _T_87783 = _T_87782[13:0]; // @[Modules.scala 160:64:@35132.4]
  assign buffer_10_494 = $signed(_T_87783); // @[Modules.scala 160:64:@35133.4]
  assign _T_87785 = $signed(buffer_10_374) + $signed(buffer_10_375); // @[Modules.scala 160:64:@35135.4]
  assign _T_87786 = _T_87785[13:0]; // @[Modules.scala 160:64:@35136.4]
  assign buffer_10_495 = $signed(_T_87786); // @[Modules.scala 160:64:@35137.4]
  assign _T_87788 = $signed(buffer_10_376) + $signed(buffer_1_373); // @[Modules.scala 160:64:@35139.4]
  assign _T_87789 = _T_87788[13:0]; // @[Modules.scala 160:64:@35140.4]
  assign buffer_10_496 = $signed(_T_87789); // @[Modules.scala 160:64:@35141.4]
  assign _T_87791 = $signed(buffer_10_378) + $signed(buffer_7_379); // @[Modules.scala 160:64:@35143.4]
  assign _T_87792 = _T_87791[13:0]; // @[Modules.scala 160:64:@35144.4]
  assign buffer_10_497 = $signed(_T_87792); // @[Modules.scala 160:64:@35145.4]
  assign _T_87794 = $signed(buffer_10_380) + $signed(buffer_10_381); // @[Modules.scala 160:64:@35147.4]
  assign _T_87795 = _T_87794[13:0]; // @[Modules.scala 160:64:@35148.4]
  assign buffer_10_498 = $signed(_T_87795); // @[Modules.scala 160:64:@35149.4]
  assign _T_87797 = $signed(buffer_3_391) + $signed(buffer_10_383); // @[Modules.scala 160:64:@35151.4]
  assign _T_87798 = _T_87797[13:0]; // @[Modules.scala 160:64:@35152.4]
  assign buffer_10_499 = $signed(_T_87798); // @[Modules.scala 160:64:@35153.4]
  assign _T_87800 = $signed(buffer_5_389) + $signed(buffer_10_385); // @[Modules.scala 160:64:@35155.4]
  assign _T_87801 = _T_87800[13:0]; // @[Modules.scala 160:64:@35156.4]
  assign buffer_10_500 = $signed(_T_87801); // @[Modules.scala 160:64:@35157.4]
  assign _T_87803 = $signed(buffer_4_375) + $signed(buffer_10_387); // @[Modules.scala 160:64:@35159.4]
  assign _T_87804 = _T_87803[13:0]; // @[Modules.scala 160:64:@35160.4]
  assign buffer_10_501 = $signed(_T_87804); // @[Modules.scala 160:64:@35161.4]
  assign _T_87806 = $signed(buffer_10_388) + $signed(buffer_7_389); // @[Modules.scala 160:64:@35163.4]
  assign _T_87807 = _T_87806[13:0]; // @[Modules.scala 160:64:@35164.4]
  assign buffer_10_502 = $signed(_T_87807); // @[Modules.scala 160:64:@35165.4]
  assign _T_87809 = $signed(buffer_10_390) + $signed(buffer_10_391); // @[Modules.scala 160:64:@35167.4]
  assign _T_87810 = _T_87809[13:0]; // @[Modules.scala 160:64:@35168.4]
  assign buffer_10_503 = $signed(_T_87810); // @[Modules.scala 160:64:@35169.4]
  assign _T_87812 = $signed(buffer_10_392) + $signed(buffer_10_393); // @[Modules.scala 160:64:@35171.4]
  assign _T_87813 = _T_87812[13:0]; // @[Modules.scala 160:64:@35172.4]
  assign buffer_10_504 = $signed(_T_87813); // @[Modules.scala 160:64:@35173.4]
  assign _T_87815 = $signed(buffer_10_394) + $signed(buffer_3_402); // @[Modules.scala 160:64:@35175.4]
  assign _T_87816 = _T_87815[13:0]; // @[Modules.scala 160:64:@35176.4]
  assign buffer_10_505 = $signed(_T_87816); // @[Modules.scala 160:64:@35177.4]
  assign _T_87818 = $signed(buffer_10_396) + $signed(buffer_10_397); // @[Modules.scala 160:64:@35179.4]
  assign _T_87819 = _T_87818[13:0]; // @[Modules.scala 160:64:@35180.4]
  assign buffer_10_506 = $signed(_T_87819); // @[Modules.scala 160:64:@35181.4]
  assign _T_87821 = $signed(buffer_10_398) + $signed(buffer_10_399); // @[Modules.scala 160:64:@35183.4]
  assign _T_87822 = _T_87821[13:0]; // @[Modules.scala 160:64:@35184.4]
  assign buffer_10_507 = $signed(_T_87822); // @[Modules.scala 160:64:@35185.4]
  assign _T_87824 = $signed(buffer_10_400) + $signed(buffer_10_401); // @[Modules.scala 160:64:@35187.4]
  assign _T_87825 = _T_87824[13:0]; // @[Modules.scala 160:64:@35188.4]
  assign buffer_10_508 = $signed(_T_87825); // @[Modules.scala 160:64:@35189.4]
  assign _T_87827 = $signed(buffer_10_402) + $signed(buffer_10_403); // @[Modules.scala 160:64:@35191.4]
  assign _T_87828 = _T_87827[13:0]; // @[Modules.scala 160:64:@35192.4]
  assign buffer_10_509 = $signed(_T_87828); // @[Modules.scala 160:64:@35193.4]
  assign _T_87830 = $signed(buffer_10_404) + $signed(buffer_10_405); // @[Modules.scala 160:64:@35195.4]
  assign _T_87831 = _T_87830[13:0]; // @[Modules.scala 160:64:@35196.4]
  assign buffer_10_510 = $signed(_T_87831); // @[Modules.scala 160:64:@35197.4]
  assign _T_87833 = $signed(buffer_10_406) + $signed(buffer_10_407); // @[Modules.scala 160:64:@35199.4]
  assign _T_87834 = _T_87833[13:0]; // @[Modules.scala 160:64:@35200.4]
  assign buffer_10_511 = $signed(_T_87834); // @[Modules.scala 160:64:@35201.4]
  assign _T_87836 = $signed(buffer_10_408) + $signed(buffer_10_409); // @[Modules.scala 160:64:@35203.4]
  assign _T_87837 = _T_87836[13:0]; // @[Modules.scala 160:64:@35204.4]
  assign buffer_10_512 = $signed(_T_87837); // @[Modules.scala 160:64:@35205.4]
  assign _T_87839 = $signed(buffer_10_410) + $signed(buffer_10_411); // @[Modules.scala 160:64:@35207.4]
  assign _T_87840 = _T_87839[13:0]; // @[Modules.scala 160:64:@35208.4]
  assign buffer_10_513 = $signed(_T_87840); // @[Modules.scala 160:64:@35209.4]
  assign _T_87842 = $signed(buffer_10_412) + $signed(buffer_5_418); // @[Modules.scala 160:64:@35211.4]
  assign _T_87843 = _T_87842[13:0]; // @[Modules.scala 160:64:@35212.4]
  assign buffer_10_514 = $signed(_T_87843); // @[Modules.scala 160:64:@35213.4]
  assign _T_87845 = $signed(buffer_10_414) + $signed(buffer_4_400); // @[Modules.scala 160:64:@35215.4]
  assign _T_87846 = _T_87845[13:0]; // @[Modules.scala 160:64:@35216.4]
  assign buffer_10_515 = $signed(_T_87846); // @[Modules.scala 160:64:@35217.4]
  assign _T_87848 = $signed(buffer_0_407) + $signed(buffer_10_417); // @[Modules.scala 160:64:@35219.4]
  assign _T_87849 = _T_87848[13:0]; // @[Modules.scala 160:64:@35220.4]
  assign buffer_10_516 = $signed(_T_87849); // @[Modules.scala 160:64:@35221.4]
  assign _T_87851 = $signed(buffer_10_418) + $signed(buffer_6_430); // @[Modules.scala 160:64:@35223.4]
  assign _T_87852 = _T_87851[13:0]; // @[Modules.scala 160:64:@35224.4]
  assign buffer_10_517 = $signed(_T_87852); // @[Modules.scala 160:64:@35225.4]
  assign _T_87854 = $signed(buffer_7_423) + $signed(buffer_10_421); // @[Modules.scala 160:64:@35227.4]
  assign _T_87855 = _T_87854[13:0]; // @[Modules.scala 160:64:@35228.4]
  assign buffer_10_518 = $signed(_T_87855); // @[Modules.scala 160:64:@35229.4]
  assign _T_87857 = $signed(buffer_10_422) + $signed(buffer_10_423); // @[Modules.scala 160:64:@35231.4]
  assign _T_87858 = _T_87857[13:0]; // @[Modules.scala 160:64:@35232.4]
  assign buffer_10_519 = $signed(_T_87858); // @[Modules.scala 160:64:@35233.4]
  assign _T_87860 = $signed(buffer_10_424) + $signed(buffer_10_425); // @[Modules.scala 160:64:@35235.4]
  assign _T_87861 = _T_87860[13:0]; // @[Modules.scala 160:64:@35236.4]
  assign buffer_10_520 = $signed(_T_87861); // @[Modules.scala 160:64:@35237.4]
  assign _T_87863 = $signed(buffer_10_426) + $signed(buffer_10_427); // @[Modules.scala 160:64:@35239.4]
  assign _T_87864 = _T_87863[13:0]; // @[Modules.scala 160:64:@35240.4]
  assign buffer_10_521 = $signed(_T_87864); // @[Modules.scala 160:64:@35241.4]
  assign _T_87866 = $signed(buffer_10_428) + $signed(buffer_10_429); // @[Modules.scala 160:64:@35243.4]
  assign _T_87867 = _T_87866[13:0]; // @[Modules.scala 160:64:@35244.4]
  assign buffer_10_522 = $signed(_T_87867); // @[Modules.scala 160:64:@35245.4]
  assign _T_87869 = $signed(buffer_10_430) + $signed(buffer_10_431); // @[Modules.scala 160:64:@35247.4]
  assign _T_87870 = _T_87869[13:0]; // @[Modules.scala 160:64:@35248.4]
  assign buffer_10_523 = $signed(_T_87870); // @[Modules.scala 160:64:@35249.4]
  assign _T_87872 = $signed(buffer_3_440) + $signed(buffer_10_433); // @[Modules.scala 160:64:@35251.4]
  assign _T_87873 = _T_87872[13:0]; // @[Modules.scala 160:64:@35252.4]
  assign buffer_10_524 = $signed(_T_87873); // @[Modules.scala 160:64:@35253.4]
  assign _T_87875 = $signed(buffer_10_434) + $signed(buffer_10_435); // @[Modules.scala 160:64:@35255.4]
  assign _T_87876 = _T_87875[13:0]; // @[Modules.scala 160:64:@35256.4]
  assign buffer_10_525 = $signed(_T_87876); // @[Modules.scala 160:64:@35257.4]
  assign _T_87878 = $signed(buffer_10_436) + $signed(buffer_10_437); // @[Modules.scala 160:64:@35259.4]
  assign _T_87879 = _T_87878[13:0]; // @[Modules.scala 160:64:@35260.4]
  assign buffer_10_526 = $signed(_T_87879); // @[Modules.scala 160:64:@35261.4]
  assign _T_87881 = $signed(buffer_2_441) + $signed(buffer_10_439); // @[Modules.scala 160:64:@35263.4]
  assign _T_87882 = _T_87881[13:0]; // @[Modules.scala 160:64:@35264.4]
  assign buffer_10_527 = $signed(_T_87882); // @[Modules.scala 160:64:@35265.4]
  assign _T_87884 = $signed(buffer_10_440) + $signed(buffer_3_449); // @[Modules.scala 160:64:@35267.4]
  assign _T_87885 = _T_87884[13:0]; // @[Modules.scala 160:64:@35268.4]
  assign buffer_10_528 = $signed(_T_87885); // @[Modules.scala 160:64:@35269.4]
  assign _T_87887 = $signed(buffer_3_450) + $signed(buffer_10_443); // @[Modules.scala 160:64:@35271.4]
  assign _T_87888 = _T_87887[13:0]; // @[Modules.scala 160:64:@35272.4]
  assign buffer_10_529 = $signed(_T_87888); // @[Modules.scala 160:64:@35273.4]
  assign _T_87890 = $signed(buffer_10_444) + $signed(buffer_10_445); // @[Modules.scala 160:64:@35275.4]
  assign _T_87891 = _T_87890[13:0]; // @[Modules.scala 160:64:@35276.4]
  assign buffer_10_530 = $signed(_T_87891); // @[Modules.scala 160:64:@35277.4]
  assign _T_87893 = $signed(buffer_10_446) + $signed(buffer_10_447); // @[Modules.scala 160:64:@35279.4]
  assign _T_87894 = _T_87893[13:0]; // @[Modules.scala 160:64:@35280.4]
  assign buffer_10_531 = $signed(_T_87894); // @[Modules.scala 160:64:@35281.4]
  assign _T_87896 = $signed(buffer_10_448) + $signed(buffer_4_436); // @[Modules.scala 160:64:@35283.4]
  assign _T_87897 = _T_87896[13:0]; // @[Modules.scala 160:64:@35284.4]
  assign buffer_10_532 = $signed(_T_87897); // @[Modules.scala 160:64:@35285.4]
  assign _T_87899 = $signed(buffer_4_437) + $signed(buffer_10_451); // @[Modules.scala 160:64:@35287.4]
  assign _T_87900 = _T_87899[13:0]; // @[Modules.scala 160:64:@35288.4]
  assign buffer_10_533 = $signed(_T_87900); // @[Modules.scala 160:64:@35289.4]
  assign _T_87902 = $signed(buffer_10_452) + $signed(buffer_10_453); // @[Modules.scala 160:64:@35291.4]
  assign _T_87903 = _T_87902[13:0]; // @[Modules.scala 160:64:@35292.4]
  assign buffer_10_534 = $signed(_T_87903); // @[Modules.scala 160:64:@35293.4]
  assign _T_87905 = $signed(buffer_10_454) + $signed(buffer_10_455); // @[Modules.scala 160:64:@35295.4]
  assign _T_87906 = _T_87905[13:0]; // @[Modules.scala 160:64:@35296.4]
  assign buffer_10_535 = $signed(_T_87906); // @[Modules.scala 160:64:@35297.4]
  assign _T_87908 = $signed(buffer_10_456) + $signed(buffer_10_457); // @[Modules.scala 160:64:@35299.4]
  assign _T_87909 = _T_87908[13:0]; // @[Modules.scala 160:64:@35300.4]
  assign buffer_10_536 = $signed(_T_87909); // @[Modules.scala 160:64:@35301.4]
  assign _T_87911 = $signed(buffer_10_458) + $signed(buffer_10_459); // @[Modules.scala 160:64:@35303.4]
  assign _T_87912 = _T_87911[13:0]; // @[Modules.scala 160:64:@35304.4]
  assign buffer_10_537 = $signed(_T_87912); // @[Modules.scala 160:64:@35305.4]
  assign _T_87917 = $signed(buffer_10_462) + $signed(buffer_10_463); // @[Modules.scala 166:64:@35311.4]
  assign _T_87918 = _T_87917[13:0]; // @[Modules.scala 166:64:@35312.4]
  assign buffer_10_539 = $signed(_T_87918); // @[Modules.scala 166:64:@35313.4]
  assign _T_87920 = $signed(buffer_10_464) + $signed(buffer_0_456); // @[Modules.scala 166:64:@35315.4]
  assign _T_87921 = _T_87920[13:0]; // @[Modules.scala 166:64:@35316.4]
  assign buffer_10_540 = $signed(_T_87921); // @[Modules.scala 166:64:@35317.4]
  assign _T_87923 = $signed(buffer_0_457) + $signed(buffer_10_467); // @[Modules.scala 166:64:@35319.4]
  assign _T_87924 = _T_87923[13:0]; // @[Modules.scala 166:64:@35320.4]
  assign buffer_10_541 = $signed(_T_87924); // @[Modules.scala 166:64:@35321.4]
  assign _T_87926 = $signed(buffer_10_468) + $signed(buffer_10_469); // @[Modules.scala 166:64:@35323.4]
  assign _T_87927 = _T_87926[13:0]; // @[Modules.scala 166:64:@35324.4]
  assign buffer_10_542 = $signed(_T_87927); // @[Modules.scala 166:64:@35325.4]
  assign _T_87929 = $signed(buffer_10_470) + $signed(buffer_10_471); // @[Modules.scala 166:64:@35327.4]
  assign _T_87930 = _T_87929[13:0]; // @[Modules.scala 166:64:@35328.4]
  assign buffer_10_543 = $signed(_T_87930); // @[Modules.scala 166:64:@35329.4]
  assign _T_87932 = $signed(buffer_10_472) + $signed(buffer_10_473); // @[Modules.scala 166:64:@35331.4]
  assign _T_87933 = _T_87932[13:0]; // @[Modules.scala 166:64:@35332.4]
  assign buffer_10_544 = $signed(_T_87933); // @[Modules.scala 166:64:@35333.4]
  assign _T_87935 = $signed(buffer_10_474) + $signed(buffer_4_463); // @[Modules.scala 166:64:@35335.4]
  assign _T_87936 = _T_87935[13:0]; // @[Modules.scala 166:64:@35336.4]
  assign buffer_10_545 = $signed(_T_87936); // @[Modules.scala 166:64:@35337.4]
  assign _T_87938 = $signed(buffer_10_476) + $signed(buffer_10_477); // @[Modules.scala 166:64:@35339.4]
  assign _T_87939 = _T_87938[13:0]; // @[Modules.scala 166:64:@35340.4]
  assign buffer_10_546 = $signed(_T_87939); // @[Modules.scala 166:64:@35341.4]
  assign _T_87941 = $signed(buffer_10_478) + $signed(buffer_10_479); // @[Modules.scala 166:64:@35343.4]
  assign _T_87942 = _T_87941[13:0]; // @[Modules.scala 166:64:@35344.4]
  assign buffer_10_547 = $signed(_T_87942); // @[Modules.scala 166:64:@35345.4]
  assign _T_87944 = $signed(buffer_10_480) + $signed(buffer_10_481); // @[Modules.scala 166:64:@35347.4]
  assign _T_87945 = _T_87944[13:0]; // @[Modules.scala 166:64:@35348.4]
  assign buffer_10_548 = $signed(_T_87945); // @[Modules.scala 166:64:@35349.4]
  assign _T_87947 = $signed(buffer_10_482) + $signed(buffer_10_483); // @[Modules.scala 166:64:@35351.4]
  assign _T_87948 = _T_87947[13:0]; // @[Modules.scala 166:64:@35352.4]
  assign buffer_10_549 = $signed(_T_87948); // @[Modules.scala 166:64:@35353.4]
  assign _T_87950 = $signed(buffer_10_484) + $signed(buffer_10_485); // @[Modules.scala 166:64:@35355.4]
  assign _T_87951 = _T_87950[13:0]; // @[Modules.scala 166:64:@35356.4]
  assign buffer_10_550 = $signed(_T_87951); // @[Modules.scala 166:64:@35357.4]
  assign _T_87953 = $signed(buffer_10_486) + $signed(buffer_10_487); // @[Modules.scala 166:64:@35359.4]
  assign _T_87954 = _T_87953[13:0]; // @[Modules.scala 166:64:@35360.4]
  assign buffer_10_551 = $signed(_T_87954); // @[Modules.scala 166:64:@35361.4]
  assign _T_87956 = $signed(buffer_10_488) + $signed(buffer_10_489); // @[Modules.scala 166:64:@35363.4]
  assign _T_87957 = _T_87956[13:0]; // @[Modules.scala 166:64:@35364.4]
  assign buffer_10_552 = $signed(_T_87957); // @[Modules.scala 166:64:@35365.4]
  assign _T_87959 = $signed(buffer_10_490) + $signed(buffer_10_491); // @[Modules.scala 166:64:@35367.4]
  assign _T_87960 = _T_87959[13:0]; // @[Modules.scala 166:64:@35368.4]
  assign buffer_10_553 = $signed(_T_87960); // @[Modules.scala 166:64:@35369.4]
  assign _T_87962 = $signed(buffer_10_492) + $signed(buffer_10_493); // @[Modules.scala 166:64:@35371.4]
  assign _T_87963 = _T_87962[13:0]; // @[Modules.scala 166:64:@35372.4]
  assign buffer_10_554 = $signed(_T_87963); // @[Modules.scala 166:64:@35373.4]
  assign _T_87965 = $signed(buffer_10_494) + $signed(buffer_10_495); // @[Modules.scala 166:64:@35375.4]
  assign _T_87966 = _T_87965[13:0]; // @[Modules.scala 166:64:@35376.4]
  assign buffer_10_555 = $signed(_T_87966); // @[Modules.scala 166:64:@35377.4]
  assign _T_87968 = $signed(buffer_10_496) + $signed(buffer_10_497); // @[Modules.scala 166:64:@35379.4]
  assign _T_87969 = _T_87968[13:0]; // @[Modules.scala 166:64:@35380.4]
  assign buffer_10_556 = $signed(_T_87969); // @[Modules.scala 166:64:@35381.4]
  assign _T_87971 = $signed(buffer_10_498) + $signed(buffer_10_499); // @[Modules.scala 166:64:@35383.4]
  assign _T_87972 = _T_87971[13:0]; // @[Modules.scala 166:64:@35384.4]
  assign buffer_10_557 = $signed(_T_87972); // @[Modules.scala 166:64:@35385.4]
  assign _T_87974 = $signed(buffer_10_500) + $signed(buffer_10_501); // @[Modules.scala 166:64:@35387.4]
  assign _T_87975 = _T_87974[13:0]; // @[Modules.scala 166:64:@35388.4]
  assign buffer_10_558 = $signed(_T_87975); // @[Modules.scala 166:64:@35389.4]
  assign _T_87977 = $signed(buffer_10_502) + $signed(buffer_10_503); // @[Modules.scala 166:64:@35391.4]
  assign _T_87978 = _T_87977[13:0]; // @[Modules.scala 166:64:@35392.4]
  assign buffer_10_559 = $signed(_T_87978); // @[Modules.scala 166:64:@35393.4]
  assign _T_87980 = $signed(buffer_10_504) + $signed(buffer_10_505); // @[Modules.scala 166:64:@35395.4]
  assign _T_87981 = _T_87980[13:0]; // @[Modules.scala 166:64:@35396.4]
  assign buffer_10_560 = $signed(_T_87981); // @[Modules.scala 166:64:@35397.4]
  assign _T_87983 = $signed(buffer_10_506) + $signed(buffer_10_507); // @[Modules.scala 166:64:@35399.4]
  assign _T_87984 = _T_87983[13:0]; // @[Modules.scala 166:64:@35400.4]
  assign buffer_10_561 = $signed(_T_87984); // @[Modules.scala 166:64:@35401.4]
  assign _T_87986 = $signed(buffer_10_508) + $signed(buffer_10_509); // @[Modules.scala 166:64:@35403.4]
  assign _T_87987 = _T_87986[13:0]; // @[Modules.scala 166:64:@35404.4]
  assign buffer_10_562 = $signed(_T_87987); // @[Modules.scala 166:64:@35405.4]
  assign _T_87989 = $signed(buffer_10_510) + $signed(buffer_10_511); // @[Modules.scala 166:64:@35407.4]
  assign _T_87990 = _T_87989[13:0]; // @[Modules.scala 166:64:@35408.4]
  assign buffer_10_563 = $signed(_T_87990); // @[Modules.scala 166:64:@35409.4]
  assign _T_87992 = $signed(buffer_10_512) + $signed(buffer_10_513); // @[Modules.scala 166:64:@35411.4]
  assign _T_87993 = _T_87992[13:0]; // @[Modules.scala 166:64:@35412.4]
  assign buffer_10_564 = $signed(_T_87993); // @[Modules.scala 166:64:@35413.4]
  assign _T_87995 = $signed(buffer_10_514) + $signed(buffer_10_515); // @[Modules.scala 166:64:@35415.4]
  assign _T_87996 = _T_87995[13:0]; // @[Modules.scala 166:64:@35416.4]
  assign buffer_10_565 = $signed(_T_87996); // @[Modules.scala 166:64:@35417.4]
  assign _T_87998 = $signed(buffer_10_516) + $signed(buffer_10_517); // @[Modules.scala 166:64:@35419.4]
  assign _T_87999 = _T_87998[13:0]; // @[Modules.scala 166:64:@35420.4]
  assign buffer_10_566 = $signed(_T_87999); // @[Modules.scala 166:64:@35421.4]
  assign _T_88001 = $signed(buffer_10_518) + $signed(buffer_10_519); // @[Modules.scala 166:64:@35423.4]
  assign _T_88002 = _T_88001[13:0]; // @[Modules.scala 166:64:@35424.4]
  assign buffer_10_567 = $signed(_T_88002); // @[Modules.scala 166:64:@35425.4]
  assign _T_88004 = $signed(buffer_10_520) + $signed(buffer_10_521); // @[Modules.scala 166:64:@35427.4]
  assign _T_88005 = _T_88004[13:0]; // @[Modules.scala 166:64:@35428.4]
  assign buffer_10_568 = $signed(_T_88005); // @[Modules.scala 166:64:@35429.4]
  assign _T_88007 = $signed(buffer_10_522) + $signed(buffer_10_523); // @[Modules.scala 166:64:@35431.4]
  assign _T_88008 = _T_88007[13:0]; // @[Modules.scala 166:64:@35432.4]
  assign buffer_10_569 = $signed(_T_88008); // @[Modules.scala 166:64:@35433.4]
  assign _T_88010 = $signed(buffer_10_524) + $signed(buffer_10_525); // @[Modules.scala 166:64:@35435.4]
  assign _T_88011 = _T_88010[13:0]; // @[Modules.scala 166:64:@35436.4]
  assign buffer_10_570 = $signed(_T_88011); // @[Modules.scala 166:64:@35437.4]
  assign _T_88013 = $signed(buffer_10_526) + $signed(buffer_10_527); // @[Modules.scala 166:64:@35439.4]
  assign _T_88014 = _T_88013[13:0]; // @[Modules.scala 166:64:@35440.4]
  assign buffer_10_571 = $signed(_T_88014); // @[Modules.scala 166:64:@35441.4]
  assign _T_88016 = $signed(buffer_10_528) + $signed(buffer_10_529); // @[Modules.scala 166:64:@35443.4]
  assign _T_88017 = _T_88016[13:0]; // @[Modules.scala 166:64:@35444.4]
  assign buffer_10_572 = $signed(_T_88017); // @[Modules.scala 166:64:@35445.4]
  assign _T_88019 = $signed(buffer_10_530) + $signed(buffer_10_531); // @[Modules.scala 166:64:@35447.4]
  assign _T_88020 = _T_88019[13:0]; // @[Modules.scala 166:64:@35448.4]
  assign buffer_10_573 = $signed(_T_88020); // @[Modules.scala 166:64:@35449.4]
  assign _T_88022 = $signed(buffer_10_532) + $signed(buffer_10_533); // @[Modules.scala 166:64:@35451.4]
  assign _T_88023 = _T_88022[13:0]; // @[Modules.scala 166:64:@35452.4]
  assign buffer_10_574 = $signed(_T_88023); // @[Modules.scala 166:64:@35453.4]
  assign _T_88025 = $signed(buffer_10_534) + $signed(buffer_10_535); // @[Modules.scala 166:64:@35455.4]
  assign _T_88026 = _T_88025[13:0]; // @[Modules.scala 166:64:@35456.4]
  assign buffer_10_575 = $signed(_T_88026); // @[Modules.scala 166:64:@35457.4]
  assign _T_88028 = $signed(buffer_10_536) + $signed(buffer_10_537); // @[Modules.scala 166:64:@35459.4]
  assign _T_88029 = _T_88028[13:0]; // @[Modules.scala 166:64:@35460.4]
  assign buffer_10_576 = $signed(_T_88029); // @[Modules.scala 166:64:@35461.4]
  assign _T_88031 = $signed(buffer_10_539) + $signed(buffer_10_540); // @[Modules.scala 160:64:@35463.4]
  assign _T_88032 = _T_88031[13:0]; // @[Modules.scala 160:64:@35464.4]
  assign buffer_10_577 = $signed(_T_88032); // @[Modules.scala 160:64:@35465.4]
  assign _T_88034 = $signed(buffer_10_541) + $signed(buffer_10_542); // @[Modules.scala 160:64:@35467.4]
  assign _T_88035 = _T_88034[13:0]; // @[Modules.scala 160:64:@35468.4]
  assign buffer_10_578 = $signed(_T_88035); // @[Modules.scala 160:64:@35469.4]
  assign _T_88037 = $signed(buffer_10_543) + $signed(buffer_10_544); // @[Modules.scala 160:64:@35471.4]
  assign _T_88038 = _T_88037[13:0]; // @[Modules.scala 160:64:@35472.4]
  assign buffer_10_579 = $signed(_T_88038); // @[Modules.scala 160:64:@35473.4]
  assign _T_88040 = $signed(buffer_10_545) + $signed(buffer_10_546); // @[Modules.scala 160:64:@35475.4]
  assign _T_88041 = _T_88040[13:0]; // @[Modules.scala 160:64:@35476.4]
  assign buffer_10_580 = $signed(_T_88041); // @[Modules.scala 160:64:@35477.4]
  assign _T_88043 = $signed(buffer_10_547) + $signed(buffer_10_548); // @[Modules.scala 160:64:@35479.4]
  assign _T_88044 = _T_88043[13:0]; // @[Modules.scala 160:64:@35480.4]
  assign buffer_10_581 = $signed(_T_88044); // @[Modules.scala 160:64:@35481.4]
  assign _T_88046 = $signed(buffer_10_549) + $signed(buffer_10_550); // @[Modules.scala 160:64:@35483.4]
  assign _T_88047 = _T_88046[13:0]; // @[Modules.scala 160:64:@35484.4]
  assign buffer_10_582 = $signed(_T_88047); // @[Modules.scala 160:64:@35485.4]
  assign _T_88049 = $signed(buffer_10_551) + $signed(buffer_10_552); // @[Modules.scala 160:64:@35487.4]
  assign _T_88050 = _T_88049[13:0]; // @[Modules.scala 160:64:@35488.4]
  assign buffer_10_583 = $signed(_T_88050); // @[Modules.scala 160:64:@35489.4]
  assign _T_88052 = $signed(buffer_10_553) + $signed(buffer_10_554); // @[Modules.scala 160:64:@35491.4]
  assign _T_88053 = _T_88052[13:0]; // @[Modules.scala 160:64:@35492.4]
  assign buffer_10_584 = $signed(_T_88053); // @[Modules.scala 160:64:@35493.4]
  assign _T_88055 = $signed(buffer_10_555) + $signed(buffer_10_556); // @[Modules.scala 160:64:@35495.4]
  assign _T_88056 = _T_88055[13:0]; // @[Modules.scala 160:64:@35496.4]
  assign buffer_10_585 = $signed(_T_88056); // @[Modules.scala 160:64:@35497.4]
  assign _T_88058 = $signed(buffer_10_557) + $signed(buffer_10_558); // @[Modules.scala 160:64:@35499.4]
  assign _T_88059 = _T_88058[13:0]; // @[Modules.scala 160:64:@35500.4]
  assign buffer_10_586 = $signed(_T_88059); // @[Modules.scala 160:64:@35501.4]
  assign _T_88061 = $signed(buffer_10_559) + $signed(buffer_10_560); // @[Modules.scala 160:64:@35503.4]
  assign _T_88062 = _T_88061[13:0]; // @[Modules.scala 160:64:@35504.4]
  assign buffer_10_587 = $signed(_T_88062); // @[Modules.scala 160:64:@35505.4]
  assign _T_88064 = $signed(buffer_10_561) + $signed(buffer_10_562); // @[Modules.scala 160:64:@35507.4]
  assign _T_88065 = _T_88064[13:0]; // @[Modules.scala 160:64:@35508.4]
  assign buffer_10_588 = $signed(_T_88065); // @[Modules.scala 160:64:@35509.4]
  assign _T_88067 = $signed(buffer_10_563) + $signed(buffer_10_564); // @[Modules.scala 160:64:@35511.4]
  assign _T_88068 = _T_88067[13:0]; // @[Modules.scala 160:64:@35512.4]
  assign buffer_10_589 = $signed(_T_88068); // @[Modules.scala 160:64:@35513.4]
  assign _T_88070 = $signed(buffer_10_565) + $signed(buffer_10_566); // @[Modules.scala 160:64:@35515.4]
  assign _T_88071 = _T_88070[13:0]; // @[Modules.scala 160:64:@35516.4]
  assign buffer_10_590 = $signed(_T_88071); // @[Modules.scala 160:64:@35517.4]
  assign _T_88073 = $signed(buffer_10_567) + $signed(buffer_10_568); // @[Modules.scala 160:64:@35519.4]
  assign _T_88074 = _T_88073[13:0]; // @[Modules.scala 160:64:@35520.4]
  assign buffer_10_591 = $signed(_T_88074); // @[Modules.scala 160:64:@35521.4]
  assign _T_88076 = $signed(buffer_10_569) + $signed(buffer_10_570); // @[Modules.scala 160:64:@35523.4]
  assign _T_88077 = _T_88076[13:0]; // @[Modules.scala 160:64:@35524.4]
  assign buffer_10_592 = $signed(_T_88077); // @[Modules.scala 160:64:@35525.4]
  assign _T_88079 = $signed(buffer_10_571) + $signed(buffer_10_572); // @[Modules.scala 160:64:@35527.4]
  assign _T_88080 = _T_88079[13:0]; // @[Modules.scala 160:64:@35528.4]
  assign buffer_10_593 = $signed(_T_88080); // @[Modules.scala 160:64:@35529.4]
  assign _T_88082 = $signed(buffer_10_573) + $signed(buffer_10_574); // @[Modules.scala 160:64:@35531.4]
  assign _T_88083 = _T_88082[13:0]; // @[Modules.scala 160:64:@35532.4]
  assign buffer_10_594 = $signed(_T_88083); // @[Modules.scala 160:64:@35533.4]
  assign _T_88085 = $signed(buffer_10_575) + $signed(buffer_10_576); // @[Modules.scala 160:64:@35535.4]
  assign _T_88086 = _T_88085[13:0]; // @[Modules.scala 160:64:@35536.4]
  assign buffer_10_595 = $signed(_T_88086); // @[Modules.scala 160:64:@35537.4]
  assign _T_88088 = $signed(buffer_10_577) + $signed(buffer_10_578); // @[Modules.scala 166:64:@35539.4]
  assign _T_88089 = _T_88088[13:0]; // @[Modules.scala 166:64:@35540.4]
  assign buffer_10_596 = $signed(_T_88089); // @[Modules.scala 166:64:@35541.4]
  assign _T_88091 = $signed(buffer_10_579) + $signed(buffer_10_580); // @[Modules.scala 166:64:@35543.4]
  assign _T_88092 = _T_88091[13:0]; // @[Modules.scala 166:64:@35544.4]
  assign buffer_10_597 = $signed(_T_88092); // @[Modules.scala 166:64:@35545.4]
  assign _T_88094 = $signed(buffer_10_581) + $signed(buffer_10_582); // @[Modules.scala 166:64:@35547.4]
  assign _T_88095 = _T_88094[13:0]; // @[Modules.scala 166:64:@35548.4]
  assign buffer_10_598 = $signed(_T_88095); // @[Modules.scala 166:64:@35549.4]
  assign _T_88097 = $signed(buffer_10_583) + $signed(buffer_10_584); // @[Modules.scala 166:64:@35551.4]
  assign _T_88098 = _T_88097[13:0]; // @[Modules.scala 166:64:@35552.4]
  assign buffer_10_599 = $signed(_T_88098); // @[Modules.scala 166:64:@35553.4]
  assign _T_88100 = $signed(buffer_10_585) + $signed(buffer_10_586); // @[Modules.scala 166:64:@35555.4]
  assign _T_88101 = _T_88100[13:0]; // @[Modules.scala 166:64:@35556.4]
  assign buffer_10_600 = $signed(_T_88101); // @[Modules.scala 166:64:@35557.4]
  assign _T_88103 = $signed(buffer_10_587) + $signed(buffer_10_588); // @[Modules.scala 166:64:@35559.4]
  assign _T_88104 = _T_88103[13:0]; // @[Modules.scala 166:64:@35560.4]
  assign buffer_10_601 = $signed(_T_88104); // @[Modules.scala 166:64:@35561.4]
  assign _T_88106 = $signed(buffer_10_589) + $signed(buffer_10_590); // @[Modules.scala 166:64:@35563.4]
  assign _T_88107 = _T_88106[13:0]; // @[Modules.scala 166:64:@35564.4]
  assign buffer_10_602 = $signed(_T_88107); // @[Modules.scala 166:64:@35565.4]
  assign _T_88109 = $signed(buffer_10_591) + $signed(buffer_10_592); // @[Modules.scala 166:64:@35567.4]
  assign _T_88110 = _T_88109[13:0]; // @[Modules.scala 166:64:@35568.4]
  assign buffer_10_603 = $signed(_T_88110); // @[Modules.scala 166:64:@35569.4]
  assign _T_88112 = $signed(buffer_10_593) + $signed(buffer_10_594); // @[Modules.scala 166:64:@35571.4]
  assign _T_88113 = _T_88112[13:0]; // @[Modules.scala 166:64:@35572.4]
  assign buffer_10_604 = $signed(_T_88113); // @[Modules.scala 166:64:@35573.4]
  assign _T_88115 = $signed(buffer_10_595) + $signed(buffer_4_524); // @[Modules.scala 172:66:@35575.4]
  assign _T_88116 = _T_88115[13:0]; // @[Modules.scala 172:66:@35576.4]
  assign buffer_10_605 = $signed(_T_88116); // @[Modules.scala 172:66:@35577.4]
  assign _T_88118 = $signed(buffer_10_596) + $signed(buffer_10_597); // @[Modules.scala 160:64:@35579.4]
  assign _T_88119 = _T_88118[13:0]; // @[Modules.scala 160:64:@35580.4]
  assign buffer_10_606 = $signed(_T_88119); // @[Modules.scala 160:64:@35581.4]
  assign _T_88121 = $signed(buffer_10_598) + $signed(buffer_10_599); // @[Modules.scala 160:64:@35583.4]
  assign _T_88122 = _T_88121[13:0]; // @[Modules.scala 160:64:@35584.4]
  assign buffer_10_607 = $signed(_T_88122); // @[Modules.scala 160:64:@35585.4]
  assign _T_88124 = $signed(buffer_10_600) + $signed(buffer_10_601); // @[Modules.scala 160:64:@35587.4]
  assign _T_88125 = _T_88124[13:0]; // @[Modules.scala 160:64:@35588.4]
  assign buffer_10_608 = $signed(_T_88125); // @[Modules.scala 160:64:@35589.4]
  assign _T_88127 = $signed(buffer_10_602) + $signed(buffer_10_603); // @[Modules.scala 160:64:@35591.4]
  assign _T_88128 = _T_88127[13:0]; // @[Modules.scala 160:64:@35592.4]
  assign buffer_10_609 = $signed(_T_88128); // @[Modules.scala 160:64:@35593.4]
  assign _T_88130 = $signed(buffer_10_604) + $signed(buffer_10_605); // @[Modules.scala 160:64:@35595.4]
  assign _T_88131 = _T_88130[13:0]; // @[Modules.scala 160:64:@35596.4]
  assign buffer_10_610 = $signed(_T_88131); // @[Modules.scala 160:64:@35597.4]
  assign _T_88133 = $signed(buffer_10_606) + $signed(buffer_10_607); // @[Modules.scala 166:64:@35599.4]
  assign _T_88134 = _T_88133[13:0]; // @[Modules.scala 166:64:@35600.4]
  assign buffer_10_611 = $signed(_T_88134); // @[Modules.scala 166:64:@35601.4]
  assign _T_88136 = $signed(buffer_10_608) + $signed(buffer_10_609); // @[Modules.scala 166:64:@35603.4]
  assign _T_88137 = _T_88136[13:0]; // @[Modules.scala 166:64:@35604.4]
  assign buffer_10_612 = $signed(_T_88137); // @[Modules.scala 166:64:@35605.4]
  assign _T_88139 = $signed(buffer_10_611) + $signed(buffer_10_612); // @[Modules.scala 160:64:@35607.4]
  assign _T_88140 = _T_88139[13:0]; // @[Modules.scala 160:64:@35608.4]
  assign buffer_10_613 = $signed(_T_88140); // @[Modules.scala 160:64:@35609.4]
  assign _T_88142 = $signed(buffer_10_613) + $signed(buffer_10_610); // @[Modules.scala 172:66:@35611.4]
  assign _T_88143 = _T_88142[13:0]; // @[Modules.scala 172:66:@35612.4]
  assign buffer_10_614 = $signed(_T_88143); // @[Modules.scala 172:66:@35613.4]
  assign _T_88146 = $signed(4'sh1) * $signed(io_in_3); // @[Modules.scala 150:74:@35784.4]
  assign _T_88149 = $signed(_T_88146) + $signed(_T_54199); // @[Modules.scala 150:103:@35786.4]
  assign _T_88150 = _T_88149[5:0]; // @[Modules.scala 150:103:@35787.4]
  assign _T_88151 = $signed(_T_88150); // @[Modules.scala 150:103:@35788.4]
  assign _T_88156 = $signed(_T_54201) + $signed(_T_54206); // @[Modules.scala 150:103:@35792.4]
  assign _T_88157 = _T_88156[5:0]; // @[Modules.scala 150:103:@35793.4]
  assign _T_88158 = $signed(_T_88157); // @[Modules.scala 150:103:@35794.4]
  assign _T_88163 = $signed(_T_54208) + $signed(_T_54215); // @[Modules.scala 150:103:@35798.4]
  assign _T_88164 = _T_88163[5:0]; // @[Modules.scala 150:103:@35799.4]
  assign _T_88165 = $signed(_T_88164); // @[Modules.scala 150:103:@35800.4]
  assign _T_88170 = $signed(_T_54220) + $signed(_T_57232); // @[Modules.scala 150:103:@35804.4]
  assign _T_88171 = _T_88170[5:0]; // @[Modules.scala 150:103:@35805.4]
  assign _T_88172 = $signed(_T_88171); // @[Modules.scala 150:103:@35806.4]
  assign _T_88205 = $signed(_T_54250) + $signed(_GEN_359); // @[Modules.scala 150:103:@35834.4]
  assign _T_88206 = _T_88205[5:0]; // @[Modules.scala 150:103:@35835.4]
  assign _T_88207 = $signed(_T_88206); // @[Modules.scala 150:103:@35836.4]
  assign _T_88226 = $signed(_T_54278) + $signed(_T_63429); // @[Modules.scala 150:103:@35852.4]
  assign _T_88227 = _T_88226[5:0]; // @[Modules.scala 150:103:@35853.4]
  assign _T_88228 = $signed(_T_88227); // @[Modules.scala 150:103:@35854.4]
  assign _T_88302 = $signed(4'sh1) * $signed(io_in_82); // @[Modules.scala 151:80:@35917.4]
  assign _T_88303 = $signed(_GEN_571) + $signed(_T_88302); // @[Modules.scala 150:103:@35918.4]
  assign _T_88304 = _T_88303[5:0]; // @[Modules.scala 150:103:@35919.4]
  assign _T_88305 = $signed(_T_88304); // @[Modules.scala 150:103:@35920.4]
  assign _T_88387 = $signed(_T_54432) + $signed(_T_57442); // @[Modules.scala 150:103:@35990.4]
  assign _T_88388 = _T_88387[5:0]; // @[Modules.scala 150:103:@35991.4]
  assign _T_88389 = $signed(_T_88388); // @[Modules.scala 150:103:@35992.4]
  assign _GEN_766 = {{1{_T_69765[4]}},_T_69765}; // @[Modules.scala 150:103:@36038.4]
  assign _T_88443 = $signed(_T_57498) + $signed(_GEN_766); // @[Modules.scala 150:103:@36038.4]
  assign _T_88444 = _T_88443[5:0]; // @[Modules.scala 150:103:@36039.4]
  assign _T_88445 = $signed(_T_88444); // @[Modules.scala 150:103:@36040.4]
  assign _T_88457 = $signed(_GEN_366) + $signed(_T_54516); // @[Modules.scala 150:103:@36050.4]
  assign _T_88458 = _T_88457[5:0]; // @[Modules.scala 150:103:@36051.4]
  assign _T_88459 = $signed(_T_88458); // @[Modules.scala 150:103:@36052.4]
  assign _T_88463 = $signed(4'sh1) * $signed(io_in_140); // @[Modules.scala 151:80:@36055.4]
  assign _T_88464 = $signed(_GEN_86) + $signed(_T_88463); // @[Modules.scala 150:103:@36056.4]
  assign _T_88465 = _T_88464[5:0]; // @[Modules.scala 150:103:@36057.4]
  assign _T_88466 = $signed(_T_88465); // @[Modules.scala 150:103:@36058.4]
  assign _T_88485 = $signed(_T_57540) + $signed(_GEN_578); // @[Modules.scala 150:103:@36074.4]
  assign _T_88486 = _T_88485[5:0]; // @[Modules.scala 150:103:@36075.4]
  assign _T_88487 = $signed(_T_88486); // @[Modules.scala 150:103:@36076.4]
  assign _T_88541 = $signed(_GEN_12) + $signed(_T_60633); // @[Modules.scala 150:103:@36122.4]
  assign _T_88542 = _T_88541[5:0]; // @[Modules.scala 150:103:@36123.4]
  assign _T_88543 = $signed(_T_88542); // @[Modules.scala 150:103:@36124.4]
  assign _T_88562 = $signed(_T_54600) + $signed(_GEN_14); // @[Modules.scala 150:103:@36140.4]
  assign _T_88563 = _T_88562[5:0]; // @[Modules.scala 150:103:@36141.4]
  assign _T_88564 = $signed(_T_88563); // @[Modules.scala 150:103:@36142.4]
  assign _T_88580 = $signed(4'sh1) * $signed(io_in_187); // @[Modules.scala 150:74:@36156.4]
  assign _T_88583 = $signed(_T_88580) + $signed(_T_69924); // @[Modules.scala 150:103:@36158.4]
  assign _T_88584 = _T_88583[5:0]; // @[Modules.scala 150:103:@36159.4]
  assign _T_88585 = $signed(_T_88584); // @[Modules.scala 150:103:@36160.4]
  assign _T_88590 = $signed(_T_54635) + $signed(_T_54642); // @[Modules.scala 150:103:@36164.4]
  assign _T_88591 = _T_88590[4:0]; // @[Modules.scala 150:103:@36165.4]
  assign _T_88592 = $signed(_T_88591); // @[Modules.scala 150:103:@36166.4]
  assign _T_88597 = $signed(_T_63823) + $signed(_GEN_15); // @[Modules.scala 150:103:@36170.4]
  assign _T_88598 = _T_88597[5:0]; // @[Modules.scala 150:103:@36171.4]
  assign _T_88599 = $signed(_T_88598); // @[Modules.scala 150:103:@36172.4]
  assign _T_88604 = $signed(_T_69947) + $signed(_T_63835); // @[Modules.scala 150:103:@36176.4]
  assign _T_88605 = _T_88604[4:0]; // @[Modules.scala 150:103:@36177.4]
  assign _T_88606 = $signed(_T_88605); // @[Modules.scala 150:103:@36178.4]
  assign _GEN_776 = {{1{_T_60726[4]}},_T_60726}; // @[Modules.scala 150:103:@36188.4]
  assign _T_88618 = $signed(_T_54675) + $signed(_GEN_776); // @[Modules.scala 150:103:@36188.4]
  assign _T_88619 = _T_88618[5:0]; // @[Modules.scala 150:103:@36189.4]
  assign _T_88620 = $signed(_T_88619); // @[Modules.scala 150:103:@36190.4]
  assign _T_88639 = $signed(_T_57722) + $signed(_T_63884); // @[Modules.scala 150:103:@36206.4]
  assign _T_88640 = _T_88639[5:0]; // @[Modules.scala 150:103:@36207.4]
  assign _T_88641 = $signed(_T_88640); // @[Modules.scala 150:103:@36208.4]
  assign _T_88653 = $signed(_T_70010) + $signed(_T_63898); // @[Modules.scala 150:103:@36218.4]
  assign _T_88654 = _T_88653[5:0]; // @[Modules.scala 150:103:@36219.4]
  assign _T_88655 = $signed(_T_88654); // @[Modules.scala 150:103:@36220.4]
  assign _T_88681 = $signed(_T_60810) + $signed(_T_60815); // @[Modules.scala 150:103:@36242.4]
  assign _T_88682 = _T_88681[4:0]; // @[Modules.scala 150:103:@36243.4]
  assign _T_88683 = $signed(_T_88682); // @[Modules.scala 150:103:@36244.4]
  assign _GEN_777 = {{1{_T_60829[4]}},_T_60829}; // @[Modules.scala 150:103:@36254.4]
  assign _T_88695 = $signed(_GEN_777) + $signed(_T_70057); // @[Modules.scala 150:103:@36254.4]
  assign _T_88696 = _T_88695[5:0]; // @[Modules.scala 150:103:@36255.4]
  assign _T_88697 = $signed(_T_88696); // @[Modules.scala 150:103:@36256.4]
  assign _T_88702 = $signed(_T_70059) + $signed(_T_57813); // @[Modules.scala 150:103:@36260.4]
  assign _T_88703 = _T_88702[5:0]; // @[Modules.scala 150:103:@36261.4]
  assign _T_88704 = $signed(_T_88703); // @[Modules.scala 150:103:@36262.4]
  assign _T_88709 = $signed(_T_57815) + $signed(_T_63968); // @[Modules.scala 150:103:@36266.4]
  assign _T_88710 = _T_88709[5:0]; // @[Modules.scala 150:103:@36267.4]
  assign _T_88711 = $signed(_T_88710); // @[Modules.scala 150:103:@36268.4]
  assign _T_88716 = $signed(_GEN_592) + $signed(_T_70099); // @[Modules.scala 150:103:@36272.4]
  assign _T_88717 = _T_88716[5:0]; // @[Modules.scala 150:103:@36273.4]
  assign _T_88718 = $signed(_T_88717); // @[Modules.scala 150:103:@36274.4]
  assign _GEN_779 = {{1{_T_54796[4]}},_T_54796}; // @[Modules.scala 150:103:@36284.4]
  assign _T_88730 = $signed(_GEN_779) + $signed(_T_63989); // @[Modules.scala 150:103:@36284.4]
  assign _T_88731 = _T_88730[5:0]; // @[Modules.scala 150:103:@36285.4]
  assign _T_88732 = $signed(_T_88731); // @[Modules.scala 150:103:@36286.4]
  assign _T_88765 = $signed(_T_57869) + $signed(_T_60920); // @[Modules.scala 150:103:@36314.4]
  assign _T_88766 = _T_88765[4:0]; // @[Modules.scala 150:103:@36315.4]
  assign _T_88767 = $signed(_T_88766); // @[Modules.scala 150:103:@36316.4]
  assign _GEN_781 = {{1{_T_60936[4]}},_T_60936}; // @[Modules.scala 150:103:@36332.4]
  assign _T_88786 = $signed(_GEN_781) + $signed(_T_57890); // @[Modules.scala 150:103:@36332.4]
  assign _T_88787 = _T_88786[5:0]; // @[Modules.scala 150:103:@36333.4]
  assign _T_88788 = $signed(_T_88787); // @[Modules.scala 150:103:@36334.4]
  assign _GEN_782 = {{1{_T_54866[4]}},_T_54866}; // @[Modules.scala 150:103:@36344.4]
  assign _T_88800 = $signed(_T_57899) + $signed(_GEN_782); // @[Modules.scala 150:103:@36344.4]
  assign _T_88801 = _T_88800[5:0]; // @[Modules.scala 150:103:@36345.4]
  assign _T_88802 = $signed(_T_88801); // @[Modules.scala 150:103:@36346.4]
  assign _T_88814 = $signed(_T_54885) + $signed(_T_54892); // @[Modules.scala 150:103:@36356.4]
  assign _T_88815 = _T_88814[4:0]; // @[Modules.scala 150:103:@36357.4]
  assign _T_88816 = $signed(_T_88815); // @[Modules.scala 150:103:@36358.4]
  assign _T_88835 = $signed(_T_54915) + $signed(_T_54927); // @[Modules.scala 150:103:@36374.4]
  assign _T_88836 = _T_88835[4:0]; // @[Modules.scala 150:103:@36375.4]
  assign _T_88837 = $signed(_T_88836); // @[Modules.scala 150:103:@36376.4]
  assign _GEN_783 = {{1{_T_61013[4]}},_T_61013}; // @[Modules.scala 150:103:@36392.4]
  assign _T_88856 = $signed(_GEN_783) + $signed(_T_54948); // @[Modules.scala 150:103:@36392.4]
  assign _T_88857 = _T_88856[5:0]; // @[Modules.scala 150:103:@36393.4]
  assign _T_88858 = $signed(_T_88857); // @[Modules.scala 150:103:@36394.4]
  assign _T_88940 = $signed(_T_55027) + $signed(_T_55032); // @[Modules.scala 150:103:@36464.4]
  assign _T_88941 = _T_88940[4:0]; // @[Modules.scala 150:103:@36465.4]
  assign _T_88942 = $signed(_T_88941); // @[Modules.scala 150:103:@36466.4]
  assign _T_88975 = $signed(_T_67324) + $signed(_T_70351); // @[Modules.scala 150:103:@36494.4]
  assign _T_88976 = _T_88975[5:0]; // @[Modules.scala 150:103:@36495.4]
  assign _T_88977 = $signed(_T_88976); // @[Modules.scala 150:103:@36496.4]
  assign _GEN_787 = {{1{_T_55069[4]}},_T_55069}; // @[Modules.scala 150:103:@36500.4]
  assign _T_88982 = $signed(_T_70353) + $signed(_GEN_787); // @[Modules.scala 150:103:@36500.4]
  assign _T_88983 = _T_88982[5:0]; // @[Modules.scala 150:103:@36501.4]
  assign _T_88984 = $signed(_T_88983); // @[Modules.scala 150:103:@36502.4]
  assign _T_89045 = $signed(_T_58158) + $signed(_T_58163); // @[Modules.scala 150:103:@36554.4]
  assign _T_89046 = _T_89045[5:0]; // @[Modules.scala 150:103:@36555.4]
  assign _T_89047 = $signed(_T_89046); // @[Modules.scala 150:103:@36556.4]
  assign _T_89052 = $signed(_T_55137) + $signed(_T_58170); // @[Modules.scala 150:103:@36560.4]
  assign _T_89053 = _T_89052[5:0]; // @[Modules.scala 150:103:@36561.4]
  assign _T_89054 = $signed(_T_89053); // @[Modules.scala 150:103:@36562.4]
  assign _T_89066 = $signed(_T_55151) + $signed(_T_58177); // @[Modules.scala 150:103:@36572.4]
  assign _T_89067 = _T_89066[5:0]; // @[Modules.scala 150:103:@36573.4]
  assign _T_89068 = $signed(_T_89067); // @[Modules.scala 150:103:@36574.4]
  assign _T_89073 = $signed(_T_64355) + $signed(_GEN_240); // @[Modules.scala 150:103:@36578.4]
  assign _T_89074 = _T_89073[5:0]; // @[Modules.scala 150:103:@36579.4]
  assign _T_89075 = $signed(_T_89074); // @[Modules.scala 150:103:@36580.4]
  assign _T_89101 = $signed(_T_55188) + $signed(_T_55200); // @[Modules.scala 150:103:@36602.4]
  assign _T_89102 = _T_89101[4:0]; // @[Modules.scala 150:103:@36603.4]
  assign _T_89103 = $signed(_T_89102); // @[Modules.scala 150:103:@36604.4]
  assign _GEN_792 = {{1{_T_55202[4]}},_T_55202}; // @[Modules.scala 150:103:@36608.4]
  assign _T_89108 = $signed(_GEN_792) + $signed(_T_58226); // @[Modules.scala 150:103:@36608.4]
  assign _T_89109 = _T_89108[5:0]; // @[Modules.scala 150:103:@36609.4]
  assign _T_89110 = $signed(_T_89109); // @[Modules.scala 150:103:@36610.4]
  assign _T_89164 = $signed(_T_58277) + $signed(_T_64458); // @[Modules.scala 150:103:@36656.4]
  assign _T_89165 = _T_89164[4:0]; // @[Modules.scala 150:103:@36657.4]
  assign _T_89166 = $signed(_T_89165); // @[Modules.scala 150:103:@36658.4]
  assign _T_89220 = $signed(_T_55312) + $signed(_T_61391); // @[Modules.scala 150:103:@36704.4]
  assign _T_89221 = _T_89220[5:0]; // @[Modules.scala 150:103:@36705.4]
  assign _T_89222 = $signed(_T_89221); // @[Modules.scala 150:103:@36706.4]
  assign _T_89241 = $signed(_GEN_42) + $signed(_T_55326); // @[Modules.scala 150:103:@36722.4]
  assign _T_89242 = _T_89241[5:0]; // @[Modules.scala 150:103:@36723.4]
  assign _T_89243 = $signed(_T_89242); // @[Modules.scala 150:103:@36724.4]
  assign _T_89248 = $signed(_T_67585) + $signed(_GEN_469); // @[Modules.scala 150:103:@36728.4]
  assign _T_89249 = _T_89248[5:0]; // @[Modules.scala 150:103:@36729.4]
  assign _T_89250 = $signed(_T_89249); // @[Modules.scala 150:103:@36730.4]
  assign _T_89262 = $signed(_T_58361) + $signed(_T_61431); // @[Modules.scala 150:103:@36740.4]
  assign _T_89263 = _T_89262[5:0]; // @[Modules.scala 150:103:@36741.4]
  assign _T_89264 = $signed(_T_89263); // @[Modules.scala 150:103:@36742.4]
  assign _T_89276 = $signed(_T_61440) + $signed(_GEN_45); // @[Modules.scala 150:103:@36752.4]
  assign _T_89277 = _T_89276[5:0]; // @[Modules.scala 150:103:@36753.4]
  assign _T_89278 = $signed(_T_89277); // @[Modules.scala 150:103:@36754.4]
  assign _T_89283 = $signed(_T_61447) + $signed(_T_55363); // @[Modules.scala 150:103:@36758.4]
  assign _T_89284 = _T_89283[5:0]; // @[Modules.scala 150:103:@36759.4]
  assign _T_89285 = $signed(_T_89284); // @[Modules.scala 150:103:@36760.4]
  assign _T_89332 = $signed(_T_55410) + $signed(_GEN_179); // @[Modules.scala 150:103:@36800.4]
  assign _T_89333 = _T_89332[5:0]; // @[Modules.scala 150:103:@36801.4]
  assign _T_89334 = $signed(_T_89333); // @[Modules.scala 150:103:@36802.4]
  assign _T_89339 = $signed(_GEN_112) + $signed(_T_55426); // @[Modules.scala 150:103:@36806.4]
  assign _T_89340 = _T_89339[5:0]; // @[Modules.scala 150:103:@36807.4]
  assign _T_89341 = $signed(_T_89340); // @[Modules.scala 150:103:@36808.4]
  assign _T_89345 = $signed(4'sh1) * $signed(io_in_453); // @[Modules.scala 151:80:@36811.4]
  assign _T_89346 = $signed(_T_58438) + $signed(_T_89345); // @[Modules.scala 150:103:@36812.4]
  assign _T_89347 = _T_89346[5:0]; // @[Modules.scala 150:103:@36813.4]
  assign _T_89348 = $signed(_T_89347); // @[Modules.scala 150:103:@36814.4]
  assign _T_89381 = $signed(_T_61545) + $signed(_T_58478); // @[Modules.scala 150:103:@36842.4]
  assign _T_89382 = _T_89381[5:0]; // @[Modules.scala 150:103:@36843.4]
  assign _T_89383 = $signed(_T_89382); // @[Modules.scala 150:103:@36844.4]
  assign _T_89451 = $signed(_GEN_330) + $signed(_T_55510); // @[Modules.scala 150:103:@36902.4]
  assign _T_89452 = _T_89451[5:0]; // @[Modules.scala 150:103:@36903.4]
  assign _T_89453 = $signed(_T_89452); // @[Modules.scala 150:103:@36904.4]
  assign _T_89486 = $signed(_GEN_116) + $signed(_T_55545); // @[Modules.scala 150:103:@36932.4]
  assign _T_89487 = _T_89486[5:0]; // @[Modules.scala 150:103:@36933.4]
  assign _T_89488 = $signed(_T_89487); // @[Modules.scala 150:103:@36934.4]
  assign _T_89514 = $signed(_T_55573) + $signed(_T_55578); // @[Modules.scala 150:103:@36956.4]
  assign _T_89515 = _T_89514[5:0]; // @[Modules.scala 150:103:@36957.4]
  assign _T_89516 = $signed(_T_89515); // @[Modules.scala 150:103:@36958.4]
  assign _T_89521 = $signed(_T_70876) + $signed(_T_55587); // @[Modules.scala 150:103:@36962.4]
  assign _T_89522 = _T_89521[5:0]; // @[Modules.scala 150:103:@36963.4]
  assign _T_89523 = $signed(_T_89522); // @[Modules.scala 150:103:@36964.4]
  assign _T_89542 = $signed(_T_55606) + $signed(_GEN_60); // @[Modules.scala 150:103:@36980.4]
  assign _T_89543 = _T_89542[5:0]; // @[Modules.scala 150:103:@36981.4]
  assign _T_89544 = $signed(_T_89543); // @[Modules.scala 150:103:@36982.4]
  assign _T_89556 = $signed(_T_64831) + $signed(_T_64838); // @[Modules.scala 150:103:@36992.4]
  assign _T_89557 = _T_89556[4:0]; // @[Modules.scala 150:103:@36993.4]
  assign _T_89558 = $signed(_T_89557); // @[Modules.scala 150:103:@36994.4]
  assign _T_89563 = $signed(_GEN_190) + $signed(_T_55629); // @[Modules.scala 150:103:@36998.4]
  assign _T_89564 = _T_89563[5:0]; // @[Modules.scala 150:103:@36999.4]
  assign _T_89565 = $signed(_T_89564); // @[Modules.scala 150:103:@37000.4]
  assign _T_89577 = $signed(_T_55641) + $signed(_GEN_191); // @[Modules.scala 150:103:@37010.4]
  assign _T_89578 = _T_89577[5:0]; // @[Modules.scala 150:103:@37011.4]
  assign _T_89579 = $signed(_T_89578); // @[Modules.scala 150:103:@37012.4]
  assign _T_89584 = $signed(_T_55648) + $signed(_T_58660); // @[Modules.scala 150:103:@37016.4]
  assign _T_89585 = _T_89584[4:0]; // @[Modules.scala 150:103:@37017.4]
  assign _T_89586 = $signed(_T_89585); // @[Modules.scala 150:103:@37018.4]
  assign _T_89598 = $signed(_GEN_612) + $signed(_T_55669); // @[Modules.scala 150:103:@37028.4]
  assign _T_89599 = _T_89598[5:0]; // @[Modules.scala 150:103:@37029.4]
  assign _T_89600 = $signed(_T_89599); // @[Modules.scala 150:103:@37030.4]
  assign _T_89605 = $signed(_T_55671) + $signed(_GEN_192); // @[Modules.scala 150:103:@37034.4]
  assign _T_89606 = _T_89605[5:0]; // @[Modules.scala 150:103:@37035.4]
  assign _T_89607 = $signed(_T_89606); // @[Modules.scala 150:103:@37036.4]
  assign _T_89633 = $signed(_T_58704) + $signed(_T_64920); // @[Modules.scala 150:103:@37058.4]
  assign _T_89634 = _T_89633[4:0]; // @[Modules.scala 150:103:@37059.4]
  assign _T_89635 = $signed(_T_89634); // @[Modules.scala 150:103:@37060.4]
  assign _T_89640 = $signed(_T_67928) + $signed(_T_58723); // @[Modules.scala 150:103:@37064.4]
  assign _T_89641 = _T_89640[4:0]; // @[Modules.scala 150:103:@37065.4]
  assign _T_89642 = $signed(_T_89641); // @[Modules.scala 150:103:@37066.4]
  assign _GEN_814 = {{1{_T_58758[4]}},_T_58758}; // @[Modules.scala 150:103:@37100.4]
  assign _T_89682 = $signed(_GEN_814) + $signed(_T_64969); // @[Modules.scala 150:103:@37100.4]
  assign _T_89683 = _T_89682[5:0]; // @[Modules.scala 150:103:@37101.4]
  assign _T_89684 = $signed(_T_89683); // @[Modules.scala 150:103:@37102.4]
  assign _T_89710 = $signed(_T_67991) + $signed(_T_58774); // @[Modules.scala 150:103:@37124.4]
  assign _T_89711 = _T_89710[4:0]; // @[Modules.scala 150:103:@37125.4]
  assign _T_89712 = $signed(_T_89711); // @[Modules.scala 150:103:@37126.4]
  assign _T_89766 = $signed(_T_55811) + $signed(_T_55816); // @[Modules.scala 150:103:@37172.4]
  assign _T_89767 = _T_89766[5:0]; // @[Modules.scala 150:103:@37173.4]
  assign _T_89768 = $signed(_T_89767); // @[Modules.scala 150:103:@37174.4]
  assign _T_89773 = $signed(_T_61916) + $signed(_T_61921); // @[Modules.scala 150:103:@37178.4]
  assign _T_89774 = _T_89773[4:0]; // @[Modules.scala 150:103:@37179.4]
  assign _T_89775 = $signed(_T_89774); // @[Modules.scala 150:103:@37180.4]
  assign _T_89780 = $signed(_T_71151) + $signed(_T_58844); // @[Modules.scala 150:103:@37184.4]
  assign _T_89781 = _T_89780[4:0]; // @[Modules.scala 150:103:@37185.4]
  assign _T_89782 = $signed(_T_89781); // @[Modules.scala 150:103:@37186.4]
  assign _T_89794 = $signed(_T_68075) + $signed(_T_58851); // @[Modules.scala 150:103:@37196.4]
  assign _T_89795 = _T_89794[4:0]; // @[Modules.scala 150:103:@37197.4]
  assign _T_89796 = $signed(_T_89795); // @[Modules.scala 150:103:@37198.4]
  assign _T_89801 = $signed(_T_74330) + $signed(_GEN_65); // @[Modules.scala 150:103:@37202.4]
  assign _T_89802 = _T_89801[5:0]; // @[Modules.scala 150:103:@37203.4]
  assign _T_89803 = $signed(_T_89802); // @[Modules.scala 150:103:@37204.4]
  assign _T_89808 = $signed(_T_55844) + $signed(_T_55851); // @[Modules.scala 150:103:@37208.4]
  assign _T_89809 = _T_89808[5:0]; // @[Modules.scala 150:103:@37209.4]
  assign _T_89810 = $signed(_T_89809); // @[Modules.scala 150:103:@37210.4]
  assign _T_89815 = $signed(_T_55853) + $signed(_T_55860); // @[Modules.scala 150:103:@37214.4]
  assign _T_89816 = _T_89815[5:0]; // @[Modules.scala 150:103:@37215.4]
  assign _T_89817 = $signed(_T_89816); // @[Modules.scala 150:103:@37216.4]
  assign _T_89836 = $signed(_T_55881) + $signed(_T_71221); // @[Modules.scala 150:103:@37232.4]
  assign _T_89837 = _T_89836[5:0]; // @[Modules.scala 150:103:@37233.4]
  assign _T_89838 = $signed(_T_89837); // @[Modules.scala 150:103:@37234.4]
  assign _T_89843 = $signed(_T_62000) + $signed(_T_55893); // @[Modules.scala 150:103:@37238.4]
  assign _T_89844 = _T_89843[4:0]; // @[Modules.scala 150:103:@37239.4]
  assign _T_89845 = $signed(_T_89844); // @[Modules.scala 150:103:@37240.4]
  assign _GEN_818 = {{1{_T_55902[4]}},_T_55902}; // @[Modules.scala 150:103:@37250.4]
  assign _T_89857 = $signed(_GEN_818) + $signed(_T_62026); // @[Modules.scala 150:103:@37250.4]
  assign _T_89858 = _T_89857[5:0]; // @[Modules.scala 150:103:@37251.4]
  assign _T_89859 = $signed(_T_89858); // @[Modules.scala 150:103:@37252.4]
  assign _GEN_819 = {{1{_T_65165[4]}},_T_65165}; // @[Modules.scala 150:103:@37274.4]
  assign _T_89885 = $signed(_T_55942) + $signed(_GEN_819); // @[Modules.scala 150:103:@37274.4]
  assign _T_89886 = _T_89885[5:0]; // @[Modules.scala 150:103:@37275.4]
  assign _T_89887 = $signed(_T_89886); // @[Modules.scala 150:103:@37276.4]
  assign _T_89927 = $signed(_T_71317) + $signed(_GEN_348); // @[Modules.scala 150:103:@37310.4]
  assign _T_89928 = _T_89927[5:0]; // @[Modules.scala 150:103:@37311.4]
  assign _T_89929 = $signed(_T_89928); // @[Modules.scala 150:103:@37312.4]
  assign _GEN_821 = {{1{_T_62126[4]}},_T_62126}; // @[Modules.scala 150:103:@37322.4]
  assign _T_89941 = $signed(_T_68257) + $signed(_GEN_821); // @[Modules.scala 150:103:@37322.4]
  assign _T_89942 = _T_89941[5:0]; // @[Modules.scala 150:103:@37323.4]
  assign _T_89943 = $signed(_T_89942); // @[Modules.scala 150:103:@37324.4]
  assign _T_89947 = $signed(4'sh1) * $signed(io_in_673); // @[Modules.scala 151:80:@37327.4]
  assign _GEN_822 = {{1{_T_65230[4]}},_T_65230}; // @[Modules.scala 150:103:@37328.4]
  assign _T_89948 = $signed(_GEN_822) + $signed(_T_89947); // @[Modules.scala 150:103:@37328.4]
  assign _T_89949 = _T_89948[5:0]; // @[Modules.scala 150:103:@37329.4]
  assign _T_89950 = $signed(_T_89949); // @[Modules.scala 150:103:@37330.4]
  assign _T_89983 = $signed(_T_56056) + $signed(_T_56068); // @[Modules.scala 150:103:@37358.4]
  assign _T_89984 = _T_89983[4:0]; // @[Modules.scala 150:103:@37359.4]
  assign _T_89985 = $signed(_T_89984); // @[Modules.scala 150:103:@37360.4]
  assign _T_90018 = $signed(_GEN_423) + $signed(_T_56110); // @[Modules.scala 150:103:@37388.4]
  assign _T_90019 = _T_90018[5:0]; // @[Modules.scala 150:103:@37389.4]
  assign _T_90020 = $signed(_T_90019); // @[Modules.scala 150:103:@37390.4]
  assign _T_90025 = $signed(_GEN_138) + $signed(_T_56117); // @[Modules.scala 150:103:@37394.4]
  assign _T_90026 = _T_90025[5:0]; // @[Modules.scala 150:103:@37395.4]
  assign _T_90027 = $signed(_T_90026); // @[Modules.scala 150:103:@37396.4]
  assign _T_90032 = $signed(_T_59124) + $signed(_GEN_70); // @[Modules.scala 150:103:@37400.4]
  assign _T_90033 = _T_90032[5:0]; // @[Modules.scala 150:103:@37401.4]
  assign _T_90034 = $signed(_T_90033); // @[Modules.scala 150:103:@37402.4]
  assign _T_90039 = $signed(_T_56124) + $signed(_T_65340); // @[Modules.scala 150:103:@37406.4]
  assign _T_90040 = _T_90039[4:0]; // @[Modules.scala 150:103:@37407.4]
  assign _T_90041 = $signed(_T_90040); // @[Modules.scala 150:103:@37408.4]
  assign _T_90046 = $signed(_T_65342) + $signed(_T_65347); // @[Modules.scala 150:103:@37412.4]
  assign _T_90047 = _T_90046[4:0]; // @[Modules.scala 150:103:@37413.4]
  assign _T_90048 = $signed(_T_90047); // @[Modules.scala 150:103:@37414.4]
  assign _T_90053 = $signed(_T_62231) + $signed(_T_56145); // @[Modules.scala 150:103:@37418.4]
  assign _T_90054 = _T_90053[4:0]; // @[Modules.scala 150:103:@37419.4]
  assign _T_90055 = $signed(_T_90054); // @[Modules.scala 150:103:@37420.4]
  assign _GEN_828 = {{1{_T_56154[4]}},_T_56154}; // @[Modules.scala 150:103:@37430.4]
  assign _T_90067 = $signed(_GEN_828) + $signed(_T_59166); // @[Modules.scala 150:103:@37430.4]
  assign _T_90068 = _T_90067[5:0]; // @[Modules.scala 150:103:@37431.4]
  assign _T_90069 = $signed(_T_90068); // @[Modules.scala 150:103:@37432.4]
  assign _T_90116 = $signed(_T_77802) + $signed(_T_65410); // @[Modules.scala 150:103:@37472.4]
  assign _T_90117 = _T_90116[4:0]; // @[Modules.scala 150:103:@37473.4]
  assign _T_90118 = $signed(_T_90117); // @[Modules.scala 150:103:@37474.4]
  assign _T_90172 = $signed(_GEN_562) + $signed(_T_59264); // @[Modules.scala 150:103:@37520.4]
  assign _T_90173 = _T_90172[5:0]; // @[Modules.scala 150:103:@37521.4]
  assign _T_90174 = $signed(_T_90173); // @[Modules.scala 150:103:@37522.4]
  assign _GEN_831 = {{1{_T_56259[4]}},_T_56259}; // @[Modules.scala 150:103:@37532.4]
  assign _T_90186 = $signed(_T_59276) + $signed(_GEN_831); // @[Modules.scala 150:103:@37532.4]
  assign _T_90187 = _T_90186[5:0]; // @[Modules.scala 150:103:@37533.4]
  assign _T_90188 = $signed(_T_90187); // @[Modules.scala 150:103:@37534.4]
  assign _T_90214 = $signed(_T_62392) + $signed(_T_62399); // @[Modules.scala 150:103:@37556.4]
  assign _T_90215 = _T_90214[4:0]; // @[Modules.scala 150:103:@37557.4]
  assign _T_90216 = $signed(_T_90215); // @[Modules.scala 150:103:@37558.4]
  assign buffer_11_0 = {{8{_T_88151[5]}},_T_88151}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_1 = {{8{_T_88158[5]}},_T_88158}; // @[Modules.scala 112:22:@8.4]
  assign _T_90233 = $signed(buffer_11_0) + $signed(buffer_11_1); // @[Modules.scala 166:64:@37574.4]
  assign _T_90234 = _T_90233[13:0]; // @[Modules.scala 166:64:@37575.4]
  assign buffer_11_299 = $signed(_T_90234); // @[Modules.scala 166:64:@37576.4]
  assign buffer_11_2 = {{8{_T_88165[5]}},_T_88165}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_3 = {{8{_T_88172[5]}},_T_88172}; // @[Modules.scala 112:22:@8.4]
  assign _T_90236 = $signed(buffer_11_2) + $signed(buffer_11_3); // @[Modules.scala 166:64:@37578.4]
  assign _T_90237 = _T_90236[13:0]; // @[Modules.scala 166:64:@37579.4]
  assign buffer_11_300 = $signed(_T_90237); // @[Modules.scala 166:64:@37580.4]
  assign _T_90239 = $signed(buffer_1_4) + $signed(buffer_5_6); // @[Modules.scala 166:64:@37582.4]
  assign _T_90240 = _T_90239[13:0]; // @[Modules.scala 166:64:@37583.4]
  assign buffer_11_301 = $signed(_T_90240); // @[Modules.scala 166:64:@37584.4]
  assign _T_90242 = $signed(buffer_2_6) + $signed(buffer_8_8); // @[Modules.scala 166:64:@37586.4]
  assign _T_90243 = _T_90242[13:0]; // @[Modules.scala 166:64:@37587.4]
  assign buffer_11_302 = $signed(_T_90243); // @[Modules.scala 166:64:@37588.4]
  assign buffer_11_8 = {{8{_T_88207[5]}},_T_88207}; // @[Modules.scala 112:22:@8.4]
  assign _T_90245 = $signed(buffer_11_8) + $signed(buffer_3_9); // @[Modules.scala 166:64:@37590.4]
  assign _T_90246 = _T_90245[13:0]; // @[Modules.scala 166:64:@37591.4]
  assign buffer_11_303 = $signed(_T_90246); // @[Modules.scala 166:64:@37592.4]
  assign buffer_11_11 = {{8{_T_88228[5]}},_T_88228}; // @[Modules.scala 112:22:@8.4]
  assign _T_90248 = $signed(buffer_4_9) + $signed(buffer_11_11); // @[Modules.scala 166:64:@37594.4]
  assign _T_90249 = _T_90248[13:0]; // @[Modules.scala 166:64:@37595.4]
  assign buffer_11_304 = $signed(_T_90249); // @[Modules.scala 166:64:@37596.4]
  assign _T_90263 = $signed(buffer_6_21) + $signed(buffer_3_20); // @[Modules.scala 166:64:@37614.4]
  assign _T_90264 = _T_90263[13:0]; // @[Modules.scala 166:64:@37615.4]
  assign buffer_11_309 = $signed(_T_90264); // @[Modules.scala 166:64:@37616.4]
  assign buffer_11_22 = {{8{_T_88305[5]}},_T_88305}; // @[Modules.scala 112:22:@8.4]
  assign _T_90266 = $signed(buffer_11_22) + $signed(buffer_1_22); // @[Modules.scala 166:64:@37618.4]
  assign _T_90267 = _T_90266[13:0]; // @[Modules.scala 166:64:@37619.4]
  assign buffer_11_310 = $signed(_T_90267); // @[Modules.scala 166:64:@37620.4]
  assign _T_90269 = $signed(buffer_2_22) + $signed(buffer_1_24); // @[Modules.scala 166:64:@37622.4]
  assign _T_90270 = _T_90269[13:0]; // @[Modules.scala 166:64:@37623.4]
  assign buffer_11_311 = $signed(_T_90270); // @[Modules.scala 166:64:@37624.4]
  assign _T_90272 = $signed(buffer_6_25) + $signed(buffer_1_26); // @[Modules.scala 166:64:@37626.4]
  assign _T_90273 = _T_90272[13:0]; // @[Modules.scala 166:64:@37627.4]
  assign buffer_11_312 = $signed(_T_90273); // @[Modules.scala 166:64:@37628.4]
  assign _T_90275 = $signed(buffer_1_27) + $signed(buffer_5_27); // @[Modules.scala 166:64:@37630.4]
  assign _T_90276 = _T_90275[13:0]; // @[Modules.scala 166:64:@37631.4]
  assign buffer_11_313 = $signed(_T_90276); // @[Modules.scala 166:64:@37632.4]
  assign buffer_11_34 = {{8{_T_88389[5]}},_T_88389}; // @[Modules.scala 112:22:@8.4]
  assign _T_90284 = $signed(buffer_11_34) + $signed(buffer_5_33); // @[Modules.scala 166:64:@37642.4]
  assign _T_90285 = _T_90284[13:0]; // @[Modules.scala 166:64:@37643.4]
  assign buffer_11_316 = $signed(_T_90285); // @[Modules.scala 166:64:@37644.4]
  assign _T_90287 = $signed(buffer_5_34) + $signed(buffer_3_36); // @[Modules.scala 166:64:@37646.4]
  assign _T_90288 = _T_90287[13:0]; // @[Modules.scala 166:64:@37647.4]
  assign buffer_11_317 = $signed(_T_90288); // @[Modules.scala 166:64:@37648.4]
  assign _T_90290 = $signed(buffer_4_37) + $signed(buffer_1_38); // @[Modules.scala 166:64:@37650.4]
  assign _T_90291 = _T_90290[13:0]; // @[Modules.scala 166:64:@37651.4]
  assign buffer_11_318 = $signed(_T_90291); // @[Modules.scala 166:64:@37652.4]
  assign _T_90293 = $signed(buffer_10_40) + $signed(buffer_0_42); // @[Modules.scala 166:64:@37654.4]
  assign _T_90294 = _T_90293[13:0]; // @[Modules.scala 166:64:@37655.4]
  assign buffer_11_319 = $signed(_T_90294); // @[Modules.scala 166:64:@37656.4]
  assign buffer_11_42 = {{8{_T_88445[5]}},_T_88445}; // @[Modules.scala 112:22:@8.4]
  assign _T_90296 = $signed(buffer_11_42) + $signed(buffer_5_43); // @[Modules.scala 166:64:@37658.4]
  assign _T_90297 = _T_90296[13:0]; // @[Modules.scala 166:64:@37659.4]
  assign buffer_11_320 = $signed(_T_90297); // @[Modules.scala 166:64:@37660.4]
  assign buffer_11_44 = {{8{_T_88459[5]}},_T_88459}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_45 = {{8{_T_88466[5]}},_T_88466}; // @[Modules.scala 112:22:@8.4]
  assign _T_90299 = $signed(buffer_11_44) + $signed(buffer_11_45); // @[Modules.scala 166:64:@37662.4]
  assign _T_90300 = _T_90299[13:0]; // @[Modules.scala 166:64:@37663.4]
  assign buffer_11_321 = $signed(_T_90300); // @[Modules.scala 166:64:@37664.4]
  assign _T_90302 = $signed(buffer_1_45) + $signed(buffer_1_46); // @[Modules.scala 166:64:@37666.4]
  assign _T_90303 = _T_90302[13:0]; // @[Modules.scala 166:64:@37667.4]
  assign buffer_11_322 = $signed(_T_90303); // @[Modules.scala 166:64:@37668.4]
  assign buffer_11_48 = {{8{_T_88487[5]}},_T_88487}; // @[Modules.scala 112:22:@8.4]
  assign _T_90305 = $signed(buffer_11_48) + $signed(buffer_8_47); // @[Modules.scala 166:64:@37670.4]
  assign _T_90306 = _T_90305[13:0]; // @[Modules.scala 166:64:@37671.4]
  assign buffer_11_323 = $signed(_T_90306); // @[Modules.scala 166:64:@37672.4]
  assign _T_90308 = $signed(buffer_1_49) + $signed(buffer_6_50); // @[Modules.scala 166:64:@37674.4]
  assign _T_90309 = _T_90308[13:0]; // @[Modules.scala 166:64:@37675.4]
  assign buffer_11_324 = $signed(_T_90309); // @[Modules.scala 166:64:@37676.4]
  assign _T_90311 = $signed(buffer_0_50) + $signed(buffer_1_53); // @[Modules.scala 166:64:@37678.4]
  assign _T_90312 = _T_90311[13:0]; // @[Modules.scala 166:64:@37679.4]
  assign buffer_11_325 = $signed(_T_90312); // @[Modules.scala 166:64:@37680.4]
  assign _T_90314 = $signed(buffer_5_55) + $signed(buffer_3_57); // @[Modules.scala 166:64:@37682.4]
  assign _T_90315 = _T_90314[13:0]; // @[Modules.scala 166:64:@37683.4]
  assign buffer_11_326 = $signed(_T_90315); // @[Modules.scala 166:64:@37684.4]
  assign buffer_11_56 = {{8{_T_88543[5]}},_T_88543}; // @[Modules.scala 112:22:@8.4]
  assign _T_90317 = $signed(buffer_11_56) + $signed(buffer_6_56); // @[Modules.scala 166:64:@37686.4]
  assign _T_90318 = _T_90317[13:0]; // @[Modules.scala 166:64:@37687.4]
  assign buffer_11_327 = $signed(_T_90318); // @[Modules.scala 166:64:@37688.4]
  assign buffer_11_59 = {{8{_T_88564[5]}},_T_88564}; // @[Modules.scala 112:22:@8.4]
  assign _T_90320 = $signed(buffer_6_57) + $signed(buffer_11_59); // @[Modules.scala 166:64:@37690.4]
  assign _T_90321 = _T_90320[13:0]; // @[Modules.scala 166:64:@37691.4]
  assign buffer_11_328 = $signed(_T_90321); // @[Modules.scala 166:64:@37692.4]
  assign _T_90323 = $signed(buffer_6_60) + $signed(buffer_5_63); // @[Modules.scala 166:64:@37694.4]
  assign _T_90324 = _T_90323[13:0]; // @[Modules.scala 166:64:@37695.4]
  assign buffer_11_329 = $signed(_T_90324); // @[Modules.scala 166:64:@37696.4]
  assign buffer_11_62 = {{8{_T_88585[5]}},_T_88585}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_63 = {{9{_T_88592[4]}},_T_88592}; // @[Modules.scala 112:22:@8.4]
  assign _T_90326 = $signed(buffer_11_62) + $signed(buffer_11_63); // @[Modules.scala 166:64:@37698.4]
  assign _T_90327 = _T_90326[13:0]; // @[Modules.scala 166:64:@37699.4]
  assign buffer_11_330 = $signed(_T_90327); // @[Modules.scala 166:64:@37700.4]
  assign buffer_11_64 = {{8{_T_88599[5]}},_T_88599}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_65 = {{9{_T_88606[4]}},_T_88606}; // @[Modules.scala 112:22:@8.4]
  assign _T_90329 = $signed(buffer_11_64) + $signed(buffer_11_65); // @[Modules.scala 166:64:@37702.4]
  assign _T_90330 = _T_90329[13:0]; // @[Modules.scala 166:64:@37703.4]
  assign buffer_11_331 = $signed(_T_90330); // @[Modules.scala 166:64:@37704.4]
  assign buffer_11_67 = {{8{_T_88620[5]}},_T_88620}; // @[Modules.scala 112:22:@8.4]
  assign _T_90332 = $signed(buffer_0_67) + $signed(buffer_11_67); // @[Modules.scala 166:64:@37706.4]
  assign _T_90333 = _T_90332[13:0]; // @[Modules.scala 166:64:@37707.4]
  assign buffer_11_332 = $signed(_T_90333); // @[Modules.scala 166:64:@37708.4]
  assign buffer_11_70 = {{8{_T_88641[5]}},_T_88641}; // @[Modules.scala 112:22:@8.4]
  assign _T_90338 = $signed(buffer_11_70) + $signed(buffer_1_75); // @[Modules.scala 166:64:@37714.4]
  assign _T_90339 = _T_90338[13:0]; // @[Modules.scala 166:64:@37715.4]
  assign buffer_11_334 = $signed(_T_90339); // @[Modules.scala 166:64:@37716.4]
  assign buffer_11_72 = {{8{_T_88655[5]}},_T_88655}; // @[Modules.scala 112:22:@8.4]
  assign _T_90341 = $signed(buffer_11_72) + $signed(buffer_0_74); // @[Modules.scala 166:64:@37718.4]
  assign _T_90342 = _T_90341[13:0]; // @[Modules.scala 166:64:@37719.4]
  assign buffer_11_335 = $signed(_T_90342); // @[Modules.scala 166:64:@37720.4]
  assign _T_90344 = $signed(buffer_7_77) + $signed(buffer_10_77); // @[Modules.scala 166:64:@37722.4]
  assign _T_90345 = _T_90344[13:0]; // @[Modules.scala 166:64:@37723.4]
  assign buffer_11_336 = $signed(_T_90345); // @[Modules.scala 166:64:@37724.4]
  assign buffer_11_76 = {{9{_T_88683[4]}},_T_88683}; // @[Modules.scala 112:22:@8.4]
  assign _T_90347 = $signed(buffer_11_76) + $signed(buffer_2_82); // @[Modules.scala 166:64:@37726.4]
  assign _T_90348 = _T_90347[13:0]; // @[Modules.scala 166:64:@37727.4]
  assign buffer_11_337 = $signed(_T_90348); // @[Modules.scala 166:64:@37728.4]
  assign buffer_11_78 = {{8{_T_88697[5]}},_T_88697}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_79 = {{8{_T_88704[5]}},_T_88704}; // @[Modules.scala 112:22:@8.4]
  assign _T_90350 = $signed(buffer_11_78) + $signed(buffer_11_79); // @[Modules.scala 166:64:@37730.4]
  assign _T_90351 = _T_90350[13:0]; // @[Modules.scala 166:64:@37731.4]
  assign buffer_11_338 = $signed(_T_90351); // @[Modules.scala 166:64:@37732.4]
  assign buffer_11_80 = {{8{_T_88711[5]}},_T_88711}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_81 = {{8{_T_88718[5]}},_T_88718}; // @[Modules.scala 112:22:@8.4]
  assign _T_90353 = $signed(buffer_11_80) + $signed(buffer_11_81); // @[Modules.scala 166:64:@37734.4]
  assign _T_90354 = _T_90353[13:0]; // @[Modules.scala 166:64:@37735.4]
  assign buffer_11_339 = $signed(_T_90354); // @[Modules.scala 166:64:@37736.4]
  assign buffer_11_83 = {{8{_T_88732[5]}},_T_88732}; // @[Modules.scala 112:22:@8.4]
  assign _T_90356 = $signed(buffer_2_89) + $signed(buffer_11_83); // @[Modules.scala 166:64:@37738.4]
  assign _T_90357 = _T_90356[13:0]; // @[Modules.scala 166:64:@37739.4]
  assign buffer_11_340 = $signed(_T_90357); // @[Modules.scala 166:64:@37740.4]
  assign _T_90359 = $signed(buffer_0_87) + $signed(buffer_3_93); // @[Modules.scala 166:64:@37742.4]
  assign _T_90360 = _T_90359[13:0]; // @[Modules.scala 166:64:@37743.4]
  assign buffer_11_341 = $signed(_T_90360); // @[Modules.scala 166:64:@37744.4]
  assign buffer_11_88 = {{9{_T_88767[4]}},_T_88767}; // @[Modules.scala 112:22:@8.4]
  assign _T_90365 = $signed(buffer_11_88) + $signed(buffer_0_91); // @[Modules.scala 166:64:@37750.4]
  assign _T_90366 = _T_90365[13:0]; // @[Modules.scala 166:64:@37751.4]
  assign buffer_11_343 = $signed(_T_90366); // @[Modules.scala 166:64:@37752.4]
  assign buffer_11_91 = {{8{_T_88788[5]}},_T_88788}; // @[Modules.scala 112:22:@8.4]
  assign _T_90368 = $signed(buffer_3_98) + $signed(buffer_11_91); // @[Modules.scala 166:64:@37754.4]
  assign _T_90369 = _T_90368[13:0]; // @[Modules.scala 166:64:@37755.4]
  assign buffer_11_344 = $signed(_T_90369); // @[Modules.scala 166:64:@37756.4]
  assign buffer_11_93 = {{8{_T_88802[5]}},_T_88802}; // @[Modules.scala 112:22:@8.4]
  assign _T_90371 = $signed(buffer_4_96) + $signed(buffer_11_93); // @[Modules.scala 166:64:@37758.4]
  assign _T_90372 = _T_90371[13:0]; // @[Modules.scala 166:64:@37759.4]
  assign buffer_11_345 = $signed(_T_90372); // @[Modules.scala 166:64:@37760.4]
  assign buffer_11_95 = {{9{_T_88816[4]}},_T_88816}; // @[Modules.scala 112:22:@8.4]
  assign _T_90374 = $signed(buffer_0_97) + $signed(buffer_11_95); // @[Modules.scala 166:64:@37762.4]
  assign _T_90375 = _T_90374[13:0]; // @[Modules.scala 166:64:@37763.4]
  assign buffer_11_346 = $signed(_T_90375); // @[Modules.scala 166:64:@37764.4]
  assign buffer_11_98 = {{9{_T_88837[4]}},_T_88837}; // @[Modules.scala 112:22:@8.4]
  assign _T_90380 = $signed(buffer_11_98) + $signed(buffer_1_106); // @[Modules.scala 166:64:@37770.4]
  assign _T_90381 = _T_90380[13:0]; // @[Modules.scala 166:64:@37771.4]
  assign buffer_11_348 = $signed(_T_90381); // @[Modules.scala 166:64:@37772.4]
  assign buffer_11_101 = {{8{_T_88858[5]}},_T_88858}; // @[Modules.scala 112:22:@8.4]
  assign _T_90383 = $signed(buffer_9_113) + $signed(buffer_11_101); // @[Modules.scala 166:64:@37774.4]
  assign _T_90384 = _T_90383[13:0]; // @[Modules.scala 166:64:@37775.4]
  assign buffer_11_349 = $signed(_T_90384); // @[Modules.scala 166:64:@37776.4]
  assign _T_90386 = $signed(buffer_1_109) + $signed(buffer_1_110); // @[Modules.scala 166:64:@37778.4]
  assign _T_90387 = _T_90386[13:0]; // @[Modules.scala 166:64:@37779.4]
  assign buffer_11_350 = $signed(_T_90387); // @[Modules.scala 166:64:@37780.4]
  assign _T_90389 = $signed(buffer_1_111) + $signed(buffer_4_110); // @[Modules.scala 166:64:@37782.4]
  assign _T_90390 = _T_90389[13:0]; // @[Modules.scala 166:64:@37783.4]
  assign buffer_11_351 = $signed(_T_90390); // @[Modules.scala 166:64:@37784.4]
  assign _T_90392 = $signed(buffer_0_111) + $signed(buffer_4_112); // @[Modules.scala 166:64:@37786.4]
  assign _T_90393 = _T_90392[13:0]; // @[Modules.scala 166:64:@37787.4]
  assign buffer_11_352 = $signed(_T_90393); // @[Modules.scala 166:64:@37788.4]
  assign _T_90395 = $signed(buffer_9_120) + $signed(buffer_10_115); // @[Modules.scala 166:64:@37790.4]
  assign _T_90396 = _T_90395[13:0]; // @[Modules.scala 166:64:@37791.4]
  assign buffer_11_353 = $signed(_T_90396); // @[Modules.scala 166:64:@37792.4]
  assign buffer_11_113 = {{9{_T_88942[4]}},_T_88942}; // @[Modules.scala 112:22:@8.4]
  assign _T_90401 = $signed(buffer_1_119) + $signed(buffer_11_113); // @[Modules.scala 166:64:@37798.4]
  assign _T_90402 = _T_90401[13:0]; // @[Modules.scala 166:64:@37799.4]
  assign buffer_11_355 = $signed(_T_90402); // @[Modules.scala 166:64:@37800.4]
  assign _T_90404 = $signed(buffer_1_121) + $signed(buffer_1_122); // @[Modules.scala 166:64:@37802.4]
  assign _T_90405 = _T_90404[13:0]; // @[Modules.scala 166:64:@37803.4]
  assign buffer_11_356 = $signed(_T_90405); // @[Modules.scala 166:64:@37804.4]
  assign _T_90407 = $signed(buffer_1_123) + $signed(buffer_1_124); // @[Modules.scala 166:64:@37806.4]
  assign _T_90408 = _T_90407[13:0]; // @[Modules.scala 166:64:@37807.4]
  assign buffer_11_357 = $signed(_T_90408); // @[Modules.scala 166:64:@37808.4]
  assign buffer_11_118 = {{8{_T_88977[5]}},_T_88977}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_119 = {{8{_T_88984[5]}},_T_88984}; // @[Modules.scala 112:22:@8.4]
  assign _T_90410 = $signed(buffer_11_118) + $signed(buffer_11_119); // @[Modules.scala 166:64:@37810.4]
  assign _T_90411 = _T_90410[13:0]; // @[Modules.scala 166:64:@37811.4]
  assign buffer_11_358 = $signed(_T_90411); // @[Modules.scala 166:64:@37812.4]
  assign _T_90413 = $signed(buffer_4_123) + $signed(buffer_0_125); // @[Modules.scala 166:64:@37814.4]
  assign _T_90414 = _T_90413[13:0]; // @[Modules.scala 166:64:@37815.4]
  assign buffer_11_359 = $signed(_T_90414); // @[Modules.scala 166:64:@37816.4]
  assign _T_90419 = $signed(buffer_0_130) + $signed(buffer_10_132); // @[Modules.scala 166:64:@37822.4]
  assign _T_90420 = _T_90419[13:0]; // @[Modules.scala 166:64:@37823.4]
  assign buffer_11_361 = $signed(_T_90420); // @[Modules.scala 166:64:@37824.4]
  assign _T_90422 = $signed(buffer_0_132) + $signed(buffer_6_136); // @[Modules.scala 166:64:@37826.4]
  assign _T_90423 = _T_90422[13:0]; // @[Modules.scala 166:64:@37827.4]
  assign buffer_11_362 = $signed(_T_90423); // @[Modules.scala 166:64:@37828.4]
  assign buffer_11_128 = {{8{_T_89047[5]}},_T_89047}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_129 = {{8{_T_89054[5]}},_T_89054}; // @[Modules.scala 112:22:@8.4]
  assign _T_90425 = $signed(buffer_11_128) + $signed(buffer_11_129); // @[Modules.scala 166:64:@37830.4]
  assign _T_90426 = _T_90425[13:0]; // @[Modules.scala 166:64:@37831.4]
  assign buffer_11_363 = $signed(_T_90426); // @[Modules.scala 166:64:@37832.4]
  assign buffer_11_131 = {{8{_T_89068[5]}},_T_89068}; // @[Modules.scala 112:22:@8.4]
  assign _T_90428 = $signed(buffer_0_135) + $signed(buffer_11_131); // @[Modules.scala 166:64:@37834.4]
  assign _T_90429 = _T_90428[13:0]; // @[Modules.scala 166:64:@37835.4]
  assign buffer_11_364 = $signed(_T_90429); // @[Modules.scala 166:64:@37836.4]
  assign buffer_11_132 = {{8{_T_89075[5]}},_T_89075}; // @[Modules.scala 112:22:@8.4]
  assign _T_90431 = $signed(buffer_11_132) + $signed(buffer_0_138); // @[Modules.scala 166:64:@37838.4]
  assign _T_90432 = _T_90431[13:0]; // @[Modules.scala 166:64:@37839.4]
  assign buffer_11_365 = $signed(_T_90432); // @[Modules.scala 166:64:@37840.4]
  assign _T_90434 = $signed(buffer_4_137) + $signed(buffer_5_143); // @[Modules.scala 166:64:@37842.4]
  assign _T_90435 = _T_90434[13:0]; // @[Modules.scala 166:64:@37843.4]
  assign buffer_11_366 = $signed(_T_90435); // @[Modules.scala 166:64:@37844.4]
  assign buffer_11_136 = {{9{_T_89103[4]}},_T_89103}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_137 = {{8{_T_89110[5]}},_T_89110}; // @[Modules.scala 112:22:@8.4]
  assign _T_90437 = $signed(buffer_11_136) + $signed(buffer_11_137); // @[Modules.scala 166:64:@37846.4]
  assign _T_90438 = _T_90437[13:0]; // @[Modules.scala 166:64:@37847.4]
  assign buffer_11_367 = $signed(_T_90438); // @[Modules.scala 166:64:@37848.4]
  assign _T_90443 = $signed(buffer_2_150) + $signed(buffer_5_147); // @[Modules.scala 166:64:@37854.4]
  assign _T_90444 = _T_90443[13:0]; // @[Modules.scala 166:64:@37855.4]
  assign buffer_11_369 = $signed(_T_90444); // @[Modules.scala 166:64:@37856.4]
  assign buffer_11_145 = {{9{_T_89166[4]}},_T_89166}; // @[Modules.scala 112:22:@8.4]
  assign _T_90449 = $signed(buffer_5_150) + $signed(buffer_11_145); // @[Modules.scala 166:64:@37862.4]
  assign _T_90450 = _T_90449[13:0]; // @[Modules.scala 166:64:@37863.4]
  assign buffer_11_371 = $signed(_T_90450); // @[Modules.scala 166:64:@37864.4]
  assign _T_90455 = $signed(buffer_5_154) + $signed(buffer_8_153); // @[Modules.scala 166:64:@37870.4]
  assign _T_90456 = _T_90455[13:0]; // @[Modules.scala 166:64:@37871.4]
  assign buffer_11_373 = $signed(_T_90456); // @[Modules.scala 166:64:@37872.4]
  assign buffer_11_153 = {{8{_T_89222[5]}},_T_89222}; // @[Modules.scala 112:22:@8.4]
  assign _T_90461 = $signed(buffer_8_156) + $signed(buffer_11_153); // @[Modules.scala 166:64:@37878.4]
  assign _T_90462 = _T_90461[13:0]; // @[Modules.scala 166:64:@37879.4]
  assign buffer_11_375 = $signed(_T_90462); // @[Modules.scala 166:64:@37880.4]
  assign buffer_11_156 = {{8{_T_89243[5]}},_T_89243}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_157 = {{8{_T_89250[5]}},_T_89250}; // @[Modules.scala 112:22:@8.4]
  assign _T_90467 = $signed(buffer_11_156) + $signed(buffer_11_157); // @[Modules.scala 166:64:@37886.4]
  assign _T_90468 = _T_90467[13:0]; // @[Modules.scala 166:64:@37887.4]
  assign buffer_11_377 = $signed(_T_90468); // @[Modules.scala 166:64:@37888.4]
  assign buffer_11_159 = {{8{_T_89264[5]}},_T_89264}; // @[Modules.scala 112:22:@8.4]
  assign _T_90470 = $signed(buffer_7_164) + $signed(buffer_11_159); // @[Modules.scala 166:64:@37890.4]
  assign _T_90471 = _T_90470[13:0]; // @[Modules.scala 166:64:@37891.4]
  assign buffer_11_378 = $signed(_T_90471); // @[Modules.scala 166:64:@37892.4]
  assign buffer_11_161 = {{8{_T_89278[5]}},_T_89278}; // @[Modules.scala 112:22:@8.4]
  assign _T_90473 = $signed(buffer_5_167) + $signed(buffer_11_161); // @[Modules.scala 166:64:@37894.4]
  assign _T_90474 = _T_90473[13:0]; // @[Modules.scala 166:64:@37895.4]
  assign buffer_11_379 = $signed(_T_90474); // @[Modules.scala 166:64:@37896.4]
  assign buffer_11_162 = {{8{_T_89285[5]}},_T_89285}; // @[Modules.scala 112:22:@8.4]
  assign _T_90476 = $signed(buffer_11_162) + $signed(buffer_0_167); // @[Modules.scala 166:64:@37898.4]
  assign _T_90477 = _T_90476[13:0]; // @[Modules.scala 166:64:@37899.4]
  assign buffer_11_380 = $signed(_T_90477); // @[Modules.scala 166:64:@37900.4]
  assign _T_90479 = $signed(buffer_8_167) + $signed(buffer_4_165); // @[Modules.scala 166:64:@37902.4]
  assign _T_90480 = _T_90479[13:0]; // @[Modules.scala 166:64:@37903.4]
  assign buffer_11_381 = $signed(_T_90480); // @[Modules.scala 166:64:@37904.4]
  assign buffer_11_169 = {{8{_T_89334[5]}},_T_89334}; // @[Modules.scala 112:22:@8.4]
  assign _T_90485 = $signed(buffer_1_171) + $signed(buffer_11_169); // @[Modules.scala 166:64:@37910.4]
  assign _T_90486 = _T_90485[13:0]; // @[Modules.scala 166:64:@37911.4]
  assign buffer_11_383 = $signed(_T_90486); // @[Modules.scala 166:64:@37912.4]
  assign buffer_11_170 = {{8{_T_89341[5]}},_T_89341}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_171 = {{8{_T_89348[5]}},_T_89348}; // @[Modules.scala 112:22:@8.4]
  assign _T_90488 = $signed(buffer_11_170) + $signed(buffer_11_171); // @[Modules.scala 166:64:@37914.4]
  assign _T_90489 = _T_90488[13:0]; // @[Modules.scala 166:64:@37915.4]
  assign buffer_11_384 = $signed(_T_90489); // @[Modules.scala 166:64:@37916.4]
  assign _T_90491 = $signed(buffer_6_183) + $signed(buffer_0_178); // @[Modules.scala 166:64:@37918.4]
  assign _T_90492 = _T_90491[13:0]; // @[Modules.scala 166:64:@37919.4]
  assign buffer_11_385 = $signed(_T_90492); // @[Modules.scala 166:64:@37920.4]
  assign _T_90494 = $signed(buffer_6_185) + $signed(buffer_8_180); // @[Modules.scala 166:64:@37922.4]
  assign _T_90495 = _T_90494[13:0]; // @[Modules.scala 166:64:@37923.4]
  assign buffer_11_386 = $signed(_T_90495); // @[Modules.scala 166:64:@37924.4]
  assign buffer_11_176 = {{8{_T_89383[5]}},_T_89383}; // @[Modules.scala 112:22:@8.4]
  assign _T_90497 = $signed(buffer_11_176) + $signed(buffer_3_189); // @[Modules.scala 166:64:@37926.4]
  assign _T_90498 = _T_90497[13:0]; // @[Modules.scala 166:64:@37927.4]
  assign buffer_11_387 = $signed(_T_90498); // @[Modules.scala 166:64:@37928.4]
  assign _T_90503 = $signed(buffer_7_189) + $signed(buffer_1_184); // @[Modules.scala 166:64:@37934.4]
  assign _T_90504 = _T_90503[13:0]; // @[Modules.scala 166:64:@37935.4]
  assign buffer_11_389 = $signed(_T_90504); // @[Modules.scala 166:64:@37936.4]
  assign _T_90509 = $signed(buffer_6_195) + $signed(buffer_4_181); // @[Modules.scala 166:64:@37942.4]
  assign _T_90510 = _T_90509[13:0]; // @[Modules.scala 166:64:@37943.4]
  assign buffer_11_391 = $signed(_T_90510); // @[Modules.scala 166:64:@37944.4]
  assign buffer_11_186 = {{8{_T_89453[5]}},_T_89453}; // @[Modules.scala 112:22:@8.4]
  assign _T_90512 = $signed(buffer_11_186) + $signed(buffer_0_188); // @[Modules.scala 166:64:@37946.4]
  assign _T_90513 = _T_90512[13:0]; // @[Modules.scala 166:64:@37947.4]
  assign buffer_11_392 = $signed(_T_90513); // @[Modules.scala 166:64:@37948.4]
  assign _T_90515 = $signed(buffer_0_189) + $signed(buffer_10_198); // @[Modules.scala 166:64:@37950.4]
  assign _T_90516 = _T_90515[13:0]; // @[Modules.scala 166:64:@37951.4]
  assign buffer_11_393 = $signed(_T_90516); // @[Modules.scala 166:64:@37952.4]
  assign buffer_11_191 = {{8{_T_89488[5]}},_T_89488}; // @[Modules.scala 112:22:@8.4]
  assign _T_90518 = $signed(buffer_7_200) + $signed(buffer_11_191); // @[Modules.scala 166:64:@37954.4]
  assign _T_90519 = _T_90518[13:0]; // @[Modules.scala 166:64:@37955.4]
  assign buffer_11_394 = $signed(_T_90519); // @[Modules.scala 166:64:@37956.4]
  assign buffer_11_195 = {{8{_T_89516[5]}},_T_89516}; // @[Modules.scala 112:22:@8.4]
  assign _T_90524 = $signed(buffer_8_199) + $signed(buffer_11_195); // @[Modules.scala 166:64:@37962.4]
  assign _T_90525 = _T_90524[13:0]; // @[Modules.scala 166:64:@37963.4]
  assign buffer_11_396 = $signed(_T_90525); // @[Modules.scala 166:64:@37964.4]
  assign buffer_11_196 = {{8{_T_89523[5]}},_T_89523}; // @[Modules.scala 112:22:@8.4]
  assign _T_90527 = $signed(buffer_11_196) + $signed(buffer_0_199); // @[Modules.scala 166:64:@37966.4]
  assign _T_90528 = _T_90527[13:0]; // @[Modules.scala 166:64:@37967.4]
  assign buffer_11_397 = $signed(_T_90528); // @[Modules.scala 166:64:@37968.4]
  assign buffer_11_199 = {{8{_T_89544[5]}},_T_89544}; // @[Modules.scala 112:22:@8.4]
  assign _T_90530 = $signed(buffer_0_200) + $signed(buffer_11_199); // @[Modules.scala 166:64:@37970.4]
  assign _T_90531 = _T_90530[13:0]; // @[Modules.scala 166:64:@37971.4]
  assign buffer_11_398 = $signed(_T_90531); // @[Modules.scala 166:64:@37972.4]
  assign buffer_11_201 = {{9{_T_89558[4]}},_T_89558}; // @[Modules.scala 112:22:@8.4]
  assign _T_90533 = $signed(buffer_7_211) + $signed(buffer_11_201); // @[Modules.scala 166:64:@37974.4]
  assign _T_90534 = _T_90533[13:0]; // @[Modules.scala 166:64:@37975.4]
  assign buffer_11_399 = $signed(_T_90534); // @[Modules.scala 166:64:@37976.4]
  assign buffer_11_202 = {{8{_T_89565[5]}},_T_89565}; // @[Modules.scala 112:22:@8.4]
  assign _T_90536 = $signed(buffer_11_202) + $signed(buffer_0_205); // @[Modules.scala 166:64:@37978.4]
  assign _T_90537 = _T_90536[13:0]; // @[Modules.scala 166:64:@37979.4]
  assign buffer_11_400 = $signed(_T_90537); // @[Modules.scala 166:64:@37980.4]
  assign buffer_11_204 = {{8{_T_89579[5]}},_T_89579}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_205 = {{9{_T_89586[4]}},_T_89586}; // @[Modules.scala 112:22:@8.4]
  assign _T_90539 = $signed(buffer_11_204) + $signed(buffer_11_205); // @[Modules.scala 166:64:@37982.4]
  assign _T_90540 = _T_90539[13:0]; // @[Modules.scala 166:64:@37983.4]
  assign buffer_11_401 = $signed(_T_90540); // @[Modules.scala 166:64:@37984.4]
  assign buffer_11_207 = {{8{_T_89600[5]}},_T_89600}; // @[Modules.scala 112:22:@8.4]
  assign _T_90542 = $signed(buffer_1_208) + $signed(buffer_11_207); // @[Modules.scala 166:64:@37986.4]
  assign _T_90543 = _T_90542[13:0]; // @[Modules.scala 166:64:@37987.4]
  assign buffer_11_402 = $signed(_T_90543); // @[Modules.scala 166:64:@37988.4]
  assign buffer_11_208 = {{8{_T_89607[5]}},_T_89607}; // @[Modules.scala 112:22:@8.4]
  assign _T_90545 = $signed(buffer_11_208) + $signed(buffer_1_211); // @[Modules.scala 166:64:@37990.4]
  assign _T_90546 = _T_90545[13:0]; // @[Modules.scala 166:64:@37991.4]
  assign buffer_11_403 = $signed(_T_90546); // @[Modules.scala 166:64:@37992.4]
  assign buffer_11_212 = {{9{_T_89635[4]}},_T_89635}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_213 = {{9{_T_89642[4]}},_T_89642}; // @[Modules.scala 112:22:@8.4]
  assign _T_90551 = $signed(buffer_11_212) + $signed(buffer_11_213); // @[Modules.scala 166:64:@37998.4]
  assign _T_90552 = _T_90551[13:0]; // @[Modules.scala 166:64:@37999.4]
  assign buffer_11_405 = $signed(_T_90552); // @[Modules.scala 166:64:@38000.4]
  assign buffer_11_219 = {{8{_T_89684[5]}},_T_89684}; // @[Modules.scala 112:22:@8.4]
  assign _T_90560 = $signed(buffer_1_220) + $signed(buffer_11_219); // @[Modules.scala 166:64:@38010.4]
  assign _T_90561 = _T_90560[13:0]; // @[Modules.scala 166:64:@38011.4]
  assign buffer_11_408 = $signed(_T_90561); // @[Modules.scala 166:64:@38012.4]
  assign _T_90563 = $signed(buffer_2_227) + $signed(buffer_3_233); // @[Modules.scala 166:64:@38014.4]
  assign _T_90564 = _T_90563[13:0]; // @[Modules.scala 166:64:@38015.4]
  assign buffer_11_409 = $signed(_T_90564); // @[Modules.scala 166:64:@38016.4]
  assign buffer_11_223 = {{9{_T_89712[4]}},_T_89712}; // @[Modules.scala 112:22:@8.4]
  assign _T_90566 = $signed(buffer_3_234) + $signed(buffer_11_223); // @[Modules.scala 166:64:@38018.4]
  assign _T_90567 = _T_90566[13:0]; // @[Modules.scala 166:64:@38019.4]
  assign buffer_11_410 = $signed(_T_90567); // @[Modules.scala 166:64:@38020.4]
  assign _T_90569 = $signed(buffer_5_230) + $signed(buffer_7_236); // @[Modules.scala 166:64:@38022.4]
  assign _T_90570 = _T_90569[13:0]; // @[Modules.scala 166:64:@38023.4]
  assign buffer_11_411 = $signed(_T_90570); // @[Modules.scala 166:64:@38024.4]
  assign _T_90572 = $signed(buffer_7_237) + $signed(buffer_7_238); // @[Modules.scala 166:64:@38026.4]
  assign _T_90573 = _T_90572[13:0]; // @[Modules.scala 166:64:@38027.4]
  assign buffer_11_412 = $signed(_T_90573); // @[Modules.scala 166:64:@38028.4]
  assign _T_90575 = $signed(buffer_0_227) + $signed(buffer_6_241); // @[Modules.scala 166:64:@38030.4]
  assign _T_90576 = _T_90575[13:0]; // @[Modules.scala 166:64:@38031.4]
  assign buffer_11_413 = $signed(_T_90576); // @[Modules.scala 166:64:@38032.4]
  assign buffer_11_231 = {{8{_T_89768[5]}},_T_89768}; // @[Modules.scala 112:22:@8.4]
  assign _T_90578 = $signed(buffer_0_229) + $signed(buffer_11_231); // @[Modules.scala 166:64:@38034.4]
  assign _T_90579 = _T_90578[13:0]; // @[Modules.scala 166:64:@38035.4]
  assign buffer_11_414 = $signed(_T_90579); // @[Modules.scala 166:64:@38036.4]
  assign buffer_11_232 = {{9{_T_89775[4]}},_T_89775}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_233 = {{9{_T_89782[4]}},_T_89782}; // @[Modules.scala 112:22:@8.4]
  assign _T_90581 = $signed(buffer_11_232) + $signed(buffer_11_233); // @[Modules.scala 166:64:@38038.4]
  assign _T_90582 = _T_90581[13:0]; // @[Modules.scala 166:64:@38039.4]
  assign buffer_11_415 = $signed(_T_90582); // @[Modules.scala 166:64:@38040.4]
  assign buffer_11_235 = {{9{_T_89796[4]}},_T_89796}; // @[Modules.scala 112:22:@8.4]
  assign _T_90584 = $signed(buffer_6_244) + $signed(buffer_11_235); // @[Modules.scala 166:64:@38042.4]
  assign _T_90585 = _T_90584[13:0]; // @[Modules.scala 166:64:@38043.4]
  assign buffer_11_416 = $signed(_T_90585); // @[Modules.scala 166:64:@38044.4]
  assign buffer_11_236 = {{8{_T_89803[5]}},_T_89803}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_237 = {{8{_T_89810[5]}},_T_89810}; // @[Modules.scala 112:22:@8.4]
  assign _T_90587 = $signed(buffer_11_236) + $signed(buffer_11_237); // @[Modules.scala 166:64:@38046.4]
  assign _T_90588 = _T_90587[13:0]; // @[Modules.scala 166:64:@38047.4]
  assign buffer_11_417 = $signed(_T_90588); // @[Modules.scala 166:64:@38048.4]
  assign buffer_11_238 = {{8{_T_89817[5]}},_T_89817}; // @[Modules.scala 112:22:@8.4]
  assign _T_90590 = $signed(buffer_11_238) + $signed(buffer_6_251); // @[Modules.scala 166:64:@38050.4]
  assign _T_90591 = _T_90590[13:0]; // @[Modules.scala 166:64:@38051.4]
  assign buffer_11_418 = $signed(_T_90591); // @[Modules.scala 166:64:@38052.4]
  assign buffer_11_241 = {{8{_T_89838[5]}},_T_89838}; // @[Modules.scala 112:22:@8.4]
  assign _T_90593 = $signed(buffer_6_252) + $signed(buffer_11_241); // @[Modules.scala 166:64:@38054.4]
  assign _T_90594 = _T_90593[13:0]; // @[Modules.scala 166:64:@38055.4]
  assign buffer_11_419 = $signed(_T_90594); // @[Modules.scala 166:64:@38056.4]
  assign buffer_11_242 = {{9{_T_89845[4]}},_T_89845}; // @[Modules.scala 112:22:@8.4]
  assign _T_90596 = $signed(buffer_11_242) + $signed(buffer_4_239); // @[Modules.scala 166:64:@38058.4]
  assign _T_90597 = _T_90596[13:0]; // @[Modules.scala 166:64:@38059.4]
  assign buffer_11_420 = $signed(_T_90597); // @[Modules.scala 166:64:@38060.4]
  assign buffer_11_244 = {{8{_T_89859[5]}},_T_89859}; // @[Modules.scala 112:22:@8.4]
  assign _T_90599 = $signed(buffer_11_244) + $signed(buffer_4_242); // @[Modules.scala 166:64:@38062.4]
  assign _T_90600 = _T_90599[13:0]; // @[Modules.scala 166:64:@38063.4]
  assign buffer_11_421 = $signed(_T_90600); // @[Modules.scala 166:64:@38064.4]
  assign _T_90602 = $signed(buffer_0_247) + $signed(buffer_0_248); // @[Modules.scala 166:64:@38066.4]
  assign _T_90603 = _T_90602[13:0]; // @[Modules.scala 166:64:@38067.4]
  assign buffer_11_422 = $signed(_T_90603); // @[Modules.scala 166:64:@38068.4]
  assign buffer_11_248 = {{8{_T_89887[5]}},_T_89887}; // @[Modules.scala 112:22:@8.4]
  assign _T_90605 = $signed(buffer_11_248) + $signed(buffer_5_259); // @[Modules.scala 166:64:@38070.4]
  assign _T_90606 = _T_90605[13:0]; // @[Modules.scala 166:64:@38071.4]
  assign buffer_11_423 = $signed(_T_90606); // @[Modules.scala 166:64:@38072.4]
  assign _T_90608 = $signed(buffer_6_263) + $signed(buffer_5_261); // @[Modules.scala 166:64:@38074.4]
  assign _T_90609 = _T_90608[13:0]; // @[Modules.scala 166:64:@38075.4]
  assign buffer_11_424 = $signed(_T_90609); // @[Modules.scala 166:64:@38076.4]
  assign _T_90611 = $signed(buffer_7_262) + $signed(buffer_6_265); // @[Modules.scala 166:64:@38078.4]
  assign _T_90612 = _T_90611[13:0]; // @[Modules.scala 166:64:@38079.4]
  assign buffer_11_425 = $signed(_T_90612); // @[Modules.scala 166:64:@38080.4]
  assign buffer_11_254 = {{8{_T_89929[5]}},_T_89929}; // @[Modules.scala 112:22:@8.4]
  assign _T_90614 = $signed(buffer_11_254) + $signed(buffer_6_270); // @[Modules.scala 166:64:@38082.4]
  assign _T_90615 = _T_90614[13:0]; // @[Modules.scala 166:64:@38083.4]
  assign buffer_11_426 = $signed(_T_90615); // @[Modules.scala 166:64:@38084.4]
  assign buffer_11_256 = {{8{_T_89943[5]}},_T_89943}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_257 = {{8{_T_89950[5]}},_T_89950}; // @[Modules.scala 112:22:@8.4]
  assign _T_90617 = $signed(buffer_11_256) + $signed(buffer_11_257); // @[Modules.scala 166:64:@38086.4]
  assign _T_90618 = _T_90617[13:0]; // @[Modules.scala 166:64:@38087.4]
  assign buffer_11_427 = $signed(_T_90618); // @[Modules.scala 166:64:@38088.4]
  assign _T_90620 = $signed(buffer_3_270) + $signed(buffer_6_273); // @[Modules.scala 166:64:@38090.4]
  assign _T_90621 = _T_90620[13:0]; // @[Modules.scala 166:64:@38091.4]
  assign buffer_11_428 = $signed(_T_90621); // @[Modules.scala 166:64:@38092.4]
  assign buffer_11_262 = {{9{_T_89985[4]}},_T_89985}; // @[Modules.scala 112:22:@8.4]
  assign _T_90626 = $signed(buffer_11_262) + $signed(buffer_1_268); // @[Modules.scala 166:64:@38098.4]
  assign _T_90627 = _T_90626[13:0]; // @[Modules.scala 166:64:@38099.4]
  assign buffer_11_430 = $signed(_T_90627); // @[Modules.scala 166:64:@38100.4]
  assign buffer_11_267 = {{8{_T_90020[5]}},_T_90020}; // @[Modules.scala 112:22:@8.4]
  assign _T_90632 = $signed(buffer_3_281) + $signed(buffer_11_267); // @[Modules.scala 166:64:@38106.4]
  assign _T_90633 = _T_90632[13:0]; // @[Modules.scala 166:64:@38107.4]
  assign buffer_11_432 = $signed(_T_90633); // @[Modules.scala 166:64:@38108.4]
  assign buffer_11_268 = {{8{_T_90027[5]}},_T_90027}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_269 = {{8{_T_90034[5]}},_T_90034}; // @[Modules.scala 112:22:@8.4]
  assign _T_90635 = $signed(buffer_11_268) + $signed(buffer_11_269); // @[Modules.scala 166:64:@38110.4]
  assign _T_90636 = _T_90635[13:0]; // @[Modules.scala 166:64:@38111.4]
  assign buffer_11_433 = $signed(_T_90636); // @[Modules.scala 166:64:@38112.4]
  assign buffer_11_270 = {{9{_T_90041[4]}},_T_90041}; // @[Modules.scala 112:22:@8.4]
  assign buffer_11_271 = {{9{_T_90048[4]}},_T_90048}; // @[Modules.scala 112:22:@8.4]
  assign _T_90638 = $signed(buffer_11_270) + $signed(buffer_11_271); // @[Modules.scala 166:64:@38114.4]
  assign _T_90639 = _T_90638[13:0]; // @[Modules.scala 166:64:@38115.4]
  assign buffer_11_434 = $signed(_T_90639); // @[Modules.scala 166:64:@38116.4]
  assign buffer_11_272 = {{9{_T_90055[4]}},_T_90055}; // @[Modules.scala 112:22:@8.4]
  assign _T_90641 = $signed(buffer_11_272) + $signed(buffer_2_284); // @[Modules.scala 166:64:@38118.4]
  assign _T_90642 = _T_90641[13:0]; // @[Modules.scala 166:64:@38119.4]
  assign buffer_11_435 = $signed(_T_90642); // @[Modules.scala 166:64:@38120.4]
  assign buffer_11_274 = {{8{_T_90069[5]}},_T_90069}; // @[Modules.scala 112:22:@8.4]
  assign _T_90644 = $signed(buffer_11_274) + $signed(buffer_1_280); // @[Modules.scala 166:64:@38122.4]
  assign _T_90645 = _T_90644[13:0]; // @[Modules.scala 166:64:@38123.4]
  assign buffer_11_436 = $signed(_T_90645); // @[Modules.scala 166:64:@38124.4]
  assign _T_90650 = $signed(buffer_3_292) + $signed(buffer_4_279); // @[Modules.scala 166:64:@38130.4]
  assign _T_90651 = _T_90650[13:0]; // @[Modules.scala 166:64:@38131.4]
  assign buffer_11_438 = $signed(_T_90651); // @[Modules.scala 166:64:@38132.4]
  assign buffer_11_281 = {{9{_T_90118[4]}},_T_90118}; // @[Modules.scala 112:22:@8.4]
  assign _T_90653 = $signed(buffer_3_294) + $signed(buffer_11_281); // @[Modules.scala 166:64:@38134.4]
  assign _T_90654 = _T_90653[13:0]; // @[Modules.scala 166:64:@38135.4]
  assign buffer_11_439 = $signed(_T_90654); // @[Modules.scala 166:64:@38136.4]
  assign _T_90659 = $signed(buffer_9_298) + $signed(buffer_2_296); // @[Modules.scala 166:64:@38142.4]
  assign _T_90660 = _T_90659[13:0]; // @[Modules.scala 166:64:@38143.4]
  assign buffer_11_441 = $signed(_T_90660); // @[Modules.scala 166:64:@38144.4]
  assign buffer_11_289 = {{8{_T_90174[5]}},_T_90174}; // @[Modules.scala 112:22:@8.4]
  assign _T_90665 = $signed(buffer_4_289) + $signed(buffer_11_289); // @[Modules.scala 166:64:@38150.4]
  assign _T_90666 = _T_90665[13:0]; // @[Modules.scala 166:64:@38151.4]
  assign buffer_11_443 = $signed(_T_90666); // @[Modules.scala 166:64:@38152.4]
  assign buffer_11_291 = {{8{_T_90188[5]}},_T_90188}; // @[Modules.scala 112:22:@8.4]
  assign _T_90668 = $signed(buffer_3_304) + $signed(buffer_11_291); // @[Modules.scala 166:64:@38154.4]
  assign _T_90669 = _T_90668[13:0]; // @[Modules.scala 166:64:@38155.4]
  assign buffer_11_444 = $signed(_T_90669); // @[Modules.scala 166:64:@38156.4]
  assign _T_90671 = $signed(buffer_9_307) + $signed(buffer_1_297); // @[Modules.scala 166:64:@38158.4]
  assign _T_90672 = _T_90671[13:0]; // @[Modules.scala 166:64:@38159.4]
  assign buffer_11_445 = $signed(_T_90672); // @[Modules.scala 166:64:@38160.4]
  assign buffer_11_295 = {{9{_T_90216[4]}},_T_90216}; // @[Modules.scala 112:22:@8.4]
  assign _T_90674 = $signed(buffer_9_309) + $signed(buffer_11_295); // @[Modules.scala 166:64:@38162.4]
  assign _T_90675 = _T_90674[13:0]; // @[Modules.scala 166:64:@38163.4]
  assign buffer_11_446 = $signed(_T_90675); // @[Modules.scala 166:64:@38164.4]
  assign _T_90677 = $signed(buffer_5_311) + $signed(buffer_2_309); // @[Modules.scala 166:64:@38166.4]
  assign _T_90678 = _T_90677[13:0]; // @[Modules.scala 166:64:@38167.4]
  assign buffer_11_447 = $signed(_T_90678); // @[Modules.scala 166:64:@38168.4]
  assign _T_90680 = $signed(buffer_11_299) + $signed(buffer_11_300); // @[Modules.scala 166:64:@38170.4]
  assign _T_90681 = _T_90680[13:0]; // @[Modules.scala 166:64:@38171.4]
  assign buffer_11_448 = $signed(_T_90681); // @[Modules.scala 166:64:@38172.4]
  assign _T_90683 = $signed(buffer_11_301) + $signed(buffer_11_302); // @[Modules.scala 166:64:@38174.4]
  assign _T_90684 = _T_90683[13:0]; // @[Modules.scala 166:64:@38175.4]
  assign buffer_11_449 = $signed(_T_90684); // @[Modules.scala 166:64:@38176.4]
  assign _T_90686 = $signed(buffer_11_303) + $signed(buffer_11_304); // @[Modules.scala 166:64:@38178.4]
  assign _T_90687 = _T_90686[13:0]; // @[Modules.scala 166:64:@38179.4]
  assign buffer_11_450 = $signed(_T_90687); // @[Modules.scala 166:64:@38180.4]
  assign _T_90689 = $signed(buffer_8_316) + $signed(buffer_7_316); // @[Modules.scala 166:64:@38182.4]
  assign _T_90690 = _T_90689[13:0]; // @[Modules.scala 166:64:@38183.4]
  assign buffer_11_451 = $signed(_T_90690); // @[Modules.scala 166:64:@38184.4]
  assign _T_90695 = $signed(buffer_11_309) + $signed(buffer_11_310); // @[Modules.scala 166:64:@38190.4]
  assign _T_90696 = _T_90695[13:0]; // @[Modules.scala 166:64:@38191.4]
  assign buffer_11_453 = $signed(_T_90696); // @[Modules.scala 166:64:@38192.4]
  assign _T_90698 = $signed(buffer_11_311) + $signed(buffer_11_312); // @[Modules.scala 166:64:@38194.4]
  assign _T_90699 = _T_90698[13:0]; // @[Modules.scala 166:64:@38195.4]
  assign buffer_11_454 = $signed(_T_90699); // @[Modules.scala 166:64:@38196.4]
  assign _T_90701 = $signed(buffer_11_313) + $signed(buffer_5_328); // @[Modules.scala 166:64:@38198.4]
  assign _T_90702 = _T_90701[13:0]; // @[Modules.scala 166:64:@38199.4]
  assign buffer_11_455 = $signed(_T_90702); // @[Modules.scala 166:64:@38200.4]
  assign _T_90704 = $signed(buffer_1_319) + $signed(buffer_11_316); // @[Modules.scala 166:64:@38202.4]
  assign _T_90705 = _T_90704[13:0]; // @[Modules.scala 166:64:@38203.4]
  assign buffer_11_456 = $signed(_T_90705); // @[Modules.scala 166:64:@38204.4]
  assign _T_90707 = $signed(buffer_11_317) + $signed(buffer_11_318); // @[Modules.scala 166:64:@38206.4]
  assign _T_90708 = _T_90707[13:0]; // @[Modules.scala 166:64:@38207.4]
  assign buffer_11_457 = $signed(_T_90708); // @[Modules.scala 166:64:@38208.4]
  assign _T_90710 = $signed(buffer_11_319) + $signed(buffer_11_320); // @[Modules.scala 166:64:@38210.4]
  assign _T_90711 = _T_90710[13:0]; // @[Modules.scala 166:64:@38211.4]
  assign buffer_11_458 = $signed(_T_90711); // @[Modules.scala 166:64:@38212.4]
  assign _T_90713 = $signed(buffer_11_321) + $signed(buffer_11_322); // @[Modules.scala 166:64:@38214.4]
  assign _T_90714 = _T_90713[13:0]; // @[Modules.scala 166:64:@38215.4]
  assign buffer_11_459 = $signed(_T_90714); // @[Modules.scala 166:64:@38216.4]
  assign _T_90716 = $signed(buffer_11_323) + $signed(buffer_11_324); // @[Modules.scala 166:64:@38218.4]
  assign _T_90717 = _T_90716[13:0]; // @[Modules.scala 166:64:@38219.4]
  assign buffer_11_460 = $signed(_T_90717); // @[Modules.scala 166:64:@38220.4]
  assign _T_90719 = $signed(buffer_11_325) + $signed(buffer_11_326); // @[Modules.scala 166:64:@38222.4]
  assign _T_90720 = _T_90719[13:0]; // @[Modules.scala 166:64:@38223.4]
  assign buffer_11_461 = $signed(_T_90720); // @[Modules.scala 166:64:@38224.4]
  assign _T_90722 = $signed(buffer_11_327) + $signed(buffer_11_328); // @[Modules.scala 166:64:@38226.4]
  assign _T_90723 = _T_90722[13:0]; // @[Modules.scala 166:64:@38227.4]
  assign buffer_11_462 = $signed(_T_90723); // @[Modules.scala 166:64:@38228.4]
  assign _T_90725 = $signed(buffer_11_329) + $signed(buffer_11_330); // @[Modules.scala 166:64:@38230.4]
  assign _T_90726 = _T_90725[13:0]; // @[Modules.scala 166:64:@38231.4]
  assign buffer_11_463 = $signed(_T_90726); // @[Modules.scala 166:64:@38232.4]
  assign _T_90728 = $signed(buffer_11_331) + $signed(buffer_11_332); // @[Modules.scala 166:64:@38234.4]
  assign _T_90729 = _T_90728[13:0]; // @[Modules.scala 166:64:@38235.4]
  assign buffer_11_464 = $signed(_T_90729); // @[Modules.scala 166:64:@38236.4]
  assign _T_90731 = $signed(buffer_10_343) + $signed(buffer_11_334); // @[Modules.scala 166:64:@38238.4]
  assign _T_90732 = _T_90731[13:0]; // @[Modules.scala 166:64:@38239.4]
  assign buffer_11_465 = $signed(_T_90732); // @[Modules.scala 166:64:@38240.4]
  assign _T_90734 = $signed(buffer_11_335) + $signed(buffer_11_336); // @[Modules.scala 166:64:@38242.4]
  assign _T_90735 = _T_90734[13:0]; // @[Modules.scala 166:64:@38243.4]
  assign buffer_11_466 = $signed(_T_90735); // @[Modules.scala 166:64:@38244.4]
  assign _T_90737 = $signed(buffer_11_337) + $signed(buffer_11_338); // @[Modules.scala 166:64:@38246.4]
  assign _T_90738 = _T_90737[13:0]; // @[Modules.scala 166:64:@38247.4]
  assign buffer_11_467 = $signed(_T_90738); // @[Modules.scala 166:64:@38248.4]
  assign _T_90740 = $signed(buffer_11_339) + $signed(buffer_11_340); // @[Modules.scala 166:64:@38250.4]
  assign _T_90741 = _T_90740[13:0]; // @[Modules.scala 166:64:@38251.4]
  assign buffer_11_468 = $signed(_T_90741); // @[Modules.scala 166:64:@38252.4]
  assign _T_90743 = $signed(buffer_11_341) + $signed(buffer_3_361); // @[Modules.scala 166:64:@38254.4]
  assign _T_90744 = _T_90743[13:0]; // @[Modules.scala 166:64:@38255.4]
  assign buffer_11_469 = $signed(_T_90744); // @[Modules.scala 166:64:@38256.4]
  assign _T_90746 = $signed(buffer_11_343) + $signed(buffer_11_344); // @[Modules.scala 166:64:@38258.4]
  assign _T_90747 = _T_90746[13:0]; // @[Modules.scala 166:64:@38259.4]
  assign buffer_11_470 = $signed(_T_90747); // @[Modules.scala 166:64:@38260.4]
  assign _T_90749 = $signed(buffer_11_345) + $signed(buffer_11_346); // @[Modules.scala 166:64:@38262.4]
  assign _T_90750 = _T_90749[13:0]; // @[Modules.scala 166:64:@38263.4]
  assign buffer_11_471 = $signed(_T_90750); // @[Modules.scala 166:64:@38264.4]
  assign _T_90752 = $signed(buffer_9_368) + $signed(buffer_11_348); // @[Modules.scala 166:64:@38266.4]
  assign _T_90753 = _T_90752[13:0]; // @[Modules.scala 166:64:@38267.4]
  assign buffer_11_472 = $signed(_T_90753); // @[Modules.scala 166:64:@38268.4]
  assign _T_90755 = $signed(buffer_11_349) + $signed(buffer_11_350); // @[Modules.scala 166:64:@38270.4]
  assign _T_90756 = _T_90755[13:0]; // @[Modules.scala 166:64:@38271.4]
  assign buffer_11_473 = $signed(_T_90756); // @[Modules.scala 166:64:@38272.4]
  assign _T_90758 = $signed(buffer_11_351) + $signed(buffer_11_352); // @[Modules.scala 166:64:@38274.4]
  assign _T_90759 = _T_90758[13:0]; // @[Modules.scala 166:64:@38275.4]
  assign buffer_11_474 = $signed(_T_90759); // @[Modules.scala 166:64:@38276.4]
  assign _T_90761 = $signed(buffer_11_353) + $signed(buffer_6_375); // @[Modules.scala 166:64:@38278.4]
  assign _T_90762 = _T_90761[13:0]; // @[Modules.scala 166:64:@38279.4]
  assign buffer_11_475 = $signed(_T_90762); // @[Modules.scala 166:64:@38280.4]
  assign _T_90764 = $signed(buffer_11_355) + $signed(buffer_11_356); // @[Modules.scala 166:64:@38282.4]
  assign _T_90765 = _T_90764[13:0]; // @[Modules.scala 166:64:@38283.4]
  assign buffer_11_476 = $signed(_T_90765); // @[Modules.scala 166:64:@38284.4]
  assign _T_90767 = $signed(buffer_11_357) + $signed(buffer_11_358); // @[Modules.scala 166:64:@38286.4]
  assign _T_90768 = _T_90767[13:0]; // @[Modules.scala 166:64:@38287.4]
  assign buffer_11_477 = $signed(_T_90768); // @[Modules.scala 166:64:@38288.4]
  assign _T_90770 = $signed(buffer_11_359) + $signed(buffer_0_366); // @[Modules.scala 166:64:@38290.4]
  assign _T_90771 = _T_90770[13:0]; // @[Modules.scala 166:64:@38291.4]
  assign buffer_11_478 = $signed(_T_90771); // @[Modules.scala 166:64:@38292.4]
  assign _T_90773 = $signed(buffer_11_361) + $signed(buffer_11_362); // @[Modules.scala 166:64:@38294.4]
  assign _T_90774 = _T_90773[13:0]; // @[Modules.scala 166:64:@38295.4]
  assign buffer_11_479 = $signed(_T_90774); // @[Modules.scala 166:64:@38296.4]
  assign _T_90776 = $signed(buffer_11_363) + $signed(buffer_11_364); // @[Modules.scala 166:64:@38298.4]
  assign _T_90777 = _T_90776[13:0]; // @[Modules.scala 166:64:@38299.4]
  assign buffer_11_480 = $signed(_T_90777); // @[Modules.scala 166:64:@38300.4]
  assign _T_90779 = $signed(buffer_11_365) + $signed(buffer_11_366); // @[Modules.scala 166:64:@38302.4]
  assign _T_90780 = _T_90779[13:0]; // @[Modules.scala 166:64:@38303.4]
  assign buffer_11_481 = $signed(_T_90780); // @[Modules.scala 166:64:@38304.4]
  assign _T_90782 = $signed(buffer_11_367) + $signed(buffer_3_390); // @[Modules.scala 166:64:@38306.4]
  assign _T_90783 = _T_90782[13:0]; // @[Modules.scala 166:64:@38307.4]
  assign buffer_11_482 = $signed(_T_90783); // @[Modules.scala 166:64:@38308.4]
  assign _T_90785 = $signed(buffer_11_369) + $signed(buffer_5_388); // @[Modules.scala 166:64:@38310.4]
  assign _T_90786 = _T_90785[13:0]; // @[Modules.scala 166:64:@38311.4]
  assign buffer_11_483 = $signed(_T_90786); // @[Modules.scala 166:64:@38312.4]
  assign _T_90788 = $signed(buffer_11_371) + $signed(buffer_7_385); // @[Modules.scala 166:64:@38314.4]
  assign _T_90789 = _T_90788[13:0]; // @[Modules.scala 166:64:@38315.4]
  assign buffer_11_484 = $signed(_T_90789); // @[Modules.scala 166:64:@38316.4]
  assign _T_90791 = $signed(buffer_11_373) + $signed(buffer_8_386); // @[Modules.scala 166:64:@38318.4]
  assign _T_90792 = _T_90791[13:0]; // @[Modules.scala 166:64:@38319.4]
  assign buffer_11_485 = $signed(_T_90792); // @[Modules.scala 166:64:@38320.4]
  assign _T_90794 = $signed(buffer_11_375) + $signed(buffer_1_384); // @[Modules.scala 166:64:@38322.4]
  assign _T_90795 = _T_90794[13:0]; // @[Modules.scala 166:64:@38323.4]
  assign buffer_11_486 = $signed(_T_90795); // @[Modules.scala 166:64:@38324.4]
  assign _T_90797 = $signed(buffer_11_377) + $signed(buffer_11_378); // @[Modules.scala 166:64:@38326.4]
  assign _T_90798 = _T_90797[13:0]; // @[Modules.scala 166:64:@38327.4]
  assign buffer_11_487 = $signed(_T_90798); // @[Modules.scala 166:64:@38328.4]
  assign _T_90800 = $signed(buffer_11_379) + $signed(buffer_11_380); // @[Modules.scala 166:64:@38330.4]
  assign _T_90801 = _T_90800[13:0]; // @[Modules.scala 166:64:@38331.4]
  assign buffer_11_488 = $signed(_T_90801); // @[Modules.scala 166:64:@38332.4]
  assign _T_90803 = $signed(buffer_11_381) + $signed(buffer_3_402); // @[Modules.scala 166:64:@38334.4]
  assign _T_90804 = _T_90803[13:0]; // @[Modules.scala 166:64:@38335.4]
  assign buffer_11_489 = $signed(_T_90804); // @[Modules.scala 166:64:@38336.4]
  assign _T_90806 = $signed(buffer_11_383) + $signed(buffer_11_384); // @[Modules.scala 166:64:@38338.4]
  assign _T_90807 = _T_90806[13:0]; // @[Modules.scala 166:64:@38339.4]
  assign buffer_11_490 = $signed(_T_90807); // @[Modules.scala 166:64:@38340.4]
  assign _T_90809 = $signed(buffer_11_385) + $signed(buffer_11_386); // @[Modules.scala 166:64:@38342.4]
  assign _T_90810 = _T_90809[13:0]; // @[Modules.scala 166:64:@38343.4]
  assign buffer_11_491 = $signed(_T_90810); // @[Modules.scala 166:64:@38344.4]
  assign _T_90812 = $signed(buffer_11_387) + $signed(buffer_3_409); // @[Modules.scala 166:64:@38346.4]
  assign _T_90813 = _T_90812[13:0]; // @[Modules.scala 166:64:@38347.4]
  assign buffer_11_492 = $signed(_T_90813); // @[Modules.scala 166:64:@38348.4]
  assign _T_90815 = $signed(buffer_11_389) + $signed(buffer_0_394); // @[Modules.scala 166:64:@38350.4]
  assign _T_90816 = _T_90815[13:0]; // @[Modules.scala 166:64:@38351.4]
  assign buffer_11_493 = $signed(_T_90816); // @[Modules.scala 166:64:@38352.4]
  assign _T_90818 = $signed(buffer_11_391) + $signed(buffer_11_392); // @[Modules.scala 166:64:@38354.4]
  assign _T_90819 = _T_90818[13:0]; // @[Modules.scala 166:64:@38355.4]
  assign buffer_11_494 = $signed(_T_90819); // @[Modules.scala 166:64:@38356.4]
  assign _T_90821 = $signed(buffer_11_393) + $signed(buffer_11_394); // @[Modules.scala 166:64:@38358.4]
  assign _T_90822 = _T_90821[13:0]; // @[Modules.scala 166:64:@38359.4]
  assign buffer_11_495 = $signed(_T_90822); // @[Modules.scala 166:64:@38360.4]
  assign _T_90824 = $signed(buffer_7_410) + $signed(buffer_11_396); // @[Modules.scala 166:64:@38362.4]
  assign _T_90825 = _T_90824[13:0]; // @[Modules.scala 166:64:@38363.4]
  assign buffer_11_496 = $signed(_T_90825); // @[Modules.scala 166:64:@38364.4]
  assign _T_90827 = $signed(buffer_11_397) + $signed(buffer_11_398); // @[Modules.scala 166:64:@38366.4]
  assign _T_90828 = _T_90827[13:0]; // @[Modules.scala 166:64:@38367.4]
  assign buffer_11_497 = $signed(_T_90828); // @[Modules.scala 166:64:@38368.4]
  assign _T_90830 = $signed(buffer_11_399) + $signed(buffer_11_400); // @[Modules.scala 166:64:@38370.4]
  assign _T_90831 = _T_90830[13:0]; // @[Modules.scala 166:64:@38371.4]
  assign buffer_11_498 = $signed(_T_90831); // @[Modules.scala 166:64:@38372.4]
  assign _T_90833 = $signed(buffer_11_401) + $signed(buffer_11_402); // @[Modules.scala 166:64:@38374.4]
  assign _T_90834 = _T_90833[13:0]; // @[Modules.scala 166:64:@38375.4]
  assign buffer_11_499 = $signed(_T_90834); // @[Modules.scala 166:64:@38376.4]
  assign _T_90836 = $signed(buffer_11_403) + $signed(buffer_8_417); // @[Modules.scala 166:64:@38378.4]
  assign _T_90837 = _T_90836[13:0]; // @[Modules.scala 166:64:@38379.4]
  assign buffer_11_500 = $signed(_T_90837); // @[Modules.scala 166:64:@38380.4]
  assign _T_90839 = $signed(buffer_11_405) + $signed(buffer_5_424); // @[Modules.scala 166:64:@38382.4]
  assign _T_90840 = _T_90839[13:0]; // @[Modules.scala 166:64:@38383.4]
  assign buffer_11_501 = $signed(_T_90840); // @[Modules.scala 166:64:@38384.4]
  assign _T_90842 = $signed(buffer_5_425) + $signed(buffer_11_408); // @[Modules.scala 166:64:@38386.4]
  assign _T_90843 = _T_90842[13:0]; // @[Modules.scala 166:64:@38387.4]
  assign buffer_11_502 = $signed(_T_90843); // @[Modules.scala 166:64:@38388.4]
  assign _T_90845 = $signed(buffer_11_409) + $signed(buffer_11_410); // @[Modules.scala 166:64:@38390.4]
  assign _T_90846 = _T_90845[13:0]; // @[Modules.scala 166:64:@38391.4]
  assign buffer_11_503 = $signed(_T_90846); // @[Modules.scala 166:64:@38392.4]
  assign _T_90848 = $signed(buffer_11_411) + $signed(buffer_11_412); // @[Modules.scala 166:64:@38394.4]
  assign _T_90849 = _T_90848[13:0]; // @[Modules.scala 166:64:@38395.4]
  assign buffer_11_504 = $signed(_T_90849); // @[Modules.scala 166:64:@38396.4]
  assign _T_90851 = $signed(buffer_11_413) + $signed(buffer_11_414); // @[Modules.scala 166:64:@38398.4]
  assign _T_90852 = _T_90851[13:0]; // @[Modules.scala 166:64:@38399.4]
  assign buffer_11_505 = $signed(_T_90852); // @[Modules.scala 166:64:@38400.4]
  assign _T_90854 = $signed(buffer_11_415) + $signed(buffer_11_416); // @[Modules.scala 166:64:@38402.4]
  assign _T_90855 = _T_90854[13:0]; // @[Modules.scala 166:64:@38403.4]
  assign buffer_11_506 = $signed(_T_90855); // @[Modules.scala 166:64:@38404.4]
  assign _T_90857 = $signed(buffer_11_417) + $signed(buffer_11_418); // @[Modules.scala 166:64:@38406.4]
  assign _T_90858 = _T_90857[13:0]; // @[Modules.scala 166:64:@38407.4]
  assign buffer_11_507 = $signed(_T_90858); // @[Modules.scala 166:64:@38408.4]
  assign _T_90860 = $signed(buffer_11_419) + $signed(buffer_11_420); // @[Modules.scala 166:64:@38410.4]
  assign _T_90861 = _T_90860[13:0]; // @[Modules.scala 166:64:@38411.4]
  assign buffer_11_508 = $signed(_T_90861); // @[Modules.scala 166:64:@38412.4]
  assign _T_90863 = $signed(buffer_11_421) + $signed(buffer_11_422); // @[Modules.scala 166:64:@38414.4]
  assign _T_90864 = _T_90863[13:0]; // @[Modules.scala 166:64:@38415.4]
  assign buffer_11_509 = $signed(_T_90864); // @[Modules.scala 166:64:@38416.4]
  assign _T_90866 = $signed(buffer_11_423) + $signed(buffer_11_424); // @[Modules.scala 166:64:@38418.4]
  assign _T_90867 = _T_90866[13:0]; // @[Modules.scala 166:64:@38419.4]
  assign buffer_11_510 = $signed(_T_90867); // @[Modules.scala 166:64:@38420.4]
  assign _T_90869 = $signed(buffer_11_425) + $signed(buffer_11_426); // @[Modules.scala 166:64:@38422.4]
  assign _T_90870 = _T_90869[13:0]; // @[Modules.scala 166:64:@38423.4]
  assign buffer_11_511 = $signed(_T_90870); // @[Modules.scala 166:64:@38424.4]
  assign _T_90872 = $signed(buffer_11_427) + $signed(buffer_11_428); // @[Modules.scala 166:64:@38426.4]
  assign _T_90873 = _T_90872[13:0]; // @[Modules.scala 166:64:@38427.4]
  assign buffer_11_512 = $signed(_T_90873); // @[Modules.scala 166:64:@38428.4]
  assign _T_90875 = $signed(buffer_3_450) + $signed(buffer_11_430); // @[Modules.scala 166:64:@38430.4]
  assign _T_90876 = _T_90875[13:0]; // @[Modules.scala 166:64:@38431.4]
  assign buffer_11_513 = $signed(_T_90876); // @[Modules.scala 166:64:@38432.4]
  assign _T_90878 = $signed(buffer_10_445) + $signed(buffer_11_432); // @[Modules.scala 166:64:@38434.4]
  assign _T_90879 = _T_90878[13:0]; // @[Modules.scala 166:64:@38435.4]
  assign buffer_11_514 = $signed(_T_90879); // @[Modules.scala 166:64:@38436.4]
  assign _T_90881 = $signed(buffer_11_433) + $signed(buffer_11_434); // @[Modules.scala 166:64:@38438.4]
  assign _T_90882 = _T_90881[13:0]; // @[Modules.scala 166:64:@38439.4]
  assign buffer_11_515 = $signed(_T_90882); // @[Modules.scala 166:64:@38440.4]
  assign _T_90884 = $signed(buffer_11_435) + $signed(buffer_11_436); // @[Modules.scala 166:64:@38442.4]
  assign _T_90885 = _T_90884[13:0]; // @[Modules.scala 166:64:@38443.4]
  assign buffer_11_516 = $signed(_T_90885); // @[Modules.scala 166:64:@38444.4]
  assign _T_90887 = $signed(buffer_3_459) + $signed(buffer_11_438); // @[Modules.scala 166:64:@38446.4]
  assign _T_90888 = _T_90887[13:0]; // @[Modules.scala 166:64:@38447.4]
  assign buffer_11_517 = $signed(_T_90888); // @[Modules.scala 166:64:@38448.4]
  assign _T_90890 = $signed(buffer_11_439) + $signed(buffer_9_462); // @[Modules.scala 166:64:@38450.4]
  assign _T_90891 = _T_90890[13:0]; // @[Modules.scala 166:64:@38451.4]
  assign buffer_11_518 = $signed(_T_90891); // @[Modules.scala 166:64:@38452.4]
  assign _T_90893 = $signed(buffer_11_441) + $signed(buffer_10_456); // @[Modules.scala 166:64:@38454.4]
  assign _T_90894 = _T_90893[13:0]; // @[Modules.scala 166:64:@38455.4]
  assign buffer_11_519 = $signed(_T_90894); // @[Modules.scala 166:64:@38456.4]
  assign _T_90896 = $signed(buffer_11_443) + $signed(buffer_11_444); // @[Modules.scala 166:64:@38458.4]
  assign _T_90897 = _T_90896[13:0]; // @[Modules.scala 166:64:@38459.4]
  assign buffer_11_520 = $signed(_T_90897); // @[Modules.scala 166:64:@38460.4]
  assign _T_90899 = $signed(buffer_11_445) + $signed(buffer_11_446); // @[Modules.scala 166:64:@38462.4]
  assign _T_90900 = _T_90899[13:0]; // @[Modules.scala 166:64:@38463.4]
  assign buffer_11_521 = $signed(_T_90900); // @[Modules.scala 166:64:@38464.4]
  assign buffer_11_298 = {{8{_T_56301[5]}},_T_56301}; // @[Modules.scala 112:22:@8.4]
  assign _T_90902 = $signed(buffer_11_447) + $signed(buffer_11_298); // @[Modules.scala 172:66:@38466.4]
  assign _T_90903 = _T_90902[13:0]; // @[Modules.scala 172:66:@38467.4]
  assign buffer_11_522 = $signed(_T_90903); // @[Modules.scala 172:66:@38468.4]
  assign _T_90905 = $signed(buffer_11_448) + $signed(buffer_11_449); // @[Modules.scala 166:64:@38470.4]
  assign _T_90906 = _T_90905[13:0]; // @[Modules.scala 166:64:@38471.4]
  assign buffer_11_523 = $signed(_T_90906); // @[Modules.scala 166:64:@38472.4]
  assign _T_90908 = $signed(buffer_11_450) + $signed(buffer_11_451); // @[Modules.scala 166:64:@38474.4]
  assign _T_90909 = _T_90908[13:0]; // @[Modules.scala 166:64:@38475.4]
  assign buffer_11_524 = $signed(_T_90909); // @[Modules.scala 166:64:@38476.4]
  assign _T_90911 = $signed(buffer_7_467) + $signed(buffer_11_453); // @[Modules.scala 166:64:@38478.4]
  assign _T_90912 = _T_90911[13:0]; // @[Modules.scala 166:64:@38479.4]
  assign buffer_11_525 = $signed(_T_90912); // @[Modules.scala 166:64:@38480.4]
  assign _T_90914 = $signed(buffer_11_454) + $signed(buffer_11_455); // @[Modules.scala 166:64:@38482.4]
  assign _T_90915 = _T_90914[13:0]; // @[Modules.scala 166:64:@38483.4]
  assign buffer_11_526 = $signed(_T_90915); // @[Modules.scala 166:64:@38484.4]
  assign _T_90917 = $signed(buffer_11_456) + $signed(buffer_11_457); // @[Modules.scala 166:64:@38486.4]
  assign _T_90918 = _T_90917[13:0]; // @[Modules.scala 166:64:@38487.4]
  assign buffer_11_527 = $signed(_T_90918); // @[Modules.scala 166:64:@38488.4]
  assign _T_90920 = $signed(buffer_11_458) + $signed(buffer_11_459); // @[Modules.scala 166:64:@38490.4]
  assign _T_90921 = _T_90920[13:0]; // @[Modules.scala 166:64:@38491.4]
  assign buffer_11_528 = $signed(_T_90921); // @[Modules.scala 166:64:@38492.4]
  assign _T_90923 = $signed(buffer_11_460) + $signed(buffer_11_461); // @[Modules.scala 166:64:@38494.4]
  assign _T_90924 = _T_90923[13:0]; // @[Modules.scala 166:64:@38495.4]
  assign buffer_11_529 = $signed(_T_90924); // @[Modules.scala 166:64:@38496.4]
  assign _T_90926 = $signed(buffer_11_462) + $signed(buffer_11_463); // @[Modules.scala 166:64:@38498.4]
  assign _T_90927 = _T_90926[13:0]; // @[Modules.scala 166:64:@38499.4]
  assign buffer_11_530 = $signed(_T_90927); // @[Modules.scala 166:64:@38500.4]
  assign _T_90929 = $signed(buffer_11_464) + $signed(buffer_11_465); // @[Modules.scala 166:64:@38502.4]
  assign _T_90930 = _T_90929[13:0]; // @[Modules.scala 166:64:@38503.4]
  assign buffer_11_531 = $signed(_T_90930); // @[Modules.scala 166:64:@38504.4]
  assign _T_90932 = $signed(buffer_11_466) + $signed(buffer_11_467); // @[Modules.scala 166:64:@38506.4]
  assign _T_90933 = _T_90932[13:0]; // @[Modules.scala 166:64:@38507.4]
  assign buffer_11_532 = $signed(_T_90933); // @[Modules.scala 166:64:@38508.4]
  assign _T_90935 = $signed(buffer_11_468) + $signed(buffer_11_469); // @[Modules.scala 166:64:@38510.4]
  assign _T_90936 = _T_90935[13:0]; // @[Modules.scala 166:64:@38511.4]
  assign buffer_11_533 = $signed(_T_90936); // @[Modules.scala 166:64:@38512.4]
  assign _T_90938 = $signed(buffer_11_470) + $signed(buffer_11_471); // @[Modules.scala 166:64:@38514.4]
  assign _T_90939 = _T_90938[13:0]; // @[Modules.scala 166:64:@38515.4]
  assign buffer_11_534 = $signed(_T_90939); // @[Modules.scala 166:64:@38516.4]
  assign _T_90941 = $signed(buffer_11_472) + $signed(buffer_11_473); // @[Modules.scala 166:64:@38518.4]
  assign _T_90942 = _T_90941[13:0]; // @[Modules.scala 166:64:@38519.4]
  assign buffer_11_535 = $signed(_T_90942); // @[Modules.scala 166:64:@38520.4]
  assign _T_90944 = $signed(buffer_11_474) + $signed(buffer_11_475); // @[Modules.scala 166:64:@38522.4]
  assign _T_90945 = _T_90944[13:0]; // @[Modules.scala 166:64:@38523.4]
  assign buffer_11_536 = $signed(_T_90945); // @[Modules.scala 166:64:@38524.4]
  assign _T_90947 = $signed(buffer_11_476) + $signed(buffer_11_477); // @[Modules.scala 166:64:@38526.4]
  assign _T_90948 = _T_90947[13:0]; // @[Modules.scala 166:64:@38527.4]
  assign buffer_11_537 = $signed(_T_90948); // @[Modules.scala 166:64:@38528.4]
  assign _T_90950 = $signed(buffer_11_478) + $signed(buffer_11_479); // @[Modules.scala 166:64:@38530.4]
  assign _T_90951 = _T_90950[13:0]; // @[Modules.scala 166:64:@38531.4]
  assign buffer_11_538 = $signed(_T_90951); // @[Modules.scala 166:64:@38532.4]
  assign _T_90953 = $signed(buffer_11_480) + $signed(buffer_11_481); // @[Modules.scala 166:64:@38534.4]
  assign _T_90954 = _T_90953[13:0]; // @[Modules.scala 166:64:@38535.4]
  assign buffer_11_539 = $signed(_T_90954); // @[Modules.scala 166:64:@38536.4]
  assign _T_90956 = $signed(buffer_11_482) + $signed(buffer_11_483); // @[Modules.scala 166:64:@38538.4]
  assign _T_90957 = _T_90956[13:0]; // @[Modules.scala 166:64:@38539.4]
  assign buffer_11_540 = $signed(_T_90957); // @[Modules.scala 166:64:@38540.4]
  assign _T_90959 = $signed(buffer_11_484) + $signed(buffer_11_485); // @[Modules.scala 166:64:@38542.4]
  assign _T_90960 = _T_90959[13:0]; // @[Modules.scala 166:64:@38543.4]
  assign buffer_11_541 = $signed(_T_90960); // @[Modules.scala 166:64:@38544.4]
  assign _T_90962 = $signed(buffer_11_486) + $signed(buffer_11_487); // @[Modules.scala 166:64:@38546.4]
  assign _T_90963 = _T_90962[13:0]; // @[Modules.scala 166:64:@38547.4]
  assign buffer_11_542 = $signed(_T_90963); // @[Modules.scala 166:64:@38548.4]
  assign _T_90965 = $signed(buffer_11_488) + $signed(buffer_11_489); // @[Modules.scala 166:64:@38550.4]
  assign _T_90966 = _T_90965[13:0]; // @[Modules.scala 166:64:@38551.4]
  assign buffer_11_543 = $signed(_T_90966); // @[Modules.scala 166:64:@38552.4]
  assign _T_90968 = $signed(buffer_11_490) + $signed(buffer_11_491); // @[Modules.scala 166:64:@38554.4]
  assign _T_90969 = _T_90968[13:0]; // @[Modules.scala 166:64:@38555.4]
  assign buffer_11_544 = $signed(_T_90969); // @[Modules.scala 166:64:@38556.4]
  assign _T_90971 = $signed(buffer_11_492) + $signed(buffer_11_493); // @[Modules.scala 166:64:@38558.4]
  assign _T_90972 = _T_90971[13:0]; // @[Modules.scala 166:64:@38559.4]
  assign buffer_11_545 = $signed(_T_90972); // @[Modules.scala 166:64:@38560.4]
  assign _T_90974 = $signed(buffer_11_494) + $signed(buffer_11_495); // @[Modules.scala 166:64:@38562.4]
  assign _T_90975 = _T_90974[13:0]; // @[Modules.scala 166:64:@38563.4]
  assign buffer_11_546 = $signed(_T_90975); // @[Modules.scala 166:64:@38564.4]
  assign _T_90977 = $signed(buffer_11_496) + $signed(buffer_11_497); // @[Modules.scala 166:64:@38566.4]
  assign _T_90978 = _T_90977[13:0]; // @[Modules.scala 166:64:@38567.4]
  assign buffer_11_547 = $signed(_T_90978); // @[Modules.scala 166:64:@38568.4]
  assign _T_90980 = $signed(buffer_11_498) + $signed(buffer_11_499); // @[Modules.scala 166:64:@38570.4]
  assign _T_90981 = _T_90980[13:0]; // @[Modules.scala 166:64:@38571.4]
  assign buffer_11_548 = $signed(_T_90981); // @[Modules.scala 166:64:@38572.4]
  assign _T_90983 = $signed(buffer_11_500) + $signed(buffer_11_501); // @[Modules.scala 166:64:@38574.4]
  assign _T_90984 = _T_90983[13:0]; // @[Modules.scala 166:64:@38575.4]
  assign buffer_11_549 = $signed(_T_90984); // @[Modules.scala 166:64:@38576.4]
  assign _T_90986 = $signed(buffer_11_502) + $signed(buffer_11_503); // @[Modules.scala 166:64:@38578.4]
  assign _T_90987 = _T_90986[13:0]; // @[Modules.scala 166:64:@38579.4]
  assign buffer_11_550 = $signed(_T_90987); // @[Modules.scala 166:64:@38580.4]
  assign _T_90989 = $signed(buffer_11_504) + $signed(buffer_11_505); // @[Modules.scala 166:64:@38582.4]
  assign _T_90990 = _T_90989[13:0]; // @[Modules.scala 166:64:@38583.4]
  assign buffer_11_551 = $signed(_T_90990); // @[Modules.scala 166:64:@38584.4]
  assign _T_90992 = $signed(buffer_11_506) + $signed(buffer_11_507); // @[Modules.scala 166:64:@38586.4]
  assign _T_90993 = _T_90992[13:0]; // @[Modules.scala 166:64:@38587.4]
  assign buffer_11_552 = $signed(_T_90993); // @[Modules.scala 166:64:@38588.4]
  assign _T_90995 = $signed(buffer_11_508) + $signed(buffer_11_509); // @[Modules.scala 166:64:@38590.4]
  assign _T_90996 = _T_90995[13:0]; // @[Modules.scala 166:64:@38591.4]
  assign buffer_11_553 = $signed(_T_90996); // @[Modules.scala 166:64:@38592.4]
  assign _T_90998 = $signed(buffer_11_510) + $signed(buffer_11_511); // @[Modules.scala 166:64:@38594.4]
  assign _T_90999 = _T_90998[13:0]; // @[Modules.scala 166:64:@38595.4]
  assign buffer_11_554 = $signed(_T_90999); // @[Modules.scala 166:64:@38596.4]
  assign _T_91001 = $signed(buffer_11_512) + $signed(buffer_11_513); // @[Modules.scala 166:64:@38598.4]
  assign _T_91002 = _T_91001[13:0]; // @[Modules.scala 166:64:@38599.4]
  assign buffer_11_555 = $signed(_T_91002); // @[Modules.scala 166:64:@38600.4]
  assign _T_91004 = $signed(buffer_11_514) + $signed(buffer_11_515); // @[Modules.scala 166:64:@38602.4]
  assign _T_91005 = _T_91004[13:0]; // @[Modules.scala 166:64:@38603.4]
  assign buffer_11_556 = $signed(_T_91005); // @[Modules.scala 166:64:@38604.4]
  assign _T_91007 = $signed(buffer_11_516) + $signed(buffer_11_517); // @[Modules.scala 166:64:@38606.4]
  assign _T_91008 = _T_91007[13:0]; // @[Modules.scala 166:64:@38607.4]
  assign buffer_11_557 = $signed(_T_91008); // @[Modules.scala 166:64:@38608.4]
  assign _T_91010 = $signed(buffer_11_518) + $signed(buffer_11_519); // @[Modules.scala 166:64:@38610.4]
  assign _T_91011 = _T_91010[13:0]; // @[Modules.scala 166:64:@38611.4]
  assign buffer_11_558 = $signed(_T_91011); // @[Modules.scala 166:64:@38612.4]
  assign _T_91013 = $signed(buffer_11_520) + $signed(buffer_11_521); // @[Modules.scala 166:64:@38614.4]
  assign _T_91014 = _T_91013[13:0]; // @[Modules.scala 166:64:@38615.4]
  assign buffer_11_559 = $signed(_T_91014); // @[Modules.scala 166:64:@38616.4]
  assign _T_91016 = $signed(buffer_11_523) + $signed(buffer_11_524); // @[Modules.scala 166:64:@38618.4]
  assign _T_91017 = _T_91016[13:0]; // @[Modules.scala 166:64:@38619.4]
  assign buffer_11_560 = $signed(_T_91017); // @[Modules.scala 166:64:@38620.4]
  assign _T_91019 = $signed(buffer_11_525) + $signed(buffer_11_526); // @[Modules.scala 166:64:@38622.4]
  assign _T_91020 = _T_91019[13:0]; // @[Modules.scala 166:64:@38623.4]
  assign buffer_11_561 = $signed(_T_91020); // @[Modules.scala 166:64:@38624.4]
  assign _T_91022 = $signed(buffer_11_527) + $signed(buffer_11_528); // @[Modules.scala 166:64:@38626.4]
  assign _T_91023 = _T_91022[13:0]; // @[Modules.scala 166:64:@38627.4]
  assign buffer_11_562 = $signed(_T_91023); // @[Modules.scala 166:64:@38628.4]
  assign _T_91025 = $signed(buffer_11_529) + $signed(buffer_11_530); // @[Modules.scala 166:64:@38630.4]
  assign _T_91026 = _T_91025[13:0]; // @[Modules.scala 166:64:@38631.4]
  assign buffer_11_563 = $signed(_T_91026); // @[Modules.scala 166:64:@38632.4]
  assign _T_91028 = $signed(buffer_11_531) + $signed(buffer_11_532); // @[Modules.scala 166:64:@38634.4]
  assign _T_91029 = _T_91028[13:0]; // @[Modules.scala 166:64:@38635.4]
  assign buffer_11_564 = $signed(_T_91029); // @[Modules.scala 166:64:@38636.4]
  assign _T_91031 = $signed(buffer_11_533) + $signed(buffer_11_534); // @[Modules.scala 166:64:@38638.4]
  assign _T_91032 = _T_91031[13:0]; // @[Modules.scala 166:64:@38639.4]
  assign buffer_11_565 = $signed(_T_91032); // @[Modules.scala 166:64:@38640.4]
  assign _T_91034 = $signed(buffer_11_535) + $signed(buffer_11_536); // @[Modules.scala 166:64:@38642.4]
  assign _T_91035 = _T_91034[13:0]; // @[Modules.scala 166:64:@38643.4]
  assign buffer_11_566 = $signed(_T_91035); // @[Modules.scala 166:64:@38644.4]
  assign _T_91037 = $signed(buffer_11_537) + $signed(buffer_11_538); // @[Modules.scala 166:64:@38646.4]
  assign _T_91038 = _T_91037[13:0]; // @[Modules.scala 166:64:@38647.4]
  assign buffer_11_567 = $signed(_T_91038); // @[Modules.scala 166:64:@38648.4]
  assign _T_91040 = $signed(buffer_11_539) + $signed(buffer_11_540); // @[Modules.scala 166:64:@38650.4]
  assign _T_91041 = _T_91040[13:0]; // @[Modules.scala 166:64:@38651.4]
  assign buffer_11_568 = $signed(_T_91041); // @[Modules.scala 166:64:@38652.4]
  assign _T_91043 = $signed(buffer_11_541) + $signed(buffer_11_542); // @[Modules.scala 166:64:@38654.4]
  assign _T_91044 = _T_91043[13:0]; // @[Modules.scala 166:64:@38655.4]
  assign buffer_11_569 = $signed(_T_91044); // @[Modules.scala 166:64:@38656.4]
  assign _T_91046 = $signed(buffer_11_543) + $signed(buffer_11_544); // @[Modules.scala 166:64:@38658.4]
  assign _T_91047 = _T_91046[13:0]; // @[Modules.scala 166:64:@38659.4]
  assign buffer_11_570 = $signed(_T_91047); // @[Modules.scala 166:64:@38660.4]
  assign _T_91049 = $signed(buffer_11_545) + $signed(buffer_11_546); // @[Modules.scala 166:64:@38662.4]
  assign _T_91050 = _T_91049[13:0]; // @[Modules.scala 166:64:@38663.4]
  assign buffer_11_571 = $signed(_T_91050); // @[Modules.scala 166:64:@38664.4]
  assign _T_91052 = $signed(buffer_11_547) + $signed(buffer_11_548); // @[Modules.scala 166:64:@38666.4]
  assign _T_91053 = _T_91052[13:0]; // @[Modules.scala 166:64:@38667.4]
  assign buffer_11_572 = $signed(_T_91053); // @[Modules.scala 166:64:@38668.4]
  assign _T_91055 = $signed(buffer_11_549) + $signed(buffer_11_550); // @[Modules.scala 166:64:@38670.4]
  assign _T_91056 = _T_91055[13:0]; // @[Modules.scala 166:64:@38671.4]
  assign buffer_11_573 = $signed(_T_91056); // @[Modules.scala 166:64:@38672.4]
  assign _T_91058 = $signed(buffer_11_551) + $signed(buffer_11_552); // @[Modules.scala 166:64:@38674.4]
  assign _T_91059 = _T_91058[13:0]; // @[Modules.scala 166:64:@38675.4]
  assign buffer_11_574 = $signed(_T_91059); // @[Modules.scala 166:64:@38676.4]
  assign _T_91061 = $signed(buffer_11_553) + $signed(buffer_11_554); // @[Modules.scala 166:64:@38678.4]
  assign _T_91062 = _T_91061[13:0]; // @[Modules.scala 166:64:@38679.4]
  assign buffer_11_575 = $signed(_T_91062); // @[Modules.scala 166:64:@38680.4]
  assign _T_91064 = $signed(buffer_11_555) + $signed(buffer_11_556); // @[Modules.scala 166:64:@38682.4]
  assign _T_91065 = _T_91064[13:0]; // @[Modules.scala 166:64:@38683.4]
  assign buffer_11_576 = $signed(_T_91065); // @[Modules.scala 166:64:@38684.4]
  assign _T_91067 = $signed(buffer_11_557) + $signed(buffer_11_558); // @[Modules.scala 166:64:@38686.4]
  assign _T_91068 = _T_91067[13:0]; // @[Modules.scala 166:64:@38687.4]
  assign buffer_11_577 = $signed(_T_91068); // @[Modules.scala 166:64:@38688.4]
  assign _T_91070 = $signed(buffer_11_559) + $signed(buffer_11_522); // @[Modules.scala 172:66:@38690.4]
  assign _T_91071 = _T_91070[13:0]; // @[Modules.scala 172:66:@38691.4]
  assign buffer_11_578 = $signed(_T_91071); // @[Modules.scala 172:66:@38692.4]
  assign _T_91073 = $signed(buffer_11_560) + $signed(buffer_11_561); // @[Modules.scala 166:64:@38694.4]
  assign _T_91074 = _T_91073[13:0]; // @[Modules.scala 166:64:@38695.4]
  assign buffer_11_579 = $signed(_T_91074); // @[Modules.scala 166:64:@38696.4]
  assign _T_91076 = $signed(buffer_11_562) + $signed(buffer_11_563); // @[Modules.scala 166:64:@38698.4]
  assign _T_91077 = _T_91076[13:0]; // @[Modules.scala 166:64:@38699.4]
  assign buffer_11_580 = $signed(_T_91077); // @[Modules.scala 166:64:@38700.4]
  assign _T_91079 = $signed(buffer_11_564) + $signed(buffer_11_565); // @[Modules.scala 166:64:@38702.4]
  assign _T_91080 = _T_91079[13:0]; // @[Modules.scala 166:64:@38703.4]
  assign buffer_11_581 = $signed(_T_91080); // @[Modules.scala 166:64:@38704.4]
  assign _T_91082 = $signed(buffer_11_566) + $signed(buffer_11_567); // @[Modules.scala 166:64:@38706.4]
  assign _T_91083 = _T_91082[13:0]; // @[Modules.scala 166:64:@38707.4]
  assign buffer_11_582 = $signed(_T_91083); // @[Modules.scala 166:64:@38708.4]
  assign _T_91085 = $signed(buffer_11_568) + $signed(buffer_11_569); // @[Modules.scala 166:64:@38710.4]
  assign _T_91086 = _T_91085[13:0]; // @[Modules.scala 166:64:@38711.4]
  assign buffer_11_583 = $signed(_T_91086); // @[Modules.scala 166:64:@38712.4]
  assign _T_91088 = $signed(buffer_11_570) + $signed(buffer_11_571); // @[Modules.scala 166:64:@38714.4]
  assign _T_91089 = _T_91088[13:0]; // @[Modules.scala 166:64:@38715.4]
  assign buffer_11_584 = $signed(_T_91089); // @[Modules.scala 166:64:@38716.4]
  assign _T_91091 = $signed(buffer_11_572) + $signed(buffer_11_573); // @[Modules.scala 166:64:@38718.4]
  assign _T_91092 = _T_91091[13:0]; // @[Modules.scala 166:64:@38719.4]
  assign buffer_11_585 = $signed(_T_91092); // @[Modules.scala 166:64:@38720.4]
  assign _T_91094 = $signed(buffer_11_574) + $signed(buffer_11_575); // @[Modules.scala 166:64:@38722.4]
  assign _T_91095 = _T_91094[13:0]; // @[Modules.scala 166:64:@38723.4]
  assign buffer_11_586 = $signed(_T_91095); // @[Modules.scala 166:64:@38724.4]
  assign _T_91097 = $signed(buffer_11_576) + $signed(buffer_11_577); // @[Modules.scala 166:64:@38726.4]
  assign _T_91098 = _T_91097[13:0]; // @[Modules.scala 166:64:@38727.4]
  assign buffer_11_587 = $signed(_T_91098); // @[Modules.scala 166:64:@38728.4]
  assign _T_91100 = $signed(buffer_11_579) + $signed(buffer_11_580); // @[Modules.scala 166:64:@38730.4]
  assign _T_91101 = _T_91100[13:0]; // @[Modules.scala 166:64:@38731.4]
  assign buffer_11_588 = $signed(_T_91101); // @[Modules.scala 166:64:@38732.4]
  assign _T_91103 = $signed(buffer_11_581) + $signed(buffer_11_582); // @[Modules.scala 166:64:@38734.4]
  assign _T_91104 = _T_91103[13:0]; // @[Modules.scala 166:64:@38735.4]
  assign buffer_11_589 = $signed(_T_91104); // @[Modules.scala 166:64:@38736.4]
  assign _T_91106 = $signed(buffer_11_583) + $signed(buffer_11_584); // @[Modules.scala 166:64:@38738.4]
  assign _T_91107 = _T_91106[13:0]; // @[Modules.scala 166:64:@38739.4]
  assign buffer_11_590 = $signed(_T_91107); // @[Modules.scala 166:64:@38740.4]
  assign _T_91109 = $signed(buffer_11_585) + $signed(buffer_11_586); // @[Modules.scala 166:64:@38742.4]
  assign _T_91110 = _T_91109[13:0]; // @[Modules.scala 166:64:@38743.4]
  assign buffer_11_591 = $signed(_T_91110); // @[Modules.scala 166:64:@38744.4]
  assign _T_91112 = $signed(buffer_11_587) + $signed(buffer_11_578); // @[Modules.scala 172:66:@38746.4]
  assign _T_91113 = _T_91112[13:0]; // @[Modules.scala 172:66:@38747.4]
  assign buffer_11_592 = $signed(_T_91113); // @[Modules.scala 172:66:@38748.4]
  assign _T_91115 = $signed(buffer_11_588) + $signed(buffer_11_589); // @[Modules.scala 166:64:@38750.4]
  assign _T_91116 = _T_91115[13:0]; // @[Modules.scala 166:64:@38751.4]
  assign buffer_11_593 = $signed(_T_91116); // @[Modules.scala 166:64:@38752.4]
  assign _T_91118 = $signed(buffer_11_590) + $signed(buffer_11_591); // @[Modules.scala 166:64:@38754.4]
  assign _T_91119 = _T_91118[13:0]; // @[Modules.scala 166:64:@38755.4]
  assign buffer_11_594 = $signed(_T_91119); // @[Modules.scala 166:64:@38756.4]
  assign _T_91121 = $signed(buffer_11_593) + $signed(buffer_11_594); // @[Modules.scala 160:64:@38758.4]
  assign _T_91122 = _T_91121[13:0]; // @[Modules.scala 160:64:@38759.4]
  assign buffer_11_595 = $signed(_T_91122); // @[Modules.scala 160:64:@38760.4]
  assign _T_91124 = $signed(buffer_11_595) + $signed(buffer_11_592); // @[Modules.scala 172:66:@38762.4]
  assign _T_91125 = _T_91124[13:0]; // @[Modules.scala 172:66:@38763.4]
  assign buffer_11_596 = $signed(_T_91125); // @[Modules.scala 172:66:@38764.4]
  assign _T_91128 = $signed(4'sh1) * $signed(io_in_10); // @[Modules.scala 143:74:@38953.4]
  assign _GEN_832 = {{1{_T_60248[4]}},_T_60248}; // @[Modules.scala 143:103:@38955.4]
  assign _T_91131 = $signed(_T_91128) + $signed(_GEN_832); // @[Modules.scala 143:103:@38955.4]
  assign _T_91132 = _T_91131[5:0]; // @[Modules.scala 143:103:@38956.4]
  assign _T_91133 = $signed(_T_91132); // @[Modules.scala 143:103:@38957.4]
  assign _GEN_833 = {{1{_T_60250[4]}},_T_60250}; // @[Modules.scala 143:103:@38961.4]
  assign _T_91138 = $signed(_GEN_833) + $signed(_T_54206); // @[Modules.scala 143:103:@38961.4]
  assign _T_91139 = _T_91138[5:0]; // @[Modules.scala 143:103:@38962.4]
  assign _T_91140 = $signed(_T_91139); // @[Modules.scala 143:103:@38963.4]
  assign _T_91166 = $signed(_T_54227) + $signed(_T_54234); // @[Modules.scala 143:103:@38985.4]
  assign _T_91167 = _T_91166[5:0]; // @[Modules.scala 143:103:@38986.4]
  assign _T_91168 = $signed(_T_91167); // @[Modules.scala 143:103:@38987.4]
  assign _GEN_834 = {{1{_T_63408[4]}},_T_63408}; // @[Modules.scala 143:103:@39009.4]
  assign _T_91194 = $signed(_T_54262) + $signed(_GEN_834); // @[Modules.scala 143:103:@39009.4]
  assign _T_91195 = _T_91194[5:0]; // @[Modules.scala 143:103:@39010.4]
  assign _T_91196 = $signed(_T_91195); // @[Modules.scala 143:103:@39011.4]
  assign _T_91207 = $signed(4'sh1) * $signed(io_in_56); // @[Modules.scala 144:80:@39020.4]
  assign _T_91208 = $signed(_T_54276) + $signed(_T_91207); // @[Modules.scala 143:103:@39021.4]
  assign _T_91209 = _T_91208[5:0]; // @[Modules.scala 143:103:@39022.4]
  assign _T_91210 = $signed(_T_91209); // @[Modules.scala 143:103:@39023.4]
  assign _T_91222 = $signed(_T_60334) + $signed(_T_57302); // @[Modules.scala 143:103:@39033.4]
  assign _T_91223 = _T_91222[4:0]; // @[Modules.scala 143:103:@39034.4]
  assign _T_91224 = $signed(_T_91223); // @[Modules.scala 143:103:@39035.4]
  assign _GEN_835 = {{1{_T_57304[4]}},_T_57304}; // @[Modules.scala 143:103:@39039.4]
  assign _T_91229 = $signed(_GEN_835) + $signed(_T_54299); // @[Modules.scala 143:103:@39039.4]
  assign _T_91230 = _T_91229[5:0]; // @[Modules.scala 143:103:@39040.4]
  assign _T_91231 = $signed(_T_91230); // @[Modules.scala 143:103:@39041.4]
  assign _GEN_836 = {{1{_T_57316[4]}},_T_57316}; // @[Modules.scala 143:103:@39045.4]
  assign _T_91236 = $signed(_T_54304) + $signed(_GEN_836); // @[Modules.scala 143:103:@39045.4]
  assign _T_91237 = _T_91236[5:0]; // @[Modules.scala 143:103:@39046.4]
  assign _T_91238 = $signed(_T_91237); // @[Modules.scala 143:103:@39047.4]
  assign _GEN_837 = {{1{_T_57318[4]}},_T_57318}; // @[Modules.scala 143:103:@39051.4]
  assign _T_91243 = $signed(_GEN_837) + $signed(_T_54320); // @[Modules.scala 143:103:@39051.4]
  assign _T_91244 = _T_91243[5:0]; // @[Modules.scala 143:103:@39052.4]
  assign _T_91245 = $signed(_T_91244); // @[Modules.scala 143:103:@39053.4]
  assign _GEN_838 = {{1{_T_66603[4]}},_T_66603}; // @[Modules.scala 143:103:@39057.4]
  assign _T_91250 = $signed(_GEN_838) + $signed(_T_54341); // @[Modules.scala 143:103:@39057.4]
  assign _T_91251 = _T_91250[5:0]; // @[Modules.scala 143:103:@39058.4]
  assign _T_91252 = $signed(_T_91251); // @[Modules.scala 143:103:@39059.4]
  assign _T_91320 = $signed(_T_57409) + $signed(_T_57421); // @[Modules.scala 143:103:@39117.4]
  assign _T_91321 = _T_91320[4:0]; // @[Modules.scala 143:103:@39118.4]
  assign _T_91322 = $signed(_T_91321); // @[Modules.scala 143:103:@39119.4]
  assign _T_91362 = $signed(_T_57456) + $signed(_GEN_5); // @[Modules.scala 143:103:@39153.4]
  assign _T_91363 = _T_91362[5:0]; // @[Modules.scala 143:103:@39154.4]
  assign _T_91364 = $signed(_T_91363); // @[Modules.scala 143:103:@39155.4]
  assign _GEN_843 = {{1{_T_60502[4]}},_T_60502}; // @[Modules.scala 143:103:@39165.4]
  assign _T_91376 = $signed(_GEN_843) + $signed(_T_69749); // @[Modules.scala 143:103:@39165.4]
  assign _T_91377 = _T_91376[5:0]; // @[Modules.scala 143:103:@39166.4]
  assign _T_91378 = $signed(_T_91377); // @[Modules.scala 143:103:@39167.4]
  assign _T_91383 = $signed(_T_57486) + $signed(_T_66750); // @[Modules.scala 143:103:@39171.4]
  assign _T_91384 = _T_91383[4:0]; // @[Modules.scala 143:103:@39172.4]
  assign _T_91385 = $signed(_T_91384); // @[Modules.scala 143:103:@39173.4]
  assign _T_91397 = $signed(_GEN_639) + $signed(_T_54500); // @[Modules.scala 143:103:@39183.4]
  assign _T_91398 = _T_91397[5:0]; // @[Modules.scala 143:103:@39184.4]
  assign _T_91399 = $signed(_T_91398); // @[Modules.scala 143:103:@39185.4]
  assign _T_91418 = $signed(_T_54516) + $signed(_T_60549); // @[Modules.scala 143:103:@39201.4]
  assign _T_91419 = _T_91418[5:0]; // @[Modules.scala 143:103:@39202.4]
  assign _T_91420 = $signed(_T_91419); // @[Modules.scala 143:103:@39203.4]
  assign _T_91432 = $signed(_T_57533) + $signed(_T_57542); // @[Modules.scala 143:103:@39213.4]
  assign _T_91433 = _T_91432[5:0]; // @[Modules.scala 143:103:@39214.4]
  assign _T_91434 = $signed(_T_91433); // @[Modules.scala 143:103:@39215.4]
  assign _T_91439 = $signed(_T_60577) + $signed(_T_60586); // @[Modules.scala 143:103:@39219.4]
  assign _T_91440 = _T_91439[4:0]; // @[Modules.scala 143:103:@39220.4]
  assign _T_91441 = $signed(_T_91440); // @[Modules.scala 143:103:@39221.4]
  assign _GEN_845 = {{1{_T_57563[4]}},_T_57563}; // @[Modules.scala 143:103:@39225.4]
  assign _T_91446 = $signed(_GEN_845) + $signed(_T_69833); // @[Modules.scala 143:103:@39225.4]
  assign _T_91447 = _T_91446[5:0]; // @[Modules.scala 143:103:@39226.4]
  assign _T_91448 = $signed(_T_91447); // @[Modules.scala 143:103:@39227.4]
  assign _T_91453 = $signed(_T_60605) + $signed(_T_63723); // @[Modules.scala 143:103:@39231.4]
  assign _T_91454 = _T_91453[5:0]; // @[Modules.scala 143:103:@39232.4]
  assign _T_91455 = $signed(_T_91454); // @[Modules.scala 143:103:@39233.4]
  assign _T_91481 = $signed(_T_54577) + $signed(_T_60628); // @[Modules.scala 143:103:@39255.4]
  assign _T_91482 = _T_91481[5:0]; // @[Modules.scala 143:103:@39256.4]
  assign _T_91483 = $signed(_T_91482); // @[Modules.scala 143:103:@39257.4]
  assign _T_91488 = $signed(_GEN_13) + $signed(_T_54591); // @[Modules.scala 143:103:@39261.4]
  assign _T_91489 = _T_91488[5:0]; // @[Modules.scala 143:103:@39262.4]
  assign _T_91490 = $signed(_T_91489); // @[Modules.scala 143:103:@39263.4]
  assign _T_91502 = $signed(_GEN_373) + $signed(_T_73021); // @[Modules.scala 143:103:@39273.4]
  assign _T_91503 = _T_91502[5:0]; // @[Modules.scala 143:103:@39274.4]
  assign _T_91504 = $signed(_T_91503); // @[Modules.scala 143:103:@39275.4]
  assign _T_91530 = $signed(_T_73049) + $signed(_T_63814); // @[Modules.scala 143:103:@39297.4]
  assign _T_91531 = _T_91530[5:0]; // @[Modules.scala 143:103:@39298.4]
  assign _T_91532 = $signed(_T_91531); // @[Modules.scala 143:103:@39299.4]
  assign _T_91551 = $signed(_T_54654) + $signed(_T_57675); // @[Modules.scala 143:103:@39315.4]
  assign _T_91552 = _T_91551[5:0]; // @[Modules.scala 143:103:@39316.4]
  assign _T_91553 = $signed(_T_91552); // @[Modules.scala 143:103:@39317.4]
  assign _T_91558 = $signed(_T_54661) + $signed(_GEN_646); // @[Modules.scala 143:103:@39321.4]
  assign _T_91559 = _T_91558[5:0]; // @[Modules.scala 143:103:@39322.4]
  assign _T_91560 = $signed(_T_91559); // @[Modules.scala 143:103:@39323.4]
  assign _GEN_850 = {{1{_T_60717[4]}},_T_60717}; // @[Modules.scala 143:103:@39327.4]
  assign _T_91565 = $signed(_GEN_850) + $signed(_T_54670); // @[Modules.scala 143:103:@39327.4]
  assign _T_91566 = _T_91565[5:0]; // @[Modules.scala 143:103:@39328.4]
  assign _T_91567 = $signed(_T_91566); // @[Modules.scala 143:103:@39329.4]
  assign _T_91600 = $signed(_T_57738) + $signed(_T_63898); // @[Modules.scala 143:103:@39357.4]
  assign _T_91601 = _T_91600[5:0]; // @[Modules.scala 143:103:@39358.4]
  assign _T_91602 = $signed(_T_91601); // @[Modules.scala 143:103:@39359.4]
  assign _T_91621 = $signed(_T_57764) + $signed(_GEN_379); // @[Modules.scala 143:103:@39375.4]
  assign _T_91622 = _T_91621[5:0]; // @[Modules.scala 143:103:@39376.4]
  assign _T_91623 = $signed(_T_91622); // @[Modules.scala 143:103:@39377.4]
  assign _T_91642 = $signed(_T_57787) + $signed(_T_60831); // @[Modules.scala 143:103:@39393.4]
  assign _T_91643 = _T_91642[4:0]; // @[Modules.scala 143:103:@39394.4]
  assign _T_91644 = $signed(_T_91643); // @[Modules.scala 143:103:@39395.4]
  assign _GEN_854 = {{1{_T_57794[4]}},_T_57794}; // @[Modules.scala 143:103:@39399.4]
  assign _T_91649 = $signed(_GEN_854) + $signed(_T_57799); // @[Modules.scala 143:103:@39399.4]
  assign _T_91650 = _T_91649[5:0]; // @[Modules.scala 143:103:@39400.4]
  assign _T_91651 = $signed(_T_91650); // @[Modules.scala 143:103:@39401.4]
  assign _GEN_855 = {{1{_T_60850[4]}},_T_60850}; // @[Modules.scala 143:103:@39405.4]
  assign _T_91656 = $signed(_T_54766) + $signed(_GEN_855); // @[Modules.scala 143:103:@39405.4]
  assign _T_91657 = _T_91656[5:0]; // @[Modules.scala 143:103:@39406.4]
  assign _T_91658 = $signed(_T_91657); // @[Modules.scala 143:103:@39407.4]
  assign _T_91663 = $signed(_T_57815) + $signed(_GEN_592); // @[Modules.scala 143:103:@39411.4]
  assign _T_91664 = _T_91663[5:0]; // @[Modules.scala 143:103:@39412.4]
  assign _T_91665 = $signed(_T_91664); // @[Modules.scala 143:103:@39413.4]
  assign _T_91698 = $signed(_GEN_593) + $signed(_T_54822); // @[Modules.scala 143:103:@39441.4]
  assign _T_91699 = _T_91698[5:0]; // @[Modules.scala 143:103:@39442.4]
  assign _T_91700 = $signed(_T_91699); // @[Modules.scala 143:103:@39443.4]
  assign _GEN_858 = {{1{_T_54864[4]}},_T_54864}; // @[Modules.scala 143:103:@39483.4]
  assign _T_91747 = $signed(_GEN_858) + $signed(_T_57904); // @[Modules.scala 143:103:@39483.4]
  assign _T_91748 = _T_91747[5:0]; // @[Modules.scala 143:103:@39484.4]
  assign _T_91749 = $signed(_T_91748); // @[Modules.scala 143:103:@39485.4]
  assign _T_91768 = $signed(_T_70213) + $signed(_GEN_654); // @[Modules.scala 143:103:@39501.4]
  assign _T_91769 = _T_91768[5:0]; // @[Modules.scala 143:103:@39502.4]
  assign _T_91770 = $signed(_T_91769); // @[Modules.scala 143:103:@39503.4]
  assign _T_91775 = $signed(_T_70220) + $signed(_T_60983); // @[Modules.scala 143:103:@39507.4]
  assign _T_91776 = _T_91775[4:0]; // @[Modules.scala 143:103:@39508.4]
  assign _T_91777 = $signed(_T_91776); // @[Modules.scala 143:103:@39509.4]
  assign _GEN_860 = {{1{_T_54915[4]}},_T_54915}; // @[Modules.scala 143:103:@39519.4]
  assign _T_91789 = $signed(_GEN_860) + $signed(_T_64115); // @[Modules.scala 143:103:@39519.4]
  assign _T_91790 = _T_91789[5:0]; // @[Modules.scala 143:103:@39520.4]
  assign _T_91791 = $signed(_T_91790); // @[Modules.scala 143:103:@39521.4]
  assign _T_91859 = $signed(_GEN_26) + $signed(_T_58025); // @[Modules.scala 143:103:@39579.4]
  assign _T_91860 = _T_91859[5:0]; // @[Modules.scala 143:103:@39580.4]
  assign _T_91861 = $signed(_T_91860); // @[Modules.scala 143:103:@39581.4]
  assign _T_91866 = $signed(_GEN_100) + $signed(_T_61088); // @[Modules.scala 143:103:@39585.4]
  assign _T_91867 = _T_91866[5:0]; // @[Modules.scala 143:103:@39586.4]
  assign _T_91868 = $signed(_T_91867); // @[Modules.scala 143:103:@39587.4]
  assign _T_91873 = $signed(_GEN_658) + $signed(_T_61095); // @[Modules.scala 143:103:@39591.4]
  assign _T_91874 = _T_91873[5:0]; // @[Modules.scala 143:103:@39592.4]
  assign _T_91875 = $signed(_T_91874); // @[Modules.scala 143:103:@39593.4]
  assign _T_91950 = $signed(_T_55090) + $signed(_T_55095); // @[Modules.scala 143:103:@39657.4]
  assign _T_91951 = _T_91950[4:0]; // @[Modules.scala 143:103:@39658.4]
  assign _T_91952 = $signed(_T_91951); // @[Modules.scala 143:103:@39659.4]
  assign _T_91957 = $signed(_T_55102) + $signed(_T_55109); // @[Modules.scala 143:103:@39663.4]
  assign _T_91958 = _T_91957[4:0]; // @[Modules.scala 143:103:@39664.4]
  assign _T_91959 = $signed(_T_91958); // @[Modules.scala 143:103:@39665.4]
  assign _GEN_865 = {{1{_T_76696[4]}},_T_76696}; // @[Modules.scala 143:103:@39687.4]
  assign _T_91985 = $signed(_T_58158) + $signed(_GEN_865); // @[Modules.scala 143:103:@39687.4]
  assign _T_91986 = _T_91985[5:0]; // @[Modules.scala 143:103:@39688.4]
  assign _T_91987 = $signed(_T_91986); // @[Modules.scala 143:103:@39689.4]
  assign _T_92013 = $signed(_GEN_32) + $signed(_T_55165); // @[Modules.scala 143:103:@39711.4]
  assign _T_92014 = _T_92013[5:0]; // @[Modules.scala 143:103:@39712.4]
  assign _T_92015 = $signed(_T_92014); // @[Modules.scala 143:103:@39713.4]
  assign _T_92027 = $signed(_T_61244) + $signed(_T_55179); // @[Modules.scala 143:103:@39723.4]
  assign _T_92028 = _T_92027[4:0]; // @[Modules.scala 143:103:@39724.4]
  assign _T_92029 = $signed(_T_92028); // @[Modules.scala 143:103:@39725.4]
  assign _T_92048 = $signed(_T_55195) + $signed(_T_55200); // @[Modules.scala 143:103:@39741.4]
  assign _T_92049 = _T_92048[4:0]; // @[Modules.scala 143:103:@39742.4]
  assign _T_92050 = $signed(_T_92049); // @[Modules.scala 143:103:@39743.4]
  assign _GEN_872 = {{1{_T_61412[4]}},_T_61412}; // @[Modules.scala 143:103:@39855.4]
  assign _T_92181 = $signed(_GEN_872) + $signed(_T_55328); // @[Modules.scala 143:103:@39855.4]
  assign _T_92182 = _T_92181[5:0]; // @[Modules.scala 143:103:@39856.4]
  assign _T_92183 = $signed(_T_92182); // @[Modules.scala 143:103:@39857.4]
  assign _T_92251 = $signed(_T_64579) + $signed(_T_58401); // @[Modules.scala 143:103:@39915.4]
  assign _T_92252 = _T_92251[4:0]; // @[Modules.scala 143:103:@39916.4]
  assign _T_92253 = $signed(_T_92252); // @[Modules.scala 143:103:@39917.4]
  assign _GEN_874 = {{1{_T_55433[4]}},_T_55433}; // @[Modules.scala 143:103:@39951.4]
  assign _T_92293 = $signed(_T_58438) + $signed(_GEN_874); // @[Modules.scala 143:103:@39951.4]
  assign _T_92294 = _T_92293[5:0]; // @[Modules.scala 143:103:@39952.4]
  assign _T_92295 = $signed(_T_92294); // @[Modules.scala 143:103:@39953.4]
  assign _T_92321 = $signed(_GEN_181) + $signed(_T_55452); // @[Modules.scala 143:103:@39975.4]
  assign _T_92322 = _T_92321[5:0]; // @[Modules.scala 143:103:@39976.4]
  assign _T_92323 = $signed(_T_92322); // @[Modules.scala 143:103:@39977.4]
  assign _GEN_876 = {{1{_T_58471[4]}},_T_58471}; // @[Modules.scala 143:103:@39981.4]
  assign _T_92328 = $signed(_T_55454) + $signed(_GEN_876); // @[Modules.scala 143:103:@39981.4]
  assign _T_92329 = _T_92328[5:0]; // @[Modules.scala 143:103:@39982.4]
  assign _T_92330 = $signed(_T_92329); // @[Modules.scala 143:103:@39983.4]
  assign _T_92335 = $signed(_T_58473) + $signed(_T_55461); // @[Modules.scala 143:103:@39987.4]
  assign _T_92336 = _T_92335[4:0]; // @[Modules.scala 143:103:@39988.4]
  assign _T_92337 = $signed(_T_92336); // @[Modules.scala 143:103:@39989.4]
  assign _T_92349 = $signed(_T_55475) + $signed(_T_58492); // @[Modules.scala 143:103:@39999.4]
  assign _T_92350 = _T_92349[4:0]; // @[Modules.scala 143:103:@40000.4]
  assign _T_92351 = $signed(_T_92350); // @[Modules.scala 143:103:@40001.4]
  assign _GEN_878 = {{1{_T_58520[4]}},_T_58520}; // @[Modules.scala 143:103:@40023.4]
  assign _T_92377 = $signed(_T_55496) + $signed(_GEN_878); // @[Modules.scala 143:103:@40023.4]
  assign _T_92378 = _T_92377[5:0]; // @[Modules.scala 143:103:@40024.4]
  assign _T_92379 = $signed(_T_92378); // @[Modules.scala 143:103:@40025.4]
  assign _T_92405 = $signed(_T_58543) + $signed(_T_70815); // @[Modules.scala 143:103:@40047.4]
  assign _T_92406 = _T_92405[4:0]; // @[Modules.scala 143:103:@40048.4]
  assign _T_92407 = $signed(_T_92406); // @[Modules.scala 143:103:@40049.4]
  assign _T_92503 = $signed(_T_70904) + $signed(_T_70918); // @[Modules.scala 143:103:@40131.4]
  assign _T_92504 = _T_92503[5:0]; // @[Modules.scala 143:103:@40132.4]
  assign _T_92505 = $signed(_T_92504); // @[Modules.scala 143:103:@40133.4]
  assign _T_92510 = $signed(_T_55627) + $signed(_GEN_672); // @[Modules.scala 143:103:@40137.4]
  assign _T_92511 = _T_92510[5:0]; // @[Modules.scala 143:103:@40138.4]
  assign _T_92512 = $signed(_T_92511); // @[Modules.scala 143:103:@40139.4]
  assign _T_92573 = $signed(_GEN_194) + $signed(_T_55699); // @[Modules.scala 143:103:@40191.4]
  assign _T_92574 = _T_92573[5:0]; // @[Modules.scala 143:103:@40192.4]
  assign _T_92575 = $signed(_T_92574); // @[Modules.scala 143:103:@40193.4]
  assign _T_92580 = $signed(_T_70990) + $signed(_GEN_121); // @[Modules.scala 143:103:@40197.4]
  assign _T_92581 = _T_92580[5:0]; // @[Modules.scala 143:103:@40198.4]
  assign _T_92582 = $signed(_T_92581); // @[Modules.scala 143:103:@40199.4]
  assign _GEN_884 = {{1{_T_58725[4]}},_T_58725}; // @[Modules.scala 143:103:@40203.4]
  assign _T_92587 = $signed(_T_71004) + $signed(_GEN_884); // @[Modules.scala 143:103:@40203.4]
  assign _T_92588 = _T_92587[5:0]; // @[Modules.scala 143:103:@40204.4]
  assign _T_92589 = $signed(_T_92588); // @[Modules.scala 143:103:@40205.4]
  assign _T_92636 = $signed(_T_77382) + $signed(_T_55748); // @[Modules.scala 143:103:@40245.4]
  assign _T_92637 = _T_92636[5:0]; // @[Modules.scala 143:103:@40246.4]
  assign _T_92638 = $signed(_T_92637); // @[Modules.scala 143:103:@40247.4]
  assign _T_92643 = $signed(_T_55753) + $signed(_GEN_742); // @[Modules.scala 143:103:@40251.4]
  assign _T_92644 = _T_92643[5:0]; // @[Modules.scala 143:103:@40252.4]
  assign _T_92645 = $signed(_T_92644); // @[Modules.scala 143:103:@40253.4]
  assign _GEN_886 = {{1{_T_58793[4]}},_T_58793}; // @[Modules.scala 143:103:@40275.4]
  assign _T_92671 = $signed(_T_58788) + $signed(_GEN_886); // @[Modules.scala 143:103:@40275.4]
  assign _T_92672 = _T_92671[5:0]; // @[Modules.scala 143:103:@40276.4]
  assign _T_92673 = $signed(_T_92672); // @[Modules.scala 143:103:@40277.4]
  assign _T_92720 = $signed(_T_71137) + $signed(_T_55816); // @[Modules.scala 143:103:@40317.4]
  assign _T_92721 = _T_92720[5:0]; // @[Modules.scala 143:103:@40318.4]
  assign _T_92722 = $signed(_T_92721); // @[Modules.scala 143:103:@40319.4]
  assign _T_92727 = $signed(_T_77464) + $signed(_T_55818); // @[Modules.scala 143:103:@40323.4]
  assign _T_92728 = _T_92727[5:0]; // @[Modules.scala 143:103:@40324.4]
  assign _T_92729 = $signed(_T_92728); // @[Modules.scala 143:103:@40325.4]
  assign _T_92734 = $signed(_T_55823) + $signed(_T_61923); // @[Modules.scala 143:103:@40329.4]
  assign _T_92735 = _T_92734[5:0]; // @[Modules.scala 143:103:@40330.4]
  assign _T_92736 = $signed(_T_92735); // @[Modules.scala 143:103:@40331.4]
  assign _GEN_888 = {{1{_T_71163[4]}},_T_71163}; // @[Modules.scala 143:103:@40335.4]
  assign _T_92741 = $signed(_T_55825) + $signed(_GEN_888); // @[Modules.scala 143:103:@40335.4]
  assign _T_92742 = _T_92741[5:0]; // @[Modules.scala 143:103:@40336.4]
  assign _T_92743 = $signed(_T_92742); // @[Modules.scala 143:103:@40337.4]
  assign _GEN_889 = {{1{_T_58851[4]}},_T_58851}; // @[Modules.scala 143:103:@40341.4]
  assign _T_92748 = $signed(_GEN_889) + $signed(_T_58858); // @[Modules.scala 143:103:@40341.4]
  assign _T_92749 = _T_92748[5:0]; // @[Modules.scala 143:103:@40342.4]
  assign _T_92750 = $signed(_T_92749); // @[Modules.scala 143:103:@40343.4]
  assign _GEN_891 = {{1{_T_62000[4]}},_T_62000}; // @[Modules.scala 143:103:@40383.4]
  assign _T_92797 = $signed(_T_55879) + $signed(_GEN_891); // @[Modules.scala 143:103:@40383.4]
  assign _T_92798 = _T_92797[5:0]; // @[Modules.scala 143:103:@40384.4]
  assign _T_92799 = $signed(_T_92798); // @[Modules.scala 143:103:@40385.4]
  assign _T_92804 = $signed(_T_71235) + $signed(_T_71240); // @[Modules.scala 143:103:@40389.4]
  assign _T_92805 = _T_92804[5:0]; // @[Modules.scala 143:103:@40390.4]
  assign _T_92806 = $signed(_T_92805); // @[Modules.scala 143:103:@40391.4]
  assign _T_92811 = $signed(_T_71242) + $signed(_GEN_818); // @[Modules.scala 143:103:@40395.4]
  assign _T_92812 = _T_92811[5:0]; // @[Modules.scala 143:103:@40396.4]
  assign _T_92813 = $signed(_T_92812); // @[Modules.scala 143:103:@40397.4]
  assign _T_92825 = $signed(_GEN_419) + $signed(_T_55923); // @[Modules.scala 143:103:@40407.4]
  assign _T_92826 = _T_92825[5:0]; // @[Modules.scala 143:103:@40408.4]
  assign _T_92827 = $signed(_T_92826); // @[Modules.scala 143:103:@40409.4]
  assign _T_92846 = $signed(_GEN_819) + $signed(_T_55949); // @[Modules.scala 143:103:@40425.4]
  assign _T_92847 = _T_92846[5:0]; // @[Modules.scala 143:103:@40426.4]
  assign _T_92848 = $signed(_T_92847); // @[Modules.scala 143:103:@40427.4]
  assign _T_92888 = $signed(_T_71317) + $signed(_T_65195); // @[Modules.scala 143:103:@40461.4]
  assign _T_92889 = _T_92888[5:0]; // @[Modules.scala 143:103:@40462.4]
  assign _T_92890 = $signed(_T_92889); // @[Modules.scala 143:103:@40463.4]
  assign _T_92902 = $signed(_T_59005) + $signed(_T_62110); // @[Modules.scala 143:103:@40473.4]
  assign _T_92903 = _T_92902[5:0]; // @[Modules.scala 143:103:@40474.4]
  assign _T_92904 = $signed(_T_92903); // @[Modules.scala 143:103:@40475.4]
  assign _T_92909 = $signed(_T_56014) + $signed(_T_59017); // @[Modules.scala 143:103:@40479.4]
  assign _T_92910 = _T_92909[4:0]; // @[Modules.scala 143:103:@40480.4]
  assign _T_92911 = $signed(_T_92910); // @[Modules.scala 143:103:@40481.4]
  assign _T_92916 = $signed(_T_59019) + $signed(_T_59024); // @[Modules.scala 143:103:@40485.4]
  assign _T_92917 = _T_92916[4:0]; // @[Modules.scala 143:103:@40486.4]
  assign _T_92918 = $signed(_T_92917); // @[Modules.scala 143:103:@40487.4]
  assign _T_92923 = $signed(_GEN_821) + $signed(_T_56026); // @[Modules.scala 143:103:@40491.4]
  assign _T_92924 = _T_92923[5:0]; // @[Modules.scala 143:103:@40492.4]
  assign _T_92925 = $signed(_T_92924); // @[Modules.scala 143:103:@40493.4]
  assign _T_92958 = $signed(_T_62159) + $signed(_T_59061); // @[Modules.scala 143:103:@40521.4]
  assign _T_92959 = _T_92958[5:0]; // @[Modules.scala 143:103:@40522.4]
  assign _T_92960 = $signed(_T_92959); // @[Modules.scala 143:103:@40523.4]
  assign _T_92972 = $signed(_T_59080) + $signed(_GEN_353); // @[Modules.scala 143:103:@40533.4]
  assign _T_92973 = _T_92972[5:0]; // @[Modules.scala 143:103:@40534.4]
  assign _T_92974 = $signed(_T_92973); // @[Modules.scala 143:103:@40535.4]
  assign _T_92993 = $signed(_T_62189) + $signed(_GEN_69); // @[Modules.scala 143:103:@40551.4]
  assign _T_92994 = _T_92993[5:0]; // @[Modules.scala 143:103:@40552.4]
  assign _T_92995 = $signed(_T_92994); // @[Modules.scala 143:103:@40553.4]
  assign _T_93007 = $signed(_GEN_208) + $signed(_T_56117); // @[Modules.scala 143:103:@40563.4]
  assign _T_93008 = _T_93007[5:0]; // @[Modules.scala 143:103:@40564.4]
  assign _T_93009 = $signed(_T_93008); // @[Modules.scala 143:103:@40565.4]
  assign _GEN_903 = {{1{_T_56152[4]}},_T_56152}; // @[Modules.scala 143:103:@40593.4]
  assign _T_93042 = $signed(_T_59157) + $signed(_GEN_903); // @[Modules.scala 143:103:@40593.4]
  assign _T_93043 = _T_93042[5:0]; // @[Modules.scala 143:103:@40594.4]
  assign _T_93044 = $signed(_T_93043); // @[Modules.scala 143:103:@40595.4]
  assign _GEN_904 = {{1{_T_56168[4]}},_T_56168}; // @[Modules.scala 143:103:@40611.4]
  assign _T_93063 = $signed(_GEN_904) + $signed(_T_59180); // @[Modules.scala 143:103:@40611.4]
  assign _T_93064 = _T_93063[5:0]; // @[Modules.scala 143:103:@40612.4]
  assign _T_93065 = $signed(_T_93064); // @[Modules.scala 143:103:@40613.4]
  assign _T_93077 = $signed(_T_56182) + $signed(_T_56189); // @[Modules.scala 143:103:@40623.4]
  assign _T_93078 = _T_93077[4:0]; // @[Modules.scala 143:103:@40624.4]
  assign _T_93079 = $signed(_T_93078); // @[Modules.scala 143:103:@40625.4]
  assign _T_93091 = $signed(_GEN_140) + $signed(_T_59206); // @[Modules.scala 143:103:@40635.4]
  assign _T_93092 = _T_93091[5:0]; // @[Modules.scala 143:103:@40636.4]
  assign _T_93093 = $signed(_T_93092); // @[Modules.scala 143:103:@40637.4]
  assign _T_93154 = $signed(_T_65475) + $signed(_T_62362); // @[Modules.scala 143:103:@40689.4]
  assign _T_93155 = _T_93154[4:0]; // @[Modules.scala 143:103:@40690.4]
  assign _T_93156 = $signed(_T_93155); // @[Modules.scala 143:103:@40691.4]
  assign _T_93203 = $signed(_GEN_497) + $signed(_T_56299); // @[Modules.scala 143:103:@40731.4]
  assign _T_93204 = _T_93203[5:0]; // @[Modules.scala 143:103:@40732.4]
  assign _T_93205 = $signed(_T_93204); // @[Modules.scala 143:103:@40733.4]
  assign buffer_12_0 = {{8{_T_91133[5]}},_T_91133}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_1 = {{8{_T_91140[5]}},_T_91140}; // @[Modules.scala 112:22:@8.4]
  assign _T_93213 = $signed(buffer_12_0) + $signed(buffer_12_1); // @[Modules.scala 160:64:@40741.4]
  assign _T_93214 = _T_93213[13:0]; // @[Modules.scala 160:64:@40742.4]
  assign buffer_12_298 = $signed(_T_93214); // @[Modules.scala 160:64:@40743.4]
  assign buffer_12_5 = {{8{_T_91168[5]}},_T_91168}; // @[Modules.scala 112:22:@8.4]
  assign _T_93219 = $signed(buffer_10_3) + $signed(buffer_12_5); // @[Modules.scala 160:64:@40749.4]
  assign _T_93220 = _T_93219[13:0]; // @[Modules.scala 160:64:@40750.4]
  assign buffer_12_300 = $signed(_T_93220); // @[Modules.scala 160:64:@40751.4]
  assign buffer_12_9 = {{8{_T_91196[5]}},_T_91196}; // @[Modules.scala 112:22:@8.4]
  assign _T_93225 = $signed(buffer_0_8) + $signed(buffer_12_9); // @[Modules.scala 160:64:@40757.4]
  assign _T_93226 = _T_93225[13:0]; // @[Modules.scala 160:64:@40758.4]
  assign buffer_12_302 = $signed(_T_93226); // @[Modules.scala 160:64:@40759.4]
  assign buffer_12_11 = {{8{_T_91210[5]}},_T_91210}; // @[Modules.scala 112:22:@8.4]
  assign _T_93228 = $signed(buffer_1_9) + $signed(buffer_12_11); // @[Modules.scala 160:64:@40761.4]
  assign _T_93229 = _T_93228[13:0]; // @[Modules.scala 160:64:@40762.4]
  assign buffer_12_303 = $signed(_T_93229); // @[Modules.scala 160:64:@40763.4]
  assign buffer_12_13 = {{9{_T_91224[4]}},_T_91224}; // @[Modules.scala 112:22:@8.4]
  assign _T_93231 = $signed(buffer_3_12) + $signed(buffer_12_13); // @[Modules.scala 160:64:@40765.4]
  assign _T_93232 = _T_93231[13:0]; // @[Modules.scala 160:64:@40766.4]
  assign buffer_12_304 = $signed(_T_93232); // @[Modules.scala 160:64:@40767.4]
  assign buffer_12_14 = {{8{_T_91231[5]}},_T_91231}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_15 = {{8{_T_91238[5]}},_T_91238}; // @[Modules.scala 112:22:@8.4]
  assign _T_93234 = $signed(buffer_12_14) + $signed(buffer_12_15); // @[Modules.scala 160:64:@40769.4]
  assign _T_93235 = _T_93234[13:0]; // @[Modules.scala 160:64:@40770.4]
  assign buffer_12_305 = $signed(_T_93235); // @[Modules.scala 160:64:@40771.4]
  assign buffer_12_16 = {{8{_T_91245[5]}},_T_91245}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_17 = {{8{_T_91252[5]}},_T_91252}; // @[Modules.scala 112:22:@8.4]
  assign _T_93237 = $signed(buffer_12_16) + $signed(buffer_12_17); // @[Modules.scala 160:64:@40773.4]
  assign _T_93238 = _T_93237[13:0]; // @[Modules.scala 160:64:@40774.4]
  assign buffer_12_306 = $signed(_T_93238); // @[Modules.scala 160:64:@40775.4]
  assign _T_93240 = $signed(buffer_9_22) + $signed(buffer_8_24); // @[Modules.scala 160:64:@40777.4]
  assign _T_93241 = _T_93240[13:0]; // @[Modules.scala 160:64:@40778.4]
  assign buffer_12_307 = $signed(_T_93241); // @[Modules.scala 160:64:@40779.4]
  assign _T_93243 = $signed(buffer_0_23) + $signed(buffer_3_23); // @[Modules.scala 160:64:@40781.4]
  assign _T_93244 = _T_93243[13:0]; // @[Modules.scala 160:64:@40782.4]
  assign buffer_12_308 = $signed(_T_93244); // @[Modules.scala 160:64:@40783.4]
  assign buffer_12_27 = {{9{_T_91322[4]}},_T_91322}; // @[Modules.scala 112:22:@8.4]
  assign _T_93252 = $signed(buffer_3_28) + $signed(buffer_12_27); // @[Modules.scala 160:64:@40793.4]
  assign _T_93253 = _T_93252[13:0]; // @[Modules.scala 160:64:@40794.4]
  assign buffer_12_311 = $signed(_T_93253); // @[Modules.scala 160:64:@40795.4]
  assign _T_93255 = $signed(buffer_0_32) + $signed(buffer_8_34); // @[Modules.scala 160:64:@40797.4]
  assign _T_93256 = _T_93255[13:0]; // @[Modules.scala 160:64:@40798.4]
  assign buffer_12_312 = $signed(_T_93256); // @[Modules.scala 160:64:@40799.4]
  assign _T_93258 = $signed(buffer_8_35) + $signed(buffer_4_33); // @[Modules.scala 160:64:@40801.4]
  assign _T_93259 = _T_93258[13:0]; // @[Modules.scala 160:64:@40802.4]
  assign buffer_12_313 = $signed(_T_93259); // @[Modules.scala 160:64:@40803.4]
  assign buffer_12_33 = {{8{_T_91364[5]}},_T_91364}; // @[Modules.scala 112:22:@8.4]
  assign _T_93261 = $signed(buffer_4_34) + $signed(buffer_12_33); // @[Modules.scala 160:64:@40805.4]
  assign _T_93262 = _T_93261[13:0]; // @[Modules.scala 160:64:@40806.4]
  assign buffer_12_314 = $signed(_T_93262); // @[Modules.scala 160:64:@40807.4]
  assign buffer_12_35 = {{8{_T_91378[5]}},_T_91378}; // @[Modules.scala 112:22:@8.4]
  assign _T_93264 = $signed(buffer_1_36) + $signed(buffer_12_35); // @[Modules.scala 160:64:@40809.4]
  assign _T_93265 = _T_93264[13:0]; // @[Modules.scala 160:64:@40810.4]
  assign buffer_12_315 = $signed(_T_93265); // @[Modules.scala 160:64:@40811.4]
  assign buffer_12_36 = {{9{_T_91385[4]}},_T_91385}; // @[Modules.scala 112:22:@8.4]
  assign _T_93267 = $signed(buffer_12_36) + $signed(buffer_0_42); // @[Modules.scala 160:64:@40813.4]
  assign _T_93268 = _T_93267[13:0]; // @[Modules.scala 160:64:@40814.4]
  assign buffer_12_316 = $signed(_T_93268); // @[Modules.scala 160:64:@40815.4]
  assign buffer_12_38 = {{8{_T_91399[5]}},_T_91399}; // @[Modules.scala 112:22:@8.4]
  assign _T_93270 = $signed(buffer_12_38) + $signed(buffer_1_42); // @[Modules.scala 160:64:@40817.4]
  assign _T_93271 = _T_93270[13:0]; // @[Modules.scala 160:64:@40818.4]
  assign buffer_12_317 = $signed(_T_93271); // @[Modules.scala 160:64:@40819.4]
  assign buffer_12_41 = {{8{_T_91420[5]}},_T_91420}; // @[Modules.scala 112:22:@8.4]
  assign _T_93273 = $signed(buffer_1_43) + $signed(buffer_12_41); // @[Modules.scala 160:64:@40821.4]
  assign _T_93274 = _T_93273[13:0]; // @[Modules.scala 160:64:@40822.4]
  assign buffer_12_318 = $signed(_T_93274); // @[Modules.scala 160:64:@40823.4]
  assign buffer_12_43 = {{8{_T_91434[5]}},_T_91434}; // @[Modules.scala 112:22:@8.4]
  assign _T_93276 = $signed(buffer_1_45) + $signed(buffer_12_43); // @[Modules.scala 160:64:@40825.4]
  assign _T_93277 = _T_93276[13:0]; // @[Modules.scala 160:64:@40826.4]
  assign buffer_12_319 = $signed(_T_93277); // @[Modules.scala 160:64:@40827.4]
  assign buffer_12_44 = {{9{_T_91441[4]}},_T_91441}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_45 = {{8{_T_91448[5]}},_T_91448}; // @[Modules.scala 112:22:@8.4]
  assign _T_93279 = $signed(buffer_12_44) + $signed(buffer_12_45); // @[Modules.scala 160:64:@40829.4]
  assign _T_93280 = _T_93279[13:0]; // @[Modules.scala 160:64:@40830.4]
  assign buffer_12_320 = $signed(_T_93280); // @[Modules.scala 160:64:@40831.4]
  assign buffer_12_46 = {{8{_T_91455[5]}},_T_91455}; // @[Modules.scala 112:22:@8.4]
  assign _T_93282 = $signed(buffer_12_46) + $signed(buffer_7_52); // @[Modules.scala 160:64:@40833.4]
  assign _T_93283 = _T_93282[13:0]; // @[Modules.scala 160:64:@40834.4]
  assign buffer_12_321 = $signed(_T_93283); // @[Modules.scala 160:64:@40835.4]
  assign _T_93285 = $signed(buffer_7_53) + $signed(buffer_7_54); // @[Modules.scala 160:64:@40837.4]
  assign _T_93286 = _T_93285[13:0]; // @[Modules.scala 160:64:@40838.4]
  assign buffer_12_322 = $signed(_T_93286); // @[Modules.scala 160:64:@40839.4]
  assign buffer_12_50 = {{8{_T_91483[5]}},_T_91483}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_51 = {{8{_T_91490[5]}},_T_91490}; // @[Modules.scala 112:22:@8.4]
  assign _T_93288 = $signed(buffer_12_50) + $signed(buffer_12_51); // @[Modules.scala 160:64:@40841.4]
  assign _T_93289 = _T_93288[13:0]; // @[Modules.scala 160:64:@40842.4]
  assign buffer_12_323 = $signed(_T_93289); // @[Modules.scala 160:64:@40843.4]
  assign buffer_12_53 = {{8{_T_91504[5]}},_T_91504}; // @[Modules.scala 112:22:@8.4]
  assign _T_93291 = $signed(buffer_3_60) + $signed(buffer_12_53); // @[Modules.scala 160:64:@40845.4]
  assign _T_93292 = _T_93291[13:0]; // @[Modules.scala 160:64:@40846.4]
  assign buffer_12_324 = $signed(_T_93292); // @[Modules.scala 160:64:@40847.4]
  assign _T_93294 = $signed(buffer_5_61) + $signed(buffer_1_61); // @[Modules.scala 160:64:@40849.4]
  assign _T_93295 = _T_93294[13:0]; // @[Modules.scala 160:64:@40850.4]
  assign buffer_12_325 = $signed(_T_93295); // @[Modules.scala 160:64:@40851.4]
  assign buffer_12_57 = {{8{_T_91532[5]}},_T_91532}; // @[Modules.scala 112:22:@8.4]
  assign _T_93297 = $signed(buffer_8_59) + $signed(buffer_12_57); // @[Modules.scala 160:64:@40853.4]
  assign _T_93298 = _T_93297[13:0]; // @[Modules.scala 160:64:@40854.4]
  assign buffer_12_326 = $signed(_T_93298); // @[Modules.scala 160:64:@40855.4]
  assign _T_93300 = $signed(buffer_8_61) + $signed(buffer_8_62); // @[Modules.scala 160:64:@40857.4]
  assign _T_93301 = _T_93300[13:0]; // @[Modules.scala 160:64:@40858.4]
  assign buffer_12_327 = $signed(_T_93301); // @[Modules.scala 160:64:@40859.4]
  assign buffer_12_60 = {{8{_T_91553[5]}},_T_91553}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_61 = {{8{_T_91560[5]}},_T_91560}; // @[Modules.scala 112:22:@8.4]
  assign _T_93303 = $signed(buffer_12_60) + $signed(buffer_12_61); // @[Modules.scala 160:64:@40861.4]
  assign _T_93304 = _T_93303[13:0]; // @[Modules.scala 160:64:@40862.4]
  assign buffer_12_328 = $signed(_T_93304); // @[Modules.scala 160:64:@40863.4]
  assign buffer_12_62 = {{8{_T_91567[5]}},_T_91567}; // @[Modules.scala 112:22:@8.4]
  assign _T_93306 = $signed(buffer_12_62) + $signed(buffer_3_72); // @[Modules.scala 160:64:@40865.4]
  assign _T_93307 = _T_93306[13:0]; // @[Modules.scala 160:64:@40866.4]
  assign buffer_12_329 = $signed(_T_93307); // @[Modules.scala 160:64:@40867.4]
  assign _T_93309 = $signed(buffer_9_74) + $signed(buffer_3_75); // @[Modules.scala 160:64:@40869.4]
  assign _T_93310 = _T_93309[13:0]; // @[Modules.scala 160:64:@40870.4]
  assign buffer_12_330 = $signed(_T_93310); // @[Modules.scala 160:64:@40871.4]
  assign buffer_12_67 = {{8{_T_91602[5]}},_T_91602}; // @[Modules.scala 112:22:@8.4]
  assign _T_93312 = $signed(buffer_5_76) + $signed(buffer_12_67); // @[Modules.scala 160:64:@40873.4]
  assign _T_93313 = _T_93312[13:0]; // @[Modules.scala 160:64:@40874.4]
  assign buffer_12_331 = $signed(_T_93313); // @[Modules.scala 160:64:@40875.4]
  assign buffer_12_70 = {{8{_T_91623[5]}},_T_91623}; // @[Modules.scala 112:22:@8.4]
  assign _T_93318 = $signed(buffer_12_70) + $signed(buffer_2_80); // @[Modules.scala 160:64:@40881.4]
  assign _T_93319 = _T_93318[13:0]; // @[Modules.scala 160:64:@40882.4]
  assign buffer_12_333 = $signed(_T_93319); // @[Modules.scala 160:64:@40883.4]
  assign buffer_12_73 = {{9{_T_91644[4]}},_T_91644}; // @[Modules.scala 112:22:@8.4]
  assign _T_93321 = $signed(buffer_1_81) + $signed(buffer_12_73); // @[Modules.scala 160:64:@40885.4]
  assign _T_93322 = _T_93321[13:0]; // @[Modules.scala 160:64:@40886.4]
  assign buffer_12_334 = $signed(_T_93322); // @[Modules.scala 160:64:@40887.4]
  assign buffer_12_74 = {{8{_T_91651[5]}},_T_91651}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_75 = {{8{_T_91658[5]}},_T_91658}; // @[Modules.scala 112:22:@8.4]
  assign _T_93324 = $signed(buffer_12_74) + $signed(buffer_12_75); // @[Modules.scala 160:64:@40889.4]
  assign _T_93325 = _T_93324[13:0]; // @[Modules.scala 160:64:@40890.4]
  assign buffer_12_335 = $signed(_T_93325); // @[Modules.scala 160:64:@40891.4]
  assign buffer_12_76 = {{8{_T_91665[5]}},_T_91665}; // @[Modules.scala 112:22:@8.4]
  assign _T_93327 = $signed(buffer_12_76) + $signed(buffer_3_90); // @[Modules.scala 160:64:@40893.4]
  assign _T_93328 = _T_93327[13:0]; // @[Modules.scala 160:64:@40894.4]
  assign buffer_12_336 = $signed(_T_93328); // @[Modules.scala 160:64:@40895.4]
  assign buffer_12_81 = {{8{_T_91700[5]}},_T_91700}; // @[Modules.scala 112:22:@8.4]
  assign _T_93333 = $signed(buffer_8_86) + $signed(buffer_12_81); // @[Modules.scala 160:64:@40901.4]
  assign _T_93334 = _T_93333[13:0]; // @[Modules.scala 160:64:@40902.4]
  assign buffer_12_338 = $signed(_T_93334); // @[Modules.scala 160:64:@40903.4]
  assign _T_93336 = $signed(buffer_8_89) + $signed(buffer_0_90); // @[Modules.scala 160:64:@40905.4]
  assign _T_93337 = _T_93336[13:0]; // @[Modules.scala 160:64:@40906.4]
  assign buffer_12_339 = $signed(_T_93337); // @[Modules.scala 160:64:@40907.4]
  assign _T_93339 = $signed(buffer_0_91) + $signed(buffer_3_98); // @[Modules.scala 160:64:@40909.4]
  assign _T_93340 = _T_93339[13:0]; // @[Modules.scala 160:64:@40910.4]
  assign buffer_12_340 = $signed(_T_93340); // @[Modules.scala 160:64:@40911.4]
  assign _T_93342 = $signed(buffer_3_99) + $signed(buffer_0_94); // @[Modules.scala 160:64:@40913.4]
  assign _T_93343 = _T_93342[13:0]; // @[Modules.scala 160:64:@40914.4]
  assign buffer_12_341 = $signed(_T_93343); // @[Modules.scala 160:64:@40915.4]
  assign buffer_12_88 = {{8{_T_91749[5]}},_T_91749}; // @[Modules.scala 112:22:@8.4]
  assign _T_93345 = $signed(buffer_12_88) + $signed(buffer_3_103); // @[Modules.scala 160:64:@40917.4]
  assign _T_93346 = _T_93345[13:0]; // @[Modules.scala 160:64:@40918.4]
  assign buffer_12_342 = $signed(_T_93346); // @[Modules.scala 160:64:@40919.4]
  assign buffer_12_91 = {{8{_T_91770[5]}},_T_91770}; // @[Modules.scala 112:22:@8.4]
  assign _T_93348 = $signed(buffer_3_104) + $signed(buffer_12_91); // @[Modules.scala 160:64:@40921.4]
  assign _T_93349 = _T_93348[13:0]; // @[Modules.scala 160:64:@40922.4]
  assign buffer_12_343 = $signed(_T_93349); // @[Modules.scala 160:64:@40923.4]
  assign buffer_12_92 = {{9{_T_91777[4]}},_T_91777}; // @[Modules.scala 112:22:@8.4]
  assign _T_93351 = $signed(buffer_12_92) + $signed(buffer_1_104); // @[Modules.scala 160:64:@40925.4]
  assign _T_93352 = _T_93351[13:0]; // @[Modules.scala 160:64:@40926.4]
  assign buffer_12_344 = $signed(_T_93352); // @[Modules.scala 160:64:@40927.4]
  assign buffer_12_94 = {{8{_T_91791[5]}},_T_91791}; // @[Modules.scala 112:22:@8.4]
  assign _T_93354 = $signed(buffer_12_94) + $signed(buffer_0_105); // @[Modules.scala 160:64:@40929.4]
  assign _T_93355 = _T_93354[13:0]; // @[Modules.scala 160:64:@40930.4]
  assign buffer_12_345 = $signed(_T_93355); // @[Modules.scala 160:64:@40931.4]
  assign _T_93357 = $signed(buffer_1_108) + $signed(buffer_3_113); // @[Modules.scala 160:64:@40933.4]
  assign _T_93358 = _T_93357[13:0]; // @[Modules.scala 160:64:@40934.4]
  assign buffer_12_346 = $signed(_T_93358); // @[Modules.scala 160:64:@40935.4]
  assign buffer_12_104 = {{8{_T_91861[5]}},_T_91861}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_105 = {{8{_T_91868[5]}},_T_91868}; // @[Modules.scala 112:22:@8.4]
  assign _T_93369 = $signed(buffer_12_104) + $signed(buffer_12_105); // @[Modules.scala 160:64:@40949.4]
  assign _T_93370 = _T_93369[13:0]; // @[Modules.scala 160:64:@40950.4]
  assign buffer_12_350 = $signed(_T_93370); // @[Modules.scala 160:64:@40951.4]
  assign buffer_12_106 = {{8{_T_91875[5]}},_T_91875}; // @[Modules.scala 112:22:@8.4]
  assign _T_93372 = $signed(buffer_12_106) + $signed(buffer_3_125); // @[Modules.scala 160:64:@40953.4]
  assign _T_93373 = _T_93372[13:0]; // @[Modules.scala 160:64:@40954.4]
  assign buffer_12_351 = $signed(_T_93373); // @[Modules.scala 160:64:@40955.4]
  assign _T_93375 = $signed(buffer_1_121) + $signed(buffer_9_127); // @[Modules.scala 160:64:@40957.4]
  assign _T_93376 = _T_93375[13:0]; // @[Modules.scala 160:64:@40958.4]
  assign buffer_12_352 = $signed(_T_93376); // @[Modules.scala 160:64:@40959.4]
  assign buffer_12_117 = {{9{_T_91952[4]}},_T_91952}; // @[Modules.scala 112:22:@8.4]
  assign _T_93387 = $signed(buffer_9_134) + $signed(buffer_12_117); // @[Modules.scala 160:64:@40973.4]
  assign _T_93388 = _T_93387[13:0]; // @[Modules.scala 160:64:@40974.4]
  assign buffer_12_356 = $signed(_T_93388); // @[Modules.scala 160:64:@40975.4]
  assign buffer_12_118 = {{9{_T_91959[4]}},_T_91959}; // @[Modules.scala 112:22:@8.4]
  assign _T_93390 = $signed(buffer_12_118) + $signed(buffer_2_133); // @[Modules.scala 160:64:@40977.4]
  assign _T_93391 = _T_93390[13:0]; // @[Modules.scala 160:64:@40978.4]
  assign buffer_12_357 = $signed(_T_93391); // @[Modules.scala 160:64:@40979.4]
  assign buffer_12_122 = {{8{_T_91987[5]}},_T_91987}; // @[Modules.scala 112:22:@8.4]
  assign _T_93396 = $signed(buffer_12_122) + $signed(buffer_9_142); // @[Modules.scala 160:64:@40985.4]
  assign _T_93397 = _T_93396[13:0]; // @[Modules.scala 160:64:@40986.4]
  assign buffer_12_359 = $signed(_T_93397); // @[Modules.scala 160:64:@40987.4]
  assign _T_93399 = $signed(buffer_0_135) + $signed(buffer_2_139); // @[Modules.scala 160:64:@40989.4]
  assign _T_93400 = _T_93399[13:0]; // @[Modules.scala 160:64:@40990.4]
  assign buffer_12_360 = $signed(_T_93400); // @[Modules.scala 160:64:@40991.4]
  assign buffer_12_126 = {{8{_T_92015[5]}},_T_92015}; // @[Modules.scala 112:22:@8.4]
  assign _T_93402 = $signed(buffer_12_126) + $signed(buffer_1_140); // @[Modules.scala 160:64:@40993.4]
  assign _T_93403 = _T_93402[13:0]; // @[Modules.scala 160:64:@40994.4]
  assign buffer_12_361 = $signed(_T_93403); // @[Modules.scala 160:64:@40995.4]
  assign buffer_12_128 = {{9{_T_92029[4]}},_T_92029}; // @[Modules.scala 112:22:@8.4]
  assign _T_93405 = $signed(buffer_12_128) + $signed(buffer_5_143); // @[Modules.scala 160:64:@40997.4]
  assign _T_93406 = _T_93405[13:0]; // @[Modules.scala 160:64:@40998.4]
  assign buffer_12_362 = $signed(_T_93406); // @[Modules.scala 160:64:@40999.4]
  assign buffer_12_131 = {{9{_T_92050[4]}},_T_92050}; // @[Modules.scala 112:22:@8.4]
  assign _T_93408 = $signed(buffer_5_144) + $signed(buffer_12_131); // @[Modules.scala 160:64:@41001.4]
  assign _T_93409 = _T_93408[13:0]; // @[Modules.scala 160:64:@41002.4]
  assign buffer_12_363 = $signed(_T_93409); // @[Modules.scala 160:64:@41003.4]
  assign _T_93414 = $signed(buffer_0_146) + $signed(buffer_1_149); // @[Modules.scala 160:64:@41009.4]
  assign _T_93415 = _T_93414[13:0]; // @[Modules.scala 160:64:@41010.4]
  assign buffer_12_365 = $signed(_T_93415); // @[Modules.scala 160:64:@41011.4]
  assign _T_93417 = $signed(buffer_1_150) + $signed(buffer_2_153); // @[Modules.scala 160:64:@41013.4]
  assign _T_93418 = _T_93417[13:0]; // @[Modules.scala 160:64:@41014.4]
  assign buffer_12_366 = $signed(_T_93418); // @[Modules.scala 160:64:@41015.4]
  assign _T_93420 = $signed(buffer_2_154) + $signed(buffer_8_150); // @[Modules.scala 160:64:@41017.4]
  assign _T_93421 = _T_93420[13:0]; // @[Modules.scala 160:64:@41018.4]
  assign buffer_12_367 = $signed(_T_93421); // @[Modules.scala 160:64:@41019.4]
  assign _T_93426 = $signed(buffer_5_154) + $signed(buffer_2_160); // @[Modules.scala 160:64:@41025.4]
  assign _T_93427 = _T_93426[13:0]; // @[Modules.scala 160:64:@41026.4]
  assign buffer_12_369 = $signed(_T_93427); // @[Modules.scala 160:64:@41027.4]
  assign _T_93429 = $signed(buffer_1_157) + $signed(buffer_0_157); // @[Modules.scala 160:64:@41029.4]
  assign _T_93430 = _T_93429[13:0]; // @[Modules.scala 160:64:@41030.4]
  assign buffer_12_370 = $signed(_T_93430); // @[Modules.scala 160:64:@41031.4]
  assign _T_93432 = $signed(buffer_1_159) + $signed(buffer_1_160); // @[Modules.scala 160:64:@41033.4]
  assign _T_93433 = _T_93432[13:0]; // @[Modules.scala 160:64:@41034.4]
  assign buffer_12_371 = $signed(_T_93433); // @[Modules.scala 160:64:@41035.4]
  assign _T_93435 = $signed(buffer_1_161) + $signed(buffer_1_162); // @[Modules.scala 160:64:@41037.4]
  assign _T_93436 = _T_93435[13:0]; // @[Modules.scala 160:64:@41038.4]
  assign buffer_12_372 = $signed(_T_93436); // @[Modules.scala 160:64:@41039.4]
  assign buffer_12_150 = {{8{_T_92183[5]}},_T_92183}; // @[Modules.scala 112:22:@8.4]
  assign _T_93438 = $signed(buffer_12_150) + $signed(buffer_9_169); // @[Modules.scala 160:64:@41041.4]
  assign _T_93439 = _T_93438[13:0]; // @[Modules.scala 160:64:@41042.4]
  assign buffer_12_373 = $signed(_T_93439); // @[Modules.scala 160:64:@41043.4]
  assign _T_93441 = $signed(buffer_0_163) + $signed(buffer_0_164); // @[Modules.scala 160:64:@41045.4]
  assign _T_93442 = _T_93441[13:0]; // @[Modules.scala 160:64:@41046.4]
  assign buffer_12_374 = $signed(_T_93442); // @[Modules.scala 160:64:@41047.4]
  assign _T_93444 = $signed(buffer_1_166) + $signed(buffer_7_168); // @[Modules.scala 160:64:@41049.4]
  assign _T_93445 = _T_93444[13:0]; // @[Modules.scala 160:64:@41050.4]
  assign buffer_12_375 = $signed(_T_93445); // @[Modules.scala 160:64:@41051.4]
  assign _T_93450 = $signed(buffer_7_171) + $signed(buffer_3_175); // @[Modules.scala 160:64:@41057.4]
  assign _T_93451 = _T_93450[13:0]; // @[Modules.scala 160:64:@41058.4]
  assign buffer_12_377 = $signed(_T_93451); // @[Modules.scala 160:64:@41059.4]
  assign buffer_12_160 = {{9{_T_92253[4]}},_T_92253}; // @[Modules.scala 112:22:@8.4]
  assign _T_93453 = $signed(buffer_12_160) + $signed(buffer_6_177); // @[Modules.scala 160:64:@41061.4]
  assign _T_93454 = _T_93453[13:0]; // @[Modules.scala 160:64:@41062.4]
  assign buffer_12_378 = $signed(_T_93454); // @[Modules.scala 160:64:@41063.4]
  assign _T_93456 = $signed(buffer_8_171) + $signed(buffer_2_178); // @[Modules.scala 160:64:@41065.4]
  assign _T_93457 = _T_93456[13:0]; // @[Modules.scala 160:64:@41066.4]
  assign buffer_12_379 = $signed(_T_93457); // @[Modules.scala 160:64:@41067.4]
  assign _T_93459 = $signed(buffer_8_173) + $signed(buffer_0_175); // @[Modules.scala 160:64:@41069.4]
  assign _T_93460 = _T_93459[13:0]; // @[Modules.scala 160:64:@41070.4]
  assign buffer_12_380 = $signed(_T_93460); // @[Modules.scala 160:64:@41071.4]
  assign buffer_12_166 = {{8{_T_92295[5]}},_T_92295}; // @[Modules.scala 112:22:@8.4]
  assign _T_93462 = $signed(buffer_12_166) + $signed(buffer_8_176); // @[Modules.scala 160:64:@41073.4]
  assign _T_93463 = _T_93462[13:0]; // @[Modules.scala 160:64:@41074.4]
  assign buffer_12_381 = $signed(_T_93463); // @[Modules.scala 160:64:@41075.4]
  assign _T_93465 = $signed(buffer_8_177) + $signed(buffer_4_172); // @[Modules.scala 160:64:@41077.4]
  assign _T_93466 = _T_93465[13:0]; // @[Modules.scala 160:64:@41078.4]
  assign buffer_12_382 = $signed(_T_93466); // @[Modules.scala 160:64:@41079.4]
  assign buffer_12_170 = {{8{_T_92323[5]}},_T_92323}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_171 = {{8{_T_92330[5]}},_T_92330}; // @[Modules.scala 112:22:@8.4]
  assign _T_93468 = $signed(buffer_12_170) + $signed(buffer_12_171); // @[Modules.scala 160:64:@41081.4]
  assign _T_93469 = _T_93468[13:0]; // @[Modules.scala 160:64:@41082.4]
  assign buffer_12_383 = $signed(_T_93469); // @[Modules.scala 160:64:@41083.4]
  assign buffer_12_172 = {{9{_T_92337[4]}},_T_92337}; // @[Modules.scala 112:22:@8.4]
  assign _T_93471 = $signed(buffer_12_172) + $signed(buffer_6_189); // @[Modules.scala 160:64:@41085.4]
  assign _T_93472 = _T_93471[13:0]; // @[Modules.scala 160:64:@41086.4]
  assign buffer_12_384 = $signed(_T_93472); // @[Modules.scala 160:64:@41087.4]
  assign buffer_12_174 = {{9{_T_92351[4]}},_T_92351}; // @[Modules.scala 112:22:@8.4]
  assign _T_93474 = $signed(buffer_12_174) + $signed(buffer_9_192); // @[Modules.scala 160:64:@41089.4]
  assign _T_93475 = _T_93474[13:0]; // @[Modules.scala 160:64:@41090.4]
  assign buffer_12_385 = $signed(_T_93475); // @[Modules.scala 160:64:@41091.4]
  assign _T_93477 = $signed(buffer_2_190) + $signed(buffer_6_193); // @[Modules.scala 160:64:@41093.4]
  assign _T_93478 = _T_93477[13:0]; // @[Modules.scala 160:64:@41094.4]
  assign buffer_12_386 = $signed(_T_93478); // @[Modules.scala 160:64:@41095.4]
  assign buffer_12_178 = {{8{_T_92379[5]}},_T_92379}; // @[Modules.scala 112:22:@8.4]
  assign _T_93480 = $signed(buffer_12_178) + $signed(buffer_8_188); // @[Modules.scala 160:64:@41097.4]
  assign _T_93481 = _T_93480[13:0]; // @[Modules.scala 160:64:@41098.4]
  assign buffer_12_387 = $signed(_T_93481); // @[Modules.scala 160:64:@41099.4]
  assign _T_93483 = $signed(buffer_8_189) + $signed(buffer_8_190); // @[Modules.scala 160:64:@41101.4]
  assign _T_93484 = _T_93483[13:0]; // @[Modules.scala 160:64:@41102.4]
  assign buffer_12_388 = $signed(_T_93484); // @[Modules.scala 160:64:@41103.4]
  assign buffer_12_182 = {{9{_T_92407[4]}},_T_92407}; // @[Modules.scala 112:22:@8.4]
  assign _T_93486 = $signed(buffer_12_182) + $signed(buffer_1_191); // @[Modules.scala 160:64:@41105.4]
  assign _T_93487 = _T_93486[13:0]; // @[Modules.scala 160:64:@41106.4]
  assign buffer_12_389 = $signed(_T_93487); // @[Modules.scala 160:64:@41107.4]
  assign _T_93489 = $signed(buffer_0_190) + $signed(buffer_6_202); // @[Modules.scala 160:64:@41109.4]
  assign _T_93490 = _T_93489[13:0]; // @[Modules.scala 160:64:@41110.4]
  assign buffer_12_390 = $signed(_T_93490); // @[Modules.scala 160:64:@41111.4]
  assign _T_93492 = $signed(buffer_9_203) + $signed(buffer_3_203); // @[Modules.scala 160:64:@41113.4]
  assign _T_93493 = _T_93492[13:0]; // @[Modules.scala 160:64:@41114.4]
  assign buffer_12_391 = $signed(_T_93493); // @[Modules.scala 160:64:@41115.4]
  assign _T_93495 = $signed(buffer_9_205) + $signed(buffer_0_195); // @[Modules.scala 160:64:@41117.4]
  assign _T_93496 = _T_93495[13:0]; // @[Modules.scala 160:64:@41118.4]
  assign buffer_12_392 = $signed(_T_93496); // @[Modules.scala 160:64:@41119.4]
  assign _T_93498 = $signed(buffer_0_196) + $signed(buffer_4_191); // @[Modules.scala 160:64:@41121.4]
  assign _T_93499 = _T_93498[13:0]; // @[Modules.scala 160:64:@41122.4]
  assign buffer_12_393 = $signed(_T_93499); // @[Modules.scala 160:64:@41123.4]
  assign _T_93504 = $signed(buffer_8_203) + $signed(buffer_8_204); // @[Modules.scala 160:64:@41129.4]
  assign _T_93505 = _T_93504[13:0]; // @[Modules.scala 160:64:@41130.4]
  assign buffer_12_395 = $signed(_T_93505); // @[Modules.scala 160:64:@41131.4]
  assign buffer_12_196 = {{8{_T_92505[5]}},_T_92505}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_197 = {{8{_T_92512[5]}},_T_92512}; // @[Modules.scala 112:22:@8.4]
  assign _T_93507 = $signed(buffer_12_196) + $signed(buffer_12_197); // @[Modules.scala 160:64:@41133.4]
  assign _T_93508 = _T_93507[13:0]; // @[Modules.scala 160:64:@41134.4]
  assign buffer_12_396 = $signed(_T_93508); // @[Modules.scala 160:64:@41135.4]
  assign _T_93510 = $signed(buffer_1_205) + $signed(buffer_8_211); // @[Modules.scala 160:64:@41137.4]
  assign _T_93511 = _T_93510[13:0]; // @[Modules.scala 160:64:@41138.4]
  assign buffer_12_397 = $signed(_T_93511); // @[Modules.scala 160:64:@41139.4]
  assign _T_93516 = $signed(buffer_5_213) + $signed(buffer_11_208); // @[Modules.scala 160:64:@41145.4]
  assign _T_93517 = _T_93516[13:0]; // @[Modules.scala 160:64:@41146.4]
  assign buffer_12_399 = $signed(_T_93517); // @[Modules.scala 160:64:@41147.4]
  assign _T_93519 = $signed(buffer_1_211) + $signed(buffer_1_212); // @[Modules.scala 160:64:@41149.4]
  assign _T_93520 = _T_93519[13:0]; // @[Modules.scala 160:64:@41150.4]
  assign buffer_12_400 = $signed(_T_93520); // @[Modules.scala 160:64:@41151.4]
  assign buffer_12_206 = {{8{_T_92575[5]}},_T_92575}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_207 = {{8{_T_92582[5]}},_T_92582}; // @[Modules.scala 112:22:@8.4]
  assign _T_93522 = $signed(buffer_12_206) + $signed(buffer_12_207); // @[Modules.scala 160:64:@41153.4]
  assign _T_93523 = _T_93522[13:0]; // @[Modules.scala 160:64:@41154.4]
  assign buffer_12_401 = $signed(_T_93523); // @[Modules.scala 160:64:@41155.4]
  assign buffer_12_208 = {{8{_T_92589[5]}},_T_92589}; // @[Modules.scala 112:22:@8.4]
  assign _T_93525 = $signed(buffer_12_208) + $signed(buffer_1_217); // @[Modules.scala 160:64:@41157.4]
  assign _T_93526 = _T_93525[13:0]; // @[Modules.scala 160:64:@41158.4]
  assign buffer_12_402 = $signed(_T_93526); // @[Modules.scala 160:64:@41159.4]
  assign _T_93531 = $signed(buffer_0_219) + $signed(buffer_0_220); // @[Modules.scala 160:64:@41165.4]
  assign _T_93532 = _T_93531[13:0]; // @[Modules.scala 160:64:@41166.4]
  assign buffer_12_404 = $signed(_T_93532); // @[Modules.scala 160:64:@41167.4]
  assign buffer_12_215 = {{8{_T_92638[5]}},_T_92638}; // @[Modules.scala 112:22:@8.4]
  assign _T_93534 = $signed(buffer_8_226) + $signed(buffer_12_215); // @[Modules.scala 160:64:@41169.4]
  assign _T_93535 = _T_93534[13:0]; // @[Modules.scala 160:64:@41170.4]
  assign buffer_12_405 = $signed(_T_93535); // @[Modules.scala 160:64:@41171.4]
  assign buffer_12_216 = {{8{_T_92645[5]}},_T_92645}; // @[Modules.scala 112:22:@8.4]
  assign _T_93537 = $signed(buffer_12_216) + $signed(buffer_5_228); // @[Modules.scala 160:64:@41173.4]
  assign _T_93538 = _T_93537[13:0]; // @[Modules.scala 160:64:@41174.4]
  assign buffer_12_406 = $signed(_T_93538); // @[Modules.scala 160:64:@41175.4]
  assign buffer_12_220 = {{8{_T_92673[5]}},_T_92673}; // @[Modules.scala 112:22:@8.4]
  assign _T_93543 = $signed(buffer_12_220) + $signed(buffer_1_227); // @[Modules.scala 160:64:@41181.4]
  assign _T_93544 = _T_93543[13:0]; // @[Modules.scala 160:64:@41182.4]
  assign buffer_12_408 = $signed(_T_93544); // @[Modules.scala 160:64:@41183.4]
  assign _T_93546 = $signed(buffer_9_237) + $signed(buffer_9_238); // @[Modules.scala 160:64:@41185.4]
  assign _T_93547 = _T_93546[13:0]; // @[Modules.scala 160:64:@41186.4]
  assign buffer_12_409 = $signed(_T_93547); // @[Modules.scala 160:64:@41187.4]
  assign buffer_12_227 = {{8{_T_92722[5]}},_T_92722}; // @[Modules.scala 112:22:@8.4]
  assign _T_93552 = $signed(buffer_0_230) + $signed(buffer_12_227); // @[Modules.scala 160:64:@41193.4]
  assign _T_93553 = _T_93552[13:0]; // @[Modules.scala 160:64:@41194.4]
  assign buffer_12_411 = $signed(_T_93553); // @[Modules.scala 160:64:@41195.4]
  assign buffer_12_228 = {{8{_T_92729[5]}},_T_92729}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_229 = {{8{_T_92736[5]}},_T_92736}; // @[Modules.scala 112:22:@8.4]
  assign _T_93555 = $signed(buffer_12_228) + $signed(buffer_12_229); // @[Modules.scala 160:64:@41197.4]
  assign _T_93556 = _T_93555[13:0]; // @[Modules.scala 160:64:@41198.4]
  assign buffer_12_412 = $signed(_T_93556); // @[Modules.scala 160:64:@41199.4]
  assign buffer_12_230 = {{8{_T_92743[5]}},_T_92743}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_231 = {{8{_T_92750[5]}},_T_92750}; // @[Modules.scala 112:22:@8.4]
  assign _T_93558 = $signed(buffer_12_230) + $signed(buffer_12_231); // @[Modules.scala 160:64:@41201.4]
  assign _T_93559 = _T_93558[13:0]; // @[Modules.scala 160:64:@41202.4]
  assign buffer_12_413 = $signed(_T_93559); // @[Modules.scala 160:64:@41203.4]
  assign buffer_12_238 = {{8{_T_92799[5]}},_T_92799}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_239 = {{8{_T_92806[5]}},_T_92806}; // @[Modules.scala 112:22:@8.4]
  assign _T_93570 = $signed(buffer_12_238) + $signed(buffer_12_239); // @[Modules.scala 160:64:@41217.4]
  assign _T_93571 = _T_93570[13:0]; // @[Modules.scala 160:64:@41218.4]
  assign buffer_12_417 = $signed(_T_93571); // @[Modules.scala 160:64:@41219.4]
  assign buffer_12_240 = {{8{_T_92813[5]}},_T_92813}; // @[Modules.scala 112:22:@8.4]
  assign _T_93573 = $signed(buffer_12_240) + $signed(buffer_0_244); // @[Modules.scala 160:64:@41221.4]
  assign _T_93574 = _T_93573[13:0]; // @[Modules.scala 160:64:@41222.4]
  assign buffer_12_418 = $signed(_T_93574); // @[Modules.scala 160:64:@41223.4]
  assign buffer_12_242 = {{8{_T_92827[5]}},_T_92827}; // @[Modules.scala 112:22:@8.4]
  assign _T_93576 = $signed(buffer_12_242) + $signed(buffer_1_248); // @[Modules.scala 160:64:@41225.4]
  assign _T_93577 = _T_93576[13:0]; // @[Modules.scala 160:64:@41226.4]
  assign buffer_12_419 = $signed(_T_93577); // @[Modules.scala 160:64:@41227.4]
  assign buffer_12_245 = {{8{_T_92848[5]}},_T_92848}; // @[Modules.scala 112:22:@8.4]
  assign _T_93579 = $signed(buffer_3_259) + $signed(buffer_12_245); // @[Modules.scala 160:64:@41229.4]
  assign _T_93580 = _T_93579[13:0]; // @[Modules.scala 160:64:@41230.4]
  assign buffer_12_420 = $signed(_T_93580); // @[Modules.scala 160:64:@41231.4]
  assign _T_93585 = $signed(buffer_9_263) + $signed(buffer_5_262); // @[Modules.scala 160:64:@41237.4]
  assign _T_93586 = _T_93585[13:0]; // @[Modules.scala 160:64:@41238.4]
  assign buffer_12_422 = $signed(_T_93586); // @[Modules.scala 160:64:@41239.4]
  assign buffer_12_251 = {{8{_T_92890[5]}},_T_92890}; // @[Modules.scala 112:22:@8.4]
  assign _T_93588 = $signed(buffer_3_263) + $signed(buffer_12_251); // @[Modules.scala 160:64:@41241.4]
  assign _T_93589 = _T_93588[13:0]; // @[Modules.scala 160:64:@41242.4]
  assign buffer_12_423 = $signed(_T_93589); // @[Modules.scala 160:64:@41243.4]
  assign buffer_12_253 = {{8{_T_92904[5]}},_T_92904}; // @[Modules.scala 112:22:@8.4]
  assign _T_93591 = $signed(buffer_4_252) + $signed(buffer_12_253); // @[Modules.scala 160:64:@41245.4]
  assign _T_93592 = _T_93591[13:0]; // @[Modules.scala 160:64:@41246.4]
  assign buffer_12_424 = $signed(_T_93592); // @[Modules.scala 160:64:@41247.4]
  assign buffer_12_254 = {{9{_T_92911[4]}},_T_92911}; // @[Modules.scala 112:22:@8.4]
  assign buffer_12_255 = {{9{_T_92918[4]}},_T_92918}; // @[Modules.scala 112:22:@8.4]
  assign _T_93594 = $signed(buffer_12_254) + $signed(buffer_12_255); // @[Modules.scala 160:64:@41249.4]
  assign _T_93595 = _T_93594[13:0]; // @[Modules.scala 160:64:@41250.4]
  assign buffer_12_425 = $signed(_T_93595); // @[Modules.scala 160:64:@41251.4]
  assign buffer_12_256 = {{8{_T_92925[5]}},_T_92925}; // @[Modules.scala 112:22:@8.4]
  assign _T_93597 = $signed(buffer_12_256) + $signed(buffer_5_270); // @[Modules.scala 160:64:@41253.4]
  assign _T_93598 = _T_93597[13:0]; // @[Modules.scala 160:64:@41254.4]
  assign buffer_12_426 = $signed(_T_93598); // @[Modules.scala 160:64:@41255.4]
  assign buffer_12_261 = {{8{_T_92960[5]}},_T_92960}; // @[Modules.scala 112:22:@8.4]
  assign _T_93603 = $signed(buffer_2_272) + $signed(buffer_12_261); // @[Modules.scala 160:64:@41261.4]
  assign _T_93604 = _T_93603[13:0]; // @[Modules.scala 160:64:@41262.4]
  assign buffer_12_428 = $signed(_T_93604); // @[Modules.scala 160:64:@41263.4]
  assign buffer_12_263 = {{8{_T_92974[5]}},_T_92974}; // @[Modules.scala 112:22:@8.4]
  assign _T_93606 = $signed(buffer_7_273) + $signed(buffer_12_263); // @[Modules.scala 160:64:@41265.4]
  assign _T_93607 = _T_93606[13:0]; // @[Modules.scala 160:64:@41266.4]
  assign buffer_12_429 = $signed(_T_93607); // @[Modules.scala 160:64:@41267.4]
  assign _T_93609 = $signed(buffer_9_278) + $signed(buffer_3_279); // @[Modules.scala 160:64:@41269.4]
  assign _T_93610 = _T_93609[13:0]; // @[Modules.scala 160:64:@41270.4]
  assign buffer_12_430 = $signed(_T_93610); // @[Modules.scala 160:64:@41271.4]
  assign buffer_12_266 = {{8{_T_92995[5]}},_T_92995}; // @[Modules.scala 112:22:@8.4]
  assign _T_93612 = $signed(buffer_12_266) + $signed(buffer_7_278); // @[Modules.scala 160:64:@41273.4]
  assign _T_93613 = _T_93612[13:0]; // @[Modules.scala 160:64:@41274.4]
  assign buffer_12_431 = $signed(_T_93613); // @[Modules.scala 160:64:@41275.4]
  assign buffer_12_268 = {{8{_T_93009[5]}},_T_93009}; // @[Modules.scala 112:22:@8.4]
  assign _T_93615 = $signed(buffer_12_268) + $signed(buffer_7_281); // @[Modules.scala 160:64:@41277.4]
  assign _T_93616 = _T_93615[13:0]; // @[Modules.scala 160:64:@41278.4]
  assign buffer_12_432 = $signed(_T_93616); // @[Modules.scala 160:64:@41279.4]
  assign buffer_12_273 = {{8{_T_93044[5]}},_T_93044}; // @[Modules.scala 112:22:@8.4]
  assign _T_93621 = $signed(buffer_0_277) + $signed(buffer_12_273); // @[Modules.scala 160:64:@41285.4]
  assign _T_93622 = _T_93621[13:0]; // @[Modules.scala 160:64:@41286.4]
  assign buffer_12_434 = $signed(_T_93622); // @[Modules.scala 160:64:@41287.4]
  assign _T_93624 = $signed(buffer_2_285) + $signed(buffer_6_291); // @[Modules.scala 160:64:@41289.4]
  assign _T_93625 = _T_93624[13:0]; // @[Modules.scala 160:64:@41290.4]
  assign buffer_12_435 = $signed(_T_93625); // @[Modules.scala 160:64:@41291.4]
  assign buffer_12_276 = {{8{_T_93065[5]}},_T_93065}; // @[Modules.scala 112:22:@8.4]
  assign _T_93627 = $signed(buffer_12_276) + $signed(buffer_3_291); // @[Modules.scala 160:64:@41293.4]
  assign _T_93628 = _T_93627[13:0]; // @[Modules.scala 160:64:@41294.4]
  assign buffer_12_436 = $signed(_T_93628); // @[Modules.scala 160:64:@41295.4]
  assign buffer_12_278 = {{9{_T_93079[4]}},_T_93079}; // @[Modules.scala 112:22:@8.4]
  assign _T_93630 = $signed(buffer_12_278) + $signed(buffer_1_283); // @[Modules.scala 160:64:@41297.4]
  assign _T_93631 = _T_93630[13:0]; // @[Modules.scala 160:64:@41298.4]
  assign buffer_12_437 = $signed(_T_93631); // @[Modules.scala 160:64:@41299.4]
  assign buffer_12_280 = {{8{_T_93093[5]}},_T_93093}; // @[Modules.scala 112:22:@8.4]
  assign _T_93633 = $signed(buffer_12_280) + $signed(buffer_9_297); // @[Modules.scala 160:64:@41301.4]
  assign _T_93634 = _T_93633[13:0]; // @[Modules.scala 160:64:@41302.4]
  assign buffer_12_438 = $signed(_T_93634); // @[Modules.scala 160:64:@41303.4]
  assign buffer_12_289 = {{9{_T_93156[4]}},_T_93156}; // @[Modules.scala 112:22:@8.4]
  assign _T_93645 = $signed(buffer_5_304) + $signed(buffer_12_289); // @[Modules.scala 160:64:@41317.4]
  assign _T_93646 = _T_93645[13:0]; // @[Modules.scala 160:64:@41318.4]
  assign buffer_12_442 = $signed(_T_93646); // @[Modules.scala 160:64:@41319.4]
  assign _T_93648 = $signed(buffer_0_294) + $signed(buffer_2_304); // @[Modules.scala 160:64:@41321.4]
  assign _T_93649 = _T_93648[13:0]; // @[Modules.scala 160:64:@41322.4]
  assign buffer_12_443 = $signed(_T_93649); // @[Modules.scala 160:64:@41323.4]
  assign buffer_12_296 = {{8{_T_93205[5]}},_T_93205}; // @[Modules.scala 112:22:@8.4]
  assign _T_93657 = $signed(buffer_12_296) + $signed(buffer_7_308); // @[Modules.scala 160:64:@41333.4]
  assign _T_93658 = _T_93657[13:0]; // @[Modules.scala 160:64:@41334.4]
  assign buffer_12_446 = $signed(_T_93658); // @[Modules.scala 160:64:@41335.4]
  assign _T_93660 = $signed(buffer_12_298) + $signed(buffer_11_300); // @[Modules.scala 166:64:@41337.4]
  assign _T_93661 = _T_93660[13:0]; // @[Modules.scala 166:64:@41338.4]
  assign buffer_12_447 = $signed(_T_93661); // @[Modules.scala 166:64:@41339.4]
  assign _T_93663 = $signed(buffer_12_300) + $signed(buffer_0_305); // @[Modules.scala 166:64:@41341.4]
  assign _T_93664 = _T_93663[13:0]; // @[Modules.scala 166:64:@41342.4]
  assign buffer_12_448 = $signed(_T_93664); // @[Modules.scala 166:64:@41343.4]
  assign _T_93666 = $signed(buffer_12_302) + $signed(buffer_12_303); // @[Modules.scala 166:64:@41345.4]
  assign _T_93667 = _T_93666[13:0]; // @[Modules.scala 166:64:@41346.4]
  assign buffer_12_449 = $signed(_T_93667); // @[Modules.scala 166:64:@41347.4]
  assign _T_93669 = $signed(buffer_12_304) + $signed(buffer_12_305); // @[Modules.scala 166:64:@41349.4]
  assign _T_93670 = _T_93669[13:0]; // @[Modules.scala 166:64:@41350.4]
  assign buffer_12_450 = $signed(_T_93670); // @[Modules.scala 166:64:@41351.4]
  assign _T_93672 = $signed(buffer_12_306) + $signed(buffer_12_307); // @[Modules.scala 166:64:@41353.4]
  assign _T_93673 = _T_93672[13:0]; // @[Modules.scala 166:64:@41354.4]
  assign buffer_12_451 = $signed(_T_93673); // @[Modules.scala 166:64:@41355.4]
  assign _T_93675 = $signed(buffer_12_308) + $signed(buffer_3_326); // @[Modules.scala 166:64:@41357.4]
  assign _T_93676 = _T_93675[13:0]; // @[Modules.scala 166:64:@41358.4]
  assign buffer_12_452 = $signed(_T_93676); // @[Modules.scala 166:64:@41359.4]
  assign _T_93678 = $signed(buffer_3_327) + $signed(buffer_12_311); // @[Modules.scala 166:64:@41361.4]
  assign _T_93679 = _T_93678[13:0]; // @[Modules.scala 166:64:@41362.4]
  assign buffer_12_453 = $signed(_T_93679); // @[Modules.scala 166:64:@41363.4]
  assign _T_93681 = $signed(buffer_12_312) + $signed(buffer_12_313); // @[Modules.scala 166:64:@41365.4]
  assign _T_93682 = _T_93681[13:0]; // @[Modules.scala 166:64:@41366.4]
  assign buffer_12_454 = $signed(_T_93682); // @[Modules.scala 166:64:@41367.4]
  assign _T_93684 = $signed(buffer_12_314) + $signed(buffer_12_315); // @[Modules.scala 166:64:@41369.4]
  assign _T_93685 = _T_93684[13:0]; // @[Modules.scala 166:64:@41370.4]
  assign buffer_12_455 = $signed(_T_93685); // @[Modules.scala 166:64:@41371.4]
  assign _T_93687 = $signed(buffer_12_316) + $signed(buffer_12_317); // @[Modules.scala 166:64:@41373.4]
  assign _T_93688 = _T_93687[13:0]; // @[Modules.scala 166:64:@41374.4]
  assign buffer_12_456 = $signed(_T_93688); // @[Modules.scala 166:64:@41375.4]
  assign _T_93690 = $signed(buffer_12_318) + $signed(buffer_12_319); // @[Modules.scala 166:64:@41377.4]
  assign _T_93691 = _T_93690[13:0]; // @[Modules.scala 166:64:@41378.4]
  assign buffer_12_457 = $signed(_T_93691); // @[Modules.scala 166:64:@41379.4]
  assign _T_93693 = $signed(buffer_12_320) + $signed(buffer_12_321); // @[Modules.scala 166:64:@41381.4]
  assign _T_93694 = _T_93693[13:0]; // @[Modules.scala 166:64:@41382.4]
  assign buffer_12_458 = $signed(_T_93694); // @[Modules.scala 166:64:@41383.4]
  assign _T_93696 = $signed(buffer_12_322) + $signed(buffer_12_323); // @[Modules.scala 166:64:@41385.4]
  assign _T_93697 = _T_93696[13:0]; // @[Modules.scala 166:64:@41386.4]
  assign buffer_12_459 = $signed(_T_93697); // @[Modules.scala 166:64:@41387.4]
  assign _T_93699 = $signed(buffer_12_324) + $signed(buffer_12_325); // @[Modules.scala 166:64:@41389.4]
  assign _T_93700 = _T_93699[13:0]; // @[Modules.scala 166:64:@41390.4]
  assign buffer_12_460 = $signed(_T_93700); // @[Modules.scala 166:64:@41391.4]
  assign _T_93702 = $signed(buffer_12_326) + $signed(buffer_12_327); // @[Modules.scala 166:64:@41393.4]
  assign _T_93703 = _T_93702[13:0]; // @[Modules.scala 166:64:@41394.4]
  assign buffer_12_461 = $signed(_T_93703); // @[Modules.scala 166:64:@41395.4]
  assign _T_93705 = $signed(buffer_12_328) + $signed(buffer_12_329); // @[Modules.scala 166:64:@41397.4]
  assign _T_93706 = _T_93705[13:0]; // @[Modules.scala 166:64:@41398.4]
  assign buffer_12_462 = $signed(_T_93706); // @[Modules.scala 166:64:@41399.4]
  assign _T_93708 = $signed(buffer_12_330) + $signed(buffer_12_331); // @[Modules.scala 166:64:@41401.4]
  assign _T_93709 = _T_93708[13:0]; // @[Modules.scala 166:64:@41402.4]
  assign buffer_12_463 = $signed(_T_93709); // @[Modules.scala 166:64:@41403.4]
  assign _T_93711 = $signed(buffer_7_347) + $signed(buffer_12_333); // @[Modules.scala 166:64:@41405.4]
  assign _T_93712 = _T_93711[13:0]; // @[Modules.scala 166:64:@41406.4]
  assign buffer_12_464 = $signed(_T_93712); // @[Modules.scala 166:64:@41407.4]
  assign _T_93714 = $signed(buffer_12_334) + $signed(buffer_12_335); // @[Modules.scala 166:64:@41409.4]
  assign _T_93715 = _T_93714[13:0]; // @[Modules.scala 166:64:@41410.4]
  assign buffer_12_465 = $signed(_T_93715); // @[Modules.scala 166:64:@41411.4]
  assign _T_93717 = $signed(buffer_12_336) + $signed(buffer_8_351); // @[Modules.scala 166:64:@41413.4]
  assign _T_93718 = _T_93717[13:0]; // @[Modules.scala 166:64:@41414.4]
  assign buffer_12_466 = $signed(_T_93718); // @[Modules.scala 166:64:@41415.4]
  assign _T_93720 = $signed(buffer_12_338) + $signed(buffer_12_339); // @[Modules.scala 166:64:@41417.4]
  assign _T_93721 = _T_93720[13:0]; // @[Modules.scala 166:64:@41418.4]
  assign buffer_12_467 = $signed(_T_93721); // @[Modules.scala 166:64:@41419.4]
  assign _T_93723 = $signed(buffer_12_340) + $signed(buffer_12_341); // @[Modules.scala 166:64:@41421.4]
  assign _T_93724 = _T_93723[13:0]; // @[Modules.scala 166:64:@41422.4]
  assign buffer_12_468 = $signed(_T_93724); // @[Modules.scala 166:64:@41423.4]
  assign _T_93726 = $signed(buffer_12_342) + $signed(buffer_12_343); // @[Modules.scala 166:64:@41425.4]
  assign _T_93727 = _T_93726[13:0]; // @[Modules.scala 166:64:@41426.4]
  assign buffer_12_469 = $signed(_T_93727); // @[Modules.scala 166:64:@41427.4]
  assign _T_93729 = $signed(buffer_12_344) + $signed(buffer_12_345); // @[Modules.scala 166:64:@41429.4]
  assign _T_93730 = _T_93729[13:0]; // @[Modules.scala 166:64:@41430.4]
  assign buffer_12_470 = $signed(_T_93730); // @[Modules.scala 166:64:@41431.4]
  assign _T_93732 = $signed(buffer_12_346) + $signed(buffer_0_356); // @[Modules.scala 166:64:@41433.4]
  assign _T_93733 = _T_93732[13:0]; // @[Modules.scala 166:64:@41434.4]
  assign buffer_12_471 = $signed(_T_93733); // @[Modules.scala 166:64:@41435.4]
  assign _T_93738 = $signed(buffer_12_350) + $signed(buffer_12_351); // @[Modules.scala 166:64:@41441.4]
  assign _T_93739 = _T_93738[13:0]; // @[Modules.scala 166:64:@41442.4]
  assign buffer_12_473 = $signed(_T_93739); // @[Modules.scala 166:64:@41443.4]
  assign _T_93741 = $signed(buffer_12_352) + $signed(buffer_9_378); // @[Modules.scala 166:64:@41445.4]
  assign _T_93742 = _T_93741[13:0]; // @[Modules.scala 166:64:@41446.4]
  assign buffer_12_474 = $signed(_T_93742); // @[Modules.scala 166:64:@41447.4]
  assign _T_93744 = $signed(buffer_9_379) + $signed(buffer_10_371); // @[Modules.scala 166:64:@41449.4]
  assign _T_93745 = _T_93744[13:0]; // @[Modules.scala 166:64:@41450.4]
  assign buffer_12_475 = $signed(_T_93745); // @[Modules.scala 166:64:@41451.4]
  assign _T_93747 = $signed(buffer_12_356) + $signed(buffer_12_357); // @[Modules.scala 166:64:@41453.4]
  assign _T_93748 = _T_93747[13:0]; // @[Modules.scala 166:64:@41454.4]
  assign buffer_12_476 = $signed(_T_93748); // @[Modules.scala 166:64:@41455.4]
  assign _T_93750 = $signed(buffer_8_374) + $signed(buffer_12_359); // @[Modules.scala 166:64:@41457.4]
  assign _T_93751 = _T_93750[13:0]; // @[Modules.scala 166:64:@41458.4]
  assign buffer_12_477 = $signed(_T_93751); // @[Modules.scala 166:64:@41459.4]
  assign _T_93753 = $signed(buffer_12_360) + $signed(buffer_12_361); // @[Modules.scala 166:64:@41461.4]
  assign _T_93754 = _T_93753[13:0]; // @[Modules.scala 166:64:@41462.4]
  assign buffer_12_478 = $signed(_T_93754); // @[Modules.scala 166:64:@41463.4]
  assign _T_93756 = $signed(buffer_12_362) + $signed(buffer_12_363); // @[Modules.scala 166:64:@41465.4]
  assign _T_93757 = _T_93756[13:0]; // @[Modules.scala 166:64:@41466.4]
  assign buffer_12_479 = $signed(_T_93757); // @[Modules.scala 166:64:@41467.4]
  assign _T_93759 = $signed(buffer_8_380) + $signed(buffer_12_365); // @[Modules.scala 166:64:@41469.4]
  assign _T_93760 = _T_93759[13:0]; // @[Modules.scala 166:64:@41470.4]
  assign buffer_12_480 = $signed(_T_93760); // @[Modules.scala 166:64:@41471.4]
  assign _T_93762 = $signed(buffer_12_366) + $signed(buffer_12_367); // @[Modules.scala 166:64:@41473.4]
  assign _T_93763 = _T_93762[13:0]; // @[Modules.scala 166:64:@41474.4]
  assign buffer_12_481 = $signed(_T_93763); // @[Modules.scala 166:64:@41475.4]
  assign _T_93765 = $signed(buffer_7_385) + $signed(buffer_12_369); // @[Modules.scala 166:64:@41477.4]
  assign _T_93766 = _T_93765[13:0]; // @[Modules.scala 166:64:@41478.4]
  assign buffer_12_482 = $signed(_T_93766); // @[Modules.scala 166:64:@41479.4]
  assign _T_93768 = $signed(buffer_12_370) + $signed(buffer_12_371); // @[Modules.scala 166:64:@41481.4]
  assign _T_93769 = _T_93768[13:0]; // @[Modules.scala 166:64:@41482.4]
  assign buffer_12_483 = $signed(_T_93769); // @[Modules.scala 166:64:@41483.4]
  assign _T_93771 = $signed(buffer_12_372) + $signed(buffer_12_373); // @[Modules.scala 166:64:@41485.4]
  assign _T_93772 = _T_93771[13:0]; // @[Modules.scala 166:64:@41486.4]
  assign buffer_12_484 = $signed(_T_93772); // @[Modules.scala 166:64:@41487.4]
  assign _T_93774 = $signed(buffer_12_374) + $signed(buffer_12_375); // @[Modules.scala 166:64:@41489.4]
  assign _T_93775 = _T_93774[13:0]; // @[Modules.scala 166:64:@41490.4]
  assign buffer_12_485 = $signed(_T_93775); // @[Modules.scala 166:64:@41491.4]
  assign _T_93777 = $signed(buffer_11_380) + $signed(buffer_12_377); // @[Modules.scala 166:64:@41493.4]
  assign _T_93778 = _T_93777[13:0]; // @[Modules.scala 166:64:@41494.4]
  assign buffer_12_486 = $signed(_T_93778); // @[Modules.scala 166:64:@41495.4]
  assign _T_93780 = $signed(buffer_12_378) + $signed(buffer_12_379); // @[Modules.scala 166:64:@41497.4]
  assign _T_93781 = _T_93780[13:0]; // @[Modules.scala 166:64:@41498.4]
  assign buffer_12_487 = $signed(_T_93781); // @[Modules.scala 166:64:@41499.4]
  assign _T_93783 = $signed(buffer_12_380) + $signed(buffer_12_381); // @[Modules.scala 166:64:@41501.4]
  assign _T_93784 = _T_93783[13:0]; // @[Modules.scala 166:64:@41502.4]
  assign buffer_12_488 = $signed(_T_93784); // @[Modules.scala 166:64:@41503.4]
  assign _T_93786 = $signed(buffer_12_382) + $signed(buffer_12_383); // @[Modules.scala 166:64:@41505.4]
  assign _T_93787 = _T_93786[13:0]; // @[Modules.scala 166:64:@41506.4]
  assign buffer_12_489 = $signed(_T_93787); // @[Modules.scala 166:64:@41507.4]
  assign _T_93789 = $signed(buffer_12_384) + $signed(buffer_12_385); // @[Modules.scala 166:64:@41509.4]
  assign _T_93790 = _T_93789[13:0]; // @[Modules.scala 166:64:@41510.4]
  assign buffer_12_490 = $signed(_T_93790); // @[Modules.scala 166:64:@41511.4]
  assign _T_93792 = $signed(buffer_12_386) + $signed(buffer_12_387); // @[Modules.scala 166:64:@41513.4]
  assign _T_93793 = _T_93792[13:0]; // @[Modules.scala 166:64:@41514.4]
  assign buffer_12_491 = $signed(_T_93793); // @[Modules.scala 166:64:@41515.4]
  assign _T_93795 = $signed(buffer_12_388) + $signed(buffer_12_389); // @[Modules.scala 166:64:@41517.4]
  assign _T_93796 = _T_93795[13:0]; // @[Modules.scala 166:64:@41518.4]
  assign buffer_12_492 = $signed(_T_93796); // @[Modules.scala 166:64:@41519.4]
  assign _T_93798 = $signed(buffer_12_390) + $signed(buffer_12_391); // @[Modules.scala 166:64:@41521.4]
  assign _T_93799 = _T_93798[13:0]; // @[Modules.scala 166:64:@41522.4]
  assign buffer_12_493 = $signed(_T_93799); // @[Modules.scala 166:64:@41523.4]
  assign _T_93801 = $signed(buffer_12_392) + $signed(buffer_12_393); // @[Modules.scala 166:64:@41525.4]
  assign _T_93802 = _T_93801[13:0]; // @[Modules.scala 166:64:@41526.4]
  assign buffer_12_494 = $signed(_T_93802); // @[Modules.scala 166:64:@41527.4]
  assign _T_93804 = $signed(buffer_4_396) + $signed(buffer_12_395); // @[Modules.scala 166:64:@41529.4]
  assign _T_93805 = _T_93804[13:0]; // @[Modules.scala 166:64:@41530.4]
  assign buffer_12_495 = $signed(_T_93805); // @[Modules.scala 166:64:@41531.4]
  assign _T_93807 = $signed(buffer_12_396) + $signed(buffer_12_397); // @[Modules.scala 166:64:@41533.4]
  assign _T_93808 = _T_93807[13:0]; // @[Modules.scala 166:64:@41534.4]
  assign buffer_12_496 = $signed(_T_93808); // @[Modules.scala 166:64:@41535.4]
  assign _T_93810 = $signed(buffer_0_406) + $signed(buffer_12_399); // @[Modules.scala 166:64:@41537.4]
  assign _T_93811 = _T_93810[13:0]; // @[Modules.scala 166:64:@41538.4]
  assign buffer_12_497 = $signed(_T_93811); // @[Modules.scala 166:64:@41539.4]
  assign _T_93813 = $signed(buffer_12_400) + $signed(buffer_12_401); // @[Modules.scala 166:64:@41541.4]
  assign _T_93814 = _T_93813[13:0]; // @[Modules.scala 166:64:@41542.4]
  assign buffer_12_498 = $signed(_T_93814); // @[Modules.scala 166:64:@41543.4]
  assign _T_93816 = $signed(buffer_12_402) + $signed(buffer_2_421); // @[Modules.scala 166:64:@41545.4]
  assign _T_93817 = _T_93816[13:0]; // @[Modules.scala 166:64:@41546.4]
  assign buffer_12_499 = $signed(_T_93817); // @[Modules.scala 166:64:@41547.4]
  assign _T_93819 = $signed(buffer_12_404) + $signed(buffer_12_405); // @[Modules.scala 166:64:@41549.4]
  assign _T_93820 = _T_93819[13:0]; // @[Modules.scala 166:64:@41550.4]
  assign buffer_12_500 = $signed(_T_93820); // @[Modules.scala 166:64:@41551.4]
  assign _T_93822 = $signed(buffer_12_406) + $signed(buffer_6_434); // @[Modules.scala 166:64:@41553.4]
  assign _T_93823 = _T_93822[13:0]; // @[Modules.scala 166:64:@41554.4]
  assign buffer_12_501 = $signed(_T_93823); // @[Modules.scala 166:64:@41555.4]
  assign _T_93825 = $signed(buffer_12_408) + $signed(buffer_12_409); // @[Modules.scala 166:64:@41557.4]
  assign _T_93826 = _T_93825[13:0]; // @[Modules.scala 166:64:@41558.4]
  assign buffer_12_502 = $signed(_T_93826); // @[Modules.scala 166:64:@41559.4]
  assign _T_93828 = $signed(buffer_0_416) + $signed(buffer_12_411); // @[Modules.scala 166:64:@41561.4]
  assign _T_93829 = _T_93828[13:0]; // @[Modules.scala 166:64:@41562.4]
  assign buffer_12_503 = $signed(_T_93829); // @[Modules.scala 166:64:@41563.4]
  assign _T_93831 = $signed(buffer_12_412) + $signed(buffer_12_413); // @[Modules.scala 166:64:@41565.4]
  assign _T_93832 = _T_93831[13:0]; // @[Modules.scala 166:64:@41566.4]
  assign buffer_12_504 = $signed(_T_93832); // @[Modules.scala 166:64:@41567.4]
  assign _T_93837 = $signed(buffer_1_424) + $signed(buffer_12_417); // @[Modules.scala 166:64:@41573.4]
  assign _T_93838 = _T_93837[13:0]; // @[Modules.scala 166:64:@41574.4]
  assign buffer_12_506 = $signed(_T_93838); // @[Modules.scala 166:64:@41575.4]
  assign _T_93840 = $signed(buffer_12_418) + $signed(buffer_12_419); // @[Modules.scala 166:64:@41577.4]
  assign _T_93841 = _T_93840[13:0]; // @[Modules.scala 166:64:@41578.4]
  assign buffer_12_507 = $signed(_T_93841); // @[Modules.scala 166:64:@41579.4]
  assign _T_93843 = $signed(buffer_12_420) + $signed(buffer_6_447); // @[Modules.scala 166:64:@41581.4]
  assign _T_93844 = _T_93843[13:0]; // @[Modules.scala 166:64:@41582.4]
  assign buffer_12_508 = $signed(_T_93844); // @[Modules.scala 166:64:@41583.4]
  assign _T_93846 = $signed(buffer_12_422) + $signed(buffer_12_423); // @[Modules.scala 166:64:@41585.4]
  assign _T_93847 = _T_93846[13:0]; // @[Modules.scala 166:64:@41586.4]
  assign buffer_12_509 = $signed(_T_93847); // @[Modules.scala 166:64:@41587.4]
  assign _T_93849 = $signed(buffer_12_424) + $signed(buffer_12_425); // @[Modules.scala 166:64:@41589.4]
  assign _T_93850 = _T_93849[13:0]; // @[Modules.scala 166:64:@41590.4]
  assign buffer_12_510 = $signed(_T_93850); // @[Modules.scala 166:64:@41591.4]
  assign _T_93852 = $signed(buffer_12_426) + $signed(buffer_9_450); // @[Modules.scala 166:64:@41593.4]
  assign _T_93853 = _T_93852[13:0]; // @[Modules.scala 166:64:@41594.4]
  assign buffer_12_511 = $signed(_T_93853); // @[Modules.scala 166:64:@41595.4]
  assign _T_93855 = $signed(buffer_12_428) + $signed(buffer_12_429); // @[Modules.scala 166:64:@41597.4]
  assign _T_93856 = _T_93855[13:0]; // @[Modules.scala 166:64:@41598.4]
  assign buffer_12_512 = $signed(_T_93856); // @[Modules.scala 166:64:@41599.4]
  assign _T_93858 = $signed(buffer_12_430) + $signed(buffer_12_431); // @[Modules.scala 166:64:@41601.4]
  assign _T_93859 = _T_93858[13:0]; // @[Modules.scala 166:64:@41602.4]
  assign buffer_12_513 = $signed(_T_93859); // @[Modules.scala 166:64:@41603.4]
  assign _T_93861 = $signed(buffer_12_432) + $signed(buffer_6_459); // @[Modules.scala 166:64:@41605.4]
  assign _T_93862 = _T_93861[13:0]; // @[Modules.scala 166:64:@41606.4]
  assign buffer_12_514 = $signed(_T_93862); // @[Modules.scala 166:64:@41607.4]
  assign _T_93864 = $signed(buffer_12_434) + $signed(buffer_12_435); // @[Modules.scala 166:64:@41609.4]
  assign _T_93865 = _T_93864[13:0]; // @[Modules.scala 166:64:@41610.4]
  assign buffer_12_515 = $signed(_T_93865); // @[Modules.scala 166:64:@41611.4]
  assign _T_93867 = $signed(buffer_12_436) + $signed(buffer_12_437); // @[Modules.scala 166:64:@41613.4]
  assign _T_93868 = _T_93867[13:0]; // @[Modules.scala 166:64:@41614.4]
  assign buffer_12_516 = $signed(_T_93868); // @[Modules.scala 166:64:@41615.4]
  assign _T_93870 = $signed(buffer_12_438) + $signed(buffer_9_463); // @[Modules.scala 166:64:@41617.4]
  assign _T_93871 = _T_93870[13:0]; // @[Modules.scala 166:64:@41618.4]
  assign buffer_12_517 = $signed(_T_93871); // @[Modules.scala 166:64:@41619.4]
  assign _T_93873 = $signed(buffer_9_464) + $signed(buffer_5_465); // @[Modules.scala 166:64:@41621.4]
  assign _T_93874 = _T_93873[13:0]; // @[Modules.scala 166:64:@41622.4]
  assign buffer_12_518 = $signed(_T_93874); // @[Modules.scala 166:64:@41623.4]
  assign _T_93876 = $signed(buffer_12_442) + $signed(buffer_12_443); // @[Modules.scala 166:64:@41625.4]
  assign _T_93877 = _T_93876[13:0]; // @[Modules.scala 166:64:@41626.4]
  assign buffer_12_519 = $signed(_T_93877); // @[Modules.scala 166:64:@41627.4]
  assign _T_93882 = $signed(buffer_12_447) + $signed(buffer_12_448); // @[Modules.scala 160:64:@41633.4]
  assign _T_93883 = _T_93882[13:0]; // @[Modules.scala 160:64:@41634.4]
  assign buffer_12_521 = $signed(_T_93883); // @[Modules.scala 160:64:@41635.4]
  assign _T_93885 = $signed(buffer_12_449) + $signed(buffer_12_450); // @[Modules.scala 160:64:@41637.4]
  assign _T_93886 = _T_93885[13:0]; // @[Modules.scala 160:64:@41638.4]
  assign buffer_12_522 = $signed(_T_93886); // @[Modules.scala 160:64:@41639.4]
  assign _T_93888 = $signed(buffer_12_451) + $signed(buffer_12_452); // @[Modules.scala 160:64:@41641.4]
  assign _T_93889 = _T_93888[13:0]; // @[Modules.scala 160:64:@41642.4]
  assign buffer_12_523 = $signed(_T_93889); // @[Modules.scala 160:64:@41643.4]
  assign _T_93891 = $signed(buffer_12_453) + $signed(buffer_12_454); // @[Modules.scala 160:64:@41645.4]
  assign _T_93892 = _T_93891[13:0]; // @[Modules.scala 160:64:@41646.4]
  assign buffer_12_524 = $signed(_T_93892); // @[Modules.scala 160:64:@41647.4]
  assign _T_93894 = $signed(buffer_12_455) + $signed(buffer_12_456); // @[Modules.scala 160:64:@41649.4]
  assign _T_93895 = _T_93894[13:0]; // @[Modules.scala 160:64:@41650.4]
  assign buffer_12_525 = $signed(_T_93895); // @[Modules.scala 160:64:@41651.4]
  assign _T_93897 = $signed(buffer_12_457) + $signed(buffer_12_458); // @[Modules.scala 160:64:@41653.4]
  assign _T_93898 = _T_93897[13:0]; // @[Modules.scala 160:64:@41654.4]
  assign buffer_12_526 = $signed(_T_93898); // @[Modules.scala 160:64:@41655.4]
  assign _T_93900 = $signed(buffer_12_459) + $signed(buffer_12_460); // @[Modules.scala 160:64:@41657.4]
  assign _T_93901 = _T_93900[13:0]; // @[Modules.scala 160:64:@41658.4]
  assign buffer_12_527 = $signed(_T_93901); // @[Modules.scala 160:64:@41659.4]
  assign _T_93903 = $signed(buffer_12_461) + $signed(buffer_12_462); // @[Modules.scala 160:64:@41661.4]
  assign _T_93904 = _T_93903[13:0]; // @[Modules.scala 160:64:@41662.4]
  assign buffer_12_528 = $signed(_T_93904); // @[Modules.scala 160:64:@41663.4]
  assign _T_93906 = $signed(buffer_12_463) + $signed(buffer_12_464); // @[Modules.scala 160:64:@41665.4]
  assign _T_93907 = _T_93906[13:0]; // @[Modules.scala 160:64:@41666.4]
  assign buffer_12_529 = $signed(_T_93907); // @[Modules.scala 160:64:@41667.4]
  assign _T_93909 = $signed(buffer_12_465) + $signed(buffer_12_466); // @[Modules.scala 160:64:@41669.4]
  assign _T_93910 = _T_93909[13:0]; // @[Modules.scala 160:64:@41670.4]
  assign buffer_12_530 = $signed(_T_93910); // @[Modules.scala 160:64:@41671.4]
  assign _T_93912 = $signed(buffer_12_467) + $signed(buffer_12_468); // @[Modules.scala 160:64:@41673.4]
  assign _T_93913 = _T_93912[13:0]; // @[Modules.scala 160:64:@41674.4]
  assign buffer_12_531 = $signed(_T_93913); // @[Modules.scala 160:64:@41675.4]
  assign _T_93915 = $signed(buffer_12_469) + $signed(buffer_12_470); // @[Modules.scala 160:64:@41677.4]
  assign _T_93916 = _T_93915[13:0]; // @[Modules.scala 160:64:@41678.4]
  assign buffer_12_532 = $signed(_T_93916); // @[Modules.scala 160:64:@41679.4]
  assign _T_93918 = $signed(buffer_12_471) + $signed(buffer_3_500); // @[Modules.scala 160:64:@41681.4]
  assign _T_93919 = _T_93918[13:0]; // @[Modules.scala 160:64:@41682.4]
  assign buffer_12_533 = $signed(_T_93919); // @[Modules.scala 160:64:@41683.4]
  assign _T_93921 = $signed(buffer_12_473) + $signed(buffer_12_474); // @[Modules.scala 160:64:@41685.4]
  assign _T_93922 = _T_93921[13:0]; // @[Modules.scala 160:64:@41686.4]
  assign buffer_12_534 = $signed(_T_93922); // @[Modules.scala 160:64:@41687.4]
  assign _T_93924 = $signed(buffer_12_475) + $signed(buffer_12_476); // @[Modules.scala 160:64:@41689.4]
  assign _T_93925 = _T_93924[13:0]; // @[Modules.scala 160:64:@41690.4]
  assign buffer_12_535 = $signed(_T_93925); // @[Modules.scala 160:64:@41691.4]
  assign _T_93927 = $signed(buffer_12_477) + $signed(buffer_12_478); // @[Modules.scala 160:64:@41693.4]
  assign _T_93928 = _T_93927[13:0]; // @[Modules.scala 160:64:@41694.4]
  assign buffer_12_536 = $signed(_T_93928); // @[Modules.scala 160:64:@41695.4]
  assign _T_93930 = $signed(buffer_12_479) + $signed(buffer_12_480); // @[Modules.scala 160:64:@41697.4]
  assign _T_93931 = _T_93930[13:0]; // @[Modules.scala 160:64:@41698.4]
  assign buffer_12_537 = $signed(_T_93931); // @[Modules.scala 160:64:@41699.4]
  assign _T_93933 = $signed(buffer_12_481) + $signed(buffer_12_482); // @[Modules.scala 160:64:@41701.4]
  assign _T_93934 = _T_93933[13:0]; // @[Modules.scala 160:64:@41702.4]
  assign buffer_12_538 = $signed(_T_93934); // @[Modules.scala 160:64:@41703.4]
  assign _T_93936 = $signed(buffer_12_483) + $signed(buffer_12_484); // @[Modules.scala 160:64:@41705.4]
  assign _T_93937 = _T_93936[13:0]; // @[Modules.scala 160:64:@41706.4]
  assign buffer_12_539 = $signed(_T_93937); // @[Modules.scala 160:64:@41707.4]
  assign _T_93939 = $signed(buffer_12_485) + $signed(buffer_12_486); // @[Modules.scala 160:64:@41709.4]
  assign _T_93940 = _T_93939[13:0]; // @[Modules.scala 160:64:@41710.4]
  assign buffer_12_540 = $signed(_T_93940); // @[Modules.scala 160:64:@41711.4]
  assign _T_93942 = $signed(buffer_12_487) + $signed(buffer_12_488); // @[Modules.scala 160:64:@41713.4]
  assign _T_93943 = _T_93942[13:0]; // @[Modules.scala 160:64:@41714.4]
  assign buffer_12_541 = $signed(_T_93943); // @[Modules.scala 160:64:@41715.4]
  assign _T_93945 = $signed(buffer_12_489) + $signed(buffer_12_490); // @[Modules.scala 160:64:@41717.4]
  assign _T_93946 = _T_93945[13:0]; // @[Modules.scala 160:64:@41718.4]
  assign buffer_12_542 = $signed(_T_93946); // @[Modules.scala 160:64:@41719.4]
  assign _T_93948 = $signed(buffer_12_491) + $signed(buffer_12_492); // @[Modules.scala 160:64:@41721.4]
  assign _T_93949 = _T_93948[13:0]; // @[Modules.scala 160:64:@41722.4]
  assign buffer_12_543 = $signed(_T_93949); // @[Modules.scala 160:64:@41723.4]
  assign _T_93951 = $signed(buffer_12_493) + $signed(buffer_12_494); // @[Modules.scala 160:64:@41725.4]
  assign _T_93952 = _T_93951[13:0]; // @[Modules.scala 160:64:@41726.4]
  assign buffer_12_544 = $signed(_T_93952); // @[Modules.scala 160:64:@41727.4]
  assign _T_93954 = $signed(buffer_12_495) + $signed(buffer_12_496); // @[Modules.scala 160:64:@41729.4]
  assign _T_93955 = _T_93954[13:0]; // @[Modules.scala 160:64:@41730.4]
  assign buffer_12_545 = $signed(_T_93955); // @[Modules.scala 160:64:@41731.4]
  assign _T_93957 = $signed(buffer_12_497) + $signed(buffer_12_498); // @[Modules.scala 160:64:@41733.4]
  assign _T_93958 = _T_93957[13:0]; // @[Modules.scala 160:64:@41734.4]
  assign buffer_12_546 = $signed(_T_93958); // @[Modules.scala 160:64:@41735.4]
  assign _T_93960 = $signed(buffer_12_499) + $signed(buffer_12_500); // @[Modules.scala 160:64:@41737.4]
  assign _T_93961 = _T_93960[13:0]; // @[Modules.scala 160:64:@41738.4]
  assign buffer_12_547 = $signed(_T_93961); // @[Modules.scala 160:64:@41739.4]
  assign _T_93963 = $signed(buffer_12_501) + $signed(buffer_12_502); // @[Modules.scala 160:64:@41741.4]
  assign _T_93964 = _T_93963[13:0]; // @[Modules.scala 160:64:@41742.4]
  assign buffer_12_548 = $signed(_T_93964); // @[Modules.scala 160:64:@41743.4]
  assign _T_93966 = $signed(buffer_12_503) + $signed(buffer_12_504); // @[Modules.scala 160:64:@41745.4]
  assign _T_93967 = _T_93966[13:0]; // @[Modules.scala 160:64:@41746.4]
  assign buffer_12_549 = $signed(_T_93967); // @[Modules.scala 160:64:@41747.4]
  assign _T_93969 = $signed(buffer_8_524) + $signed(buffer_12_506); // @[Modules.scala 160:64:@41749.4]
  assign _T_93970 = _T_93969[13:0]; // @[Modules.scala 160:64:@41750.4]
  assign buffer_12_550 = $signed(_T_93970); // @[Modules.scala 160:64:@41751.4]
  assign _T_93972 = $signed(buffer_12_507) + $signed(buffer_12_508); // @[Modules.scala 160:64:@41753.4]
  assign _T_93973 = _T_93972[13:0]; // @[Modules.scala 160:64:@41754.4]
  assign buffer_12_551 = $signed(_T_93973); // @[Modules.scala 160:64:@41755.4]
  assign _T_93975 = $signed(buffer_12_509) + $signed(buffer_12_510); // @[Modules.scala 160:64:@41757.4]
  assign _T_93976 = _T_93975[13:0]; // @[Modules.scala 160:64:@41758.4]
  assign buffer_12_552 = $signed(_T_93976); // @[Modules.scala 160:64:@41759.4]
  assign _T_93978 = $signed(buffer_12_511) + $signed(buffer_12_512); // @[Modules.scala 160:64:@41761.4]
  assign _T_93979 = _T_93978[13:0]; // @[Modules.scala 160:64:@41762.4]
  assign buffer_12_553 = $signed(_T_93979); // @[Modules.scala 160:64:@41763.4]
  assign _T_93981 = $signed(buffer_12_513) + $signed(buffer_12_514); // @[Modules.scala 160:64:@41765.4]
  assign _T_93982 = _T_93981[13:0]; // @[Modules.scala 160:64:@41766.4]
  assign buffer_12_554 = $signed(_T_93982); // @[Modules.scala 160:64:@41767.4]
  assign _T_93984 = $signed(buffer_12_515) + $signed(buffer_12_516); // @[Modules.scala 160:64:@41769.4]
  assign _T_93985 = _T_93984[13:0]; // @[Modules.scala 160:64:@41770.4]
  assign buffer_12_555 = $signed(_T_93985); // @[Modules.scala 160:64:@41771.4]
  assign _T_93987 = $signed(buffer_12_517) + $signed(buffer_12_518); // @[Modules.scala 160:64:@41773.4]
  assign _T_93988 = _T_93987[13:0]; // @[Modules.scala 160:64:@41774.4]
  assign buffer_12_556 = $signed(_T_93988); // @[Modules.scala 160:64:@41775.4]
  assign _T_93990 = $signed(buffer_12_519) + $signed(buffer_3_548); // @[Modules.scala 160:64:@41777.4]
  assign _T_93991 = _T_93990[13:0]; // @[Modules.scala 160:64:@41778.4]
  assign buffer_12_557 = $signed(_T_93991); // @[Modules.scala 160:64:@41779.4]
  assign _T_93993 = $signed(buffer_12_521) + $signed(buffer_12_522); // @[Modules.scala 166:64:@41781.4]
  assign _T_93994 = _T_93993[13:0]; // @[Modules.scala 166:64:@41782.4]
  assign buffer_12_558 = $signed(_T_93994); // @[Modules.scala 166:64:@41783.4]
  assign _T_93996 = $signed(buffer_12_523) + $signed(buffer_12_524); // @[Modules.scala 166:64:@41785.4]
  assign _T_93997 = _T_93996[13:0]; // @[Modules.scala 166:64:@41786.4]
  assign buffer_12_559 = $signed(_T_93997); // @[Modules.scala 166:64:@41787.4]
  assign _T_93999 = $signed(buffer_12_525) + $signed(buffer_12_526); // @[Modules.scala 166:64:@41789.4]
  assign _T_94000 = _T_93999[13:0]; // @[Modules.scala 166:64:@41790.4]
  assign buffer_12_560 = $signed(_T_94000); // @[Modules.scala 166:64:@41791.4]
  assign _T_94002 = $signed(buffer_12_527) + $signed(buffer_12_528); // @[Modules.scala 166:64:@41793.4]
  assign _T_94003 = _T_94002[13:0]; // @[Modules.scala 166:64:@41794.4]
  assign buffer_12_561 = $signed(_T_94003); // @[Modules.scala 166:64:@41795.4]
  assign _T_94005 = $signed(buffer_12_529) + $signed(buffer_12_530); // @[Modules.scala 166:64:@41797.4]
  assign _T_94006 = _T_94005[13:0]; // @[Modules.scala 166:64:@41798.4]
  assign buffer_12_562 = $signed(_T_94006); // @[Modules.scala 166:64:@41799.4]
  assign _T_94008 = $signed(buffer_12_531) + $signed(buffer_12_532); // @[Modules.scala 166:64:@41801.4]
  assign _T_94009 = _T_94008[13:0]; // @[Modules.scala 166:64:@41802.4]
  assign buffer_12_563 = $signed(_T_94009); // @[Modules.scala 166:64:@41803.4]
  assign _T_94011 = $signed(buffer_12_533) + $signed(buffer_12_534); // @[Modules.scala 166:64:@41805.4]
  assign _T_94012 = _T_94011[13:0]; // @[Modules.scala 166:64:@41806.4]
  assign buffer_12_564 = $signed(_T_94012); // @[Modules.scala 166:64:@41807.4]
  assign _T_94014 = $signed(buffer_12_535) + $signed(buffer_12_536); // @[Modules.scala 166:64:@41809.4]
  assign _T_94015 = _T_94014[13:0]; // @[Modules.scala 166:64:@41810.4]
  assign buffer_12_565 = $signed(_T_94015); // @[Modules.scala 166:64:@41811.4]
  assign _T_94017 = $signed(buffer_12_537) + $signed(buffer_12_538); // @[Modules.scala 166:64:@41813.4]
  assign _T_94018 = _T_94017[13:0]; // @[Modules.scala 166:64:@41814.4]
  assign buffer_12_566 = $signed(_T_94018); // @[Modules.scala 166:64:@41815.4]
  assign _T_94020 = $signed(buffer_12_539) + $signed(buffer_12_540); // @[Modules.scala 166:64:@41817.4]
  assign _T_94021 = _T_94020[13:0]; // @[Modules.scala 166:64:@41818.4]
  assign buffer_12_567 = $signed(_T_94021); // @[Modules.scala 166:64:@41819.4]
  assign _T_94023 = $signed(buffer_12_541) + $signed(buffer_12_542); // @[Modules.scala 166:64:@41821.4]
  assign _T_94024 = _T_94023[13:0]; // @[Modules.scala 166:64:@41822.4]
  assign buffer_12_568 = $signed(_T_94024); // @[Modules.scala 166:64:@41823.4]
  assign _T_94026 = $signed(buffer_12_543) + $signed(buffer_12_544); // @[Modules.scala 166:64:@41825.4]
  assign _T_94027 = _T_94026[13:0]; // @[Modules.scala 166:64:@41826.4]
  assign buffer_12_569 = $signed(_T_94027); // @[Modules.scala 166:64:@41827.4]
  assign _T_94029 = $signed(buffer_12_545) + $signed(buffer_12_546); // @[Modules.scala 166:64:@41829.4]
  assign _T_94030 = _T_94029[13:0]; // @[Modules.scala 166:64:@41830.4]
  assign buffer_12_570 = $signed(_T_94030); // @[Modules.scala 166:64:@41831.4]
  assign _T_94032 = $signed(buffer_12_547) + $signed(buffer_12_548); // @[Modules.scala 166:64:@41833.4]
  assign _T_94033 = _T_94032[13:0]; // @[Modules.scala 166:64:@41834.4]
  assign buffer_12_571 = $signed(_T_94033); // @[Modules.scala 166:64:@41835.4]
  assign _T_94035 = $signed(buffer_12_549) + $signed(buffer_12_550); // @[Modules.scala 166:64:@41837.4]
  assign _T_94036 = _T_94035[13:0]; // @[Modules.scala 166:64:@41838.4]
  assign buffer_12_572 = $signed(_T_94036); // @[Modules.scala 166:64:@41839.4]
  assign _T_94038 = $signed(buffer_12_551) + $signed(buffer_12_552); // @[Modules.scala 166:64:@41841.4]
  assign _T_94039 = _T_94038[13:0]; // @[Modules.scala 166:64:@41842.4]
  assign buffer_12_573 = $signed(_T_94039); // @[Modules.scala 166:64:@41843.4]
  assign _T_94041 = $signed(buffer_12_553) + $signed(buffer_12_554); // @[Modules.scala 166:64:@41845.4]
  assign _T_94042 = _T_94041[13:0]; // @[Modules.scala 166:64:@41846.4]
  assign buffer_12_574 = $signed(_T_94042); // @[Modules.scala 166:64:@41847.4]
  assign _T_94044 = $signed(buffer_12_555) + $signed(buffer_12_556); // @[Modules.scala 166:64:@41849.4]
  assign _T_94045 = _T_94044[13:0]; // @[Modules.scala 166:64:@41850.4]
  assign buffer_12_575 = $signed(_T_94045); // @[Modules.scala 166:64:@41851.4]
  assign _T_94047 = $signed(buffer_12_557) + $signed(buffer_12_446); // @[Modules.scala 172:66:@41853.4]
  assign _T_94048 = _T_94047[13:0]; // @[Modules.scala 172:66:@41854.4]
  assign buffer_12_576 = $signed(_T_94048); // @[Modules.scala 172:66:@41855.4]
  assign _T_94050 = $signed(buffer_12_558) + $signed(buffer_12_559); // @[Modules.scala 166:64:@41857.4]
  assign _T_94051 = _T_94050[13:0]; // @[Modules.scala 166:64:@41858.4]
  assign buffer_12_577 = $signed(_T_94051); // @[Modules.scala 166:64:@41859.4]
  assign _T_94053 = $signed(buffer_12_560) + $signed(buffer_12_561); // @[Modules.scala 166:64:@41861.4]
  assign _T_94054 = _T_94053[13:0]; // @[Modules.scala 166:64:@41862.4]
  assign buffer_12_578 = $signed(_T_94054); // @[Modules.scala 166:64:@41863.4]
  assign _T_94056 = $signed(buffer_12_562) + $signed(buffer_12_563); // @[Modules.scala 166:64:@41865.4]
  assign _T_94057 = _T_94056[13:0]; // @[Modules.scala 166:64:@41866.4]
  assign buffer_12_579 = $signed(_T_94057); // @[Modules.scala 166:64:@41867.4]
  assign _T_94059 = $signed(buffer_12_564) + $signed(buffer_12_565); // @[Modules.scala 166:64:@41869.4]
  assign _T_94060 = _T_94059[13:0]; // @[Modules.scala 166:64:@41870.4]
  assign buffer_12_580 = $signed(_T_94060); // @[Modules.scala 166:64:@41871.4]
  assign _T_94062 = $signed(buffer_12_566) + $signed(buffer_12_567); // @[Modules.scala 166:64:@41873.4]
  assign _T_94063 = _T_94062[13:0]; // @[Modules.scala 166:64:@41874.4]
  assign buffer_12_581 = $signed(_T_94063); // @[Modules.scala 166:64:@41875.4]
  assign _T_94065 = $signed(buffer_12_568) + $signed(buffer_12_569); // @[Modules.scala 166:64:@41877.4]
  assign _T_94066 = _T_94065[13:0]; // @[Modules.scala 166:64:@41878.4]
  assign buffer_12_582 = $signed(_T_94066); // @[Modules.scala 166:64:@41879.4]
  assign _T_94068 = $signed(buffer_12_570) + $signed(buffer_12_571); // @[Modules.scala 166:64:@41881.4]
  assign _T_94069 = _T_94068[13:0]; // @[Modules.scala 166:64:@41882.4]
  assign buffer_12_583 = $signed(_T_94069); // @[Modules.scala 166:64:@41883.4]
  assign _T_94071 = $signed(buffer_12_572) + $signed(buffer_12_573); // @[Modules.scala 166:64:@41885.4]
  assign _T_94072 = _T_94071[13:0]; // @[Modules.scala 166:64:@41886.4]
  assign buffer_12_584 = $signed(_T_94072); // @[Modules.scala 166:64:@41887.4]
  assign _T_94074 = $signed(buffer_12_574) + $signed(buffer_12_575); // @[Modules.scala 166:64:@41889.4]
  assign _T_94075 = _T_94074[13:0]; // @[Modules.scala 166:64:@41890.4]
  assign buffer_12_585 = $signed(_T_94075); // @[Modules.scala 166:64:@41891.4]
  assign _T_94077 = $signed(buffer_12_577) + $signed(buffer_12_578); // @[Modules.scala 166:64:@41893.4]
  assign _T_94078 = _T_94077[13:0]; // @[Modules.scala 166:64:@41894.4]
  assign buffer_12_586 = $signed(_T_94078); // @[Modules.scala 166:64:@41895.4]
  assign _T_94080 = $signed(buffer_12_579) + $signed(buffer_12_580); // @[Modules.scala 166:64:@41897.4]
  assign _T_94081 = _T_94080[13:0]; // @[Modules.scala 166:64:@41898.4]
  assign buffer_12_587 = $signed(_T_94081); // @[Modules.scala 166:64:@41899.4]
  assign _T_94083 = $signed(buffer_12_581) + $signed(buffer_12_582); // @[Modules.scala 166:64:@41901.4]
  assign _T_94084 = _T_94083[13:0]; // @[Modules.scala 166:64:@41902.4]
  assign buffer_12_588 = $signed(_T_94084); // @[Modules.scala 166:64:@41903.4]
  assign _T_94086 = $signed(buffer_12_583) + $signed(buffer_12_584); // @[Modules.scala 166:64:@41905.4]
  assign _T_94087 = _T_94086[13:0]; // @[Modules.scala 166:64:@41906.4]
  assign buffer_12_589 = $signed(_T_94087); // @[Modules.scala 166:64:@41907.4]
  assign _T_94089 = $signed(buffer_12_585) + $signed(buffer_12_576); // @[Modules.scala 172:66:@41909.4]
  assign _T_94090 = _T_94089[13:0]; // @[Modules.scala 172:66:@41910.4]
  assign buffer_12_590 = $signed(_T_94090); // @[Modules.scala 172:66:@41911.4]
  assign _T_94092 = $signed(buffer_12_586) + $signed(buffer_12_587); // @[Modules.scala 166:64:@41913.4]
  assign _T_94093 = _T_94092[13:0]; // @[Modules.scala 166:64:@41914.4]
  assign buffer_12_591 = $signed(_T_94093); // @[Modules.scala 166:64:@41915.4]
  assign _T_94095 = $signed(buffer_12_588) + $signed(buffer_12_589); // @[Modules.scala 166:64:@41917.4]
  assign _T_94096 = _T_94095[13:0]; // @[Modules.scala 166:64:@41918.4]
  assign buffer_12_592 = $signed(_T_94096); // @[Modules.scala 166:64:@41919.4]
  assign _T_94098 = $signed(buffer_12_591) + $signed(buffer_12_592); // @[Modules.scala 160:64:@41921.4]
  assign _T_94099 = _T_94098[13:0]; // @[Modules.scala 160:64:@41922.4]
  assign buffer_12_593 = $signed(_T_94099); // @[Modules.scala 160:64:@41923.4]
  assign _T_94101 = $signed(buffer_12_593) + $signed(buffer_12_590); // @[Modules.scala 172:66:@41925.4]
  assign _T_94102 = _T_94101[13:0]; // @[Modules.scala 172:66:@41926.4]
  assign buffer_12_594 = $signed(_T_94102); // @[Modules.scala 172:66:@41927.4]
  assign _T_94105 = $signed(-4'sh1) * $signed(io_in_10); // @[Modules.scala 143:74:@42118.4]
  assign _T_94108 = $signed(_T_94105) + $signed(_T_60255); // @[Modules.scala 143:103:@42120.4]
  assign _T_94109 = _T_94108[4:0]; // @[Modules.scala 143:103:@42121.4]
  assign _T_94110 = $signed(_T_94109); // @[Modules.scala 143:103:@42122.4]
  assign _T_94114 = $signed(-4'sh1) * $signed(io_in_23); // @[Modules.scala 144:80:@42125.4]
  assign _T_94115 = $signed(_T_60257) + $signed(_T_94114); // @[Modules.scala 143:103:@42126.4]
  assign _T_94116 = _T_94115[4:0]; // @[Modules.scala 143:103:@42127.4]
  assign _T_94117 = $signed(_T_94116); // @[Modules.scala 143:103:@42128.4]
  assign _T_94143 = $signed(_GEN_498) + $signed(_T_54234); // @[Modules.scala 143:103:@42150.4]
  assign _T_94144 = _T_94143[5:0]; // @[Modules.scala 143:103:@42151.4]
  assign _T_94145 = $signed(_T_94144); // @[Modules.scala 143:103:@42152.4]
  assign _T_94150 = $signed(_T_54236) + $signed(_T_54243); // @[Modules.scala 143:103:@42156.4]
  assign _T_94151 = _T_94150[5:0]; // @[Modules.scala 143:103:@42157.4]
  assign _T_94152 = $signed(_T_94151); // @[Modules.scala 143:103:@42158.4]
  assign _T_94164 = $signed(_T_57262) + $signed(_T_63403); // @[Modules.scala 143:103:@42168.4]
  assign _T_94165 = _T_94164[4:0]; // @[Modules.scala 143:103:@42169.4]
  assign _T_94166 = $signed(_T_94165); // @[Modules.scala 143:103:@42170.4]
  assign _T_94178 = $signed(_T_54276) + $signed(_GEN_281); // @[Modules.scala 143:103:@42180.4]
  assign _T_94179 = _T_94178[5:0]; // @[Modules.scala 143:103:@42181.4]
  assign _T_94180 = $signed(_T_94179); // @[Modules.scala 143:103:@42182.4]
  assign _T_94185 = $signed(_T_57288) + $signed(_T_60332); // @[Modules.scala 143:103:@42186.4]
  assign _T_94186 = _T_94185[4:0]; // @[Modules.scala 143:103:@42187.4]
  assign _T_94187 = $signed(_T_94186); // @[Modules.scala 143:103:@42188.4]
  assign _GEN_909 = {{1{_T_57302[4]}},_T_57302}; // @[Modules.scala 143:103:@42192.4]
  assign _T_94192 = $signed(_T_54285) + $signed(_GEN_909); // @[Modules.scala 143:103:@42192.4]
  assign _T_94193 = _T_94192[5:0]; // @[Modules.scala 143:103:@42193.4]
  assign _T_94194 = $signed(_T_94193); // @[Modules.scala 143:103:@42194.4]
  assign _T_94254 = $signed(-4'sh1) * $signed(io_in_83); // @[Modules.scala 144:80:@42245.4]
  assign _GEN_910 = {{1{_T_94254[4]}},_T_94254}; // @[Modules.scala 143:103:@42246.4]
  assign _T_94255 = $signed(_T_54353) + $signed(_GEN_910); // @[Modules.scala 143:103:@42246.4]
  assign _T_94256 = _T_94255[5:0]; // @[Modules.scala 143:103:@42247.4]
  assign _T_94257 = $signed(_T_94256); // @[Modules.scala 143:103:@42248.4]
  assign _GEN_911 = {{1{_T_60402[4]}},_T_60402}; // @[Modules.scala 143:103:@42258.4]
  assign _T_94269 = $signed(_GEN_911) + $signed(_T_54367); // @[Modules.scala 143:103:@42258.4]
  assign _T_94270 = _T_94269[5:0]; // @[Modules.scala 143:103:@42259.4]
  assign _T_94271 = $signed(_T_94270); // @[Modules.scala 143:103:@42260.4]
  assign _T_94360 = $signed(_T_54451) + $signed(_T_57456); // @[Modules.scala 143:103:@42336.4]
  assign _T_94361 = _T_94360[5:0]; // @[Modules.scala 143:103:@42337.4]
  assign _T_94362 = $signed(_T_94361); // @[Modules.scala 143:103:@42338.4]
  assign _T_94395 = $signed(_GEN_151) + $signed(_T_54486); // @[Modules.scala 143:103:@42366.4]
  assign _T_94396 = _T_94395[5:0]; // @[Modules.scala 143:103:@42367.4]
  assign _T_94397 = $signed(_T_94396); // @[Modules.scala 143:103:@42368.4]
  assign _T_94402 = $signed(_T_54493) + $signed(_GEN_639); // @[Modules.scala 143:103:@42372.4]
  assign _T_94403 = _T_94402[5:0]; // @[Modules.scala 143:103:@42373.4]
  assign _T_94404 = $signed(_T_94403); // @[Modules.scala 143:103:@42374.4]
  assign _T_94423 = $signed(_GEN_152) + $signed(_T_57526); // @[Modules.scala 143:103:@42390.4]
  assign _T_94424 = _T_94423[5:0]; // @[Modules.scala 143:103:@42391.4]
  assign _T_94425 = $signed(_T_94424); // @[Modules.scala 143:103:@42392.4]
  assign _T_94444 = $signed(_T_54530) + $signed(_T_54535); // @[Modules.scala 143:103:@42408.4]
  assign _T_94445 = _T_94444[5:0]; // @[Modules.scala 143:103:@42409.4]
  assign _T_94446 = $signed(_T_94445); // @[Modules.scala 143:103:@42410.4]
  assign _T_94451 = $signed(_T_54537) + $signed(_GEN_642); // @[Modules.scala 143:103:@42414.4]
  assign _T_94452 = _T_94451[5:0]; // @[Modules.scala 143:103:@42415.4]
  assign _T_94453 = $signed(_T_94452); // @[Modules.scala 143:103:@42416.4]
  assign _T_94493 = $signed(_T_57596) + $signed(_T_63746); // @[Modules.scala 143:103:@42450.4]
  assign _T_94494 = _T_94493[4:0]; // @[Modules.scala 143:103:@42451.4]
  assign _T_94495 = $signed(_T_94494); // @[Modules.scala 143:103:@42452.4]
  assign _GEN_916 = {{1{_T_54612[4]}},_T_54612}; // @[Modules.scala 143:103:@42486.4]
  assign _T_94535 = $signed(_T_57626) + $signed(_GEN_916); // @[Modules.scala 143:103:@42486.4]
  assign _T_94536 = _T_94535[5:0]; // @[Modules.scala 143:103:@42487.4]
  assign _T_94537 = $signed(_T_94536); // @[Modules.scala 143:103:@42488.4]
  assign _T_94563 = $signed(_T_54633) + $signed(_T_60689); // @[Modules.scala 143:103:@42510.4]
  assign _T_94564 = _T_94563[4:0]; // @[Modules.scala 143:103:@42511.4]
  assign _T_94565 = $signed(_T_94564); // @[Modules.scala 143:103:@42512.4]
  assign _GEN_918 = {{1{_T_60745[4]}},_T_60745}; // @[Modules.scala 143:103:@42558.4]
  assign _T_94619 = $signed(_T_54689) + $signed(_GEN_918); // @[Modules.scala 143:103:@42558.4]
  assign _T_94620 = _T_94619[5:0]; // @[Modules.scala 143:103:@42559.4]
  assign _T_94621 = $signed(_T_94620); // @[Modules.scala 143:103:@42560.4]
  assign _T_94626 = $signed(_T_60747) + $signed(_T_60752); // @[Modules.scala 143:103:@42564.4]
  assign _T_94627 = _T_94626[4:0]; // @[Modules.scala 143:103:@42565.4]
  assign _T_94628 = $signed(_T_94627); // @[Modules.scala 143:103:@42566.4]
  assign _T_94647 = $signed(_T_54698) + $signed(_T_60773); // @[Modules.scala 143:103:@42582.4]
  assign _T_94648 = _T_94647[4:0]; // @[Modules.scala 143:103:@42583.4]
  assign _T_94649 = $signed(_T_94648); // @[Modules.scala 143:103:@42584.4]
  assign _GEN_920 = {{1{_T_54719[4]}},_T_54719}; // @[Modules.scala 143:103:@42594.4]
  assign _T_94661 = $signed(_T_63900) + $signed(_GEN_920); // @[Modules.scala 143:103:@42594.4]
  assign _T_94662 = _T_94661[5:0]; // @[Modules.scala 143:103:@42595.4]
  assign _T_94663 = $signed(_T_94662); // @[Modules.scala 143:103:@42596.4]
  assign _T_94675 = $signed(_GEN_18) + $signed(_T_54738); // @[Modules.scala 143:103:@42606.4]
  assign _T_94676 = _T_94675[5:0]; // @[Modules.scala 143:103:@42607.4]
  assign _T_94677 = $signed(_T_94676); // @[Modules.scala 143:103:@42608.4]
  assign _T_94696 = $signed(_T_60829) + $signed(_T_57794); // @[Modules.scala 143:103:@42624.4]
  assign _T_94697 = _T_94696[4:0]; // @[Modules.scala 143:103:@42625.4]
  assign _T_94698 = $signed(_T_94697); // @[Modules.scala 143:103:@42626.4]
  assign _T_94703 = $signed(_T_60838) + $signed(_T_60843); // @[Modules.scala 143:103:@42630.4]
  assign _T_94704 = _T_94703[4:0]; // @[Modules.scala 143:103:@42631.4]
  assign _T_94705 = $signed(_T_94704); // @[Modules.scala 143:103:@42632.4]
  assign _T_94717 = $signed(_T_54768) + $signed(_T_54773); // @[Modules.scala 143:103:@42642.4]
  assign _T_94718 = _T_94717[4:0]; // @[Modules.scala 143:103:@42643.4]
  assign _T_94719 = $signed(_T_94718); // @[Modules.scala 143:103:@42644.4]
  assign _GEN_923 = {{1{_T_54775[4]}},_T_54775}; // @[Modules.scala 143:103:@42648.4]
  assign _T_94724 = $signed(_GEN_923) + $signed(_T_70099); // @[Modules.scala 143:103:@42648.4]
  assign _T_94725 = _T_94724[5:0]; // @[Modules.scala 143:103:@42649.4]
  assign _T_94726 = $signed(_T_94725); // @[Modules.scala 143:103:@42650.4]
  assign _GEN_924 = {{1{_T_54801[4]}},_T_54801}; // @[Modules.scala 143:103:@42660.4]
  assign _T_94738 = $signed(_GEN_924) + $signed(_T_63989); // @[Modules.scala 143:103:@42660.4]
  assign _T_94739 = _T_94738[5:0]; // @[Modules.scala 143:103:@42661.4]
  assign _T_94740 = $signed(_T_94739); // @[Modules.scala 143:103:@42662.4]
  assign _T_94773 = $signed(_T_70148) + $signed(_GEN_167); // @[Modules.scala 143:103:@42690.4]
  assign _T_94774 = _T_94773[5:0]; // @[Modules.scala 143:103:@42691.4]
  assign _T_94775 = $signed(_T_94774); // @[Modules.scala 143:103:@42692.4]
  assign _T_94780 = $signed(_T_54829) + $signed(_T_54836); // @[Modules.scala 143:103:@42696.4]
  assign _T_94781 = _T_94780[4:0]; // @[Modules.scala 143:103:@42697.4]
  assign _T_94782 = $signed(_T_94781); // @[Modules.scala 143:103:@42698.4]
  assign _GEN_927 = {{1{_T_54885[4]}},_T_54885}; // @[Modules.scala 143:103:@42738.4]
  assign _T_94829 = $signed(_GEN_927) + $signed(_T_64075); // @[Modules.scala 143:103:@42738.4]
  assign _T_94830 = _T_94829[5:0]; // @[Modules.scala 143:103:@42739.4]
  assign _T_94831 = $signed(_T_94830); // @[Modules.scala 143:103:@42740.4]
  assign _T_94836 = $signed(_T_54894) + $signed(_T_70220); // @[Modules.scala 143:103:@42744.4]
  assign _T_94837 = _T_94836[4:0]; // @[Modules.scala 143:103:@42745.4]
  assign _T_94838 = $signed(_T_94837); // @[Modules.scala 143:103:@42746.4]
  assign _T_94843 = $signed(_T_54901) + $signed(_T_54906); // @[Modules.scala 143:103:@42750.4]
  assign _T_94844 = _T_94843[5:0]; // @[Modules.scala 143:103:@42751.4]
  assign _T_94845 = $signed(_T_94844); // @[Modules.scala 143:103:@42752.4]
  assign _T_94850 = $signed(_T_57941) + $signed(_T_67200); // @[Modules.scala 143:103:@42756.4]
  assign _T_94851 = _T_94850[5:0]; // @[Modules.scala 143:103:@42757.4]
  assign _T_94852 = $signed(_T_94851); // @[Modules.scala 143:103:@42758.4]
  assign _GEN_928 = {{1{_T_54922[4]}},_T_54922}; // @[Modules.scala 143:103:@42762.4]
  assign _T_94857 = $signed(_T_64103) + $signed(_GEN_928); // @[Modules.scala 143:103:@42762.4]
  assign _T_94858 = _T_94857[5:0]; // @[Modules.scala 143:103:@42763.4]
  assign _T_94859 = $signed(_T_94858); // @[Modules.scala 143:103:@42764.4]
  assign _T_94864 = $signed(_T_54927) + $signed(_T_54934); // @[Modules.scala 143:103:@42768.4]
  assign _T_94865 = _T_94864[4:0]; // @[Modules.scala 143:103:@42769.4]
  assign _T_94866 = $signed(_T_94865); // @[Modules.scala 143:103:@42770.4]
  assign _GEN_929 = {{1{_T_54964[4]}},_T_54964}; // @[Modules.scala 143:103:@42792.4]
  assign _T_94892 = $signed(_T_57981) + $signed(_GEN_929); // @[Modules.scala 143:103:@42792.4]
  assign _T_94893 = _T_94892[5:0]; // @[Modules.scala 143:103:@42793.4]
  assign _T_94894 = $signed(_T_94893); // @[Modules.scala 143:103:@42794.4]
  assign _T_94899 = $signed(_T_67247) + $signed(_T_70281); // @[Modules.scala 143:103:@42798.4]
  assign _T_94900 = _T_94899[5:0]; // @[Modules.scala 143:103:@42799.4]
  assign _T_94901 = $signed(_T_94900); // @[Modules.scala 143:103:@42800.4]
  assign _GEN_930 = {{1{_T_54983[4]}},_T_54983}; // @[Modules.scala 143:103:@42810.4]
  assign _T_94913 = $signed(_GEN_930) + $signed(_T_54997); // @[Modules.scala 143:103:@42810.4]
  assign _T_94914 = _T_94913[5:0]; // @[Modules.scala 143:103:@42811.4]
  assign _T_94915 = $signed(_T_94914); // @[Modules.scala 143:103:@42812.4]
  assign _T_94920 = $signed(_T_58025) + $signed(_GEN_100); // @[Modules.scala 143:103:@42816.4]
  assign _T_94921 = _T_94920[5:0]; // @[Modules.scala 143:103:@42817.4]
  assign _T_94922 = $signed(_T_94921); // @[Modules.scala 143:103:@42818.4]
  assign _T_94927 = $signed(_T_55006) + $signed(_T_55011); // @[Modules.scala 143:103:@42822.4]
  assign _T_94928 = _T_94927[4:0]; // @[Modules.scala 143:103:@42823.4]
  assign _T_94929 = $signed(_T_94928); // @[Modules.scala 143:103:@42824.4]
  assign _T_94955 = $signed(_T_61104) + $signed(_T_61109); // @[Modules.scala 143:103:@42846.4]
  assign _T_94956 = _T_94955[4:0]; // @[Modules.scala 143:103:@42847.4]
  assign _T_94957 = $signed(_T_94956); // @[Modules.scala 143:103:@42848.4]
  assign _T_94962 = $signed(_T_58067) + $signed(_T_58074); // @[Modules.scala 143:103:@42852.4]
  assign _T_94963 = _T_94962[5:0]; // @[Modules.scala 143:103:@42853.4]
  assign _T_94964 = $signed(_T_94963); // @[Modules.scala 143:103:@42854.4]
  assign _T_94976 = $signed(_T_70351) + $signed(_GEN_521); // @[Modules.scala 143:103:@42864.4]
  assign _T_94977 = _T_94976[5:0]; // @[Modules.scala 143:103:@42865.4]
  assign _T_94978 = $signed(_T_94977); // @[Modules.scala 143:103:@42866.4]
  assign _GEN_934 = {{1{_T_67340[4]}},_T_67340}; // @[Modules.scala 143:103:@42876.4]
  assign _T_94990 = $signed(_GEN_934) + $signed(_T_55076); // @[Modules.scala 143:103:@42876.4]
  assign _T_94991 = _T_94990[5:0]; // @[Modules.scala 143:103:@42877.4]
  assign _T_94992 = $signed(_T_94991); // @[Modules.scala 143:103:@42878.4]
  assign _T_95032 = $signed(_T_58142) + $signed(_T_58151); // @[Modules.scala 143:103:@42912.4]
  assign _T_95033 = _T_95032[5:0]; // @[Modules.scala 143:103:@42913.4]
  assign _T_95034 = $signed(_T_95033); // @[Modules.scala 143:103:@42914.4]
  assign _T_95039 = $signed(_T_55132) + $signed(_T_73565); // @[Modules.scala 143:103:@42918.4]
  assign _T_95040 = _T_95039[4:0]; // @[Modules.scala 143:103:@42919.4]
  assign _T_95041 = $signed(_T_95040); // @[Modules.scala 143:103:@42920.4]
  assign _GEN_935 = {{1{_T_55146[4]}},_T_55146}; // @[Modules.scala 143:103:@42930.4]
  assign _T_95053 = $signed(_GEN_935) + $signed(_T_55151); // @[Modules.scala 143:103:@42930.4]
  assign _T_95054 = _T_95053[5:0]; // @[Modules.scala 143:103:@42931.4]
  assign _T_95055 = $signed(_T_95054); // @[Modules.scala 143:103:@42932.4]
  assign _GEN_936 = {{1{_T_61244[4]}},_T_61244}; // @[Modules.scala 143:103:@42948.4]
  assign _T_95074 = $signed(_T_55172) + $signed(_GEN_936); // @[Modules.scala 143:103:@42948.4]
  assign _T_95075 = _T_95074[5:0]; // @[Modules.scala 143:103:@42949.4]
  assign _T_95076 = $signed(_T_95075); // @[Modules.scala 143:103:@42950.4]
  assign _T_95102 = $signed(_GEN_105) + $signed(_T_61272); // @[Modules.scala 143:103:@42972.4]
  assign _T_95103 = _T_95102[5:0]; // @[Modules.scala 143:103:@42973.4]
  assign _T_95104 = $signed(_T_95103); // @[Modules.scala 143:103:@42974.4]
  assign _GEN_938 = {{1{_T_73663[4]}},_T_73663}; // @[Modules.scala 143:103:@42990.4]
  assign _T_95123 = $signed(_T_58240) + $signed(_GEN_938); // @[Modules.scala 143:103:@42990.4]
  assign _T_95124 = _T_95123[5:0]; // @[Modules.scala 143:103:@42991.4]
  assign _T_95125 = $signed(_T_95124); // @[Modules.scala 143:103:@42992.4]
  assign _GEN_939 = {{1{_T_76787[4]}},_T_76787}; // @[Modules.scala 143:103:@42996.4]
  assign _T_95130 = $signed(_GEN_939) + $signed(_T_61307); // @[Modules.scala 143:103:@42996.4]
  assign _T_95131 = _T_95130[5:0]; // @[Modules.scala 143:103:@42997.4]
  assign _T_95132 = $signed(_T_95131); // @[Modules.scala 143:103:@42998.4]
  assign _T_95151 = $signed(_T_55249) + $signed(_T_58282); // @[Modules.scala 143:103:@43014.4]
  assign _T_95152 = _T_95151[5:0]; // @[Modules.scala 143:103:@43015.4]
  assign _T_95153 = $signed(_T_95152); // @[Modules.scala 143:103:@43016.4]
  assign _T_95172 = $signed(_T_55270) + $signed(_T_55277); // @[Modules.scala 143:103:@43032.4]
  assign _T_95173 = _T_95172[4:0]; // @[Modules.scala 143:103:@43033.4]
  assign _T_95174 = $signed(_T_95173); // @[Modules.scala 143:103:@43034.4]
  assign _T_95214 = $signed(_T_70589) + $signed(_T_58326); // @[Modules.scala 143:103:@43068.4]
  assign _T_95215 = _T_95214[4:0]; // @[Modules.scala 143:103:@43069.4]
  assign _T_95216 = $signed(_T_95215); // @[Modules.scala 143:103:@43070.4]
  assign _GEN_940 = {{1{_T_58338[4]}},_T_58338}; // @[Modules.scala 143:103:@43080.4]
  assign _T_95228 = $signed(_GEN_940) + $signed(_T_55319); // @[Modules.scala 143:103:@43080.4]
  assign _T_95229 = _T_95228[5:0]; // @[Modules.scala 143:103:@43081.4]
  assign _T_95230 = $signed(_T_95229); // @[Modules.scala 143:103:@43082.4]
  assign _T_95235 = $signed(_T_70605) + $signed(_T_55326); // @[Modules.scala 143:103:@43086.4]
  assign _T_95236 = _T_95235[5:0]; // @[Modules.scala 143:103:@43087.4]
  assign _T_95237 = $signed(_T_95236); // @[Modules.scala 143:103:@43088.4]
  assign _T_95242 = $signed(_T_67585) + $signed(_T_55328); // @[Modules.scala 143:103:@43092.4]
  assign _T_95243 = _T_95242[5:0]; // @[Modules.scala 143:103:@43093.4]
  assign _T_95244 = $signed(_T_95243); // @[Modules.scala 143:103:@43094.4]
  assign _T_95270 = $signed(_T_61438) + $signed(_GEN_394); // @[Modules.scala 143:103:@43116.4]
  assign _T_95271 = _T_95270[5:0]; // @[Modules.scala 143:103:@43117.4]
  assign _T_95272 = $signed(_T_95271); // @[Modules.scala 143:103:@43118.4]
  assign _T_95277 = $signed(_T_61440) + $signed(_T_61445); // @[Modules.scala 143:103:@43122.4]
  assign _T_95278 = _T_95277[5:0]; // @[Modules.scala 143:103:@43123.4]
  assign _T_95279 = $signed(_T_95278); // @[Modules.scala 143:103:@43124.4]
  assign _GEN_942 = {{1{_T_61475[4]}},_T_61475}; // @[Modules.scala 143:103:@43146.4]
  assign _T_95305 = $signed(_T_61468) + $signed(_GEN_942); // @[Modules.scala 143:103:@43146.4]
  assign _T_95306 = _T_95305[5:0]; // @[Modules.scala 143:103:@43147.4]
  assign _T_95307 = $signed(_T_95306); // @[Modules.scala 143:103:@43148.4]
  assign _T_95312 = $signed(_T_64579) + $signed(_T_55398); // @[Modules.scala 143:103:@43152.4]
  assign _T_95313 = _T_95312[4:0]; // @[Modules.scala 143:103:@43153.4]
  assign _T_95314 = $signed(_T_95313); // @[Modules.scala 143:103:@43154.4]
  assign _T_95326 = $signed(_T_55410) + $signed(_T_58424); // @[Modules.scala 143:103:@43164.4]
  assign _T_95327 = _T_95326[5:0]; // @[Modules.scala 143:103:@43165.4]
  assign _T_95328 = $signed(_T_95327); // @[Modules.scala 143:103:@43166.4]
  assign _T_95375 = $signed(_T_61545) + $signed(_GEN_51); // @[Modules.scala 143:103:@43206.4]
  assign _T_95376 = _T_95375[5:0]; // @[Modules.scala 143:103:@43207.4]
  assign _T_95377 = $signed(_T_95376); // @[Modules.scala 143:103:@43208.4]
  assign _T_95389 = $signed(_T_70766) + $signed(_T_55480); // @[Modules.scala 143:103:@43218.4]
  assign _T_95390 = _T_95389[5:0]; // @[Modules.scala 143:103:@43219.4]
  assign _T_95391 = $signed(_T_95390); // @[Modules.scala 143:103:@43220.4]
  assign _T_95410 = $signed(_T_55494) + $signed(_T_70799); // @[Modules.scala 143:103:@43236.4]
  assign _T_95411 = _T_95410[5:0]; // @[Modules.scala 143:103:@43237.4]
  assign _T_95412 = $signed(_T_95411); // @[Modules.scala 143:103:@43238.4]
  assign _T_95452 = $signed(_T_61622) + $signed(_GEN_55); // @[Modules.scala 143:103:@43272.4]
  assign _T_95453 = _T_95452[5:0]; // @[Modules.scala 143:103:@43273.4]
  assign _T_95454 = $signed(_T_95453); // @[Modules.scala 143:103:@43274.4]
  assign _GEN_946 = {{1{_T_58562[4]}},_T_58562}; // @[Modules.scala 143:103:@43278.4]
  assign _T_95459 = $signed(_GEN_946) + $signed(_T_67767); // @[Modules.scala 143:103:@43278.4]
  assign _T_95460 = _T_95459[5:0]; // @[Modules.scala 143:103:@43279.4]
  assign _T_95461 = $signed(_T_95460); // @[Modules.scala 143:103:@43280.4]
  assign _T_95494 = $signed(_T_70855) + $signed(_T_64782); // @[Modules.scala 143:103:@43308.4]
  assign _T_95495 = _T_95494[4:0]; // @[Modules.scala 143:103:@43309.4]
  assign _T_95496 = $signed(_T_95495); // @[Modules.scala 143:103:@43310.4]
  assign _T_95508 = $signed(_T_55578) + $signed(_T_70876); // @[Modules.scala 143:103:@43320.4]
  assign _T_95509 = _T_95508[5:0]; // @[Modules.scala 143:103:@43321.4]
  assign _T_95510 = $signed(_T_95509); // @[Modules.scala 143:103:@43322.4]
  assign _T_95536 = $signed(_T_55606) + $signed(_T_55629); // @[Modules.scala 143:103:@43344.4]
  assign _T_95537 = _T_95536[5:0]; // @[Modules.scala 143:103:@43345.4]
  assign _T_95538 = $signed(_T_95537); // @[Modules.scala 143:103:@43346.4]
  assign _GEN_951 = {{1{_T_61753[4]}},_T_61753}; // @[Modules.scala 143:103:@43374.4]
  assign _T_95571 = $signed(_T_55664) + $signed(_GEN_951); // @[Modules.scala 143:103:@43374.4]
  assign _T_95572 = _T_95571[5:0]; // @[Modules.scala 143:103:@43375.4]
  assign _T_95573 = $signed(_T_95572); // @[Modules.scala 143:103:@43376.4]
  assign _T_95578 = $signed(_GEN_478) + $signed(_T_55676); // @[Modules.scala 143:103:@43380.4]
  assign _T_95579 = _T_95578[5:0]; // @[Modules.scala 143:103:@43381.4]
  assign _T_95580 = $signed(_T_95579); // @[Modules.scala 143:103:@43382.4]
  assign _T_95585 = $signed(_T_55678) + $signed(_T_55683); // @[Modules.scala 143:103:@43386.4]
  assign _T_95586 = _T_95585[5:0]; // @[Modules.scala 143:103:@43387.4]
  assign _T_95587 = $signed(_T_95586); // @[Modules.scala 143:103:@43388.4]
  assign _T_95592 = $signed(_T_55685) + $signed(_T_55690); // @[Modules.scala 143:103:@43392.4]
  assign _T_95593 = _T_95592[5:0]; // @[Modules.scala 143:103:@43393.4]
  assign _T_95594 = $signed(_T_95593); // @[Modules.scala 143:103:@43394.4]
  assign _T_95620 = $signed(_GEN_739) + $signed(_T_71002); // @[Modules.scala 143:103:@43416.4]
  assign _T_95621 = _T_95620[5:0]; // @[Modules.scala 143:103:@43417.4]
  assign _T_95622 = $signed(_T_95621); // @[Modules.scala 143:103:@43418.4]
  assign _T_95627 = $signed(_T_71004) + $signed(_T_71009); // @[Modules.scala 143:103:@43422.4]
  assign _T_95628 = _T_95627[5:0]; // @[Modules.scala 143:103:@43423.4]
  assign _T_95629 = $signed(_T_95628); // @[Modules.scala 143:103:@43424.4]
  assign _T_95704 = $signed(_T_55776) + $signed(_T_55781); // @[Modules.scala 143:103:@43488.4]
  assign _T_95705 = _T_95704[5:0]; // @[Modules.scala 143:103:@43489.4]
  assign _T_95706 = $signed(_T_95705); // @[Modules.scala 143:103:@43490.4]
  assign _GEN_957 = {{1{_T_61914[4]}},_T_61914}; // @[Modules.scala 143:103:@43524.4]
  assign _T_95746 = $signed(_GEN_957) + $signed(_T_77464); // @[Modules.scala 143:103:@43524.4]
  assign _T_95747 = _T_95746[5:0]; // @[Modules.scala 143:103:@43525.4]
  assign _T_95748 = $signed(_T_95747); // @[Modules.scala 143:103:@43526.4]
  assign _T_95781 = $signed(_GEN_545) + $signed(_T_55839); // @[Modules.scala 143:103:@43554.4]
  assign _T_95782 = _T_95781[5:0]; // @[Modules.scala 143:103:@43555.4]
  assign _T_95783 = $signed(_T_95782); // @[Modules.scala 143:103:@43556.4]
  assign _T_95823 = $signed(_T_55888) + $signed(_T_58919); // @[Modules.scala 143:103:@43590.4]
  assign _T_95824 = _T_95823[5:0]; // @[Modules.scala 143:103:@43591.4]
  assign _T_95825 = $signed(_T_95824); // @[Modules.scala 143:103:@43592.4]
  assign _T_95844 = $signed(_T_58933) + $signed(_T_62026); // @[Modules.scala 143:103:@43608.4]
  assign _T_95845 = _T_95844[5:0]; // @[Modules.scala 143:103:@43609.4]
  assign _T_95846 = $signed(_T_95845); // @[Modules.scala 143:103:@43610.4]
  assign _GEN_964 = {{1{_T_68171[4]}},_T_68171}; // @[Modules.scala 143:103:@43614.4]
  assign _T_95851 = $signed(_GEN_964) + $signed(_T_55923); // @[Modules.scala 143:103:@43614.4]
  assign _T_95852 = _T_95851[5:0]; // @[Modules.scala 143:103:@43615.4]
  assign _T_95853 = $signed(_T_95852); // @[Modules.scala 143:103:@43616.4]
  assign _GEN_965 = {{1{_T_62061[4]}},_T_62061}; // @[Modules.scala 143:103:@43650.4]
  assign _T_95893 = $signed(_GEN_965) + $signed(_T_55965); // @[Modules.scala 143:103:@43650.4]
  assign _T_95894 = _T_95893[5:0]; // @[Modules.scala 143:103:@43651.4]
  assign _T_95895 = $signed(_T_95894); // @[Modules.scala 143:103:@43652.4]
  assign _T_95900 = $signed(_T_58982) + $signed(_T_71303); // @[Modules.scala 143:103:@43656.4]
  assign _T_95901 = _T_95900[5:0]; // @[Modules.scala 143:103:@43657.4]
  assign _T_95902 = $signed(_T_95901); // @[Modules.scala 143:103:@43658.4]
  assign _T_95907 = $signed(_T_65188) + $signed(_T_71317); // @[Modules.scala 143:103:@43662.4]
  assign _T_95908 = _T_95907[5:0]; // @[Modules.scala 143:103:@43663.4]
  assign _T_95909 = $signed(_T_95908); // @[Modules.scala 143:103:@43664.4]
  assign _GEN_966 = {{1{_T_55998[4]}},_T_55998}; // @[Modules.scala 143:103:@43674.4]
  assign _T_95921 = $signed(_GEN_966) + $signed(_T_62103); // @[Modules.scala 143:103:@43674.4]
  assign _T_95922 = _T_95921[5:0]; // @[Modules.scala 143:103:@43675.4]
  assign _T_95923 = $signed(_T_95922); // @[Modules.scala 143:103:@43676.4]
  assign _GEN_968 = {{1{_T_56061[4]}},_T_56061}; // @[Modules.scala 143:103:@43734.4]
  assign _T_95991 = $signed(_T_71389) + $signed(_GEN_968); // @[Modules.scala 143:103:@43734.4]
  assign _T_95992 = _T_95991[5:0]; // @[Modules.scala 143:103:@43735.4]
  assign _T_95993 = $signed(_T_95992); // @[Modules.scala 143:103:@43736.4]
  assign _T_95998 = $signed(_T_71396) + $signed(_T_59075); // @[Modules.scala 143:103:@43740.4]
  assign _T_95999 = _T_95998[5:0]; // @[Modules.scala 143:103:@43741.4]
  assign _T_96000 = $signed(_T_95999); // @[Modules.scala 143:103:@43742.4]
  assign _T_96075 = $signed(_T_62231) + $signed(_T_65354); // @[Modules.scala 143:103:@43806.4]
  assign _T_96076 = _T_96075[4:0]; // @[Modules.scala 143:103:@43807.4]
  assign _T_96077 = $signed(_T_96076); // @[Modules.scala 143:103:@43808.4]
  assign _T_96138 = $signed(_T_59199) + $signed(_T_65410); // @[Modules.scala 143:103:@43860.4]
  assign _T_96139 = _T_96138[4:0]; // @[Modules.scala 143:103:@43861.4]
  assign _T_96140 = $signed(_T_96139); // @[Modules.scala 143:103:@43862.4]
  assign _T_96215 = $signed(_GEN_564) + $signed(_T_56266); // @[Modules.scala 143:103:@43926.4]
  assign _T_96216 = _T_96215[5:0]; // @[Modules.scala 143:103:@43927.4]
  assign _T_96217 = $signed(_T_96216); // @[Modules.scala 143:103:@43928.4]
  assign _GEN_974 = {{1{_T_62390[4]}},_T_62390}; // @[Modules.scala 143:103:@43938.4]
  assign _T_96229 = $signed(_GEN_974) + $signed(_T_56280); // @[Modules.scala 143:103:@43938.4]
  assign _T_96230 = _T_96229[5:0]; // @[Modules.scala 143:103:@43939.4]
  assign _T_96231 = $signed(_T_96230); // @[Modules.scala 143:103:@43940.4]
  assign buffer_13_0 = {{9{_T_94110[4]}},_T_94110}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_1 = {{9{_T_94117[4]}},_T_94117}; // @[Modules.scala 112:22:@8.4]
  assign _T_96253 = $signed(buffer_13_0) + $signed(buffer_13_1); // @[Modules.scala 166:64:@43960.4]
  assign _T_96254 = _T_96253[13:0]; // @[Modules.scala 166:64:@43961.4]
  assign buffer_13_307 = $signed(_T_96254); // @[Modules.scala 166:64:@43962.4]
  assign _T_96256 = $signed(buffer_3_2) + $signed(buffer_1_3); // @[Modules.scala 166:64:@43964.4]
  assign _T_96257 = _T_96256[13:0]; // @[Modules.scala 166:64:@43965.4]
  assign buffer_13_308 = $signed(_T_96257); // @[Modules.scala 166:64:@43966.4]
  assign buffer_13_5 = {{8{_T_94145[5]}},_T_94145}; // @[Modules.scala 112:22:@8.4]
  assign _T_96259 = $signed(buffer_2_4) + $signed(buffer_13_5); // @[Modules.scala 166:64:@43968.4]
  assign _T_96260 = _T_96259[13:0]; // @[Modules.scala 166:64:@43969.4]
  assign buffer_13_309 = $signed(_T_96260); // @[Modules.scala 166:64:@43970.4]
  assign buffer_13_6 = {{8{_T_94152[5]}},_T_94152}; // @[Modules.scala 112:22:@8.4]
  assign _T_96262 = $signed(buffer_13_6) + $signed(buffer_0_7); // @[Modules.scala 166:64:@43972.4]
  assign _T_96263 = _T_96262[13:0]; // @[Modules.scala 166:64:@43973.4]
  assign buffer_13_310 = $signed(_T_96263); // @[Modules.scala 166:64:@43974.4]
  assign buffer_13_8 = {{9{_T_94166[4]}},_T_94166}; // @[Modules.scala 112:22:@8.4]
  assign _T_96265 = $signed(buffer_13_8) + $signed(buffer_0_10); // @[Modules.scala 166:64:@43976.4]
  assign _T_96266 = _T_96265[13:0]; // @[Modules.scala 166:64:@43977.4]
  assign buffer_13_311 = $signed(_T_96266); // @[Modules.scala 166:64:@43978.4]
  assign buffer_13_10 = {{8{_T_94180[5]}},_T_94180}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_11 = {{9{_T_94187[4]}},_T_94187}; // @[Modules.scala 112:22:@8.4]
  assign _T_96268 = $signed(buffer_13_10) + $signed(buffer_13_11); // @[Modules.scala 166:64:@43980.4]
  assign _T_96269 = _T_96268[13:0]; // @[Modules.scala 166:64:@43981.4]
  assign buffer_13_312 = $signed(_T_96269); // @[Modules.scala 166:64:@43982.4]
  assign buffer_13_12 = {{8{_T_94194[5]}},_T_94194}; // @[Modules.scala 112:22:@8.4]
  assign _T_96271 = $signed(buffer_13_12) + $signed(buffer_0_14); // @[Modules.scala 166:64:@43984.4]
  assign _T_96272 = _T_96271[13:0]; // @[Modules.scala 166:64:@43985.4]
  assign buffer_13_313 = $signed(_T_96272); // @[Modules.scala 166:64:@43986.4]
  assign buffer_13_21 = {{8{_T_94257[5]}},_T_94257}; // @[Modules.scala 112:22:@8.4]
  assign _T_96283 = $signed(buffer_0_21) + $signed(buffer_13_21); // @[Modules.scala 166:64:@44000.4]
  assign _T_96284 = _T_96283[13:0]; // @[Modules.scala 166:64:@44001.4]
  assign buffer_13_317 = $signed(_T_96284); // @[Modules.scala 166:64:@44002.4]
  assign buffer_13_23 = {{8{_T_94271[5]}},_T_94271}; // @[Modules.scala 112:22:@8.4]
  assign _T_96286 = $signed(buffer_10_22) + $signed(buffer_13_23); // @[Modules.scala 166:64:@44004.4]
  assign _T_96287 = _T_96286[13:0]; // @[Modules.scala 166:64:@44005.4]
  assign buffer_13_318 = $signed(_T_96287); // @[Modules.scala 166:64:@44006.4]
  assign _T_96304 = $signed(buffer_2_32) + $signed(buffer_3_34); // @[Modules.scala 166:64:@44028.4]
  assign _T_96305 = _T_96304[13:0]; // @[Modules.scala 166:64:@44029.4]
  assign buffer_13_324 = $signed(_T_96305); // @[Modules.scala 166:64:@44030.4]
  assign buffer_13_36 = {{8{_T_94362[5]}},_T_94362}; // @[Modules.scala 112:22:@8.4]
  assign _T_96307 = $signed(buffer_13_36) + $signed(buffer_2_34); // @[Modules.scala 166:64:@44032.4]
  assign _T_96308 = _T_96307[13:0]; // @[Modules.scala 166:64:@44033.4]
  assign buffer_13_325 = $signed(_T_96308); // @[Modules.scala 166:64:@44034.4]
  assign _T_96310 = $signed(buffer_1_36) + $signed(buffer_2_36); // @[Modules.scala 166:64:@44036.4]
  assign _T_96311 = _T_96310[13:0]; // @[Modules.scala 166:64:@44037.4]
  assign buffer_13_326 = $signed(_T_96311); // @[Modules.scala 166:64:@44038.4]
  assign buffer_13_41 = {{8{_T_94397[5]}},_T_94397}; // @[Modules.scala 112:22:@8.4]
  assign _T_96313 = $signed(buffer_2_37) + $signed(buffer_13_41); // @[Modules.scala 166:64:@44040.4]
  assign _T_96314 = _T_96313[13:0]; // @[Modules.scala 166:64:@44041.4]
  assign buffer_13_327 = $signed(_T_96314); // @[Modules.scala 166:64:@44042.4]
  assign buffer_13_42 = {{8{_T_94404[5]}},_T_94404}; // @[Modules.scala 112:22:@8.4]
  assign _T_96316 = $signed(buffer_13_42) + $signed(buffer_5_43); // @[Modules.scala 166:64:@44044.4]
  assign _T_96317 = _T_96316[13:0]; // @[Modules.scala 166:64:@44045.4]
  assign buffer_13_328 = $signed(_T_96317); // @[Modules.scala 166:64:@44046.4]
  assign buffer_13_45 = {{8{_T_94425[5]}},_T_94425}; // @[Modules.scala 112:22:@8.4]
  assign _T_96319 = $signed(buffer_4_42) + $signed(buffer_13_45); // @[Modules.scala 166:64:@44048.4]
  assign _T_96320 = _T_96319[13:0]; // @[Modules.scala 166:64:@44049.4]
  assign buffer_13_329 = $signed(_T_96320); // @[Modules.scala 166:64:@44050.4]
  assign buffer_13_48 = {{8{_T_94446[5]}},_T_94446}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_49 = {{8{_T_94453[5]}},_T_94453}; // @[Modules.scala 112:22:@8.4]
  assign _T_96325 = $signed(buffer_13_48) + $signed(buffer_13_49); // @[Modules.scala 166:64:@44056.4]
  assign _T_96326 = _T_96325[13:0]; // @[Modules.scala 166:64:@44057.4]
  assign buffer_13_331 = $signed(_T_96326); // @[Modules.scala 166:64:@44058.4]
  assign _T_96331 = $signed(buffer_7_51) + $signed(buffer_12_46); // @[Modules.scala 166:64:@44064.4]
  assign _T_96332 = _T_96331[13:0]; // @[Modules.scala 166:64:@44065.4]
  assign buffer_13_333 = $signed(_T_96332); // @[Modules.scala 166:64:@44066.4]
  assign buffer_13_55 = {{9{_T_94495[4]}},_T_94495}; // @[Modules.scala 112:22:@8.4]
  assign _T_96334 = $signed(buffer_4_53) + $signed(buffer_13_55); // @[Modules.scala 166:64:@44068.4]
  assign _T_96335 = _T_96334[13:0]; // @[Modules.scala 166:64:@44069.4]
  assign buffer_13_334 = $signed(_T_96335); // @[Modules.scala 166:64:@44070.4]
  assign _T_96337 = $signed(buffer_10_56) + $signed(buffer_6_56); // @[Modules.scala 166:64:@44072.4]
  assign _T_96338 = _T_96337[13:0]; // @[Modules.scala 166:64:@44073.4]
  assign buffer_13_335 = $signed(_T_96338); // @[Modules.scala 166:64:@44074.4]
  assign _T_96340 = $signed(buffer_6_57) + $signed(buffer_6_58); // @[Modules.scala 166:64:@44076.4]
  assign _T_96341 = _T_96340[13:0]; // @[Modules.scala 166:64:@44077.4]
  assign buffer_13_336 = $signed(_T_96341); // @[Modules.scala 166:64:@44078.4]
  assign buffer_13_61 = {{8{_T_94537[5]}},_T_94537}; // @[Modules.scala 112:22:@8.4]
  assign _T_96343 = $signed(buffer_6_59) + $signed(buffer_13_61); // @[Modules.scala 166:64:@44080.4]
  assign _T_96344 = _T_96343[13:0]; // @[Modules.scala 166:64:@44081.4]
  assign buffer_13_337 = $signed(_T_96344); // @[Modules.scala 166:64:@44082.4]
  assign buffer_13_65 = {{9{_T_94565[4]}},_T_94565}; // @[Modules.scala 112:22:@8.4]
  assign _T_96349 = $signed(buffer_0_61) + $signed(buffer_13_65); // @[Modules.scala 166:64:@44088.4]
  assign _T_96350 = _T_96349[13:0]; // @[Modules.scala 166:64:@44089.4]
  assign buffer_13_339 = $signed(_T_96350); // @[Modules.scala 166:64:@44090.4]
  assign _T_96352 = $signed(buffer_10_64) + $signed(buffer_8_61); // @[Modules.scala 166:64:@44092.4]
  assign _T_96353 = _T_96352[13:0]; // @[Modules.scala 166:64:@44093.4]
  assign buffer_13_340 = $signed(_T_96353); // @[Modules.scala 166:64:@44094.4]
  assign _T_96355 = $signed(buffer_11_64) + $signed(buffer_5_69); // @[Modules.scala 166:64:@44096.4]
  assign _T_96356 = _T_96355[13:0]; // @[Modules.scala 166:64:@44097.4]
  assign buffer_13_341 = $signed(_T_96356); // @[Modules.scala 166:64:@44098.4]
  assign _T_96358 = $signed(buffer_6_69) + $signed(buffer_6_70); // @[Modules.scala 166:64:@44100.4]
  assign _T_96359 = _T_96358[13:0]; // @[Modules.scala 166:64:@44101.4]
  assign buffer_13_342 = $signed(_T_96359); // @[Modules.scala 166:64:@44102.4]
  assign buffer_13_73 = {{8{_T_94621[5]}},_T_94621}; // @[Modules.scala 112:22:@8.4]
  assign _T_96361 = $signed(buffer_6_71) + $signed(buffer_13_73); // @[Modules.scala 166:64:@44104.4]
  assign _T_96362 = _T_96361[13:0]; // @[Modules.scala 166:64:@44105.4]
  assign buffer_13_343 = $signed(_T_96362); // @[Modules.scala 166:64:@44106.4]
  assign buffer_13_74 = {{9{_T_94628[4]}},_T_94628}; // @[Modules.scala 112:22:@8.4]
  assign _T_96364 = $signed(buffer_13_74) + $signed(buffer_6_73); // @[Modules.scala 166:64:@44108.4]
  assign _T_96365 = _T_96364[13:0]; // @[Modules.scala 166:64:@44109.4]
  assign buffer_13_344 = $signed(_T_96365); // @[Modules.scala 166:64:@44110.4]
  assign buffer_13_77 = {{9{_T_94649[4]}},_T_94649}; // @[Modules.scala 112:22:@8.4]
  assign _T_96367 = $signed(buffer_9_77) + $signed(buffer_13_77); // @[Modules.scala 166:64:@44112.4]
  assign _T_96368 = _T_96367[13:0]; // @[Modules.scala 166:64:@44113.4]
  assign buffer_13_345 = $signed(_T_96368); // @[Modules.scala 166:64:@44114.4]
  assign buffer_13_79 = {{8{_T_94663[5]}},_T_94663}; // @[Modules.scala 112:22:@8.4]
  assign _T_96370 = $signed(buffer_3_78) + $signed(buffer_13_79); // @[Modules.scala 166:64:@44116.4]
  assign _T_96371 = _T_96370[13:0]; // @[Modules.scala 166:64:@44117.4]
  assign buffer_13_346 = $signed(_T_96371); // @[Modules.scala 166:64:@44118.4]
  assign buffer_13_81 = {{8{_T_94677[5]}},_T_94677}; // @[Modules.scala 112:22:@8.4]
  assign _T_96373 = $signed(buffer_4_78) + $signed(buffer_13_81); // @[Modules.scala 166:64:@44120.4]
  assign _T_96374 = _T_96373[13:0]; // @[Modules.scala 166:64:@44121.4]
  assign buffer_13_347 = $signed(_T_96374); // @[Modules.scala 166:64:@44122.4]
  assign buffer_13_84 = {{9{_T_94698[4]}},_T_94698}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_85 = {{9{_T_94705[4]}},_T_94705}; // @[Modules.scala 112:22:@8.4]
  assign _T_96379 = $signed(buffer_13_84) + $signed(buffer_13_85); // @[Modules.scala 166:64:@44128.4]
  assign _T_96380 = _T_96379[13:0]; // @[Modules.scala 166:64:@44129.4]
  assign buffer_13_349 = $signed(_T_96380); // @[Modules.scala 166:64:@44130.4]
  assign buffer_13_87 = {{9{_T_94719[4]}},_T_94719}; // @[Modules.scala 112:22:@8.4]
  assign _T_96382 = $signed(buffer_8_80) + $signed(buffer_13_87); // @[Modules.scala 166:64:@44132.4]
  assign _T_96383 = _T_96382[13:0]; // @[Modules.scala 166:64:@44133.4]
  assign buffer_13_350 = $signed(_T_96383); // @[Modules.scala 166:64:@44134.4]
  assign buffer_13_88 = {{8{_T_94726[5]}},_T_94726}; // @[Modules.scala 112:22:@8.4]
  assign _T_96385 = $signed(buffer_13_88) + $signed(buffer_0_85); // @[Modules.scala 166:64:@44136.4]
  assign _T_96386 = _T_96385[13:0]; // @[Modules.scala 166:64:@44137.4]
  assign buffer_13_351 = $signed(_T_96386); // @[Modules.scala 166:64:@44138.4]
  assign buffer_13_90 = {{8{_T_94740[5]}},_T_94740}; // @[Modules.scala 112:22:@8.4]
  assign _T_96388 = $signed(buffer_13_90) + $signed(buffer_0_87); // @[Modules.scala 166:64:@44140.4]
  assign _T_96389 = _T_96388[13:0]; // @[Modules.scala 166:64:@44141.4]
  assign buffer_13_352 = $signed(_T_96389); // @[Modules.scala 166:64:@44142.4]
  assign _T_96391 = $signed(buffer_3_93) + $signed(buffer_5_95); // @[Modules.scala 166:64:@44144.4]
  assign _T_96392 = _T_96391[13:0]; // @[Modules.scala 166:64:@44145.4]
  assign buffer_13_353 = $signed(_T_96392); // @[Modules.scala 166:64:@44146.4]
  assign buffer_13_95 = {{8{_T_94775[5]}},_T_94775}; // @[Modules.scala 112:22:@8.4]
  assign _T_96394 = $signed(buffer_5_96) + $signed(buffer_13_95); // @[Modules.scala 166:64:@44148.4]
  assign _T_96395 = _T_96394[13:0]; // @[Modules.scala 166:64:@44149.4]
  assign buffer_13_354 = $signed(_T_96395); // @[Modules.scala 166:64:@44150.4]
  assign buffer_13_96 = {{9{_T_94782[4]}},_T_94782}; // @[Modules.scala 112:22:@8.4]
  assign _T_96397 = $signed(buffer_13_96) + $signed(buffer_2_97); // @[Modules.scala 166:64:@44152.4]
  assign _T_96398 = _T_96397[13:0]; // @[Modules.scala 166:64:@44153.4]
  assign buffer_13_355 = $signed(_T_96398); // @[Modules.scala 166:64:@44154.4]
  assign buffer_13_103 = {{8{_T_94831[5]}},_T_94831}; // @[Modules.scala 112:22:@8.4]
  assign _T_96406 = $signed(buffer_0_97) + $signed(buffer_13_103); // @[Modules.scala 166:64:@44164.4]
  assign _T_96407 = _T_96406[13:0]; // @[Modules.scala 166:64:@44165.4]
  assign buffer_13_358 = $signed(_T_96407); // @[Modules.scala 166:64:@44166.4]
  assign buffer_13_104 = {{9{_T_94838[4]}},_T_94838}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_105 = {{8{_T_94845[5]}},_T_94845}; // @[Modules.scala 112:22:@8.4]
  assign _T_96409 = $signed(buffer_13_104) + $signed(buffer_13_105); // @[Modules.scala 166:64:@44168.4]
  assign _T_96410 = _T_96409[13:0]; // @[Modules.scala 166:64:@44169.4]
  assign buffer_13_359 = $signed(_T_96410); // @[Modules.scala 166:64:@44170.4]
  assign buffer_13_106 = {{8{_T_94852[5]}},_T_94852}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_107 = {{8{_T_94859[5]}},_T_94859}; // @[Modules.scala 112:22:@8.4]
  assign _T_96412 = $signed(buffer_13_106) + $signed(buffer_13_107); // @[Modules.scala 166:64:@44172.4]
  assign _T_96413 = _T_96412[13:0]; // @[Modules.scala 166:64:@44173.4]
  assign buffer_13_360 = $signed(_T_96413); // @[Modules.scala 166:64:@44174.4]
  assign buffer_13_108 = {{9{_T_94866[4]}},_T_94866}; // @[Modules.scala 112:22:@8.4]
  assign _T_96415 = $signed(buffer_13_108) + $signed(buffer_9_113); // @[Modules.scala 166:64:@44176.4]
  assign _T_96416 = _T_96415[13:0]; // @[Modules.scala 166:64:@44177.4]
  assign buffer_13_361 = $signed(_T_96416); // @[Modules.scala 166:64:@44178.4]
  assign buffer_13_112 = {{8{_T_94894[5]}},_T_94894}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_113 = {{8{_T_94901[5]}},_T_94901}; // @[Modules.scala 112:22:@8.4]
  assign _T_96421 = $signed(buffer_13_112) + $signed(buffer_13_113); // @[Modules.scala 166:64:@44184.4]
  assign _T_96422 = _T_96421[13:0]; // @[Modules.scala 166:64:@44185.4]
  assign buffer_13_363 = $signed(_T_96422); // @[Modules.scala 166:64:@44186.4]
  assign buffer_13_115 = {{8{_T_94915[5]}},_T_94915}; // @[Modules.scala 112:22:@8.4]
  assign _T_96424 = $signed(buffer_0_111) + $signed(buffer_13_115); // @[Modules.scala 166:64:@44188.4]
  assign _T_96425 = _T_96424[13:0]; // @[Modules.scala 166:64:@44189.4]
  assign buffer_13_364 = $signed(_T_96425); // @[Modules.scala 166:64:@44190.4]
  assign buffer_13_116 = {{8{_T_94922[5]}},_T_94922}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_117 = {{9{_T_94929[4]}},_T_94929}; // @[Modules.scala 112:22:@8.4]
  assign _T_96427 = $signed(buffer_13_116) + $signed(buffer_13_117); // @[Modules.scala 166:64:@44192.4]
  assign _T_96428 = _T_96427[13:0]; // @[Modules.scala 166:64:@44193.4]
  assign buffer_13_365 = $signed(_T_96428); // @[Modules.scala 166:64:@44194.4]
  assign buffer_13_121 = {{9{_T_94957[4]}},_T_94957}; // @[Modules.scala 112:22:@8.4]
  assign _T_96433 = $signed(buffer_7_120) + $signed(buffer_13_121); // @[Modules.scala 166:64:@44200.4]
  assign _T_96434 = _T_96433[13:0]; // @[Modules.scala 166:64:@44201.4]
  assign buffer_13_367 = $signed(_T_96434); // @[Modules.scala 166:64:@44202.4]
  assign buffer_13_122 = {{8{_T_94964[5]}},_T_94964}; // @[Modules.scala 112:22:@8.4]
  assign _T_96436 = $signed(buffer_13_122) + $signed(buffer_10_123); // @[Modules.scala 166:64:@44204.4]
  assign _T_96437 = _T_96436[13:0]; // @[Modules.scala 166:64:@44205.4]
  assign buffer_13_368 = $signed(_T_96437); // @[Modules.scala 166:64:@44206.4]
  assign buffer_13_124 = {{8{_T_94978[5]}},_T_94978}; // @[Modules.scala 112:22:@8.4]
  assign _T_96439 = $signed(buffer_13_124) + $signed(buffer_1_126); // @[Modules.scala 166:64:@44208.4]
  assign _T_96440 = _T_96439[13:0]; // @[Modules.scala 166:64:@44209.4]
  assign buffer_13_369 = $signed(_T_96440); // @[Modules.scala 166:64:@44210.4]
  assign buffer_13_126 = {{8{_T_94992[5]}},_T_94992}; // @[Modules.scala 112:22:@8.4]
  assign _T_96442 = $signed(buffer_13_126) + $signed(buffer_2_129); // @[Modules.scala 166:64:@44212.4]
  assign _T_96443 = _T_96442[13:0]; // @[Modules.scala 166:64:@44213.4]
  assign buffer_13_370 = $signed(_T_96443); // @[Modules.scala 166:64:@44214.4]
  assign _T_96445 = $signed(buffer_0_127) + $signed(buffer_0_128); // @[Modules.scala 166:64:@44216.4]
  assign _T_96446 = _T_96445[13:0]; // @[Modules.scala 166:64:@44217.4]
  assign buffer_13_371 = $signed(_T_96446); // @[Modules.scala 166:64:@44218.4]
  assign _T_96448 = $signed(buffer_0_129) + $signed(buffer_2_133); // @[Modules.scala 166:64:@44220.4]
  assign _T_96449 = _T_96448[13:0]; // @[Modules.scala 166:64:@44221.4]
  assign buffer_13_372 = $signed(_T_96449); // @[Modules.scala 166:64:@44222.4]
  assign buffer_13_132 = {{8{_T_95034[5]}},_T_95034}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_133 = {{9{_T_95041[4]}},_T_95041}; // @[Modules.scala 112:22:@8.4]
  assign _T_96451 = $signed(buffer_13_132) + $signed(buffer_13_133); // @[Modules.scala 166:64:@44224.4]
  assign _T_96452 = _T_96451[13:0]; // @[Modules.scala 166:64:@44225.4]
  assign buffer_13_373 = $signed(_T_96452); // @[Modules.scala 166:64:@44226.4]
  assign buffer_13_135 = {{8{_T_95055[5]}},_T_95055}; // @[Modules.scala 112:22:@8.4]
  assign _T_96454 = $signed(buffer_4_133) + $signed(buffer_13_135); // @[Modules.scala 166:64:@44228.4]
  assign _T_96455 = _T_96454[13:0]; // @[Modules.scala 166:64:@44229.4]
  assign buffer_13_374 = $signed(_T_96455); // @[Modules.scala 166:64:@44230.4]
  assign _T_96457 = $signed(buffer_3_144) + $signed(buffer_0_138); // @[Modules.scala 166:64:@44232.4]
  assign _T_96458 = _T_96457[13:0]; // @[Modules.scala 166:64:@44233.4]
  assign buffer_13_375 = $signed(_T_96458); // @[Modules.scala 166:64:@44234.4]
  assign buffer_13_138 = {{8{_T_95076[5]}},_T_95076}; // @[Modules.scala 112:22:@8.4]
  assign _T_96460 = $signed(buffer_13_138) + $signed(buffer_0_140); // @[Modules.scala 166:64:@44236.4]
  assign _T_96461 = _T_96460[13:0]; // @[Modules.scala 166:64:@44237.4]
  assign buffer_13_376 = $signed(_T_96461); // @[Modules.scala 166:64:@44238.4]
  assign buffer_13_142 = {{8{_T_95104[5]}},_T_95104}; // @[Modules.scala 112:22:@8.4]
  assign _T_96466 = $signed(buffer_13_142) + $signed(buffer_2_147); // @[Modules.scala 166:64:@44244.4]
  assign _T_96467 = _T_96466[13:0]; // @[Modules.scala 166:64:@44245.4]
  assign buffer_13_378 = $signed(_T_96467); // @[Modules.scala 166:64:@44246.4]
  assign buffer_13_145 = {{8{_T_95125[5]}},_T_95125}; // @[Modules.scala 112:22:@8.4]
  assign _T_96469 = $signed(buffer_1_146) + $signed(buffer_13_145); // @[Modules.scala 166:64:@44248.4]
  assign _T_96470 = _T_96469[13:0]; // @[Modules.scala 166:64:@44249.4]
  assign buffer_13_379 = $signed(_T_96470); // @[Modules.scala 166:64:@44250.4]
  assign buffer_13_146 = {{8{_T_95132[5]}},_T_95132}; // @[Modules.scala 112:22:@8.4]
  assign _T_96472 = $signed(buffer_13_146) + $signed(buffer_10_151); // @[Modules.scala 166:64:@44252.4]
  assign _T_96473 = _T_96472[13:0]; // @[Modules.scala 166:64:@44253.4]
  assign buffer_13_380 = $signed(_T_96473); // @[Modules.scala 166:64:@44254.4]
  assign buffer_13_149 = {{8{_T_95153[5]}},_T_95153}; // @[Modules.scala 112:22:@8.4]
  assign _T_96475 = $signed(buffer_5_150) + $signed(buffer_13_149); // @[Modules.scala 166:64:@44256.4]
  assign _T_96476 = _T_96475[13:0]; // @[Modules.scala 166:64:@44257.4]
  assign buffer_13_381 = $signed(_T_96476); // @[Modules.scala 166:64:@44258.4]
  assign _T_96478 = $signed(buffer_0_151) + $signed(buffer_0_152); // @[Modules.scala 166:64:@44260.4]
  assign _T_96479 = _T_96478[13:0]; // @[Modules.scala 166:64:@44261.4]
  assign buffer_13_382 = $signed(_T_96479); // @[Modules.scala 166:64:@44262.4]
  assign buffer_13_152 = {{9{_T_95174[4]}},_T_95174}; // @[Modules.scala 112:22:@8.4]
  assign _T_96481 = $signed(buffer_13_152) + $signed(buffer_2_159); // @[Modules.scala 166:64:@44264.4]
  assign _T_96482 = _T_96481[13:0]; // @[Modules.scala 166:64:@44265.4]
  assign buffer_13_383 = $signed(_T_96482); // @[Modules.scala 166:64:@44266.4]
  assign _T_96484 = $signed(buffer_2_160) + $signed(buffer_1_157); // @[Modules.scala 166:64:@44268.4]
  assign _T_96485 = _T_96484[13:0]; // @[Modules.scala 166:64:@44269.4]
  assign buffer_13_384 = $signed(_T_96485); // @[Modules.scala 166:64:@44270.4]
  assign _T_96487 = $signed(buffer_8_155) + $signed(buffer_8_156); // @[Modules.scala 166:64:@44272.4]
  assign _T_96488 = _T_96487[13:0]; // @[Modules.scala 166:64:@44273.4]
  assign buffer_13_385 = $signed(_T_96488); // @[Modules.scala 166:64:@44274.4]
  assign buffer_13_158 = {{9{_T_95216[4]}},_T_95216}; // @[Modules.scala 112:22:@8.4]
  assign _T_96490 = $signed(buffer_13_158) + $signed(buffer_1_160); // @[Modules.scala 166:64:@44276.4]
  assign _T_96491 = _T_96490[13:0]; // @[Modules.scala 166:64:@44277.4]
  assign buffer_13_386 = $signed(_T_96491); // @[Modules.scala 166:64:@44278.4]
  assign buffer_13_160 = {{8{_T_95230[5]}},_T_95230}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_161 = {{8{_T_95237[5]}},_T_95237}; // @[Modules.scala 112:22:@8.4]
  assign _T_96493 = $signed(buffer_13_160) + $signed(buffer_13_161); // @[Modules.scala 166:64:@44280.4]
  assign _T_96494 = _T_96493[13:0]; // @[Modules.scala 166:64:@44281.4]
  assign buffer_13_387 = $signed(_T_96494); // @[Modules.scala 166:64:@44282.4]
  assign buffer_13_162 = {{8{_T_95244[5]}},_T_95244}; // @[Modules.scala 112:22:@8.4]
  assign _T_96496 = $signed(buffer_13_162) + $signed(buffer_9_169); // @[Modules.scala 166:64:@44284.4]
  assign _T_96497 = _T_96496[13:0]; // @[Modules.scala 166:64:@44285.4]
  assign buffer_13_388 = $signed(_T_96497); // @[Modules.scala 166:64:@44286.4]
  assign buffer_13_166 = {{8{_T_95272[5]}},_T_95272}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_167 = {{8{_T_95279[5]}},_T_95279}; // @[Modules.scala 112:22:@8.4]
  assign _T_96502 = $signed(buffer_13_166) + $signed(buffer_13_167); // @[Modules.scala 166:64:@44292.4]
  assign _T_96503 = _T_96502[13:0]; // @[Modules.scala 166:64:@44293.4]
  assign buffer_13_390 = $signed(_T_96503); // @[Modules.scala 166:64:@44294.4]
  assign buffer_13_171 = {{8{_T_95307[5]}},_T_95307}; // @[Modules.scala 112:22:@8.4]
  assign _T_96508 = $signed(buffer_8_167) + $signed(buffer_13_171); // @[Modules.scala 166:64:@44300.4]
  assign _T_96509 = _T_96508[13:0]; // @[Modules.scala 166:64:@44301.4]
  assign buffer_13_392 = $signed(_T_96509); // @[Modules.scala 166:64:@44302.4]
  assign buffer_13_172 = {{9{_T_95314[4]}},_T_95314}; // @[Modules.scala 112:22:@8.4]
  assign _T_96511 = $signed(buffer_13_172) + $signed(buffer_0_172); // @[Modules.scala 166:64:@44304.4]
  assign _T_96512 = _T_96511[13:0]; // @[Modules.scala 166:64:@44305.4]
  assign buffer_13_393 = $signed(_T_96512); // @[Modules.scala 166:64:@44306.4]
  assign buffer_13_174 = {{8{_T_95328[5]}},_T_95328}; // @[Modules.scala 112:22:@8.4]
  assign _T_96514 = $signed(buffer_13_174) + $signed(buffer_3_181); // @[Modules.scala 166:64:@44308.4]
  assign _T_96515 = _T_96514[13:0]; // @[Modules.scala 166:64:@44309.4]
  assign buffer_13_394 = $signed(_T_96515); // @[Modules.scala 166:64:@44310.4]
  assign _T_96517 = $signed(buffer_1_175) + $signed(buffer_0_177); // @[Modules.scala 166:64:@44312.4]
  assign _T_96518 = _T_96517[13:0]; // @[Modules.scala 166:64:@44313.4]
  assign buffer_13_395 = $signed(_T_96518); // @[Modules.scala 166:64:@44314.4]
  assign _T_96520 = $signed(buffer_0_178) + $signed(buffer_6_185); // @[Modules.scala 166:64:@44316.4]
  assign _T_96521 = _T_96520[13:0]; // @[Modules.scala 166:64:@44317.4]
  assign buffer_13_396 = $signed(_T_96521); // @[Modules.scala 166:64:@44318.4]
  assign buffer_13_181 = {{8{_T_95377[5]}},_T_95377}; // @[Modules.scala 112:22:@8.4]
  assign _T_96523 = $signed(buffer_8_180) + $signed(buffer_13_181); // @[Modules.scala 166:64:@44320.4]
  assign _T_96524 = _T_96523[13:0]; // @[Modules.scala 166:64:@44321.4]
  assign buffer_13_397 = $signed(_T_96524); // @[Modules.scala 166:64:@44322.4]
  assign buffer_13_183 = {{8{_T_95391[5]}},_T_95391}; // @[Modules.scala 112:22:@8.4]
  assign _T_96526 = $signed(buffer_2_187) + $signed(buffer_13_183); // @[Modules.scala 166:64:@44324.4]
  assign _T_96527 = _T_96526[13:0]; // @[Modules.scala 166:64:@44325.4]
  assign buffer_13_398 = $signed(_T_96527); // @[Modules.scala 166:64:@44326.4]
  assign buffer_13_186 = {{8{_T_95412[5]}},_T_95412}; // @[Modules.scala 112:22:@8.4]
  assign _T_96532 = $signed(buffer_13_186) + $signed(buffer_6_195); // @[Modules.scala 166:64:@44332.4]
  assign _T_96533 = _T_96532[13:0]; // @[Modules.scala 166:64:@44333.4]
  assign buffer_13_400 = $signed(_T_96533); // @[Modules.scala 166:64:@44334.4]
  assign buffer_13_192 = {{8{_T_95454[5]}},_T_95454}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_193 = {{8{_T_95461[5]}},_T_95461}; // @[Modules.scala 112:22:@8.4]
  assign _T_96541 = $signed(buffer_13_192) + $signed(buffer_13_193); // @[Modules.scala 166:64:@44344.4]
  assign _T_96542 = _T_96541[13:0]; // @[Modules.scala 166:64:@44345.4]
  assign buffer_13_403 = $signed(_T_96542); // @[Modules.scala 166:64:@44346.4]
  assign _T_96544 = $signed(buffer_4_185) + $signed(buffer_0_192); // @[Modules.scala 166:64:@44348.4]
  assign _T_96545 = _T_96544[13:0]; // @[Modules.scala 166:64:@44349.4]
  assign buffer_13_404 = $signed(_T_96545); // @[Modules.scala 166:64:@44350.4]
  assign buffer_13_198 = {{9{_T_95496[4]}},_T_95496}; // @[Modules.scala 112:22:@8.4]
  assign _T_96550 = $signed(buffer_13_198) + $signed(buffer_9_207); // @[Modules.scala 166:64:@44356.4]
  assign _T_96551 = _T_96550[13:0]; // @[Modules.scala 166:64:@44357.4]
  assign buffer_13_406 = $signed(_T_96551); // @[Modules.scala 166:64:@44358.4]
  assign buffer_13_200 = {{8{_T_95510[5]}},_T_95510}; // @[Modules.scala 112:22:@8.4]
  assign _T_96553 = $signed(buffer_13_200) + $signed(buffer_2_204); // @[Modules.scala 166:64:@44360.4]
  assign _T_96554 = _T_96553[13:0]; // @[Modules.scala 166:64:@44361.4]
  assign buffer_13_407 = $signed(_T_96554); // @[Modules.scala 166:64:@44362.4]
  assign buffer_13_204 = {{8{_T_95538[5]}},_T_95538}; // @[Modules.scala 112:22:@8.4]
  assign _T_96559 = $signed(buffer_13_204) + $signed(buffer_0_205); // @[Modules.scala 166:64:@44368.4]
  assign _T_96560 = _T_96559[13:0]; // @[Modules.scala 166:64:@44369.4]
  assign buffer_13_409 = $signed(_T_96560); // @[Modules.scala 166:64:@44370.4]
  assign _T_96562 = $signed(buffer_11_204) + $signed(buffer_3_217); // @[Modules.scala 166:64:@44372.4]
  assign _T_96563 = _T_96562[13:0]; // @[Modules.scala 166:64:@44373.4]
  assign buffer_13_410 = $signed(_T_96563); // @[Modules.scala 166:64:@44374.4]
  assign buffer_13_209 = {{8{_T_95573[5]}},_T_95573}; // @[Modules.scala 112:22:@8.4]
  assign _T_96565 = $signed(buffer_0_208) + $signed(buffer_13_209); // @[Modules.scala 166:64:@44376.4]
  assign _T_96566 = _T_96565[13:0]; // @[Modules.scala 166:64:@44377.4]
  assign buffer_13_411 = $signed(_T_96566); // @[Modules.scala 166:64:@44378.4]
  assign buffer_13_210 = {{8{_T_95580[5]}},_T_95580}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_211 = {{8{_T_95587[5]}},_T_95587}; // @[Modules.scala 112:22:@8.4]
  assign _T_96568 = $signed(buffer_13_210) + $signed(buffer_13_211); // @[Modules.scala 166:64:@44380.4]
  assign _T_96569 = _T_96568[13:0]; // @[Modules.scala 166:64:@44381.4]
  assign buffer_13_412 = $signed(_T_96569); // @[Modules.scala 166:64:@44382.4]
  assign buffer_13_212 = {{8{_T_95594[5]}},_T_95594}; // @[Modules.scala 112:22:@8.4]
  assign _T_96571 = $signed(buffer_13_212) + $signed(buffer_6_223); // @[Modules.scala 166:64:@44384.4]
  assign _T_96572 = _T_96571[13:0]; // @[Modules.scala 166:64:@44385.4]
  assign buffer_13_413 = $signed(_T_96572); // @[Modules.scala 166:64:@44386.4]
  assign buffer_13_216 = {{8{_T_95622[5]}},_T_95622}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_217 = {{8{_T_95629[5]}},_T_95629}; // @[Modules.scala 112:22:@8.4]
  assign _T_96577 = $signed(buffer_13_216) + $signed(buffer_13_217); // @[Modules.scala 166:64:@44392.4]
  assign _T_96578 = _T_96577[13:0]; // @[Modules.scala 166:64:@44393.4]
  assign buffer_13_415 = $signed(_T_96578); // @[Modules.scala 166:64:@44394.4]
  assign _T_96580 = $signed(buffer_6_228) + $signed(buffer_5_222); // @[Modules.scala 166:64:@44396.4]
  assign _T_96581 = _T_96580[13:0]; // @[Modules.scala 166:64:@44397.4]
  assign buffer_13_416 = $signed(_T_96581); // @[Modules.scala 166:64:@44398.4]
  assign _T_96589 = $signed(buffer_2_228) + $signed(buffer_6_236); // @[Modules.scala 166:64:@44408.4]
  assign _T_96590 = _T_96589[13:0]; // @[Modules.scala 166:64:@44409.4]
  assign buffer_13_419 = $signed(_T_96590); // @[Modules.scala 166:64:@44410.4]
  assign _T_96592 = $signed(buffer_5_230) + $signed(buffer_10_231); // @[Modules.scala 166:64:@44412.4]
  assign _T_96593 = _T_96592[13:0]; // @[Modules.scala 166:64:@44413.4]
  assign buffer_13_420 = $signed(_T_96593); // @[Modules.scala 166:64:@44414.4]
  assign buffer_13_228 = {{8{_T_95706[5]}},_T_95706}; // @[Modules.scala 112:22:@8.4]
  assign _T_96595 = $signed(buffer_13_228) + $signed(buffer_7_238); // @[Modules.scala 166:64:@44416.4]
  assign _T_96596 = _T_96595[13:0]; // @[Modules.scala 166:64:@44417.4]
  assign buffer_13_421 = $signed(_T_96596); // @[Modules.scala 166:64:@44418.4]
  assign _T_96598 = $signed(buffer_9_238) + $signed(buffer_6_241); // @[Modules.scala 166:64:@44420.4]
  assign _T_96599 = _T_96598[13:0]; // @[Modules.scala 166:64:@44421.4]
  assign buffer_13_422 = $signed(_T_96599); // @[Modules.scala 166:64:@44422.4]
  assign _T_96601 = $signed(buffer_0_229) + $signed(buffer_1_232); // @[Modules.scala 166:64:@44424.4]
  assign _T_96602 = _T_96601[13:0]; // @[Modules.scala 166:64:@44425.4]
  assign buffer_13_423 = $signed(_T_96602); // @[Modules.scala 166:64:@44426.4]
  assign buffer_13_234 = {{8{_T_95748[5]}},_T_95748}; // @[Modules.scala 112:22:@8.4]
  assign _T_96604 = $signed(buffer_13_234) + $signed(buffer_5_240); // @[Modules.scala 166:64:@44428.4]
  assign _T_96605 = _T_96604[13:0]; // @[Modules.scala 166:64:@44429.4]
  assign buffer_13_424 = $signed(_T_96605); // @[Modules.scala 166:64:@44430.4]
  assign _T_96607 = $signed(buffer_12_230) + $signed(buffer_6_245); // @[Modules.scala 166:64:@44432.4]
  assign _T_96608 = _T_96607[13:0]; // @[Modules.scala 166:64:@44433.4]
  assign buffer_13_425 = $signed(_T_96608); // @[Modules.scala 166:64:@44434.4]
  assign buffer_13_239 = {{8{_T_95783[5]}},_T_95783}; // @[Modules.scala 112:22:@8.4]
  assign _T_96610 = $signed(buffer_6_246) + $signed(buffer_13_239); // @[Modules.scala 166:64:@44436.4]
  assign _T_96611 = _T_96610[13:0]; // @[Modules.scala 166:64:@44437.4]
  assign buffer_13_426 = $signed(_T_96611); // @[Modules.scala 166:64:@44438.4]
  assign _T_96613 = $signed(buffer_0_235) + $signed(buffer_1_239); // @[Modules.scala 166:64:@44440.4]
  assign _T_96614 = _T_96613[13:0]; // @[Modules.scala 166:64:@44441.4]
  assign buffer_13_427 = $signed(_T_96614); // @[Modules.scala 166:64:@44442.4]
  assign buffer_13_245 = {{8{_T_95825[5]}},_T_95825}; // @[Modules.scala 112:22:@8.4]
  assign _T_96619 = $signed(buffer_8_250) + $signed(buffer_13_245); // @[Modules.scala 166:64:@44448.4]
  assign _T_96620 = _T_96619[13:0]; // @[Modules.scala 166:64:@44449.4]
  assign buffer_13_429 = $signed(_T_96620); // @[Modules.scala 166:64:@44450.4]
  assign _T_96622 = $signed(buffer_12_239) + $signed(buffer_8_253); // @[Modules.scala 166:64:@44452.4]
  assign _T_96623 = _T_96622[13:0]; // @[Modules.scala 166:64:@44453.4]
  assign buffer_13_430 = $signed(_T_96623); // @[Modules.scala 166:64:@44454.4]
  assign buffer_13_248 = {{8{_T_95846[5]}},_T_95846}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_249 = {{8{_T_95853[5]}},_T_95853}; // @[Modules.scala 112:22:@8.4]
  assign _T_96625 = $signed(buffer_13_248) + $signed(buffer_13_249); // @[Modules.scala 166:64:@44456.4]
  assign _T_96626 = _T_96625[13:0]; // @[Modules.scala 166:64:@44457.4]
  assign buffer_13_431 = $signed(_T_96626); // @[Modules.scala 166:64:@44458.4]
  assign _T_96631 = $signed(buffer_0_249) + $signed(buffer_0_250); // @[Modules.scala 166:64:@44464.4]
  assign _T_96632 = _T_96631[13:0]; // @[Modules.scala 166:64:@44465.4]
  assign buffer_13_433 = $signed(_T_96632); // @[Modules.scala 166:64:@44466.4]
  assign buffer_13_255 = {{8{_T_95895[5]}},_T_95895}; // @[Modules.scala 112:22:@8.4]
  assign _T_96634 = $signed(buffer_2_258) + $signed(buffer_13_255); // @[Modules.scala 166:64:@44468.4]
  assign _T_96635 = _T_96634[13:0]; // @[Modules.scala 166:64:@44469.4]
  assign buffer_13_434 = $signed(_T_96635); // @[Modules.scala 166:64:@44470.4]
  assign buffer_13_256 = {{8{_T_95902[5]}},_T_95902}; // @[Modules.scala 112:22:@8.4]
  assign buffer_13_257 = {{8{_T_95909[5]}},_T_95909}; // @[Modules.scala 112:22:@8.4]
  assign _T_96637 = $signed(buffer_13_256) + $signed(buffer_13_257); // @[Modules.scala 166:64:@44472.4]
  assign _T_96638 = _T_96637[13:0]; // @[Modules.scala 166:64:@44473.4]
  assign buffer_13_435 = $signed(_T_96638); // @[Modules.scala 166:64:@44474.4]
  assign buffer_13_259 = {{8{_T_95923[5]}},_T_95923}; // @[Modules.scala 112:22:@8.4]
  assign _T_96640 = $signed(buffer_3_264) + $signed(buffer_13_259); // @[Modules.scala 166:64:@44476.4]
  assign _T_96641 = _T_96640[13:0]; // @[Modules.scala 166:64:@44477.4]
  assign buffer_13_436 = $signed(_T_96641); // @[Modules.scala 166:64:@44478.4]
  assign _T_96643 = $signed(buffer_12_253) + $signed(buffer_10_263); // @[Modules.scala 166:64:@44480.4]
  assign _T_96644 = _T_96643[13:0]; // @[Modules.scala 166:64:@44481.4]
  assign buffer_13_437 = $signed(_T_96644); // @[Modules.scala 166:64:@44482.4]
  assign _T_96652 = $signed(buffer_3_272) + $signed(buffer_2_272); // @[Modules.scala 166:64:@44492.4]
  assign _T_96653 = _T_96652[13:0]; // @[Modules.scala 166:64:@44493.4]
  assign buffer_13_440 = $signed(_T_96653); // @[Modules.scala 166:64:@44494.4]
  assign buffer_13_269 = {{8{_T_95993[5]}},_T_95993}; // @[Modules.scala 112:22:@8.4]
  assign _T_96655 = $signed(buffer_12_261) + $signed(buffer_13_269); // @[Modules.scala 166:64:@44496.4]
  assign _T_96656 = _T_96655[13:0]; // @[Modules.scala 166:64:@44497.4]
  assign buffer_13_441 = $signed(_T_96656); // @[Modules.scala 166:64:@44498.4]
  assign buffer_13_270 = {{8{_T_96000[5]}},_T_96000}; // @[Modules.scala 112:22:@8.4]
  assign _T_96658 = $signed(buffer_13_270) + $signed(buffer_12_263); // @[Modules.scala 166:64:@44500.4]
  assign _T_96659 = _T_96658[13:0]; // @[Modules.scala 166:64:@44501.4]
  assign buffer_13_442 = $signed(_T_96659); // @[Modules.scala 166:64:@44502.4]
  assign _T_96661 = $signed(buffer_6_279) + $signed(buffer_6_280); // @[Modules.scala 166:64:@44504.4]
  assign _T_96662 = _T_96661[13:0]; // @[Modules.scala 166:64:@44505.4]
  assign buffer_13_443 = $signed(_T_96662); // @[Modules.scala 166:64:@44506.4]
  assign _T_96664 = $signed(buffer_1_270) + $signed(buffer_3_281); // @[Modules.scala 166:64:@44508.4]
  assign _T_96665 = _T_96664[13:0]; // @[Modules.scala 166:64:@44509.4]
  assign buffer_13_444 = $signed(_T_96665); // @[Modules.scala 166:64:@44510.4]
  assign _T_96667 = $signed(buffer_11_267) + $signed(buffer_2_280); // @[Modules.scala 166:64:@44512.4]
  assign _T_96668 = _T_96667[13:0]; // @[Modules.scala 166:64:@44513.4]
  assign buffer_13_445 = $signed(_T_96668); // @[Modules.scala 166:64:@44514.4]
  assign _T_96670 = $signed(buffer_7_281) + $signed(buffer_11_270); // @[Modules.scala 166:64:@44516.4]
  assign _T_96671 = _T_96670[13:0]; // @[Modules.scala 166:64:@44517.4]
  assign buffer_13_446 = $signed(_T_96671); // @[Modules.scala 166:64:@44518.4]
  assign buffer_13_281 = {{9{_T_96077[4]}},_T_96077}; // @[Modules.scala 112:22:@8.4]
  assign _T_96673 = $signed(buffer_11_271) + $signed(buffer_13_281); // @[Modules.scala 166:64:@44520.4]
  assign _T_96674 = _T_96673[13:0]; // @[Modules.scala 166:64:@44521.4]
  assign buffer_13_447 = $signed(_T_96674); // @[Modules.scala 166:64:@44522.4]
  assign _T_96685 = $signed(buffer_2_289) + $signed(buffer_1_283); // @[Modules.scala 166:64:@44536.4]
  assign _T_96686 = _T_96685[13:0]; // @[Modules.scala 166:64:@44537.4]
  assign buffer_13_451 = $signed(_T_96686); // @[Modules.scala 166:64:@44538.4]
  assign buffer_13_290 = {{9{_T_96140[4]}},_T_96140}; // @[Modules.scala 112:22:@8.4]
  assign _T_96688 = $signed(buffer_13_290) + $signed(buffer_9_296); // @[Modules.scala 166:64:@44540.4]
  assign _T_96689 = _T_96688[13:0]; // @[Modules.scala 166:64:@44541.4]
  assign buffer_13_452 = $signed(_T_96689); // @[Modules.scala 166:64:@44542.4]
  assign _T_96691 = $signed(buffer_9_297) + $signed(buffer_9_298); // @[Modules.scala 166:64:@44544.4]
  assign _T_96692 = _T_96691[13:0]; // @[Modules.scala 166:64:@44545.4]
  assign buffer_13_453 = $signed(_T_96692); // @[Modules.scala 166:64:@44546.4]
  assign _T_96694 = $signed(buffer_9_299) + $signed(buffer_9_300); // @[Modules.scala 166:64:@44548.4]
  assign _T_96695 = _T_96694[13:0]; // @[Modules.scala 166:64:@44549.4]
  assign buffer_13_454 = $signed(_T_96695); // @[Modules.scala 166:64:@44550.4]
  assign _T_96697 = $signed(buffer_9_301) + $signed(buffer_6_304); // @[Modules.scala 166:64:@44552.4]
  assign _T_96698 = _T_96697[13:0]; // @[Modules.scala 166:64:@44553.4]
  assign buffer_13_455 = $signed(_T_96698); // @[Modules.scala 166:64:@44554.4]
  assign _T_96700 = $signed(buffer_10_298) + $signed(buffer_5_304); // @[Modules.scala 166:64:@44556.4]
  assign _T_96701 = _T_96700[13:0]; // @[Modules.scala 166:64:@44557.4]
  assign buffer_13_456 = $signed(_T_96701); // @[Modules.scala 166:64:@44558.4]
  assign buffer_13_301 = {{8{_T_96217[5]}},_T_96217}; // @[Modules.scala 112:22:@8.4]
  assign _T_96703 = $signed(buffer_12_289) + $signed(buffer_13_301); // @[Modules.scala 166:64:@44560.4]
  assign _T_96704 = _T_96703[13:0]; // @[Modules.scala 166:64:@44561.4]
  assign buffer_13_457 = $signed(_T_96704); // @[Modules.scala 166:64:@44562.4]
  assign buffer_13_303 = {{8{_T_96231[5]}},_T_96231}; // @[Modules.scala 112:22:@8.4]
  assign _T_96706 = $signed(buffer_7_303) + $signed(buffer_13_303); // @[Modules.scala 166:64:@44564.4]
  assign _T_96707 = _T_96706[13:0]; // @[Modules.scala 166:64:@44565.4]
  assign buffer_13_458 = $signed(_T_96707); // @[Modules.scala 166:64:@44566.4]
  assign _T_96709 = $signed(buffer_9_311) + $signed(buffer_0_299); // @[Modules.scala 166:64:@44568.4]
  assign _T_96710 = _T_96709[13:0]; // @[Modules.scala 166:64:@44569.4]
  assign buffer_13_459 = $signed(_T_96710); // @[Modules.scala 166:64:@44570.4]
  assign _T_96712 = $signed(buffer_13_307) + $signed(buffer_13_308); // @[Modules.scala 166:64:@44572.4]
  assign _T_96713 = _T_96712[13:0]; // @[Modules.scala 166:64:@44573.4]
  assign buffer_13_460 = $signed(_T_96713); // @[Modules.scala 166:64:@44574.4]
  assign _T_96715 = $signed(buffer_13_309) + $signed(buffer_13_310); // @[Modules.scala 166:64:@44576.4]
  assign _T_96716 = _T_96715[13:0]; // @[Modules.scala 166:64:@44577.4]
  assign buffer_13_461 = $signed(_T_96716); // @[Modules.scala 166:64:@44578.4]
  assign _T_96718 = $signed(buffer_13_311) + $signed(buffer_13_312); // @[Modules.scala 166:64:@44580.4]
  assign _T_96719 = _T_96718[13:0]; // @[Modules.scala 166:64:@44581.4]
  assign buffer_13_462 = $signed(_T_96719); // @[Modules.scala 166:64:@44582.4]
  assign _T_96721 = $signed(buffer_13_313) + $signed(buffer_9_322); // @[Modules.scala 166:64:@44584.4]
  assign _T_96722 = _T_96721[13:0]; // @[Modules.scala 166:64:@44585.4]
  assign buffer_13_463 = $signed(_T_96722); // @[Modules.scala 166:64:@44586.4]
  assign _T_96724 = $signed(buffer_9_323) + $signed(buffer_9_324); // @[Modules.scala 166:64:@44588.4]
  assign _T_96725 = _T_96724[13:0]; // @[Modules.scala 166:64:@44589.4]
  assign buffer_13_464 = $signed(_T_96725); // @[Modules.scala 166:64:@44590.4]
  assign _T_96727 = $signed(buffer_13_317) + $signed(buffer_13_318); // @[Modules.scala 166:64:@44592.4]
  assign _T_96728 = _T_96727[13:0]; // @[Modules.scala 166:64:@44593.4]
  assign buffer_13_465 = $signed(_T_96728); // @[Modules.scala 166:64:@44594.4]
  assign _T_96736 = $signed(buffer_2_325) + $signed(buffer_13_324); // @[Modules.scala 166:64:@44604.4]
  assign _T_96737 = _T_96736[13:0]; // @[Modules.scala 166:64:@44605.4]
  assign buffer_13_468 = $signed(_T_96737); // @[Modules.scala 166:64:@44606.4]
  assign _T_96739 = $signed(buffer_13_325) + $signed(buffer_13_326); // @[Modules.scala 166:64:@44608.4]
  assign _T_96740 = _T_96739[13:0]; // @[Modules.scala 166:64:@44609.4]
  assign buffer_13_469 = $signed(_T_96740); // @[Modules.scala 166:64:@44610.4]
  assign _T_96742 = $signed(buffer_13_327) + $signed(buffer_13_328); // @[Modules.scala 166:64:@44612.4]
  assign _T_96743 = _T_96742[13:0]; // @[Modules.scala 166:64:@44613.4]
  assign buffer_13_470 = $signed(_T_96743); // @[Modules.scala 166:64:@44614.4]
  assign _T_96745 = $signed(buffer_13_329) + $signed(buffer_1_327); // @[Modules.scala 166:64:@44616.4]
  assign _T_96746 = _T_96745[13:0]; // @[Modules.scala 166:64:@44617.4]
  assign buffer_13_471 = $signed(_T_96746); // @[Modules.scala 166:64:@44618.4]
  assign _T_96748 = $signed(buffer_13_331) + $signed(buffer_5_339); // @[Modules.scala 166:64:@44620.4]
  assign _T_96749 = _T_96748[13:0]; // @[Modules.scala 166:64:@44621.4]
  assign buffer_13_472 = $signed(_T_96749); // @[Modules.scala 166:64:@44622.4]
  assign _T_96751 = $signed(buffer_13_333) + $signed(buffer_13_334); // @[Modules.scala 166:64:@44624.4]
  assign _T_96752 = _T_96751[13:0]; // @[Modules.scala 166:64:@44625.4]
  assign buffer_13_473 = $signed(_T_96752); // @[Modules.scala 166:64:@44626.4]
  assign _T_96754 = $signed(buffer_13_335) + $signed(buffer_13_336); // @[Modules.scala 166:64:@44628.4]
  assign _T_96755 = _T_96754[13:0]; // @[Modules.scala 166:64:@44629.4]
  assign buffer_13_474 = $signed(_T_96755); // @[Modules.scala 166:64:@44630.4]
  assign _T_96757 = $signed(buffer_13_337) + $signed(buffer_3_346); // @[Modules.scala 166:64:@44632.4]
  assign _T_96758 = _T_96757[13:0]; // @[Modules.scala 166:64:@44633.4]
  assign buffer_13_475 = $signed(_T_96758); // @[Modules.scala 166:64:@44634.4]
  assign _T_96760 = $signed(buffer_13_339) + $signed(buffer_13_340); // @[Modules.scala 166:64:@44636.4]
  assign _T_96761 = _T_96760[13:0]; // @[Modules.scala 166:64:@44637.4]
  assign buffer_13_476 = $signed(_T_96761); // @[Modules.scala 166:64:@44638.4]
  assign _T_96763 = $signed(buffer_13_341) + $signed(buffer_13_342); // @[Modules.scala 166:64:@44640.4]
  assign _T_96764 = _T_96763[13:0]; // @[Modules.scala 166:64:@44641.4]
  assign buffer_13_477 = $signed(_T_96764); // @[Modules.scala 166:64:@44642.4]
  assign _T_96766 = $signed(buffer_13_343) + $signed(buffer_13_344); // @[Modules.scala 166:64:@44644.4]
  assign _T_96767 = _T_96766[13:0]; // @[Modules.scala 166:64:@44645.4]
  assign buffer_13_478 = $signed(_T_96767); // @[Modules.scala 166:64:@44646.4]
  assign _T_96769 = $signed(buffer_13_345) + $signed(buffer_13_346); // @[Modules.scala 166:64:@44648.4]
  assign _T_96770 = _T_96769[13:0]; // @[Modules.scala 166:64:@44649.4]
  assign buffer_13_479 = $signed(_T_96770); // @[Modules.scala 166:64:@44650.4]
  assign _T_96772 = $signed(buffer_13_347) + $signed(buffer_6_356); // @[Modules.scala 166:64:@44652.4]
  assign _T_96773 = _T_96772[13:0]; // @[Modules.scala 166:64:@44653.4]
  assign buffer_13_480 = $signed(_T_96773); // @[Modules.scala 166:64:@44654.4]
  assign _T_96775 = $signed(buffer_13_349) + $signed(buffer_13_350); // @[Modules.scala 166:64:@44656.4]
  assign _T_96776 = _T_96775[13:0]; // @[Modules.scala 166:64:@44657.4]
  assign buffer_13_481 = $signed(_T_96776); // @[Modules.scala 166:64:@44658.4]
  assign _T_96778 = $signed(buffer_13_351) + $signed(buffer_13_352); // @[Modules.scala 166:64:@44660.4]
  assign _T_96779 = _T_96778[13:0]; // @[Modules.scala 166:64:@44661.4]
  assign buffer_13_482 = $signed(_T_96779); // @[Modules.scala 166:64:@44662.4]
  assign _T_96781 = $signed(buffer_13_353) + $signed(buffer_13_354); // @[Modules.scala 166:64:@44664.4]
  assign _T_96782 = _T_96781[13:0]; // @[Modules.scala 166:64:@44665.4]
  assign buffer_13_483 = $signed(_T_96782); // @[Modules.scala 166:64:@44666.4]
  assign _T_96784 = $signed(buffer_13_355) + $signed(buffer_2_359); // @[Modules.scala 166:64:@44668.4]
  assign _T_96785 = _T_96784[13:0]; // @[Modules.scala 166:64:@44669.4]
  assign buffer_13_484 = $signed(_T_96785); // @[Modules.scala 166:64:@44670.4]
  assign _T_96787 = $signed(buffer_2_360) + $signed(buffer_13_358); // @[Modules.scala 166:64:@44672.4]
  assign _T_96788 = _T_96787[13:0]; // @[Modules.scala 166:64:@44673.4]
  assign buffer_13_485 = $signed(_T_96788); // @[Modules.scala 166:64:@44674.4]
  assign _T_96790 = $signed(buffer_13_359) + $signed(buffer_13_360); // @[Modules.scala 166:64:@44676.4]
  assign _T_96791 = _T_96790[13:0]; // @[Modules.scala 166:64:@44677.4]
  assign buffer_13_486 = $signed(_T_96791); // @[Modules.scala 166:64:@44678.4]
  assign _T_96793 = $signed(buffer_13_361) + $signed(buffer_3_370); // @[Modules.scala 166:64:@44680.4]
  assign _T_96794 = _T_96793[13:0]; // @[Modules.scala 166:64:@44681.4]
  assign buffer_13_487 = $signed(_T_96794); // @[Modules.scala 166:64:@44682.4]
  assign _T_96796 = $signed(buffer_13_363) + $signed(buffer_13_364); // @[Modules.scala 166:64:@44684.4]
  assign _T_96797 = _T_96796[13:0]; // @[Modules.scala 166:64:@44685.4]
  assign buffer_13_488 = $signed(_T_96797); // @[Modules.scala 166:64:@44686.4]
  assign _T_96799 = $signed(buffer_13_365) + $signed(buffer_1_363); // @[Modules.scala 166:64:@44688.4]
  assign _T_96800 = _T_96799[13:0]; // @[Modules.scala 166:64:@44689.4]
  assign buffer_13_489 = $signed(_T_96800); // @[Modules.scala 166:64:@44690.4]
  assign _T_96802 = $signed(buffer_13_367) + $signed(buffer_13_368); // @[Modules.scala 166:64:@44692.4]
  assign _T_96803 = _T_96802[13:0]; // @[Modules.scala 166:64:@44693.4]
  assign buffer_13_490 = $signed(_T_96803); // @[Modules.scala 166:64:@44694.4]
  assign _T_96805 = $signed(buffer_13_369) + $signed(buffer_13_370); // @[Modules.scala 166:64:@44696.4]
  assign _T_96806 = _T_96805[13:0]; // @[Modules.scala 166:64:@44697.4]
  assign buffer_13_491 = $signed(_T_96806); // @[Modules.scala 166:64:@44698.4]
  assign _T_96808 = $signed(buffer_13_371) + $signed(buffer_13_372); // @[Modules.scala 166:64:@44700.4]
  assign _T_96809 = _T_96808[13:0]; // @[Modules.scala 166:64:@44701.4]
  assign buffer_13_492 = $signed(_T_96809); // @[Modules.scala 166:64:@44702.4]
  assign _T_96811 = $signed(buffer_13_373) + $signed(buffer_13_374); // @[Modules.scala 166:64:@44704.4]
  assign _T_96812 = _T_96811[13:0]; // @[Modules.scala 166:64:@44705.4]
  assign buffer_13_493 = $signed(_T_96812); // @[Modules.scala 166:64:@44706.4]
  assign _T_96814 = $signed(buffer_13_375) + $signed(buffer_13_376); // @[Modules.scala 166:64:@44708.4]
  assign _T_96815 = _T_96814[13:0]; // @[Modules.scala 166:64:@44709.4]
  assign buffer_13_494 = $signed(_T_96815); // @[Modules.scala 166:64:@44710.4]
  assign _T_96817 = $signed(buffer_7_379) + $signed(buffer_13_378); // @[Modules.scala 166:64:@44712.4]
  assign _T_96818 = _T_96817[13:0]; // @[Modules.scala 166:64:@44713.4]
  assign buffer_13_495 = $signed(_T_96818); // @[Modules.scala 166:64:@44714.4]
  assign _T_96820 = $signed(buffer_13_379) + $signed(buffer_13_380); // @[Modules.scala 166:64:@44716.4]
  assign _T_96821 = _T_96820[13:0]; // @[Modules.scala 166:64:@44717.4]
  assign buffer_13_496 = $signed(_T_96821); // @[Modules.scala 166:64:@44718.4]
  assign _T_96823 = $signed(buffer_13_381) + $signed(buffer_13_382); // @[Modules.scala 166:64:@44720.4]
  assign _T_96824 = _T_96823[13:0]; // @[Modules.scala 166:64:@44721.4]
  assign buffer_13_497 = $signed(_T_96824); // @[Modules.scala 166:64:@44722.4]
  assign _T_96826 = $signed(buffer_13_383) + $signed(buffer_13_384); // @[Modules.scala 166:64:@44724.4]
  assign _T_96827 = _T_96826[13:0]; // @[Modules.scala 166:64:@44725.4]
  assign buffer_13_498 = $signed(_T_96827); // @[Modules.scala 166:64:@44726.4]
  assign _T_96829 = $signed(buffer_13_385) + $signed(buffer_13_386); // @[Modules.scala 166:64:@44728.4]
  assign _T_96830 = _T_96829[13:0]; // @[Modules.scala 166:64:@44729.4]
  assign buffer_13_499 = $signed(_T_96830); // @[Modules.scala 166:64:@44730.4]
  assign _T_96832 = $signed(buffer_13_387) + $signed(buffer_13_388); // @[Modules.scala 166:64:@44732.4]
  assign _T_96833 = _T_96832[13:0]; // @[Modules.scala 166:64:@44733.4]
  assign buffer_13_500 = $signed(_T_96833); // @[Modules.scala 166:64:@44734.4]
  assign _T_96835 = $signed(buffer_1_386) + $signed(buffer_13_390); // @[Modules.scala 166:64:@44736.4]
  assign _T_96836 = _T_96835[13:0]; // @[Modules.scala 166:64:@44737.4]
  assign buffer_13_501 = $signed(_T_96836); // @[Modules.scala 166:64:@44738.4]
  assign _T_96838 = $signed(buffer_11_380) + $signed(buffer_13_392); // @[Modules.scala 166:64:@44740.4]
  assign _T_96839 = _T_96838[13:0]; // @[Modules.scala 166:64:@44741.4]
  assign buffer_13_502 = $signed(_T_96839); // @[Modules.scala 166:64:@44742.4]
  assign _T_96841 = $signed(buffer_13_393) + $signed(buffer_13_394); // @[Modules.scala 166:64:@44744.4]
  assign _T_96842 = _T_96841[13:0]; // @[Modules.scala 166:64:@44745.4]
  assign buffer_13_503 = $signed(_T_96842); // @[Modules.scala 166:64:@44746.4]
  assign _T_96844 = $signed(buffer_13_395) + $signed(buffer_13_396); // @[Modules.scala 166:64:@44748.4]
  assign _T_96845 = _T_96844[13:0]; // @[Modules.scala 166:64:@44749.4]
  assign buffer_13_504 = $signed(_T_96845); // @[Modules.scala 166:64:@44750.4]
  assign _T_96847 = $signed(buffer_13_397) + $signed(buffer_13_398); // @[Modules.scala 166:64:@44752.4]
  assign _T_96848 = _T_96847[13:0]; // @[Modules.scala 166:64:@44753.4]
  assign buffer_13_505 = $signed(_T_96848); // @[Modules.scala 166:64:@44754.4]
  assign _T_96850 = $signed(buffer_7_404) + $signed(buffer_13_400); // @[Modules.scala 166:64:@44756.4]
  assign _T_96851 = _T_96850[13:0]; // @[Modules.scala 166:64:@44757.4]
  assign buffer_13_506 = $signed(_T_96851); // @[Modules.scala 166:64:@44758.4]
  assign _T_96853 = $signed(buffer_10_405) + $signed(buffer_0_396); // @[Modules.scala 166:64:@44760.4]
  assign _T_96854 = _T_96853[13:0]; // @[Modules.scala 166:64:@44761.4]
  assign buffer_13_507 = $signed(_T_96854); // @[Modules.scala 166:64:@44762.4]
  assign _T_96856 = $signed(buffer_13_403) + $signed(buffer_13_404); // @[Modules.scala 166:64:@44764.4]
  assign _T_96857 = _T_96856[13:0]; // @[Modules.scala 166:64:@44765.4]
  assign buffer_13_508 = $signed(_T_96857); // @[Modules.scala 166:64:@44766.4]
  assign _T_96859 = $signed(buffer_6_418) + $signed(buffer_13_406); // @[Modules.scala 166:64:@44768.4]
  assign _T_96860 = _T_96859[13:0]; // @[Modules.scala 166:64:@44769.4]
  assign buffer_13_509 = $signed(_T_96860); // @[Modules.scala 166:64:@44770.4]
  assign _T_96862 = $signed(buffer_13_407) + $signed(buffer_10_411); // @[Modules.scala 166:64:@44772.4]
  assign _T_96863 = _T_96862[13:0]; // @[Modules.scala 166:64:@44773.4]
  assign buffer_13_510 = $signed(_T_96863); // @[Modules.scala 166:64:@44774.4]
  assign _T_96865 = $signed(buffer_13_409) + $signed(buffer_13_410); // @[Modules.scala 166:64:@44776.4]
  assign _T_96866 = _T_96865[13:0]; // @[Modules.scala 166:64:@44777.4]
  assign buffer_13_511 = $signed(_T_96866); // @[Modules.scala 166:64:@44778.4]
  assign _T_96868 = $signed(buffer_13_411) + $signed(buffer_13_412); // @[Modules.scala 166:64:@44780.4]
  assign _T_96869 = _T_96868[13:0]; // @[Modules.scala 166:64:@44781.4]
  assign buffer_13_512 = $signed(_T_96869); // @[Modules.scala 166:64:@44782.4]
  assign _T_96871 = $signed(buffer_13_413) + $signed(buffer_6_428); // @[Modules.scala 166:64:@44784.4]
  assign _T_96872 = _T_96871[13:0]; // @[Modules.scala 166:64:@44785.4]
  assign buffer_13_513 = $signed(_T_96872); // @[Modules.scala 166:64:@44786.4]
  assign _T_96874 = $signed(buffer_13_415) + $signed(buffer_13_416); // @[Modules.scala 166:64:@44788.4]
  assign _T_96875 = _T_96874[13:0]; // @[Modules.scala 166:64:@44789.4]
  assign buffer_13_514 = $signed(_T_96875); // @[Modules.scala 166:64:@44790.4]
  assign _T_96877 = $signed(buffer_8_421) + $signed(buffer_11_409); // @[Modules.scala 166:64:@44792.4]
  assign _T_96878 = _T_96877[13:0]; // @[Modules.scala 166:64:@44793.4]
  assign buffer_13_515 = $signed(_T_96878); // @[Modules.scala 166:64:@44794.4]
  assign _T_96880 = $signed(buffer_13_419) + $signed(buffer_13_420); // @[Modules.scala 166:64:@44796.4]
  assign _T_96881 = _T_96880[13:0]; // @[Modules.scala 166:64:@44797.4]
  assign buffer_13_516 = $signed(_T_96881); // @[Modules.scala 166:64:@44798.4]
  assign _T_96883 = $signed(buffer_13_421) + $signed(buffer_13_422); // @[Modules.scala 166:64:@44800.4]
  assign _T_96884 = _T_96883[13:0]; // @[Modules.scala 166:64:@44801.4]
  assign buffer_13_517 = $signed(_T_96884); // @[Modules.scala 166:64:@44802.4]
  assign _T_96886 = $signed(buffer_13_423) + $signed(buffer_13_424); // @[Modules.scala 166:64:@44804.4]
  assign _T_96887 = _T_96886[13:0]; // @[Modules.scala 166:64:@44805.4]
  assign buffer_13_518 = $signed(_T_96887); // @[Modules.scala 166:64:@44806.4]
  assign _T_96889 = $signed(buffer_13_425) + $signed(buffer_13_426); // @[Modules.scala 166:64:@44808.4]
  assign _T_96890 = _T_96889[13:0]; // @[Modules.scala 166:64:@44809.4]
  assign buffer_13_519 = $signed(_T_96890); // @[Modules.scala 166:64:@44810.4]
  assign _T_96892 = $signed(buffer_13_427) + $signed(buffer_8_433); // @[Modules.scala 166:64:@44812.4]
  assign _T_96893 = _T_96892[13:0]; // @[Modules.scala 166:64:@44813.4]
  assign buffer_13_520 = $signed(_T_96893); // @[Modules.scala 166:64:@44814.4]
  assign _T_96895 = $signed(buffer_13_429) + $signed(buffer_13_430); // @[Modules.scala 166:64:@44816.4]
  assign _T_96896 = _T_96895[13:0]; // @[Modules.scala 166:64:@44817.4]
  assign buffer_13_521 = $signed(_T_96896); // @[Modules.scala 166:64:@44818.4]
  assign _T_96898 = $signed(buffer_13_431) + $signed(buffer_11_422); // @[Modules.scala 166:64:@44820.4]
  assign _T_96899 = _T_96898[13:0]; // @[Modules.scala 166:64:@44821.4]
  assign buffer_13_522 = $signed(_T_96899); // @[Modules.scala 166:64:@44822.4]
  assign _T_96901 = $signed(buffer_13_433) + $signed(buffer_13_434); // @[Modules.scala 166:64:@44824.4]
  assign _T_96902 = _T_96901[13:0]; // @[Modules.scala 166:64:@44825.4]
  assign buffer_13_523 = $signed(_T_96902); // @[Modules.scala 166:64:@44826.4]
  assign _T_96904 = $signed(buffer_13_435) + $signed(buffer_13_436); // @[Modules.scala 166:64:@44828.4]
  assign _T_96905 = _T_96904[13:0]; // @[Modules.scala 166:64:@44829.4]
  assign buffer_13_524 = $signed(_T_96905); // @[Modules.scala 166:64:@44830.4]
  assign _T_96907 = $signed(buffer_13_437) + $signed(buffer_10_440); // @[Modules.scala 166:64:@44832.4]
  assign _T_96908 = _T_96907[13:0]; // @[Modules.scala 166:64:@44833.4]
  assign buffer_13_525 = $signed(_T_96908); // @[Modules.scala 166:64:@44834.4]
  assign _T_96910 = $signed(buffer_3_449) + $signed(buffer_13_440); // @[Modules.scala 166:64:@44836.4]
  assign _T_96911 = _T_96910[13:0]; // @[Modules.scala 166:64:@44837.4]
  assign buffer_13_526 = $signed(_T_96911); // @[Modules.scala 166:64:@44838.4]
  assign _T_96913 = $signed(buffer_13_441) + $signed(buffer_13_442); // @[Modules.scala 166:64:@44840.4]
  assign _T_96914 = _T_96913[13:0]; // @[Modules.scala 166:64:@44841.4]
  assign buffer_13_527 = $signed(_T_96914); // @[Modules.scala 166:64:@44842.4]
  assign _T_96916 = $signed(buffer_13_443) + $signed(buffer_13_444); // @[Modules.scala 166:64:@44844.4]
  assign _T_96917 = _T_96916[13:0]; // @[Modules.scala 166:64:@44845.4]
  assign buffer_13_528 = $signed(_T_96917); // @[Modules.scala 166:64:@44846.4]
  assign _T_96919 = $signed(buffer_13_445) + $signed(buffer_13_446); // @[Modules.scala 166:64:@44848.4]
  assign _T_96920 = _T_96919[13:0]; // @[Modules.scala 166:64:@44849.4]
  assign buffer_13_529 = $signed(_T_96920); // @[Modules.scala 166:64:@44850.4]
  assign _T_96922 = $signed(buffer_13_447) + $signed(buffer_0_441); // @[Modules.scala 166:64:@44852.4]
  assign _T_96923 = _T_96922[13:0]; // @[Modules.scala 166:64:@44853.4]
  assign buffer_13_530 = $signed(_T_96923); // @[Modules.scala 166:64:@44854.4]
  assign _T_96928 = $signed(buffer_13_451) + $signed(buffer_13_452); // @[Modules.scala 166:64:@44860.4]
  assign _T_96929 = _T_96928[13:0]; // @[Modules.scala 166:64:@44861.4]
  assign buffer_13_532 = $signed(_T_96929); // @[Modules.scala 166:64:@44862.4]
  assign _T_96931 = $signed(buffer_13_453) + $signed(buffer_13_454); // @[Modules.scala 166:64:@44864.4]
  assign _T_96932 = _T_96931[13:0]; // @[Modules.scala 166:64:@44865.4]
  assign buffer_13_533 = $signed(_T_96932); // @[Modules.scala 166:64:@44866.4]
  assign _T_96934 = $signed(buffer_13_455) + $signed(buffer_13_456); // @[Modules.scala 166:64:@44868.4]
  assign _T_96935 = _T_96934[13:0]; // @[Modules.scala 166:64:@44869.4]
  assign buffer_13_534 = $signed(_T_96935); // @[Modules.scala 166:64:@44870.4]
  assign _T_96937 = $signed(buffer_13_457) + $signed(buffer_13_458); // @[Modules.scala 166:64:@44872.4]
  assign _T_96938 = _T_96937[13:0]; // @[Modules.scala 166:64:@44873.4]
  assign buffer_13_535 = $signed(_T_96938); // @[Modules.scala 166:64:@44874.4]
  assign _T_96940 = $signed(buffer_13_459) + $signed(buffer_0_300); // @[Modules.scala 172:66:@44876.4]
  assign _T_96941 = _T_96940[13:0]; // @[Modules.scala 172:66:@44877.4]
  assign buffer_13_536 = $signed(_T_96941); // @[Modules.scala 172:66:@44878.4]
  assign _T_96943 = $signed(buffer_13_460) + $signed(buffer_13_461); // @[Modules.scala 166:64:@44880.4]
  assign _T_96944 = _T_96943[13:0]; // @[Modules.scala 166:64:@44881.4]
  assign buffer_13_537 = $signed(_T_96944); // @[Modules.scala 166:64:@44882.4]
  assign _T_96946 = $signed(buffer_13_462) + $signed(buffer_13_463); // @[Modules.scala 166:64:@44884.4]
  assign _T_96947 = _T_96946[13:0]; // @[Modules.scala 166:64:@44885.4]
  assign buffer_13_538 = $signed(_T_96947); // @[Modules.scala 166:64:@44886.4]
  assign _T_96949 = $signed(buffer_13_464) + $signed(buffer_13_465); // @[Modules.scala 166:64:@44888.4]
  assign _T_96950 = _T_96949[13:0]; // @[Modules.scala 166:64:@44889.4]
  assign buffer_13_539 = $signed(_T_96950); // @[Modules.scala 166:64:@44890.4]
  assign _T_96955 = $signed(buffer_13_468) + $signed(buffer_13_469); // @[Modules.scala 166:64:@44896.4]
  assign _T_96956 = _T_96955[13:0]; // @[Modules.scala 166:64:@44897.4]
  assign buffer_13_541 = $signed(_T_96956); // @[Modules.scala 166:64:@44898.4]
  assign _T_96958 = $signed(buffer_13_470) + $signed(buffer_13_471); // @[Modules.scala 166:64:@44900.4]
  assign _T_96959 = _T_96958[13:0]; // @[Modules.scala 166:64:@44901.4]
  assign buffer_13_542 = $signed(_T_96959); // @[Modules.scala 166:64:@44902.4]
  assign _T_96961 = $signed(buffer_13_472) + $signed(buffer_13_473); // @[Modules.scala 166:64:@44904.4]
  assign _T_96962 = _T_96961[13:0]; // @[Modules.scala 166:64:@44905.4]
  assign buffer_13_543 = $signed(_T_96962); // @[Modules.scala 166:64:@44906.4]
  assign _T_96964 = $signed(buffer_13_474) + $signed(buffer_13_475); // @[Modules.scala 166:64:@44908.4]
  assign _T_96965 = _T_96964[13:0]; // @[Modules.scala 166:64:@44909.4]
  assign buffer_13_544 = $signed(_T_96965); // @[Modules.scala 166:64:@44910.4]
  assign _T_96967 = $signed(buffer_13_476) + $signed(buffer_13_477); // @[Modules.scala 166:64:@44912.4]
  assign _T_96968 = _T_96967[13:0]; // @[Modules.scala 166:64:@44913.4]
  assign buffer_13_545 = $signed(_T_96968); // @[Modules.scala 166:64:@44914.4]
  assign _T_96970 = $signed(buffer_13_478) + $signed(buffer_13_479); // @[Modules.scala 166:64:@44916.4]
  assign _T_96971 = _T_96970[13:0]; // @[Modules.scala 166:64:@44917.4]
  assign buffer_13_546 = $signed(_T_96971); // @[Modules.scala 166:64:@44918.4]
  assign _T_96973 = $signed(buffer_13_480) + $signed(buffer_13_481); // @[Modules.scala 166:64:@44920.4]
  assign _T_96974 = _T_96973[13:0]; // @[Modules.scala 166:64:@44921.4]
  assign buffer_13_547 = $signed(_T_96974); // @[Modules.scala 166:64:@44922.4]
  assign _T_96976 = $signed(buffer_13_482) + $signed(buffer_13_483); // @[Modules.scala 166:64:@44924.4]
  assign _T_96977 = _T_96976[13:0]; // @[Modules.scala 166:64:@44925.4]
  assign buffer_13_548 = $signed(_T_96977); // @[Modules.scala 166:64:@44926.4]
  assign _T_96979 = $signed(buffer_13_484) + $signed(buffer_13_485); // @[Modules.scala 166:64:@44928.4]
  assign _T_96980 = _T_96979[13:0]; // @[Modules.scala 166:64:@44929.4]
  assign buffer_13_549 = $signed(_T_96980); // @[Modules.scala 166:64:@44930.4]
  assign _T_96982 = $signed(buffer_13_486) + $signed(buffer_13_487); // @[Modules.scala 166:64:@44932.4]
  assign _T_96983 = _T_96982[13:0]; // @[Modules.scala 166:64:@44933.4]
  assign buffer_13_550 = $signed(_T_96983); // @[Modules.scala 166:64:@44934.4]
  assign _T_96985 = $signed(buffer_13_488) + $signed(buffer_13_489); // @[Modules.scala 166:64:@44936.4]
  assign _T_96986 = _T_96985[13:0]; // @[Modules.scala 166:64:@44937.4]
  assign buffer_13_551 = $signed(_T_96986); // @[Modules.scala 166:64:@44938.4]
  assign _T_96988 = $signed(buffer_13_490) + $signed(buffer_13_491); // @[Modules.scala 166:64:@44940.4]
  assign _T_96989 = _T_96988[13:0]; // @[Modules.scala 166:64:@44941.4]
  assign buffer_13_552 = $signed(_T_96989); // @[Modules.scala 166:64:@44942.4]
  assign _T_96991 = $signed(buffer_13_492) + $signed(buffer_13_493); // @[Modules.scala 166:64:@44944.4]
  assign _T_96992 = _T_96991[13:0]; // @[Modules.scala 166:64:@44945.4]
  assign buffer_13_553 = $signed(_T_96992); // @[Modules.scala 166:64:@44946.4]
  assign _T_96994 = $signed(buffer_13_494) + $signed(buffer_13_495); // @[Modules.scala 166:64:@44948.4]
  assign _T_96995 = _T_96994[13:0]; // @[Modules.scala 166:64:@44949.4]
  assign buffer_13_554 = $signed(_T_96995); // @[Modules.scala 166:64:@44950.4]
  assign _T_96997 = $signed(buffer_13_496) + $signed(buffer_13_497); // @[Modules.scala 166:64:@44952.4]
  assign _T_96998 = _T_96997[13:0]; // @[Modules.scala 166:64:@44953.4]
  assign buffer_13_555 = $signed(_T_96998); // @[Modules.scala 166:64:@44954.4]
  assign _T_97000 = $signed(buffer_13_498) + $signed(buffer_13_499); // @[Modules.scala 166:64:@44956.4]
  assign _T_97001 = _T_97000[13:0]; // @[Modules.scala 166:64:@44957.4]
  assign buffer_13_556 = $signed(_T_97001); // @[Modules.scala 166:64:@44958.4]
  assign _T_97003 = $signed(buffer_13_500) + $signed(buffer_13_501); // @[Modules.scala 166:64:@44960.4]
  assign _T_97004 = _T_97003[13:0]; // @[Modules.scala 166:64:@44961.4]
  assign buffer_13_557 = $signed(_T_97004); // @[Modules.scala 166:64:@44962.4]
  assign _T_97006 = $signed(buffer_13_502) + $signed(buffer_13_503); // @[Modules.scala 166:64:@44964.4]
  assign _T_97007 = _T_97006[13:0]; // @[Modules.scala 166:64:@44965.4]
  assign buffer_13_558 = $signed(_T_97007); // @[Modules.scala 166:64:@44966.4]
  assign _T_97009 = $signed(buffer_13_504) + $signed(buffer_13_505); // @[Modules.scala 166:64:@44968.4]
  assign _T_97010 = _T_97009[13:0]; // @[Modules.scala 166:64:@44969.4]
  assign buffer_13_559 = $signed(_T_97010); // @[Modules.scala 166:64:@44970.4]
  assign _T_97012 = $signed(buffer_13_506) + $signed(buffer_13_507); // @[Modules.scala 166:64:@44972.4]
  assign _T_97013 = _T_97012[13:0]; // @[Modules.scala 166:64:@44973.4]
  assign buffer_13_560 = $signed(_T_97013); // @[Modules.scala 166:64:@44974.4]
  assign _T_97015 = $signed(buffer_13_508) + $signed(buffer_13_509); // @[Modules.scala 166:64:@44976.4]
  assign _T_97016 = _T_97015[13:0]; // @[Modules.scala 166:64:@44977.4]
  assign buffer_13_561 = $signed(_T_97016); // @[Modules.scala 166:64:@44978.4]
  assign _T_97018 = $signed(buffer_13_510) + $signed(buffer_13_511); // @[Modules.scala 166:64:@44980.4]
  assign _T_97019 = _T_97018[13:0]; // @[Modules.scala 166:64:@44981.4]
  assign buffer_13_562 = $signed(_T_97019); // @[Modules.scala 166:64:@44982.4]
  assign _T_97021 = $signed(buffer_13_512) + $signed(buffer_13_513); // @[Modules.scala 166:64:@44984.4]
  assign _T_97022 = _T_97021[13:0]; // @[Modules.scala 166:64:@44985.4]
  assign buffer_13_563 = $signed(_T_97022); // @[Modules.scala 166:64:@44986.4]
  assign _T_97024 = $signed(buffer_13_514) + $signed(buffer_13_515); // @[Modules.scala 166:64:@44988.4]
  assign _T_97025 = _T_97024[13:0]; // @[Modules.scala 166:64:@44989.4]
  assign buffer_13_564 = $signed(_T_97025); // @[Modules.scala 166:64:@44990.4]
  assign _T_97027 = $signed(buffer_13_516) + $signed(buffer_13_517); // @[Modules.scala 166:64:@44992.4]
  assign _T_97028 = _T_97027[13:0]; // @[Modules.scala 166:64:@44993.4]
  assign buffer_13_565 = $signed(_T_97028); // @[Modules.scala 166:64:@44994.4]
  assign _T_97030 = $signed(buffer_13_518) + $signed(buffer_13_519); // @[Modules.scala 166:64:@44996.4]
  assign _T_97031 = _T_97030[13:0]; // @[Modules.scala 166:64:@44997.4]
  assign buffer_13_566 = $signed(_T_97031); // @[Modules.scala 166:64:@44998.4]
  assign _T_97033 = $signed(buffer_13_520) + $signed(buffer_13_521); // @[Modules.scala 166:64:@45000.4]
  assign _T_97034 = _T_97033[13:0]; // @[Modules.scala 166:64:@45001.4]
  assign buffer_13_567 = $signed(_T_97034); // @[Modules.scala 166:64:@45002.4]
  assign _T_97036 = $signed(buffer_13_522) + $signed(buffer_13_523); // @[Modules.scala 166:64:@45004.4]
  assign _T_97037 = _T_97036[13:0]; // @[Modules.scala 166:64:@45005.4]
  assign buffer_13_568 = $signed(_T_97037); // @[Modules.scala 166:64:@45006.4]
  assign _T_97039 = $signed(buffer_13_524) + $signed(buffer_13_525); // @[Modules.scala 166:64:@45008.4]
  assign _T_97040 = _T_97039[13:0]; // @[Modules.scala 166:64:@45009.4]
  assign buffer_13_569 = $signed(_T_97040); // @[Modules.scala 166:64:@45010.4]
  assign _T_97042 = $signed(buffer_13_526) + $signed(buffer_13_527); // @[Modules.scala 166:64:@45012.4]
  assign _T_97043 = _T_97042[13:0]; // @[Modules.scala 166:64:@45013.4]
  assign buffer_13_570 = $signed(_T_97043); // @[Modules.scala 166:64:@45014.4]
  assign _T_97045 = $signed(buffer_13_528) + $signed(buffer_13_529); // @[Modules.scala 166:64:@45016.4]
  assign _T_97046 = _T_97045[13:0]; // @[Modules.scala 166:64:@45017.4]
  assign buffer_13_571 = $signed(_T_97046); // @[Modules.scala 166:64:@45018.4]
  assign _T_97048 = $signed(buffer_13_530) + $signed(buffer_0_523); // @[Modules.scala 166:64:@45020.4]
  assign _T_97049 = _T_97048[13:0]; // @[Modules.scala 166:64:@45021.4]
  assign buffer_13_572 = $signed(_T_97049); // @[Modules.scala 166:64:@45022.4]
  assign _T_97051 = $signed(buffer_13_532) + $signed(buffer_13_533); // @[Modules.scala 166:64:@45024.4]
  assign _T_97052 = _T_97051[13:0]; // @[Modules.scala 166:64:@45025.4]
  assign buffer_13_573 = $signed(_T_97052); // @[Modules.scala 166:64:@45026.4]
  assign _T_97054 = $signed(buffer_13_534) + $signed(buffer_13_535); // @[Modules.scala 166:64:@45028.4]
  assign _T_97055 = _T_97054[13:0]; // @[Modules.scala 166:64:@45029.4]
  assign buffer_13_574 = $signed(_T_97055); // @[Modules.scala 166:64:@45030.4]
  assign _T_97057 = $signed(buffer_13_537) + $signed(buffer_13_538); // @[Modules.scala 160:64:@45032.4]
  assign _T_97058 = _T_97057[13:0]; // @[Modules.scala 160:64:@45033.4]
  assign buffer_13_575 = $signed(_T_97058); // @[Modules.scala 160:64:@45034.4]
  assign _T_97060 = $signed(buffer_13_539) + $signed(buffer_10_542); // @[Modules.scala 160:64:@45036.4]
  assign _T_97061 = _T_97060[13:0]; // @[Modules.scala 160:64:@45037.4]
  assign buffer_13_576 = $signed(_T_97061); // @[Modules.scala 160:64:@45038.4]
  assign _T_97063 = $signed(buffer_13_541) + $signed(buffer_13_542); // @[Modules.scala 160:64:@45040.4]
  assign _T_97064 = _T_97063[13:0]; // @[Modules.scala 160:64:@45041.4]
  assign buffer_13_577 = $signed(_T_97064); // @[Modules.scala 160:64:@45042.4]
  assign _T_97066 = $signed(buffer_13_543) + $signed(buffer_13_544); // @[Modules.scala 160:64:@45044.4]
  assign _T_97067 = _T_97066[13:0]; // @[Modules.scala 160:64:@45045.4]
  assign buffer_13_578 = $signed(_T_97067); // @[Modules.scala 160:64:@45046.4]
  assign _T_97069 = $signed(buffer_13_545) + $signed(buffer_13_546); // @[Modules.scala 160:64:@45048.4]
  assign _T_97070 = _T_97069[13:0]; // @[Modules.scala 160:64:@45049.4]
  assign buffer_13_579 = $signed(_T_97070); // @[Modules.scala 160:64:@45050.4]
  assign _T_97072 = $signed(buffer_13_547) + $signed(buffer_13_548); // @[Modules.scala 160:64:@45052.4]
  assign _T_97073 = _T_97072[13:0]; // @[Modules.scala 160:64:@45053.4]
  assign buffer_13_580 = $signed(_T_97073); // @[Modules.scala 160:64:@45054.4]
  assign _T_97075 = $signed(buffer_13_549) + $signed(buffer_13_550); // @[Modules.scala 160:64:@45056.4]
  assign _T_97076 = _T_97075[13:0]; // @[Modules.scala 160:64:@45057.4]
  assign buffer_13_581 = $signed(_T_97076); // @[Modules.scala 160:64:@45058.4]
  assign _T_97078 = $signed(buffer_13_551) + $signed(buffer_13_552); // @[Modules.scala 160:64:@45060.4]
  assign _T_97079 = _T_97078[13:0]; // @[Modules.scala 160:64:@45061.4]
  assign buffer_13_582 = $signed(_T_97079); // @[Modules.scala 160:64:@45062.4]
  assign _T_97081 = $signed(buffer_13_553) + $signed(buffer_13_554); // @[Modules.scala 160:64:@45064.4]
  assign _T_97082 = _T_97081[13:0]; // @[Modules.scala 160:64:@45065.4]
  assign buffer_13_583 = $signed(_T_97082); // @[Modules.scala 160:64:@45066.4]
  assign _T_97084 = $signed(buffer_13_555) + $signed(buffer_13_556); // @[Modules.scala 160:64:@45068.4]
  assign _T_97085 = _T_97084[13:0]; // @[Modules.scala 160:64:@45069.4]
  assign buffer_13_584 = $signed(_T_97085); // @[Modules.scala 160:64:@45070.4]
  assign _T_97087 = $signed(buffer_13_557) + $signed(buffer_13_558); // @[Modules.scala 160:64:@45072.4]
  assign _T_97088 = _T_97087[13:0]; // @[Modules.scala 160:64:@45073.4]
  assign buffer_13_585 = $signed(_T_97088); // @[Modules.scala 160:64:@45074.4]
  assign _T_97090 = $signed(buffer_13_559) + $signed(buffer_13_560); // @[Modules.scala 160:64:@45076.4]
  assign _T_97091 = _T_97090[13:0]; // @[Modules.scala 160:64:@45077.4]
  assign buffer_13_586 = $signed(_T_97091); // @[Modules.scala 160:64:@45078.4]
  assign _T_97093 = $signed(buffer_13_561) + $signed(buffer_13_562); // @[Modules.scala 160:64:@45080.4]
  assign _T_97094 = _T_97093[13:0]; // @[Modules.scala 160:64:@45081.4]
  assign buffer_13_587 = $signed(_T_97094); // @[Modules.scala 160:64:@45082.4]
  assign _T_97096 = $signed(buffer_13_563) + $signed(buffer_13_564); // @[Modules.scala 160:64:@45084.4]
  assign _T_97097 = _T_97096[13:0]; // @[Modules.scala 160:64:@45085.4]
  assign buffer_13_588 = $signed(_T_97097); // @[Modules.scala 160:64:@45086.4]
  assign _T_97099 = $signed(buffer_13_565) + $signed(buffer_13_566); // @[Modules.scala 160:64:@45088.4]
  assign _T_97100 = _T_97099[13:0]; // @[Modules.scala 160:64:@45089.4]
  assign buffer_13_589 = $signed(_T_97100); // @[Modules.scala 160:64:@45090.4]
  assign _T_97102 = $signed(buffer_13_567) + $signed(buffer_13_568); // @[Modules.scala 160:64:@45092.4]
  assign _T_97103 = _T_97102[13:0]; // @[Modules.scala 160:64:@45093.4]
  assign buffer_13_590 = $signed(_T_97103); // @[Modules.scala 160:64:@45094.4]
  assign _T_97105 = $signed(buffer_13_569) + $signed(buffer_13_570); // @[Modules.scala 160:64:@45096.4]
  assign _T_97106 = _T_97105[13:0]; // @[Modules.scala 160:64:@45097.4]
  assign buffer_13_591 = $signed(_T_97106); // @[Modules.scala 160:64:@45098.4]
  assign _T_97108 = $signed(buffer_13_571) + $signed(buffer_13_572); // @[Modules.scala 160:64:@45100.4]
  assign _T_97109 = _T_97108[13:0]; // @[Modules.scala 160:64:@45101.4]
  assign buffer_13_592 = $signed(_T_97109); // @[Modules.scala 160:64:@45102.4]
  assign _T_97111 = $signed(buffer_13_573) + $signed(buffer_13_574); // @[Modules.scala 160:64:@45104.4]
  assign _T_97112 = _T_97111[13:0]; // @[Modules.scala 160:64:@45105.4]
  assign buffer_13_593 = $signed(_T_97112); // @[Modules.scala 160:64:@45106.4]
  assign _T_97114 = $signed(buffer_13_575) + $signed(buffer_13_576); // @[Modules.scala 166:64:@45108.4]
  assign _T_97115 = _T_97114[13:0]; // @[Modules.scala 166:64:@45109.4]
  assign buffer_13_594 = $signed(_T_97115); // @[Modules.scala 166:64:@45110.4]
  assign _T_97117 = $signed(buffer_13_577) + $signed(buffer_13_578); // @[Modules.scala 166:64:@45112.4]
  assign _T_97118 = _T_97117[13:0]; // @[Modules.scala 166:64:@45113.4]
  assign buffer_13_595 = $signed(_T_97118); // @[Modules.scala 166:64:@45114.4]
  assign _T_97120 = $signed(buffer_13_579) + $signed(buffer_13_580); // @[Modules.scala 166:64:@45116.4]
  assign _T_97121 = _T_97120[13:0]; // @[Modules.scala 166:64:@45117.4]
  assign buffer_13_596 = $signed(_T_97121); // @[Modules.scala 166:64:@45118.4]
  assign _T_97123 = $signed(buffer_13_581) + $signed(buffer_13_582); // @[Modules.scala 166:64:@45120.4]
  assign _T_97124 = _T_97123[13:0]; // @[Modules.scala 166:64:@45121.4]
  assign buffer_13_597 = $signed(_T_97124); // @[Modules.scala 166:64:@45122.4]
  assign _T_97126 = $signed(buffer_13_583) + $signed(buffer_13_584); // @[Modules.scala 166:64:@45124.4]
  assign _T_97127 = _T_97126[13:0]; // @[Modules.scala 166:64:@45125.4]
  assign buffer_13_598 = $signed(_T_97127); // @[Modules.scala 166:64:@45126.4]
  assign _T_97129 = $signed(buffer_13_585) + $signed(buffer_13_586); // @[Modules.scala 166:64:@45128.4]
  assign _T_97130 = _T_97129[13:0]; // @[Modules.scala 166:64:@45129.4]
  assign buffer_13_599 = $signed(_T_97130); // @[Modules.scala 166:64:@45130.4]
  assign _T_97132 = $signed(buffer_13_587) + $signed(buffer_13_588); // @[Modules.scala 166:64:@45132.4]
  assign _T_97133 = _T_97132[13:0]; // @[Modules.scala 166:64:@45133.4]
  assign buffer_13_600 = $signed(_T_97133); // @[Modules.scala 166:64:@45134.4]
  assign _T_97135 = $signed(buffer_13_589) + $signed(buffer_13_590); // @[Modules.scala 166:64:@45136.4]
  assign _T_97136 = _T_97135[13:0]; // @[Modules.scala 166:64:@45137.4]
  assign buffer_13_601 = $signed(_T_97136); // @[Modules.scala 166:64:@45138.4]
  assign _T_97138 = $signed(buffer_13_591) + $signed(buffer_13_592); // @[Modules.scala 166:64:@45140.4]
  assign _T_97139 = _T_97138[13:0]; // @[Modules.scala 166:64:@45141.4]
  assign buffer_13_602 = $signed(_T_97139); // @[Modules.scala 166:64:@45142.4]
  assign _T_97141 = $signed(buffer_13_593) + $signed(buffer_13_536); // @[Modules.scala 172:66:@45144.4]
  assign _T_97142 = _T_97141[13:0]; // @[Modules.scala 172:66:@45145.4]
  assign buffer_13_603 = $signed(_T_97142); // @[Modules.scala 172:66:@45146.4]
  assign _T_97144 = $signed(buffer_13_594) + $signed(buffer_13_595); // @[Modules.scala 160:64:@45148.4]
  assign _T_97145 = _T_97144[13:0]; // @[Modules.scala 160:64:@45149.4]
  assign buffer_13_604 = $signed(_T_97145); // @[Modules.scala 160:64:@45150.4]
  assign _T_97147 = $signed(buffer_13_596) + $signed(buffer_13_597); // @[Modules.scala 160:64:@45152.4]
  assign _T_97148 = _T_97147[13:0]; // @[Modules.scala 160:64:@45153.4]
  assign buffer_13_605 = $signed(_T_97148); // @[Modules.scala 160:64:@45154.4]
  assign _T_97150 = $signed(buffer_13_598) + $signed(buffer_13_599); // @[Modules.scala 160:64:@45156.4]
  assign _T_97151 = _T_97150[13:0]; // @[Modules.scala 160:64:@45157.4]
  assign buffer_13_606 = $signed(_T_97151); // @[Modules.scala 160:64:@45158.4]
  assign _T_97153 = $signed(buffer_13_600) + $signed(buffer_13_601); // @[Modules.scala 160:64:@45160.4]
  assign _T_97154 = _T_97153[13:0]; // @[Modules.scala 160:64:@45161.4]
  assign buffer_13_607 = $signed(_T_97154); // @[Modules.scala 160:64:@45162.4]
  assign _T_97156 = $signed(buffer_13_602) + $signed(buffer_13_603); // @[Modules.scala 160:64:@45164.4]
  assign _T_97157 = _T_97156[13:0]; // @[Modules.scala 160:64:@45165.4]
  assign buffer_13_608 = $signed(_T_97157); // @[Modules.scala 160:64:@45166.4]
  assign _T_97159 = $signed(buffer_13_604) + $signed(buffer_13_605); // @[Modules.scala 166:64:@45168.4]
  assign _T_97160 = _T_97159[13:0]; // @[Modules.scala 166:64:@45169.4]
  assign buffer_13_609 = $signed(_T_97160); // @[Modules.scala 166:64:@45170.4]
  assign _T_97162 = $signed(buffer_13_606) + $signed(buffer_13_607); // @[Modules.scala 166:64:@45172.4]
  assign _T_97163 = _T_97162[13:0]; // @[Modules.scala 166:64:@45173.4]
  assign buffer_13_610 = $signed(_T_97163); // @[Modules.scala 166:64:@45174.4]
  assign _T_97165 = $signed(buffer_13_609) + $signed(buffer_13_610); // @[Modules.scala 160:64:@45176.4]
  assign _T_97166 = _T_97165[13:0]; // @[Modules.scala 160:64:@45177.4]
  assign buffer_13_611 = $signed(_T_97166); // @[Modules.scala 160:64:@45178.4]
  assign _T_97168 = $signed(buffer_13_611) + $signed(buffer_13_608); // @[Modules.scala 172:66:@45180.4]
  assign _T_97169 = _T_97168[13:0]; // @[Modules.scala 172:66:@45181.4]
  assign buffer_13_612 = $signed(_T_97169); // @[Modules.scala 172:66:@45182.4]
  assign _GEN_976 = {{1{_T_60257[4]}},_T_60257}; // @[Modules.scala 143:103:@45363.4]
  assign _T_97182 = $signed(_GEN_976) + $signed(_T_54215); // @[Modules.scala 143:103:@45363.4]
  assign _T_97183 = _T_97182[5:0]; // @[Modules.scala 143:103:@45364.4]
  assign _T_97184 = $signed(_T_97183); // @[Modules.scala 143:103:@45365.4]
  assign _GEN_977 = {{1{_T_60332[4]}},_T_60332}; // @[Modules.scala 143:103:@45429.4]
  assign _T_97259 = $signed(_T_63429) + $signed(_GEN_977); // @[Modules.scala 143:103:@45429.4]
  assign _T_97260 = _T_97259[5:0]; // @[Modules.scala 143:103:@45430.4]
  assign _T_97261 = $signed(_T_97260); // @[Modules.scala 143:103:@45431.4]
  assign _T_97273 = $signed(_T_54292) + $signed(_T_54297); // @[Modules.scala 143:103:@45441.4]
  assign _T_97274 = _T_97273[5:0]; // @[Modules.scala 143:103:@45442.4]
  assign _T_97275 = $signed(_T_97274); // @[Modules.scala 143:103:@45443.4]
  assign _T_97280 = $signed(_T_54299) + $signed(_T_54304); // @[Modules.scala 143:103:@45447.4]
  assign _T_97281 = _T_97280[5:0]; // @[Modules.scala 143:103:@45448.4]
  assign _T_97282 = $signed(_T_97281); // @[Modules.scala 143:103:@45449.4]
  assign _T_97287 = $signed(_T_54306) + $signed(_T_54311); // @[Modules.scala 143:103:@45453.4]
  assign _T_97288 = _T_97287[5:0]; // @[Modules.scala 143:103:@45454.4]
  assign _T_97289 = $signed(_T_97288); // @[Modules.scala 143:103:@45455.4]
  assign _T_97294 = $signed(_T_54313) + $signed(_T_54318); // @[Modules.scala 143:103:@45459.4]
  assign _T_97295 = _T_97294[5:0]; // @[Modules.scala 143:103:@45460.4]
  assign _T_97296 = $signed(_T_97295); // @[Modules.scala 143:103:@45461.4]
  assign _T_97301 = $signed(_T_54320) + $signed(_T_54325); // @[Modules.scala 143:103:@45465.4]
  assign _T_97302 = _T_97301[5:0]; // @[Modules.scala 143:103:@45466.4]
  assign _T_97303 = $signed(_T_97302); // @[Modules.scala 143:103:@45467.4]
  assign _T_97308 = $signed(_T_54327) + $signed(_T_54332); // @[Modules.scala 143:103:@45471.4]
  assign _T_97309 = _T_97308[5:0]; // @[Modules.scala 143:103:@45472.4]
  assign _T_97310 = $signed(_T_97309); // @[Modules.scala 143:103:@45473.4]
  assign _GEN_978 = {{1{_T_60404[4]}},_T_60404}; // @[Modules.scala 143:103:@45501.4]
  assign _T_97343 = $signed(_T_54362) + $signed(_GEN_978); // @[Modules.scala 143:103:@45501.4]
  assign _T_97344 = _T_97343[5:0]; // @[Modules.scala 143:103:@45502.4]
  assign _T_97345 = $signed(_T_97344); // @[Modules.scala 143:103:@45503.4]
  assign _GEN_979 = {{1{_T_57379[4]}},_T_57379}; // @[Modules.scala 143:103:@45507.4]
  assign _T_97350 = $signed(_GEN_979) + $signed(_T_54374); // @[Modules.scala 143:103:@45507.4]
  assign _T_97351 = _T_97350[5:0]; // @[Modules.scala 143:103:@45508.4]
  assign _T_97352 = $signed(_T_97351); // @[Modules.scala 143:103:@45509.4]
  assign _T_97420 = $signed(_GEN_2) + $signed(_T_54444); // @[Modules.scala 143:103:@45567.4]
  assign _T_97421 = _T_97420[5:0]; // @[Modules.scala 143:103:@45568.4]
  assign _T_97422 = $signed(_T_97421); // @[Modules.scala 143:103:@45569.4]
  assign _T_97441 = $signed(_T_63599) + $signed(_T_63606); // @[Modules.scala 143:103:@45585.4]
  assign _T_97442 = _T_97441[4:0]; // @[Modules.scala 143:103:@45586.4]
  assign _T_97443 = $signed(_T_97442); // @[Modules.scala 143:103:@45587.4]
  assign _T_97469 = $signed(_T_57498) + $signed(_GEN_507); // @[Modules.scala 143:103:@45609.4]
  assign _T_97470 = _T_97469[5:0]; // @[Modules.scala 143:103:@45610.4]
  assign _T_97471 = $signed(_T_97470); // @[Modules.scala 143:103:@45611.4]
  assign _T_97476 = $signed(_T_54507) + $signed(_T_54514); // @[Modules.scala 143:103:@45615.4]
  assign _T_97477 = _T_97476[4:0]; // @[Modules.scala 143:103:@45616.4]
  assign _T_97478 = $signed(_T_97477); // @[Modules.scala 143:103:@45617.4]
  assign _T_97483 = $signed(_GEN_152) + $signed(_T_54521); // @[Modules.scala 143:103:@45621.4]
  assign _T_97484 = _T_97483[5:0]; // @[Modules.scala 143:103:@45622.4]
  assign _T_97485 = $signed(_T_97484); // @[Modules.scala 143:103:@45623.4]
  assign _T_97518 = $signed(_T_69819) + $signed(_GEN_845); // @[Modules.scala 143:103:@45651.4]
  assign _T_97519 = _T_97518[5:0]; // @[Modules.scala 143:103:@45652.4]
  assign _T_97520 = $signed(_T_97519); // @[Modules.scala 143:103:@45653.4]
  assign _GEN_990 = {{1{_T_63774[4]}},_T_63774}; // @[Modules.scala 143:103:@45705.4]
  assign _T_97581 = $signed(_GEN_990) + $signed(_T_73021); // @[Modules.scala 143:103:@45705.4]
  assign _T_97582 = _T_97581[5:0]; // @[Modules.scala 143:103:@45706.4]
  assign _T_97583 = $signed(_T_97582); // @[Modules.scala 143:103:@45707.4]
  assign _GEN_991 = {{1{_T_54619[4]}},_T_54619}; // @[Modules.scala 143:103:@45717.4]
  assign _T_97595 = $signed(_GEN_991) + $signed(_T_66925); // @[Modules.scala 143:103:@45717.4]
  assign _T_97596 = _T_97595[5:0]; // @[Modules.scala 143:103:@45718.4]
  assign _T_97597 = $signed(_T_97596); // @[Modules.scala 143:103:@45719.4]
  assign _T_97623 = $signed(_T_69938) + $signed(_GEN_15); // @[Modules.scala 143:103:@45741.4]
  assign _T_97624 = _T_97623[5:0]; // @[Modules.scala 143:103:@45742.4]
  assign _T_97625 = $signed(_T_97624); // @[Modules.scala 143:103:@45743.4]
  assign _T_97630 = $signed(_GEN_704) + $signed(_T_54663); // @[Modules.scala 143:103:@45747.4]
  assign _T_97631 = _T_97630[5:0]; // @[Modules.scala 143:103:@45748.4]
  assign _T_97632 = $signed(_T_97631); // @[Modules.scala 143:103:@45749.4]
  assign _T_97651 = $signed(_GEN_587) + $signed(_T_69973); // @[Modules.scala 143:103:@45765.4]
  assign _T_97652 = _T_97651[5:0]; // @[Modules.scala 143:103:@45766.4]
  assign _T_97653 = $signed(_T_97652); // @[Modules.scala 143:103:@45767.4]
  assign _T_97658 = $signed(_T_54689) + $signed(_T_57715); // @[Modules.scala 143:103:@45771.4]
  assign _T_97659 = _T_97658[5:0]; // @[Modules.scala 143:103:@45772.4]
  assign _T_97660 = $signed(_T_97659); // @[Modules.scala 143:103:@45773.4]
  assign _T_97672 = $signed(_T_57738) + $signed(_T_63893); // @[Modules.scala 143:103:@45783.4]
  assign _T_97673 = _T_97672[5:0]; // @[Modules.scala 143:103:@45784.4]
  assign _T_97674 = $signed(_T_97673); // @[Modules.scala 143:103:@45785.4]
  assign _T_97686 = $signed(_T_63905) + $signed(_T_54724); // @[Modules.scala 143:103:@45795.4]
  assign _T_97687 = _T_97686[5:0]; // @[Modules.scala 143:103:@45796.4]
  assign _T_97688 = $signed(_T_97687); // @[Modules.scala 143:103:@45797.4]
  assign _GEN_997 = {{1{_T_60808[4]}},_T_60808}; // @[Modules.scala 143:103:@45807.4]
  assign _T_97700 = $signed(_GEN_997) + $signed(_T_54738); // @[Modules.scala 143:103:@45807.4]
  assign _T_97701 = _T_97700[5:0]; // @[Modules.scala 143:103:@45808.4]
  assign _T_97702 = $signed(_T_97701); // @[Modules.scala 143:103:@45809.4]
  assign _T_97721 = $signed(_T_70059) + $signed(_T_67053); // @[Modules.scala 143:103:@45825.4]
  assign _T_97722 = _T_97721[5:0]; // @[Modules.scala 143:103:@45826.4]
  assign _T_97723 = $signed(_T_97722); // @[Modules.scala 143:103:@45827.4]
  assign _GEN_999 = {{1{_T_60843[4]}},_T_60843}; // @[Modules.scala 143:103:@45831.4]
  assign _T_97728 = $signed(_GEN_999) + $signed(_T_54766); // @[Modules.scala 143:103:@45831.4]
  assign _T_97729 = _T_97728[5:0]; // @[Modules.scala 143:103:@45832.4]
  assign _T_97730 = $signed(_T_97729); // @[Modules.scala 143:103:@45833.4]
  assign _GEN_1000 = {{1{_T_60908[4]}},_T_60908}; // @[Modules.scala 143:103:@45879.4]
  assign _T_97784 = $signed(_T_54822) + $signed(_GEN_1000); // @[Modules.scala 143:103:@45879.4]
  assign _T_97785 = _T_97784[5:0]; // @[Modules.scala 143:103:@45880.4]
  assign _T_97786 = $signed(_T_97785); // @[Modules.scala 143:103:@45881.4]
  assign _GEN_1001 = {{1{_T_54831[4]}},_T_54831}; // @[Modules.scala 143:103:@45885.4]
  assign _T_97791 = $signed(_T_70148) + $signed(_GEN_1001); // @[Modules.scala 143:103:@45885.4]
  assign _T_97792 = _T_97791[5:0]; // @[Modules.scala 143:103:@45886.4]
  assign _T_97793 = $signed(_T_97792); // @[Modules.scala 143:103:@45887.4]
  assign _GEN_1002 = {{1{_T_54859[4]}},_T_54859}; // @[Modules.scala 143:103:@45909.4]
  assign _T_97819 = $signed(_GEN_1002) + $signed(_T_57904); // @[Modules.scala 143:103:@45909.4]
  assign _T_97820 = _T_97819[5:0]; // @[Modules.scala 143:103:@45910.4]
  assign _T_97821 = $signed(_T_97820); // @[Modules.scala 143:103:@45911.4]
  assign _T_97847 = $signed(_T_54894) + $signed(_T_60985); // @[Modules.scala 143:103:@45933.4]
  assign _T_97848 = _T_97847[4:0]; // @[Modules.scala 143:103:@45934.4]
  assign _T_97849 = $signed(_T_97848); // @[Modules.scala 143:103:@45935.4]
  assign _T_97854 = $signed(_T_57941) + $signed(_GEN_860); // @[Modules.scala 143:103:@45939.4]
  assign _T_97855 = _T_97854[5:0]; // @[Modules.scala 143:103:@45940.4]
  assign _T_97856 = $signed(_T_97855); // @[Modules.scala 143:103:@45941.4]
  assign _T_97861 = $signed(_T_54922) + $signed(_T_54934); // @[Modules.scala 143:103:@45945.4]
  assign _T_97862 = _T_97861[4:0]; // @[Modules.scala 143:103:@45946.4]
  assign _T_97863 = $signed(_T_97862); // @[Modules.scala 143:103:@45947.4]
  assign _T_97882 = $signed(_T_54955) + $signed(_T_54962); // @[Modules.scala 143:103:@45963.4]
  assign _T_97883 = _T_97882[4:0]; // @[Modules.scala 143:103:@45964.4]
  assign _T_97884 = $signed(_T_97883); // @[Modules.scala 143:103:@45965.4]
  assign _T_97910 = $signed(_T_64173) + $signed(_T_61062); // @[Modules.scala 143:103:@45987.4]
  assign _T_97911 = _T_97910[4:0]; // @[Modules.scala 143:103:@45988.4]
  assign _T_97912 = $signed(_T_97911); // @[Modules.scala 143:103:@45989.4]
  assign _T_97931 = $signed(_T_58032) + $signed(_GEN_657); // @[Modules.scala 143:103:@46005.4]
  assign _T_97932 = _T_97931[5:0]; // @[Modules.scala 143:103:@46006.4]
  assign _T_97933 = $signed(_T_97932); // @[Modules.scala 143:103:@46007.4]
  assign _GEN_1006 = {{1{_T_55039[4]}},_T_55039}; // @[Modules.scala 143:103:@46029.4]
  assign _T_97959 = $signed(_T_58058) + $signed(_GEN_1006); // @[Modules.scala 143:103:@46029.4]
  assign _T_97960 = _T_97959[5:0]; // @[Modules.scala 143:103:@46030.4]
  assign _T_97961 = $signed(_T_97960); // @[Modules.scala 143:103:@46031.4]
  assign _T_97987 = $signed(_T_70353) + $signed(_T_64262); // @[Modules.scala 143:103:@46053.4]
  assign _T_97988 = _T_97987[5:0]; // @[Modules.scala 143:103:@46054.4]
  assign _T_97989 = $signed(_T_97988); // @[Modules.scala 143:103:@46055.4]
  assign _GEN_1008 = {{1{_T_55097[4]}},_T_55097}; // @[Modules.scala 143:103:@46077.4]
  assign _T_98015 = $signed(_T_61160) + $signed(_GEN_1008); // @[Modules.scala 143:103:@46077.4]
  assign _T_98016 = _T_98015[5:0]; // @[Modules.scala 143:103:@46078.4]
  assign _T_98017 = $signed(_T_98016); // @[Modules.scala 143:103:@46079.4]
  assign _T_98057 = $signed(_T_76696) + $signed(_T_64334); // @[Modules.scala 143:103:@46113.4]
  assign _T_98058 = _T_98057[4:0]; // @[Modules.scala 143:103:@46114.4]
  assign _T_98059 = $signed(_T_98058); // @[Modules.scala 143:103:@46115.4]
  assign _T_98085 = $signed(_T_58193) + $signed(_T_55179); // @[Modules.scala 143:103:@46137.4]
  assign _T_98086 = _T_98085[4:0]; // @[Modules.scala 143:103:@46138.4]
  assign _T_98087 = $signed(_T_98086); // @[Modules.scala 143:103:@46139.4]
  assign _T_98092 = $signed(_GEN_466) + $signed(_T_58207); // @[Modules.scala 143:103:@46143.4]
  assign _T_98093 = _T_98092[5:0]; // @[Modules.scala 143:103:@46144.4]
  assign _T_98094 = $signed(_T_98093); // @[Modules.scala 143:103:@46145.4]
  assign _T_98099 = $signed(_T_61265) + $signed(_T_61272); // @[Modules.scala 143:103:@46149.4]
  assign _T_98100 = _T_98099[5:0]; // @[Modules.scala 143:103:@46150.4]
  assign _T_98101 = $signed(_T_98100); // @[Modules.scala 143:103:@46151.4]
  assign _T_98127 = $signed(_T_55223) + $signed(_T_58254); // @[Modules.scala 143:103:@46173.4]
  assign _T_98128 = _T_98127[4:0]; // @[Modules.scala 143:103:@46174.4]
  assign _T_98129 = $signed(_T_98128); // @[Modules.scala 143:103:@46175.4]
  assign _GEN_1013 = {{1{_T_70533[4]}},_T_70533}; // @[Modules.scala 143:103:@46197.4]
  assign _T_98155 = $signed(_T_58282) + $signed(_GEN_1013); // @[Modules.scala 143:103:@46197.4]
  assign _T_98156 = _T_98155[5:0]; // @[Modules.scala 143:103:@46198.4]
  assign _T_98157 = $signed(_T_98156); // @[Modules.scala 143:103:@46199.4]
  assign _GEN_1014 = {{1{_T_55270[4]}},_T_55270}; // @[Modules.scala 143:103:@46209.4]
  assign _T_98169 = $signed(_GEN_1014) + $signed(_T_61354); // @[Modules.scala 143:103:@46209.4]
  assign _T_98170 = _T_98169[5:0]; // @[Modules.scala 143:103:@46210.4]
  assign _T_98171 = $signed(_T_98170); // @[Modules.scala 143:103:@46211.4]
  assign _GEN_1015 = {{1{_T_55286[4]}},_T_55286}; // @[Modules.scala 143:103:@46215.4]
  assign _T_98176 = $signed(_T_58296) + $signed(_GEN_1015); // @[Modules.scala 143:103:@46215.4]
  assign _T_98177 = _T_98176[5:0]; // @[Modules.scala 143:103:@46216.4]
  assign _T_98178 = $signed(_T_98177); // @[Modules.scala 143:103:@46217.4]
  assign _T_98183 = $signed(_GEN_39) + $signed(_T_58310); // @[Modules.scala 143:103:@46221.4]
  assign _T_98184 = _T_98183[5:0]; // @[Modules.scala 143:103:@46222.4]
  assign _T_98185 = $signed(_T_98184); // @[Modules.scala 143:103:@46223.4]
  assign _T_98190 = $signed(_T_55293) + $signed(_GEN_390); // @[Modules.scala 143:103:@46227.4]
  assign _T_98191 = _T_98190[5:0]; // @[Modules.scala 143:103:@46228.4]
  assign _T_98192 = $signed(_T_98191); // @[Modules.scala 143:103:@46229.4]
  assign _T_98211 = $signed(_T_58326) + $signed(_T_58333); // @[Modules.scala 143:103:@46245.4]
  assign _T_98212 = _T_98211[4:0]; // @[Modules.scala 143:103:@46246.4]
  assign _T_98213 = $signed(_T_98212); // @[Modules.scala 143:103:@46247.4]
  assign _T_98239 = $signed(_T_61419) + $signed(_GEN_321); // @[Modules.scala 143:103:@46269.4]
  assign _T_98240 = _T_98239[5:0]; // @[Modules.scala 143:103:@46270.4]
  assign _T_98241 = $signed(_T_98240); // @[Modules.scala 143:103:@46271.4]
  assign _T_98260 = $signed(_GEN_726) + $signed(_T_61445); // @[Modules.scala 143:103:@46287.4]
  assign _T_98261 = _T_98260[5:0]; // @[Modules.scala 143:103:@46288.4]
  assign _T_98262 = $signed(_T_98261); // @[Modules.scala 143:103:@46289.4]
  assign _T_98302 = $signed(_T_55396) + $signed(_T_83183); // @[Modules.scala 143:103:@46323.4]
  assign _T_98303 = _T_98302[5:0]; // @[Modules.scala 143:103:@46324.4]
  assign _T_98304 = $signed(_T_98303); // @[Modules.scala 143:103:@46325.4]
  assign _T_98309 = $signed(_T_61489) + $signed(_GEN_664); // @[Modules.scala 143:103:@46329.4]
  assign _T_98310 = _T_98309[5:0]; // @[Modules.scala 143:103:@46330.4]
  assign _T_98311 = $signed(_T_98310); // @[Modules.scala 143:103:@46331.4]
  assign _T_98344 = $signed(_GEN_731) + $signed(_T_55445); // @[Modules.scala 143:103:@46359.4]
  assign _T_98345 = _T_98344[5:0]; // @[Modules.scala 143:103:@46360.4]
  assign _T_98346 = $signed(_T_98345); // @[Modules.scala 143:103:@46361.4]
  assign _T_98358 = $signed(_T_55452) + $signed(_GEN_876); // @[Modules.scala 143:103:@46371.4]
  assign _T_98359 = _T_98358[5:0]; // @[Modules.scala 143:103:@46372.4]
  assign _T_98360 = $signed(_T_98359); // @[Modules.scala 143:103:@46373.4]
  assign _T_98372 = $signed(_T_55466) + $signed(_T_64675); // @[Modules.scala 143:103:@46383.4]
  assign _T_98373 = _T_98372[4:0]; // @[Modules.scala 143:103:@46384.4]
  assign _T_98374 = $signed(_T_98373); // @[Modules.scala 143:103:@46385.4]
  assign _T_98393 = $signed(_T_61578) + $signed(_T_70780); // @[Modules.scala 143:103:@46401.4]
  assign _T_98394 = _T_98393[4:0]; // @[Modules.scala 143:103:@46402.4]
  assign _T_98395 = $signed(_T_98394); // @[Modules.scala 143:103:@46403.4]
  assign _T_98407 = $signed(_T_55494) + $signed(_GEN_185); // @[Modules.scala 143:103:@46413.4]
  assign _T_98408 = _T_98407[5:0]; // @[Modules.scala 143:103:@46414.4]
  assign _T_98409 = $signed(_T_98408); // @[Modules.scala 143:103:@46415.4]
  assign _T_98421 = $signed(_T_55510) + $signed(_GEN_473); // @[Modules.scala 143:103:@46425.4]
  assign _T_98422 = _T_98421[5:0]; // @[Modules.scala 143:103:@46426.4]
  assign _T_98423 = $signed(_T_98422); // @[Modules.scala 143:103:@46427.4]
  assign _T_98442 = $signed(_GEN_55) + $signed(_T_67765); // @[Modules.scala 143:103:@46443.4]
  assign _T_98443 = _T_98442[5:0]; // @[Modules.scala 143:103:@46444.4]
  assign _T_98444 = $signed(_T_98443); // @[Modules.scala 143:103:@46445.4]
  assign _T_98449 = $signed(_T_67767) + $signed(_GEN_186); // @[Modules.scala 143:103:@46449.4]
  assign _T_98450 = _T_98449[5:0]; // @[Modules.scala 143:103:@46450.4]
  assign _T_98451 = $signed(_T_98450); // @[Modules.scala 143:103:@46451.4]
  assign _T_98491 = $signed(_T_64796) + $signed(_T_55592); // @[Modules.scala 143:103:@46485.4]
  assign _T_98492 = _T_98491[5:0]; // @[Modules.scala 143:103:@46486.4]
  assign _T_98493 = $signed(_T_98492); // @[Modules.scala 143:103:@46487.4]
  assign _T_98498 = $signed(_T_55594) + $signed(_GEN_408); // @[Modules.scala 143:103:@46491.4]
  assign _T_98499 = _T_98498[5:0]; // @[Modules.scala 143:103:@46492.4]
  assign _T_98500 = $signed(_T_98499); // @[Modules.scala 143:103:@46493.4]
  assign _T_98512 = $signed(_T_55615) + $signed(_T_70911); // @[Modules.scala 143:103:@46503.4]
  assign _T_98513 = _T_98512[5:0]; // @[Modules.scala 143:103:@46504.4]
  assign _T_98514 = $signed(_T_98513); // @[Modules.scala 143:103:@46505.4]
  assign _T_98533 = $signed(_T_55629) + $signed(_GEN_191); // @[Modules.scala 143:103:@46521.4]
  assign _T_98534 = _T_98533[5:0]; // @[Modules.scala 143:103:@46522.4]
  assign _T_98535 = $signed(_T_98534); // @[Modules.scala 143:103:@46523.4]
  assign _GEN_1038 = {{1{_T_61739[4]}},_T_61739}; // @[Modules.scala 143:103:@46533.4]
  assign _T_98547 = $signed(_T_55655) + $signed(_GEN_1038); // @[Modules.scala 143:103:@46533.4]
  assign _T_98548 = _T_98547[5:0]; // @[Modules.scala 143:103:@46534.4]
  assign _T_98549 = $signed(_T_98548); // @[Modules.scala 143:103:@46535.4]
  assign _GEN_1039 = {{1{_T_61741[4]}},_T_61741}; // @[Modules.scala 143:103:@46539.4]
  assign _T_98554 = $signed(_GEN_1039) + $signed(_T_55664); // @[Modules.scala 143:103:@46539.4]
  assign _T_98555 = _T_98554[5:0]; // @[Modules.scala 143:103:@46540.4]
  assign _T_98556 = $signed(_T_98555); // @[Modules.scala 143:103:@46541.4]
  assign _T_98568 = $signed(_T_55671) + $signed(_T_55676); // @[Modules.scala 143:103:@46551.4]
  assign _T_98569 = _T_98568[5:0]; // @[Modules.scala 143:103:@46552.4]
  assign _T_98570 = $signed(_T_98569); // @[Modules.scala 143:103:@46553.4]
  assign _T_98610 = $signed(_T_55711) + $signed(_T_71002); // @[Modules.scala 143:103:@46587.4]
  assign _T_98611 = _T_98610[5:0]; // @[Modules.scala 143:103:@46588.4]
  assign _T_98612 = $signed(_T_98611); // @[Modules.scala 143:103:@46589.4]
  assign _T_98729 = $signed(_T_61895) + $signed(_T_61902); // @[Modules.scala 143:103:@46689.4]
  assign _T_98730 = _T_98729[4:0]; // @[Modules.scala 143:103:@46690.4]
  assign _T_98731 = $signed(_T_98730); // @[Modules.scala 143:103:@46691.4]
  assign _T_98743 = $signed(_T_55816) + $signed(_T_77464); // @[Modules.scala 143:103:@46701.4]
  assign _T_98744 = _T_98743[5:0]; // @[Modules.scala 143:103:@46702.4]
  assign _T_98745 = $signed(_T_98744); // @[Modules.scala 143:103:@46703.4]
  assign _T_98750 = $signed(_T_55818) + $signed(_T_55823); // @[Modules.scala 143:103:@46707.4]
  assign _T_98751 = _T_98750[5:0]; // @[Modules.scala 143:103:@46708.4]
  assign _T_98752 = $signed(_T_98751); // @[Modules.scala 143:103:@46709.4]
  assign _T_98757 = $signed(_T_61923) + $signed(_T_55825); // @[Modules.scala 143:103:@46713.4]
  assign _T_98758 = _T_98757[5:0]; // @[Modules.scala 143:103:@46714.4]
  assign _T_98759 = $signed(_T_98758); // @[Modules.scala 143:103:@46715.4]
  assign _T_98778 = $signed(_T_74330) + $signed(_T_58858); // @[Modules.scala 143:103:@46731.4]
  assign _T_98779 = _T_98778[5:0]; // @[Modules.scala 143:103:@46732.4]
  assign _T_98780 = $signed(_T_98779); // @[Modules.scala 143:103:@46733.4]
  assign _GEN_1045 = {{1{_T_58872[4]}},_T_58872}; // @[Modules.scala 143:103:@46743.4]
  assign _T_98792 = $signed(_T_55844) + $signed(_GEN_1045); // @[Modules.scala 143:103:@46743.4]
  assign _T_98793 = _T_98792[5:0]; // @[Modules.scala 143:103:@46744.4]
  assign _T_98794 = $signed(_T_98793); // @[Modules.scala 143:103:@46745.4]
  assign _T_98799 = $signed(_GEN_201) + $signed(_T_55853); // @[Modules.scala 143:103:@46749.4]
  assign _T_98800 = _T_98799[5:0]; // @[Modules.scala 143:103:@46750.4]
  assign _T_98801 = $signed(_T_98800); // @[Modules.scala 143:103:@46751.4]
  assign _T_98813 = $signed(_T_58891) + $signed(_T_61979); // @[Modules.scala 143:103:@46761.4]
  assign _T_98814 = _T_98813[4:0]; // @[Modules.scala 143:103:@46762.4]
  assign _T_98815 = $signed(_T_98814); // @[Modules.scala 143:103:@46763.4]
  assign _T_98834 = $signed(_GEN_617) + $signed(_T_58919); // @[Modules.scala 143:103:@46779.4]
  assign _T_98835 = _T_98834[5:0]; // @[Modules.scala 143:103:@46780.4]
  assign _T_98836 = $signed(_T_98835); // @[Modules.scala 143:103:@46781.4]
  assign _T_98848 = $signed(_T_71242) + $signed(_T_71247); // @[Modules.scala 143:103:@46791.4]
  assign _T_98849 = _T_98848[5:0]; // @[Modules.scala 143:103:@46792.4]
  assign _T_98850 = $signed(_T_98849); // @[Modules.scala 143:103:@46793.4]
  assign _T_98855 = $signed(_T_65125) + $signed(_T_65130); // @[Modules.scala 143:103:@46797.4]
  assign _T_98856 = _T_98855[5:0]; // @[Modules.scala 143:103:@46798.4]
  assign _T_98857 = $signed(_T_98856); // @[Modules.scala 143:103:@46799.4]
  assign _GEN_1048 = {{1{_T_58947[4]}},_T_58947}; // @[Modules.scala 143:103:@46815.4]
  assign _T_98876 = $signed(_T_55928) + $signed(_GEN_1048); // @[Modules.scala 143:103:@46815.4]
  assign _T_98877 = _T_98876[5:0]; // @[Modules.scala 143:103:@46816.4]
  assign _T_98878 = $signed(_T_98877); // @[Modules.scala 143:103:@46817.4]
  assign _T_98890 = $signed(_GEN_344) + $signed(_T_55944); // @[Modules.scala 143:103:@46827.4]
  assign _T_98891 = _T_98890[5:0]; // @[Modules.scala 143:103:@46828.4]
  assign _T_98892 = $signed(_T_98891); // @[Modules.scala 143:103:@46829.4]
  assign _T_98925 = $signed(_T_68220) + $signed(_T_58984); // @[Modules.scala 143:103:@46857.4]
  assign _T_98926 = _T_98925[5:0]; // @[Modules.scala 143:103:@46858.4]
  assign _T_98927 = $signed(_T_98926); // @[Modules.scala 143:103:@46859.4]
  assign _GEN_1050 = {{1{_T_59017[4]}},_T_59017}; // @[Modules.scala 143:103:@46887.4]
  assign _T_98960 = $signed(_T_62110) + $signed(_GEN_1050); // @[Modules.scala 143:103:@46887.4]
  assign _T_98961 = _T_98960[5:0]; // @[Modules.scala 143:103:@46888.4]
  assign _T_98962 = $signed(_T_98961); // @[Modules.scala 143:103:@46889.4]
  assign _GEN_1051 = {{1{_T_62145[4]}},_T_62145}; // @[Modules.scala 143:103:@46911.4]
  assign _T_98988 = $signed(_GEN_1051) + $signed(_T_56047); // @[Modules.scala 143:103:@46911.4]
  assign _T_98989 = _T_98988[5:0]; // @[Modules.scala 143:103:@46912.4]
  assign _T_98990 = $signed(_T_98989); // @[Modules.scala 143:103:@46913.4]
  assign _T_99023 = $signed(_T_59080) + $signed(_GEN_690); // @[Modules.scala 143:103:@46941.4]
  assign _T_99024 = _T_99023[5:0]; // @[Modules.scala 143:103:@46942.4]
  assign _T_99025 = $signed(_T_99024); // @[Modules.scala 143:103:@46943.4]
  assign _GEN_1053 = {{1{_T_56084[4]}},_T_56084}; // @[Modules.scala 143:103:@46947.4]
  assign _T_99030 = $signed(_T_59089) + $signed(_GEN_1053); // @[Modules.scala 143:103:@46947.4]
  assign _T_99031 = _T_99030[5:0]; // @[Modules.scala 143:103:@46948.4]
  assign _T_99032 = $signed(_T_99031); // @[Modules.scala 143:103:@46949.4]
  assign _T_99044 = $signed(_T_56096) + $signed(_T_59108); // @[Modules.scala 143:103:@46959.4]
  assign _T_99045 = _T_99044[4:0]; // @[Modules.scala 143:103:@46960.4]
  assign _T_99046 = $signed(_T_99045); // @[Modules.scala 143:103:@46961.4]
  assign _T_99107 = $signed(_T_59164) + $signed(_GEN_277); // @[Modules.scala 143:103:@47013.4]
  assign _T_99108 = _T_99107[5:0]; // @[Modules.scala 143:103:@47014.4]
  assign _T_99109 = $signed(_T_99108); // @[Modules.scala 143:103:@47015.4]
  assign _T_99128 = $signed(_T_65382) + $signed(_T_68423); // @[Modules.scala 143:103:@47031.4]
  assign _T_99129 = _T_99128[5:0]; // @[Modules.scala 143:103:@47032.4]
  assign _T_99130 = $signed(_T_99129); // @[Modules.scala 143:103:@47033.4]
  assign _T_99219 = $signed(_T_59264) + $signed(_T_56250); // @[Modules.scala 143:103:@47109.4]
  assign _T_99220 = _T_99219[5:0]; // @[Modules.scala 143:103:@47110.4]
  assign _T_99221 = $signed(_T_99220); // @[Modules.scala 143:103:@47111.4]
  assign _T_99233 = $signed(_T_68523) + $signed(_T_59278); // @[Modules.scala 143:103:@47121.4]
  assign _T_99234 = _T_99233[5:0]; // @[Modules.scala 143:103:@47122.4]
  assign _T_99235 = $signed(_T_99234); // @[Modules.scala 143:103:@47123.4]
  assign _GEN_1057 = {{1{_T_62376[4]}},_T_62376}; // @[Modules.scala 143:103:@47127.4]
  assign _T_99240 = $signed(_T_56264) + $signed(_GEN_1057); // @[Modules.scala 143:103:@47127.4]
  assign _T_99241 = _T_99240[5:0]; // @[Modules.scala 143:103:@47128.4]
  assign _T_99242 = $signed(_T_99241); // @[Modules.scala 143:103:@47129.4]
  assign _T_99247 = $signed(_T_59290) + $signed(_T_62385); // @[Modules.scala 143:103:@47133.4]
  assign _T_99248 = _T_99247[4:0]; // @[Modules.scala 143:103:@47134.4]
  assign _T_99249 = $signed(_T_99248); // @[Modules.scala 143:103:@47135.4]
  assign _T_99275 = $signed(_T_56294) + $signed(_T_65529); // @[Modules.scala 143:103:@47157.4]
  assign _T_99276 = _T_99275[4:0]; // @[Modules.scala 143:103:@47158.4]
  assign _T_99277 = $signed(_T_99276); // @[Modules.scala 143:103:@47159.4]
  assign buffer_14_1 = {{8{_T_97184[5]}},_T_97184}; // @[Modules.scala 112:22:@8.4]
  assign _T_99285 = $signed(buffer_10_0) + $signed(buffer_14_1); // @[Modules.scala 160:64:@47167.4]
  assign _T_99286 = _T_99285[13:0]; // @[Modules.scala 160:64:@47168.4]
  assign buffer_14_302 = $signed(_T_99286); // @[Modules.scala 160:64:@47169.4]
  assign _T_99288 = $signed(buffer_11_3) + $signed(buffer_10_3); // @[Modules.scala 160:64:@47171.4]
  assign _T_99289 = _T_99288[13:0]; // @[Modules.scala 160:64:@47172.4]
  assign buffer_14_303 = $signed(_T_99289); // @[Modules.scala 160:64:@47173.4]
  assign buffer_14_12 = {{8{_T_97261[5]}},_T_97261}; // @[Modules.scala 112:22:@8.4]
  assign _T_99303 = $signed(buffer_14_12) + $signed(buffer_7_13); // @[Modules.scala 160:64:@47191.4]
  assign _T_99304 = _T_99303[13:0]; // @[Modules.scala 160:64:@47192.4]
  assign buffer_14_308 = $signed(_T_99304); // @[Modules.scala 160:64:@47193.4]
  assign buffer_14_14 = {{8{_T_97275[5]}},_T_97275}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_15 = {{8{_T_97282[5]}},_T_97282}; // @[Modules.scala 112:22:@8.4]
  assign _T_99306 = $signed(buffer_14_14) + $signed(buffer_14_15); // @[Modules.scala 160:64:@47195.4]
  assign _T_99307 = _T_99306[13:0]; // @[Modules.scala 160:64:@47196.4]
  assign buffer_14_309 = $signed(_T_99307); // @[Modules.scala 160:64:@47197.4]
  assign buffer_14_16 = {{8{_T_97289[5]}},_T_97289}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_17 = {{8{_T_97296[5]}},_T_97296}; // @[Modules.scala 112:22:@8.4]
  assign _T_99309 = $signed(buffer_14_16) + $signed(buffer_14_17); // @[Modules.scala 160:64:@47199.4]
  assign _T_99310 = _T_99309[13:0]; // @[Modules.scala 160:64:@47200.4]
  assign buffer_14_310 = $signed(_T_99310); // @[Modules.scala 160:64:@47201.4]
  assign buffer_14_18 = {{8{_T_97303[5]}},_T_97303}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_19 = {{8{_T_97310[5]}},_T_97310}; // @[Modules.scala 112:22:@8.4]
  assign _T_99312 = $signed(buffer_14_18) + $signed(buffer_14_19); // @[Modules.scala 160:64:@47203.4]
  assign _T_99313 = _T_99312[13:0]; // @[Modules.scala 160:64:@47204.4]
  assign buffer_14_311 = $signed(_T_99313); // @[Modules.scala 160:64:@47205.4]
  assign _T_99318 = $signed(buffer_1_21) + $signed(buffer_7_22); // @[Modules.scala 160:64:@47211.4]
  assign _T_99319 = _T_99318[13:0]; // @[Modules.scala 160:64:@47212.4]
  assign buffer_14_313 = $signed(_T_99319); // @[Modules.scala 160:64:@47213.4]
  assign buffer_14_24 = {{8{_T_97345[5]}},_T_97345}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_25 = {{8{_T_97352[5]}},_T_97352}; // @[Modules.scala 112:22:@8.4]
  assign _T_99321 = $signed(buffer_14_24) + $signed(buffer_14_25); // @[Modules.scala 160:64:@47215.4]
  assign _T_99322 = _T_99321[13:0]; // @[Modules.scala 160:64:@47216.4]
  assign buffer_14_314 = $signed(_T_99322); // @[Modules.scala 160:64:@47217.4]
  assign _T_99324 = $signed(buffer_10_25) + $signed(buffer_6_26); // @[Modules.scala 160:64:@47219.4]
  assign _T_99325 = _T_99324[13:0]; // @[Modules.scala 160:64:@47220.4]
  assign buffer_14_315 = $signed(_T_99325); // @[Modules.scala 160:64:@47221.4]
  assign _T_99327 = $signed(buffer_10_27) + $signed(buffer_9_29); // @[Modules.scala 160:64:@47223.4]
  assign _T_99328 = _T_99327[13:0]; // @[Modules.scala 160:64:@47224.4]
  assign buffer_14_316 = $signed(_T_99328); // @[Modules.scala 160:64:@47225.4]
  assign buffer_14_35 = {{8{_T_97422[5]}},_T_97422}; // @[Modules.scala 112:22:@8.4]
  assign _T_99336 = $signed(buffer_7_33) + $signed(buffer_14_35); // @[Modules.scala 160:64:@47235.4]
  assign _T_99337 = _T_99336[13:0]; // @[Modules.scala 160:64:@47236.4]
  assign buffer_14_319 = $signed(_T_99337); // @[Modules.scala 160:64:@47237.4]
  assign _T_99339 = $signed(buffer_5_34) + $signed(buffer_4_35); // @[Modules.scala 160:64:@47239.4]
  assign _T_99340 = _T_99339[13:0]; // @[Modules.scala 160:64:@47240.4]
  assign buffer_14_320 = $signed(_T_99340); // @[Modules.scala 160:64:@47241.4]
  assign buffer_14_38 = {{9{_T_97443[4]}},_T_97443}; // @[Modules.scala 112:22:@8.4]
  assign _T_99342 = $signed(buffer_14_38) + $signed(buffer_10_40); // @[Modules.scala 160:64:@47243.4]
  assign _T_99343 = _T_99342[13:0]; // @[Modules.scala 160:64:@47244.4]
  assign buffer_14_321 = $signed(_T_99343); // @[Modules.scala 160:64:@47245.4]
  assign _T_99345 = $signed(buffer_8_41) + $signed(buffer_0_42); // @[Modules.scala 160:64:@47247.4]
  assign _T_99346 = _T_99345[13:0]; // @[Modules.scala 160:64:@47248.4]
  assign buffer_14_322 = $signed(_T_99346); // @[Modules.scala 160:64:@47249.4]
  assign buffer_14_42 = {{8{_T_97471[5]}},_T_97471}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_43 = {{9{_T_97478[4]}},_T_97478}; // @[Modules.scala 112:22:@8.4]
  assign _T_99348 = $signed(buffer_14_42) + $signed(buffer_14_43); // @[Modules.scala 160:64:@47251.4]
  assign _T_99349 = _T_99348[13:0]; // @[Modules.scala 160:64:@47252.4]
  assign buffer_14_323 = $signed(_T_99349); // @[Modules.scala 160:64:@47253.4]
  assign buffer_14_44 = {{8{_T_97485[5]}},_T_97485}; // @[Modules.scala 112:22:@8.4]
  assign _T_99351 = $signed(buffer_14_44) + $signed(buffer_2_45); // @[Modules.scala 160:64:@47255.4]
  assign _T_99352 = _T_99351[13:0]; // @[Modules.scala 160:64:@47256.4]
  assign buffer_14_324 = $signed(_T_99352); // @[Modules.scala 160:64:@47257.4]
  assign buffer_14_49 = {{8{_T_97520[5]}},_T_97520}; // @[Modules.scala 112:22:@8.4]
  assign _T_99357 = $signed(buffer_1_49) + $signed(buffer_14_49); // @[Modules.scala 160:64:@47263.4]
  assign _T_99358 = _T_99357[13:0]; // @[Modules.scala 160:64:@47264.4]
  assign buffer_14_326 = $signed(_T_99358); // @[Modules.scala 160:64:@47265.4]
  assign _T_99366 = $signed(buffer_0_53) + $signed(buffer_11_56); // @[Modules.scala 160:64:@47275.4]
  assign _T_99367 = _T_99366[13:0]; // @[Modules.scala 160:64:@47276.4]
  assign buffer_14_329 = $signed(_T_99367); // @[Modules.scala 160:64:@47277.4]
  assign buffer_14_58 = {{8{_T_97583[5]}},_T_97583}; // @[Modules.scala 112:22:@8.4]
  assign _T_99372 = $signed(buffer_14_58) + $signed(buffer_1_60); // @[Modules.scala 160:64:@47283.4]
  assign _T_99373 = _T_99372[13:0]; // @[Modules.scala 160:64:@47284.4]
  assign buffer_14_331 = $signed(_T_99373); // @[Modules.scala 160:64:@47285.4]
  assign buffer_14_60 = {{8{_T_97597[5]}},_T_97597}; // @[Modules.scala 112:22:@8.4]
  assign _T_99375 = $signed(buffer_14_60) + $signed(buffer_11_62); // @[Modules.scala 160:64:@47287.4]
  assign _T_99376 = _T_99375[13:0]; // @[Modules.scala 160:64:@47288.4]
  assign buffer_14_332 = $signed(_T_99376); // @[Modules.scala 160:64:@47289.4]
  assign _T_99378 = $signed(buffer_2_64) + $signed(buffer_3_68); // @[Modules.scala 160:64:@47291.4]
  assign _T_99379 = _T_99378[13:0]; // @[Modules.scala 160:64:@47292.4]
  assign buffer_14_333 = $signed(_T_99379); // @[Modules.scala 160:64:@47293.4]
  assign buffer_14_64 = {{8{_T_97625[5]}},_T_97625}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_65 = {{8{_T_97632[5]}},_T_97632}; // @[Modules.scala 112:22:@8.4]
  assign _T_99381 = $signed(buffer_14_64) + $signed(buffer_14_65); // @[Modules.scala 160:64:@47295.4]
  assign _T_99382 = _T_99381[13:0]; // @[Modules.scala 160:64:@47296.4]
  assign buffer_14_334 = $signed(_T_99382); // @[Modules.scala 160:64:@47297.4]
  assign _T_99384 = $signed(buffer_2_67) + $signed(buffer_2_68); // @[Modules.scala 160:64:@47299.4]
  assign _T_99385 = _T_99384[13:0]; // @[Modules.scala 160:64:@47300.4]
  assign buffer_14_335 = $signed(_T_99385); // @[Modules.scala 160:64:@47301.4]
  assign buffer_14_68 = {{8{_T_97653[5]}},_T_97653}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_69 = {{8{_T_97660[5]}},_T_97660}; // @[Modules.scala 112:22:@8.4]
  assign _T_99387 = $signed(buffer_14_68) + $signed(buffer_14_69); // @[Modules.scala 160:64:@47303.4]
  assign _T_99388 = _T_99387[13:0]; // @[Modules.scala 160:64:@47304.4]
  assign buffer_14_336 = $signed(_T_99388); // @[Modules.scala 160:64:@47305.4]
  assign buffer_14_71 = {{8{_T_97674[5]}},_T_97674}; // @[Modules.scala 112:22:@8.4]
  assign _T_99390 = $signed(buffer_6_74) + $signed(buffer_14_71); // @[Modules.scala 160:64:@47307.4]
  assign _T_99391 = _T_99390[13:0]; // @[Modules.scala 160:64:@47308.4]
  assign buffer_14_337 = $signed(_T_99391); // @[Modules.scala 160:64:@47309.4]
  assign buffer_14_73 = {{8{_T_97688[5]}},_T_97688}; // @[Modules.scala 112:22:@8.4]
  assign _T_99393 = $signed(buffer_3_79) + $signed(buffer_14_73); // @[Modules.scala 160:64:@47311.4]
  assign _T_99394 = _T_99393[13:0]; // @[Modules.scala 160:64:@47312.4]
  assign buffer_14_338 = $signed(_T_99394); // @[Modules.scala 160:64:@47313.4]
  assign buffer_14_75 = {{8{_T_97702[5]}},_T_97702}; // @[Modules.scala 112:22:@8.4]
  assign _T_99396 = $signed(buffer_8_74) + $signed(buffer_14_75); // @[Modules.scala 160:64:@47315.4]
  assign _T_99397 = _T_99396[13:0]; // @[Modules.scala 160:64:@47316.4]
  assign buffer_14_339 = $signed(_T_99397); // @[Modules.scala 160:64:@47317.4]
  assign _T_99399 = $signed(buffer_2_81) + $signed(buffer_8_77); // @[Modules.scala 160:64:@47319.4]
  assign _T_99400 = _T_99399[13:0]; // @[Modules.scala 160:64:@47320.4]
  assign buffer_14_340 = $signed(_T_99400); // @[Modules.scala 160:64:@47321.4]
  assign buffer_14_78 = {{8{_T_97723[5]}},_T_97723}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_79 = {{8{_T_97730[5]}},_T_97730}; // @[Modules.scala 112:22:@8.4]
  assign _T_99402 = $signed(buffer_14_78) + $signed(buffer_14_79); // @[Modules.scala 160:64:@47323.4]
  assign _T_99403 = _T_99402[13:0]; // @[Modules.scala 160:64:@47324.4]
  assign buffer_14_341 = $signed(_T_99403); // @[Modules.scala 160:64:@47325.4]
  assign _T_99405 = $signed(buffer_1_85) + $signed(buffer_11_80); // @[Modules.scala 160:64:@47327.4]
  assign _T_99406 = _T_99405[13:0]; // @[Modules.scala 160:64:@47328.4]
  assign buffer_14_342 = $signed(_T_99406); // @[Modules.scala 160:64:@47329.4]
  assign _T_99411 = $signed(buffer_8_85) + $signed(buffer_8_86); // @[Modules.scala 160:64:@47335.4]
  assign _T_99412 = _T_99411[13:0]; // @[Modules.scala 160:64:@47336.4]
  assign buffer_14_344 = $signed(_T_99412); // @[Modules.scala 160:64:@47337.4]
  assign buffer_14_87 = {{8{_T_97786[5]}},_T_97786}; // @[Modules.scala 112:22:@8.4]
  assign _T_99414 = $signed(buffer_2_93) + $signed(buffer_14_87); // @[Modules.scala 160:64:@47339.4]
  assign _T_99415 = _T_99414[13:0]; // @[Modules.scala 160:64:@47340.4]
  assign buffer_14_345 = $signed(_T_99415); // @[Modules.scala 160:64:@47341.4]
  assign buffer_14_88 = {{8{_T_97793[5]}},_T_97793}; // @[Modules.scala 112:22:@8.4]
  assign _T_99417 = $signed(buffer_14_88) + $signed(buffer_2_97); // @[Modules.scala 160:64:@47343.4]
  assign _T_99418 = _T_99417[13:0]; // @[Modules.scala 160:64:@47344.4]
  assign buffer_14_346 = $signed(_T_99418); // @[Modules.scala 160:64:@47345.4]
  assign buffer_14_92 = {{8{_T_97821[5]}},_T_97821}; // @[Modules.scala 112:22:@8.4]
  assign _T_99423 = $signed(buffer_14_92) + $signed(buffer_5_104); // @[Modules.scala 160:64:@47351.4]
  assign _T_99424 = _T_99423[13:0]; // @[Modules.scala 160:64:@47352.4]
  assign buffer_14_348 = $signed(_T_99424); // @[Modules.scala 160:64:@47353.4]
  assign _T_99426 = $signed(buffer_5_105) + $signed(buffer_5_106); // @[Modules.scala 160:64:@47355.4]
  assign _T_99427 = _T_99426[13:0]; // @[Modules.scala 160:64:@47356.4]
  assign buffer_14_349 = $signed(_T_99427); // @[Modules.scala 160:64:@47357.4]
  assign buffer_14_96 = {{9{_T_97849[4]}},_T_97849}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_97 = {{8{_T_97856[5]}},_T_97856}; // @[Modules.scala 112:22:@8.4]
  assign _T_99429 = $signed(buffer_14_96) + $signed(buffer_14_97); // @[Modules.scala 160:64:@47359.4]
  assign _T_99430 = _T_99429[13:0]; // @[Modules.scala 160:64:@47360.4]
  assign buffer_14_350 = $signed(_T_99430); // @[Modules.scala 160:64:@47361.4]
  assign buffer_14_98 = {{9{_T_97863[4]}},_T_97863}; // @[Modules.scala 112:22:@8.4]
  assign _T_99432 = $signed(buffer_14_98) + $signed(buffer_4_106); // @[Modules.scala 160:64:@47363.4]
  assign _T_99433 = _T_99432[13:0]; // @[Modules.scala 160:64:@47364.4]
  assign buffer_14_351 = $signed(_T_99433); // @[Modules.scala 160:64:@47365.4]
  assign buffer_14_101 = {{9{_T_97884[4]}},_T_97884}; // @[Modules.scala 112:22:@8.4]
  assign _T_99435 = $signed(buffer_3_113) + $signed(buffer_14_101); // @[Modules.scala 160:64:@47367.4]
  assign _T_99436 = _T_99435[13:0]; // @[Modules.scala 160:64:@47368.4]
  assign buffer_14_352 = $signed(_T_99436); // @[Modules.scala 160:64:@47369.4]
  assign _T_99438 = $signed(buffer_5_115) + $signed(buffer_5_116); // @[Modules.scala 160:64:@47371.4]
  assign _T_99439 = _T_99438[13:0]; // @[Modules.scala 160:64:@47372.4]
  assign buffer_14_353 = $signed(_T_99439); // @[Modules.scala 160:64:@47373.4]
  assign buffer_14_105 = {{9{_T_97912[4]}},_T_97912}; // @[Modules.scala 112:22:@8.4]
  assign _T_99441 = $signed(buffer_5_117) + $signed(buffer_14_105); // @[Modules.scala 160:64:@47375.4]
  assign _T_99442 = _T_99441[13:0]; // @[Modules.scala 160:64:@47376.4]
  assign buffer_14_354 = $signed(_T_99442); // @[Modules.scala 160:64:@47377.4]
  assign _T_99444 = $signed(buffer_2_117) + $signed(buffer_2_118); // @[Modules.scala 160:64:@47379.4]
  assign _T_99445 = _T_99444[13:0]; // @[Modules.scala 160:64:@47380.4]
  assign buffer_14_355 = $signed(_T_99445); // @[Modules.scala 160:64:@47381.4]
  assign buffer_14_108 = {{8{_T_97933[5]}},_T_97933}; // @[Modules.scala 112:22:@8.4]
  assign _T_99447 = $signed(buffer_14_108) + $signed(buffer_1_118); // @[Modules.scala 160:64:@47383.4]
  assign _T_99448 = _T_99447[13:0]; // @[Modules.scala 160:64:@47384.4]
  assign buffer_14_356 = $signed(_T_99448); // @[Modules.scala 160:64:@47385.4]
  assign _T_99450 = $signed(buffer_1_119) + $signed(buffer_1_120); // @[Modules.scala 160:64:@47387.4]
  assign _T_99451 = _T_99450[13:0]; // @[Modules.scala 160:64:@47388.4]
  assign buffer_14_357 = $signed(_T_99451); // @[Modules.scala 160:64:@47389.4]
  assign buffer_14_112 = {{8{_T_97961[5]}},_T_97961}; // @[Modules.scala 112:22:@8.4]
  assign _T_99453 = $signed(buffer_14_112) + $signed(buffer_9_127); // @[Modules.scala 160:64:@47391.4]
  assign _T_99454 = _T_99453[13:0]; // @[Modules.scala 160:64:@47392.4]
  assign buffer_14_358 = $signed(_T_99454); // @[Modules.scala 160:64:@47393.4]
  assign _T_99456 = $signed(buffer_9_128) + $signed(buffer_11_118); // @[Modules.scala 160:64:@47395.4]
  assign _T_99457 = _T_99456[13:0]; // @[Modules.scala 160:64:@47396.4]
  assign buffer_14_359 = $signed(_T_99457); // @[Modules.scala 160:64:@47397.4]
  assign buffer_14_116 = {{8{_T_97989[5]}},_T_97989}; // @[Modules.scala 112:22:@8.4]
  assign _T_99459 = $signed(buffer_14_116) + $signed(buffer_7_126); // @[Modules.scala 160:64:@47399.4]
  assign _T_99460 = _T_99459[13:0]; // @[Modules.scala 160:64:@47400.4]
  assign buffer_14_360 = $signed(_T_99460); // @[Modules.scala 160:64:@47401.4]
  assign _T_99462 = $signed(buffer_4_124) + $signed(buffer_9_134); // @[Modules.scala 160:64:@47403.4]
  assign _T_99463 = _T_99462[13:0]; // @[Modules.scala 160:64:@47404.4]
  assign buffer_14_361 = $signed(_T_99463); // @[Modules.scala 160:64:@47405.4]
  assign buffer_14_120 = {{8{_T_98017[5]}},_T_98017}; // @[Modules.scala 112:22:@8.4]
  assign _T_99465 = $signed(buffer_14_120) + $signed(buffer_12_118); // @[Modules.scala 160:64:@47407.4]
  assign _T_99466 = _T_99465[13:0]; // @[Modules.scala 160:64:@47408.4]
  assign buffer_14_362 = $signed(_T_99466); // @[Modules.scala 160:64:@47409.4]
  assign _T_99468 = $signed(buffer_5_133) + $signed(buffer_1_133); // @[Modules.scala 160:64:@47411.4]
  assign _T_99469 = _T_99468[13:0]; // @[Modules.scala 160:64:@47412.4]
  assign buffer_14_363 = $signed(_T_99469); // @[Modules.scala 160:64:@47413.4]
  assign _T_99471 = $signed(buffer_5_135) + $signed(buffer_13_133); // @[Modules.scala 160:64:@47415.4]
  assign _T_99472 = _T_99471[13:0]; // @[Modules.scala 160:64:@47416.4]
  assign buffer_14_364 = $signed(_T_99472); // @[Modules.scala 160:64:@47417.4]
  assign buffer_14_126 = {{9{_T_98059[4]}},_T_98059}; // @[Modules.scala 112:22:@8.4]
  assign _T_99474 = $signed(buffer_14_126) + $signed(buffer_10_137); // @[Modules.scala 160:64:@47419.4]
  assign _T_99475 = _T_99474[13:0]; // @[Modules.scala 160:64:@47420.4]
  assign buffer_14_365 = $signed(_T_99475); // @[Modules.scala 160:64:@47421.4]
  assign buffer_14_130 = {{9{_T_98087[4]}},_T_98087}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_131 = {{8{_T_98094[5]}},_T_98094}; // @[Modules.scala 112:22:@8.4]
  assign _T_99480 = $signed(buffer_14_130) + $signed(buffer_14_131); // @[Modules.scala 160:64:@47427.4]
  assign _T_99481 = _T_99480[13:0]; // @[Modules.scala 160:64:@47428.4]
  assign buffer_14_367 = $signed(_T_99481); // @[Modules.scala 160:64:@47429.4]
  assign buffer_14_132 = {{8{_T_98101[5]}},_T_98101}; // @[Modules.scala 112:22:@8.4]
  assign _T_99483 = $signed(buffer_14_132) + $signed(buffer_1_145); // @[Modules.scala 160:64:@47431.4]
  assign _T_99484 = _T_99483[13:0]; // @[Modules.scala 160:64:@47432.4]
  assign buffer_14_368 = $signed(_T_99484); // @[Modules.scala 160:64:@47433.4]
  assign _T_99486 = $signed(buffer_7_145) + $signed(buffer_7_146); // @[Modules.scala 160:64:@47435.4]
  assign _T_99487 = _T_99486[13:0]; // @[Modules.scala 160:64:@47436.4]
  assign buffer_14_369 = $signed(_T_99487); // @[Modules.scala 160:64:@47437.4]
  assign buffer_14_136 = {{9{_T_98129[4]}},_T_98129}; // @[Modules.scala 112:22:@8.4]
  assign _T_99489 = $signed(buffer_14_136) + $signed(buffer_2_152); // @[Modules.scala 160:64:@47439.4]
  assign _T_99490 = _T_99489[13:0]; // @[Modules.scala 160:64:@47440.4]
  assign buffer_14_370 = $signed(_T_99490); // @[Modules.scala 160:64:@47441.4]
  assign _T_99492 = $signed(buffer_2_153) + $signed(buffer_2_154); // @[Modules.scala 160:64:@47443.4]
  assign _T_99493 = _T_99492[13:0]; // @[Modules.scala 160:64:@47444.4]
  assign buffer_14_371 = $signed(_T_99493); // @[Modules.scala 160:64:@47445.4]
  assign buffer_14_140 = {{8{_T_98157[5]}},_T_98157}; // @[Modules.scala 112:22:@8.4]
  assign _T_99495 = $signed(buffer_14_140) + $signed(buffer_0_152); // @[Modules.scala 160:64:@47447.4]
  assign _T_99496 = _T_99495[13:0]; // @[Modules.scala 160:64:@47448.4]
  assign buffer_14_372 = $signed(_T_99496); // @[Modules.scala 160:64:@47449.4]
  assign buffer_14_142 = {{8{_T_98171[5]}},_T_98171}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_143 = {{8{_T_98178[5]}},_T_98178}; // @[Modules.scala 112:22:@8.4]
  assign _T_99498 = $signed(buffer_14_142) + $signed(buffer_14_143); // @[Modules.scala 160:64:@47451.4]
  assign _T_99499 = _T_99498[13:0]; // @[Modules.scala 160:64:@47452.4]
  assign buffer_14_373 = $signed(_T_99499); // @[Modules.scala 160:64:@47453.4]
  assign buffer_14_144 = {{8{_T_98185[5]}},_T_98185}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_145 = {{8{_T_98192[5]}},_T_98192}; // @[Modules.scala 112:22:@8.4]
  assign _T_99501 = $signed(buffer_14_144) + $signed(buffer_14_145); // @[Modules.scala 160:64:@47455.4]
  assign _T_99502 = _T_99501[13:0]; // @[Modules.scala 160:64:@47456.4]
  assign buffer_14_374 = $signed(_T_99502); // @[Modules.scala 160:64:@47457.4]
  assign buffer_14_148 = {{9{_T_98213[4]}},_T_98213}; // @[Modules.scala 112:22:@8.4]
  assign _T_99507 = $signed(buffer_14_148) + $signed(buffer_2_165); // @[Modules.scala 160:64:@47463.4]
  assign _T_99508 = _T_99507[13:0]; // @[Modules.scala 160:64:@47464.4]
  assign buffer_14_376 = $signed(_T_99508); // @[Modules.scala 160:64:@47465.4]
  assign _T_99510 = $signed(buffer_1_162) + $signed(buffer_12_150); // @[Modules.scala 160:64:@47467.4]
  assign _T_99511 = _T_99510[13:0]; // @[Modules.scala 160:64:@47468.4]
  assign buffer_14_377 = $signed(_T_99511); // @[Modules.scala 160:64:@47469.4]
  assign buffer_14_152 = {{8{_T_98241[5]}},_T_98241}; // @[Modules.scala 112:22:@8.4]
  assign _T_99513 = $signed(buffer_14_152) + $signed(buffer_7_165); // @[Modules.scala 160:64:@47471.4]
  assign _T_99514 = _T_99513[13:0]; // @[Modules.scala 160:64:@47472.4]
  assign buffer_14_378 = $signed(_T_99514); // @[Modules.scala 160:64:@47473.4]
  assign buffer_14_155 = {{8{_T_98262[5]}},_T_98262}; // @[Modules.scala 112:22:@8.4]
  assign _T_99516 = $signed(buffer_0_164) + $signed(buffer_14_155); // @[Modules.scala 160:64:@47475.4]
  assign _T_99517 = _T_99516[13:0]; // @[Modules.scala 160:64:@47476.4]
  assign buffer_14_379 = $signed(_T_99517); // @[Modules.scala 160:64:@47477.4]
  assign _T_99519 = $signed(buffer_8_165) + $signed(buffer_0_167); // @[Modules.scala 160:64:@47479.4]
  assign _T_99520 = _T_99519[13:0]; // @[Modules.scala 160:64:@47480.4]
  assign buffer_14_380 = $signed(_T_99520); // @[Modules.scala 160:64:@47481.4]
  assign buffer_14_161 = {{8{_T_98304[5]}},_T_98304}; // @[Modules.scala 112:22:@8.4]
  assign _T_99525 = $signed(buffer_3_176) + $signed(buffer_14_161); // @[Modules.scala 160:64:@47487.4]
  assign _T_99526 = _T_99525[13:0]; // @[Modules.scala 160:64:@47488.4]
  assign buffer_14_382 = $signed(_T_99526); // @[Modules.scala 160:64:@47489.4]
  assign buffer_14_162 = {{8{_T_98311[5]}},_T_98311}; // @[Modules.scala 112:22:@8.4]
  assign _T_99528 = $signed(buffer_14_162) + $signed(buffer_4_169); // @[Modules.scala 160:64:@47491.4]
  assign _T_99529 = _T_99528[13:0]; // @[Modules.scala 160:64:@47492.4]
  assign buffer_14_383 = $signed(_T_99529); // @[Modules.scala 160:64:@47493.4]
  assign _T_99531 = $signed(buffer_10_179) + $signed(buffer_0_176); // @[Modules.scala 160:64:@47495.4]
  assign _T_99532 = _T_99531[13:0]; // @[Modules.scala 160:64:@47496.4]
  assign buffer_14_384 = $signed(_T_99532); // @[Modules.scala 160:64:@47497.4]
  assign buffer_14_167 = {{8{_T_98346[5]}},_T_98346}; // @[Modules.scala 112:22:@8.4]
  assign _T_99534 = $signed(buffer_8_176) + $signed(buffer_14_167); // @[Modules.scala 160:64:@47499.4]
  assign _T_99535 = _T_99534[13:0]; // @[Modules.scala 160:64:@47500.4]
  assign buffer_14_385 = $signed(_T_99535); // @[Modules.scala 160:64:@47501.4]
  assign buffer_14_169 = {{8{_T_98360[5]}},_T_98360}; // @[Modules.scala 112:22:@8.4]
  assign _T_99537 = $signed(buffer_5_180) + $signed(buffer_14_169); // @[Modules.scala 160:64:@47503.4]
  assign _T_99538 = _T_99537[13:0]; // @[Modules.scala 160:64:@47504.4]
  assign buffer_14_386 = $signed(_T_99538); // @[Modules.scala 160:64:@47505.4]
  assign buffer_14_171 = {{9{_T_98374[4]}},_T_98374}; // @[Modules.scala 112:22:@8.4]
  assign _T_99540 = $signed(buffer_12_172) + $signed(buffer_14_171); // @[Modules.scala 160:64:@47507.4]
  assign _T_99541 = _T_99540[13:0]; // @[Modules.scala 160:64:@47508.4]
  assign buffer_14_387 = $signed(_T_99541); // @[Modules.scala 160:64:@47509.4]
  assign _T_99543 = $signed(buffer_1_182) + $signed(buffer_9_192); // @[Modules.scala 160:64:@47511.4]
  assign _T_99544 = _T_99543[13:0]; // @[Modules.scala 160:64:@47512.4]
  assign buffer_14_388 = $signed(_T_99544); // @[Modules.scala 160:64:@47513.4]
  assign buffer_14_174 = {{9{_T_98395[4]}},_T_98395}; // @[Modules.scala 112:22:@8.4]
  assign _T_99546 = $signed(buffer_14_174) + $signed(buffer_0_184); // @[Modules.scala 160:64:@47515.4]
  assign _T_99547 = _T_99546[13:0]; // @[Modules.scala 160:64:@47516.4]
  assign buffer_14_389 = $signed(_T_99547); // @[Modules.scala 160:64:@47517.4]
  assign buffer_14_176 = {{8{_T_98409[5]}},_T_98409}; // @[Modules.scala 112:22:@8.4]
  assign _T_99549 = $signed(buffer_14_176) + $signed(buffer_1_188); // @[Modules.scala 160:64:@47519.4]
  assign _T_99550 = _T_99549[13:0]; // @[Modules.scala 160:64:@47520.4]
  assign buffer_14_390 = $signed(_T_99550); // @[Modules.scala 160:64:@47521.4]
  assign buffer_14_178 = {{8{_T_98423[5]}},_T_98423}; // @[Modules.scala 112:22:@8.4]
  assign _T_99552 = $signed(buffer_14_178) + $signed(buffer_1_191); // @[Modules.scala 160:64:@47523.4]
  assign _T_99553 = _T_99552[13:0]; // @[Modules.scala 160:64:@47524.4]
  assign buffer_14_391 = $signed(_T_99553); // @[Modules.scala 160:64:@47525.4]
  assign buffer_14_181 = {{8{_T_98444[5]}},_T_98444}; // @[Modules.scala 112:22:@8.4]
  assign _T_99555 = $signed(buffer_0_190) + $signed(buffer_14_181); // @[Modules.scala 160:64:@47527.4]
  assign _T_99556 = _T_99555[13:0]; // @[Modules.scala 160:64:@47528.4]
  assign buffer_14_392 = $signed(_T_99556); // @[Modules.scala 160:64:@47529.4]
  assign buffer_14_182 = {{8{_T_98451[5]}},_T_98451}; // @[Modules.scala 112:22:@8.4]
  assign _T_99558 = $signed(buffer_14_182) + $signed(buffer_2_198); // @[Modules.scala 160:64:@47531.4]
  assign _T_99559 = _T_99558[13:0]; // @[Modules.scala 160:64:@47532.4]
  assign buffer_14_393 = $signed(_T_99559); // @[Modules.scala 160:64:@47533.4]
  assign _T_99561 = $signed(buffer_3_203) + $signed(buffer_0_194); // @[Modules.scala 160:64:@47535.4]
  assign _T_99562 = _T_99561[13:0]; // @[Modules.scala 160:64:@47536.4]
  assign buffer_14_394 = $signed(_T_99562); // @[Modules.scala 160:64:@47537.4]
  assign _T_99564 = $signed(buffer_5_198) + $signed(buffer_3_206); // @[Modules.scala 160:64:@47539.4]
  assign _T_99565 = _T_99564[13:0]; // @[Modules.scala 160:64:@47540.4]
  assign buffer_14_395 = $signed(_T_99565); // @[Modules.scala 160:64:@47541.4]
  assign buffer_14_188 = {{8{_T_98493[5]}},_T_98493}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_189 = {{8{_T_98500[5]}},_T_98500}; // @[Modules.scala 112:22:@8.4]
  assign _T_99567 = $signed(buffer_14_188) + $signed(buffer_14_189); // @[Modules.scala 160:64:@47543.4]
  assign _T_99568 = _T_99567[13:0]; // @[Modules.scala 160:64:@47544.4]
  assign buffer_14_396 = $signed(_T_99568); // @[Modules.scala 160:64:@47545.4]
  assign buffer_14_191 = {{8{_T_98514[5]}},_T_98514}; // @[Modules.scala 112:22:@8.4]
  assign _T_99570 = $signed(buffer_8_205) + $signed(buffer_14_191); // @[Modules.scala 160:64:@47547.4]
  assign _T_99571 = _T_99570[13:0]; // @[Modules.scala 160:64:@47548.4]
  assign buffer_14_397 = $signed(_T_99571); // @[Modules.scala 160:64:@47549.4]
  assign _T_99573 = $signed(buffer_0_203) + $signed(buffer_5_207); // @[Modules.scala 160:64:@47551.4]
  assign _T_99574 = _T_99573[13:0]; // @[Modules.scala 160:64:@47552.4]
  assign buffer_14_398 = $signed(_T_99574); // @[Modules.scala 160:64:@47553.4]
  assign buffer_14_194 = {{8{_T_98535[5]}},_T_98535}; // @[Modules.scala 112:22:@8.4]
  assign _T_99576 = $signed(buffer_14_194) + $signed(buffer_11_205); // @[Modules.scala 160:64:@47555.4]
  assign _T_99577 = _T_99576[13:0]; // @[Modules.scala 160:64:@47556.4]
  assign buffer_14_399 = $signed(_T_99577); // @[Modules.scala 160:64:@47557.4]
  assign buffer_14_196 = {{8{_T_98549[5]}},_T_98549}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_197 = {{8{_T_98556[5]}},_T_98556}; // @[Modules.scala 112:22:@8.4]
  assign _T_99579 = $signed(buffer_14_196) + $signed(buffer_14_197); // @[Modules.scala 160:64:@47559.4]
  assign _T_99580 = _T_99579[13:0]; // @[Modules.scala 160:64:@47560.4]
  assign buffer_14_400 = $signed(_T_99580); // @[Modules.scala 160:64:@47561.4]
  assign buffer_14_199 = {{8{_T_98570[5]}},_T_98570}; // @[Modules.scala 112:22:@8.4]
  assign _T_99582 = $signed(buffer_11_207) + $signed(buffer_14_199); // @[Modules.scala 160:64:@47563.4]
  assign _T_99583 = _T_99582[13:0]; // @[Modules.scala 160:64:@47564.4]
  assign buffer_14_401 = $signed(_T_99583); // @[Modules.scala 160:64:@47565.4]
  assign _T_99585 = $signed(buffer_13_211) + $signed(buffer_13_212); // @[Modules.scala 160:64:@47567.4]
  assign _T_99586 = _T_99585[13:0]; // @[Modules.scala 160:64:@47568.4]
  assign buffer_14_402 = $signed(_T_99586); // @[Modules.scala 160:64:@47569.4]
  assign _T_99588 = $signed(buffer_6_223) + $signed(buffer_6_224); // @[Modules.scala 160:64:@47571.4]
  assign _T_99589 = _T_99588[13:0]; // @[Modules.scala 160:64:@47572.4]
  assign buffer_14_403 = $signed(_T_99589); // @[Modules.scala 160:64:@47573.4]
  assign buffer_14_205 = {{8{_T_98612[5]}},_T_98612}; // @[Modules.scala 112:22:@8.4]
  assign _T_99591 = $signed(buffer_6_225) + $signed(buffer_14_205); // @[Modules.scala 160:64:@47575.4]
  assign _T_99592 = _T_99591[13:0]; // @[Modules.scala 160:64:@47576.4]
  assign buffer_14_404 = $signed(_T_99592); // @[Modules.scala 160:64:@47577.4]
  assign _T_99594 = $signed(buffer_13_217) + $signed(buffer_1_217); // @[Modules.scala 160:64:@47579.4]
  assign _T_99595 = _T_99594[13:0]; // @[Modules.scala 160:64:@47580.4]
  assign buffer_14_405 = $signed(_T_99595); // @[Modules.scala 160:64:@47581.4]
  assign _T_99597 = $signed(buffer_6_229) + $signed(buffer_2_224); // @[Modules.scala 160:64:@47583.4]
  assign _T_99598 = _T_99597[13:0]; // @[Modules.scala 160:64:@47584.4]
  assign buffer_14_406 = $signed(_T_99598); // @[Modules.scala 160:64:@47585.4]
  assign _T_99612 = $signed(buffer_5_232) + $signed(buffer_8_234); // @[Modules.scala 160:64:@47603.4]
  assign _T_99613 = _T_99612[13:0]; // @[Modules.scala 160:64:@47604.4]
  assign buffer_14_411 = $signed(_T_99613); // @[Modules.scala 160:64:@47605.4]
  assign buffer_14_222 = {{9{_T_98731[4]}},_T_98731}; // @[Modules.scala 112:22:@8.4]
  assign _T_99618 = $signed(buffer_14_222) + $signed(buffer_5_238); // @[Modules.scala 160:64:@47611.4]
  assign _T_99619 = _T_99618[13:0]; // @[Modules.scala 160:64:@47612.4]
  assign buffer_14_413 = $signed(_T_99619); // @[Modules.scala 160:64:@47613.4]
  assign buffer_14_224 = {{8{_T_98745[5]}},_T_98745}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_225 = {{8{_T_98752[5]}},_T_98752}; // @[Modules.scala 112:22:@8.4]
  assign _T_99621 = $signed(buffer_14_224) + $signed(buffer_14_225); // @[Modules.scala 160:64:@47615.4]
  assign _T_99622 = _T_99621[13:0]; // @[Modules.scala 160:64:@47616.4]
  assign buffer_14_414 = $signed(_T_99622); // @[Modules.scala 160:64:@47617.4]
  assign buffer_14_226 = {{8{_T_98759[5]}},_T_98759}; // @[Modules.scala 112:22:@8.4]
  assign _T_99624 = $signed(buffer_14_226) + $signed(buffer_0_233); // @[Modules.scala 160:64:@47619.4]
  assign _T_99625 = _T_99624[13:0]; // @[Modules.scala 160:64:@47620.4]
  assign buffer_14_415 = $signed(_T_99625); // @[Modules.scala 160:64:@47621.4]
  assign buffer_14_229 = {{8{_T_98780[5]}},_T_98780}; // @[Modules.scala 112:22:@8.4]
  assign _T_99627 = $signed(buffer_9_245) + $signed(buffer_14_229); // @[Modules.scala 160:64:@47623.4]
  assign _T_99628 = _T_99627[13:0]; // @[Modules.scala 160:64:@47624.4]
  assign buffer_14_416 = $signed(_T_99628); // @[Modules.scala 160:64:@47625.4]
  assign buffer_14_231 = {{8{_T_98794[5]}},_T_98794}; // @[Modules.scala 112:22:@8.4]
  assign _T_99630 = $signed(buffer_6_247) + $signed(buffer_14_231); // @[Modules.scala 160:64:@47627.4]
  assign _T_99631 = _T_99630[13:0]; // @[Modules.scala 160:64:@47628.4]
  assign buffer_14_417 = $signed(_T_99631); // @[Modules.scala 160:64:@47629.4]
  assign buffer_14_232 = {{8{_T_98801[5]}},_T_98801}; // @[Modules.scala 112:22:@8.4]
  assign _T_99633 = $signed(buffer_14_232) + $signed(buffer_4_233); // @[Modules.scala 160:64:@47631.4]
  assign _T_99634 = _T_99633[13:0]; // @[Modules.scala 160:64:@47632.4]
  assign buffer_14_418 = $signed(_T_99634); // @[Modules.scala 160:64:@47633.4]
  assign buffer_14_234 = {{9{_T_98815[4]}},_T_98815}; // @[Modules.scala 112:22:@8.4]
  assign _T_99636 = $signed(buffer_14_234) + $signed(buffer_6_252); // @[Modules.scala 160:64:@47635.4]
  assign _T_99637 = _T_99636[13:0]; // @[Modules.scala 160:64:@47636.4]
  assign buffer_14_419 = $signed(_T_99637); // @[Modules.scala 160:64:@47637.4]
  assign buffer_14_237 = {{8{_T_98836[5]}},_T_98836}; // @[Modules.scala 112:22:@8.4]
  assign _T_99639 = $signed(buffer_11_241) + $signed(buffer_14_237); // @[Modules.scala 160:64:@47639.4]
  assign _T_99640 = _T_99639[13:0]; // @[Modules.scala 160:64:@47640.4]
  assign buffer_14_420 = $signed(_T_99640); // @[Modules.scala 160:64:@47641.4]
  assign buffer_14_239 = {{8{_T_98850[5]}},_T_98850}; // @[Modules.scala 112:22:@8.4]
  assign _T_99642 = $signed(buffer_12_239) + $signed(buffer_14_239); // @[Modules.scala 160:64:@47643.4]
  assign _T_99643 = _T_99642[13:0]; // @[Modules.scala 160:64:@47644.4]
  assign buffer_14_421 = $signed(_T_99643); // @[Modules.scala 160:64:@47645.4]
  assign buffer_14_240 = {{8{_T_98857[5]}},_T_98857}; // @[Modules.scala 112:22:@8.4]
  assign _T_99645 = $signed(buffer_14_240) + $signed(buffer_13_248); // @[Modules.scala 160:64:@47647.4]
  assign _T_99646 = _T_99645[13:0]; // @[Modules.scala 160:64:@47648.4]
  assign buffer_14_422 = $signed(_T_99646); // @[Modules.scala 160:64:@47649.4]
  assign buffer_14_243 = {{8{_T_98878[5]}},_T_98878}; // @[Modules.scala 112:22:@8.4]
  assign _T_99648 = $signed(buffer_0_246) + $signed(buffer_14_243); // @[Modules.scala 160:64:@47651.4]
  assign _T_99649 = _T_99648[13:0]; // @[Modules.scala 160:64:@47652.4]
  assign buffer_14_423 = $signed(_T_99649); // @[Modules.scala 160:64:@47653.4]
  assign buffer_14_245 = {{8{_T_98892[5]}},_T_98892}; // @[Modules.scala 112:22:@8.4]
  assign _T_99651 = $signed(buffer_9_259) + $signed(buffer_14_245); // @[Modules.scala 160:64:@47655.4]
  assign _T_99652 = _T_99651[13:0]; // @[Modules.scala 160:64:@47656.4]
  assign buffer_14_424 = $signed(_T_99652); // @[Modules.scala 160:64:@47657.4]
  assign _T_99657 = $signed(buffer_0_252) + $signed(buffer_13_256); // @[Modules.scala 160:64:@47663.4]
  assign _T_99658 = _T_99657[13:0]; // @[Modules.scala 160:64:@47664.4]
  assign buffer_14_426 = $signed(_T_99658); // @[Modules.scala 160:64:@47665.4]
  assign buffer_14_250 = {{8{_T_98927[5]}},_T_98927}; // @[Modules.scala 112:22:@8.4]
  assign _T_99660 = $signed(buffer_14_250) + $signed(buffer_13_257); // @[Modules.scala 160:64:@47667.4]
  assign _T_99661 = _T_99660[13:0]; // @[Modules.scala 160:64:@47668.4]
  assign buffer_14_427 = $signed(_T_99661); // @[Modules.scala 160:64:@47669.4]
  assign buffer_14_255 = {{8{_T_98962[5]}},_T_98962}; // @[Modules.scala 112:22:@8.4]
  assign _T_99666 = $signed(buffer_2_265) + $signed(buffer_14_255); // @[Modules.scala 160:64:@47675.4]
  assign _T_99667 = _T_99666[13:0]; // @[Modules.scala 160:64:@47676.4]
  assign buffer_14_429 = $signed(_T_99667); // @[Modules.scala 160:64:@47677.4]
  assign _T_99669 = $signed(buffer_12_255) + $signed(buffer_3_269); // @[Modules.scala 160:64:@47679.4]
  assign _T_99670 = _T_99669[13:0]; // @[Modules.scala 160:64:@47680.4]
  assign buffer_14_430 = $signed(_T_99670); // @[Modules.scala 160:64:@47681.4]
  assign buffer_14_259 = {{8{_T_98990[5]}},_T_98990}; // @[Modules.scala 112:22:@8.4]
  assign _T_99672 = $signed(buffer_6_272) + $signed(buffer_14_259); // @[Modules.scala 160:64:@47683.4]
  assign _T_99673 = _T_99672[13:0]; // @[Modules.scala 160:64:@47684.4]
  assign buffer_14_431 = $signed(_T_99673); // @[Modules.scala 160:64:@47685.4]
  assign _T_99678 = $signed(buffer_10_271) + $signed(buffer_13_270); // @[Modules.scala 160:64:@47691.4]
  assign _T_99679 = _T_99678[13:0]; // @[Modules.scala 160:64:@47692.4]
  assign buffer_14_433 = $signed(_T_99679); // @[Modules.scala 160:64:@47693.4]
  assign buffer_14_264 = {{8{_T_99025[5]}},_T_99025}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_265 = {{8{_T_99032[5]}},_T_99032}; // @[Modules.scala 112:22:@8.4]
  assign _T_99681 = $signed(buffer_14_264) + $signed(buffer_14_265); // @[Modules.scala 160:64:@47695.4]
  assign _T_99682 = _T_99681[13:0]; // @[Modules.scala 160:64:@47696.4]
  assign buffer_14_434 = $signed(_T_99682); // @[Modules.scala 160:64:@47697.4]
  assign buffer_14_267 = {{9{_T_99046[4]}},_T_99046}; // @[Modules.scala 112:22:@8.4]
  assign _T_99684 = $signed(buffer_0_270) + $signed(buffer_14_267); // @[Modules.scala 160:64:@47699.4]
  assign _T_99685 = _T_99684[13:0]; // @[Modules.scala 160:64:@47700.4]
  assign buffer_14_435 = $signed(_T_99685); // @[Modules.scala 160:64:@47701.4]
  assign _T_99687 = $signed(buffer_4_266) + $signed(buffer_0_273); // @[Modules.scala 160:64:@47703.4]
  assign _T_99688 = _T_99687[13:0]; // @[Modules.scala 160:64:@47704.4]
  assign buffer_14_436 = $signed(_T_99688); // @[Modules.scala 160:64:@47705.4]
  assign _T_99696 = $signed(buffer_3_287) + $signed(buffer_12_273); // @[Modules.scala 160:64:@47715.4]
  assign _T_99697 = _T_99696[13:0]; // @[Modules.scala 160:64:@47716.4]
  assign buffer_14_439 = $signed(_T_99697); // @[Modules.scala 160:64:@47717.4]
  assign buffer_14_276 = {{8{_T_99109[5]}},_T_99109}; // @[Modules.scala 112:22:@8.4]
  assign _T_99699 = $signed(buffer_14_276) + $signed(buffer_6_291); // @[Modules.scala 160:64:@47719.4]
  assign _T_99700 = _T_99699[13:0]; // @[Modules.scala 160:64:@47720.4]
  assign buffer_14_440 = $signed(_T_99700); // @[Modules.scala 160:64:@47721.4]
  assign buffer_14_279 = {{8{_T_99130[5]}},_T_99130}; // @[Modules.scala 112:22:@8.4]
  assign _T_99702 = $signed(buffer_6_292) + $signed(buffer_14_279); // @[Modules.scala 160:64:@47723.4]
  assign _T_99703 = _T_99702[13:0]; // @[Modules.scala 160:64:@47724.4]
  assign buffer_14_441 = $signed(_T_99703); // @[Modules.scala 160:64:@47725.4]
  assign _T_99705 = $signed(buffer_0_284) + $signed(buffer_1_283); // @[Modules.scala 160:64:@47727.4]
  assign _T_99706 = _T_99705[13:0]; // @[Modules.scala 160:64:@47728.4]
  assign buffer_14_442 = $signed(_T_99706); // @[Modules.scala 160:64:@47729.4]
  assign _T_99708 = $signed(buffer_7_291) + $signed(buffer_3_295); // @[Modules.scala 160:64:@47731.4]
  assign _T_99709 = _T_99708[13:0]; // @[Modules.scala 160:64:@47732.4]
  assign buffer_14_443 = $signed(_T_99709); // @[Modules.scala 160:64:@47733.4]
  assign _T_99717 = $signed(buffer_2_297) + $signed(buffer_2_298); // @[Modules.scala 160:64:@47743.4]
  assign _T_99718 = _T_99717[13:0]; // @[Modules.scala 160:64:@47744.4]
  assign buffer_14_446 = $signed(_T_99718); // @[Modules.scala 160:64:@47745.4]
  assign buffer_14_292 = {{8{_T_99221[5]}},_T_99221}; // @[Modules.scala 112:22:@8.4]
  assign _T_99723 = $signed(buffer_14_292) + $signed(buffer_5_305); // @[Modules.scala 160:64:@47751.4]
  assign _T_99724 = _T_99723[13:0]; // @[Modules.scala 160:64:@47752.4]
  assign buffer_14_448 = $signed(_T_99724); // @[Modules.scala 160:64:@47753.4]
  assign buffer_14_294 = {{8{_T_99235[5]}},_T_99235}; // @[Modules.scala 112:22:@8.4]
  assign buffer_14_295 = {{8{_T_99242[5]}},_T_99242}; // @[Modules.scala 112:22:@8.4]
  assign _T_99726 = $signed(buffer_14_294) + $signed(buffer_14_295); // @[Modules.scala 160:64:@47755.4]
  assign _T_99727 = _T_99726[13:0]; // @[Modules.scala 160:64:@47756.4]
  assign buffer_14_449 = $signed(_T_99727); // @[Modules.scala 160:64:@47757.4]
  assign buffer_14_296 = {{9{_T_99249[4]}},_T_99249}; // @[Modules.scala 112:22:@8.4]
  assign _T_99729 = $signed(buffer_14_296) + $signed(buffer_2_306); // @[Modules.scala 160:64:@47759.4]
  assign _T_99730 = _T_99729[13:0]; // @[Modules.scala 160:64:@47760.4]
  assign buffer_14_450 = $signed(_T_99730); // @[Modules.scala 160:64:@47761.4]
  assign buffer_14_300 = {{9{_T_99277[4]}},_T_99277}; // @[Modules.scala 112:22:@8.4]
  assign _T_99735 = $signed(buffer_14_300) + $signed(buffer_7_308); // @[Modules.scala 160:64:@47767.4]
  assign _T_99736 = _T_99735[13:0]; // @[Modules.scala 160:64:@47768.4]
  assign buffer_14_452 = $signed(_T_99736); // @[Modules.scala 160:64:@47769.4]
  assign _T_99738 = $signed(buffer_14_302) + $signed(buffer_14_303); // @[Modules.scala 166:64:@47771.4]
  assign _T_99739 = _T_99738[13:0]; // @[Modules.scala 166:64:@47772.4]
  assign buffer_14_453 = $signed(_T_99739); // @[Modules.scala 166:64:@47773.4]
  assign _T_99747 = $signed(buffer_14_308) + $signed(buffer_14_309); // @[Modules.scala 166:64:@47783.4]
  assign _T_99748 = _T_99747[13:0]; // @[Modules.scala 166:64:@47784.4]
  assign buffer_14_456 = $signed(_T_99748); // @[Modules.scala 166:64:@47785.4]
  assign _T_99750 = $signed(buffer_14_310) + $signed(buffer_14_311); // @[Modules.scala 166:64:@47787.4]
  assign _T_99751 = _T_99750[13:0]; // @[Modules.scala 166:64:@47788.4]
  assign buffer_14_457 = $signed(_T_99751); // @[Modules.scala 166:64:@47789.4]
  assign _T_99753 = $signed(buffer_2_319) + $signed(buffer_14_313); // @[Modules.scala 166:64:@47791.4]
  assign _T_99754 = _T_99753[13:0]; // @[Modules.scala 166:64:@47792.4]
  assign buffer_14_458 = $signed(_T_99754); // @[Modules.scala 166:64:@47793.4]
  assign _T_99756 = $signed(buffer_14_314) + $signed(buffer_14_315); // @[Modules.scala 166:64:@47795.4]
  assign _T_99757 = _T_99756[13:0]; // @[Modules.scala 166:64:@47796.4]
  assign buffer_14_459 = $signed(_T_99757); // @[Modules.scala 166:64:@47797.4]
  assign _T_99759 = $signed(buffer_14_316) + $signed(buffer_9_329); // @[Modules.scala 166:64:@47799.4]
  assign _T_99760 = _T_99759[13:0]; // @[Modules.scala 166:64:@47800.4]
  assign buffer_14_460 = $signed(_T_99760); // @[Modules.scala 166:64:@47801.4]
  assign _T_99762 = $signed(buffer_9_330) + $signed(buffer_14_319); // @[Modules.scala 166:64:@47803.4]
  assign _T_99763 = _T_99762[13:0]; // @[Modules.scala 166:64:@47804.4]
  assign buffer_14_461 = $signed(_T_99763); // @[Modules.scala 166:64:@47805.4]
  assign _T_99765 = $signed(buffer_14_320) + $signed(buffer_14_321); // @[Modules.scala 166:64:@47807.4]
  assign _T_99766 = _T_99765[13:0]; // @[Modules.scala 166:64:@47808.4]
  assign buffer_14_462 = $signed(_T_99766); // @[Modules.scala 166:64:@47809.4]
  assign _T_99768 = $signed(buffer_14_322) + $signed(buffer_14_323); // @[Modules.scala 166:64:@47811.4]
  assign _T_99769 = _T_99768[13:0]; // @[Modules.scala 166:64:@47812.4]
  assign buffer_14_463 = $signed(_T_99769); // @[Modules.scala 166:64:@47813.4]
  assign _T_99771 = $signed(buffer_14_324) + $signed(buffer_3_338); // @[Modules.scala 166:64:@47815.4]
  assign _T_99772 = _T_99771[13:0]; // @[Modules.scala 166:64:@47816.4]
  assign buffer_14_464 = $signed(_T_99772); // @[Modules.scala 166:64:@47817.4]
  assign _T_99774 = $signed(buffer_14_326) + $signed(buffer_13_333); // @[Modules.scala 166:64:@47819.4]
  assign _T_99775 = _T_99774[13:0]; // @[Modules.scala 166:64:@47820.4]
  assign buffer_14_465 = $signed(_T_99775); // @[Modules.scala 166:64:@47821.4]
  assign _T_99777 = $signed(buffer_6_342) + $signed(buffer_14_329); // @[Modules.scala 166:64:@47823.4]
  assign _T_99778 = _T_99777[13:0]; // @[Modules.scala 166:64:@47824.4]
  assign buffer_14_466 = $signed(_T_99778); // @[Modules.scala 166:64:@47825.4]
  assign _T_99780 = $signed(buffer_8_336) + $signed(buffer_14_331); // @[Modules.scala 166:64:@47827.4]
  assign _T_99781 = _T_99780[13:0]; // @[Modules.scala 166:64:@47828.4]
  assign buffer_14_467 = $signed(_T_99781); // @[Modules.scala 166:64:@47829.4]
  assign _T_99783 = $signed(buffer_14_332) + $signed(buffer_14_333); // @[Modules.scala 166:64:@47831.4]
  assign _T_99784 = _T_99783[13:0]; // @[Modules.scala 166:64:@47832.4]
  assign buffer_14_468 = $signed(_T_99784); // @[Modules.scala 166:64:@47833.4]
  assign _T_99786 = $signed(buffer_14_334) + $signed(buffer_14_335); // @[Modules.scala 166:64:@47835.4]
  assign _T_99787 = _T_99786[13:0]; // @[Modules.scala 166:64:@47836.4]
  assign buffer_14_469 = $signed(_T_99787); // @[Modules.scala 166:64:@47837.4]
  assign _T_99789 = $signed(buffer_14_336) + $signed(buffer_14_337); // @[Modules.scala 166:64:@47839.4]
  assign _T_99790 = _T_99789[13:0]; // @[Modules.scala 166:64:@47840.4]
  assign buffer_14_470 = $signed(_T_99790); // @[Modules.scala 166:64:@47841.4]
  assign _T_99792 = $signed(buffer_14_338) + $signed(buffer_14_339); // @[Modules.scala 166:64:@47843.4]
  assign _T_99793 = _T_99792[13:0]; // @[Modules.scala 166:64:@47844.4]
  assign buffer_14_471 = $signed(_T_99793); // @[Modules.scala 166:64:@47845.4]
  assign _T_99795 = $signed(buffer_14_340) + $signed(buffer_14_341); // @[Modules.scala 166:64:@47847.4]
  assign _T_99796 = _T_99795[13:0]; // @[Modules.scala 166:64:@47848.4]
  assign buffer_14_472 = $signed(_T_99796); // @[Modules.scala 166:64:@47849.4]
  assign _T_99798 = $signed(buffer_14_342) + $signed(buffer_3_359); // @[Modules.scala 166:64:@47851.4]
  assign _T_99799 = _T_99798[13:0]; // @[Modules.scala 166:64:@47852.4]
  assign buffer_14_473 = $signed(_T_99799); // @[Modules.scala 166:64:@47853.4]
  assign _T_99801 = $signed(buffer_14_344) + $signed(buffer_14_345); // @[Modules.scala 166:64:@47855.4]
  assign _T_99802 = _T_99801[13:0]; // @[Modules.scala 166:64:@47856.4]
  assign buffer_14_474 = $signed(_T_99802); // @[Modules.scala 166:64:@47857.4]
  assign _T_99804 = $signed(buffer_14_346) + $signed(buffer_10_355); // @[Modules.scala 166:64:@47859.4]
  assign _T_99805 = _T_99804[13:0]; // @[Modules.scala 166:64:@47860.4]
  assign buffer_14_475 = $signed(_T_99805); // @[Modules.scala 166:64:@47861.4]
  assign _T_99807 = $signed(buffer_14_348) + $signed(buffer_14_349); // @[Modules.scala 166:64:@47863.4]
  assign _T_99808 = _T_99807[13:0]; // @[Modules.scala 166:64:@47864.4]
  assign buffer_14_476 = $signed(_T_99808); // @[Modules.scala 166:64:@47865.4]
  assign _T_99810 = $signed(buffer_14_350) + $signed(buffer_14_351); // @[Modules.scala 166:64:@47867.4]
  assign _T_99811 = _T_99810[13:0]; // @[Modules.scala 166:64:@47868.4]
  assign buffer_14_477 = $signed(_T_99811); // @[Modules.scala 166:64:@47869.4]
  assign _T_99813 = $signed(buffer_14_352) + $signed(buffer_14_353); // @[Modules.scala 166:64:@47871.4]
  assign _T_99814 = _T_99813[13:0]; // @[Modules.scala 166:64:@47872.4]
  assign buffer_14_478 = $signed(_T_99814); // @[Modules.scala 166:64:@47873.4]
  assign _T_99816 = $signed(buffer_14_354) + $signed(buffer_14_355); // @[Modules.scala 166:64:@47875.4]
  assign _T_99817 = _T_99816[13:0]; // @[Modules.scala 166:64:@47876.4]
  assign buffer_14_479 = $signed(_T_99817); // @[Modules.scala 166:64:@47877.4]
  assign _T_99819 = $signed(buffer_14_356) + $signed(buffer_14_357); // @[Modules.scala 166:64:@47879.4]
  assign _T_99820 = _T_99819[13:0]; // @[Modules.scala 166:64:@47880.4]
  assign buffer_14_480 = $signed(_T_99820); // @[Modules.scala 166:64:@47881.4]
  assign _T_99822 = $signed(buffer_14_358) + $signed(buffer_14_359); // @[Modules.scala 166:64:@47883.4]
  assign _T_99823 = _T_99822[13:0]; // @[Modules.scala 166:64:@47884.4]
  assign buffer_14_481 = $signed(_T_99823); // @[Modules.scala 166:64:@47885.4]
  assign _T_99825 = $signed(buffer_14_360) + $signed(buffer_14_361); // @[Modules.scala 166:64:@47887.4]
  assign _T_99826 = _T_99825[13:0]; // @[Modules.scala 166:64:@47888.4]
  assign buffer_14_482 = $signed(_T_99826); // @[Modules.scala 166:64:@47889.4]
  assign _T_99828 = $signed(buffer_14_362) + $signed(buffer_14_363); // @[Modules.scala 166:64:@47891.4]
  assign _T_99829 = _T_99828[13:0]; // @[Modules.scala 166:64:@47892.4]
  assign buffer_14_483 = $signed(_T_99829); // @[Modules.scala 166:64:@47893.4]
  assign _T_99831 = $signed(buffer_14_364) + $signed(buffer_14_365); // @[Modules.scala 166:64:@47895.4]
  assign _T_99832 = _T_99831[13:0]; // @[Modules.scala 166:64:@47896.4]
  assign buffer_14_484 = $signed(_T_99832); // @[Modules.scala 166:64:@47897.4]
  assign _T_99834 = $signed(buffer_3_386) + $signed(buffer_14_367); // @[Modules.scala 166:64:@47899.4]
  assign _T_99835 = _T_99834[13:0]; // @[Modules.scala 166:64:@47900.4]
  assign buffer_14_485 = $signed(_T_99835); // @[Modules.scala 166:64:@47901.4]
  assign _T_99837 = $signed(buffer_14_368) + $signed(buffer_14_369); // @[Modules.scala 166:64:@47903.4]
  assign _T_99838 = _T_99837[13:0]; // @[Modules.scala 166:64:@47904.4]
  assign buffer_14_486 = $signed(_T_99838); // @[Modules.scala 166:64:@47905.4]
  assign _T_99840 = $signed(buffer_14_370) + $signed(buffer_14_371); // @[Modules.scala 166:64:@47907.4]
  assign _T_99841 = _T_99840[13:0]; // @[Modules.scala 166:64:@47908.4]
  assign buffer_14_487 = $signed(_T_99841); // @[Modules.scala 166:64:@47909.4]
  assign _T_99843 = $signed(buffer_14_372) + $signed(buffer_14_373); // @[Modules.scala 166:64:@47911.4]
  assign _T_99844 = _T_99843[13:0]; // @[Modules.scala 166:64:@47912.4]
  assign buffer_14_488 = $signed(_T_99844); // @[Modules.scala 166:64:@47913.4]
  assign _T_99846 = $signed(buffer_14_374) + $signed(buffer_7_388); // @[Modules.scala 166:64:@47915.4]
  assign _T_99847 = _T_99846[13:0]; // @[Modules.scala 166:64:@47916.4]
  assign buffer_14_489 = $signed(_T_99847); // @[Modules.scala 166:64:@47917.4]
  assign _T_99849 = $signed(buffer_14_376) + $signed(buffer_14_377); // @[Modules.scala 166:64:@47919.4]
  assign _T_99850 = _T_99849[13:0]; // @[Modules.scala 166:64:@47920.4]
  assign buffer_14_490 = $signed(_T_99850); // @[Modules.scala 166:64:@47921.4]
  assign _T_99852 = $signed(buffer_14_378) + $signed(buffer_14_379); // @[Modules.scala 166:64:@47923.4]
  assign _T_99853 = _T_99852[13:0]; // @[Modules.scala 166:64:@47924.4]
  assign buffer_14_491 = $signed(_T_99853); // @[Modules.scala 166:64:@47925.4]
  assign _T_99855 = $signed(buffer_14_380) + $signed(buffer_12_377); // @[Modules.scala 166:64:@47927.4]
  assign _T_99856 = _T_99855[13:0]; // @[Modules.scala 166:64:@47928.4]
  assign buffer_14_492 = $signed(_T_99856); // @[Modules.scala 166:64:@47929.4]
  assign _T_99858 = $signed(buffer_14_382) + $signed(buffer_14_383); // @[Modules.scala 166:64:@47931.4]
  assign _T_99859 = _T_99858[13:0]; // @[Modules.scala 166:64:@47932.4]
  assign buffer_14_493 = $signed(_T_99859); // @[Modules.scala 166:64:@47933.4]
  assign _T_99861 = $signed(buffer_14_384) + $signed(buffer_14_385); // @[Modules.scala 166:64:@47935.4]
  assign _T_99862 = _T_99861[13:0]; // @[Modules.scala 166:64:@47936.4]
  assign buffer_14_494 = $signed(_T_99862); // @[Modules.scala 166:64:@47937.4]
  assign _T_99864 = $signed(buffer_14_386) + $signed(buffer_14_387); // @[Modules.scala 166:64:@47939.4]
  assign _T_99865 = _T_99864[13:0]; // @[Modules.scala 166:64:@47940.4]
  assign buffer_14_495 = $signed(_T_99865); // @[Modules.scala 166:64:@47941.4]
  assign _T_99867 = $signed(buffer_14_388) + $signed(buffer_14_389); // @[Modules.scala 166:64:@47943.4]
  assign _T_99868 = _T_99867[13:0]; // @[Modules.scala 166:64:@47944.4]
  assign buffer_14_496 = $signed(_T_99868); // @[Modules.scala 166:64:@47945.4]
  assign _T_99870 = $signed(buffer_14_390) + $signed(buffer_14_391); // @[Modules.scala 166:64:@47947.4]
  assign _T_99871 = _T_99870[13:0]; // @[Modules.scala 166:64:@47948.4]
  assign buffer_14_497 = $signed(_T_99871); // @[Modules.scala 166:64:@47949.4]
  assign _T_99873 = $signed(buffer_14_392) + $signed(buffer_14_393); // @[Modules.scala 166:64:@47951.4]
  assign _T_99874 = _T_99873[13:0]; // @[Modules.scala 166:64:@47952.4]
  assign buffer_14_498 = $signed(_T_99874); // @[Modules.scala 166:64:@47953.4]
  assign _T_99876 = $signed(buffer_14_394) + $signed(buffer_14_395); // @[Modules.scala 166:64:@47955.4]
  assign _T_99877 = _T_99876[13:0]; // @[Modules.scala 166:64:@47956.4]
  assign buffer_14_499 = $signed(_T_99877); // @[Modules.scala 166:64:@47957.4]
  assign _T_99879 = $signed(buffer_14_396) + $signed(buffer_14_397); // @[Modules.scala 166:64:@47959.4]
  assign _T_99880 = _T_99879[13:0]; // @[Modules.scala 166:64:@47960.4]
  assign buffer_14_500 = $signed(_T_99880); // @[Modules.scala 166:64:@47961.4]
  assign _T_99882 = $signed(buffer_14_398) + $signed(buffer_14_399); // @[Modules.scala 166:64:@47963.4]
  assign _T_99883 = _T_99882[13:0]; // @[Modules.scala 166:64:@47964.4]
  assign buffer_14_501 = $signed(_T_99883); // @[Modules.scala 166:64:@47965.4]
  assign _T_99885 = $signed(buffer_14_400) + $signed(buffer_14_401); // @[Modules.scala 166:64:@47967.4]
  assign _T_99886 = _T_99885[13:0]; // @[Modules.scala 166:64:@47968.4]
  assign buffer_14_502 = $signed(_T_99886); // @[Modules.scala 166:64:@47969.4]
  assign _T_99888 = $signed(buffer_14_402) + $signed(buffer_14_403); // @[Modules.scala 166:64:@47971.4]
  assign _T_99889 = _T_99888[13:0]; // @[Modules.scala 166:64:@47972.4]
  assign buffer_14_503 = $signed(_T_99889); // @[Modules.scala 166:64:@47973.4]
  assign _T_99891 = $signed(buffer_14_404) + $signed(buffer_14_405); // @[Modules.scala 166:64:@47975.4]
  assign _T_99892 = _T_99891[13:0]; // @[Modules.scala 166:64:@47976.4]
  assign buffer_14_504 = $signed(_T_99892); // @[Modules.scala 166:64:@47977.4]
  assign _T_99894 = $signed(buffer_14_406) + $signed(buffer_10_421); // @[Modules.scala 166:64:@47979.4]
  assign _T_99895 = _T_99894[13:0]; // @[Modules.scala 166:64:@47980.4]
  assign buffer_14_505 = $signed(_T_99895); // @[Modules.scala 166:64:@47981.4]
  assign _T_99897 = $signed(buffer_7_425) + $signed(buffer_13_419); // @[Modules.scala 166:64:@47983.4]
  assign _T_99898 = _T_99897[13:0]; // @[Modules.scala 166:64:@47984.4]
  assign buffer_14_506 = $signed(_T_99898); // @[Modules.scala 166:64:@47985.4]
  assign _T_99900 = $signed(buffer_5_429) + $signed(buffer_14_411); // @[Modules.scala 166:64:@47987.4]
  assign _T_99901 = _T_99900[13:0]; // @[Modules.scala 166:64:@47988.4]
  assign buffer_14_507 = $signed(_T_99901); // @[Modules.scala 166:64:@47989.4]
  assign _T_99903 = $signed(buffer_13_422) + $signed(buffer_14_413); // @[Modules.scala 166:64:@47991.4]
  assign _T_99904 = _T_99903[13:0]; // @[Modules.scala 166:64:@47992.4]
  assign buffer_14_508 = $signed(_T_99904); // @[Modules.scala 166:64:@47993.4]
  assign _T_99906 = $signed(buffer_14_414) + $signed(buffer_14_415); // @[Modules.scala 166:64:@47995.4]
  assign _T_99907 = _T_99906[13:0]; // @[Modules.scala 166:64:@47996.4]
  assign buffer_14_509 = $signed(_T_99907); // @[Modules.scala 166:64:@47997.4]
  assign _T_99909 = $signed(buffer_14_416) + $signed(buffer_14_417); // @[Modules.scala 166:64:@47999.4]
  assign _T_99910 = _T_99909[13:0]; // @[Modules.scala 166:64:@48000.4]
  assign buffer_14_510 = $signed(_T_99910); // @[Modules.scala 166:64:@48001.4]
  assign _T_99912 = $signed(buffer_14_418) + $signed(buffer_14_419); // @[Modules.scala 166:64:@48003.4]
  assign _T_99913 = _T_99912[13:0]; // @[Modules.scala 166:64:@48004.4]
  assign buffer_14_511 = $signed(_T_99913); // @[Modules.scala 166:64:@48005.4]
  assign _T_99915 = $signed(buffer_14_420) + $signed(buffer_14_421); // @[Modules.scala 166:64:@48007.4]
  assign _T_99916 = _T_99915[13:0]; // @[Modules.scala 166:64:@48008.4]
  assign buffer_14_512 = $signed(_T_99916); // @[Modules.scala 166:64:@48009.4]
  assign _T_99918 = $signed(buffer_14_422) + $signed(buffer_14_423); // @[Modules.scala 166:64:@48011.4]
  assign _T_99919 = _T_99918[13:0]; // @[Modules.scala 166:64:@48012.4]
  assign buffer_14_513 = $signed(_T_99919); // @[Modules.scala 166:64:@48013.4]
  assign _T_99921 = $signed(buffer_14_424) + $signed(buffer_0_427); // @[Modules.scala 166:64:@48015.4]
  assign _T_99922 = _T_99921[13:0]; // @[Modules.scala 166:64:@48016.4]
  assign buffer_14_514 = $signed(_T_99922); // @[Modules.scala 166:64:@48017.4]
  assign _T_99924 = $signed(buffer_14_426) + $signed(buffer_14_427); // @[Modules.scala 166:64:@48019.4]
  assign _T_99925 = _T_99924[13:0]; // @[Modules.scala 166:64:@48020.4]
  assign buffer_14_515 = $signed(_T_99925); // @[Modules.scala 166:64:@48021.4]
  assign _T_99927 = $signed(buffer_3_446) + $signed(buffer_14_429); // @[Modules.scala 166:64:@48023.4]
  assign _T_99928 = _T_99927[13:0]; // @[Modules.scala 166:64:@48024.4]
  assign buffer_14_516 = $signed(_T_99928); // @[Modules.scala 166:64:@48025.4]
  assign _T_99930 = $signed(buffer_14_430) + $signed(buffer_14_431); // @[Modules.scala 166:64:@48027.4]
  assign _T_99931 = _T_99930[13:0]; // @[Modules.scala 166:64:@48028.4]
  assign buffer_14_517 = $signed(_T_99931); // @[Modules.scala 166:64:@48029.4]
  assign _T_99933 = $signed(buffer_12_428) + $signed(buffer_14_433); // @[Modules.scala 166:64:@48031.4]
  assign _T_99934 = _T_99933[13:0]; // @[Modules.scala 166:64:@48032.4]
  assign buffer_14_518 = $signed(_T_99934); // @[Modules.scala 166:64:@48033.4]
  assign _T_99936 = $signed(buffer_14_434) + $signed(buffer_14_435); // @[Modules.scala 166:64:@48035.4]
  assign _T_99937 = _T_99936[13:0]; // @[Modules.scala 166:64:@48036.4]
  assign buffer_14_519 = $signed(_T_99937); // @[Modules.scala 166:64:@48037.4]
  assign _T_99939 = $signed(buffer_14_436) + $signed(buffer_10_447); // @[Modules.scala 166:64:@48039.4]
  assign _T_99940 = _T_99939[13:0]; // @[Modules.scala 166:64:@48040.4]
  assign buffer_14_520 = $signed(_T_99940); // @[Modules.scala 166:64:@48041.4]
  assign _T_99942 = $signed(buffer_10_448) + $signed(buffer_14_439); // @[Modules.scala 166:64:@48043.4]
  assign _T_99943 = _T_99942[13:0]; // @[Modules.scala 166:64:@48044.4]
  assign buffer_14_521 = $signed(_T_99943); // @[Modules.scala 166:64:@48045.4]
  assign _T_99945 = $signed(buffer_14_440) + $signed(buffer_14_441); // @[Modules.scala 166:64:@48047.4]
  assign _T_99946 = _T_99945[13:0]; // @[Modules.scala 166:64:@48048.4]
  assign buffer_14_522 = $signed(_T_99946); // @[Modules.scala 166:64:@48049.4]
  assign _T_99948 = $signed(buffer_14_442) + $signed(buffer_14_443); // @[Modules.scala 166:64:@48051.4]
  assign _T_99949 = _T_99948[13:0]; // @[Modules.scala 166:64:@48052.4]
  assign buffer_14_523 = $signed(_T_99949); // @[Modules.scala 166:64:@48053.4]
  assign _T_99954 = $signed(buffer_14_446) + $signed(buffer_5_465); // @[Modules.scala 166:64:@48059.4]
  assign _T_99955 = _T_99954[13:0]; // @[Modules.scala 166:64:@48060.4]
  assign buffer_14_525 = $signed(_T_99955); // @[Modules.scala 166:64:@48061.4]
  assign _T_99957 = $signed(buffer_14_448) + $signed(buffer_14_449); // @[Modules.scala 166:64:@48063.4]
  assign _T_99958 = _T_99957[13:0]; // @[Modules.scala 166:64:@48064.4]
  assign buffer_14_526 = $signed(_T_99958); // @[Modules.scala 166:64:@48065.4]
  assign _T_99960 = $signed(buffer_14_450) + $signed(buffer_3_469); // @[Modules.scala 166:64:@48067.4]
  assign _T_99961 = _T_99960[13:0]; // @[Modules.scala 166:64:@48068.4]
  assign buffer_14_527 = $signed(_T_99961); // @[Modules.scala 166:64:@48069.4]
  assign _T_99963 = $signed(buffer_14_453) + $signed(buffer_0_454); // @[Modules.scala 166:64:@48071.4]
  assign _T_99964 = _T_99963[13:0]; // @[Modules.scala 166:64:@48072.4]
  assign buffer_14_528 = $signed(_T_99964); // @[Modules.scala 166:64:@48073.4]
  assign _T_99966 = $signed(buffer_0_455) + $signed(buffer_14_456); // @[Modules.scala 166:64:@48075.4]
  assign _T_99967 = _T_99966[13:0]; // @[Modules.scala 166:64:@48076.4]
  assign buffer_14_529 = $signed(_T_99967); // @[Modules.scala 166:64:@48077.4]
  assign _T_99969 = $signed(buffer_14_457) + $signed(buffer_14_458); // @[Modules.scala 166:64:@48079.4]
  assign _T_99970 = _T_99969[13:0]; // @[Modules.scala 166:64:@48080.4]
  assign buffer_14_530 = $signed(_T_99970); // @[Modules.scala 166:64:@48081.4]
  assign _T_99972 = $signed(buffer_14_459) + $signed(buffer_14_460); // @[Modules.scala 166:64:@48083.4]
  assign _T_99973 = _T_99972[13:0]; // @[Modules.scala 166:64:@48084.4]
  assign buffer_14_531 = $signed(_T_99973); // @[Modules.scala 166:64:@48085.4]
  assign _T_99975 = $signed(buffer_14_461) + $signed(buffer_14_462); // @[Modules.scala 166:64:@48087.4]
  assign _T_99976 = _T_99975[13:0]; // @[Modules.scala 166:64:@48088.4]
  assign buffer_14_532 = $signed(_T_99976); // @[Modules.scala 166:64:@48089.4]
  assign _T_99978 = $signed(buffer_14_463) + $signed(buffer_14_464); // @[Modules.scala 166:64:@48091.4]
  assign _T_99979 = _T_99978[13:0]; // @[Modules.scala 166:64:@48092.4]
  assign buffer_14_533 = $signed(_T_99979); // @[Modules.scala 166:64:@48093.4]
  assign _T_99981 = $signed(buffer_14_465) + $signed(buffer_14_466); // @[Modules.scala 166:64:@48095.4]
  assign _T_99982 = _T_99981[13:0]; // @[Modules.scala 166:64:@48096.4]
  assign buffer_14_534 = $signed(_T_99982); // @[Modules.scala 166:64:@48097.4]
  assign _T_99984 = $signed(buffer_14_467) + $signed(buffer_14_468); // @[Modules.scala 166:64:@48099.4]
  assign _T_99985 = _T_99984[13:0]; // @[Modules.scala 166:64:@48100.4]
  assign buffer_14_535 = $signed(_T_99985); // @[Modules.scala 166:64:@48101.4]
  assign _T_99987 = $signed(buffer_14_469) + $signed(buffer_14_470); // @[Modules.scala 166:64:@48103.4]
  assign _T_99988 = _T_99987[13:0]; // @[Modules.scala 166:64:@48104.4]
  assign buffer_14_536 = $signed(_T_99988); // @[Modules.scala 166:64:@48105.4]
  assign _T_99990 = $signed(buffer_14_471) + $signed(buffer_14_472); // @[Modules.scala 166:64:@48107.4]
  assign _T_99991 = _T_99990[13:0]; // @[Modules.scala 166:64:@48108.4]
  assign buffer_14_537 = $signed(_T_99991); // @[Modules.scala 166:64:@48109.4]
  assign _T_99993 = $signed(buffer_14_473) + $signed(buffer_14_474); // @[Modules.scala 166:64:@48111.4]
  assign _T_99994 = _T_99993[13:0]; // @[Modules.scala 166:64:@48112.4]
  assign buffer_14_538 = $signed(_T_99994); // @[Modules.scala 166:64:@48113.4]
  assign _T_99996 = $signed(buffer_14_475) + $signed(buffer_14_476); // @[Modules.scala 166:64:@48115.4]
  assign _T_99997 = _T_99996[13:0]; // @[Modules.scala 166:64:@48116.4]
  assign buffer_14_539 = $signed(_T_99997); // @[Modules.scala 166:64:@48117.4]
  assign _T_99999 = $signed(buffer_14_477) + $signed(buffer_14_478); // @[Modules.scala 166:64:@48119.4]
  assign _T_100000 = _T_99999[13:0]; // @[Modules.scala 166:64:@48120.4]
  assign buffer_14_540 = $signed(_T_100000); // @[Modules.scala 166:64:@48121.4]
  assign _T_100002 = $signed(buffer_14_479) + $signed(buffer_14_480); // @[Modules.scala 166:64:@48123.4]
  assign _T_100003 = _T_100002[13:0]; // @[Modules.scala 166:64:@48124.4]
  assign buffer_14_541 = $signed(_T_100003); // @[Modules.scala 166:64:@48125.4]
  assign _T_100005 = $signed(buffer_14_481) + $signed(buffer_14_482); // @[Modules.scala 166:64:@48127.4]
  assign _T_100006 = _T_100005[13:0]; // @[Modules.scala 166:64:@48128.4]
  assign buffer_14_542 = $signed(_T_100006); // @[Modules.scala 166:64:@48129.4]
  assign _T_100008 = $signed(buffer_14_483) + $signed(buffer_14_484); // @[Modules.scala 166:64:@48131.4]
  assign _T_100009 = _T_100008[13:0]; // @[Modules.scala 166:64:@48132.4]
  assign buffer_14_543 = $signed(_T_100009); // @[Modules.scala 166:64:@48133.4]
  assign _T_100011 = $signed(buffer_14_485) + $signed(buffer_14_486); // @[Modules.scala 166:64:@48135.4]
  assign _T_100012 = _T_100011[13:0]; // @[Modules.scala 166:64:@48136.4]
  assign buffer_14_544 = $signed(_T_100012); // @[Modules.scala 166:64:@48137.4]
  assign _T_100014 = $signed(buffer_14_487) + $signed(buffer_14_488); // @[Modules.scala 166:64:@48139.4]
  assign _T_100015 = _T_100014[13:0]; // @[Modules.scala 166:64:@48140.4]
  assign buffer_14_545 = $signed(_T_100015); // @[Modules.scala 166:64:@48141.4]
  assign _T_100017 = $signed(buffer_14_489) + $signed(buffer_14_490); // @[Modules.scala 166:64:@48143.4]
  assign _T_100018 = _T_100017[13:0]; // @[Modules.scala 166:64:@48144.4]
  assign buffer_14_546 = $signed(_T_100018); // @[Modules.scala 166:64:@48145.4]
  assign _T_100020 = $signed(buffer_14_491) + $signed(buffer_14_492); // @[Modules.scala 166:64:@48147.4]
  assign _T_100021 = _T_100020[13:0]; // @[Modules.scala 166:64:@48148.4]
  assign buffer_14_547 = $signed(_T_100021); // @[Modules.scala 166:64:@48149.4]
  assign _T_100023 = $signed(buffer_14_493) + $signed(buffer_14_494); // @[Modules.scala 166:64:@48151.4]
  assign _T_100024 = _T_100023[13:0]; // @[Modules.scala 166:64:@48152.4]
  assign buffer_14_548 = $signed(_T_100024); // @[Modules.scala 166:64:@48153.4]
  assign _T_100026 = $signed(buffer_14_495) + $signed(buffer_14_496); // @[Modules.scala 166:64:@48155.4]
  assign _T_100027 = _T_100026[13:0]; // @[Modules.scala 166:64:@48156.4]
  assign buffer_14_549 = $signed(_T_100027); // @[Modules.scala 166:64:@48157.4]
  assign _T_100029 = $signed(buffer_14_497) + $signed(buffer_14_498); // @[Modules.scala 166:64:@48159.4]
  assign _T_100030 = _T_100029[13:0]; // @[Modules.scala 166:64:@48160.4]
  assign buffer_14_550 = $signed(_T_100030); // @[Modules.scala 166:64:@48161.4]
  assign _T_100032 = $signed(buffer_14_499) + $signed(buffer_14_500); // @[Modules.scala 166:64:@48163.4]
  assign _T_100033 = _T_100032[13:0]; // @[Modules.scala 166:64:@48164.4]
  assign buffer_14_551 = $signed(_T_100033); // @[Modules.scala 166:64:@48165.4]
  assign _T_100035 = $signed(buffer_14_501) + $signed(buffer_14_502); // @[Modules.scala 166:64:@48167.4]
  assign _T_100036 = _T_100035[13:0]; // @[Modules.scala 166:64:@48168.4]
  assign buffer_14_552 = $signed(_T_100036); // @[Modules.scala 166:64:@48169.4]
  assign _T_100038 = $signed(buffer_14_503) + $signed(buffer_14_504); // @[Modules.scala 166:64:@48171.4]
  assign _T_100039 = _T_100038[13:0]; // @[Modules.scala 166:64:@48172.4]
  assign buffer_14_553 = $signed(_T_100039); // @[Modules.scala 166:64:@48173.4]
  assign _T_100041 = $signed(buffer_14_505) + $signed(buffer_14_506); // @[Modules.scala 166:64:@48175.4]
  assign _T_100042 = _T_100041[13:0]; // @[Modules.scala 166:64:@48176.4]
  assign buffer_14_554 = $signed(_T_100042); // @[Modules.scala 166:64:@48177.4]
  assign _T_100044 = $signed(buffer_14_507) + $signed(buffer_14_508); // @[Modules.scala 166:64:@48179.4]
  assign _T_100045 = _T_100044[13:0]; // @[Modules.scala 166:64:@48180.4]
  assign buffer_14_555 = $signed(_T_100045); // @[Modules.scala 166:64:@48181.4]
  assign _T_100047 = $signed(buffer_14_509) + $signed(buffer_14_510); // @[Modules.scala 166:64:@48183.4]
  assign _T_100048 = _T_100047[13:0]; // @[Modules.scala 166:64:@48184.4]
  assign buffer_14_556 = $signed(_T_100048); // @[Modules.scala 166:64:@48185.4]
  assign _T_100050 = $signed(buffer_14_511) + $signed(buffer_14_512); // @[Modules.scala 166:64:@48187.4]
  assign _T_100051 = _T_100050[13:0]; // @[Modules.scala 166:64:@48188.4]
  assign buffer_14_557 = $signed(_T_100051); // @[Modules.scala 166:64:@48189.4]
  assign _T_100053 = $signed(buffer_14_513) + $signed(buffer_14_514); // @[Modules.scala 166:64:@48191.4]
  assign _T_100054 = _T_100053[13:0]; // @[Modules.scala 166:64:@48192.4]
  assign buffer_14_558 = $signed(_T_100054); // @[Modules.scala 166:64:@48193.4]
  assign _T_100056 = $signed(buffer_14_515) + $signed(buffer_14_516); // @[Modules.scala 166:64:@48195.4]
  assign _T_100057 = _T_100056[13:0]; // @[Modules.scala 166:64:@48196.4]
  assign buffer_14_559 = $signed(_T_100057); // @[Modules.scala 166:64:@48197.4]
  assign _T_100059 = $signed(buffer_14_517) + $signed(buffer_14_518); // @[Modules.scala 166:64:@48199.4]
  assign _T_100060 = _T_100059[13:0]; // @[Modules.scala 166:64:@48200.4]
  assign buffer_14_560 = $signed(_T_100060); // @[Modules.scala 166:64:@48201.4]
  assign _T_100062 = $signed(buffer_14_519) + $signed(buffer_14_520); // @[Modules.scala 166:64:@48203.4]
  assign _T_100063 = _T_100062[13:0]; // @[Modules.scala 166:64:@48204.4]
  assign buffer_14_561 = $signed(_T_100063); // @[Modules.scala 166:64:@48205.4]
  assign _T_100065 = $signed(buffer_14_521) + $signed(buffer_14_522); // @[Modules.scala 166:64:@48207.4]
  assign _T_100066 = _T_100065[13:0]; // @[Modules.scala 166:64:@48208.4]
  assign buffer_14_562 = $signed(_T_100066); // @[Modules.scala 166:64:@48209.4]
  assign _T_100068 = $signed(buffer_14_523) + $signed(buffer_3_545); // @[Modules.scala 166:64:@48211.4]
  assign _T_100069 = _T_100068[13:0]; // @[Modules.scala 166:64:@48212.4]
  assign buffer_14_563 = $signed(_T_100069); // @[Modules.scala 166:64:@48213.4]
  assign _T_100071 = $signed(buffer_14_525) + $signed(buffer_14_526); // @[Modules.scala 166:64:@48215.4]
  assign _T_100072 = _T_100071[13:0]; // @[Modules.scala 166:64:@48216.4]
  assign buffer_14_564 = $signed(_T_100072); // @[Modules.scala 166:64:@48217.4]
  assign _T_100074 = $signed(buffer_14_527) + $signed(buffer_14_452); // @[Modules.scala 172:66:@48219.4]
  assign _T_100075 = _T_100074[13:0]; // @[Modules.scala 172:66:@48220.4]
  assign buffer_14_565 = $signed(_T_100075); // @[Modules.scala 172:66:@48221.4]
  assign _T_100077 = $signed(buffer_14_528) + $signed(buffer_14_529); // @[Modules.scala 160:64:@48223.4]
  assign _T_100078 = _T_100077[13:0]; // @[Modules.scala 160:64:@48224.4]
  assign buffer_14_566 = $signed(_T_100078); // @[Modules.scala 160:64:@48225.4]
  assign _T_100080 = $signed(buffer_14_530) + $signed(buffer_14_531); // @[Modules.scala 160:64:@48227.4]
  assign _T_100081 = _T_100080[13:0]; // @[Modules.scala 160:64:@48228.4]
  assign buffer_14_567 = $signed(_T_100081); // @[Modules.scala 160:64:@48229.4]
  assign _T_100083 = $signed(buffer_14_532) + $signed(buffer_14_533); // @[Modules.scala 160:64:@48231.4]
  assign _T_100084 = _T_100083[13:0]; // @[Modules.scala 160:64:@48232.4]
  assign buffer_14_568 = $signed(_T_100084); // @[Modules.scala 160:64:@48233.4]
  assign _T_100086 = $signed(buffer_14_534) + $signed(buffer_14_535); // @[Modules.scala 160:64:@48235.4]
  assign _T_100087 = _T_100086[13:0]; // @[Modules.scala 160:64:@48236.4]
  assign buffer_14_569 = $signed(_T_100087); // @[Modules.scala 160:64:@48237.4]
  assign _T_100089 = $signed(buffer_14_536) + $signed(buffer_14_537); // @[Modules.scala 160:64:@48239.4]
  assign _T_100090 = _T_100089[13:0]; // @[Modules.scala 160:64:@48240.4]
  assign buffer_14_570 = $signed(_T_100090); // @[Modules.scala 160:64:@48241.4]
  assign _T_100092 = $signed(buffer_14_538) + $signed(buffer_14_539); // @[Modules.scala 160:64:@48243.4]
  assign _T_100093 = _T_100092[13:0]; // @[Modules.scala 160:64:@48244.4]
  assign buffer_14_571 = $signed(_T_100093); // @[Modules.scala 160:64:@48245.4]
  assign _T_100095 = $signed(buffer_14_540) + $signed(buffer_14_541); // @[Modules.scala 160:64:@48247.4]
  assign _T_100096 = _T_100095[13:0]; // @[Modules.scala 160:64:@48248.4]
  assign buffer_14_572 = $signed(_T_100096); // @[Modules.scala 160:64:@48249.4]
  assign _T_100098 = $signed(buffer_14_542) + $signed(buffer_14_543); // @[Modules.scala 160:64:@48251.4]
  assign _T_100099 = _T_100098[13:0]; // @[Modules.scala 160:64:@48252.4]
  assign buffer_14_573 = $signed(_T_100099); // @[Modules.scala 160:64:@48253.4]
  assign _T_100101 = $signed(buffer_14_544) + $signed(buffer_14_545); // @[Modules.scala 160:64:@48255.4]
  assign _T_100102 = _T_100101[13:0]; // @[Modules.scala 160:64:@48256.4]
  assign buffer_14_574 = $signed(_T_100102); // @[Modules.scala 160:64:@48257.4]
  assign _T_100104 = $signed(buffer_14_546) + $signed(buffer_14_547); // @[Modules.scala 160:64:@48259.4]
  assign _T_100105 = _T_100104[13:0]; // @[Modules.scala 160:64:@48260.4]
  assign buffer_14_575 = $signed(_T_100105); // @[Modules.scala 160:64:@48261.4]
  assign _T_100107 = $signed(buffer_14_548) + $signed(buffer_14_549); // @[Modules.scala 160:64:@48263.4]
  assign _T_100108 = _T_100107[13:0]; // @[Modules.scala 160:64:@48264.4]
  assign buffer_14_576 = $signed(_T_100108); // @[Modules.scala 160:64:@48265.4]
  assign _T_100110 = $signed(buffer_14_550) + $signed(buffer_14_551); // @[Modules.scala 160:64:@48267.4]
  assign _T_100111 = _T_100110[13:0]; // @[Modules.scala 160:64:@48268.4]
  assign buffer_14_577 = $signed(_T_100111); // @[Modules.scala 160:64:@48269.4]
  assign _T_100113 = $signed(buffer_14_552) + $signed(buffer_14_553); // @[Modules.scala 160:64:@48271.4]
  assign _T_100114 = _T_100113[13:0]; // @[Modules.scala 160:64:@48272.4]
  assign buffer_14_578 = $signed(_T_100114); // @[Modules.scala 160:64:@48273.4]
  assign _T_100116 = $signed(buffer_14_554) + $signed(buffer_14_555); // @[Modules.scala 160:64:@48275.4]
  assign _T_100117 = _T_100116[13:0]; // @[Modules.scala 160:64:@48276.4]
  assign buffer_14_579 = $signed(_T_100117); // @[Modules.scala 160:64:@48277.4]
  assign _T_100119 = $signed(buffer_14_556) + $signed(buffer_14_557); // @[Modules.scala 160:64:@48279.4]
  assign _T_100120 = _T_100119[13:0]; // @[Modules.scala 160:64:@48280.4]
  assign buffer_14_580 = $signed(_T_100120); // @[Modules.scala 160:64:@48281.4]
  assign _T_100122 = $signed(buffer_14_558) + $signed(buffer_14_559); // @[Modules.scala 160:64:@48283.4]
  assign _T_100123 = _T_100122[13:0]; // @[Modules.scala 160:64:@48284.4]
  assign buffer_14_581 = $signed(_T_100123); // @[Modules.scala 160:64:@48285.4]
  assign _T_100125 = $signed(buffer_14_560) + $signed(buffer_14_561); // @[Modules.scala 160:64:@48287.4]
  assign _T_100126 = _T_100125[13:0]; // @[Modules.scala 160:64:@48288.4]
  assign buffer_14_582 = $signed(_T_100126); // @[Modules.scala 160:64:@48289.4]
  assign _T_100128 = $signed(buffer_14_562) + $signed(buffer_14_563); // @[Modules.scala 160:64:@48291.4]
  assign _T_100129 = _T_100128[13:0]; // @[Modules.scala 160:64:@48292.4]
  assign buffer_14_583 = $signed(_T_100129); // @[Modules.scala 160:64:@48293.4]
  assign _T_100131 = $signed(buffer_14_564) + $signed(buffer_14_565); // @[Modules.scala 160:64:@48295.4]
  assign _T_100132 = _T_100131[13:0]; // @[Modules.scala 160:64:@48296.4]
  assign buffer_14_584 = $signed(_T_100132); // @[Modules.scala 160:64:@48297.4]
  assign _T_100134 = $signed(buffer_14_566) + $signed(buffer_14_567); // @[Modules.scala 166:64:@48299.4]
  assign _T_100135 = _T_100134[13:0]; // @[Modules.scala 166:64:@48300.4]
  assign buffer_14_585 = $signed(_T_100135); // @[Modules.scala 166:64:@48301.4]
  assign _T_100137 = $signed(buffer_14_568) + $signed(buffer_14_569); // @[Modules.scala 166:64:@48303.4]
  assign _T_100138 = _T_100137[13:0]; // @[Modules.scala 166:64:@48304.4]
  assign buffer_14_586 = $signed(_T_100138); // @[Modules.scala 166:64:@48305.4]
  assign _T_100140 = $signed(buffer_14_570) + $signed(buffer_14_571); // @[Modules.scala 166:64:@48307.4]
  assign _T_100141 = _T_100140[13:0]; // @[Modules.scala 166:64:@48308.4]
  assign buffer_14_587 = $signed(_T_100141); // @[Modules.scala 166:64:@48309.4]
  assign _T_100143 = $signed(buffer_14_572) + $signed(buffer_14_573); // @[Modules.scala 166:64:@48311.4]
  assign _T_100144 = _T_100143[13:0]; // @[Modules.scala 166:64:@48312.4]
  assign buffer_14_588 = $signed(_T_100144); // @[Modules.scala 166:64:@48313.4]
  assign _T_100146 = $signed(buffer_14_574) + $signed(buffer_14_575); // @[Modules.scala 166:64:@48315.4]
  assign _T_100147 = _T_100146[13:0]; // @[Modules.scala 166:64:@48316.4]
  assign buffer_14_589 = $signed(_T_100147); // @[Modules.scala 166:64:@48317.4]
  assign _T_100149 = $signed(buffer_14_576) + $signed(buffer_14_577); // @[Modules.scala 166:64:@48319.4]
  assign _T_100150 = _T_100149[13:0]; // @[Modules.scala 166:64:@48320.4]
  assign buffer_14_590 = $signed(_T_100150); // @[Modules.scala 166:64:@48321.4]
  assign _T_100152 = $signed(buffer_14_578) + $signed(buffer_14_579); // @[Modules.scala 166:64:@48323.4]
  assign _T_100153 = _T_100152[13:0]; // @[Modules.scala 166:64:@48324.4]
  assign buffer_14_591 = $signed(_T_100153); // @[Modules.scala 166:64:@48325.4]
  assign _T_100155 = $signed(buffer_14_580) + $signed(buffer_14_581); // @[Modules.scala 166:64:@48327.4]
  assign _T_100156 = _T_100155[13:0]; // @[Modules.scala 166:64:@48328.4]
  assign buffer_14_592 = $signed(_T_100156); // @[Modules.scala 166:64:@48329.4]
  assign _T_100158 = $signed(buffer_14_582) + $signed(buffer_14_583); // @[Modules.scala 166:64:@48331.4]
  assign _T_100159 = _T_100158[13:0]; // @[Modules.scala 166:64:@48332.4]
  assign buffer_14_593 = $signed(_T_100159); // @[Modules.scala 166:64:@48333.4]
  assign _T_100161 = $signed(buffer_14_585) + $signed(buffer_14_586); // @[Modules.scala 166:64:@48335.4]
  assign _T_100162 = _T_100161[13:0]; // @[Modules.scala 166:64:@48336.4]
  assign buffer_14_594 = $signed(_T_100162); // @[Modules.scala 166:64:@48337.4]
  assign _T_100164 = $signed(buffer_14_587) + $signed(buffer_14_588); // @[Modules.scala 166:64:@48339.4]
  assign _T_100165 = _T_100164[13:0]; // @[Modules.scala 166:64:@48340.4]
  assign buffer_14_595 = $signed(_T_100165); // @[Modules.scala 166:64:@48341.4]
  assign _T_100167 = $signed(buffer_14_589) + $signed(buffer_14_590); // @[Modules.scala 166:64:@48343.4]
  assign _T_100168 = _T_100167[13:0]; // @[Modules.scala 166:64:@48344.4]
  assign buffer_14_596 = $signed(_T_100168); // @[Modules.scala 166:64:@48345.4]
  assign _T_100170 = $signed(buffer_14_591) + $signed(buffer_14_592); // @[Modules.scala 166:64:@48347.4]
  assign _T_100171 = _T_100170[13:0]; // @[Modules.scala 166:64:@48348.4]
  assign buffer_14_597 = $signed(_T_100171); // @[Modules.scala 166:64:@48349.4]
  assign _T_100173 = $signed(buffer_14_593) + $signed(buffer_14_584); // @[Modules.scala 172:66:@48351.4]
  assign _T_100174 = _T_100173[13:0]; // @[Modules.scala 172:66:@48352.4]
  assign buffer_14_598 = $signed(_T_100174); // @[Modules.scala 172:66:@48353.4]
  assign _T_100176 = $signed(buffer_14_594) + $signed(buffer_14_595); // @[Modules.scala 166:64:@48355.4]
  assign _T_100177 = _T_100176[13:0]; // @[Modules.scala 166:64:@48356.4]
  assign buffer_14_599 = $signed(_T_100177); // @[Modules.scala 166:64:@48357.4]
  assign _T_100179 = $signed(buffer_14_596) + $signed(buffer_14_597); // @[Modules.scala 166:64:@48359.4]
  assign _T_100180 = _T_100179[13:0]; // @[Modules.scala 166:64:@48360.4]
  assign buffer_14_600 = $signed(_T_100180); // @[Modules.scala 166:64:@48361.4]
  assign _T_100182 = $signed(buffer_14_599) + $signed(buffer_14_600); // @[Modules.scala 160:64:@48363.4]
  assign _T_100183 = _T_100182[13:0]; // @[Modules.scala 160:64:@48364.4]
  assign buffer_14_601 = $signed(_T_100183); // @[Modules.scala 160:64:@48365.4]
  assign _T_100185 = $signed(buffer_14_601) + $signed(buffer_14_598); // @[Modules.scala 172:66:@48367.4]
  assign _T_100186 = _T_100185[13:0]; // @[Modules.scala 172:66:@48368.4]
  assign buffer_14_602 = $signed(_T_100186); // @[Modules.scala 172:66:@48369.4]
  assign _T_100206 = $signed(_T_54215) + $signed(_GEN_633); // @[Modules.scala 143:103:@48566.4]
  assign _T_100207 = _T_100206[5:0]; // @[Modules.scala 143:103:@48567.4]
  assign _T_100208 = $signed(_T_100207); // @[Modules.scala 143:103:@48568.4]
  assign _GEN_1060 = {{1{_T_60334[4]}},_T_60334}; // @[Modules.scala 143:103:@48632.4]
  assign _T_100283 = $signed(_GEN_1060) + $signed(_T_54290); // @[Modules.scala 143:103:@48632.4]
  assign _T_100284 = _T_100283[5:0]; // @[Modules.scala 143:103:@48633.4]
  assign _T_100285 = $signed(_T_100284); // @[Modules.scala 143:103:@48634.4]
  assign _T_100416 = $signed(_T_54423) + $signed(_T_54430); // @[Modules.scala 143:103:@48746.4]
  assign _T_100417 = _T_100416[5:0]; // @[Modules.scala 143:103:@48747.4]
  assign _T_100418 = $signed(_T_100417); // @[Modules.scala 143:103:@48748.4]
  assign _T_100437 = $signed(_GEN_3) + $signed(_T_57451); // @[Modules.scala 143:103:@48764.4]
  assign _T_100438 = _T_100437[5:0]; // @[Modules.scala 143:103:@48765.4]
  assign _T_100439 = $signed(_T_100438); // @[Modules.scala 143:103:@48766.4]
  assign _GEN_1068 = {{1{_T_60563[4]}},_T_60563}; // @[Modules.scala 143:103:@48830.4]
  assign _T_100514 = $signed(_T_54521) + $signed(_GEN_1068); // @[Modules.scala 143:103:@48830.4]
  assign _T_100515 = _T_100514[5:0]; // @[Modules.scala 143:103:@48831.4]
  assign _T_100516 = $signed(_T_100515); // @[Modules.scala 143:103:@48832.4]
  assign _T_100528 = $signed(_T_63683) + $signed(_T_63688); // @[Modules.scala 143:103:@48842.4]
  assign _T_100529 = _T_100528[4:0]; // @[Modules.scala 143:103:@48843.4]
  assign _T_100530 = $signed(_T_100529); // @[Modules.scala 143:103:@48844.4]
  assign _T_100563 = $signed(_T_60605) + $signed(_T_54556); // @[Modules.scala 143:103:@48872.4]
  assign _T_100564 = _T_100563[5:0]; // @[Modules.scala 143:103:@48873.4]
  assign _T_100565 = $signed(_T_100564); // @[Modules.scala 143:103:@48874.4]
  assign _GEN_1069 = {{1{_T_54563[4]}},_T_54563}; // @[Modules.scala 143:103:@48878.4]
  assign _T_100570 = $signed(_T_63730) + $signed(_GEN_1069); // @[Modules.scala 143:103:@48878.4]
  assign _T_100571 = _T_100570[5:0]; // @[Modules.scala 143:103:@48879.4]
  assign _T_100572 = $signed(_T_100571); // @[Modules.scala 143:103:@48880.4]
  assign _GEN_1073 = {{1{_T_63760[4]}},_T_63760}; // @[Modules.scala 143:103:@48902.4]
  assign _T_100598 = $signed(_T_54586) + $signed(_GEN_1073); // @[Modules.scala 143:103:@48902.4]
  assign _T_100599 = _T_100598[5:0]; // @[Modules.scala 143:103:@48903.4]
  assign _T_100600 = $signed(_T_100599); // @[Modules.scala 143:103:@48904.4]
  assign _T_100605 = $signed(_GEN_160) + $signed(_T_54598); // @[Modules.scala 143:103:@48908.4]
  assign _T_100606 = _T_100605[5:0]; // @[Modules.scala 143:103:@48909.4]
  assign _T_100607 = $signed(_T_100606); // @[Modules.scala 143:103:@48910.4]
  assign _T_100633 = $signed(_T_88580) + $signed(_GEN_293); // @[Modules.scala 143:103:@48932.4]
  assign _T_100634 = _T_100633[5:0]; // @[Modules.scala 143:103:@48933.4]
  assign _T_100635 = $signed(_T_100634); // @[Modules.scala 143:103:@48934.4]
  assign _T_100682 = $signed(_GEN_588) + $signed(_T_57715); // @[Modules.scala 143:103:@48974.4]
  assign _T_100683 = _T_100682[5:0]; // @[Modules.scala 143:103:@48975.4]
  assign _T_100684 = $signed(_T_100683); // @[Modules.scala 143:103:@48976.4]
  assign _T_100689 = $signed(_T_54691) + $signed(_T_54698); // @[Modules.scala 143:103:@48980.4]
  assign _T_100690 = _T_100689[4:0]; // @[Modules.scala 143:103:@48981.4]
  assign _T_100691 = $signed(_T_100690); // @[Modules.scala 143:103:@48982.4]
  assign _T_100696 = $signed(_GEN_230) + $signed(_T_63893); // @[Modules.scala 143:103:@48986.4]
  assign _T_100697 = _T_100696[5:0]; // @[Modules.scala 143:103:@48987.4]
  assign _T_100698 = $signed(_T_100697); // @[Modules.scala 143:103:@48988.4]
  assign _T_100731 = $signed(_T_60810) + $signed(_T_60817); // @[Modules.scala 143:103:@49016.4]
  assign _T_100732 = _T_100731[4:0]; // @[Modules.scala 143:103:@49017.4]
  assign _T_100733 = $signed(_T_100732); // @[Modules.scala 143:103:@49018.4]
  assign _T_100745 = $signed(_T_54759) + $signed(_T_60843); // @[Modules.scala 143:103:@49028.4]
  assign _T_100746 = _T_100745[4:0]; // @[Modules.scala 143:103:@49029.4]
  assign _T_100747 = $signed(_T_100746); // @[Modules.scala 143:103:@49030.4]
  assign _T_100752 = $signed(_T_57806) + $signed(_GEN_20); // @[Modules.scala 143:103:@49034.4]
  assign _T_100753 = _T_100752[5:0]; // @[Modules.scala 143:103:@49035.4]
  assign _T_100754 = $signed(_T_100753); // @[Modules.scala 143:103:@49036.4]
  assign _T_100759 = $signed(_T_57815) + $signed(_T_63970); // @[Modules.scala 143:103:@49040.4]
  assign _T_100760 = _T_100759[5:0]; // @[Modules.scala 143:103:@49041.4]
  assign _T_100761 = $signed(_T_100760); // @[Modules.scala 143:103:@49042.4]
  assign _T_100801 = $signed(_T_60901) + $signed(_T_60908); // @[Modules.scala 143:103:@49076.4]
  assign _T_100802 = _T_100801[4:0]; // @[Modules.scala 143:103:@49077.4]
  assign _T_100803 = $signed(_T_100802); // @[Modules.scala 143:103:@49078.4]
  assign _T_100808 = $signed(_T_70148) + $signed(_GEN_453); // @[Modules.scala 143:103:@49082.4]
  assign _T_100809 = _T_100808[5:0]; // @[Modules.scala 143:103:@49083.4]
  assign _T_100810 = $signed(_T_100809); // @[Modules.scala 143:103:@49084.4]
  assign _T_100815 = $signed(_T_54843) + $signed(_T_54852); // @[Modules.scala 143:103:@49088.4]
  assign _T_100816 = _T_100815[4:0]; // @[Modules.scala 143:103:@49089.4]
  assign _T_100817 = $signed(_T_100816); // @[Modules.scala 143:103:@49090.4]
  assign _T_100829 = $signed(_GEN_858) + $signed(_T_70192); // @[Modules.scala 143:103:@49100.4]
  assign _T_100830 = _T_100829[5:0]; // @[Modules.scala 143:103:@49101.4]
  assign _T_100831 = $signed(_T_100830); // @[Modules.scala 143:103:@49102.4]
  assign _T_100857 = $signed(_T_54894) + $signed(_T_60983); // @[Modules.scala 143:103:@49124.4]
  assign _T_100858 = _T_100857[4:0]; // @[Modules.scala 143:103:@49125.4]
  assign _T_100859 = $signed(_T_100858); // @[Modules.scala 143:103:@49126.4]
  assign _GEN_1083 = {{1{_T_54934[4]}},_T_54934}; // @[Modules.scala 143:103:@49136.4]
  assign _T_100871 = $signed(_T_64115) + $signed(_GEN_1083); // @[Modules.scala 143:103:@49136.4]
  assign _T_100872 = _T_100871[5:0]; // @[Modules.scala 143:103:@49137.4]
  assign _T_100873 = $signed(_T_100872); // @[Modules.scala 143:103:@49138.4]
  assign _GEN_1084 = {{1{_T_61018[4]}},_T_61018}; // @[Modules.scala 143:103:@49148.4]
  assign _T_100885 = $signed(_T_54943) + $signed(_GEN_1084); // @[Modules.scala 143:103:@49148.4]
  assign _T_100886 = _T_100885[5:0]; // @[Modules.scala 143:103:@49149.4]
  assign _T_100887 = $signed(_T_100886); // @[Modules.scala 143:103:@49150.4]
  assign _T_100934 = $signed(_T_54985) + $signed(_T_61069); // @[Modules.scala 143:103:@49190.4]
  assign _T_100935 = _T_100934[4:0]; // @[Modules.scala 143:103:@49191.4]
  assign _T_100936 = $signed(_T_100935); // @[Modules.scala 143:103:@49192.4]
  assign _T_101018 = $signed(_T_55081) + $signed(_GEN_239); // @[Modules.scala 143:103:@49262.4]
  assign _T_101019 = _T_101018[5:0]; // @[Modules.scala 143:103:@49263.4]
  assign _T_101020 = $signed(_T_101019); // @[Modules.scala 143:103:@49264.4]
  assign _T_101046 = $signed(_GEN_384) + $signed(_T_58142); // @[Modules.scala 143:103:@49286.4]
  assign _T_101047 = _T_101046[5:0]; // @[Modules.scala 143:103:@49287.4]
  assign _T_101048 = $signed(_T_101047); // @[Modules.scala 143:103:@49288.4]
  assign _GEN_1091 = {{1{_T_70414[4]}},_T_70414}; // @[Modules.scala 143:103:@49292.4]
  assign _T_101053 = $signed(_T_55123) + $signed(_GEN_1091); // @[Modules.scala 143:103:@49292.4]
  assign _T_101054 = _T_101053[5:0]; // @[Modules.scala 143:103:@49293.4]
  assign _T_101055 = $signed(_T_101054); // @[Modules.scala 143:103:@49294.4]
  assign _T_101067 = $signed(_T_73565) + $signed(_T_55139); // @[Modules.scala 143:103:@49304.4]
  assign _T_101068 = _T_101067[4:0]; // @[Modules.scala 143:103:@49305.4]
  assign _T_101069 = $signed(_T_101068); // @[Modules.scala 143:103:@49306.4]
  assign _GEN_1092 = {{1{_T_55144[4]}},_T_55144}; // @[Modules.scala 143:103:@49310.4]
  assign _T_101074 = $signed(_GEN_1092) + $signed(_T_61216); // @[Modules.scala 143:103:@49310.4]
  assign _T_101075 = _T_101074[5:0]; // @[Modules.scala 143:103:@49311.4]
  assign _T_101076 = $signed(_T_101075); // @[Modules.scala 143:103:@49312.4]
  assign _T_101116 = $signed(_T_55186) + $signed(_T_55195); // @[Modules.scala 143:103:@49346.4]
  assign _T_101117 = _T_101116[4:0]; // @[Modules.scala 143:103:@49347.4]
  assign _T_101118 = $signed(_T_101117); // @[Modules.scala 143:103:@49348.4]
  assign _T_101137 = $signed(_T_55214) + $signed(_GEN_387); // @[Modules.scala 143:103:@49364.4]
  assign _T_101138 = _T_101137[5:0]; // @[Modules.scala 143:103:@49365.4]
  assign _T_101139 = $signed(_T_101138); // @[Modules.scala 143:103:@49366.4]
  assign _T_101158 = $signed(_GEN_388) + $signed(_T_55230); // @[Modules.scala 143:103:@49382.4]
  assign _T_101159 = _T_101158[5:0]; // @[Modules.scala 143:103:@49383.4]
  assign _T_101160 = $signed(_T_101159); // @[Modules.scala 143:103:@49384.4]
  assign _T_101165 = $signed(_T_55235) + $signed(_GEN_37); // @[Modules.scala 143:103:@49388.4]
  assign _T_101166 = _T_101165[5:0]; // @[Modules.scala 143:103:@49389.4]
  assign _T_101167 = $signed(_T_101166); // @[Modules.scala 143:103:@49390.4]
  assign _T_101200 = $signed(_T_61363) + $signed(_T_61368); // @[Modules.scala 143:103:@49418.4]
  assign _T_101201 = _T_101200[5:0]; // @[Modules.scala 143:103:@49419.4]
  assign _T_101202 = $signed(_T_101201); // @[Modules.scala 143:103:@49420.4]
  assign _T_101242 = $signed(_GEN_243) + $signed(_T_61403); // @[Modules.scala 143:103:@49454.4]
  assign _T_101243 = _T_101242[5:0]; // @[Modules.scala 143:103:@49455.4]
  assign _T_101244 = $signed(_T_101243); // @[Modules.scala 143:103:@49456.4]
  assign _T_101368 = $signed(_T_89345) + $signed(_T_61522); // @[Modules.scala 143:103:@49562.4]
  assign _T_101369 = _T_101368[5:0]; // @[Modules.scala 143:103:@49563.4]
  assign _T_101370 = $signed(_T_101369); // @[Modules.scala 143:103:@49564.4]
  assign _T_101382 = $signed(_T_55445) + $signed(_GEN_400); // @[Modules.scala 143:103:@49574.4]
  assign _T_101383 = _T_101382[5:0]; // @[Modules.scala 143:103:@49575.4]
  assign _T_101384 = $signed(_T_101383); // @[Modules.scala 143:103:@49576.4]
  assign _T_101417 = $signed(_GEN_402) + $signed(_T_58485); // @[Modules.scala 143:103:@49604.4]
  assign _T_101418 = _T_101417[5:0]; // @[Modules.scala 143:103:@49605.4]
  assign _T_101419 = $signed(_T_101418); // @[Modules.scala 143:103:@49606.4]
  assign _T_101459 = $signed(_T_61601) + $signed(_T_55510); // @[Modules.scala 143:103:@49640.4]
  assign _T_101460 = _T_101459[5:0]; // @[Modules.scala 143:103:@49641.4]
  assign _T_101461 = $signed(_T_101460); // @[Modules.scala 143:103:@49642.4]
  assign _GEN_1110 = {{1{_T_58548[4]}},_T_58548}; // @[Modules.scala 143:103:@49646.4]
  assign _T_101466 = $signed(_T_55515) + $signed(_GEN_1110); // @[Modules.scala 143:103:@49646.4]
  assign _T_101467 = _T_101466[5:0]; // @[Modules.scala 143:103:@49647.4]
  assign _T_101468 = $signed(_T_101467); // @[Modules.scala 143:103:@49648.4]
  assign _T_101473 = $signed(_T_58550) + $signed(_T_55529); // @[Modules.scala 143:103:@49652.4]
  assign _T_101474 = _T_101473[4:0]; // @[Modules.scala 143:103:@49653.4]
  assign _T_101475 = $signed(_T_101474); // @[Modules.scala 143:103:@49654.4]
  assign _T_101480 = $signed(_GEN_331) + $signed(_T_58557); // @[Modules.scala 143:103:@49658.4]
  assign _T_101481 = _T_101480[5:0]; // @[Modules.scala 143:103:@49659.4]
  assign _T_101482 = $signed(_T_101481); // @[Modules.scala 143:103:@49660.4]
  assign _T_101536 = $signed(_T_64796) + $signed(_T_70876); // @[Modules.scala 143:103:@49706.4]
  assign _T_101537 = _T_101536[5:0]; // @[Modules.scala 143:103:@49707.4]
  assign _T_101538 = $signed(_T_101537); // @[Modules.scala 143:103:@49708.4]
  assign _T_101564 = $signed(_T_70897) + $signed(_T_55608); // @[Modules.scala 143:103:@49730.4]
  assign _T_101565 = _T_101564[4:0]; // @[Modules.scala 143:103:@49731.4]
  assign _T_101566 = $signed(_T_101565); // @[Modules.scala 143:103:@49732.4]
  assign _T_101627 = $signed(_T_55664) + $signed(_T_70960); // @[Modules.scala 143:103:@49784.4]
  assign _T_101628 = _T_101627[5:0]; // @[Modules.scala 143:103:@49785.4]
  assign _T_101629 = $signed(_T_101628); // @[Modules.scala 143:103:@49786.4]
  assign _T_101697 = $signed(_T_55718) + $signed(_GEN_261); // @[Modules.scala 143:103:@49844.4]
  assign _T_101698 = _T_101697[5:0]; // @[Modules.scala 143:103:@49845.4]
  assign _T_101699 = $signed(_T_101698); // @[Modules.scala 143:103:@49846.4]
  assign _T_101704 = $signed(_T_55725) + $signed(_T_64950); // @[Modules.scala 143:103:@49850.4]
  assign _T_101705 = _T_101704[4:0]; // @[Modules.scala 143:103:@49851.4]
  assign _T_101706 = $signed(_T_101705); // @[Modules.scala 143:103:@49852.4]
  assign _T_101753 = $signed(_T_61846) + $signed(_T_61851); // @[Modules.scala 143:103:@49892.4]
  assign _T_101754 = _T_101753[5:0]; // @[Modules.scala 143:103:@49893.4]
  assign _T_101755 = $signed(_T_101754); // @[Modules.scala 143:103:@49894.4]
  assign _T_101760 = $signed(_T_74260) + $signed(_T_55767); // @[Modules.scala 143:103:@49898.4]
  assign _T_101761 = _T_101760[5:0]; // @[Modules.scala 143:103:@49899.4]
  assign _T_101762 = $signed(_T_101761); // @[Modules.scala 143:103:@49900.4]
  assign _GEN_1118 = {{1{_T_61900[4]}},_T_61900}; // @[Modules.scala 143:103:@49940.4]
  assign _T_101809 = $signed(_T_55802) + $signed(_GEN_1118); // @[Modules.scala 143:103:@49940.4]
  assign _T_101810 = _T_101809[5:0]; // @[Modules.scala 143:103:@49941.4]
  assign _T_101811 = $signed(_T_101810); // @[Modules.scala 143:103:@49942.4]
  assign _T_101851 = $signed(_T_55832) + $signed(_T_74323); // @[Modules.scala 143:103:@49976.4]
  assign _T_101852 = _T_101851[5:0]; // @[Modules.scala 143:103:@49977.4]
  assign _T_101853 = $signed(_T_101852); // @[Modules.scala 143:103:@49978.4]
  assign _T_101879 = $signed(_T_55846) + $signed(_GEN_201); // @[Modules.scala 143:103:@50000.4]
  assign _T_101880 = _T_101879[5:0]; // @[Modules.scala 143:103:@50001.4]
  assign _T_101881 = $signed(_T_101880); // @[Modules.scala 143:103:@50002.4]
  assign _T_101890 = $signed(-4'sh1) * $signed(io_in_615); // @[Modules.scala 143:74:@50010.4]
  assign _T_101893 = $signed(_T_101890) + $signed(_T_58886); // @[Modules.scala 143:103:@50012.4]
  assign _T_101894 = _T_101893[4:0]; // @[Modules.scala 143:103:@50013.4]
  assign _T_101895 = $signed(_T_101894); // @[Modules.scala 143:103:@50014.4]
  assign _T_101928 = $signed(_T_71235) + $signed(_T_71242); // @[Modules.scala 143:103:@50042.4]
  assign _T_101929 = _T_101928[5:0]; // @[Modules.scala 143:103:@50043.4]
  assign _T_101930 = $signed(_T_101929); // @[Modules.scala 143:103:@50044.4]
  assign _T_101935 = $signed(_T_71247) + $signed(_GEN_419); // @[Modules.scala 143:103:@50048.4]
  assign _T_101936 = _T_101935[5:0]; // @[Modules.scala 143:103:@50049.4]
  assign _T_101937 = $signed(_T_101936); // @[Modules.scala 143:103:@50050.4]
  assign _T_101963 = $signed(_GEN_132) + $signed(_T_55944); // @[Modules.scala 143:103:@50072.4]
  assign _T_101964 = _T_101963[5:0]; // @[Modules.scala 143:103:@50073.4]
  assign _T_101965 = $signed(_T_101964); // @[Modules.scala 143:103:@50074.4]
  assign _GEN_1125 = {{1{_T_55970[4]}},_T_55970}; // @[Modules.scala 143:103:@50090.4]
  assign _T_101984 = $signed(_T_55963) + $signed(_GEN_1125); // @[Modules.scala 143:103:@50090.4]
  assign _T_101985 = _T_101984[5:0]; // @[Modules.scala 143:103:@50091.4]
  assign _T_101986 = $signed(_T_101985); // @[Modules.scala 143:103:@50092.4]
  assign _T_102012 = $signed(_T_65195) + $signed(_T_59003); // @[Modules.scala 143:103:@50114.4]
  assign _T_102013 = _T_102012[5:0]; // @[Modules.scala 143:103:@50115.4]
  assign _T_102014 = $signed(_T_102013); // @[Modules.scala 143:103:@50116.4]
  assign _T_102152 = $signed(_GEN_211) + $signed(_T_59152); // @[Modules.scala 143:103:@50234.4]
  assign _T_102153 = _T_102152[5:0]; // @[Modules.scala 143:103:@50235.4]
  assign _T_102154 = $signed(_T_102153); // @[Modules.scala 143:103:@50236.4]
  assign _T_102208 = $signed(_T_59194) + $signed(_T_59199); // @[Modules.scala 143:103:@50282.4]
  assign _T_102209 = _T_102208[4:0]; // @[Modules.scala 143:103:@50283.4]
  assign _T_102210 = $signed(_T_102209); // @[Modules.scala 143:103:@50284.4]
  assign _T_102313 = $signed(_T_71625) + $signed(_GEN_974); // @[Modules.scala 143:103:@50372.4]
  assign _T_102314 = _T_102313[5:0]; // @[Modules.scala 143:103:@50373.4]
  assign _T_102315 = $signed(_T_102314); // @[Modules.scala 143:103:@50374.4]
  assign _T_102341 = $signed(_GEN_693) + $signed(_T_56301); // @[Modules.scala 143:103:@50396.4]
  assign _T_102342 = _T_102341[5:0]; // @[Modules.scala 143:103:@50397.4]
  assign _T_102343 = $signed(_T_102342); // @[Modules.scala 143:103:@50398.4]
  assign _T_102344 = $signed(buffer_0_0) + $signed(buffer_2_1); // @[Modules.scala 160:64:@50400.4]
  assign _T_102345 = _T_102344[13:0]; // @[Modules.scala 160:64:@50401.4]
  assign buffer_15_308 = $signed(_T_102345); // @[Modules.scala 160:64:@50402.4]
  assign buffer_15_2 = {{8{_T_100208[5]}},_T_100208}; // @[Modules.scala 112:22:@8.4]
  assign _T_102347 = $signed(buffer_15_2) + $signed(buffer_10_3); // @[Modules.scala 160:64:@50404.4]
  assign _T_102348 = _T_102347[13:0]; // @[Modules.scala 160:64:@50405.4]
  assign buffer_15_309 = $signed(_T_102348); // @[Modules.scala 160:64:@50406.4]
  assign buffer_15_13 = {{8{_T_100285[5]}},_T_100285}; // @[Modules.scala 112:22:@8.4]
  assign _T_102362 = $signed(buffer_14_12) + $signed(buffer_15_13); // @[Modules.scala 160:64:@50424.4]
  assign _T_102363 = _T_102362[13:0]; // @[Modules.scala 160:64:@50425.4]
  assign buffer_15_314 = $signed(_T_102363); // @[Modules.scala 160:64:@50426.4]
  assign _T_102380 = $signed(buffer_14_24) + $signed(buffer_2_23); // @[Modules.scala 160:64:@50448.4]
  assign _T_102381 = _T_102380[13:0]; // @[Modules.scala 160:64:@50449.4]
  assign buffer_15_320 = $signed(_T_102381); // @[Modules.scala 160:64:@50450.4]
  assign buffer_15_32 = {{8{_T_100418[5]}},_T_100418}; // @[Modules.scala 112:22:@8.4]
  assign _T_102392 = $signed(buffer_15_32) + $signed(buffer_7_33); // @[Modules.scala 160:64:@50464.4]
  assign _T_102393 = _T_102392[13:0]; // @[Modules.scala 160:64:@50465.4]
  assign buffer_15_324 = $signed(_T_102393); // @[Modules.scala 160:64:@50466.4]
  assign buffer_15_35 = {{8{_T_100439[5]}},_T_100439}; // @[Modules.scala 112:22:@8.4]
  assign _T_102395 = $signed(buffer_14_35) + $signed(buffer_15_35); // @[Modules.scala 160:64:@50468.4]
  assign _T_102396 = _T_102395[13:0]; // @[Modules.scala 160:64:@50469.4]
  assign buffer_15_325 = $signed(_T_102396); // @[Modules.scala 160:64:@50470.4]
  assign _T_102410 = $signed(buffer_4_41) + $signed(buffer_11_44); // @[Modules.scala 160:64:@50488.4]
  assign _T_102411 = _T_102410[13:0]; // @[Modules.scala 160:64:@50489.4]
  assign buffer_15_330 = $signed(_T_102411); // @[Modules.scala 160:64:@50490.4]
  assign buffer_15_46 = {{8{_T_100516[5]}},_T_100516}; // @[Modules.scala 112:22:@8.4]
  assign _T_102413 = $signed(buffer_15_46) + $signed(buffer_10_48); // @[Modules.scala 160:64:@50492.4]
  assign _T_102414 = _T_102413[13:0]; // @[Modules.scala 160:64:@50493.4]
  assign buffer_15_331 = $signed(_T_102414); // @[Modules.scala 160:64:@50494.4]
  assign buffer_15_48 = {{9{_T_100530[4]}},_T_100530}; // @[Modules.scala 112:22:@8.4]
  assign _T_102416 = $signed(buffer_15_48) + $signed(buffer_1_49); // @[Modules.scala 160:64:@50496.4]
  assign _T_102417 = _T_102416[13:0]; // @[Modules.scala 160:64:@50497.4]
  assign buffer_15_332 = $signed(_T_102417); // @[Modules.scala 160:64:@50498.4]
  assign buffer_15_53 = {{8{_T_100565[5]}},_T_100565}; // @[Modules.scala 112:22:@8.4]
  assign _T_102422 = $signed(buffer_7_51) + $signed(buffer_15_53); // @[Modules.scala 160:64:@50504.4]
  assign _T_102423 = _T_102422[13:0]; // @[Modules.scala 160:64:@50505.4]
  assign buffer_15_334 = $signed(_T_102423); // @[Modules.scala 160:64:@50506.4]
  assign buffer_15_54 = {{8{_T_100572[5]}},_T_100572}; // @[Modules.scala 112:22:@8.4]
  assign _T_102425 = $signed(buffer_15_54) + $signed(buffer_5_55); // @[Modules.scala 160:64:@50508.4]
  assign _T_102426 = _T_102425[13:0]; // @[Modules.scala 160:64:@50509.4]
  assign buffer_15_335 = $signed(_T_102426); // @[Modules.scala 160:64:@50510.4]
  assign _T_102428 = $signed(buffer_3_57) + $signed(buffer_11_56); // @[Modules.scala 160:64:@50512.4]
  assign _T_102429 = _T_102428[13:0]; // @[Modules.scala 160:64:@50513.4]
  assign buffer_15_336 = $signed(_T_102429); // @[Modules.scala 160:64:@50514.4]
  assign buffer_15_58 = {{8{_T_100600[5]}},_T_100600}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_59 = {{8{_T_100607[5]}},_T_100607}; // @[Modules.scala 112:22:@8.4]
  assign _T_102431 = $signed(buffer_15_58) + $signed(buffer_15_59); // @[Modules.scala 160:64:@50516.4]
  assign _T_102432 = _T_102431[13:0]; // @[Modules.scala 160:64:@50517.4]
  assign buffer_15_337 = $signed(_T_102432); // @[Modules.scala 160:64:@50518.4]
  assign buffer_15_63 = {{8{_T_100635[5]}},_T_100635}; // @[Modules.scala 112:22:@8.4]
  assign _T_102437 = $signed(buffer_5_63) + $signed(buffer_15_63); // @[Modules.scala 160:64:@50524.4]
  assign _T_102438 = _T_102437[13:0]; // @[Modules.scala 160:64:@50525.4]
  assign buffer_15_339 = $signed(_T_102438); // @[Modules.scala 160:64:@50526.4]
  assign _T_102440 = $signed(buffer_1_64) + $signed(buffer_3_68); // @[Modules.scala 160:64:@50528.4]
  assign _T_102441 = _T_102440[13:0]; // @[Modules.scala 160:64:@50529.4]
  assign buffer_15_340 = $signed(_T_102441); // @[Modules.scala 160:64:@50530.4]
  assign _T_102443 = $signed(buffer_7_66) + $signed(buffer_5_68); // @[Modules.scala 160:64:@50532.4]
  assign _T_102444 = _T_102443[13:0]; // @[Modules.scala 160:64:@50533.4]
  assign buffer_15_341 = $signed(_T_102444); // @[Modules.scala 160:64:@50534.4]
  assign _T_102446 = $signed(buffer_3_70) + $signed(buffer_6_70); // @[Modules.scala 160:64:@50536.4]
  assign _T_102447 = _T_102446[13:0]; // @[Modules.scala 160:64:@50537.4]
  assign buffer_15_342 = $signed(_T_102447); // @[Modules.scala 160:64:@50538.4]
  assign buffer_15_70 = {{8{_T_100684[5]}},_T_100684}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_71 = {{9{_T_100691[4]}},_T_100691}; // @[Modules.scala 112:22:@8.4]
  assign _T_102449 = $signed(buffer_15_70) + $signed(buffer_15_71); // @[Modules.scala 160:64:@50540.4]
  assign _T_102450 = _T_102449[13:0]; // @[Modules.scala 160:64:@50541.4]
  assign buffer_15_343 = $signed(_T_102450); // @[Modules.scala 160:64:@50542.4]
  assign buffer_15_72 = {{8{_T_100698[5]}},_T_100698}; // @[Modules.scala 112:22:@8.4]
  assign _T_102452 = $signed(buffer_15_72) + $signed(buffer_3_79); // @[Modules.scala 160:64:@50544.4]
  assign _T_102453 = _T_102452[13:0]; // @[Modules.scala 160:64:@50545.4]
  assign buffer_15_344 = $signed(_T_102453); // @[Modules.scala 160:64:@50546.4]
  assign _T_102455 = $signed(buffer_3_80) + $signed(buffer_0_75); // @[Modules.scala 160:64:@50548.4]
  assign _T_102456 = _T_102455[13:0]; // @[Modules.scala 160:64:@50549.4]
  assign buffer_15_345 = $signed(_T_102456); // @[Modules.scala 160:64:@50550.4]
  assign buffer_15_77 = {{9{_T_100733[4]}},_T_100733}; // @[Modules.scala 112:22:@8.4]
  assign _T_102458 = $signed(buffer_10_77) + $signed(buffer_15_77); // @[Modules.scala 160:64:@50552.4]
  assign _T_102459 = _T_102458[13:0]; // @[Modules.scala 160:64:@50553.4]
  assign buffer_15_346 = $signed(_T_102459); // @[Modules.scala 160:64:@50554.4]
  assign buffer_15_79 = {{9{_T_100747[4]}},_T_100747}; // @[Modules.scala 112:22:@8.4]
  assign _T_102461 = $signed(buffer_9_84) + $signed(buffer_15_79); // @[Modules.scala 160:64:@50556.4]
  assign _T_102462 = _T_102461[13:0]; // @[Modules.scala 160:64:@50557.4]
  assign buffer_15_347 = $signed(_T_102462); // @[Modules.scala 160:64:@50558.4]
  assign buffer_15_80 = {{8{_T_100754[5]}},_T_100754}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_81 = {{8{_T_100761[5]}},_T_100761}; // @[Modules.scala 112:22:@8.4]
  assign _T_102464 = $signed(buffer_15_80) + $signed(buffer_15_81); // @[Modules.scala 160:64:@50560.4]
  assign _T_102465 = _T_102464[13:0]; // @[Modules.scala 160:64:@50561.4]
  assign buffer_15_348 = $signed(_T_102465); // @[Modules.scala 160:64:@50562.4]
  assign _T_102470 = $signed(buffer_5_92) + $signed(buffer_0_87); // @[Modules.scala 160:64:@50568.4]
  assign _T_102471 = _T_102470[13:0]; // @[Modules.scala 160:64:@50569.4]
  assign buffer_15_350 = $signed(_T_102471); // @[Modules.scala 160:64:@50570.4]
  assign buffer_15_87 = {{9{_T_100803[4]}},_T_100803}; // @[Modules.scala 112:22:@8.4]
  assign _T_102473 = $signed(buffer_3_93) + $signed(buffer_15_87); // @[Modules.scala 160:64:@50572.4]
  assign _T_102474 = _T_102473[13:0]; // @[Modules.scala 160:64:@50573.4]
  assign buffer_15_351 = $signed(_T_102474); // @[Modules.scala 160:64:@50574.4]
  assign buffer_15_88 = {{8{_T_100810[5]}},_T_100810}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_89 = {{9{_T_100817[4]}},_T_100817}; // @[Modules.scala 112:22:@8.4]
  assign _T_102476 = $signed(buffer_15_88) + $signed(buffer_15_89); // @[Modules.scala 160:64:@50576.4]
  assign _T_102477 = _T_102476[13:0]; // @[Modules.scala 160:64:@50577.4]
  assign buffer_15_352 = $signed(_T_102477); // @[Modules.scala 160:64:@50578.4]
  assign buffer_15_91 = {{8{_T_100831[5]}},_T_100831}; // @[Modules.scala 112:22:@8.4]
  assign _T_102479 = $signed(buffer_0_94) + $signed(buffer_15_91); // @[Modules.scala 160:64:@50580.4]
  assign _T_102480 = _T_102479[13:0]; // @[Modules.scala 160:64:@50581.4]
  assign buffer_15_353 = $signed(_T_102480); // @[Modules.scala 160:64:@50582.4]
  assign buffer_15_95 = {{9{_T_100859[4]}},_T_100859}; // @[Modules.scala 112:22:@8.4]
  assign _T_102485 = $signed(buffer_5_106) + $signed(buffer_15_95); // @[Modules.scala 160:64:@50588.4]
  assign _T_102486 = _T_102485[13:0]; // @[Modules.scala 160:64:@50589.4]
  assign buffer_15_355 = $signed(_T_102486); // @[Modules.scala 160:64:@50590.4]
  assign buffer_15_97 = {{8{_T_100873[5]}},_T_100873}; // @[Modules.scala 112:22:@8.4]
  assign _T_102488 = $signed(buffer_10_104) + $signed(buffer_15_97); // @[Modules.scala 160:64:@50592.4]
  assign _T_102489 = _T_102488[13:0]; // @[Modules.scala 160:64:@50593.4]
  assign buffer_15_356 = $signed(_T_102489); // @[Modules.scala 160:64:@50594.4]
  assign buffer_15_99 = {{8{_T_100887[5]}},_T_100887}; // @[Modules.scala 112:22:@8.4]
  assign _T_102491 = $signed(buffer_9_113) + $signed(buffer_15_99); // @[Modules.scala 160:64:@50596.4]
  assign _T_102492 = _T_102491[13:0]; // @[Modules.scala 160:64:@50597.4]
  assign buffer_15_357 = $signed(_T_102492); // @[Modules.scala 160:64:@50598.4]
  assign _T_102494 = $signed(buffer_3_113) + $signed(buffer_0_108); // @[Modules.scala 160:64:@50600.4]
  assign _T_102495 = _T_102494[13:0]; // @[Modules.scala 160:64:@50601.4]
  assign buffer_15_358 = $signed(_T_102495); // @[Modules.scala 160:64:@50602.4]
  assign _T_102497 = $signed(buffer_0_109) + $signed(buffer_13_113); // @[Modules.scala 160:64:@50604.4]
  assign _T_102498 = _T_102497[13:0]; // @[Modules.scala 160:64:@50605.4]
  assign buffer_15_359 = $signed(_T_102498); // @[Modules.scala 160:64:@50606.4]
  assign _T_102500 = $signed(buffer_3_117) + $signed(buffer_3_118); // @[Modules.scala 160:64:@50608.4]
  assign _T_102501 = _T_102500[13:0]; // @[Modules.scala 160:64:@50609.4]
  assign buffer_15_360 = $signed(_T_102501); // @[Modules.scala 160:64:@50610.4]
  assign buffer_15_106 = {{9{_T_100936[4]}},_T_100936}; // @[Modules.scala 112:22:@8.4]
  assign _T_102503 = $signed(buffer_15_106) + $signed(buffer_2_118); // @[Modules.scala 160:64:@50612.4]
  assign _T_102504 = _T_102503[13:0]; // @[Modules.scala 160:64:@50613.4]
  assign buffer_15_361 = $signed(_T_102504); // @[Modules.scala 160:64:@50614.4]
  assign _T_102506 = $signed(buffer_0_116) + $signed(buffer_1_119); // @[Modules.scala 160:64:@50616.4]
  assign _T_102507 = _T_102506[13:0]; // @[Modules.scala 160:64:@50617.4]
  assign buffer_15_362 = $signed(_T_102507); // @[Modules.scala 160:64:@50618.4]
  assign _T_102509 = $signed(buffer_1_120) + $signed(buffer_3_126); // @[Modules.scala 160:64:@50620.4]
  assign _T_102510 = _T_102509[13:0]; // @[Modules.scala 160:64:@50621.4]
  assign buffer_15_363 = $signed(_T_102510); // @[Modules.scala 160:64:@50622.4]
  assign _T_102515 = $signed(buffer_0_122) + $signed(buffer_5_126); // @[Modules.scala 160:64:@50628.4]
  assign _T_102516 = _T_102515[13:0]; // @[Modules.scala 160:64:@50629.4]
  assign buffer_15_365 = $signed(_T_102516); // @[Modules.scala 160:64:@50630.4]
  assign _T_102518 = $signed(buffer_3_131) + $signed(buffer_0_125); // @[Modules.scala 160:64:@50632.4]
  assign _T_102519 = _T_102518[13:0]; // @[Modules.scala 160:64:@50633.4]
  assign buffer_15_366 = $signed(_T_102519); // @[Modules.scala 160:64:@50634.4]
  assign buffer_15_118 = {{8{_T_101020[5]}},_T_101020}; // @[Modules.scala 112:22:@8.4]
  assign _T_102521 = $signed(buffer_15_118) + $signed(buffer_0_127); // @[Modules.scala 160:64:@50636.4]
  assign _T_102522 = _T_102521[13:0]; // @[Modules.scala 160:64:@50637.4]
  assign buffer_15_367 = $signed(_T_102522); // @[Modules.scala 160:64:@50638.4]
  assign _T_102524 = $signed(buffer_0_128) + $signed(buffer_1_131); // @[Modules.scala 160:64:@50640.4]
  assign _T_102525 = _T_102524[13:0]; // @[Modules.scala 160:64:@50641.4]
  assign buffer_15_368 = $signed(_T_102525); // @[Modules.scala 160:64:@50642.4]
  assign buffer_15_122 = {{8{_T_101048[5]}},_T_101048}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_123 = {{8{_T_101055[5]}},_T_101055}; // @[Modules.scala 112:22:@8.4]
  assign _T_102527 = $signed(buffer_15_122) + $signed(buffer_15_123); // @[Modules.scala 160:64:@50644.4]
  assign _T_102528 = _T_102527[13:0]; // @[Modules.scala 160:64:@50645.4]
  assign buffer_15_369 = $signed(_T_102528); // @[Modules.scala 160:64:@50646.4]
  assign buffer_15_125 = {{9{_T_101069[4]}},_T_101069}; // @[Modules.scala 112:22:@8.4]
  assign _T_102530 = $signed(buffer_0_133) + $signed(buffer_15_125); // @[Modules.scala 160:64:@50648.4]
  assign _T_102531 = _T_102530[13:0]; // @[Modules.scala 160:64:@50649.4]
  assign buffer_15_370 = $signed(_T_102531); // @[Modules.scala 160:64:@50650.4]
  assign buffer_15_126 = {{8{_T_101076[5]}},_T_101076}; // @[Modules.scala 112:22:@8.4]
  assign _T_102533 = $signed(buffer_15_126) + $signed(buffer_11_131); // @[Modules.scala 160:64:@50652.4]
  assign _T_102534 = _T_102533[13:0]; // @[Modules.scala 160:64:@50653.4]
  assign buffer_15_371 = $signed(_T_102534); // @[Modules.scala 160:64:@50654.4]
  assign buffer_15_132 = {{9{_T_101118[4]}},_T_101118}; // @[Modules.scala 112:22:@8.4]
  assign _T_102542 = $signed(buffer_15_132) + $signed(buffer_0_143); // @[Modules.scala 160:64:@50664.4]
  assign _T_102543 = _T_102542[13:0]; // @[Modules.scala 160:64:@50665.4]
  assign buffer_15_374 = $signed(_T_102543); // @[Modules.scala 160:64:@50666.4]
  assign buffer_15_135 = {{8{_T_101139[5]}},_T_101139}; // @[Modules.scala 112:22:@8.4]
  assign _T_102545 = $signed(buffer_2_147) + $signed(buffer_15_135); // @[Modules.scala 160:64:@50668.4]
  assign _T_102546 = _T_102545[13:0]; // @[Modules.scala 160:64:@50669.4]
  assign buffer_15_375 = $signed(_T_102546); // @[Modules.scala 160:64:@50670.4]
  assign _T_102548 = $signed(buffer_7_145) + $signed(buffer_6_151); // @[Modules.scala 160:64:@50672.4]
  assign _T_102549 = _T_102548[13:0]; // @[Modules.scala 160:64:@50673.4]
  assign buffer_15_376 = $signed(_T_102549); // @[Modules.scala 160:64:@50674.4]
  assign buffer_15_138 = {{8{_T_101160[5]}},_T_101160}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_139 = {{8{_T_101167[5]}},_T_101167}; // @[Modules.scala 112:22:@8.4]
  assign _T_102551 = $signed(buffer_15_138) + $signed(buffer_15_139); // @[Modules.scala 160:64:@50676.4]
  assign _T_102552 = _T_102551[13:0]; // @[Modules.scala 160:64:@50677.4]
  assign buffer_15_377 = $signed(_T_102552); // @[Modules.scala 160:64:@50678.4]
  assign _T_102554 = $signed(buffer_7_150) + $signed(buffer_2_155); // @[Modules.scala 160:64:@50680.4]
  assign _T_102555 = _T_102554[13:0]; // @[Modules.scala 160:64:@50681.4]
  assign buffer_15_378 = $signed(_T_102555); // @[Modules.scala 160:64:@50682.4]
  assign buffer_15_144 = {{8{_T_101202[5]}},_T_101202}; // @[Modules.scala 112:22:@8.4]
  assign _T_102560 = $signed(buffer_15_144) + $signed(buffer_3_163); // @[Modules.scala 160:64:@50688.4]
  assign _T_102561 = _T_102560[13:0]; // @[Modules.scala 160:64:@50689.4]
  assign buffer_15_380 = $signed(_T_102561); // @[Modules.scala 160:64:@50690.4]
  assign _T_102563 = $signed(buffer_14_145) + $signed(buffer_7_158); // @[Modules.scala 160:64:@50692.4]
  assign _T_102564 = _T_102563[13:0]; // @[Modules.scala 160:64:@50693.4]
  assign buffer_15_381 = $signed(_T_102564); // @[Modules.scala 160:64:@50694.4]
  assign _T_102566 = $signed(buffer_7_159) + $signed(buffer_6_165); // @[Modules.scala 160:64:@50696.4]
  assign _T_102567 = _T_102566[13:0]; // @[Modules.scala 160:64:@50697.4]
  assign buffer_15_382 = $signed(_T_102567); // @[Modules.scala 160:64:@50698.4]
  assign buffer_15_150 = {{8{_T_101244[5]}},_T_101244}; // @[Modules.scala 112:22:@8.4]
  assign _T_102569 = $signed(buffer_15_150) + $signed(buffer_10_164); // @[Modules.scala 160:64:@50700.4]
  assign _T_102570 = _T_102569[13:0]; // @[Modules.scala 160:64:@50701.4]
  assign buffer_15_383 = $signed(_T_102570); // @[Modules.scala 160:64:@50702.4]
  assign _T_102572 = $signed(buffer_5_163) + $signed(buffer_5_164); // @[Modules.scala 160:64:@50704.4]
  assign _T_102573 = _T_102572[13:0]; // @[Modules.scala 160:64:@50705.4]
  assign buffer_15_384 = $signed(_T_102573); // @[Modules.scala 160:64:@50706.4]
  assign _T_102578 = $signed(buffer_9_172) + $signed(buffer_8_165); // @[Modules.scala 160:64:@50712.4]
  assign _T_102579 = _T_102578[13:0]; // @[Modules.scala 160:64:@50713.4]
  assign buffer_15_386 = $signed(_T_102579); // @[Modules.scala 160:64:@50714.4]
  assign _T_102587 = $signed(buffer_3_177) + $signed(buffer_9_178); // @[Modules.scala 160:64:@50724.4]
  assign _T_102588 = _T_102587[13:0]; // @[Modules.scala 160:64:@50725.4]
  assign buffer_15_389 = $signed(_T_102588); // @[Modules.scala 160:64:@50726.4]
  assign _T_102590 = $signed(buffer_7_176) + $signed(buffer_1_173); // @[Modules.scala 160:64:@50728.4]
  assign _T_102591 = _T_102590[13:0]; // @[Modules.scala 160:64:@50729.4]
  assign buffer_15_390 = $signed(_T_102591); // @[Modules.scala 160:64:@50730.4]
  assign _T_102593 = $signed(buffer_1_174) + $signed(buffer_9_182); // @[Modules.scala 160:64:@50732.4]
  assign _T_102594 = _T_102593[13:0]; // @[Modules.scala 160:64:@50733.4]
  assign buffer_15_391 = $signed(_T_102594); // @[Modules.scala 160:64:@50734.4]
  assign buffer_15_168 = {{8{_T_101370[5]}},_T_101370}; // @[Modules.scala 112:22:@8.4]
  assign _T_102596 = $signed(buffer_15_168) + $signed(buffer_1_177); // @[Modules.scala 160:64:@50736.4]
  assign _T_102597 = _T_102596[13:0]; // @[Modules.scala 160:64:@50737.4]
  assign buffer_15_392 = $signed(_T_102597); // @[Modules.scala 160:64:@50738.4]
  assign buffer_15_170 = {{8{_T_101384[5]}},_T_101384}; // @[Modules.scala 112:22:@8.4]
  assign _T_102599 = $signed(buffer_15_170) + $signed(buffer_6_185); // @[Modules.scala 160:64:@50740.4]
  assign _T_102600 = _T_102599[13:0]; // @[Modules.scala 160:64:@50741.4]
  assign buffer_15_393 = $signed(_T_102600); // @[Modules.scala 160:64:@50742.4]
  assign _T_102602 = $signed(buffer_12_171) + $signed(buffer_12_172); // @[Modules.scala 160:64:@50744.4]
  assign _T_102603 = _T_102602[13:0]; // @[Modules.scala 160:64:@50745.4]
  assign buffer_15_394 = $signed(_T_102603); // @[Modules.scala 160:64:@50746.4]
  assign buffer_15_175 = {{8{_T_101419[5]}},_T_101419}; // @[Modules.scala 112:22:@8.4]
  assign _T_102605 = $signed(buffer_0_181) + $signed(buffer_15_175); // @[Modules.scala 160:64:@50748.4]
  assign _T_102606 = _T_102605[13:0]; // @[Modules.scala 160:64:@50749.4]
  assign buffer_15_395 = $signed(_T_102606); // @[Modules.scala 160:64:@50750.4]
  assign _T_102611 = $signed(buffer_10_191) + $signed(buffer_0_185); // @[Modules.scala 160:64:@50756.4]
  assign _T_102612 = _T_102611[13:0]; // @[Modules.scala 160:64:@50757.4]
  assign buffer_15_397 = $signed(_T_102612); // @[Modules.scala 160:64:@50758.4]
  assign buffer_15_181 = {{8{_T_101461[5]}},_T_101461}; // @[Modules.scala 112:22:@8.4]
  assign _T_102614 = $signed(buffer_5_190) + $signed(buffer_15_181); // @[Modules.scala 160:64:@50760.4]
  assign _T_102615 = _T_102614[13:0]; // @[Modules.scala 160:64:@50761.4]
  assign buffer_15_398 = $signed(_T_102615); // @[Modules.scala 160:64:@50762.4]
  assign buffer_15_182 = {{8{_T_101468[5]}},_T_101468}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_183 = {{9{_T_101475[4]}},_T_101475}; // @[Modules.scala 112:22:@8.4]
  assign _T_102617 = $signed(buffer_15_182) + $signed(buffer_15_183); // @[Modules.scala 160:64:@50764.4]
  assign _T_102618 = _T_102617[13:0]; // @[Modules.scala 160:64:@50765.4]
  assign buffer_15_399 = $signed(_T_102618); // @[Modules.scala 160:64:@50766.4]
  assign buffer_15_184 = {{8{_T_101482[5]}},_T_101482}; // @[Modules.scala 112:22:@8.4]
  assign _T_102620 = $signed(buffer_15_184) + $signed(buffer_4_184); // @[Modules.scala 160:64:@50768.4]
  assign _T_102621 = _T_102620[13:0]; // @[Modules.scala 160:64:@50769.4]
  assign buffer_15_400 = $signed(_T_102621); // @[Modules.scala 160:64:@50770.4]
  assign _T_102626 = $signed(buffer_0_193) + $signed(buffer_0_194); // @[Modules.scala 160:64:@50776.4]
  assign _T_102627 = _T_102626[13:0]; // @[Modules.scala 160:64:@50777.4]
  assign buffer_15_402 = $signed(_T_102627); // @[Modules.scala 160:64:@50778.4]
  assign _T_102629 = $signed(buffer_13_198) + $signed(buffer_11_195); // @[Modules.scala 160:64:@50780.4]
  assign _T_102630 = _T_102629[13:0]; // @[Modules.scala 160:64:@50781.4]
  assign buffer_15_403 = $signed(_T_102630); // @[Modules.scala 160:64:@50782.4]
  assign buffer_15_192 = {{8{_T_101538[5]}},_T_101538}; // @[Modules.scala 112:22:@8.4]
  assign _T_102632 = $signed(buffer_15_192) + $signed(buffer_2_204); // @[Modules.scala 160:64:@50784.4]
  assign _T_102633 = _T_102632[13:0]; // @[Modules.scala 160:64:@50785.4]
  assign buffer_15_404 = $signed(_T_102633); // @[Modules.scala 160:64:@50786.4]
  assign buffer_15_196 = {{9{_T_101566[4]}},_T_101566}; // @[Modules.scala 112:22:@8.4]
  assign _T_102638 = $signed(buffer_15_196) + $signed(buffer_14_191); // @[Modules.scala 160:64:@50792.4]
  assign _T_102639 = _T_102638[13:0]; // @[Modules.scala 160:64:@50793.4]
  assign buffer_15_406 = $signed(_T_102639); // @[Modules.scala 160:64:@50794.4]
  assign buffer_15_205 = {{8{_T_101629[5]}},_T_101629}; // @[Modules.scala 112:22:@8.4]
  assign _T_102650 = $signed(buffer_1_208) + $signed(buffer_15_205); // @[Modules.scala 160:64:@50808.4]
  assign _T_102651 = _T_102650[13:0]; // @[Modules.scala 160:64:@50809.4]
  assign buffer_15_410 = $signed(_T_102651); // @[Modules.scala 160:64:@50810.4]
  assign _T_102659 = $signed(buffer_0_214) + $signed(buffer_5_217); // @[Modules.scala 160:64:@50820.4]
  assign _T_102660 = _T_102659[13:0]; // @[Modules.scala 160:64:@50821.4]
  assign buffer_15_413 = $signed(_T_102660); // @[Modules.scala 160:64:@50822.4]
  assign _T_102662 = $signed(buffer_9_224) + $signed(buffer_5_219); // @[Modules.scala 160:64:@50824.4]
  assign _T_102663 = _T_102662[13:0]; // @[Modules.scala 160:64:@50825.4]
  assign buffer_15_414 = $signed(_T_102663); // @[Modules.scala 160:64:@50826.4]
  assign buffer_15_215 = {{8{_T_101699[5]}},_T_101699}; // @[Modules.scala 112:22:@8.4]
  assign _T_102665 = $signed(buffer_5_220) + $signed(buffer_15_215); // @[Modules.scala 160:64:@50828.4]
  assign _T_102666 = _T_102665[13:0]; // @[Modules.scala 160:64:@50829.4]
  assign buffer_15_415 = $signed(_T_102666); // @[Modules.scala 160:64:@50830.4]
  assign buffer_15_216 = {{9{_T_101706[4]}},_T_101706}; // @[Modules.scala 112:22:@8.4]
  assign _T_102668 = $signed(buffer_15_216) + $signed(buffer_0_219); // @[Modules.scala 160:64:@50832.4]
  assign _T_102669 = _T_102668[13:0]; // @[Modules.scala 160:64:@50833.4]
  assign buffer_15_416 = $signed(_T_102669); // @[Modules.scala 160:64:@50834.4]
  assign _T_102671 = $signed(buffer_0_220) + $signed(buffer_8_226); // @[Modules.scala 160:64:@50836.4]
  assign _T_102672 = _T_102671[13:0]; // @[Modules.scala 160:64:@50837.4]
  assign buffer_15_417 = $signed(_T_102672); // @[Modules.scala 160:64:@50838.4]
  assign _T_102674 = $signed(buffer_12_215) + $signed(buffer_0_222); // @[Modules.scala 160:64:@50840.4]
  assign _T_102675 = _T_102674[13:0]; // @[Modules.scala 160:64:@50841.4]
  assign buffer_15_418 = $signed(_T_102675); // @[Modules.scala 160:64:@50842.4]
  assign buffer_15_223 = {{8{_T_101755[5]}},_T_101755}; // @[Modules.scala 112:22:@8.4]
  assign _T_102677 = $signed(buffer_0_223) + $signed(buffer_15_223); // @[Modules.scala 160:64:@50844.4]
  assign _T_102678 = _T_102677[13:0]; // @[Modules.scala 160:64:@50845.4]
  assign buffer_15_419 = $signed(_T_102678); // @[Modules.scala 160:64:@50846.4]
  assign buffer_15_224 = {{8{_T_101762[5]}},_T_101762}; // @[Modules.scala 112:22:@8.4]
  assign _T_102680 = $signed(buffer_15_224) + $signed(buffer_1_225); // @[Modules.scala 160:64:@50848.4]
  assign _T_102681 = _T_102680[13:0]; // @[Modules.scala 160:64:@50849.4]
  assign buffer_15_420 = $signed(_T_102681); // @[Modules.scala 160:64:@50850.4]
  assign _T_102683 = $signed(buffer_10_231) + $signed(buffer_13_228); // @[Modules.scala 160:64:@50852.4]
  assign _T_102684 = _T_102683[13:0]; // @[Modules.scala 160:64:@50853.4]
  assign buffer_15_421 = $signed(_T_102684); // @[Modules.scala 160:64:@50854.4]
  assign _T_102686 = $signed(buffer_1_228) + $signed(buffer_9_238); // @[Modules.scala 160:64:@50856.4]
  assign _T_102687 = _T_102686[13:0]; // @[Modules.scala 160:64:@50857.4]
  assign buffer_15_422 = $signed(_T_102687); // @[Modules.scala 160:64:@50858.4]
  assign buffer_15_231 = {{8{_T_101811[5]}},_T_101811}; // @[Modules.scala 112:22:@8.4]
  assign _T_102689 = $signed(buffer_6_241) + $signed(buffer_15_231); // @[Modules.scala 160:64:@50860.4]
  assign _T_102690 = _T_102689[13:0]; // @[Modules.scala 160:64:@50861.4]
  assign buffer_15_423 = $signed(_T_102690); // @[Modules.scala 160:64:@50862.4]
  assign buffer_15_237 = {{8{_T_101853[5]}},_T_101853}; // @[Modules.scala 112:22:@8.4]
  assign _T_102698 = $signed(buffer_2_240) + $signed(buffer_15_237); // @[Modules.scala 160:64:@50872.4]
  assign _T_102699 = _T_102698[13:0]; // @[Modules.scala 160:64:@50873.4]
  assign buffer_15_426 = $signed(_T_102699); // @[Modules.scala 160:64:@50874.4]
  assign _T_102701 = $signed(buffer_6_246) + $signed(buffer_5_244); // @[Modules.scala 160:64:@50876.4]
  assign _T_102702 = _T_102701[13:0]; // @[Modules.scala 160:64:@50877.4]
  assign buffer_15_427 = $signed(_T_102702); // @[Modules.scala 160:64:@50878.4]
  assign buffer_15_241 = {{8{_T_101881[5]}},_T_101881}; // @[Modules.scala 112:22:@8.4]
  assign _T_102704 = $signed(buffer_5_245) + $signed(buffer_15_241); // @[Modules.scala 160:64:@50880.4]
  assign _T_102705 = _T_102704[13:0]; // @[Modules.scala 160:64:@50881.4]
  assign buffer_15_428 = $signed(_T_102705); // @[Modules.scala 160:64:@50882.4]
  assign buffer_15_243 = {{9{_T_101895[4]}},_T_101895}; // @[Modules.scala 112:22:@8.4]
  assign _T_102707 = $signed(buffer_5_247) + $signed(buffer_15_243); // @[Modules.scala 160:64:@50884.4]
  assign _T_102708 = _T_102707[13:0]; // @[Modules.scala 160:64:@50885.4]
  assign buffer_15_429 = $signed(_T_102708); // @[Modules.scala 160:64:@50886.4]
  assign buffer_15_248 = {{8{_T_101930[5]}},_T_101930}; // @[Modules.scala 112:22:@8.4]
  assign buffer_15_249 = {{8{_T_101937[5]}},_T_101937}; // @[Modules.scala 112:22:@8.4]
  assign _T_102716 = $signed(buffer_15_248) + $signed(buffer_15_249); // @[Modules.scala 160:64:@50896.4]
  assign _T_102717 = _T_102716[13:0]; // @[Modules.scala 160:64:@50897.4]
  assign buffer_15_432 = $signed(_T_102717); // @[Modules.scala 160:64:@50898.4]
  assign _T_102719 = $signed(buffer_3_256) + $signed(buffer_6_258); // @[Modules.scala 160:64:@50900.4]
  assign _T_102720 = _T_102719[13:0]; // @[Modules.scala 160:64:@50901.4]
  assign buffer_15_433 = $signed(_T_102720); // @[Modules.scala 160:64:@50902.4]
  assign buffer_15_253 = {{8{_T_101965[5]}},_T_101965}; // @[Modules.scala 112:22:@8.4]
  assign _T_102722 = $signed(buffer_3_258) + $signed(buffer_15_253); // @[Modules.scala 160:64:@50904.4]
  assign _T_102723 = _T_102722[13:0]; // @[Modules.scala 160:64:@50905.4]
  assign buffer_15_434 = $signed(_T_102723); // @[Modules.scala 160:64:@50906.4]
  assign buffer_15_256 = {{8{_T_101986[5]}},_T_101986}; // @[Modules.scala 112:22:@8.4]
  assign _T_102728 = $signed(buffer_15_256) + $signed(buffer_5_262); // @[Modules.scala 160:64:@50912.4]
  assign _T_102729 = _T_102728[13:0]; // @[Modules.scala 160:64:@50913.4]
  assign buffer_15_436 = $signed(_T_102729); // @[Modules.scala 160:64:@50914.4]
  assign _T_102731 = $signed(buffer_3_263) + $signed(buffer_5_264); // @[Modules.scala 160:64:@50916.4]
  assign _T_102732 = _T_102731[13:0]; // @[Modules.scala 160:64:@50917.4]
  assign buffer_15_437 = $signed(_T_102732); // @[Modules.scala 160:64:@50918.4]
  assign buffer_15_260 = {{8{_T_102014[5]}},_T_102014}; // @[Modules.scala 112:22:@8.4]
  assign _T_102734 = $signed(buffer_15_260) + $signed(buffer_2_265); // @[Modules.scala 160:64:@50920.4]
  assign _T_102735 = _T_102734[13:0]; // @[Modules.scala 160:64:@50921.4]
  assign buffer_15_438 = $signed(_T_102735); // @[Modules.scala 160:64:@50922.4]
  assign _T_102737 = $signed(buffer_0_259) + $signed(buffer_6_271); // @[Modules.scala 160:64:@50924.4]
  assign _T_102738 = _T_102737[13:0]; // @[Modules.scala 160:64:@50925.4]
  assign buffer_15_439 = $signed(_T_102738); // @[Modules.scala 160:64:@50926.4]
  assign _T_102743 = $signed(buffer_4_258) + $signed(buffer_2_272); // @[Modules.scala 160:64:@50932.4]
  assign _T_102744 = _T_102743[13:0]; // @[Modules.scala 160:64:@50933.4]
  assign buffer_15_441 = $signed(_T_102744); // @[Modules.scala 160:64:@50934.4]
  assign _T_102752 = $signed(buffer_0_269) + $signed(buffer_0_270); // @[Modules.scala 160:64:@50944.4]
  assign _T_102753 = _T_102752[13:0]; // @[Modules.scala 160:64:@50945.4]
  assign buffer_15_444 = $signed(_T_102753); // @[Modules.scala 160:64:@50946.4]
  assign _T_102755 = $signed(buffer_0_271) + $signed(buffer_0_272); // @[Modules.scala 160:64:@50948.4]
  assign _T_102756 = _T_102755[13:0]; // @[Modules.scala 160:64:@50949.4]
  assign buffer_15_445 = $signed(_T_102756); // @[Modules.scala 160:64:@50950.4]
  assign _T_102758 = $signed(buffer_0_273) + $signed(buffer_10_278); // @[Modules.scala 160:64:@50952.4]
  assign _T_102759 = _T_102758[13:0]; // @[Modules.scala 160:64:@50953.4]
  assign buffer_15_446 = $signed(_T_102759); // @[Modules.scala 160:64:@50954.4]
  assign buffer_15_280 = {{8{_T_102154[5]}},_T_102154}; // @[Modules.scala 112:22:@8.4]
  assign _T_102764 = $signed(buffer_15_280) + $signed(buffer_12_273); // @[Modules.scala 160:64:@50960.4]
  assign _T_102765 = _T_102764[13:0]; // @[Modules.scala 160:64:@50961.4]
  assign buffer_15_448 = $signed(_T_102765); // @[Modules.scala 160:64:@50962.4]
  assign buffer_15_288 = {{9{_T_102210[4]}},_T_102210}; // @[Modules.scala 112:22:@8.4]
  assign _T_102776 = $signed(buffer_15_288) + $signed(buffer_11_281); // @[Modules.scala 160:64:@50976.4]
  assign _T_102777 = _T_102776[13:0]; // @[Modules.scala 160:64:@50977.4]
  assign buffer_15_452 = $signed(_T_102777); // @[Modules.scala 160:64:@50978.4]
  assign buffer_15_303 = {{8{_T_102315[5]}},_T_102315}; // @[Modules.scala 112:22:@8.4]
  assign _T_102797 = $signed(buffer_2_304) + $signed(buffer_15_303); // @[Modules.scala 160:64:@51004.4]
  assign _T_102798 = _T_102797[13:0]; // @[Modules.scala 160:64:@51005.4]
  assign buffer_15_459 = $signed(_T_102798); // @[Modules.scala 160:64:@51006.4]
  assign buffer_15_307 = {{8{_T_102343[5]}},_T_102343}; // @[Modules.scala 112:22:@8.4]
  assign _T_102803 = $signed(buffer_0_299) + $signed(buffer_15_307); // @[Modules.scala 160:64:@51012.4]
  assign _T_102804 = _T_102803[13:0]; // @[Modules.scala 160:64:@51013.4]
  assign buffer_15_461 = $signed(_T_102804); // @[Modules.scala 160:64:@51014.4]
  assign _T_102806 = $signed(buffer_15_308) + $signed(buffer_15_309); // @[Modules.scala 160:64:@51016.4]
  assign _T_102807 = _T_102806[13:0]; // @[Modules.scala 160:64:@51017.4]
  assign buffer_15_462 = $signed(_T_102807); // @[Modules.scala 160:64:@51018.4]
  assign _T_102815 = $signed(buffer_15_314) + $signed(buffer_14_309); // @[Modules.scala 160:64:@51028.4]
  assign _T_102816 = _T_102815[13:0]; // @[Modules.scala 160:64:@51029.4]
  assign buffer_15_465 = $signed(_T_102816); // @[Modules.scala 160:64:@51030.4]
  assign _T_102824 = $signed(buffer_15_320) + $signed(buffer_14_315); // @[Modules.scala 160:64:@51040.4]
  assign _T_102825 = _T_102824[13:0]; // @[Modules.scala 160:64:@51041.4]
  assign buffer_15_468 = $signed(_T_102825); // @[Modules.scala 160:64:@51042.4]
  assign _T_102830 = $signed(buffer_15_324) + $signed(buffer_15_325); // @[Modules.scala 160:64:@51048.4]
  assign _T_102831 = _T_102830[13:0]; // @[Modules.scala 160:64:@51049.4]
  assign buffer_15_470 = $signed(_T_102831); // @[Modules.scala 160:64:@51050.4]
  assign _T_102836 = $signed(buffer_10_328) + $signed(buffer_1_324); // @[Modules.scala 160:64:@51056.4]
  assign _T_102837 = _T_102836[13:0]; // @[Modules.scala 160:64:@51057.4]
  assign buffer_15_472 = $signed(_T_102837); // @[Modules.scala 160:64:@51058.4]
  assign _T_102839 = $signed(buffer_15_330) + $signed(buffer_15_331); // @[Modules.scala 160:64:@51060.4]
  assign _T_102840 = _T_102839[13:0]; // @[Modules.scala 160:64:@51061.4]
  assign buffer_15_473 = $signed(_T_102840); // @[Modules.scala 160:64:@51062.4]
  assign _T_102842 = $signed(buffer_15_332) + $signed(buffer_5_339); // @[Modules.scala 160:64:@51064.4]
  assign _T_102843 = _T_102842[13:0]; // @[Modules.scala 160:64:@51065.4]
  assign buffer_15_474 = $signed(_T_102843); // @[Modules.scala 160:64:@51066.4]
  assign _T_102845 = $signed(buffer_15_334) + $signed(buffer_15_335); // @[Modules.scala 160:64:@51068.4]
  assign _T_102846 = _T_102845[13:0]; // @[Modules.scala 160:64:@51069.4]
  assign buffer_15_475 = $signed(_T_102846); // @[Modules.scala 160:64:@51070.4]
  assign _T_102848 = $signed(buffer_15_336) + $signed(buffer_15_337); // @[Modules.scala 160:64:@51072.4]
  assign _T_102849 = _T_102848[13:0]; // @[Modules.scala 160:64:@51073.4]
  assign buffer_15_476 = $signed(_T_102849); // @[Modules.scala 160:64:@51074.4]
  assign _T_102851 = $signed(buffer_10_338) + $signed(buffer_15_339); // @[Modules.scala 160:64:@51076.4]
  assign _T_102852 = _T_102851[13:0]; // @[Modules.scala 160:64:@51077.4]
  assign buffer_15_477 = $signed(_T_102852); // @[Modules.scala 160:64:@51078.4]
  assign _T_102854 = $signed(buffer_15_340) + $signed(buffer_15_341); // @[Modules.scala 160:64:@51080.4]
  assign _T_102855 = _T_102854[13:0]; // @[Modules.scala 160:64:@51081.4]
  assign buffer_15_478 = $signed(_T_102855); // @[Modules.scala 160:64:@51082.4]
  assign _T_102857 = $signed(buffer_15_342) + $signed(buffer_15_343); // @[Modules.scala 160:64:@51084.4]
  assign _T_102858 = _T_102857[13:0]; // @[Modules.scala 160:64:@51085.4]
  assign buffer_15_479 = $signed(_T_102858); // @[Modules.scala 160:64:@51086.4]
  assign _T_102860 = $signed(buffer_15_344) + $signed(buffer_15_345); // @[Modules.scala 160:64:@51088.4]
  assign _T_102861 = _T_102860[13:0]; // @[Modules.scala 160:64:@51089.4]
  assign buffer_15_480 = $signed(_T_102861); // @[Modules.scala 160:64:@51090.4]
  assign _T_102863 = $signed(buffer_15_346) + $signed(buffer_15_347); // @[Modules.scala 160:64:@51092.4]
  assign _T_102864 = _T_102863[13:0]; // @[Modules.scala 160:64:@51093.4]
  assign buffer_15_481 = $signed(_T_102864); // @[Modules.scala 160:64:@51094.4]
  assign _T_102866 = $signed(buffer_15_348) + $signed(buffer_5_359); // @[Modules.scala 160:64:@51096.4]
  assign _T_102867 = _T_102866[13:0]; // @[Modules.scala 160:64:@51097.4]
  assign buffer_15_482 = $signed(_T_102867); // @[Modules.scala 160:64:@51098.4]
  assign _T_102869 = $signed(buffer_15_350) + $signed(buffer_15_351); // @[Modules.scala 160:64:@51100.4]
  assign _T_102870 = _T_102869[13:0]; // @[Modules.scala 160:64:@51101.4]
  assign buffer_15_483 = $signed(_T_102870); // @[Modules.scala 160:64:@51102.4]
  assign _T_102872 = $signed(buffer_15_352) + $signed(buffer_15_353); // @[Modules.scala 160:64:@51104.4]
  assign _T_102873 = _T_102872[13:0]; // @[Modules.scala 160:64:@51105.4]
  assign buffer_15_484 = $signed(_T_102873); // @[Modules.scala 160:64:@51106.4]
  assign _T_102875 = $signed(buffer_5_366) + $signed(buffer_15_355); // @[Modules.scala 160:64:@51108.4]
  assign _T_102876 = _T_102875[13:0]; // @[Modules.scala 160:64:@51109.4]
  assign buffer_15_485 = $signed(_T_102876); // @[Modules.scala 160:64:@51110.4]
  assign _T_102878 = $signed(buffer_15_356) + $signed(buffer_15_357); // @[Modules.scala 160:64:@51112.4]
  assign _T_102879 = _T_102878[13:0]; // @[Modules.scala 160:64:@51113.4]
  assign buffer_15_486 = $signed(_T_102879); // @[Modules.scala 160:64:@51114.4]
  assign _T_102881 = $signed(buffer_15_358) + $signed(buffer_15_359); // @[Modules.scala 160:64:@51116.4]
  assign _T_102882 = _T_102881[13:0]; // @[Modules.scala 160:64:@51117.4]
  assign buffer_15_487 = $signed(_T_102882); // @[Modules.scala 160:64:@51118.4]
  assign _T_102884 = $signed(buffer_15_360) + $signed(buffer_15_361); // @[Modules.scala 160:64:@51120.4]
  assign _T_102885 = _T_102884[13:0]; // @[Modules.scala 160:64:@51121.4]
  assign buffer_15_488 = $signed(_T_102885); // @[Modules.scala 160:64:@51122.4]
  assign _T_102887 = $signed(buffer_15_362) + $signed(buffer_15_363); // @[Modules.scala 160:64:@51124.4]
  assign _T_102888 = _T_102887[13:0]; // @[Modules.scala 160:64:@51125.4]
  assign buffer_15_489 = $signed(_T_102888); // @[Modules.scala 160:64:@51126.4]
  assign _T_102890 = $signed(buffer_0_362) + $signed(buffer_15_365); // @[Modules.scala 160:64:@51128.4]
  assign _T_102891 = _T_102890[13:0]; // @[Modules.scala 160:64:@51129.4]
  assign buffer_15_490 = $signed(_T_102891); // @[Modules.scala 160:64:@51130.4]
  assign _T_102893 = $signed(buffer_15_366) + $signed(buffer_15_367); // @[Modules.scala 160:64:@51132.4]
  assign _T_102894 = _T_102893[13:0]; // @[Modules.scala 160:64:@51133.4]
  assign buffer_15_491 = $signed(_T_102894); // @[Modules.scala 160:64:@51134.4]
  assign _T_102896 = $signed(buffer_15_368) + $signed(buffer_15_369); // @[Modules.scala 160:64:@51136.4]
  assign _T_102897 = _T_102896[13:0]; // @[Modules.scala 160:64:@51137.4]
  assign buffer_15_492 = $signed(_T_102897); // @[Modules.scala 160:64:@51138.4]
  assign _T_102899 = $signed(buffer_15_370) + $signed(buffer_15_371); // @[Modules.scala 160:64:@51140.4]
  assign _T_102900 = _T_102899[13:0]; // @[Modules.scala 160:64:@51141.4]
  assign buffer_15_493 = $signed(_T_102900); // @[Modules.scala 160:64:@51142.4]
  assign _T_102902 = $signed(buffer_11_365) + $signed(buffer_13_376); // @[Modules.scala 160:64:@51144.4]
  assign _T_102903 = _T_102902[13:0]; // @[Modules.scala 160:64:@51145.4]
  assign buffer_15_494 = $signed(_T_102903); // @[Modules.scala 160:64:@51146.4]
  assign _T_102905 = $signed(buffer_15_374) + $signed(buffer_15_375); // @[Modules.scala 160:64:@51148.4]
  assign _T_102906 = _T_102905[13:0]; // @[Modules.scala 160:64:@51149.4]
  assign buffer_15_495 = $signed(_T_102906); // @[Modules.scala 160:64:@51150.4]
  assign _T_102908 = $signed(buffer_15_376) + $signed(buffer_15_377); // @[Modules.scala 160:64:@51152.4]
  assign _T_102909 = _T_102908[13:0]; // @[Modules.scala 160:64:@51153.4]
  assign buffer_15_496 = $signed(_T_102909); // @[Modules.scala 160:64:@51154.4]
  assign _T_102911 = $signed(buffer_15_378) + $signed(buffer_5_390); // @[Modules.scala 160:64:@51156.4]
  assign _T_102912 = _T_102911[13:0]; // @[Modules.scala 160:64:@51157.4]
  assign buffer_15_497 = $signed(_T_102912); // @[Modules.scala 160:64:@51158.4]
  assign _T_102914 = $signed(buffer_15_380) + $signed(buffer_15_381); // @[Modules.scala 160:64:@51160.4]
  assign _T_102915 = _T_102914[13:0]; // @[Modules.scala 160:64:@51161.4]
  assign buffer_15_498 = $signed(_T_102915); // @[Modules.scala 160:64:@51162.4]
  assign _T_102917 = $signed(buffer_15_382) + $signed(buffer_15_383); // @[Modules.scala 160:64:@51164.4]
  assign _T_102918 = _T_102917[13:0]; // @[Modules.scala 160:64:@51165.4]
  assign buffer_15_499 = $signed(_T_102918); // @[Modules.scala 160:64:@51166.4]
  assign _T_102920 = $signed(buffer_15_384) + $signed(buffer_12_374); // @[Modules.scala 160:64:@51168.4]
  assign _T_102921 = _T_102920[13:0]; // @[Modules.scala 160:64:@51169.4]
  assign buffer_15_500 = $signed(_T_102921); // @[Modules.scala 160:64:@51170.4]
  assign _T_102923 = $signed(buffer_15_386) + $signed(buffer_7_394); // @[Modules.scala 160:64:@51172.4]
  assign _T_102924 = _T_102923[13:0]; // @[Modules.scala 160:64:@51173.4]
  assign buffer_15_501 = $signed(_T_102924); // @[Modules.scala 160:64:@51174.4]
  assign _T_102926 = $signed(buffer_7_395) + $signed(buffer_15_389); // @[Modules.scala 160:64:@51176.4]
  assign _T_102927 = _T_102926[13:0]; // @[Modules.scala 160:64:@51177.4]
  assign buffer_15_502 = $signed(_T_102927); // @[Modules.scala 160:64:@51178.4]
  assign _T_102929 = $signed(buffer_15_390) + $signed(buffer_15_391); // @[Modules.scala 160:64:@51180.4]
  assign _T_102930 = _T_102929[13:0]; // @[Modules.scala 160:64:@51181.4]
  assign buffer_15_503 = $signed(_T_102930); // @[Modules.scala 160:64:@51182.4]
  assign _T_102932 = $signed(buffer_15_392) + $signed(buffer_15_393); // @[Modules.scala 160:64:@51184.4]
  assign _T_102933 = _T_102932[13:0]; // @[Modules.scala 160:64:@51185.4]
  assign buffer_15_504 = $signed(_T_102933); // @[Modules.scala 160:64:@51186.4]
  assign _T_102935 = $signed(buffer_15_394) + $signed(buffer_15_395); // @[Modules.scala 160:64:@51188.4]
  assign _T_102936 = _T_102935[13:0]; // @[Modules.scala 160:64:@51189.4]
  assign buffer_15_505 = $signed(_T_102936); // @[Modules.scala 160:64:@51190.4]
  assign _T_102938 = $signed(buffer_6_411) + $signed(buffer_15_397); // @[Modules.scala 160:64:@51192.4]
  assign _T_102939 = _T_102938[13:0]; // @[Modules.scala 160:64:@51193.4]
  assign buffer_15_506 = $signed(_T_102939); // @[Modules.scala 160:64:@51194.4]
  assign _T_102941 = $signed(buffer_15_398) + $signed(buffer_15_399); // @[Modules.scala 160:64:@51196.4]
  assign _T_102942 = _T_102941[13:0]; // @[Modules.scala 160:64:@51197.4]
  assign buffer_15_507 = $signed(_T_102942); // @[Modules.scala 160:64:@51198.4]
  assign _T_102944 = $signed(buffer_15_400) + $signed(buffer_6_417); // @[Modules.scala 160:64:@51200.4]
  assign _T_102945 = _T_102944[13:0]; // @[Modules.scala 160:64:@51201.4]
  assign buffer_15_508 = $signed(_T_102945); // @[Modules.scala 160:64:@51202.4]
  assign _T_102947 = $signed(buffer_15_402) + $signed(buffer_15_403); // @[Modules.scala 160:64:@51204.4]
  assign _T_102948 = _T_102947[13:0]; // @[Modules.scala 160:64:@51205.4]
  assign buffer_15_509 = $signed(_T_102948); // @[Modules.scala 160:64:@51206.4]
  assign _T_102950 = $signed(buffer_15_404) + $signed(buffer_10_411); // @[Modules.scala 160:64:@51208.4]
  assign _T_102951 = _T_102950[13:0]; // @[Modules.scala 160:64:@51209.4]
  assign buffer_15_510 = $signed(_T_102951); // @[Modules.scala 160:64:@51210.4]
  assign _T_102953 = $signed(buffer_15_406) + $signed(buffer_14_398); // @[Modules.scala 160:64:@51212.4]
  assign _T_102954 = _T_102953[13:0]; // @[Modules.scala 160:64:@51213.4]
  assign buffer_15_511 = $signed(_T_102954); // @[Modules.scala 160:64:@51214.4]
  assign _T_102956 = $signed(buffer_5_418) + $signed(buffer_10_414); // @[Modules.scala 160:64:@51216.4]
  assign _T_102957 = _T_102956[13:0]; // @[Modules.scala 160:64:@51217.4]
  assign buffer_15_512 = $signed(_T_102957); // @[Modules.scala 160:64:@51218.4]
  assign _T_102959 = $signed(buffer_15_410) + $signed(buffer_0_407); // @[Modules.scala 160:64:@51220.4]
  assign _T_102960 = _T_102959[13:0]; // @[Modules.scala 160:64:@51221.4]
  assign buffer_15_513 = $signed(_T_102960); // @[Modules.scala 160:64:@51222.4]
  assign _T_102962 = $signed(buffer_0_408) + $signed(buffer_15_413); // @[Modules.scala 160:64:@51224.4]
  assign _T_102963 = _T_102962[13:0]; // @[Modules.scala 160:64:@51225.4]
  assign buffer_15_514 = $signed(_T_102963); // @[Modules.scala 160:64:@51226.4]
  assign _T_102965 = $signed(buffer_15_414) + $signed(buffer_15_415); // @[Modules.scala 160:64:@51228.4]
  assign _T_102966 = _T_102965[13:0]; // @[Modules.scala 160:64:@51229.4]
  assign buffer_15_515 = $signed(_T_102966); // @[Modules.scala 160:64:@51230.4]
  assign _T_102968 = $signed(buffer_15_416) + $signed(buffer_15_417); // @[Modules.scala 160:64:@51232.4]
  assign _T_102969 = _T_102968[13:0]; // @[Modules.scala 160:64:@51233.4]
  assign buffer_15_516 = $signed(_T_102969); // @[Modules.scala 160:64:@51234.4]
  assign _T_102971 = $signed(buffer_15_418) + $signed(buffer_15_419); // @[Modules.scala 160:64:@51236.4]
  assign _T_102972 = _T_102971[13:0]; // @[Modules.scala 160:64:@51237.4]
  assign buffer_15_517 = $signed(_T_102972); // @[Modules.scala 160:64:@51238.4]
  assign _T_102974 = $signed(buffer_15_420) + $signed(buffer_15_421); // @[Modules.scala 160:64:@51240.4]
  assign _T_102975 = _T_102974[13:0]; // @[Modules.scala 160:64:@51241.4]
  assign buffer_15_518 = $signed(_T_102975); // @[Modules.scala 160:64:@51242.4]
  assign _T_102977 = $signed(buffer_15_422) + $signed(buffer_15_423); // @[Modules.scala 160:64:@51244.4]
  assign _T_102978 = _T_102977[13:0]; // @[Modules.scala 160:64:@51245.4]
  assign buffer_15_519 = $signed(_T_102978); // @[Modules.scala 160:64:@51246.4]
  assign _T_102980 = $signed(buffer_12_411) + $signed(buffer_12_412); // @[Modules.scala 160:64:@51248.4]
  assign _T_102981 = _T_102980[13:0]; // @[Modules.scala 160:64:@51249.4]
  assign buffer_15_520 = $signed(_T_102981); // @[Modules.scala 160:64:@51250.4]
  assign _T_102983 = $signed(buffer_15_426) + $signed(buffer_15_427); // @[Modules.scala 160:64:@51252.4]
  assign _T_102984 = _T_102983[13:0]; // @[Modules.scala 160:64:@51253.4]
  assign buffer_15_521 = $signed(_T_102984); // @[Modules.scala 160:64:@51254.4]
  assign _T_102986 = $signed(buffer_15_428) + $signed(buffer_15_429); // @[Modules.scala 160:64:@51256.4]
  assign _T_102987 = _T_102986[13:0]; // @[Modules.scala 160:64:@51257.4]
  assign buffer_15_522 = $signed(_T_102987); // @[Modules.scala 160:64:@51258.4]
  assign _T_102989 = $signed(buffer_1_424) + $signed(buffer_14_420); // @[Modules.scala 160:64:@51260.4]
  assign _T_102990 = _T_102989[13:0]; // @[Modules.scala 160:64:@51261.4]
  assign buffer_15_523 = $signed(_T_102990); // @[Modules.scala 160:64:@51262.4]
  assign _T_102992 = $signed(buffer_15_432) + $signed(buffer_15_433); // @[Modules.scala 160:64:@51264.4]
  assign _T_102993 = _T_102992[13:0]; // @[Modules.scala 160:64:@51265.4]
  assign buffer_15_524 = $signed(_T_102993); // @[Modules.scala 160:64:@51266.4]
  assign _T_102995 = $signed(buffer_15_434) + $signed(buffer_0_427); // @[Modules.scala 160:64:@51268.4]
  assign _T_102996 = _T_102995[13:0]; // @[Modules.scala 160:64:@51269.4]
  assign buffer_15_525 = $signed(_T_102996); // @[Modules.scala 160:64:@51270.4]
  assign _T_102998 = $signed(buffer_15_436) + $signed(buffer_15_437); // @[Modules.scala 160:64:@51272.4]
  assign _T_102999 = _T_102998[13:0]; // @[Modules.scala 160:64:@51273.4]
  assign buffer_15_526 = $signed(_T_102999); // @[Modules.scala 160:64:@51274.4]
  assign _T_103001 = $signed(buffer_15_438) + $signed(buffer_15_439); // @[Modules.scala 160:64:@51276.4]
  assign _T_103002 = _T_103001[13:0]; // @[Modules.scala 160:64:@51277.4]
  assign buffer_15_527 = $signed(_T_103002); // @[Modules.scala 160:64:@51278.4]
  assign _T_103004 = $signed(buffer_1_434) + $signed(buffer_15_441); // @[Modules.scala 160:64:@51280.4]
  assign _T_103005 = _T_103004[13:0]; // @[Modules.scala 160:64:@51281.4]
  assign buffer_15_528 = $signed(_T_103005); // @[Modules.scala 160:64:@51282.4]
  assign _T_103007 = $signed(buffer_5_451) + $signed(buffer_5_452); // @[Modules.scala 160:64:@51284.4]
  assign _T_103008 = _T_103007[13:0]; // @[Modules.scala 160:64:@51285.4]
  assign buffer_15_529 = $signed(_T_103008); // @[Modules.scala 160:64:@51286.4]
  assign _T_103010 = $signed(buffer_15_444) + $signed(buffer_15_445); // @[Modules.scala 160:64:@51288.4]
  assign _T_103011 = _T_103010[13:0]; // @[Modules.scala 160:64:@51289.4]
  assign buffer_15_530 = $signed(_T_103011); // @[Modules.scala 160:64:@51290.4]
  assign _T_103013 = $signed(buffer_15_446) + $signed(buffer_3_456); // @[Modules.scala 160:64:@51292.4]
  assign _T_103014 = _T_103013[13:0]; // @[Modules.scala 160:64:@51293.4]
  assign buffer_15_531 = $signed(_T_103014); // @[Modules.scala 160:64:@51294.4]
  assign _T_103016 = $signed(buffer_15_448) + $signed(buffer_12_435); // @[Modules.scala 160:64:@51296.4]
  assign _T_103017 = _T_103016[13:0]; // @[Modules.scala 160:64:@51297.4]
  assign buffer_15_532 = $signed(_T_103017); // @[Modules.scala 160:64:@51298.4]
  assign _T_103022 = $signed(buffer_15_452) + $signed(buffer_9_462); // @[Modules.scala 160:64:@51304.4]
  assign _T_103023 = _T_103022[13:0]; // @[Modules.scala 160:64:@51305.4]
  assign buffer_15_534 = $signed(_T_103023); // @[Modules.scala 160:64:@51306.4]
  assign _T_103025 = $signed(buffer_9_463) + $signed(buffer_9_464); // @[Modules.scala 160:64:@51308.4]
  assign _T_103026 = _T_103025[13:0]; // @[Modules.scala 160:64:@51309.4]
  assign buffer_15_535 = $signed(_T_103026); // @[Modules.scala 160:64:@51310.4]
  assign _T_103031 = $signed(buffer_6_470) + $signed(buffer_15_459); // @[Modules.scala 160:64:@51316.4]
  assign _T_103032 = _T_103031[13:0]; // @[Modules.scala 160:64:@51317.4]
  assign buffer_15_537 = $signed(_T_103032); // @[Modules.scala 160:64:@51318.4]
  assign _T_103034 = $signed(buffer_9_469) + $signed(buffer_15_461); // @[Modules.scala 160:64:@51320.4]
  assign _T_103035 = _T_103034[13:0]; // @[Modules.scala 160:64:@51321.4]
  assign buffer_15_538 = $signed(_T_103035); // @[Modules.scala 160:64:@51322.4]
  assign _T_103037 = $signed(buffer_15_462) + $signed(buffer_0_454); // @[Modules.scala 166:64:@51324.4]
  assign _T_103038 = _T_103037[13:0]; // @[Modules.scala 166:64:@51325.4]
  assign buffer_15_539 = $signed(_T_103038); // @[Modules.scala 166:64:@51326.4]
  assign _T_103040 = $signed(buffer_0_455) + $signed(buffer_15_465); // @[Modules.scala 166:64:@51328.4]
  assign _T_103041 = _T_103040[13:0]; // @[Modules.scala 166:64:@51329.4]
  assign buffer_15_540 = $signed(_T_103041); // @[Modules.scala 166:64:@51330.4]
  assign _T_103046 = $signed(buffer_15_468) + $signed(buffer_14_460); // @[Modules.scala 166:64:@51336.4]
  assign _T_103047 = _T_103046[13:0]; // @[Modules.scala 166:64:@51337.4]
  assign buffer_15_542 = $signed(_T_103047); // @[Modules.scala 166:64:@51338.4]
  assign _T_103049 = $signed(buffer_15_470) + $signed(buffer_10_471); // @[Modules.scala 166:64:@51340.4]
  assign _T_103050 = _T_103049[13:0]; // @[Modules.scala 166:64:@51341.4]
  assign buffer_15_543 = $signed(_T_103050); // @[Modules.scala 166:64:@51342.4]
  assign _T_103052 = $signed(buffer_15_472) + $signed(buffer_15_473); // @[Modules.scala 166:64:@51344.4]
  assign _T_103053 = _T_103052[13:0]; // @[Modules.scala 166:64:@51345.4]
  assign buffer_15_544 = $signed(_T_103053); // @[Modules.scala 166:64:@51346.4]
  assign _T_103055 = $signed(buffer_15_474) + $signed(buffer_15_475); // @[Modules.scala 166:64:@51348.4]
  assign _T_103056 = _T_103055[13:0]; // @[Modules.scala 166:64:@51349.4]
  assign buffer_15_545 = $signed(_T_103056); // @[Modules.scala 166:64:@51350.4]
  assign _T_103058 = $signed(buffer_15_476) + $signed(buffer_15_477); // @[Modules.scala 166:64:@51352.4]
  assign _T_103059 = _T_103058[13:0]; // @[Modules.scala 166:64:@51353.4]
  assign buffer_15_546 = $signed(_T_103059); // @[Modules.scala 166:64:@51354.4]
  assign _T_103061 = $signed(buffer_15_478) + $signed(buffer_15_479); // @[Modules.scala 166:64:@51356.4]
  assign _T_103062 = _T_103061[13:0]; // @[Modules.scala 166:64:@51357.4]
  assign buffer_15_547 = $signed(_T_103062); // @[Modules.scala 166:64:@51358.4]
  assign _T_103064 = $signed(buffer_15_480) + $signed(buffer_15_481); // @[Modules.scala 166:64:@51360.4]
  assign _T_103065 = _T_103064[13:0]; // @[Modules.scala 166:64:@51361.4]
  assign buffer_15_548 = $signed(_T_103065); // @[Modules.scala 166:64:@51362.4]
  assign _T_103067 = $signed(buffer_15_482) + $signed(buffer_15_483); // @[Modules.scala 166:64:@51364.4]
  assign _T_103068 = _T_103067[13:0]; // @[Modules.scala 166:64:@51365.4]
  assign buffer_15_549 = $signed(_T_103068); // @[Modules.scala 166:64:@51366.4]
  assign _T_103070 = $signed(buffer_15_484) + $signed(buffer_15_485); // @[Modules.scala 166:64:@51368.4]
  assign _T_103071 = _T_103070[13:0]; // @[Modules.scala 166:64:@51369.4]
  assign buffer_15_550 = $signed(_T_103071); // @[Modules.scala 166:64:@51370.4]
  assign _T_103073 = $signed(buffer_15_486) + $signed(buffer_15_487); // @[Modules.scala 166:64:@51372.4]
  assign _T_103074 = _T_103073[13:0]; // @[Modules.scala 166:64:@51373.4]
  assign buffer_15_551 = $signed(_T_103074); // @[Modules.scala 166:64:@51374.4]
  assign _T_103076 = $signed(buffer_15_488) + $signed(buffer_15_489); // @[Modules.scala 166:64:@51376.4]
  assign _T_103077 = _T_103076[13:0]; // @[Modules.scala 166:64:@51377.4]
  assign buffer_15_552 = $signed(_T_103077); // @[Modules.scala 166:64:@51378.4]
  assign _T_103079 = $signed(buffer_15_490) + $signed(buffer_15_491); // @[Modules.scala 166:64:@51380.4]
  assign _T_103080 = _T_103079[13:0]; // @[Modules.scala 166:64:@51381.4]
  assign buffer_15_553 = $signed(_T_103080); // @[Modules.scala 166:64:@51382.4]
  assign _T_103082 = $signed(buffer_15_492) + $signed(buffer_15_493); // @[Modules.scala 166:64:@51384.4]
  assign _T_103083 = _T_103082[13:0]; // @[Modules.scala 166:64:@51385.4]
  assign buffer_15_554 = $signed(_T_103083); // @[Modules.scala 166:64:@51386.4]
  assign _T_103085 = $signed(buffer_15_494) + $signed(buffer_15_495); // @[Modules.scala 166:64:@51388.4]
  assign _T_103086 = _T_103085[13:0]; // @[Modules.scala 166:64:@51389.4]
  assign buffer_15_555 = $signed(_T_103086); // @[Modules.scala 166:64:@51390.4]
  assign _T_103088 = $signed(buffer_15_496) + $signed(buffer_15_497); // @[Modules.scala 166:64:@51392.4]
  assign _T_103089 = _T_103088[13:0]; // @[Modules.scala 166:64:@51393.4]
  assign buffer_15_556 = $signed(_T_103089); // @[Modules.scala 166:64:@51394.4]
  assign _T_103091 = $signed(buffer_15_498) + $signed(buffer_15_499); // @[Modules.scala 166:64:@51396.4]
  assign _T_103092 = _T_103091[13:0]; // @[Modules.scala 166:64:@51397.4]
  assign buffer_15_557 = $signed(_T_103092); // @[Modules.scala 166:64:@51398.4]
  assign _T_103094 = $signed(buffer_15_500) + $signed(buffer_15_501); // @[Modules.scala 166:64:@51400.4]
  assign _T_103095 = _T_103094[13:0]; // @[Modules.scala 166:64:@51401.4]
  assign buffer_15_558 = $signed(_T_103095); // @[Modules.scala 166:64:@51402.4]
  assign _T_103097 = $signed(buffer_15_502) + $signed(buffer_15_503); // @[Modules.scala 166:64:@51404.4]
  assign _T_103098 = _T_103097[13:0]; // @[Modules.scala 166:64:@51405.4]
  assign buffer_15_559 = $signed(_T_103098); // @[Modules.scala 166:64:@51406.4]
  assign _T_103100 = $signed(buffer_15_504) + $signed(buffer_15_505); // @[Modules.scala 166:64:@51408.4]
  assign _T_103101 = _T_103100[13:0]; // @[Modules.scala 166:64:@51409.4]
  assign buffer_15_560 = $signed(_T_103101); // @[Modules.scala 166:64:@51410.4]
  assign _T_103103 = $signed(buffer_15_506) + $signed(buffer_15_507); // @[Modules.scala 166:64:@51412.4]
  assign _T_103104 = _T_103103[13:0]; // @[Modules.scala 166:64:@51413.4]
  assign buffer_15_561 = $signed(_T_103104); // @[Modules.scala 166:64:@51414.4]
  assign _T_103106 = $signed(buffer_15_508) + $signed(buffer_15_509); // @[Modules.scala 166:64:@51416.4]
  assign _T_103107 = _T_103106[13:0]; // @[Modules.scala 166:64:@51417.4]
  assign buffer_15_562 = $signed(_T_103107); // @[Modules.scala 166:64:@51418.4]
  assign _T_103109 = $signed(buffer_15_510) + $signed(buffer_15_511); // @[Modules.scala 166:64:@51420.4]
  assign _T_103110 = _T_103109[13:0]; // @[Modules.scala 166:64:@51421.4]
  assign buffer_15_563 = $signed(_T_103110); // @[Modules.scala 166:64:@51422.4]
  assign _T_103112 = $signed(buffer_15_512) + $signed(buffer_15_513); // @[Modules.scala 166:64:@51424.4]
  assign _T_103113 = _T_103112[13:0]; // @[Modules.scala 166:64:@51425.4]
  assign buffer_15_564 = $signed(_T_103113); // @[Modules.scala 166:64:@51426.4]
  assign _T_103115 = $signed(buffer_15_514) + $signed(buffer_15_515); // @[Modules.scala 166:64:@51428.4]
  assign _T_103116 = _T_103115[13:0]; // @[Modules.scala 166:64:@51429.4]
  assign buffer_15_565 = $signed(_T_103116); // @[Modules.scala 166:64:@51430.4]
  assign _T_103118 = $signed(buffer_15_516) + $signed(buffer_15_517); // @[Modules.scala 166:64:@51432.4]
  assign _T_103119 = _T_103118[13:0]; // @[Modules.scala 166:64:@51433.4]
  assign buffer_15_566 = $signed(_T_103119); // @[Modules.scala 166:64:@51434.4]
  assign _T_103121 = $signed(buffer_15_518) + $signed(buffer_15_519); // @[Modules.scala 166:64:@51436.4]
  assign _T_103122 = _T_103121[13:0]; // @[Modules.scala 166:64:@51437.4]
  assign buffer_15_567 = $signed(_T_103122); // @[Modules.scala 166:64:@51438.4]
  assign _T_103124 = $signed(buffer_15_520) + $signed(buffer_15_521); // @[Modules.scala 166:64:@51440.4]
  assign _T_103125 = _T_103124[13:0]; // @[Modules.scala 166:64:@51441.4]
  assign buffer_15_568 = $signed(_T_103125); // @[Modules.scala 166:64:@51442.4]
  assign _T_103127 = $signed(buffer_15_522) + $signed(buffer_15_523); // @[Modules.scala 166:64:@51444.4]
  assign _T_103128 = _T_103127[13:0]; // @[Modules.scala 166:64:@51445.4]
  assign buffer_15_569 = $signed(_T_103128); // @[Modules.scala 166:64:@51446.4]
  assign _T_103130 = $signed(buffer_15_524) + $signed(buffer_15_525); // @[Modules.scala 166:64:@51448.4]
  assign _T_103131 = _T_103130[13:0]; // @[Modules.scala 166:64:@51449.4]
  assign buffer_15_570 = $signed(_T_103131); // @[Modules.scala 166:64:@51450.4]
  assign _T_103133 = $signed(buffer_15_526) + $signed(buffer_15_527); // @[Modules.scala 166:64:@51452.4]
  assign _T_103134 = _T_103133[13:0]; // @[Modules.scala 166:64:@51453.4]
  assign buffer_15_571 = $signed(_T_103134); // @[Modules.scala 166:64:@51454.4]
  assign _T_103136 = $signed(buffer_15_528) + $signed(buffer_15_529); // @[Modules.scala 166:64:@51456.4]
  assign _T_103137 = _T_103136[13:0]; // @[Modules.scala 166:64:@51457.4]
  assign buffer_15_572 = $signed(_T_103137); // @[Modules.scala 166:64:@51458.4]
  assign _T_103139 = $signed(buffer_15_530) + $signed(buffer_15_531); // @[Modules.scala 166:64:@51460.4]
  assign _T_103140 = _T_103139[13:0]; // @[Modules.scala 166:64:@51461.4]
  assign buffer_15_573 = $signed(_T_103140); // @[Modules.scala 166:64:@51462.4]
  assign _T_103142 = $signed(buffer_15_532) + $signed(buffer_6_547); // @[Modules.scala 166:64:@51464.4]
  assign _T_103143 = _T_103142[13:0]; // @[Modules.scala 166:64:@51465.4]
  assign buffer_15_574 = $signed(_T_103143); // @[Modules.scala 166:64:@51466.4]
  assign _T_103145 = $signed(buffer_15_534) + $signed(buffer_15_535); // @[Modules.scala 166:64:@51468.4]
  assign _T_103146 = _T_103145[13:0]; // @[Modules.scala 166:64:@51469.4]
  assign buffer_15_575 = $signed(_T_103146); // @[Modules.scala 166:64:@51470.4]
  assign _T_103148 = $signed(buffer_6_550) + $signed(buffer_15_537); // @[Modules.scala 166:64:@51472.4]
  assign _T_103149 = _T_103148[13:0]; // @[Modules.scala 166:64:@51473.4]
  assign buffer_15_576 = $signed(_T_103149); // @[Modules.scala 166:64:@51474.4]
  assign _T_103151 = $signed(buffer_15_539) + $signed(buffer_15_540); // @[Modules.scala 160:64:@51476.4]
  assign _T_103152 = _T_103151[13:0]; // @[Modules.scala 160:64:@51477.4]
  assign buffer_15_577 = $signed(_T_103152); // @[Modules.scala 160:64:@51478.4]
  assign _T_103154 = $signed(buffer_14_530) + $signed(buffer_15_542); // @[Modules.scala 160:64:@51480.4]
  assign _T_103155 = _T_103154[13:0]; // @[Modules.scala 160:64:@51481.4]
  assign buffer_15_578 = $signed(_T_103155); // @[Modules.scala 160:64:@51482.4]
  assign _T_103157 = $signed(buffer_15_543) + $signed(buffer_15_544); // @[Modules.scala 160:64:@51484.4]
  assign _T_103158 = _T_103157[13:0]; // @[Modules.scala 160:64:@51485.4]
  assign buffer_15_579 = $signed(_T_103158); // @[Modules.scala 160:64:@51486.4]
  assign _T_103160 = $signed(buffer_15_545) + $signed(buffer_15_546); // @[Modules.scala 160:64:@51488.4]
  assign _T_103161 = _T_103160[13:0]; // @[Modules.scala 160:64:@51489.4]
  assign buffer_15_580 = $signed(_T_103161); // @[Modules.scala 160:64:@51490.4]
  assign _T_103163 = $signed(buffer_15_547) + $signed(buffer_15_548); // @[Modules.scala 160:64:@51492.4]
  assign _T_103164 = _T_103163[13:0]; // @[Modules.scala 160:64:@51493.4]
  assign buffer_15_581 = $signed(_T_103164); // @[Modules.scala 160:64:@51494.4]
  assign _T_103166 = $signed(buffer_15_549) + $signed(buffer_15_550); // @[Modules.scala 160:64:@51496.4]
  assign _T_103167 = _T_103166[13:0]; // @[Modules.scala 160:64:@51497.4]
  assign buffer_15_582 = $signed(_T_103167); // @[Modules.scala 160:64:@51498.4]
  assign _T_103169 = $signed(buffer_15_551) + $signed(buffer_15_552); // @[Modules.scala 160:64:@51500.4]
  assign _T_103170 = _T_103169[13:0]; // @[Modules.scala 160:64:@51501.4]
  assign buffer_15_583 = $signed(_T_103170); // @[Modules.scala 160:64:@51502.4]
  assign _T_103172 = $signed(buffer_15_553) + $signed(buffer_15_554); // @[Modules.scala 160:64:@51504.4]
  assign _T_103173 = _T_103172[13:0]; // @[Modules.scala 160:64:@51505.4]
  assign buffer_15_584 = $signed(_T_103173); // @[Modules.scala 160:64:@51506.4]
  assign _T_103175 = $signed(buffer_15_555) + $signed(buffer_15_556); // @[Modules.scala 160:64:@51508.4]
  assign _T_103176 = _T_103175[13:0]; // @[Modules.scala 160:64:@51509.4]
  assign buffer_15_585 = $signed(_T_103176); // @[Modules.scala 160:64:@51510.4]
  assign _T_103178 = $signed(buffer_15_557) + $signed(buffer_15_558); // @[Modules.scala 160:64:@51512.4]
  assign _T_103179 = _T_103178[13:0]; // @[Modules.scala 160:64:@51513.4]
  assign buffer_15_586 = $signed(_T_103179); // @[Modules.scala 160:64:@51514.4]
  assign _T_103181 = $signed(buffer_15_559) + $signed(buffer_15_560); // @[Modules.scala 160:64:@51516.4]
  assign _T_103182 = _T_103181[13:0]; // @[Modules.scala 160:64:@51517.4]
  assign buffer_15_587 = $signed(_T_103182); // @[Modules.scala 160:64:@51518.4]
  assign _T_103184 = $signed(buffer_15_561) + $signed(buffer_15_562); // @[Modules.scala 160:64:@51520.4]
  assign _T_103185 = _T_103184[13:0]; // @[Modules.scala 160:64:@51521.4]
  assign buffer_15_588 = $signed(_T_103185); // @[Modules.scala 160:64:@51522.4]
  assign _T_103187 = $signed(buffer_15_563) + $signed(buffer_15_564); // @[Modules.scala 160:64:@51524.4]
  assign _T_103188 = _T_103187[13:0]; // @[Modules.scala 160:64:@51525.4]
  assign buffer_15_589 = $signed(_T_103188); // @[Modules.scala 160:64:@51526.4]
  assign _T_103190 = $signed(buffer_15_565) + $signed(buffer_15_566); // @[Modules.scala 160:64:@51528.4]
  assign _T_103191 = _T_103190[13:0]; // @[Modules.scala 160:64:@51529.4]
  assign buffer_15_590 = $signed(_T_103191); // @[Modules.scala 160:64:@51530.4]
  assign _T_103193 = $signed(buffer_15_567) + $signed(buffer_15_568); // @[Modules.scala 160:64:@51532.4]
  assign _T_103194 = _T_103193[13:0]; // @[Modules.scala 160:64:@51533.4]
  assign buffer_15_591 = $signed(_T_103194); // @[Modules.scala 160:64:@51534.4]
  assign _T_103196 = $signed(buffer_15_569) + $signed(buffer_15_570); // @[Modules.scala 160:64:@51536.4]
  assign _T_103197 = _T_103196[13:0]; // @[Modules.scala 160:64:@51537.4]
  assign buffer_15_592 = $signed(_T_103197); // @[Modules.scala 160:64:@51538.4]
  assign _T_103199 = $signed(buffer_15_571) + $signed(buffer_15_572); // @[Modules.scala 160:64:@51540.4]
  assign _T_103200 = _T_103199[13:0]; // @[Modules.scala 160:64:@51541.4]
  assign buffer_15_593 = $signed(_T_103200); // @[Modules.scala 160:64:@51542.4]
  assign _T_103202 = $signed(buffer_15_573) + $signed(buffer_15_574); // @[Modules.scala 160:64:@51544.4]
  assign _T_103203 = _T_103202[13:0]; // @[Modules.scala 160:64:@51545.4]
  assign buffer_15_594 = $signed(_T_103203); // @[Modules.scala 160:64:@51546.4]
  assign _T_103205 = $signed(buffer_15_575) + $signed(buffer_15_576); // @[Modules.scala 160:64:@51548.4]
  assign _T_103206 = _T_103205[13:0]; // @[Modules.scala 160:64:@51549.4]
  assign buffer_15_595 = $signed(_T_103206); // @[Modules.scala 160:64:@51550.4]
  assign _T_103208 = $signed(buffer_15_577) + $signed(buffer_15_578); // @[Modules.scala 166:64:@51552.4]
  assign _T_103209 = _T_103208[13:0]; // @[Modules.scala 166:64:@51553.4]
  assign buffer_15_596 = $signed(_T_103209); // @[Modules.scala 166:64:@51554.4]
  assign _T_103211 = $signed(buffer_15_579) + $signed(buffer_15_580); // @[Modules.scala 166:64:@51556.4]
  assign _T_103212 = _T_103211[13:0]; // @[Modules.scala 166:64:@51557.4]
  assign buffer_15_597 = $signed(_T_103212); // @[Modules.scala 166:64:@51558.4]
  assign _T_103214 = $signed(buffer_15_581) + $signed(buffer_15_582); // @[Modules.scala 166:64:@51560.4]
  assign _T_103215 = _T_103214[13:0]; // @[Modules.scala 166:64:@51561.4]
  assign buffer_15_598 = $signed(_T_103215); // @[Modules.scala 166:64:@51562.4]
  assign _T_103217 = $signed(buffer_15_583) + $signed(buffer_15_584); // @[Modules.scala 166:64:@51564.4]
  assign _T_103218 = _T_103217[13:0]; // @[Modules.scala 166:64:@51565.4]
  assign buffer_15_599 = $signed(_T_103218); // @[Modules.scala 166:64:@51566.4]
  assign _T_103220 = $signed(buffer_15_585) + $signed(buffer_15_586); // @[Modules.scala 166:64:@51568.4]
  assign _T_103221 = _T_103220[13:0]; // @[Modules.scala 166:64:@51569.4]
  assign buffer_15_600 = $signed(_T_103221); // @[Modules.scala 166:64:@51570.4]
  assign _T_103223 = $signed(buffer_15_587) + $signed(buffer_15_588); // @[Modules.scala 166:64:@51572.4]
  assign _T_103224 = _T_103223[13:0]; // @[Modules.scala 166:64:@51573.4]
  assign buffer_15_601 = $signed(_T_103224); // @[Modules.scala 166:64:@51574.4]
  assign _T_103226 = $signed(buffer_15_589) + $signed(buffer_15_590); // @[Modules.scala 166:64:@51576.4]
  assign _T_103227 = _T_103226[13:0]; // @[Modules.scala 166:64:@51577.4]
  assign buffer_15_602 = $signed(_T_103227); // @[Modules.scala 166:64:@51578.4]
  assign _T_103229 = $signed(buffer_15_591) + $signed(buffer_15_592); // @[Modules.scala 166:64:@51580.4]
  assign _T_103230 = _T_103229[13:0]; // @[Modules.scala 166:64:@51581.4]
  assign buffer_15_603 = $signed(_T_103230); // @[Modules.scala 166:64:@51582.4]
  assign _T_103232 = $signed(buffer_15_593) + $signed(buffer_15_594); // @[Modules.scala 166:64:@51584.4]
  assign _T_103233 = _T_103232[13:0]; // @[Modules.scala 166:64:@51585.4]
  assign buffer_15_604 = $signed(_T_103233); // @[Modules.scala 166:64:@51586.4]
  assign _T_103235 = $signed(buffer_15_595) + $signed(buffer_15_538); // @[Modules.scala 172:66:@51588.4]
  assign _T_103236 = _T_103235[13:0]; // @[Modules.scala 172:66:@51589.4]
  assign buffer_15_605 = $signed(_T_103236); // @[Modules.scala 172:66:@51590.4]
  assign _T_103238 = $signed(buffer_15_596) + $signed(buffer_15_597); // @[Modules.scala 160:64:@51592.4]
  assign _T_103239 = _T_103238[13:0]; // @[Modules.scala 160:64:@51593.4]
  assign buffer_15_606 = $signed(_T_103239); // @[Modules.scala 160:64:@51594.4]
  assign _T_103241 = $signed(buffer_15_598) + $signed(buffer_15_599); // @[Modules.scala 160:64:@51596.4]
  assign _T_103242 = _T_103241[13:0]; // @[Modules.scala 160:64:@51597.4]
  assign buffer_15_607 = $signed(_T_103242); // @[Modules.scala 160:64:@51598.4]
  assign _T_103244 = $signed(buffer_15_600) + $signed(buffer_15_601); // @[Modules.scala 160:64:@51600.4]
  assign _T_103245 = _T_103244[13:0]; // @[Modules.scala 160:64:@51601.4]
  assign buffer_15_608 = $signed(_T_103245); // @[Modules.scala 160:64:@51602.4]
  assign _T_103247 = $signed(buffer_15_602) + $signed(buffer_15_603); // @[Modules.scala 160:64:@51604.4]
  assign _T_103248 = _T_103247[13:0]; // @[Modules.scala 160:64:@51605.4]
  assign buffer_15_609 = $signed(_T_103248); // @[Modules.scala 160:64:@51606.4]
  assign _T_103250 = $signed(buffer_15_604) + $signed(buffer_15_605); // @[Modules.scala 160:64:@51608.4]
  assign _T_103251 = _T_103250[13:0]; // @[Modules.scala 160:64:@51609.4]
  assign buffer_15_610 = $signed(_T_103251); // @[Modules.scala 160:64:@51610.4]
  assign _T_103253 = $signed(buffer_15_606) + $signed(buffer_15_607); // @[Modules.scala 166:64:@51612.4]
  assign _T_103254 = _T_103253[13:0]; // @[Modules.scala 166:64:@51613.4]
  assign buffer_15_611 = $signed(_T_103254); // @[Modules.scala 166:64:@51614.4]
  assign _T_103256 = $signed(buffer_15_608) + $signed(buffer_15_609); // @[Modules.scala 166:64:@51616.4]
  assign _T_103257 = _T_103256[13:0]; // @[Modules.scala 166:64:@51617.4]
  assign buffer_15_612 = $signed(_T_103257); // @[Modules.scala 166:64:@51618.4]
  assign _T_103259 = $signed(buffer_15_611) + $signed(buffer_15_612); // @[Modules.scala 160:64:@51620.4]
  assign _T_103260 = _T_103259[13:0]; // @[Modules.scala 160:64:@51621.4]
  assign buffer_15_613 = $signed(_T_103260); // @[Modules.scala 160:64:@51622.4]
  assign _T_103262 = $signed(buffer_15_613) + $signed(buffer_15_610); // @[Modules.scala 172:66:@51624.4]
  assign _T_103263 = _T_103262[13:0]; // @[Modules.scala 172:66:@51625.4]
  assign buffer_15_614 = $signed(_T_103263); // @[Modules.scala 172:66:@51626.4]
  assign io_out_0 = buffer_0_602;
  assign io_out_1 = buffer_1_606;
  assign io_out_2 = buffer_2_618;
  assign io_out_3 = buffer_3_626;
  assign io_out_4 = buffer_4_598;
  assign io_out_5 = buffer_5_626;
  assign io_out_6 = buffer_6_630;
  assign io_out_7 = buffer_7_616;
  assign io_out_8 = buffer_8_616;
  assign io_out_9 = buffer_9_626;
  assign io_out_10 = buffer_10_614;
  assign io_out_11 = buffer_11_596;
  assign io_out_12 = buffer_12_594;
  assign io_out_13 = buffer_13_612;
  assign io_out_14 = buffer_14_602;
  assign io_out_15 = buffer_15_614;
endmodule
module BN_BI( // @[:@52084.2]
  input  [13:0] io_in_0, // @[:@52087.4]
  input  [13:0] io_in_1, // @[:@52087.4]
  input  [13:0] io_in_2, // @[:@52087.4]
  input  [13:0] io_in_3, // @[:@52087.4]
  input  [13:0] io_in_4, // @[:@52087.4]
  input  [13:0] io_in_5, // @[:@52087.4]
  input  [13:0] io_in_6, // @[:@52087.4]
  input  [13:0] io_in_7, // @[:@52087.4]
  input  [13:0] io_in_8, // @[:@52087.4]
  input  [13:0] io_in_9, // @[:@52087.4]
  input  [13:0] io_in_10, // @[:@52087.4]
  input  [13:0] io_in_11, // @[:@52087.4]
  input  [13:0] io_in_12, // @[:@52087.4]
  input  [13:0] io_in_13, // @[:@52087.4]
  input  [13:0] io_in_14, // @[:@52087.4]
  input  [13:0] io_in_15, // @[:@52087.4]
  output [13:0] io_out_0, // @[:@52087.4]
  output [13:0] io_out_1, // @[:@52087.4]
  output [13:0] io_out_2, // @[:@52087.4]
  output [13:0] io_out_3, // @[:@52087.4]
  output [13:0] io_out_4, // @[:@52087.4]
  output [13:0] io_out_5, // @[:@52087.4]
  output [13:0] io_out_6, // @[:@52087.4]
  output [13:0] io_out_7, // @[:@52087.4]
  output [13:0] io_out_8, // @[:@52087.4]
  output [13:0] io_out_9, // @[:@52087.4]
  output [13:0] io_out_10, // @[:@52087.4]
  output [13:0] io_out_11, // @[:@52087.4]
  output [13:0] io_out_12, // @[:@52087.4]
  output [13:0] io_out_13, // @[:@52087.4]
  output [13:0] io_out_14, // @[:@52087.4]
  output [13:0] io_out_15 // @[:@52087.4]
);
  wire [14:0] _T_66; // @[Modules.scala 282:31:@52090.4]
  wire [13:0] _T_67; // @[Modules.scala 282:31:@52091.4]
  wire [13:0] buffer_0; // @[Modules.scala 282:31:@52092.4]
  wire  _T_70; // @[Modules.scala 283:24:@52094.4]
  wire [1:0] _GEN_0; // @[Modules.scala 283:32:@52095.4]
  wire [14:0] _T_74; // @[Modules.scala 282:31:@52101.4]
  wire [13:0] _T_75; // @[Modules.scala 282:31:@52102.4]
  wire [13:0] buffer_1; // @[Modules.scala 282:31:@52103.4]
  wire  _T_78; // @[Modules.scala 283:24:@52105.4]
  wire [1:0] _GEN_1; // @[Modules.scala 283:32:@52106.4]
  wire [14:0] _T_82; // @[Modules.scala 282:31:@52112.4]
  wire [13:0] _T_83; // @[Modules.scala 282:31:@52113.4]
  wire [13:0] buffer_2; // @[Modules.scala 282:31:@52114.4]
  wire  _T_86; // @[Modules.scala 283:24:@52116.4]
  wire [1:0] _GEN_2; // @[Modules.scala 283:32:@52117.4]
  wire [14:0] _T_90; // @[Modules.scala 282:31:@52123.4]
  wire [13:0] _T_91; // @[Modules.scala 282:31:@52124.4]
  wire [13:0] buffer_3; // @[Modules.scala 282:31:@52125.4]
  wire  _T_94; // @[Modules.scala 283:24:@52127.4]
  wire [1:0] _GEN_3; // @[Modules.scala 283:32:@52128.4]
  wire [14:0] _T_98; // @[Modules.scala 282:31:@52134.4]
  wire [13:0] _T_99; // @[Modules.scala 282:31:@52135.4]
  wire [13:0] buffer_4; // @[Modules.scala 282:31:@52136.4]
  wire  _T_102; // @[Modules.scala 283:24:@52138.4]
  wire [1:0] _GEN_4; // @[Modules.scala 283:32:@52139.4]
  wire [14:0] _T_106; // @[Modules.scala 282:31:@52145.4]
  wire [13:0] _T_107; // @[Modules.scala 282:31:@52146.4]
  wire [13:0] buffer_5; // @[Modules.scala 282:31:@52147.4]
  wire  _T_110; // @[Modules.scala 283:24:@52149.4]
  wire [1:0] _GEN_5; // @[Modules.scala 283:32:@52150.4]
  wire [14:0] _T_114; // @[Modules.scala 282:31:@52156.4]
  wire [13:0] _T_115; // @[Modules.scala 282:31:@52157.4]
  wire [13:0] buffer_6; // @[Modules.scala 282:31:@52158.4]
  wire  _T_118; // @[Modules.scala 283:24:@52160.4]
  wire [1:0] _GEN_6; // @[Modules.scala 283:32:@52161.4]
  wire [14:0] _T_122; // @[Modules.scala 282:31:@52167.4]
  wire [13:0] _T_123; // @[Modules.scala 282:31:@52168.4]
  wire [13:0] buffer_7; // @[Modules.scala 282:31:@52169.4]
  wire  _T_126; // @[Modules.scala 283:24:@52171.4]
  wire [1:0] _GEN_7; // @[Modules.scala 283:32:@52172.4]
  wire [14:0] _T_130; // @[Modules.scala 282:31:@52178.4]
  wire [13:0] _T_131; // @[Modules.scala 282:31:@52179.4]
  wire [13:0] buffer_8; // @[Modules.scala 282:31:@52180.4]
  wire  _T_134; // @[Modules.scala 283:24:@52182.4]
  wire [1:0] _GEN_8; // @[Modules.scala 283:32:@52183.4]
  wire [14:0] _T_138; // @[Modules.scala 282:31:@52189.4]
  wire [13:0] _T_139; // @[Modules.scala 282:31:@52190.4]
  wire [13:0] buffer_9; // @[Modules.scala 282:31:@52191.4]
  wire  _T_142; // @[Modules.scala 283:24:@52193.4]
  wire [1:0] _GEN_9; // @[Modules.scala 283:32:@52194.4]
  wire [14:0] _T_146; // @[Modules.scala 282:31:@52200.4]
  wire [13:0] _T_147; // @[Modules.scala 282:31:@52201.4]
  wire [13:0] buffer_10; // @[Modules.scala 282:31:@52202.4]
  wire  _T_150; // @[Modules.scala 283:24:@52204.4]
  wire [1:0] _GEN_10; // @[Modules.scala 283:32:@52205.4]
  wire [14:0] _T_154; // @[Modules.scala 282:31:@52211.4]
  wire [13:0] _T_155; // @[Modules.scala 282:31:@52212.4]
  wire [13:0] buffer_11; // @[Modules.scala 282:31:@52213.4]
  wire  _T_158; // @[Modules.scala 283:24:@52215.4]
  wire [1:0] _GEN_11; // @[Modules.scala 283:32:@52216.4]
  wire [14:0] _T_162; // @[Modules.scala 282:31:@52222.4]
  wire [13:0] _T_163; // @[Modules.scala 282:31:@52223.4]
  wire [13:0] buffer_12; // @[Modules.scala 282:31:@52224.4]
  wire  _T_166; // @[Modules.scala 283:24:@52226.4]
  wire [1:0] _GEN_12; // @[Modules.scala 283:32:@52227.4]
  wire [14:0] _T_170; // @[Modules.scala 282:31:@52233.4]
  wire [13:0] _T_171; // @[Modules.scala 282:31:@52234.4]
  wire [13:0] buffer_13; // @[Modules.scala 282:31:@52235.4]
  wire  _T_174; // @[Modules.scala 283:24:@52237.4]
  wire [1:0] _GEN_13; // @[Modules.scala 283:32:@52238.4]
  wire [14:0] _T_178; // @[Modules.scala 282:31:@52244.4]
  wire [13:0] _T_179; // @[Modules.scala 282:31:@52245.4]
  wire [13:0] buffer_14; // @[Modules.scala 282:31:@52246.4]
  wire  _T_182; // @[Modules.scala 283:24:@52248.4]
  wire [1:0] _GEN_14; // @[Modules.scala 283:32:@52249.4]
  wire [14:0] _T_186; // @[Modules.scala 282:31:@52255.4]
  wire [13:0] _T_187; // @[Modules.scala 282:31:@52256.4]
  wire [13:0] buffer_15; // @[Modules.scala 282:31:@52257.4]
  wire  _T_190; // @[Modules.scala 283:24:@52259.4]
  wire [1:0] _GEN_15; // @[Modules.scala 283:32:@52260.4]
  assign _T_66 = $signed(io_in_0) - $signed(-14'sh56); // @[Modules.scala 282:31:@52090.4]
  assign _T_67 = _T_66[13:0]; // @[Modules.scala 282:31:@52091.4]
  assign buffer_0 = $signed(_T_67); // @[Modules.scala 282:31:@52092.4]
  assign _T_70 = $signed(buffer_0) >= $signed(14'sh0); // @[Modules.scala 283:24:@52094.4]
  assign _GEN_0 = _T_70 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52095.4]
  assign _T_74 = $signed(io_in_1) - $signed(-14'sh15); // @[Modules.scala 282:31:@52101.4]
  assign _T_75 = _T_74[13:0]; // @[Modules.scala 282:31:@52102.4]
  assign buffer_1 = $signed(_T_75); // @[Modules.scala 282:31:@52103.4]
  assign _T_78 = $signed(buffer_1) >= $signed(14'sh0); // @[Modules.scala 283:24:@52105.4]
  assign _GEN_1 = _T_78 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52106.4]
  assign _T_82 = $signed(io_in_2) - $signed(14'sh90); // @[Modules.scala 282:31:@52112.4]
  assign _T_83 = _T_82[13:0]; // @[Modules.scala 282:31:@52113.4]
  assign buffer_2 = $signed(_T_83); // @[Modules.scala 282:31:@52114.4]
  assign _T_86 = $signed(buffer_2) >= $signed(14'sh0); // @[Modules.scala 283:24:@52116.4]
  assign _GEN_2 = _T_86 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52117.4]
  assign _T_90 = $signed(io_in_3) - $signed(14'sh7a); // @[Modules.scala 282:31:@52123.4]
  assign _T_91 = _T_90[13:0]; // @[Modules.scala 282:31:@52124.4]
  assign buffer_3 = $signed(_T_91); // @[Modules.scala 282:31:@52125.4]
  assign _T_94 = $signed(buffer_3) >= $signed(14'sh0); // @[Modules.scala 283:24:@52127.4]
  assign _GEN_3 = _T_94 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52128.4]
  assign _T_98 = $signed(io_in_4) - $signed(14'sh6a); // @[Modules.scala 282:31:@52134.4]
  assign _T_99 = _T_98[13:0]; // @[Modules.scala 282:31:@52135.4]
  assign buffer_4 = $signed(_T_99); // @[Modules.scala 282:31:@52136.4]
  assign _T_102 = $signed(buffer_4) >= $signed(14'sh0); // @[Modules.scala 283:24:@52138.4]
  assign _GEN_4 = _T_102 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52139.4]
  assign _T_106 = $signed(io_in_5) - $signed(-14'sh69); // @[Modules.scala 282:31:@52145.4]
  assign _T_107 = _T_106[13:0]; // @[Modules.scala 282:31:@52146.4]
  assign buffer_5 = $signed(_T_107); // @[Modules.scala 282:31:@52147.4]
  assign _T_110 = $signed(buffer_5) >= $signed(14'sh0); // @[Modules.scala 283:24:@52149.4]
  assign _GEN_5 = _T_110 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52150.4]
  assign _T_114 = $signed(io_in_6) - $signed(-14'sh34); // @[Modules.scala 282:31:@52156.4]
  assign _T_115 = _T_114[13:0]; // @[Modules.scala 282:31:@52157.4]
  assign buffer_6 = $signed(_T_115); // @[Modules.scala 282:31:@52158.4]
  assign _T_118 = $signed(buffer_6) >= $signed(14'sh0); // @[Modules.scala 283:24:@52160.4]
  assign _GEN_6 = _T_118 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52161.4]
  assign _T_122 = $signed(io_in_7) - $signed(-14'sh7); // @[Modules.scala 282:31:@52167.4]
  assign _T_123 = _T_122[13:0]; // @[Modules.scala 282:31:@52168.4]
  assign buffer_7 = $signed(_T_123); // @[Modules.scala 282:31:@52169.4]
  assign _T_126 = $signed(buffer_7) >= $signed(14'sh0); // @[Modules.scala 283:24:@52171.4]
  assign _GEN_7 = _T_126 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52172.4]
  assign _T_130 = $signed(io_in_8) - $signed(-14'she); // @[Modules.scala 282:31:@52178.4]
  assign _T_131 = _T_130[13:0]; // @[Modules.scala 282:31:@52179.4]
  assign buffer_8 = $signed(_T_131); // @[Modules.scala 282:31:@52180.4]
  assign _T_134 = $signed(buffer_8) >= $signed(14'sh0); // @[Modules.scala 283:24:@52182.4]
  assign _GEN_8 = _T_134 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52183.4]
  assign _T_138 = $signed(io_in_9) - $signed(-14'sh17); // @[Modules.scala 282:31:@52189.4]
  assign _T_139 = _T_138[13:0]; // @[Modules.scala 282:31:@52190.4]
  assign buffer_9 = $signed(_T_139); // @[Modules.scala 282:31:@52191.4]
  assign _T_142 = $signed(buffer_9) >= $signed(14'sh0); // @[Modules.scala 283:24:@52193.4]
  assign _GEN_9 = _T_142 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52194.4]
  assign _T_146 = $signed(io_in_10) - $signed(14'sh2f); // @[Modules.scala 282:31:@52200.4]
  assign _T_147 = _T_146[13:0]; // @[Modules.scala 282:31:@52201.4]
  assign buffer_10 = $signed(_T_147); // @[Modules.scala 282:31:@52202.4]
  assign _T_150 = $signed(buffer_10) >= $signed(14'sh0); // @[Modules.scala 283:24:@52204.4]
  assign _GEN_10 = _T_150 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52205.4]
  assign _T_154 = $signed(io_in_11) - $signed(14'sh3d); // @[Modules.scala 282:31:@52211.4]
  assign _T_155 = _T_154[13:0]; // @[Modules.scala 282:31:@52212.4]
  assign buffer_11 = $signed(_T_155); // @[Modules.scala 282:31:@52213.4]
  assign _T_158 = $signed(buffer_11) >= $signed(14'sh0); // @[Modules.scala 283:24:@52215.4]
  assign _GEN_11 = _T_158 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52216.4]
  assign _T_162 = $signed(io_in_12) - $signed(14'sh22); // @[Modules.scala 282:31:@52222.4]
  assign _T_163 = _T_162[13:0]; // @[Modules.scala 282:31:@52223.4]
  assign buffer_12 = $signed(_T_163); // @[Modules.scala 282:31:@52224.4]
  assign _T_166 = $signed(buffer_12) >= $signed(14'sh0); // @[Modules.scala 283:24:@52226.4]
  assign _GEN_12 = _T_166 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52227.4]
  assign _T_170 = $signed(io_in_13) - $signed(-14'sh6); // @[Modules.scala 282:31:@52233.4]
  assign _T_171 = _T_170[13:0]; // @[Modules.scala 282:31:@52234.4]
  assign buffer_13 = $signed(_T_171); // @[Modules.scala 282:31:@52235.4]
  assign _T_174 = $signed(buffer_13) >= $signed(14'sh0); // @[Modules.scala 283:24:@52237.4]
  assign _GEN_13 = _T_174 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52238.4]
  assign _T_178 = $signed(io_in_14) - $signed(-14'sh5); // @[Modules.scala 282:31:@52244.4]
  assign _T_179 = _T_178[13:0]; // @[Modules.scala 282:31:@52245.4]
  assign buffer_14 = $signed(_T_179); // @[Modules.scala 282:31:@52246.4]
  assign _T_182 = $signed(buffer_14) >= $signed(14'sh0); // @[Modules.scala 283:24:@52248.4]
  assign _GEN_14 = _T_182 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52249.4]
  assign _T_186 = $signed(io_in_15) - $signed(-14'sh6d); // @[Modules.scala 282:31:@52255.4]
  assign _T_187 = _T_186[13:0]; // @[Modules.scala 282:31:@52256.4]
  assign buffer_15 = $signed(_T_187); // @[Modules.scala 282:31:@52257.4]
  assign _T_190 = $signed(buffer_15) >= $signed(14'sh0); // @[Modules.scala 283:24:@52259.4]
  assign _GEN_15 = _T_190 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@52260.4]
  assign io_out_0 = {{12{_GEN_0[1]}},_GEN_0};
  assign io_out_1 = {{12{_GEN_1[1]}},_GEN_1};
  assign io_out_2 = {{12{_GEN_2[1]}},_GEN_2};
  assign io_out_3 = {{12{_GEN_3[1]}},_GEN_3};
  assign io_out_4 = {{12{_GEN_4[1]}},_GEN_4};
  assign io_out_5 = {{12{_GEN_5[1]}},_GEN_5};
  assign io_out_6 = {{12{_GEN_6[1]}},_GEN_6};
  assign io_out_7 = {{12{_GEN_7[1]}},_GEN_7};
  assign io_out_8 = {{12{_GEN_8[1]}},_GEN_8};
  assign io_out_9 = {{12{_GEN_9[1]}},_GEN_9};
  assign io_out_10 = {{12{_GEN_10[1]}},_GEN_10};
  assign io_out_11 = {{12{_GEN_11[1]}},_GEN_11};
  assign io_out_12 = {{12{_GEN_12[1]}},_GEN_12};
  assign io_out_13 = {{12{_GEN_13[1]}},_GEN_13};
  assign io_out_14 = {{12{_GEN_14[1]}},_GEN_14};
  assign io_out_15 = {{12{_GEN_15[1]}},_GEN_15};
endmodule
module Linear_p_1( // @[:@52267.2]
  input  [1:0] io_in_0, // @[:@52270.4]
  input  [1:0] io_in_1, // @[:@52270.4]
  input  [1:0] io_in_2, // @[:@52270.4]
  input  [1:0] io_in_3, // @[:@52270.4]
  input  [1:0] io_in_4, // @[:@52270.4]
  input  [1:0] io_in_5, // @[:@52270.4]
  input  [1:0] io_in_6, // @[:@52270.4]
  input  [1:0] io_in_7, // @[:@52270.4]
  input  [1:0] io_in_8, // @[:@52270.4]
  input  [1:0] io_in_9, // @[:@52270.4]
  input  [1:0] io_in_10, // @[:@52270.4]
  input  [1:0] io_in_11, // @[:@52270.4]
  input  [1:0] io_in_12, // @[:@52270.4]
  input  [1:0] io_in_13, // @[:@52270.4]
  input  [1:0] io_in_14, // @[:@52270.4]
  input  [1:0] io_in_15, // @[:@52270.4]
  output [5:0] io_out_0, // @[:@52270.4]
  output [5:0] io_out_1, // @[:@52270.4]
  output [5:0] io_out_2, // @[:@52270.4]
  output [5:0] io_out_3, // @[:@52270.4]
  output [5:0] io_out_4, // @[:@52270.4]
  output [5:0] io_out_5, // @[:@52270.4]
  output [5:0] io_out_6, // @[:@52270.4]
  output [5:0] io_out_7, // @[:@52270.4]
  output [5:0] io_out_8, // @[:@52270.4]
  output [5:0] io_out_9, // @[:@52270.4]
  output [5:0] io_out_10, // @[:@52270.4]
  output [5:0] io_out_11, // @[:@52270.4]
  output [5:0] io_out_12, // @[:@52270.4]
  output [5:0] io_out_13, // @[:@52270.4]
  output [5:0] io_out_14, // @[:@52270.4]
  output [5:0] io_out_15 // @[:@52270.4]
);
  wire [3:0] _T_1207; // @[Modules.scala 143:74:@52273.4]
  wire [3:0] _T_1209; // @[Modules.scala 144:80:@52274.4]
  wire [4:0] _T_1210; // @[Modules.scala 143:103:@52275.4]
  wire [3:0] _T_1211; // @[Modules.scala 143:103:@52276.4]
  wire [3:0] _T_1212; // @[Modules.scala 143:103:@52277.4]
  wire [3:0] _T_1214; // @[Modules.scala 143:74:@52279.4]
  wire [3:0] _T_1216; // @[Modules.scala 144:80:@52280.4]
  wire [4:0] _T_1217; // @[Modules.scala 143:103:@52281.4]
  wire [3:0] _T_1218; // @[Modules.scala 143:103:@52282.4]
  wire [3:0] _T_1219; // @[Modules.scala 143:103:@52283.4]
  wire [3:0] _T_1221; // @[Modules.scala 143:74:@52285.4]
  wire [2:0] _T_1223; // @[Modules.scala 144:80:@52286.4]
  wire [3:0] _GEN_0; // @[Modules.scala 143:103:@52287.4]
  wire [4:0] _T_1224; // @[Modules.scala 143:103:@52287.4]
  wire [3:0] _T_1225; // @[Modules.scala 143:103:@52288.4]
  wire [3:0] _T_1226; // @[Modules.scala 143:103:@52289.4]
  wire [3:0] _T_1228; // @[Modules.scala 143:74:@52291.4]
  wire [2:0] _T_1230; // @[Modules.scala 144:80:@52292.4]
  wire [3:0] _GEN_1; // @[Modules.scala 143:103:@52293.4]
  wire [4:0] _T_1231; // @[Modules.scala 143:103:@52293.4]
  wire [3:0] _T_1232; // @[Modules.scala 143:103:@52294.4]
  wire [3:0] _T_1233; // @[Modules.scala 143:103:@52295.4]
  wire [3:0] _T_1235; // @[Modules.scala 143:74:@52297.4]
  wire [3:0] _T_1237; // @[Modules.scala 144:80:@52298.4]
  wire [4:0] _T_1238; // @[Modules.scala 143:103:@52299.4]
  wire [3:0] _T_1239; // @[Modules.scala 143:103:@52300.4]
  wire [3:0] _T_1240; // @[Modules.scala 143:103:@52301.4]
  wire [3:0] _T_1242; // @[Modules.scala 143:74:@52303.4]
  wire [2:0] _T_1244; // @[Modules.scala 144:80:@52304.4]
  wire [3:0] _GEN_2; // @[Modules.scala 143:103:@52305.4]
  wire [4:0] _T_1245; // @[Modules.scala 143:103:@52305.4]
  wire [3:0] _T_1246; // @[Modules.scala 143:103:@52306.4]
  wire [3:0] _T_1247; // @[Modules.scala 143:103:@52307.4]
  wire [2:0] _T_1249; // @[Modules.scala 143:74:@52309.4]
  wire [2:0] _T_1251; // @[Modules.scala 144:80:@52310.4]
  wire [3:0] _T_1252; // @[Modules.scala 143:103:@52311.4]
  wire [2:0] _T_1253; // @[Modules.scala 143:103:@52312.4]
  wire [2:0] _T_1254; // @[Modules.scala 143:103:@52313.4]
  wire [5:0] buffer_0_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_0_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1255; // @[Modules.scala 166:64:@52315.4]
  wire [5:0] _T_1256; // @[Modules.scala 166:64:@52316.4]
  wire [5:0] buffer_0_7; // @[Modules.scala 166:64:@52317.4]
  wire [5:0] buffer_0_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_0_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1258; // @[Modules.scala 166:64:@52319.4]
  wire [5:0] _T_1259; // @[Modules.scala 166:64:@52320.4]
  wire [5:0] buffer_0_8; // @[Modules.scala 166:64:@52321.4]
  wire [5:0] buffer_0_4; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_0_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1261; // @[Modules.scala 166:64:@52323.4]
  wire [5:0] _T_1262; // @[Modules.scala 166:64:@52324.4]
  wire [5:0] buffer_0_9; // @[Modules.scala 166:64:@52325.4]
  wire [6:0] _T_1264; // @[Modules.scala 166:64:@52327.4]
  wire [5:0] _T_1265; // @[Modules.scala 166:64:@52328.4]
  wire [5:0] buffer_0_10; // @[Modules.scala 166:64:@52329.4]
  wire [5:0] buffer_0_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1267; // @[Modules.scala 172:66:@52331.4]
  wire [5:0] _T_1268; // @[Modules.scala 172:66:@52332.4]
  wire [5:0] buffer_0_11; // @[Modules.scala 172:66:@52333.4]
  wire [6:0] _T_1270; // @[Modules.scala 160:64:@52335.4]
  wire [5:0] _T_1271; // @[Modules.scala 160:64:@52336.4]
  wire [5:0] buffer_0_12; // @[Modules.scala 160:64:@52337.4]
  wire [2:0] _T_1274; // @[Modules.scala 143:74:@52342.4]
  wire [3:0] _GEN_3; // @[Modules.scala 143:103:@52344.4]
  wire [4:0] _T_1277; // @[Modules.scala 143:103:@52344.4]
  wire [3:0] _T_1278; // @[Modules.scala 143:103:@52345.4]
  wire [3:0] _T_1279; // @[Modules.scala 143:103:@52346.4]
  wire [2:0] _T_1283; // @[Modules.scala 144:80:@52349.4]
  wire [3:0] _GEN_4; // @[Modules.scala 143:103:@52350.4]
  wire [4:0] _T_1284; // @[Modules.scala 143:103:@52350.4]
  wire [3:0] _T_1285; // @[Modules.scala 143:103:@52351.4]
  wire [3:0] _T_1286; // @[Modules.scala 143:103:@52352.4]
  wire [3:0] _T_1288; // @[Modules.scala 143:74:@52354.4]
  wire [2:0] _T_1290; // @[Modules.scala 144:80:@52355.4]
  wire [3:0] _GEN_5; // @[Modules.scala 143:103:@52356.4]
  wire [4:0] _T_1291; // @[Modules.scala 143:103:@52356.4]
  wire [3:0] _T_1292; // @[Modules.scala 143:103:@52357.4]
  wire [3:0] _T_1293; // @[Modules.scala 143:103:@52358.4]
  wire [2:0] _T_1295; // @[Modules.scala 143:74:@52360.4]
  wire [3:0] _T_1298; // @[Modules.scala 143:103:@52362.4]
  wire [2:0] _T_1299; // @[Modules.scala 143:103:@52363.4]
  wire [2:0] _T_1300; // @[Modules.scala 143:103:@52364.4]
  wire [2:0] _T_1302; // @[Modules.scala 143:74:@52366.4]
  wire [3:0] _GEN_6; // @[Modules.scala 143:103:@52368.4]
  wire [4:0] _T_1305; // @[Modules.scala 143:103:@52368.4]
  wire [3:0] _T_1306; // @[Modules.scala 143:103:@52369.4]
  wire [3:0] _T_1307; // @[Modules.scala 143:103:@52370.4]
  wire [3:0] _T_1316; // @[Modules.scala 143:74:@52378.4]
  wire [3:0] _GEN_8; // @[Modules.scala 143:103:@52380.4]
  wire [4:0] _T_1319; // @[Modules.scala 143:103:@52380.4]
  wire [3:0] _T_1320; // @[Modules.scala 143:103:@52381.4]
  wire [3:0] _T_1321; // @[Modules.scala 143:103:@52382.4]
  wire [5:0] buffer_1_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_1_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1322; // @[Modules.scala 166:64:@52384.4]
  wire [5:0] _T_1323; // @[Modules.scala 166:64:@52385.4]
  wire [5:0] buffer_1_7; // @[Modules.scala 166:64:@52386.4]
  wire [5:0] buffer_1_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_1_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1325; // @[Modules.scala 166:64:@52388.4]
  wire [5:0] _T_1326; // @[Modules.scala 166:64:@52389.4]
  wire [5:0] buffer_1_8; // @[Modules.scala 166:64:@52390.4]
  wire [5:0] buffer_1_4; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1328; // @[Modules.scala 166:64:@52392.4]
  wire [5:0] _T_1329; // @[Modules.scala 166:64:@52393.4]
  wire [5:0] buffer_1_9; // @[Modules.scala 166:64:@52394.4]
  wire [6:0] _T_1331; // @[Modules.scala 166:64:@52396.4]
  wire [5:0] _T_1332; // @[Modules.scala 166:64:@52397.4]
  wire [5:0] buffer_1_10; // @[Modules.scala 166:64:@52398.4]
  wire [5:0] buffer_1_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1334; // @[Modules.scala 172:66:@52400.4]
  wire [5:0] _T_1335; // @[Modules.scala 172:66:@52401.4]
  wire [5:0] buffer_1_11; // @[Modules.scala 172:66:@52402.4]
  wire [6:0] _T_1337; // @[Modules.scala 160:64:@52404.4]
  wire [5:0] _T_1338; // @[Modules.scala 160:64:@52405.4]
  wire [5:0] buffer_1_12; // @[Modules.scala 160:64:@52406.4]
  wire [4:0] _T_1344; // @[Modules.scala 150:103:@52413.4]
  wire [3:0] _T_1345; // @[Modules.scala 150:103:@52414.4]
  wire [3:0] _T_1346; // @[Modules.scala 150:103:@52415.4]
  wire [4:0] _T_1351; // @[Modules.scala 150:103:@52419.4]
  wire [3:0] _T_1352; // @[Modules.scala 150:103:@52420.4]
  wire [3:0] _T_1353; // @[Modules.scala 150:103:@52421.4]
  wire [4:0] _T_1358; // @[Modules.scala 150:103:@52425.4]
  wire [3:0] _T_1359; // @[Modules.scala 150:103:@52426.4]
  wire [3:0] _T_1360; // @[Modules.scala 150:103:@52427.4]
  wire [3:0] _T_1362; // @[Modules.scala 150:74:@52429.4]
  wire [4:0] _T_1365; // @[Modules.scala 150:103:@52431.4]
  wire [3:0] _T_1366; // @[Modules.scala 150:103:@52432.4]
  wire [3:0] _T_1367; // @[Modules.scala 150:103:@52433.4]
  wire [2:0] _T_1371; // @[Modules.scala 151:80:@52436.4]
  wire [3:0] _GEN_12; // @[Modules.scala 150:103:@52437.4]
  wire [4:0] _T_1372; // @[Modules.scala 150:103:@52437.4]
  wire [3:0] _T_1373; // @[Modules.scala 150:103:@52438.4]
  wire [3:0] _T_1374; // @[Modules.scala 150:103:@52439.4]
  wire [3:0] _T_1376; // @[Modules.scala 150:74:@52441.4]
  wire [3:0] _T_1378; // @[Modules.scala 151:80:@52442.4]
  wire [4:0] _T_1379; // @[Modules.scala 150:103:@52443.4]
  wire [3:0] _T_1380; // @[Modules.scala 150:103:@52444.4]
  wire [3:0] _T_1381; // @[Modules.scala 150:103:@52445.4]
  wire [3:0] _T_1383; // @[Modules.scala 153:80:@52447.4]
  wire [5:0] buffer_2_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_2_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1384; // @[Modules.scala 166:64:@52449.4]
  wire [5:0] _T_1385; // @[Modules.scala 166:64:@52450.4]
  wire [5:0] buffer_2_7; // @[Modules.scala 166:64:@52451.4]
  wire [5:0] buffer_2_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_2_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1387; // @[Modules.scala 166:64:@52453.4]
  wire [5:0] _T_1388; // @[Modules.scala 166:64:@52454.4]
  wire [5:0] buffer_2_8; // @[Modules.scala 166:64:@52455.4]
  wire [5:0] buffer_2_4; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_2_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1390; // @[Modules.scala 166:64:@52457.4]
  wire [5:0] _T_1391; // @[Modules.scala 166:64:@52458.4]
  wire [5:0] buffer_2_9; // @[Modules.scala 166:64:@52459.4]
  wire [6:0] _T_1393; // @[Modules.scala 166:64:@52461.4]
  wire [5:0] _T_1394; // @[Modules.scala 166:64:@52462.4]
  wire [5:0] buffer_2_10; // @[Modules.scala 166:64:@52463.4]
  wire [5:0] buffer_2_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1396; // @[Modules.scala 172:66:@52465.4]
  wire [5:0] _T_1397; // @[Modules.scala 172:66:@52466.4]
  wire [5:0] buffer_2_11; // @[Modules.scala 172:66:@52467.4]
  wire [6:0] _T_1399; // @[Modules.scala 160:64:@52469.4]
  wire [5:0] _T_1400; // @[Modules.scala 160:64:@52470.4]
  wire [5:0] buffer_2_12; // @[Modules.scala 160:64:@52471.4]
  wire [2:0] _T_1405; // @[Modules.scala 144:80:@52477.4]
  wire [3:0] _GEN_13; // @[Modules.scala 143:103:@52478.4]
  wire [4:0] _T_1406; // @[Modules.scala 143:103:@52478.4]
  wire [3:0] _T_1407; // @[Modules.scala 143:103:@52479.4]
  wire [3:0] _T_1408; // @[Modules.scala 143:103:@52480.4]
  wire [4:0] _T_1413; // @[Modules.scala 143:103:@52484.4]
  wire [3:0] _T_1414; // @[Modules.scala 143:103:@52485.4]
  wire [3:0] _T_1415; // @[Modules.scala 143:103:@52486.4]
  wire [3:0] _T_1417; // @[Modules.scala 143:74:@52488.4]
  wire [4:0] _T_1420; // @[Modules.scala 143:103:@52490.4]
  wire [3:0] _T_1421; // @[Modules.scala 143:103:@52491.4]
  wire [3:0] _T_1422; // @[Modules.scala 143:103:@52492.4]
  wire [4:0] _T_1434; // @[Modules.scala 143:103:@52502.4]
  wire [3:0] _T_1435; // @[Modules.scala 143:103:@52503.4]
  wire [3:0] _T_1436; // @[Modules.scala 143:103:@52504.4]
  wire [4:0] _T_1441; // @[Modules.scala 143:103:@52508.4]
  wire [3:0] _T_1442; // @[Modules.scala 143:103:@52509.4]
  wire [3:0] _T_1443; // @[Modules.scala 143:103:@52510.4]
  wire [5:0] buffer_3_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_3_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1444; // @[Modules.scala 160:64:@52512.4]
  wire [5:0] _T_1445; // @[Modules.scala 160:64:@52513.4]
  wire [5:0] buffer_3_6; // @[Modules.scala 160:64:@52514.4]
  wire [5:0] buffer_3_2; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1447; // @[Modules.scala 160:64:@52516.4]
  wire [5:0] _T_1448; // @[Modules.scala 160:64:@52517.4]
  wire [5:0] buffer_3_7; // @[Modules.scala 160:64:@52518.4]
  wire [5:0] buffer_3_4; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_3_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1450; // @[Modules.scala 160:64:@52520.4]
  wire [5:0] _T_1451; // @[Modules.scala 160:64:@52521.4]
  wire [5:0] buffer_3_8; // @[Modules.scala 160:64:@52522.4]
  wire [6:0] _T_1453; // @[Modules.scala 166:64:@52524.4]
  wire [5:0] _T_1454; // @[Modules.scala 166:64:@52525.4]
  wire [5:0] buffer_3_9; // @[Modules.scala 166:64:@52526.4]
  wire [6:0] _T_1456; // @[Modules.scala 172:66:@52528.4]
  wire [5:0] _T_1457; // @[Modules.scala 172:66:@52529.4]
  wire [5:0] buffer_3_10; // @[Modules.scala 172:66:@52530.4]
  wire [2:0] _T_1460; // @[Modules.scala 143:74:@52537.4]
  wire [3:0] _GEN_15; // @[Modules.scala 143:103:@52539.4]
  wire [4:0] _T_1463; // @[Modules.scala 143:103:@52539.4]
  wire [3:0] _T_1464; // @[Modules.scala 143:103:@52540.4]
  wire [3:0] _T_1465; // @[Modules.scala 143:103:@52541.4]
  wire [4:0] _T_1470; // @[Modules.scala 143:103:@52545.4]
  wire [3:0] _T_1471; // @[Modules.scala 143:103:@52546.4]
  wire [3:0] _T_1472; // @[Modules.scala 143:103:@52547.4]
  wire [3:0] _T_1477; // @[Modules.scala 143:103:@52551.4]
  wire [2:0] _T_1478; // @[Modules.scala 143:103:@52552.4]
  wire [2:0] _T_1479; // @[Modules.scala 143:103:@52553.4]
  wire [4:0] _T_1484; // @[Modules.scala 143:103:@52557.4]
  wire [3:0] _T_1485; // @[Modules.scala 143:103:@52558.4]
  wire [3:0] _T_1486; // @[Modules.scala 143:103:@52559.4]
  wire [4:0] _T_1491; // @[Modules.scala 143:103:@52563.4]
  wire [3:0] _T_1492; // @[Modules.scala 143:103:@52564.4]
  wire [3:0] _T_1493; // @[Modules.scala 143:103:@52565.4]
  wire [2:0] _T_1497; // @[Modules.scala 144:80:@52568.4]
  wire [3:0] _GEN_17; // @[Modules.scala 143:103:@52569.4]
  wire [4:0] _T_1498; // @[Modules.scala 143:103:@52569.4]
  wire [3:0] _T_1499; // @[Modules.scala 143:103:@52570.4]
  wire [3:0] _T_1500; // @[Modules.scala 143:103:@52571.4]
  wire [5:0] buffer_4_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_4_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1508; // @[Modules.scala 166:64:@52579.4]
  wire [5:0] _T_1509; // @[Modules.scala 166:64:@52580.4]
  wire [5:0] buffer_4_7; // @[Modules.scala 166:64:@52581.4]
  wire [5:0] buffer_4_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_4_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1511; // @[Modules.scala 166:64:@52583.4]
  wire [5:0] _T_1512; // @[Modules.scala 166:64:@52584.4]
  wire [5:0] buffer_4_8; // @[Modules.scala 166:64:@52585.4]
  wire [5:0] buffer_4_4; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_4_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1514; // @[Modules.scala 166:64:@52587.4]
  wire [5:0] _T_1515; // @[Modules.scala 166:64:@52588.4]
  wire [5:0] buffer_4_9; // @[Modules.scala 166:64:@52589.4]
  wire [6:0] _T_1517; // @[Modules.scala 166:64:@52591.4]
  wire [5:0] _T_1518; // @[Modules.scala 166:64:@52592.4]
  wire [5:0] buffer_4_10; // @[Modules.scala 166:64:@52593.4]
  wire [6:0] _T_1520; // @[Modules.scala 172:66:@52595.4]
  wire [5:0] _T_1521; // @[Modules.scala 172:66:@52596.4]
  wire [5:0] buffer_4_11; // @[Modules.scala 172:66:@52597.4]
  wire [6:0] _T_1523; // @[Modules.scala 160:64:@52599.4]
  wire [5:0] _T_1524; // @[Modules.scala 160:64:@52600.4]
  wire [5:0] buffer_4_12; // @[Modules.scala 160:64:@52601.4]
  wire [4:0] _T_1530; // @[Modules.scala 150:103:@52608.4]
  wire [3:0] _T_1531; // @[Modules.scala 150:103:@52609.4]
  wire [3:0] _T_1532; // @[Modules.scala 150:103:@52610.4]
  wire [2:0] _T_1534; // @[Modules.scala 150:74:@52612.4]
  wire [3:0] _T_1537; // @[Modules.scala 150:103:@52614.4]
  wire [2:0] _T_1538; // @[Modules.scala 150:103:@52615.4]
  wire [2:0] _T_1539; // @[Modules.scala 150:103:@52616.4]
  wire [4:0] _T_1544; // @[Modules.scala 150:103:@52620.4]
  wire [3:0] _T_1545; // @[Modules.scala 150:103:@52621.4]
  wire [3:0] _T_1546; // @[Modules.scala 150:103:@52622.4]
  wire [2:0] _T_1557; // @[Modules.scala 151:80:@52631.4]
  wire [3:0] _GEN_19; // @[Modules.scala 150:103:@52632.4]
  wire [4:0] _T_1558; // @[Modules.scala 150:103:@52632.4]
  wire [3:0] _T_1559; // @[Modules.scala 150:103:@52633.4]
  wire [3:0] _T_1560; // @[Modules.scala 150:103:@52634.4]
  wire [5:0] buffer_5_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_5_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1577; // @[Modules.scala 160:64:@52650.4]
  wire [5:0] _T_1578; // @[Modules.scala 160:64:@52651.4]
  wire [5:0] buffer_5_8; // @[Modules.scala 160:64:@52652.4]
  wire [5:0] buffer_5_2; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1580; // @[Modules.scala 160:64:@52654.4]
  wire [5:0] _T_1581; // @[Modules.scala 160:64:@52655.4]
  wire [5:0] buffer_5_9; // @[Modules.scala 160:64:@52656.4]
  wire [5:0] buffer_5_4; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1583; // @[Modules.scala 160:64:@52658.4]
  wire [5:0] _T_1584; // @[Modules.scala 160:64:@52659.4]
  wire [5:0] buffer_5_10; // @[Modules.scala 160:64:@52660.4]
  wire [6:0] _T_1586; // @[Modules.scala 160:64:@52662.4]
  wire [5:0] _T_1587; // @[Modules.scala 160:64:@52663.4]
  wire [5:0] buffer_5_11; // @[Modules.scala 160:64:@52664.4]
  wire [6:0] _T_1589; // @[Modules.scala 160:64:@52666.4]
  wire [5:0] _T_1590; // @[Modules.scala 160:64:@52667.4]
  wire [5:0] buffer_5_12; // @[Modules.scala 160:64:@52668.4]
  wire [6:0] _T_1592; // @[Modules.scala 160:64:@52670.4]
  wire [5:0] _T_1593; // @[Modules.scala 160:64:@52671.4]
  wire [5:0] buffer_5_13; // @[Modules.scala 160:64:@52672.4]
  wire [6:0] _T_1595; // @[Modules.scala 160:64:@52674.4]
  wire [5:0] _T_1596; // @[Modules.scala 160:64:@52675.4]
  wire [5:0] buffer_5_14; // @[Modules.scala 160:64:@52676.4]
  wire [3:0] _T_1602; // @[Modules.scala 143:103:@52681.4]
  wire [2:0] _T_1603; // @[Modules.scala 143:103:@52682.4]
  wire [2:0] _T_1604; // @[Modules.scala 143:103:@52683.4]
  wire [4:0] _T_1609; // @[Modules.scala 143:103:@52687.4]
  wire [3:0] _T_1610; // @[Modules.scala 143:103:@52688.4]
  wire [3:0] _T_1611; // @[Modules.scala 143:103:@52689.4]
  wire [4:0] _T_1616; // @[Modules.scala 143:103:@52693.4]
  wire [3:0] _T_1617; // @[Modules.scala 143:103:@52694.4]
  wire [3:0] _T_1618; // @[Modules.scala 143:103:@52695.4]
  wire [4:0] _T_1623; // @[Modules.scala 143:103:@52699.4]
  wire [3:0] _T_1624; // @[Modules.scala 143:103:@52700.4]
  wire [3:0] _T_1625; // @[Modules.scala 143:103:@52701.4]
  wire [4:0] _T_1630; // @[Modules.scala 143:103:@52705.4]
  wire [3:0] _T_1631; // @[Modules.scala 143:103:@52706.4]
  wire [3:0] _T_1632; // @[Modules.scala 143:103:@52707.4]
  wire [5:0] buffer_6_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_6_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1640; // @[Modules.scala 160:64:@52715.4]
  wire [5:0] _T_1641; // @[Modules.scala 160:64:@52716.4]
  wire [5:0] buffer_6_6; // @[Modules.scala 160:64:@52717.4]
  wire [5:0] buffer_6_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_6_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1643; // @[Modules.scala 160:64:@52719.4]
  wire [5:0] _T_1644; // @[Modules.scala 160:64:@52720.4]
  wire [5:0] buffer_6_7; // @[Modules.scala 160:64:@52721.4]
  wire [5:0] buffer_6_4; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1646; // @[Modules.scala 160:64:@52723.4]
  wire [5:0] _T_1647; // @[Modules.scala 160:64:@52724.4]
  wire [5:0] buffer_6_8; // @[Modules.scala 160:64:@52725.4]
  wire [6:0] _T_1649; // @[Modules.scala 166:64:@52727.4]
  wire [5:0] _T_1650; // @[Modules.scala 166:64:@52728.4]
  wire [5:0] buffer_6_9; // @[Modules.scala 166:64:@52729.4]
  wire [6:0] _T_1652; // @[Modules.scala 172:66:@52731.4]
  wire [5:0] _T_1653; // @[Modules.scala 172:66:@52732.4]
  wire [5:0] buffer_6_10; // @[Modules.scala 172:66:@52733.4]
  wire [4:0] _T_1659; // @[Modules.scala 150:103:@52742.4]
  wire [3:0] _T_1660; // @[Modules.scala 150:103:@52743.4]
  wire [3:0] _T_1661; // @[Modules.scala 150:103:@52744.4]
  wire [3:0] _GEN_24; // @[Modules.scala 150:103:@52748.4]
  wire [4:0] _T_1666; // @[Modules.scala 150:103:@52748.4]
  wire [3:0] _T_1667; // @[Modules.scala 150:103:@52749.4]
  wire [3:0] _T_1668; // @[Modules.scala 150:103:@52750.4]
  wire [4:0] _T_1673; // @[Modules.scala 150:103:@52754.4]
  wire [3:0] _T_1674; // @[Modules.scala 150:103:@52755.4]
  wire [3:0] _T_1675; // @[Modules.scala 150:103:@52756.4]
  wire [3:0] _GEN_25; // @[Modules.scala 150:103:@52760.4]
  wire [4:0] _T_1680; // @[Modules.scala 150:103:@52760.4]
  wire [3:0] _T_1681; // @[Modules.scala 150:103:@52761.4]
  wire [3:0] _T_1682; // @[Modules.scala 150:103:@52762.4]
  wire [4:0] _T_1694; // @[Modules.scala 150:103:@52772.4]
  wire [3:0] _T_1695; // @[Modules.scala 150:103:@52773.4]
  wire [3:0] _T_1696; // @[Modules.scala 150:103:@52774.4]
  wire [5:0] buffer_7_0; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_7_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1699; // @[Modules.scala 166:64:@52778.4]
  wire [5:0] _T_1700; // @[Modules.scala 166:64:@52779.4]
  wire [5:0] buffer_7_7; // @[Modules.scala 166:64:@52780.4]
  wire [5:0] buffer_7_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_7_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1702; // @[Modules.scala 166:64:@52782.4]
  wire [5:0] _T_1703; // @[Modules.scala 166:64:@52783.4]
  wire [5:0] buffer_7_8; // @[Modules.scala 166:64:@52784.4]
  wire [5:0] buffer_7_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1705; // @[Modules.scala 166:64:@52786.4]
  wire [5:0] _T_1706; // @[Modules.scala 166:64:@52787.4]
  wire [5:0] buffer_7_9; // @[Modules.scala 166:64:@52788.4]
  wire [6:0] _T_1708; // @[Modules.scala 166:64:@52790.4]
  wire [5:0] _T_1709; // @[Modules.scala 166:64:@52791.4]
  wire [5:0] buffer_7_10; // @[Modules.scala 166:64:@52792.4]
  wire [5:0] buffer_7_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1711; // @[Modules.scala 172:66:@52794.4]
  wire [5:0] _T_1712; // @[Modules.scala 172:66:@52795.4]
  wire [5:0] buffer_7_11; // @[Modules.scala 172:66:@52796.4]
  wire [6:0] _T_1714; // @[Modules.scala 160:64:@52798.4]
  wire [5:0] _T_1715; // @[Modules.scala 160:64:@52799.4]
  wire [5:0] buffer_7_12; // @[Modules.scala 160:64:@52800.4]
  wire [4:0] _T_1742; // @[Modules.scala 150:103:@52825.4]
  wire [3:0] _T_1743; // @[Modules.scala 150:103:@52826.4]
  wire [3:0] _T_1744; // @[Modules.scala 150:103:@52827.4]
  wire [4:0] _T_1756; // @[Modules.scala 150:103:@52837.4]
  wire [3:0] _T_1757; // @[Modules.scala 150:103:@52838.4]
  wire [3:0] _T_1758; // @[Modules.scala 150:103:@52839.4]
  wire [6:0] _T_1761; // @[Modules.scala 166:64:@52843.4]
  wire [5:0] _T_1762; // @[Modules.scala 166:64:@52844.4]
  wire [5:0] buffer_8_7; // @[Modules.scala 166:64:@52845.4]
  wire [5:0] buffer_8_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1764; // @[Modules.scala 166:64:@52847.4]
  wire [5:0] _T_1765; // @[Modules.scala 166:64:@52848.4]
  wire [5:0] buffer_8_8; // @[Modules.scala 166:64:@52849.4]
  wire [5:0] buffer_8_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1767; // @[Modules.scala 166:64:@52851.4]
  wire [5:0] _T_1768; // @[Modules.scala 166:64:@52852.4]
  wire [5:0] buffer_8_9; // @[Modules.scala 166:64:@52853.4]
  wire [6:0] _T_1770; // @[Modules.scala 166:64:@52855.4]
  wire [5:0] _T_1771; // @[Modules.scala 166:64:@52856.4]
  wire [5:0] buffer_8_10; // @[Modules.scala 166:64:@52857.4]
  wire [6:0] _T_1773; // @[Modules.scala 172:66:@52859.4]
  wire [5:0] _T_1774; // @[Modules.scala 172:66:@52860.4]
  wire [5:0] buffer_8_11; // @[Modules.scala 172:66:@52861.4]
  wire [6:0] _T_1776; // @[Modules.scala 160:64:@52863.4]
  wire [5:0] _T_1777; // @[Modules.scala 160:64:@52864.4]
  wire [5:0] buffer_8_12; // @[Modules.scala 160:64:@52865.4]
  wire [3:0] _T_1790; // @[Modules.scala 150:103:@52878.4]
  wire [2:0] _T_1791; // @[Modules.scala 150:103:@52879.4]
  wire [2:0] _T_1792; // @[Modules.scala 150:103:@52880.4]
  wire [4:0] _T_1811; // @[Modules.scala 150:103:@52896.4]
  wire [3:0] _T_1812; // @[Modules.scala 150:103:@52897.4]
  wire [3:0] _T_1813; // @[Modules.scala 150:103:@52898.4]
  wire [5:0] buffer_9_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1816; // @[Modules.scala 160:64:@52902.4]
  wire [5:0] _T_1817; // @[Modules.scala 160:64:@52903.4]
  wire [5:0] buffer_9_6; // @[Modules.scala 160:64:@52904.4]
  wire [6:0] _T_1819; // @[Modules.scala 160:64:@52906.4]
  wire [5:0] _T_1820; // @[Modules.scala 160:64:@52907.4]
  wire [5:0] buffer_9_7; // @[Modules.scala 160:64:@52908.4]
  wire [5:0] buffer_9_4; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1822; // @[Modules.scala 160:64:@52910.4]
  wire [5:0] _T_1823; // @[Modules.scala 160:64:@52911.4]
  wire [5:0] buffer_9_8; // @[Modules.scala 160:64:@52912.4]
  wire [6:0] _T_1825; // @[Modules.scala 166:64:@52914.4]
  wire [5:0] _T_1826; // @[Modules.scala 166:64:@52915.4]
  wire [5:0] buffer_9_9; // @[Modules.scala 166:64:@52916.4]
  wire [6:0] _T_1828; // @[Modules.scala 172:66:@52918.4]
  wire [5:0] _T_1829; // @[Modules.scala 172:66:@52919.4]
  wire [5:0] buffer_9_10; // @[Modules.scala 172:66:@52920.4]
  wire [4:0] _T_1849; // @[Modules.scala 150:103:@52941.4]
  wire [3:0] _T_1850; // @[Modules.scala 150:103:@52942.4]
  wire [3:0] _T_1851; // @[Modules.scala 150:103:@52943.4]
  wire [3:0] _T_1863; // @[Modules.scala 150:103:@52953.4]
  wire [2:0] _T_1864; // @[Modules.scala 150:103:@52954.4]
  wire [2:0] _T_1865; // @[Modules.scala 150:103:@52955.4]
  wire [4:0] _T_1870; // @[Modules.scala 150:103:@52959.4]
  wire [3:0] _T_1871; // @[Modules.scala 150:103:@52960.4]
  wire [3:0] _T_1872; // @[Modules.scala 150:103:@52961.4]
  wire [4:0] _T_1877; // @[Modules.scala 150:103:@52965.4]
  wire [3:0] _T_1878; // @[Modules.scala 150:103:@52966.4]
  wire [3:0] _T_1879; // @[Modules.scala 150:103:@52967.4]
  wire [6:0] _T_1882; // @[Modules.scala 160:64:@52971.4]
  wire [5:0] _T_1883; // @[Modules.scala 160:64:@52972.4]
  wire [5:0] buffer_10_8; // @[Modules.scala 160:64:@52973.4]
  wire [5:0] buffer_10_2; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1885; // @[Modules.scala 160:64:@52975.4]
  wire [5:0] _T_1886; // @[Modules.scala 160:64:@52976.4]
  wire [5:0] buffer_10_9; // @[Modules.scala 160:64:@52977.4]
  wire [5:0] buffer_10_4; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_10_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1888; // @[Modules.scala 160:64:@52979.4]
  wire [5:0] _T_1889; // @[Modules.scala 160:64:@52980.4]
  wire [5:0] buffer_10_10; // @[Modules.scala 160:64:@52981.4]
  wire [5:0] buffer_10_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1891; // @[Modules.scala 160:64:@52983.4]
  wire [5:0] _T_1892; // @[Modules.scala 160:64:@52984.4]
  wire [5:0] buffer_10_11; // @[Modules.scala 160:64:@52985.4]
  wire [6:0] _T_1894; // @[Modules.scala 160:64:@52987.4]
  wire [5:0] _T_1895; // @[Modules.scala 160:64:@52988.4]
  wire [5:0] buffer_10_12; // @[Modules.scala 160:64:@52989.4]
  wire [6:0] _T_1897; // @[Modules.scala 160:64:@52991.4]
  wire [5:0] _T_1898; // @[Modules.scala 160:64:@52992.4]
  wire [5:0] buffer_10_13; // @[Modules.scala 160:64:@52993.4]
  wire [6:0] _T_1900; // @[Modules.scala 160:64:@52995.4]
  wire [5:0] _T_1901; // @[Modules.scala 160:64:@52996.4]
  wire [5:0] buffer_10_14; // @[Modules.scala 160:64:@52997.4]
  wire [3:0] _T_1935; // @[Modules.scala 143:103:@53026.4]
  wire [2:0] _T_1936; // @[Modules.scala 143:103:@53027.4]
  wire [2:0] _T_1937; // @[Modules.scala 143:103:@53028.4]
  wire [6:0] _T_1952; // @[Modules.scala 166:64:@53042.4]
  wire [5:0] _T_1953; // @[Modules.scala 166:64:@53043.4]
  wire [5:0] buffer_11_7; // @[Modules.scala 166:64:@53044.4]
  wire [6:0] _T_1955; // @[Modules.scala 166:64:@53046.4]
  wire [5:0] _T_1956; // @[Modules.scala 166:64:@53047.4]
  wire [5:0] buffer_11_8; // @[Modules.scala 166:64:@53048.4]
  wire [5:0] buffer_11_4; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_1958; // @[Modules.scala 166:64:@53050.4]
  wire [5:0] _T_1959; // @[Modules.scala 166:64:@53051.4]
  wire [5:0] buffer_11_9; // @[Modules.scala 166:64:@53052.4]
  wire [6:0] _T_1961; // @[Modules.scala 166:64:@53054.4]
  wire [5:0] _T_1962; // @[Modules.scala 166:64:@53055.4]
  wire [5:0] buffer_11_10; // @[Modules.scala 166:64:@53056.4]
  wire [6:0] _T_1964; // @[Modules.scala 172:66:@53058.4]
  wire [5:0] _T_1965; // @[Modules.scala 172:66:@53059.4]
  wire [5:0] buffer_11_11; // @[Modules.scala 172:66:@53060.4]
  wire [6:0] _T_1967; // @[Modules.scala 160:64:@53062.4]
  wire [5:0] _T_1968; // @[Modules.scala 160:64:@53063.4]
  wire [5:0] buffer_11_12; // @[Modules.scala 160:64:@53064.4]
  wire [3:0] _T_2009; // @[Modules.scala 150:103:@53101.4]
  wire [2:0] _T_2010; // @[Modules.scala 150:103:@53102.4]
  wire [2:0] _T_2011; // @[Modules.scala 150:103:@53103.4]
  wire [6:0] _T_2017; // @[Modules.scala 166:64:@53111.4]
  wire [5:0] _T_2018; // @[Modules.scala 166:64:@53112.4]
  wire [5:0] buffer_12_8; // @[Modules.scala 166:64:@53113.4]
  wire [5:0] buffer_12_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2020; // @[Modules.scala 166:64:@53115.4]
  wire [5:0] _T_2021; // @[Modules.scala 166:64:@53116.4]
  wire [5:0] buffer_12_9; // @[Modules.scala 166:64:@53117.4]
  wire [6:0] _T_2023; // @[Modules.scala 166:64:@53119.4]
  wire [5:0] _T_2024; // @[Modules.scala 166:64:@53120.4]
  wire [5:0] buffer_12_10; // @[Modules.scala 166:64:@53121.4]
  wire [5:0] buffer_12_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2026; // @[Modules.scala 172:66:@53123.4]
  wire [5:0] _T_2027; // @[Modules.scala 172:66:@53124.4]
  wire [5:0] buffer_12_11; // @[Modules.scala 172:66:@53125.4]
  wire [6:0] _T_2029; // @[Modules.scala 160:64:@53127.4]
  wire [5:0] _T_2030; // @[Modules.scala 160:64:@53128.4]
  wire [5:0] buffer_12_12; // @[Modules.scala 160:64:@53129.4]
  wire [3:0] _T_2050; // @[Modules.scala 150:103:@53148.4]
  wire [2:0] _T_2051; // @[Modules.scala 150:103:@53149.4]
  wire [2:0] _T_2052; // @[Modules.scala 150:103:@53150.4]
  wire [4:0] _T_2064; // @[Modules.scala 150:103:@53160.4]
  wire [3:0] _T_2065; // @[Modules.scala 150:103:@53161.4]
  wire [3:0] _T_2066; // @[Modules.scala 150:103:@53162.4]
  wire [3:0] _T_2071; // @[Modules.scala 150:103:@53166.4]
  wire [2:0] _T_2072; // @[Modules.scala 150:103:@53167.4]
  wire [2:0] _T_2073; // @[Modules.scala 150:103:@53168.4]
  wire [6:0] _T_2076; // @[Modules.scala 166:64:@53172.4]
  wire [5:0] _T_2077; // @[Modules.scala 166:64:@53173.4]
  wire [5:0] buffer_13_7; // @[Modules.scala 166:64:@53174.4]
  wire [5:0] buffer_13_2; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2079; // @[Modules.scala 166:64:@53176.4]
  wire [5:0] _T_2080; // @[Modules.scala 166:64:@53177.4]
  wire [5:0] buffer_13_8; // @[Modules.scala 166:64:@53178.4]
  wire [5:0] buffer_13_4; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_13_5; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2082; // @[Modules.scala 166:64:@53180.4]
  wire [5:0] _T_2083; // @[Modules.scala 166:64:@53181.4]
  wire [5:0] buffer_13_9; // @[Modules.scala 166:64:@53182.4]
  wire [6:0] _T_2085; // @[Modules.scala 166:64:@53184.4]
  wire [5:0] _T_2086; // @[Modules.scala 166:64:@53185.4]
  wire [5:0] buffer_13_10; // @[Modules.scala 166:64:@53186.4]
  wire [6:0] _T_2088; // @[Modules.scala 172:66:@53188.4]
  wire [5:0] _T_2089; // @[Modules.scala 172:66:@53189.4]
  wire [5:0] buffer_13_11; // @[Modules.scala 172:66:@53190.4]
  wire [6:0] _T_2091; // @[Modules.scala 160:64:@53192.4]
  wire [5:0] _T_2092; // @[Modules.scala 160:64:@53193.4]
  wire [5:0] buffer_13_12; // @[Modules.scala 160:64:@53194.4]
  wire [4:0] _T_2112; // @[Modules.scala 143:103:@53213.4]
  wire [3:0] _T_2113; // @[Modules.scala 143:103:@53214.4]
  wire [3:0] _T_2114; // @[Modules.scala 143:103:@53215.4]
  wire [3:0] _T_2119; // @[Modules.scala 143:103:@53219.4]
  wire [2:0] _T_2120; // @[Modules.scala 143:103:@53220.4]
  wire [2:0] _T_2121; // @[Modules.scala 143:103:@53221.4]
  wire [4:0] _T_2126; // @[Modules.scala 143:103:@53225.4]
  wire [3:0] _T_2127; // @[Modules.scala 143:103:@53226.4]
  wire [3:0] _T_2128; // @[Modules.scala 143:103:@53227.4]
  wire [5:0] buffer_14_2; // @[Modules.scala 112:22:@52272.4]
  wire [5:0] buffer_14_3; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2139; // @[Modules.scala 160:64:@53239.4]
  wire [5:0] _T_2140; // @[Modules.scala 160:64:@53240.4]
  wire [5:0] buffer_14_7; // @[Modules.scala 160:64:@53241.4]
  wire [5:0] buffer_14_4; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2142; // @[Modules.scala 160:64:@53243.4]
  wire [5:0] _T_2143; // @[Modules.scala 160:64:@53244.4]
  wire [5:0] buffer_14_8; // @[Modules.scala 160:64:@53245.4]
  wire [6:0] _T_2145; // @[Modules.scala 166:64:@53247.4]
  wire [5:0] _T_2146; // @[Modules.scala 166:64:@53248.4]
  wire [5:0] buffer_14_9; // @[Modules.scala 166:64:@53249.4]
  wire [6:0] _T_2148; // @[Modules.scala 172:66:@53251.4]
  wire [5:0] _T_2149; // @[Modules.scala 172:66:@53252.4]
  wire [5:0] buffer_14_10; // @[Modules.scala 172:66:@53253.4]
  wire [4:0] _T_2162; // @[Modules.scala 150:103:@53268.4]
  wire [3:0] _T_2163; // @[Modules.scala 150:103:@53269.4]
  wire [3:0] _T_2164; // @[Modules.scala 150:103:@53270.4]
  wire [3:0] _T_2169; // @[Modules.scala 150:103:@53274.4]
  wire [2:0] _T_2170; // @[Modules.scala 150:103:@53275.4]
  wire [2:0] _T_2171; // @[Modules.scala 150:103:@53276.4]
  wire [5:0] buffer_15_1; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2195; // @[Modules.scala 166:64:@53298.4]
  wire [5:0] _T_2196; // @[Modules.scala 166:64:@53299.4]
  wire [5:0] buffer_15_7; // @[Modules.scala 166:64:@53300.4]
  wire [5:0] buffer_15_2; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2198; // @[Modules.scala 166:64:@53302.4]
  wire [5:0] _T_2199; // @[Modules.scala 166:64:@53303.4]
  wire [5:0] buffer_15_8; // @[Modules.scala 166:64:@53304.4]
  wire [6:0] _T_2201; // @[Modules.scala 166:64:@53306.4]
  wire [5:0] _T_2202; // @[Modules.scala 166:64:@53307.4]
  wire [5:0] buffer_15_9; // @[Modules.scala 166:64:@53308.4]
  wire [6:0] _T_2204; // @[Modules.scala 166:64:@53310.4]
  wire [5:0] _T_2205; // @[Modules.scala 166:64:@53311.4]
  wire [5:0] buffer_15_10; // @[Modules.scala 166:64:@53312.4]
  wire [5:0] buffer_15_6; // @[Modules.scala 112:22:@52272.4]
  wire [6:0] _T_2207; // @[Modules.scala 172:66:@53314.4]
  wire [5:0] _T_2208; // @[Modules.scala 172:66:@53315.4]
  wire [5:0] buffer_15_11; // @[Modules.scala 172:66:@53316.4]
  wire [6:0] _T_2210; // @[Modules.scala 160:64:@53318.4]
  wire [5:0] _T_2211; // @[Modules.scala 160:64:@53319.4]
  wire [5:0] buffer_15_12; // @[Modules.scala 160:64:@53320.4]
  assign _T_1207 = $signed(2'sh1) * $signed(io_in_0); // @[Modules.scala 143:74:@52273.4]
  assign _T_1209 = $signed(2'sh1) * $signed(io_in_1); // @[Modules.scala 144:80:@52274.4]
  assign _T_1210 = $signed(_T_1207) + $signed(_T_1209); // @[Modules.scala 143:103:@52275.4]
  assign _T_1211 = _T_1210[3:0]; // @[Modules.scala 143:103:@52276.4]
  assign _T_1212 = $signed(_T_1211); // @[Modules.scala 143:103:@52277.4]
  assign _T_1214 = $signed(2'sh1) * $signed(io_in_2); // @[Modules.scala 143:74:@52279.4]
  assign _T_1216 = $signed(2'sh1) * $signed(io_in_3); // @[Modules.scala 144:80:@52280.4]
  assign _T_1217 = $signed(_T_1214) + $signed(_T_1216); // @[Modules.scala 143:103:@52281.4]
  assign _T_1218 = _T_1217[3:0]; // @[Modules.scala 143:103:@52282.4]
  assign _T_1219 = $signed(_T_1218); // @[Modules.scala 143:103:@52283.4]
  assign _T_1221 = $signed(2'sh1) * $signed(io_in_4); // @[Modules.scala 143:74:@52285.4]
  assign _T_1223 = $signed(-2'sh1) * $signed(io_in_5); // @[Modules.scala 144:80:@52286.4]
  assign _GEN_0 = {{1{_T_1223[2]}},_T_1223}; // @[Modules.scala 143:103:@52287.4]
  assign _T_1224 = $signed(_T_1221) + $signed(_GEN_0); // @[Modules.scala 143:103:@52287.4]
  assign _T_1225 = _T_1224[3:0]; // @[Modules.scala 143:103:@52288.4]
  assign _T_1226 = $signed(_T_1225); // @[Modules.scala 143:103:@52289.4]
  assign _T_1228 = $signed(2'sh1) * $signed(io_in_7); // @[Modules.scala 143:74:@52291.4]
  assign _T_1230 = $signed(-2'sh1) * $signed(io_in_8); // @[Modules.scala 144:80:@52292.4]
  assign _GEN_1 = {{1{_T_1230[2]}},_T_1230}; // @[Modules.scala 143:103:@52293.4]
  assign _T_1231 = $signed(_T_1228) + $signed(_GEN_1); // @[Modules.scala 143:103:@52293.4]
  assign _T_1232 = _T_1231[3:0]; // @[Modules.scala 143:103:@52294.4]
  assign _T_1233 = $signed(_T_1232); // @[Modules.scala 143:103:@52295.4]
  assign _T_1235 = $signed(2'sh1) * $signed(io_in_9); // @[Modules.scala 143:74:@52297.4]
  assign _T_1237 = $signed(2'sh1) * $signed(io_in_10); // @[Modules.scala 144:80:@52298.4]
  assign _T_1238 = $signed(_T_1235) + $signed(_T_1237); // @[Modules.scala 143:103:@52299.4]
  assign _T_1239 = _T_1238[3:0]; // @[Modules.scala 143:103:@52300.4]
  assign _T_1240 = $signed(_T_1239); // @[Modules.scala 143:103:@52301.4]
  assign _T_1242 = $signed(2'sh1) * $signed(io_in_11); // @[Modules.scala 143:74:@52303.4]
  assign _T_1244 = $signed(-2'sh1) * $signed(io_in_12); // @[Modules.scala 144:80:@52304.4]
  assign _GEN_2 = {{1{_T_1244[2]}},_T_1244}; // @[Modules.scala 143:103:@52305.4]
  assign _T_1245 = $signed(_T_1242) + $signed(_GEN_2); // @[Modules.scala 143:103:@52305.4]
  assign _T_1246 = _T_1245[3:0]; // @[Modules.scala 143:103:@52306.4]
  assign _T_1247 = $signed(_T_1246); // @[Modules.scala 143:103:@52307.4]
  assign _T_1249 = $signed(-2'sh1) * $signed(io_in_14); // @[Modules.scala 143:74:@52309.4]
  assign _T_1251 = $signed(-2'sh1) * $signed(io_in_15); // @[Modules.scala 144:80:@52310.4]
  assign _T_1252 = $signed(_T_1249) + $signed(_T_1251); // @[Modules.scala 143:103:@52311.4]
  assign _T_1253 = _T_1252[2:0]; // @[Modules.scala 143:103:@52312.4]
  assign _T_1254 = $signed(_T_1253); // @[Modules.scala 143:103:@52313.4]
  assign buffer_0_0 = {{2{_T_1212[3]}},_T_1212}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_0_1 = {{2{_T_1219[3]}},_T_1219}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1255 = $signed(buffer_0_0) + $signed(buffer_0_1); // @[Modules.scala 166:64:@52315.4]
  assign _T_1256 = _T_1255[5:0]; // @[Modules.scala 166:64:@52316.4]
  assign buffer_0_7 = $signed(_T_1256); // @[Modules.scala 166:64:@52317.4]
  assign buffer_0_2 = {{2{_T_1226[3]}},_T_1226}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_0_3 = {{2{_T_1233[3]}},_T_1233}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1258 = $signed(buffer_0_2) + $signed(buffer_0_3); // @[Modules.scala 166:64:@52319.4]
  assign _T_1259 = _T_1258[5:0]; // @[Modules.scala 166:64:@52320.4]
  assign buffer_0_8 = $signed(_T_1259); // @[Modules.scala 166:64:@52321.4]
  assign buffer_0_4 = {{2{_T_1240[3]}},_T_1240}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_0_5 = {{2{_T_1247[3]}},_T_1247}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1261 = $signed(buffer_0_4) + $signed(buffer_0_5); // @[Modules.scala 166:64:@52323.4]
  assign _T_1262 = _T_1261[5:0]; // @[Modules.scala 166:64:@52324.4]
  assign buffer_0_9 = $signed(_T_1262); // @[Modules.scala 166:64:@52325.4]
  assign _T_1264 = $signed(buffer_0_7) + $signed(buffer_0_8); // @[Modules.scala 166:64:@52327.4]
  assign _T_1265 = _T_1264[5:0]; // @[Modules.scala 166:64:@52328.4]
  assign buffer_0_10 = $signed(_T_1265); // @[Modules.scala 166:64:@52329.4]
  assign buffer_0_6 = {{3{_T_1254[2]}},_T_1254}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1267 = $signed(buffer_0_9) + $signed(buffer_0_6); // @[Modules.scala 172:66:@52331.4]
  assign _T_1268 = _T_1267[5:0]; // @[Modules.scala 172:66:@52332.4]
  assign buffer_0_11 = $signed(_T_1268); // @[Modules.scala 172:66:@52333.4]
  assign _T_1270 = $signed(buffer_0_10) + $signed(buffer_0_11); // @[Modules.scala 160:64:@52335.4]
  assign _T_1271 = _T_1270[5:0]; // @[Modules.scala 160:64:@52336.4]
  assign buffer_0_12 = $signed(_T_1271); // @[Modules.scala 160:64:@52337.4]
  assign _T_1274 = $signed(-2'sh1) * $signed(io_in_1); // @[Modules.scala 143:74:@52342.4]
  assign _GEN_3 = {{1{_T_1274[2]}},_T_1274}; // @[Modules.scala 143:103:@52344.4]
  assign _T_1277 = $signed(_GEN_3) + $signed(_T_1214); // @[Modules.scala 143:103:@52344.4]
  assign _T_1278 = _T_1277[3:0]; // @[Modules.scala 143:103:@52345.4]
  assign _T_1279 = $signed(_T_1278); // @[Modules.scala 143:103:@52346.4]
  assign _T_1283 = $signed(-2'sh1) * $signed(io_in_4); // @[Modules.scala 144:80:@52349.4]
  assign _GEN_4 = {{1{_T_1283[2]}},_T_1283}; // @[Modules.scala 143:103:@52350.4]
  assign _T_1284 = $signed(_T_1216) + $signed(_GEN_4); // @[Modules.scala 143:103:@52350.4]
  assign _T_1285 = _T_1284[3:0]; // @[Modules.scala 143:103:@52351.4]
  assign _T_1286 = $signed(_T_1285); // @[Modules.scala 143:103:@52352.4]
  assign _T_1288 = $signed(2'sh1) * $signed(io_in_5); // @[Modules.scala 143:74:@52354.4]
  assign _T_1290 = $signed(-2'sh1) * $signed(io_in_6); // @[Modules.scala 144:80:@52355.4]
  assign _GEN_5 = {{1{_T_1290[2]}},_T_1290}; // @[Modules.scala 143:103:@52356.4]
  assign _T_1291 = $signed(_T_1288) + $signed(_GEN_5); // @[Modules.scala 143:103:@52356.4]
  assign _T_1292 = _T_1291[3:0]; // @[Modules.scala 143:103:@52357.4]
  assign _T_1293 = $signed(_T_1292); // @[Modules.scala 143:103:@52358.4]
  assign _T_1295 = $signed(-2'sh1) * $signed(io_in_7); // @[Modules.scala 143:74:@52360.4]
  assign _T_1298 = $signed(_T_1295) + $signed(_T_1230); // @[Modules.scala 143:103:@52362.4]
  assign _T_1299 = _T_1298[2:0]; // @[Modules.scala 143:103:@52363.4]
  assign _T_1300 = $signed(_T_1299); // @[Modules.scala 143:103:@52364.4]
  assign _T_1302 = $signed(-2'sh1) * $signed(io_in_9); // @[Modules.scala 143:74:@52366.4]
  assign _GEN_6 = {{1{_T_1302[2]}},_T_1302}; // @[Modules.scala 143:103:@52368.4]
  assign _T_1305 = $signed(_GEN_6) + $signed(_T_1237); // @[Modules.scala 143:103:@52368.4]
  assign _T_1306 = _T_1305[3:0]; // @[Modules.scala 143:103:@52369.4]
  assign _T_1307 = $signed(_T_1306); // @[Modules.scala 143:103:@52370.4]
  assign _T_1316 = $signed(2'sh1) * $signed(io_in_13); // @[Modules.scala 143:74:@52378.4]
  assign _GEN_8 = {{1{_T_1249[2]}},_T_1249}; // @[Modules.scala 143:103:@52380.4]
  assign _T_1319 = $signed(_T_1316) + $signed(_GEN_8); // @[Modules.scala 143:103:@52380.4]
  assign _T_1320 = _T_1319[3:0]; // @[Modules.scala 143:103:@52381.4]
  assign _T_1321 = $signed(_T_1320); // @[Modules.scala 143:103:@52382.4]
  assign buffer_1_0 = {{2{_T_1279[3]}},_T_1279}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_1_1 = {{2{_T_1286[3]}},_T_1286}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1322 = $signed(buffer_1_0) + $signed(buffer_1_1); // @[Modules.scala 166:64:@52384.4]
  assign _T_1323 = _T_1322[5:0]; // @[Modules.scala 166:64:@52385.4]
  assign buffer_1_7 = $signed(_T_1323); // @[Modules.scala 166:64:@52386.4]
  assign buffer_1_2 = {{2{_T_1293[3]}},_T_1293}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_1_3 = {{3{_T_1300[2]}},_T_1300}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1325 = $signed(buffer_1_2) + $signed(buffer_1_3); // @[Modules.scala 166:64:@52388.4]
  assign _T_1326 = _T_1325[5:0]; // @[Modules.scala 166:64:@52389.4]
  assign buffer_1_8 = $signed(_T_1326); // @[Modules.scala 166:64:@52390.4]
  assign buffer_1_4 = {{2{_T_1307[3]}},_T_1307}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1328 = $signed(buffer_1_4) + $signed(buffer_0_5); // @[Modules.scala 166:64:@52392.4]
  assign _T_1329 = _T_1328[5:0]; // @[Modules.scala 166:64:@52393.4]
  assign buffer_1_9 = $signed(_T_1329); // @[Modules.scala 166:64:@52394.4]
  assign _T_1331 = $signed(buffer_1_7) + $signed(buffer_1_8); // @[Modules.scala 166:64:@52396.4]
  assign _T_1332 = _T_1331[5:0]; // @[Modules.scala 166:64:@52397.4]
  assign buffer_1_10 = $signed(_T_1332); // @[Modules.scala 166:64:@52398.4]
  assign buffer_1_6 = {{2{_T_1321[3]}},_T_1321}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1334 = $signed(buffer_1_9) + $signed(buffer_1_6); // @[Modules.scala 172:66:@52400.4]
  assign _T_1335 = _T_1334[5:0]; // @[Modules.scala 172:66:@52401.4]
  assign buffer_1_11 = $signed(_T_1335); // @[Modules.scala 172:66:@52402.4]
  assign _T_1337 = $signed(buffer_1_10) + $signed(buffer_1_11); // @[Modules.scala 160:64:@52404.4]
  assign _T_1338 = _T_1337[5:0]; // @[Modules.scala 160:64:@52405.4]
  assign buffer_1_12 = $signed(_T_1338); // @[Modules.scala 160:64:@52406.4]
  assign _T_1344 = $signed(_T_1207) + $signed(_GEN_3); // @[Modules.scala 150:103:@52413.4]
  assign _T_1345 = _T_1344[3:0]; // @[Modules.scala 150:103:@52414.4]
  assign _T_1346 = $signed(_T_1345); // @[Modules.scala 150:103:@52415.4]
  assign _T_1351 = $signed(_T_1216) + $signed(_GEN_0); // @[Modules.scala 150:103:@52419.4]
  assign _T_1352 = _T_1351[3:0]; // @[Modules.scala 150:103:@52420.4]
  assign _T_1353 = $signed(_T_1352); // @[Modules.scala 150:103:@52421.4]
  assign _T_1358 = $signed(_GEN_5) + $signed(_T_1228); // @[Modules.scala 150:103:@52425.4]
  assign _T_1359 = _T_1358[3:0]; // @[Modules.scala 150:103:@52426.4]
  assign _T_1360 = $signed(_T_1359); // @[Modules.scala 150:103:@52427.4]
  assign _T_1362 = $signed(2'sh1) * $signed(io_in_8); // @[Modules.scala 150:74:@52429.4]
  assign _T_1365 = $signed(_T_1362) + $signed(_T_1235); // @[Modules.scala 150:103:@52431.4]
  assign _T_1366 = _T_1365[3:0]; // @[Modules.scala 150:103:@52432.4]
  assign _T_1367 = $signed(_T_1366); // @[Modules.scala 150:103:@52433.4]
  assign _T_1371 = $signed(-2'sh1) * $signed(io_in_11); // @[Modules.scala 151:80:@52436.4]
  assign _GEN_12 = {{1{_T_1371[2]}},_T_1371}; // @[Modules.scala 150:103:@52437.4]
  assign _T_1372 = $signed(_T_1237) + $signed(_GEN_12); // @[Modules.scala 150:103:@52437.4]
  assign _T_1373 = _T_1372[3:0]; // @[Modules.scala 150:103:@52438.4]
  assign _T_1374 = $signed(_T_1373); // @[Modules.scala 150:103:@52439.4]
  assign _T_1376 = $signed(2'sh1) * $signed(io_in_12); // @[Modules.scala 150:74:@52441.4]
  assign _T_1378 = $signed(2'sh1) * $signed(io_in_14); // @[Modules.scala 151:80:@52442.4]
  assign _T_1379 = $signed(_T_1376) + $signed(_T_1378); // @[Modules.scala 150:103:@52443.4]
  assign _T_1380 = _T_1379[3:0]; // @[Modules.scala 150:103:@52444.4]
  assign _T_1381 = $signed(_T_1380); // @[Modules.scala 150:103:@52445.4]
  assign _T_1383 = $signed(2'sh1) * $signed(io_in_15); // @[Modules.scala 153:80:@52447.4]
  assign buffer_2_0 = {{2{_T_1346[3]}},_T_1346}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_2_1 = {{2{_T_1353[3]}},_T_1353}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1384 = $signed(buffer_2_0) + $signed(buffer_2_1); // @[Modules.scala 166:64:@52449.4]
  assign _T_1385 = _T_1384[5:0]; // @[Modules.scala 166:64:@52450.4]
  assign buffer_2_7 = $signed(_T_1385); // @[Modules.scala 166:64:@52451.4]
  assign buffer_2_2 = {{2{_T_1360[3]}},_T_1360}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_2_3 = {{2{_T_1367[3]}},_T_1367}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1387 = $signed(buffer_2_2) + $signed(buffer_2_3); // @[Modules.scala 166:64:@52453.4]
  assign _T_1388 = _T_1387[5:0]; // @[Modules.scala 166:64:@52454.4]
  assign buffer_2_8 = $signed(_T_1388); // @[Modules.scala 166:64:@52455.4]
  assign buffer_2_4 = {{2{_T_1374[3]}},_T_1374}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_2_5 = {{2{_T_1381[3]}},_T_1381}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1390 = $signed(buffer_2_4) + $signed(buffer_2_5); // @[Modules.scala 166:64:@52457.4]
  assign _T_1391 = _T_1390[5:0]; // @[Modules.scala 166:64:@52458.4]
  assign buffer_2_9 = $signed(_T_1391); // @[Modules.scala 166:64:@52459.4]
  assign _T_1393 = $signed(buffer_2_7) + $signed(buffer_2_8); // @[Modules.scala 166:64:@52461.4]
  assign _T_1394 = _T_1393[5:0]; // @[Modules.scala 166:64:@52462.4]
  assign buffer_2_10 = $signed(_T_1394); // @[Modules.scala 166:64:@52463.4]
  assign buffer_2_6 = {{2{_T_1383[3]}},_T_1383}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1396 = $signed(buffer_2_9) + $signed(buffer_2_6); // @[Modules.scala 172:66:@52465.4]
  assign _T_1397 = _T_1396[5:0]; // @[Modules.scala 172:66:@52466.4]
  assign buffer_2_11 = $signed(_T_1397); // @[Modules.scala 172:66:@52467.4]
  assign _T_1399 = $signed(buffer_2_10) + $signed(buffer_2_11); // @[Modules.scala 160:64:@52469.4]
  assign _T_1400 = _T_1399[5:0]; // @[Modules.scala 160:64:@52470.4]
  assign buffer_2_12 = $signed(_T_1400); // @[Modules.scala 160:64:@52471.4]
  assign _T_1405 = $signed(-2'sh1) * $signed(io_in_2); // @[Modules.scala 144:80:@52477.4]
  assign _GEN_13 = {{1{_T_1405[2]}},_T_1405}; // @[Modules.scala 143:103:@52478.4]
  assign _T_1406 = $signed(_T_1207) + $signed(_GEN_13); // @[Modules.scala 143:103:@52478.4]
  assign _T_1407 = _T_1406[3:0]; // @[Modules.scala 143:103:@52479.4]
  assign _T_1408 = $signed(_T_1407); // @[Modules.scala 143:103:@52480.4]
  assign _T_1413 = $signed(_GEN_4) + $signed(_T_1288); // @[Modules.scala 143:103:@52484.4]
  assign _T_1414 = _T_1413[3:0]; // @[Modules.scala 143:103:@52485.4]
  assign _T_1415 = $signed(_T_1414); // @[Modules.scala 143:103:@52486.4]
  assign _T_1417 = $signed(2'sh1) * $signed(io_in_6); // @[Modules.scala 143:74:@52488.4]
  assign _T_1420 = $signed(_T_1417) + $signed(_T_1228); // @[Modules.scala 143:103:@52490.4]
  assign _T_1421 = _T_1420[3:0]; // @[Modules.scala 143:103:@52491.4]
  assign _T_1422 = $signed(_T_1421); // @[Modules.scala 143:103:@52492.4]
  assign _T_1434 = $signed(_T_1242) + $signed(_T_1376); // @[Modules.scala 143:103:@52502.4]
  assign _T_1435 = _T_1434[3:0]; // @[Modules.scala 143:103:@52503.4]
  assign _T_1436 = $signed(_T_1435); // @[Modules.scala 143:103:@52504.4]
  assign _T_1441 = $signed(_T_1378) + $signed(_T_1383); // @[Modules.scala 143:103:@52508.4]
  assign _T_1442 = _T_1441[3:0]; // @[Modules.scala 143:103:@52509.4]
  assign _T_1443 = $signed(_T_1442); // @[Modules.scala 143:103:@52510.4]
  assign buffer_3_0 = {{2{_T_1408[3]}},_T_1408}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_3_1 = {{2{_T_1415[3]}},_T_1415}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1444 = $signed(buffer_3_0) + $signed(buffer_3_1); // @[Modules.scala 160:64:@52512.4]
  assign _T_1445 = _T_1444[5:0]; // @[Modules.scala 160:64:@52513.4]
  assign buffer_3_6 = $signed(_T_1445); // @[Modules.scala 160:64:@52514.4]
  assign buffer_3_2 = {{2{_T_1422[3]}},_T_1422}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1447 = $signed(buffer_3_2) + $signed(buffer_2_3); // @[Modules.scala 160:64:@52516.4]
  assign _T_1448 = _T_1447[5:0]; // @[Modules.scala 160:64:@52517.4]
  assign buffer_3_7 = $signed(_T_1448); // @[Modules.scala 160:64:@52518.4]
  assign buffer_3_4 = {{2{_T_1436[3]}},_T_1436}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_3_5 = {{2{_T_1443[3]}},_T_1443}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1450 = $signed(buffer_3_4) + $signed(buffer_3_5); // @[Modules.scala 160:64:@52520.4]
  assign _T_1451 = _T_1450[5:0]; // @[Modules.scala 160:64:@52521.4]
  assign buffer_3_8 = $signed(_T_1451); // @[Modules.scala 160:64:@52522.4]
  assign _T_1453 = $signed(buffer_3_6) + $signed(buffer_3_7); // @[Modules.scala 166:64:@52524.4]
  assign _T_1454 = _T_1453[5:0]; // @[Modules.scala 166:64:@52525.4]
  assign buffer_3_9 = $signed(_T_1454); // @[Modules.scala 166:64:@52526.4]
  assign _T_1456 = $signed(buffer_3_9) + $signed(buffer_3_8); // @[Modules.scala 172:66:@52528.4]
  assign _T_1457 = _T_1456[5:0]; // @[Modules.scala 172:66:@52529.4]
  assign buffer_3_10 = $signed(_T_1457); // @[Modules.scala 172:66:@52530.4]
  assign _T_1460 = $signed(-2'sh1) * $signed(io_in_0); // @[Modules.scala 143:74:@52537.4]
  assign _GEN_15 = {{1{_T_1460[2]}},_T_1460}; // @[Modules.scala 143:103:@52539.4]
  assign _T_1463 = $signed(_GEN_15) + $signed(_T_1209); // @[Modules.scala 143:103:@52539.4]
  assign _T_1464 = _T_1463[3:0]; // @[Modules.scala 143:103:@52540.4]
  assign _T_1465 = $signed(_T_1464); // @[Modules.scala 143:103:@52541.4]
  assign _T_1470 = $signed(_T_1216) + $signed(_T_1288); // @[Modules.scala 143:103:@52545.4]
  assign _T_1471 = _T_1470[3:0]; // @[Modules.scala 143:103:@52546.4]
  assign _T_1472 = $signed(_T_1471); // @[Modules.scala 143:103:@52547.4]
  assign _T_1477 = $signed(_T_1290) + $signed(_T_1295); // @[Modules.scala 143:103:@52551.4]
  assign _T_1478 = _T_1477[2:0]; // @[Modules.scala 143:103:@52552.4]
  assign _T_1479 = $signed(_T_1478); // @[Modules.scala 143:103:@52553.4]
  assign _T_1484 = $signed(_T_1362) + $signed(_GEN_6); // @[Modules.scala 143:103:@52557.4]
  assign _T_1485 = _T_1484[3:0]; // @[Modules.scala 143:103:@52558.4]
  assign _T_1486 = $signed(_T_1485); // @[Modules.scala 143:103:@52559.4]
  assign _T_1491 = $signed(_T_1237) + $signed(_T_1242); // @[Modules.scala 143:103:@52563.4]
  assign _T_1492 = _T_1491[3:0]; // @[Modules.scala 143:103:@52564.4]
  assign _T_1493 = $signed(_T_1492); // @[Modules.scala 143:103:@52565.4]
  assign _T_1497 = $signed(-2'sh1) * $signed(io_in_13); // @[Modules.scala 144:80:@52568.4]
  assign _GEN_17 = {{1{_T_1497[2]}},_T_1497}; // @[Modules.scala 143:103:@52569.4]
  assign _T_1498 = $signed(_T_1376) + $signed(_GEN_17); // @[Modules.scala 143:103:@52569.4]
  assign _T_1499 = _T_1498[3:0]; // @[Modules.scala 143:103:@52570.4]
  assign _T_1500 = $signed(_T_1499); // @[Modules.scala 143:103:@52571.4]
  assign buffer_4_0 = {{2{_T_1465[3]}},_T_1465}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_4_1 = {{2{_T_1472[3]}},_T_1472}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1508 = $signed(buffer_4_0) + $signed(buffer_4_1); // @[Modules.scala 166:64:@52579.4]
  assign _T_1509 = _T_1508[5:0]; // @[Modules.scala 166:64:@52580.4]
  assign buffer_4_7 = $signed(_T_1509); // @[Modules.scala 166:64:@52581.4]
  assign buffer_4_2 = {{3{_T_1479[2]}},_T_1479}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_4_3 = {{2{_T_1486[3]}},_T_1486}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1511 = $signed(buffer_4_2) + $signed(buffer_4_3); // @[Modules.scala 166:64:@52583.4]
  assign _T_1512 = _T_1511[5:0]; // @[Modules.scala 166:64:@52584.4]
  assign buffer_4_8 = $signed(_T_1512); // @[Modules.scala 166:64:@52585.4]
  assign buffer_4_4 = {{2{_T_1493[3]}},_T_1493}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_4_5 = {{2{_T_1500[3]}},_T_1500}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1514 = $signed(buffer_4_4) + $signed(buffer_4_5); // @[Modules.scala 166:64:@52587.4]
  assign _T_1515 = _T_1514[5:0]; // @[Modules.scala 166:64:@52588.4]
  assign buffer_4_9 = $signed(_T_1515); // @[Modules.scala 166:64:@52589.4]
  assign _T_1517 = $signed(buffer_4_7) + $signed(buffer_4_8); // @[Modules.scala 166:64:@52591.4]
  assign _T_1518 = _T_1517[5:0]; // @[Modules.scala 166:64:@52592.4]
  assign buffer_4_10 = $signed(_T_1518); // @[Modules.scala 166:64:@52593.4]
  assign _T_1520 = $signed(buffer_4_9) + $signed(buffer_3_5); // @[Modules.scala 172:66:@52595.4]
  assign _T_1521 = _T_1520[5:0]; // @[Modules.scala 172:66:@52596.4]
  assign buffer_4_11 = $signed(_T_1521); // @[Modules.scala 172:66:@52597.4]
  assign _T_1523 = $signed(buffer_4_10) + $signed(buffer_4_11); // @[Modules.scala 160:64:@52599.4]
  assign _T_1524 = _T_1523[5:0]; // @[Modules.scala 160:64:@52600.4]
  assign buffer_4_12 = $signed(_T_1524); // @[Modules.scala 160:64:@52601.4]
  assign _T_1530 = $signed(_T_1207) + $signed(_T_1214); // @[Modules.scala 150:103:@52608.4]
  assign _T_1531 = _T_1530[3:0]; // @[Modules.scala 150:103:@52609.4]
  assign _T_1532 = $signed(_T_1531); // @[Modules.scala 150:103:@52610.4]
  assign _T_1534 = $signed(-2'sh1) * $signed(io_in_3); // @[Modules.scala 150:74:@52612.4]
  assign _T_1537 = $signed(_T_1534) + $signed(_T_1283); // @[Modules.scala 150:103:@52614.4]
  assign _T_1538 = _T_1537[2:0]; // @[Modules.scala 150:103:@52615.4]
  assign _T_1539 = $signed(_T_1538); // @[Modules.scala 150:103:@52616.4]
  assign _T_1544 = $signed(_GEN_0) + $signed(_T_1417); // @[Modules.scala 150:103:@52620.4]
  assign _T_1545 = _T_1544[3:0]; // @[Modules.scala 150:103:@52621.4]
  assign _T_1546 = $signed(_T_1545); // @[Modules.scala 150:103:@52622.4]
  assign _T_1557 = $signed(-2'sh1) * $signed(io_in_10); // @[Modules.scala 151:80:@52631.4]
  assign _GEN_19 = {{1{_T_1557[2]}},_T_1557}; // @[Modules.scala 150:103:@52632.4]
  assign _T_1558 = $signed(_T_1235) + $signed(_GEN_19); // @[Modules.scala 150:103:@52632.4]
  assign _T_1559 = _T_1558[3:0]; // @[Modules.scala 150:103:@52633.4]
  assign _T_1560 = $signed(_T_1559); // @[Modules.scala 150:103:@52634.4]
  assign buffer_5_0 = {{2{_T_1532[3]}},_T_1532}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_5_1 = {{3{_T_1539[2]}},_T_1539}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1577 = $signed(buffer_5_0) + $signed(buffer_5_1); // @[Modules.scala 160:64:@52650.4]
  assign _T_1578 = _T_1577[5:0]; // @[Modules.scala 160:64:@52651.4]
  assign buffer_5_8 = $signed(_T_1578); // @[Modules.scala 160:64:@52652.4]
  assign buffer_5_2 = {{2{_T_1546[3]}},_T_1546}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1580 = $signed(buffer_5_2) + $signed(buffer_1_3); // @[Modules.scala 160:64:@52654.4]
  assign _T_1581 = _T_1580[5:0]; // @[Modules.scala 160:64:@52655.4]
  assign buffer_5_9 = $signed(_T_1581); // @[Modules.scala 160:64:@52656.4]
  assign buffer_5_4 = {{2{_T_1560[3]}},_T_1560}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1583 = $signed(buffer_5_4) + $signed(buffer_3_4); // @[Modules.scala 160:64:@52658.4]
  assign _T_1584 = _T_1583[5:0]; // @[Modules.scala 160:64:@52659.4]
  assign buffer_5_10 = $signed(_T_1584); // @[Modules.scala 160:64:@52660.4]
  assign _T_1586 = $signed(buffer_1_6) + $signed(buffer_2_6); // @[Modules.scala 160:64:@52662.4]
  assign _T_1587 = _T_1586[5:0]; // @[Modules.scala 160:64:@52663.4]
  assign buffer_5_11 = $signed(_T_1587); // @[Modules.scala 160:64:@52664.4]
  assign _T_1589 = $signed(buffer_5_8) + $signed(buffer_5_9); // @[Modules.scala 160:64:@52666.4]
  assign _T_1590 = _T_1589[5:0]; // @[Modules.scala 160:64:@52667.4]
  assign buffer_5_12 = $signed(_T_1590); // @[Modules.scala 160:64:@52668.4]
  assign _T_1592 = $signed(buffer_5_10) + $signed(buffer_5_11); // @[Modules.scala 160:64:@52670.4]
  assign _T_1593 = _T_1592[5:0]; // @[Modules.scala 160:64:@52671.4]
  assign buffer_5_13 = $signed(_T_1593); // @[Modules.scala 160:64:@52672.4]
  assign _T_1595 = $signed(buffer_5_12) + $signed(buffer_5_13); // @[Modules.scala 160:64:@52674.4]
  assign _T_1596 = _T_1595[5:0]; // @[Modules.scala 160:64:@52675.4]
  assign buffer_5_14 = $signed(_T_1596); // @[Modules.scala 160:64:@52676.4]
  assign _T_1602 = $signed(_T_1460) + $signed(_T_1274); // @[Modules.scala 143:103:@52681.4]
  assign _T_1603 = _T_1602[2:0]; // @[Modules.scala 143:103:@52682.4]
  assign _T_1604 = $signed(_T_1603); // @[Modules.scala 143:103:@52683.4]
  assign _T_1609 = $signed(_T_1214) + $signed(_T_1288); // @[Modules.scala 143:103:@52687.4]
  assign _T_1610 = _T_1609[3:0]; // @[Modules.scala 143:103:@52688.4]
  assign _T_1611 = $signed(_T_1610); // @[Modules.scala 143:103:@52689.4]
  assign _T_1616 = $signed(_T_1228) + $signed(_T_1362); // @[Modules.scala 143:103:@52693.4]
  assign _T_1617 = _T_1616[3:0]; // @[Modules.scala 143:103:@52694.4]
  assign _T_1618 = $signed(_T_1617); // @[Modules.scala 143:103:@52695.4]
  assign _T_1623 = $signed(_GEN_6) + $signed(_T_1242); // @[Modules.scala 143:103:@52699.4]
  assign _T_1624 = _T_1623[3:0]; // @[Modules.scala 143:103:@52700.4]
  assign _T_1625 = $signed(_T_1624); // @[Modules.scala 143:103:@52701.4]
  assign _T_1630 = $signed(_GEN_2) + $signed(_T_1316); // @[Modules.scala 143:103:@52705.4]
  assign _T_1631 = _T_1630[3:0]; // @[Modules.scala 143:103:@52706.4]
  assign _T_1632 = $signed(_T_1631); // @[Modules.scala 143:103:@52707.4]
  assign buffer_6_0 = {{3{_T_1604[2]}},_T_1604}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_6_1 = {{2{_T_1611[3]}},_T_1611}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1640 = $signed(buffer_6_0) + $signed(buffer_6_1); // @[Modules.scala 160:64:@52715.4]
  assign _T_1641 = _T_1640[5:0]; // @[Modules.scala 160:64:@52716.4]
  assign buffer_6_6 = $signed(_T_1641); // @[Modules.scala 160:64:@52717.4]
  assign buffer_6_2 = {{2{_T_1618[3]}},_T_1618}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_6_3 = {{2{_T_1625[3]}},_T_1625}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1643 = $signed(buffer_6_2) + $signed(buffer_6_3); // @[Modules.scala 160:64:@52719.4]
  assign _T_1644 = _T_1643[5:0]; // @[Modules.scala 160:64:@52720.4]
  assign buffer_6_7 = $signed(_T_1644); // @[Modules.scala 160:64:@52721.4]
  assign buffer_6_4 = {{2{_T_1632[3]}},_T_1632}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1646 = $signed(buffer_6_4) + $signed(buffer_0_6); // @[Modules.scala 160:64:@52723.4]
  assign _T_1647 = _T_1646[5:0]; // @[Modules.scala 160:64:@52724.4]
  assign buffer_6_8 = $signed(_T_1647); // @[Modules.scala 160:64:@52725.4]
  assign _T_1649 = $signed(buffer_6_6) + $signed(buffer_6_7); // @[Modules.scala 166:64:@52727.4]
  assign _T_1650 = _T_1649[5:0]; // @[Modules.scala 166:64:@52728.4]
  assign buffer_6_9 = $signed(_T_1650); // @[Modules.scala 166:64:@52729.4]
  assign _T_1652 = $signed(buffer_6_9) + $signed(buffer_6_8); // @[Modules.scala 172:66:@52731.4]
  assign _T_1653 = _T_1652[5:0]; // @[Modules.scala 172:66:@52732.4]
  assign buffer_6_10 = $signed(_T_1653); // @[Modules.scala 172:66:@52733.4]
  assign _T_1659 = $signed(_GEN_15) + $signed(_T_1214); // @[Modules.scala 150:103:@52742.4]
  assign _T_1660 = _T_1659[3:0]; // @[Modules.scala 150:103:@52743.4]
  assign _T_1661 = $signed(_T_1660); // @[Modules.scala 150:103:@52744.4]
  assign _GEN_24 = {{1{_T_1534[2]}},_T_1534}; // @[Modules.scala 150:103:@52748.4]
  assign _T_1666 = $signed(_GEN_24) + $signed(_T_1221); // @[Modules.scala 150:103:@52748.4]
  assign _T_1667 = _T_1666[3:0]; // @[Modules.scala 150:103:@52749.4]
  assign _T_1668 = $signed(_T_1667); // @[Modules.scala 150:103:@52750.4]
  assign _T_1673 = $signed(_T_1288) + $signed(_T_1417); // @[Modules.scala 150:103:@52754.4]
  assign _T_1674 = _T_1673[3:0]; // @[Modules.scala 150:103:@52755.4]
  assign _T_1675 = $signed(_T_1674); // @[Modules.scala 150:103:@52756.4]
  assign _GEN_25 = {{1{_T_1295[2]}},_T_1295}; // @[Modules.scala 150:103:@52760.4]
  assign _T_1680 = $signed(_GEN_25) + $signed(_T_1362); // @[Modules.scala 150:103:@52760.4]
  assign _T_1681 = _T_1680[3:0]; // @[Modules.scala 150:103:@52761.4]
  assign _T_1682 = $signed(_T_1681); // @[Modules.scala 150:103:@52762.4]
  assign _T_1694 = $signed(_T_1376) + $signed(_GEN_8); // @[Modules.scala 150:103:@52772.4]
  assign _T_1695 = _T_1694[3:0]; // @[Modules.scala 150:103:@52773.4]
  assign _T_1696 = $signed(_T_1695); // @[Modules.scala 150:103:@52774.4]
  assign buffer_7_0 = {{2{_T_1661[3]}},_T_1661}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_7_1 = {{2{_T_1668[3]}},_T_1668}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1699 = $signed(buffer_7_0) + $signed(buffer_7_1); // @[Modules.scala 166:64:@52778.4]
  assign _T_1700 = _T_1699[5:0]; // @[Modules.scala 166:64:@52779.4]
  assign buffer_7_7 = $signed(_T_1700); // @[Modules.scala 166:64:@52780.4]
  assign buffer_7_2 = {{2{_T_1675[3]}},_T_1675}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_7_3 = {{2{_T_1682[3]}},_T_1682}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1702 = $signed(buffer_7_2) + $signed(buffer_7_3); // @[Modules.scala 166:64:@52782.4]
  assign _T_1703 = _T_1702[5:0]; // @[Modules.scala 166:64:@52783.4]
  assign buffer_7_8 = $signed(_T_1703); // @[Modules.scala 166:64:@52784.4]
  assign buffer_7_5 = {{2{_T_1696[3]}},_T_1696}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1705 = $signed(buffer_5_4) + $signed(buffer_7_5); // @[Modules.scala 166:64:@52786.4]
  assign _T_1706 = _T_1705[5:0]; // @[Modules.scala 166:64:@52787.4]
  assign buffer_7_9 = $signed(_T_1706); // @[Modules.scala 166:64:@52788.4]
  assign _T_1708 = $signed(buffer_7_7) + $signed(buffer_7_8); // @[Modules.scala 166:64:@52790.4]
  assign _T_1709 = _T_1708[5:0]; // @[Modules.scala 166:64:@52791.4]
  assign buffer_7_10 = $signed(_T_1709); // @[Modules.scala 166:64:@52792.4]
  assign buffer_7_6 = {{3{_T_1251[2]}},_T_1251}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1711 = $signed(buffer_7_9) + $signed(buffer_7_6); // @[Modules.scala 172:66:@52794.4]
  assign _T_1712 = _T_1711[5:0]; // @[Modules.scala 172:66:@52795.4]
  assign buffer_7_11 = $signed(_T_1712); // @[Modules.scala 172:66:@52796.4]
  assign _T_1714 = $signed(buffer_7_10) + $signed(buffer_7_11); // @[Modules.scala 160:64:@52798.4]
  assign _T_1715 = _T_1714[5:0]; // @[Modules.scala 160:64:@52799.4]
  assign buffer_7_12 = $signed(_T_1715); // @[Modules.scala 160:64:@52800.4]
  assign _T_1742 = $signed(_GEN_1) + $signed(_T_1235); // @[Modules.scala 150:103:@52825.4]
  assign _T_1743 = _T_1742[3:0]; // @[Modules.scala 150:103:@52826.4]
  assign _T_1744 = $signed(_T_1743); // @[Modules.scala 150:103:@52827.4]
  assign _T_1756 = $signed(_T_1316) + $signed(_T_1378); // @[Modules.scala 150:103:@52837.4]
  assign _T_1757 = _T_1756[3:0]; // @[Modules.scala 150:103:@52838.4]
  assign _T_1758 = $signed(_T_1757); // @[Modules.scala 150:103:@52839.4]
  assign _T_1761 = $signed(buffer_0_0) + $signed(buffer_7_1); // @[Modules.scala 166:64:@52843.4]
  assign _T_1762 = _T_1761[5:0]; // @[Modules.scala 166:64:@52844.4]
  assign buffer_8_7 = $signed(_T_1762); // @[Modules.scala 166:64:@52845.4]
  assign buffer_8_3 = {{2{_T_1744[3]}},_T_1744}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1764 = $signed(buffer_5_2) + $signed(buffer_8_3); // @[Modules.scala 166:64:@52847.4]
  assign _T_1765 = _T_1764[5:0]; // @[Modules.scala 166:64:@52848.4]
  assign buffer_8_8 = $signed(_T_1765); // @[Modules.scala 166:64:@52849.4]
  assign buffer_8_5 = {{2{_T_1758[3]}},_T_1758}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1767 = $signed(buffer_4_4) + $signed(buffer_8_5); // @[Modules.scala 166:64:@52851.4]
  assign _T_1768 = _T_1767[5:0]; // @[Modules.scala 166:64:@52852.4]
  assign buffer_8_9 = $signed(_T_1768); // @[Modules.scala 166:64:@52853.4]
  assign _T_1770 = $signed(buffer_8_7) + $signed(buffer_8_8); // @[Modules.scala 166:64:@52855.4]
  assign _T_1771 = _T_1770[5:0]; // @[Modules.scala 166:64:@52856.4]
  assign buffer_8_10 = $signed(_T_1771); // @[Modules.scala 166:64:@52857.4]
  assign _T_1773 = $signed(buffer_8_9) + $signed(buffer_2_6); // @[Modules.scala 172:66:@52859.4]
  assign _T_1774 = _T_1773[5:0]; // @[Modules.scala 172:66:@52860.4]
  assign buffer_8_11 = $signed(_T_1774); // @[Modules.scala 172:66:@52861.4]
  assign _T_1776 = $signed(buffer_8_10) + $signed(buffer_8_11); // @[Modules.scala 160:64:@52863.4]
  assign _T_1777 = _T_1776[5:0]; // @[Modules.scala 160:64:@52864.4]
  assign buffer_8_12 = $signed(_T_1777); // @[Modules.scala 160:64:@52865.4]
  assign _T_1790 = $signed(_T_1405) + $signed(_T_1534); // @[Modules.scala 150:103:@52878.4]
  assign _T_1791 = _T_1790[2:0]; // @[Modules.scala 150:103:@52879.4]
  assign _T_1792 = $signed(_T_1791); // @[Modules.scala 150:103:@52880.4]
  assign _T_1811 = $signed(_GEN_12) + $signed(_T_1378); // @[Modules.scala 150:103:@52896.4]
  assign _T_1812 = _T_1811[3:0]; // @[Modules.scala 150:103:@52897.4]
  assign _T_1813 = $signed(_T_1812); // @[Modules.scala 150:103:@52898.4]
  assign buffer_9_1 = {{3{_T_1792[2]}},_T_1792}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1816 = $signed(buffer_2_0) + $signed(buffer_9_1); // @[Modules.scala 160:64:@52902.4]
  assign _T_1817 = _T_1816[5:0]; // @[Modules.scala 160:64:@52903.4]
  assign buffer_9_6 = $signed(_T_1817); // @[Modules.scala 160:64:@52904.4]
  assign _T_1819 = $signed(buffer_3_1) + $signed(buffer_1_3); // @[Modules.scala 160:64:@52906.4]
  assign _T_1820 = _T_1819[5:0]; // @[Modules.scala 160:64:@52907.4]
  assign buffer_9_7 = $signed(_T_1820); // @[Modules.scala 160:64:@52908.4]
  assign buffer_9_4 = {{2{_T_1813[3]}},_T_1813}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1822 = $signed(buffer_9_4) + $signed(buffer_2_6); // @[Modules.scala 160:64:@52910.4]
  assign _T_1823 = _T_1822[5:0]; // @[Modules.scala 160:64:@52911.4]
  assign buffer_9_8 = $signed(_T_1823); // @[Modules.scala 160:64:@52912.4]
  assign _T_1825 = $signed(buffer_9_6) + $signed(buffer_9_7); // @[Modules.scala 166:64:@52914.4]
  assign _T_1826 = _T_1825[5:0]; // @[Modules.scala 166:64:@52915.4]
  assign buffer_9_9 = $signed(_T_1826); // @[Modules.scala 166:64:@52916.4]
  assign _T_1828 = $signed(buffer_9_9) + $signed(buffer_9_8); // @[Modules.scala 172:66:@52918.4]
  assign _T_1829 = _T_1828[5:0]; // @[Modules.scala 172:66:@52919.4]
  assign buffer_9_10 = $signed(_T_1829); // @[Modules.scala 172:66:@52920.4]
  assign _T_1849 = $signed(_T_1221) + $signed(_T_1288); // @[Modules.scala 150:103:@52941.4]
  assign _T_1850 = _T_1849[3:0]; // @[Modules.scala 150:103:@52942.4]
  assign _T_1851 = $signed(_T_1850); // @[Modules.scala 150:103:@52943.4]
  assign _T_1863 = $signed(_T_1302) + $signed(_T_1557); // @[Modules.scala 150:103:@52953.4]
  assign _T_1864 = _T_1863[2:0]; // @[Modules.scala 150:103:@52954.4]
  assign _T_1865 = $signed(_T_1864); // @[Modules.scala 150:103:@52955.4]
  assign _T_1870 = $signed(_GEN_12) + $signed(_T_1376); // @[Modules.scala 150:103:@52959.4]
  assign _T_1871 = _T_1870[3:0]; // @[Modules.scala 150:103:@52960.4]
  assign _T_1872 = $signed(_T_1871); // @[Modules.scala 150:103:@52961.4]
  assign _T_1877 = $signed(_GEN_17) + $signed(_T_1378); // @[Modules.scala 150:103:@52965.4]
  assign _T_1878 = _T_1877[3:0]; // @[Modules.scala 150:103:@52966.4]
  assign _T_1879 = $signed(_T_1878); // @[Modules.scala 150:103:@52967.4]
  assign _T_1882 = $signed(buffer_4_0) + $signed(buffer_9_1); // @[Modules.scala 160:64:@52971.4]
  assign _T_1883 = _T_1882[5:0]; // @[Modules.scala 160:64:@52972.4]
  assign buffer_10_8 = $signed(_T_1883); // @[Modules.scala 160:64:@52973.4]
  assign buffer_10_2 = {{2{_T_1851[3]}},_T_1851}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1885 = $signed(buffer_10_2) + $signed(buffer_7_3); // @[Modules.scala 160:64:@52975.4]
  assign _T_1886 = _T_1885[5:0]; // @[Modules.scala 160:64:@52976.4]
  assign buffer_10_9 = $signed(_T_1886); // @[Modules.scala 160:64:@52977.4]
  assign buffer_10_4 = {{3{_T_1865[2]}},_T_1865}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_10_5 = {{2{_T_1872[3]}},_T_1872}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1888 = $signed(buffer_10_4) + $signed(buffer_10_5); // @[Modules.scala 160:64:@52979.4]
  assign _T_1889 = _T_1888[5:0]; // @[Modules.scala 160:64:@52980.4]
  assign buffer_10_10 = $signed(_T_1889); // @[Modules.scala 160:64:@52981.4]
  assign buffer_10_6 = {{2{_T_1879[3]}},_T_1879}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1891 = $signed(buffer_10_6) + $signed(buffer_7_6); // @[Modules.scala 160:64:@52983.4]
  assign _T_1892 = _T_1891[5:0]; // @[Modules.scala 160:64:@52984.4]
  assign buffer_10_11 = $signed(_T_1892); // @[Modules.scala 160:64:@52985.4]
  assign _T_1894 = $signed(buffer_10_8) + $signed(buffer_10_9); // @[Modules.scala 160:64:@52987.4]
  assign _T_1895 = _T_1894[5:0]; // @[Modules.scala 160:64:@52988.4]
  assign buffer_10_12 = $signed(_T_1895); // @[Modules.scala 160:64:@52989.4]
  assign _T_1897 = $signed(buffer_10_10) + $signed(buffer_10_11); // @[Modules.scala 160:64:@52991.4]
  assign _T_1898 = _T_1897[5:0]; // @[Modules.scala 160:64:@52992.4]
  assign buffer_10_13 = $signed(_T_1898); // @[Modules.scala 160:64:@52993.4]
  assign _T_1900 = $signed(buffer_10_12) + $signed(buffer_10_13); // @[Modules.scala 160:64:@52995.4]
  assign _T_1901 = _T_1900[5:0]; // @[Modules.scala 160:64:@52996.4]
  assign buffer_10_14 = $signed(_T_1901); // @[Modules.scala 160:64:@52997.4]
  assign _T_1935 = $signed(_T_1557) + $signed(_T_1371); // @[Modules.scala 143:103:@53026.4]
  assign _T_1936 = _T_1935[2:0]; // @[Modules.scala 143:103:@53027.4]
  assign _T_1937 = $signed(_T_1936); // @[Modules.scala 143:103:@53028.4]
  assign _T_1952 = $signed(buffer_2_0) + $signed(buffer_0_1); // @[Modules.scala 166:64:@53042.4]
  assign _T_1953 = _T_1952[5:0]; // @[Modules.scala 166:64:@53043.4]
  assign buffer_11_7 = $signed(_T_1953); // @[Modules.scala 166:64:@53044.4]
  assign _T_1955 = $signed(buffer_0_2) + $signed(buffer_2_3); // @[Modules.scala 166:64:@53046.4]
  assign _T_1956 = _T_1955[5:0]; // @[Modules.scala 166:64:@53047.4]
  assign buffer_11_8 = $signed(_T_1956); // @[Modules.scala 166:64:@53048.4]
  assign buffer_11_4 = {{3{_T_1937[2]}},_T_1937}; // @[Modules.scala 112:22:@52272.4]
  assign _T_1958 = $signed(buffer_11_4) + $signed(buffer_4_5); // @[Modules.scala 166:64:@53050.4]
  assign _T_1959 = _T_1958[5:0]; // @[Modules.scala 166:64:@53051.4]
  assign buffer_11_9 = $signed(_T_1959); // @[Modules.scala 166:64:@53052.4]
  assign _T_1961 = $signed(buffer_11_7) + $signed(buffer_11_8); // @[Modules.scala 166:64:@53054.4]
  assign _T_1962 = _T_1961[5:0]; // @[Modules.scala 166:64:@53055.4]
  assign buffer_11_10 = $signed(_T_1962); // @[Modules.scala 166:64:@53056.4]
  assign _T_1964 = $signed(buffer_11_9) + $signed(buffer_0_6); // @[Modules.scala 172:66:@53058.4]
  assign _T_1965 = _T_1964[5:0]; // @[Modules.scala 172:66:@53059.4]
  assign buffer_11_11 = $signed(_T_1965); // @[Modules.scala 172:66:@53060.4]
  assign _T_1967 = $signed(buffer_11_10) + $signed(buffer_11_11); // @[Modules.scala 160:64:@53062.4]
  assign _T_1968 = _T_1967[5:0]; // @[Modules.scala 160:64:@53063.4]
  assign buffer_11_12 = $signed(_T_1968); // @[Modules.scala 160:64:@53064.4]
  assign _T_2009 = $signed(_T_1371) + $signed(_T_1244); // @[Modules.scala 150:103:@53101.4]
  assign _T_2010 = _T_2009[2:0]; // @[Modules.scala 150:103:@53102.4]
  assign _T_2011 = $signed(_T_2010); // @[Modules.scala 150:103:@53103.4]
  assign _T_2017 = $signed(buffer_7_2) + $signed(buffer_0_3); // @[Modules.scala 166:64:@53111.4]
  assign _T_2018 = _T_2017[5:0]; // @[Modules.scala 166:64:@53112.4]
  assign buffer_12_8 = $signed(_T_2018); // @[Modules.scala 166:64:@53113.4]
  assign buffer_12_5 = {{3{_T_2011[2]}},_T_2011}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2020 = $signed(buffer_10_4) + $signed(buffer_12_5); // @[Modules.scala 166:64:@53115.4]
  assign _T_2021 = _T_2020[5:0]; // @[Modules.scala 166:64:@53116.4]
  assign buffer_12_9 = $signed(_T_2021); // @[Modules.scala 166:64:@53117.4]
  assign _T_2023 = $signed(buffer_9_6) + $signed(buffer_12_8); // @[Modules.scala 166:64:@53119.4]
  assign _T_2024 = _T_2023[5:0]; // @[Modules.scala 166:64:@53120.4]
  assign buffer_12_10 = $signed(_T_2024); // @[Modules.scala 166:64:@53121.4]
  assign buffer_12_6 = {{3{_T_1497[2]}},_T_1497}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2026 = $signed(buffer_12_9) + $signed(buffer_12_6); // @[Modules.scala 172:66:@53123.4]
  assign _T_2027 = _T_2026[5:0]; // @[Modules.scala 172:66:@53124.4]
  assign buffer_12_11 = $signed(_T_2027); // @[Modules.scala 172:66:@53125.4]
  assign _T_2029 = $signed(buffer_12_10) + $signed(buffer_12_11); // @[Modules.scala 160:64:@53127.4]
  assign _T_2030 = _T_2029[5:0]; // @[Modules.scala 160:64:@53128.4]
  assign buffer_12_12 = $signed(_T_2030); // @[Modules.scala 160:64:@53129.4]
  assign _T_2050 = $signed(_T_1283) + $signed(_T_1290); // @[Modules.scala 150:103:@53148.4]
  assign _T_2051 = _T_2050[2:0]; // @[Modules.scala 150:103:@53149.4]
  assign _T_2052 = $signed(_T_2051); // @[Modules.scala 150:103:@53150.4]
  assign _T_2064 = $signed(_T_1235) + $signed(_GEN_12); // @[Modules.scala 150:103:@53160.4]
  assign _T_2065 = _T_2064[3:0]; // @[Modules.scala 150:103:@53161.4]
  assign _T_2066 = $signed(_T_2065); // @[Modules.scala 150:103:@53162.4]
  assign _T_2071 = $signed(_T_1497) + $signed(_T_1249); // @[Modules.scala 150:103:@53166.4]
  assign _T_2072 = _T_2071[2:0]; // @[Modules.scala 150:103:@53167.4]
  assign _T_2073 = $signed(_T_2072); // @[Modules.scala 150:103:@53168.4]
  assign _T_2076 = $signed(buffer_6_0) + $signed(buffer_0_1); // @[Modules.scala 166:64:@53172.4]
  assign _T_2077 = _T_2076[5:0]; // @[Modules.scala 166:64:@53173.4]
  assign buffer_13_7 = $signed(_T_2077); // @[Modules.scala 166:64:@53174.4]
  assign buffer_13_2 = {{3{_T_2052[2]}},_T_2052}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2079 = $signed(buffer_13_2) + $signed(buffer_1_3); // @[Modules.scala 166:64:@53176.4]
  assign _T_2080 = _T_2079[5:0]; // @[Modules.scala 166:64:@53177.4]
  assign buffer_13_8 = $signed(_T_2080); // @[Modules.scala 166:64:@53178.4]
  assign buffer_13_4 = {{2{_T_2066[3]}},_T_2066}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_13_5 = {{3{_T_2073[2]}},_T_2073}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2082 = $signed(buffer_13_4) + $signed(buffer_13_5); // @[Modules.scala 166:64:@53180.4]
  assign _T_2083 = _T_2082[5:0]; // @[Modules.scala 166:64:@53181.4]
  assign buffer_13_9 = $signed(_T_2083); // @[Modules.scala 166:64:@53182.4]
  assign _T_2085 = $signed(buffer_13_7) + $signed(buffer_13_8); // @[Modules.scala 166:64:@53184.4]
  assign _T_2086 = _T_2085[5:0]; // @[Modules.scala 166:64:@53185.4]
  assign buffer_13_10 = $signed(_T_2086); // @[Modules.scala 166:64:@53186.4]
  assign _T_2088 = $signed(buffer_13_9) + $signed(buffer_7_6); // @[Modules.scala 172:66:@53188.4]
  assign _T_2089 = _T_2088[5:0]; // @[Modules.scala 172:66:@53189.4]
  assign buffer_13_11 = $signed(_T_2089); // @[Modules.scala 172:66:@53190.4]
  assign _T_2091 = $signed(buffer_13_10) + $signed(buffer_13_11); // @[Modules.scala 160:64:@53192.4]
  assign _T_2092 = _T_2091[5:0]; // @[Modules.scala 160:64:@53193.4]
  assign buffer_13_12 = $signed(_T_2092); // @[Modules.scala 160:64:@53194.4]
  assign _T_2112 = $signed(_T_1288) + $signed(_GEN_25); // @[Modules.scala 143:103:@53213.4]
  assign _T_2113 = _T_2112[3:0]; // @[Modules.scala 143:103:@53214.4]
  assign _T_2114 = $signed(_T_2113); // @[Modules.scala 143:103:@53215.4]
  assign _T_2119 = $signed(_T_1230) + $signed(_T_1302); // @[Modules.scala 143:103:@53219.4]
  assign _T_2120 = _T_2119[2:0]; // @[Modules.scala 143:103:@53220.4]
  assign _T_2121 = $signed(_T_2120); // @[Modules.scala 143:103:@53221.4]
  assign _T_2126 = $signed(_T_1237) + $signed(_GEN_2); // @[Modules.scala 143:103:@53225.4]
  assign _T_2127 = _T_2126[3:0]; // @[Modules.scala 143:103:@53226.4]
  assign _T_2128 = $signed(_T_2127); // @[Modules.scala 143:103:@53227.4]
  assign buffer_14_2 = {{2{_T_2114[3]}},_T_2114}; // @[Modules.scala 112:22:@52272.4]
  assign buffer_14_3 = {{3{_T_2121[2]}},_T_2121}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2139 = $signed(buffer_14_2) + $signed(buffer_14_3); // @[Modules.scala 160:64:@53239.4]
  assign _T_2140 = _T_2139[5:0]; // @[Modules.scala 160:64:@53240.4]
  assign buffer_14_7 = $signed(_T_2140); // @[Modules.scala 160:64:@53241.4]
  assign buffer_14_4 = {{2{_T_2128[3]}},_T_2128}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2142 = $signed(buffer_14_4) + $signed(buffer_13_5); // @[Modules.scala 160:64:@53243.4]
  assign _T_2143 = _T_2142[5:0]; // @[Modules.scala 160:64:@53244.4]
  assign buffer_14_8 = $signed(_T_2143); // @[Modules.scala 160:64:@53245.4]
  assign _T_2145 = $signed(buffer_8_7) + $signed(buffer_14_7); // @[Modules.scala 166:64:@53247.4]
  assign _T_2146 = _T_2145[5:0]; // @[Modules.scala 166:64:@53248.4]
  assign buffer_14_9 = $signed(_T_2146); // @[Modules.scala 166:64:@53249.4]
  assign _T_2148 = $signed(buffer_14_9) + $signed(buffer_14_8); // @[Modules.scala 172:66:@53251.4]
  assign _T_2149 = _T_2148[5:0]; // @[Modules.scala 172:66:@53252.4]
  assign buffer_14_10 = $signed(_T_2149); // @[Modules.scala 172:66:@53253.4]
  assign _T_2162 = $signed(_T_1214) + $signed(_GEN_4); // @[Modules.scala 150:103:@53268.4]
  assign _T_2163 = _T_2162[3:0]; // @[Modules.scala 150:103:@53269.4]
  assign _T_2164 = $signed(_T_2163); // @[Modules.scala 150:103:@53270.4]
  assign _T_2169 = $signed(_T_1223) + $signed(_T_1290); // @[Modules.scala 150:103:@53274.4]
  assign _T_2170 = _T_2169[2:0]; // @[Modules.scala 150:103:@53275.4]
  assign _T_2171 = $signed(_T_2170); // @[Modules.scala 150:103:@53276.4]
  assign buffer_15_1 = {{2{_T_2164[3]}},_T_2164}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2195 = $signed(buffer_6_0) + $signed(buffer_15_1); // @[Modules.scala 166:64:@53298.4]
  assign _T_2196 = _T_2195[5:0]; // @[Modules.scala 166:64:@53299.4]
  assign buffer_15_7 = $signed(_T_2196); // @[Modules.scala 166:64:@53300.4]
  assign buffer_15_2 = {{3{_T_2171[2]}},_T_2171}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2198 = $signed(buffer_15_2) + $signed(buffer_8_3); // @[Modules.scala 166:64:@53302.4]
  assign _T_2199 = _T_2198[5:0]; // @[Modules.scala 166:64:@53303.4]
  assign buffer_15_8 = $signed(_T_2199); // @[Modules.scala 166:64:@53304.4]
  assign _T_2201 = $signed(buffer_11_4) + $signed(buffer_6_4); // @[Modules.scala 166:64:@53306.4]
  assign _T_2202 = _T_2201[5:0]; // @[Modules.scala 166:64:@53307.4]
  assign buffer_15_9 = $signed(_T_2202); // @[Modules.scala 166:64:@53308.4]
  assign _T_2204 = $signed(buffer_15_7) + $signed(buffer_15_8); // @[Modules.scala 166:64:@53310.4]
  assign _T_2205 = _T_2204[5:0]; // @[Modules.scala 166:64:@53311.4]
  assign buffer_15_10 = $signed(_T_2205); // @[Modules.scala 166:64:@53312.4]
  assign buffer_15_6 = {{2{_T_1378[3]}},_T_1378}; // @[Modules.scala 112:22:@52272.4]
  assign _T_2207 = $signed(buffer_15_9) + $signed(buffer_15_6); // @[Modules.scala 172:66:@53314.4]
  assign _T_2208 = _T_2207[5:0]; // @[Modules.scala 172:66:@53315.4]
  assign buffer_15_11 = $signed(_T_2208); // @[Modules.scala 172:66:@53316.4]
  assign _T_2210 = $signed(buffer_15_10) + $signed(buffer_15_11); // @[Modules.scala 160:64:@53318.4]
  assign _T_2211 = _T_2210[5:0]; // @[Modules.scala 160:64:@53319.4]
  assign buffer_15_12 = $signed(_T_2211); // @[Modules.scala 160:64:@53320.4]
  assign io_out_0 = buffer_0_12;
  assign io_out_1 = buffer_1_12;
  assign io_out_2 = buffer_2_12;
  assign io_out_3 = buffer_3_10;
  assign io_out_4 = buffer_4_12;
  assign io_out_5 = buffer_5_14;
  assign io_out_6 = buffer_6_10;
  assign io_out_7 = buffer_7_12;
  assign io_out_8 = buffer_8_12;
  assign io_out_9 = buffer_9_10;
  assign io_out_10 = buffer_10_14;
  assign io_out_11 = buffer_11_12;
  assign io_out_12 = buffer_12_12;
  assign io_out_13 = buffer_13_12;
  assign io_out_14 = buffer_14_10;
  assign io_out_15 = buffer_15_12;
endmodule
module BN_BI_1( // @[:@53612.2]
  input  [5:0] io_in_0, // @[:@53615.4]
  input  [5:0] io_in_1, // @[:@53615.4]
  input  [5:0] io_in_2, // @[:@53615.4]
  input  [5:0] io_in_3, // @[:@53615.4]
  input  [5:0] io_in_4, // @[:@53615.4]
  input  [5:0] io_in_5, // @[:@53615.4]
  input  [5:0] io_in_6, // @[:@53615.4]
  input  [5:0] io_in_7, // @[:@53615.4]
  input  [5:0] io_in_8, // @[:@53615.4]
  input  [5:0] io_in_9, // @[:@53615.4]
  input  [5:0] io_in_10, // @[:@53615.4]
  input  [5:0] io_in_11, // @[:@53615.4]
  input  [5:0] io_in_12, // @[:@53615.4]
  input  [5:0] io_in_13, // @[:@53615.4]
  input  [5:0] io_in_14, // @[:@53615.4]
  input  [5:0] io_in_15, // @[:@53615.4]
  output [5:0] io_out_0, // @[:@53615.4]
  output [5:0] io_out_1, // @[:@53615.4]
  output [5:0] io_out_2, // @[:@53615.4]
  output [5:0] io_out_3, // @[:@53615.4]
  output [5:0] io_out_4, // @[:@53615.4]
  output [5:0] io_out_5, // @[:@53615.4]
  output [5:0] io_out_6, // @[:@53615.4]
  output [5:0] io_out_7, // @[:@53615.4]
  output [5:0] io_out_8, // @[:@53615.4]
  output [5:0] io_out_9, // @[:@53615.4]
  output [5:0] io_out_10, // @[:@53615.4]
  output [5:0] io_out_11, // @[:@53615.4]
  output [5:0] io_out_12, // @[:@53615.4]
  output [5:0] io_out_13, // @[:@53615.4]
  output [5:0] io_out_14, // @[:@53615.4]
  output [5:0] io_out_15 // @[:@53615.4]
);
  wire [6:0] _T_66; // @[Modules.scala 282:31:@53618.4]
  wire [5:0] _T_67; // @[Modules.scala 282:31:@53619.4]
  wire [5:0] buffer_0; // @[Modules.scala 282:31:@53620.4]
  wire  _T_70; // @[Modules.scala 283:24:@53622.4]
  wire [1:0] _GEN_0; // @[Modules.scala 283:32:@53623.4]
  wire [6:0] _T_74; // @[Modules.scala 282:31:@53629.4]
  wire [5:0] _T_75; // @[Modules.scala 282:31:@53630.4]
  wire [5:0] buffer_1; // @[Modules.scala 282:31:@53631.4]
  wire  _T_78; // @[Modules.scala 283:24:@53633.4]
  wire [1:0] _GEN_1; // @[Modules.scala 283:32:@53634.4]
  wire [6:0] _T_82; // @[Modules.scala 282:31:@53640.4]
  wire [5:0] _T_83; // @[Modules.scala 282:31:@53641.4]
  wire [5:0] buffer_2; // @[Modules.scala 282:31:@53642.4]
  wire  _T_86; // @[Modules.scala 283:24:@53644.4]
  wire [1:0] _GEN_2; // @[Modules.scala 283:32:@53645.4]
  wire [6:0] _T_90; // @[Modules.scala 282:31:@53651.4]
  wire [5:0] _T_91; // @[Modules.scala 282:31:@53652.4]
  wire [5:0] buffer_3; // @[Modules.scala 282:31:@53653.4]
  wire  _T_94; // @[Modules.scala 283:24:@53655.4]
  wire [1:0] _GEN_3; // @[Modules.scala 283:32:@53656.4]
  wire [6:0] _T_98; // @[Modules.scala 282:31:@53662.4]
  wire [5:0] _T_99; // @[Modules.scala 282:31:@53663.4]
  wire [5:0] buffer_4; // @[Modules.scala 282:31:@53664.4]
  wire  _T_102; // @[Modules.scala 283:24:@53666.4]
  wire [1:0] _GEN_4; // @[Modules.scala 283:32:@53667.4]
  wire [6:0] _T_106; // @[Modules.scala 282:31:@53673.4]
  wire [5:0] _T_107; // @[Modules.scala 282:31:@53674.4]
  wire [5:0] buffer_5; // @[Modules.scala 282:31:@53675.4]
  wire  _T_110; // @[Modules.scala 283:24:@53677.4]
  wire [1:0] _GEN_5; // @[Modules.scala 283:32:@53678.4]
  wire [6:0] _T_114; // @[Modules.scala 282:31:@53684.4]
  wire [5:0] _T_115; // @[Modules.scala 282:31:@53685.4]
  wire [5:0] buffer_6; // @[Modules.scala 282:31:@53686.4]
  wire  _T_118; // @[Modules.scala 283:24:@53688.4]
  wire [1:0] _GEN_6; // @[Modules.scala 283:32:@53689.4]
  wire [6:0] _T_122; // @[Modules.scala 282:31:@53695.4]
  wire [5:0] _T_123; // @[Modules.scala 282:31:@53696.4]
  wire [5:0] buffer_7; // @[Modules.scala 282:31:@53697.4]
  wire  _T_126; // @[Modules.scala 283:24:@53699.4]
  wire [1:0] _GEN_7; // @[Modules.scala 283:32:@53700.4]
  wire [6:0] _T_130; // @[Modules.scala 282:31:@53706.4]
  wire [5:0] _T_131; // @[Modules.scala 282:31:@53707.4]
  wire [5:0] buffer_8; // @[Modules.scala 282:31:@53708.4]
  wire  _T_134; // @[Modules.scala 283:24:@53710.4]
  wire [1:0] _GEN_8; // @[Modules.scala 283:32:@53711.4]
  wire [6:0] _T_138; // @[Modules.scala 282:31:@53717.4]
  wire [5:0] _T_139; // @[Modules.scala 282:31:@53718.4]
  wire [5:0] buffer_9; // @[Modules.scala 282:31:@53719.4]
  wire  _T_142; // @[Modules.scala 283:24:@53721.4]
  wire [1:0] _GEN_9; // @[Modules.scala 283:32:@53722.4]
  wire [6:0] _T_146; // @[Modules.scala 282:31:@53728.4]
  wire [5:0] _T_147; // @[Modules.scala 282:31:@53729.4]
  wire [5:0] buffer_10; // @[Modules.scala 282:31:@53730.4]
  wire  _T_150; // @[Modules.scala 283:24:@53732.4]
  wire [1:0] _GEN_10; // @[Modules.scala 283:32:@53733.4]
  wire [6:0] _T_154; // @[Modules.scala 282:31:@53739.4]
  wire [5:0] _T_155; // @[Modules.scala 282:31:@53740.4]
  wire [5:0] buffer_11; // @[Modules.scala 282:31:@53741.4]
  wire  _T_158; // @[Modules.scala 283:24:@53743.4]
  wire [1:0] _GEN_11; // @[Modules.scala 283:32:@53744.4]
  wire [6:0] _T_162; // @[Modules.scala 282:31:@53750.4]
  wire [5:0] _T_163; // @[Modules.scala 282:31:@53751.4]
  wire [5:0] buffer_12; // @[Modules.scala 282:31:@53752.4]
  wire  _T_166; // @[Modules.scala 283:24:@53754.4]
  wire [1:0] _GEN_12; // @[Modules.scala 283:32:@53755.4]
  wire [6:0] _T_170; // @[Modules.scala 282:31:@53761.4]
  wire [5:0] _T_171; // @[Modules.scala 282:31:@53762.4]
  wire [5:0] buffer_13; // @[Modules.scala 282:31:@53763.4]
  wire  _T_174; // @[Modules.scala 283:24:@53765.4]
  wire [1:0] _GEN_13; // @[Modules.scala 283:32:@53766.4]
  wire [6:0] _T_178; // @[Modules.scala 282:31:@53772.4]
  wire [5:0] _T_179; // @[Modules.scala 282:31:@53773.4]
  wire [5:0] buffer_14; // @[Modules.scala 282:31:@53774.4]
  wire  _T_182; // @[Modules.scala 283:24:@53776.4]
  wire [1:0] _GEN_14; // @[Modules.scala 283:32:@53777.4]
  wire [6:0] _T_186; // @[Modules.scala 282:31:@53783.4]
  wire [5:0] _T_187; // @[Modules.scala 282:31:@53784.4]
  wire [5:0] buffer_15; // @[Modules.scala 282:31:@53785.4]
  wire  _T_190; // @[Modules.scala 283:24:@53787.4]
  wire [1:0] _GEN_15; // @[Modules.scala 283:32:@53788.4]
  assign _T_66 = $signed(io_in_0) - $signed(-6'sh3); // @[Modules.scala 282:31:@53618.4]
  assign _T_67 = _T_66[5:0]; // @[Modules.scala 282:31:@53619.4]
  assign buffer_0 = $signed(_T_67); // @[Modules.scala 282:31:@53620.4]
  assign _T_70 = $signed(buffer_0) >= $signed(6'sh0); // @[Modules.scala 283:24:@53622.4]
  assign _GEN_0 = _T_70 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53623.4]
  assign _T_74 = $signed(io_in_1) - $signed(6'sh1); // @[Modules.scala 282:31:@53629.4]
  assign _T_75 = _T_74[5:0]; // @[Modules.scala 282:31:@53630.4]
  assign buffer_1 = $signed(_T_75); // @[Modules.scala 282:31:@53631.4]
  assign _T_78 = $signed(buffer_1) >= $signed(6'sh0); // @[Modules.scala 283:24:@53633.4]
  assign _GEN_1 = _T_78 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53634.4]
  assign _T_82 = $signed(io_in_2) - $signed(6'sh1); // @[Modules.scala 282:31:@53640.4]
  assign _T_83 = _T_82[5:0]; // @[Modules.scala 282:31:@53641.4]
  assign buffer_2 = $signed(_T_83); // @[Modules.scala 282:31:@53642.4]
  assign _T_86 = $signed(buffer_2) >= $signed(6'sh0); // @[Modules.scala 283:24:@53644.4]
  assign _GEN_2 = _T_86 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53645.4]
  assign _T_90 = $signed(io_in_3) - $signed(6'sh1); // @[Modules.scala 282:31:@53651.4]
  assign _T_91 = _T_90[5:0]; // @[Modules.scala 282:31:@53652.4]
  assign buffer_3 = $signed(_T_91); // @[Modules.scala 282:31:@53653.4]
  assign _T_94 = $signed(buffer_3) >= $signed(6'sh0); // @[Modules.scala 283:24:@53655.4]
  assign _GEN_3 = _T_94 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53656.4]
  assign _T_98 = $signed(io_in_4) - $signed(6'sh1); // @[Modules.scala 282:31:@53662.4]
  assign _T_99 = _T_98[5:0]; // @[Modules.scala 282:31:@53663.4]
  assign buffer_4 = $signed(_T_99); // @[Modules.scala 282:31:@53664.4]
  assign _T_102 = $signed(buffer_4) >= $signed(6'sh0); // @[Modules.scala 283:24:@53666.4]
  assign _GEN_4 = _T_102 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53667.4]
  assign _T_106 = $signed(io_in_5) - $signed(-6'sh1); // @[Modules.scala 282:31:@53673.4]
  assign _T_107 = _T_106[5:0]; // @[Modules.scala 282:31:@53674.4]
  assign buffer_5 = $signed(_T_107); // @[Modules.scala 282:31:@53675.4]
  assign _T_110 = $signed(buffer_5) >= $signed(6'sh0); // @[Modules.scala 283:24:@53677.4]
  assign _GEN_5 = _T_110 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53678.4]
  assign _T_114 = $signed(io_in_6) - $signed(6'sh0); // @[Modules.scala 282:31:@53684.4]
  assign _T_115 = _T_114[5:0]; // @[Modules.scala 282:31:@53685.4]
  assign buffer_6 = $signed(_T_115); // @[Modules.scala 282:31:@53686.4]
  assign _T_118 = $signed(buffer_6) >= $signed(6'sh0); // @[Modules.scala 283:24:@53688.4]
  assign _GEN_6 = _T_118 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53689.4]
  assign _T_122 = $signed(io_in_7) - $signed(6'sh0); // @[Modules.scala 282:31:@53695.4]
  assign _T_123 = _T_122[5:0]; // @[Modules.scala 282:31:@53696.4]
  assign buffer_7 = $signed(_T_123); // @[Modules.scala 282:31:@53697.4]
  assign _T_126 = $signed(buffer_7) >= $signed(6'sh0); // @[Modules.scala 283:24:@53699.4]
  assign _GEN_7 = _T_126 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53700.4]
  assign _T_130 = $signed(io_in_8) - $signed(6'sh0); // @[Modules.scala 282:31:@53706.4]
  assign _T_131 = _T_130[5:0]; // @[Modules.scala 282:31:@53707.4]
  assign buffer_8 = $signed(_T_131); // @[Modules.scala 282:31:@53708.4]
  assign _T_134 = $signed(buffer_8) >= $signed(6'sh0); // @[Modules.scala 283:24:@53710.4]
  assign _GEN_8 = _T_134 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53711.4]
  assign _T_138 = $signed(io_in_9) - $signed(6'sh0); // @[Modules.scala 282:31:@53717.4]
  assign _T_139 = _T_138[5:0]; // @[Modules.scala 282:31:@53718.4]
  assign buffer_9 = $signed(_T_139); // @[Modules.scala 282:31:@53719.4]
  assign _T_142 = $signed(buffer_9) >= $signed(6'sh0); // @[Modules.scala 283:24:@53721.4]
  assign _GEN_9 = _T_142 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53722.4]
  assign _T_146 = $signed(io_in_10) - $signed(6'sh1); // @[Modules.scala 282:31:@53728.4]
  assign _T_147 = _T_146[5:0]; // @[Modules.scala 282:31:@53729.4]
  assign buffer_10 = $signed(_T_147); // @[Modules.scala 282:31:@53730.4]
  assign _T_150 = $signed(buffer_10) >= $signed(6'sh0); // @[Modules.scala 283:24:@53732.4]
  assign _GEN_10 = _T_150 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53733.4]
  assign _T_154 = $signed(io_in_11) - $signed(-6'sh4); // @[Modules.scala 282:31:@53739.4]
  assign _T_155 = _T_154[5:0]; // @[Modules.scala 282:31:@53740.4]
  assign buffer_11 = $signed(_T_155); // @[Modules.scala 282:31:@53741.4]
  assign _T_158 = $signed(buffer_11) >= $signed(6'sh0); // @[Modules.scala 283:24:@53743.4]
  assign _GEN_11 = _T_158 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53744.4]
  assign _T_162 = $signed(io_in_12) - $signed(6'sh0); // @[Modules.scala 282:31:@53750.4]
  assign _T_163 = _T_162[5:0]; // @[Modules.scala 282:31:@53751.4]
  assign buffer_12 = $signed(_T_163); // @[Modules.scala 282:31:@53752.4]
  assign _T_166 = $signed(buffer_12) >= $signed(6'sh0); // @[Modules.scala 283:24:@53754.4]
  assign _GEN_12 = _T_166 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53755.4]
  assign _T_170 = $signed(io_in_13) - $signed(-6'sh1); // @[Modules.scala 282:31:@53761.4]
  assign _T_171 = _T_170[5:0]; // @[Modules.scala 282:31:@53762.4]
  assign buffer_13 = $signed(_T_171); // @[Modules.scala 282:31:@53763.4]
  assign _T_174 = $signed(buffer_13) >= $signed(6'sh0); // @[Modules.scala 283:24:@53765.4]
  assign _GEN_13 = _T_174 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53766.4]
  assign _T_178 = $signed(io_in_14) - $signed(-6'sh1); // @[Modules.scala 282:31:@53772.4]
  assign _T_179 = _T_178[5:0]; // @[Modules.scala 282:31:@53773.4]
  assign buffer_14 = $signed(_T_179); // @[Modules.scala 282:31:@53774.4]
  assign _T_182 = $signed(buffer_14) >= $signed(6'sh0); // @[Modules.scala 283:24:@53776.4]
  assign _GEN_14 = _T_182 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53777.4]
  assign _T_186 = $signed(io_in_15) - $signed(6'sh1); // @[Modules.scala 282:31:@53783.4]
  assign _T_187 = _T_186[5:0]; // @[Modules.scala 282:31:@53784.4]
  assign buffer_15 = $signed(_T_187); // @[Modules.scala 282:31:@53785.4]
  assign _T_190 = $signed(buffer_15) >= $signed(6'sh0); // @[Modules.scala 283:24:@53787.4]
  assign _GEN_15 = _T_190 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 283:32:@53788.4]
  assign io_out_0 = {{4{_GEN_0[1]}},_GEN_0};
  assign io_out_1 = {{4{_GEN_1[1]}},_GEN_1};
  assign io_out_2 = {{4{_GEN_2[1]}},_GEN_2};
  assign io_out_3 = {{4{_GEN_3[1]}},_GEN_3};
  assign io_out_4 = {{4{_GEN_4[1]}},_GEN_4};
  assign io_out_5 = {{4{_GEN_5[1]}},_GEN_5};
  assign io_out_6 = {{4{_GEN_6[1]}},_GEN_6};
  assign io_out_7 = {{4{_GEN_7[1]}},_GEN_7};
  assign io_out_8 = {{4{_GEN_8[1]}},_GEN_8};
  assign io_out_9 = {{4{_GEN_9[1]}},_GEN_9};
  assign io_out_10 = {{4{_GEN_10[1]}},_GEN_10};
  assign io_out_11 = {{4{_GEN_11[1]}},_GEN_11};
  assign io_out_12 = {{4{_GEN_12[1]}},_GEN_12};
  assign io_out_13 = {{4{_GEN_13[1]}},_GEN_13};
  assign io_out_14 = {{4{_GEN_14[1]}},_GEN_14};
  assign io_out_15 = {{4{_GEN_15[1]}},_GEN_15};
endmodule
module Linear_p_2( // @[:@53795.2]
  input  [1:0] io_in_0, // @[:@53798.4]
  input  [1:0] io_in_1, // @[:@53798.4]
  input  [1:0] io_in_2, // @[:@53798.4]
  input  [1:0] io_in_3, // @[:@53798.4]
  input  [1:0] io_in_4, // @[:@53798.4]
  input  [1:0] io_in_5, // @[:@53798.4]
  input  [1:0] io_in_6, // @[:@53798.4]
  input  [1:0] io_in_7, // @[:@53798.4]
  input  [1:0] io_in_8, // @[:@53798.4]
  input  [1:0] io_in_9, // @[:@53798.4]
  input  [1:0] io_in_10, // @[:@53798.4]
  input  [1:0] io_in_11, // @[:@53798.4]
  input  [1:0] io_in_12, // @[:@53798.4]
  input  [1:0] io_in_13, // @[:@53798.4]
  input  [1:0] io_in_14, // @[:@53798.4]
  input  [1:0] io_in_15, // @[:@53798.4]
  output [5:0] io_out_0, // @[:@53798.4]
  output [5:0] io_out_1, // @[:@53798.4]
  output [5:0] io_out_2, // @[:@53798.4]
  output [5:0] io_out_3, // @[:@53798.4]
  output [5:0] io_out_4, // @[:@53798.4]
  output [5:0] io_out_5, // @[:@53798.4]
  output [5:0] io_out_6, // @[:@53798.4]
  output [5:0] io_out_7, // @[:@53798.4]
  output [5:0] io_out_8, // @[:@53798.4]
  output [5:0] io_out_9 // @[:@53798.4]
);
  wire [2:0] _T_793; // @[Modules.scala 143:74:@53801.4]
  wire [2:0] _T_795; // @[Modules.scala 144:80:@53802.4]
  wire [3:0] _T_796; // @[Modules.scala 143:103:@53803.4]
  wire [2:0] _T_797; // @[Modules.scala 143:103:@53804.4]
  wire [2:0] _T_798; // @[Modules.scala 143:103:@53805.4]
  wire [2:0] _T_800; // @[Modules.scala 143:74:@53807.4]
  wire [2:0] _T_802; // @[Modules.scala 144:80:@53808.4]
  wire [3:0] _T_803; // @[Modules.scala 143:103:@53809.4]
  wire [2:0] _T_804; // @[Modules.scala 143:103:@53810.4]
  wire [2:0] _T_805; // @[Modules.scala 143:103:@53811.4]
  wire [2:0] _T_807; // @[Modules.scala 143:74:@53813.4]
  wire [2:0] _T_809; // @[Modules.scala 144:80:@53814.4]
  wire [3:0] _T_810; // @[Modules.scala 143:103:@53815.4]
  wire [2:0] _T_811; // @[Modules.scala 143:103:@53816.4]
  wire [2:0] _T_812; // @[Modules.scala 143:103:@53817.4]
  wire [2:0] _T_814; // @[Modules.scala 143:74:@53819.4]
  wire [3:0] _T_816; // @[Modules.scala 144:80:@53820.4]
  wire [3:0] _GEN_0; // @[Modules.scala 143:103:@53821.4]
  wire [4:0] _T_817; // @[Modules.scala 143:103:@53821.4]
  wire [3:0] _T_818; // @[Modules.scala 143:103:@53822.4]
  wire [3:0] _T_819; // @[Modules.scala 143:103:@53823.4]
  wire [3:0] _T_821; // @[Modules.scala 143:74:@53825.4]
  wire [2:0] _T_823; // @[Modules.scala 144:80:@53826.4]
  wire [3:0] _GEN_1; // @[Modules.scala 143:103:@53827.4]
  wire [4:0] _T_824; // @[Modules.scala 143:103:@53827.4]
  wire [3:0] _T_825; // @[Modules.scala 143:103:@53828.4]
  wire [3:0] _T_826; // @[Modules.scala 143:103:@53829.4]
  wire [3:0] _T_828; // @[Modules.scala 143:74:@53831.4]
  wire [3:0] _T_830; // @[Modules.scala 144:80:@53832.4]
  wire [4:0] _T_831; // @[Modules.scala 143:103:@53833.4]
  wire [3:0] _T_832; // @[Modules.scala 143:103:@53834.4]
  wire [3:0] _T_833; // @[Modules.scala 143:103:@53835.4]
  wire [3:0] _T_835; // @[Modules.scala 143:74:@53837.4]
  wire [3:0] _T_837; // @[Modules.scala 144:80:@53838.4]
  wire [4:0] _T_838; // @[Modules.scala 143:103:@53839.4]
  wire [3:0] _T_839; // @[Modules.scala 143:103:@53840.4]
  wire [3:0] _T_840; // @[Modules.scala 143:103:@53841.4]
  wire [5:0] buffer_0_0; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_0_1; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_841; // @[Modules.scala 166:64:@53843.4]
  wire [5:0] _T_842; // @[Modules.scala 166:64:@53844.4]
  wire [5:0] buffer_0_7; // @[Modules.scala 166:64:@53845.4]
  wire [5:0] buffer_0_2; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_0_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_844; // @[Modules.scala 166:64:@53847.4]
  wire [5:0] _T_845; // @[Modules.scala 166:64:@53848.4]
  wire [5:0] buffer_0_8; // @[Modules.scala 166:64:@53849.4]
  wire [5:0] buffer_0_4; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_0_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_847; // @[Modules.scala 166:64:@53851.4]
  wire [5:0] _T_848; // @[Modules.scala 166:64:@53852.4]
  wire [5:0] buffer_0_9; // @[Modules.scala 166:64:@53853.4]
  wire [6:0] _T_850; // @[Modules.scala 166:64:@53855.4]
  wire [5:0] _T_851; // @[Modules.scala 166:64:@53856.4]
  wire [5:0] buffer_0_10; // @[Modules.scala 166:64:@53857.4]
  wire [5:0] buffer_0_6; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_853; // @[Modules.scala 172:66:@53859.4]
  wire [5:0] _T_854; // @[Modules.scala 172:66:@53860.4]
  wire [5:0] buffer_0_11; // @[Modules.scala 172:66:@53861.4]
  wire [6:0] _T_856; // @[Modules.scala 160:64:@53863.4]
  wire [5:0] _T_857; // @[Modules.scala 160:64:@53864.4]
  wire [5:0] buffer_0_12; // @[Modules.scala 160:64:@53865.4]
  wire [3:0] _T_860; // @[Modules.scala 143:74:@53870.4]
  wire [2:0] _T_862; // @[Modules.scala 144:80:@53871.4]
  wire [3:0] _GEN_2; // @[Modules.scala 143:103:@53872.4]
  wire [4:0] _T_863; // @[Modules.scala 143:103:@53872.4]
  wire [3:0] _T_864; // @[Modules.scala 143:103:@53873.4]
  wire [3:0] _T_865; // @[Modules.scala 143:103:@53874.4]
  wire [3:0] _T_867; // @[Modules.scala 143:74:@53876.4]
  wire [3:0] _T_869; // @[Modules.scala 144:80:@53877.4]
  wire [4:0] _T_870; // @[Modules.scala 143:103:@53878.4]
  wire [3:0] _T_871; // @[Modules.scala 143:103:@53879.4]
  wire [3:0] _T_872; // @[Modules.scala 143:103:@53880.4]
  wire [3:0] _T_877; // @[Modules.scala 143:103:@53884.4]
  wire [2:0] _T_878; // @[Modules.scala 143:103:@53885.4]
  wire [2:0] _T_879; // @[Modules.scala 143:103:@53886.4]
  wire [3:0] _T_883; // @[Modules.scala 144:80:@53889.4]
  wire [3:0] _GEN_3; // @[Modules.scala 143:103:@53890.4]
  wire [4:0] _T_884; // @[Modules.scala 143:103:@53890.4]
  wire [3:0] _T_885; // @[Modules.scala 143:103:@53891.4]
  wire [3:0] _T_886; // @[Modules.scala 143:103:@53892.4]
  wire [2:0] _T_888; // @[Modules.scala 143:74:@53894.4]
  wire [2:0] _T_890; // @[Modules.scala 144:80:@53895.4]
  wire [3:0] _T_891; // @[Modules.scala 143:103:@53896.4]
  wire [2:0] _T_892; // @[Modules.scala 143:103:@53897.4]
  wire [2:0] _T_893; // @[Modules.scala 143:103:@53898.4]
  wire [3:0] _T_895; // @[Modules.scala 143:74:@53900.4]
  wire [2:0] _T_897; // @[Modules.scala 144:80:@53901.4]
  wire [3:0] _GEN_4; // @[Modules.scala 143:103:@53902.4]
  wire [4:0] _T_898; // @[Modules.scala 143:103:@53902.4]
  wire [3:0] _T_899; // @[Modules.scala 143:103:@53903.4]
  wire [3:0] _T_900; // @[Modules.scala 143:103:@53904.4]
  wire [2:0] _T_902; // @[Modules.scala 143:74:@53906.4]
  wire [2:0] _T_904; // @[Modules.scala 144:80:@53907.4]
  wire [3:0] _T_905; // @[Modules.scala 143:103:@53908.4]
  wire [2:0] _T_906; // @[Modules.scala 143:103:@53909.4]
  wire [2:0] _T_907; // @[Modules.scala 143:103:@53910.4]
  wire [5:0] buffer_1_0; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_1_1; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_908; // @[Modules.scala 166:64:@53912.4]
  wire [5:0] _T_909; // @[Modules.scala 166:64:@53913.4]
  wire [5:0] buffer_1_7; // @[Modules.scala 166:64:@53914.4]
  wire [5:0] buffer_1_2; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_1_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_911; // @[Modules.scala 166:64:@53916.4]
  wire [5:0] _T_912; // @[Modules.scala 166:64:@53917.4]
  wire [5:0] buffer_1_8; // @[Modules.scala 166:64:@53918.4]
  wire [5:0] buffer_1_4; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_1_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_914; // @[Modules.scala 166:64:@53920.4]
  wire [5:0] _T_915; // @[Modules.scala 166:64:@53921.4]
  wire [5:0] buffer_1_9; // @[Modules.scala 166:64:@53922.4]
  wire [6:0] _T_917; // @[Modules.scala 166:64:@53924.4]
  wire [5:0] _T_918; // @[Modules.scala 166:64:@53925.4]
  wire [5:0] buffer_1_10; // @[Modules.scala 166:64:@53926.4]
  wire [5:0] buffer_1_6; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_920; // @[Modules.scala 172:66:@53928.4]
  wire [5:0] _T_921; // @[Modules.scala 172:66:@53929.4]
  wire [5:0] buffer_1_11; // @[Modules.scala 172:66:@53930.4]
  wire [6:0] _T_923; // @[Modules.scala 160:64:@53932.4]
  wire [5:0] _T_924; // @[Modules.scala 160:64:@53933.4]
  wire [5:0] buffer_1_12; // @[Modules.scala 160:64:@53934.4]
  wire [3:0] _T_927; // @[Modules.scala 143:74:@53939.4]
  wire [4:0] _T_930; // @[Modules.scala 143:103:@53941.4]
  wire [3:0] _T_931; // @[Modules.scala 143:103:@53942.4]
  wire [3:0] _T_932; // @[Modules.scala 143:103:@53943.4]
  wire [2:0] _T_934; // @[Modules.scala 143:74:@53945.4]
  wire [3:0] _T_936; // @[Modules.scala 144:80:@53946.4]
  wire [3:0] _GEN_5; // @[Modules.scala 143:103:@53947.4]
  wire [4:0] _T_937; // @[Modules.scala 143:103:@53947.4]
  wire [3:0] _T_938; // @[Modules.scala 143:103:@53948.4]
  wire [3:0] _T_939; // @[Modules.scala 143:103:@53949.4]
  wire [3:0] _T_941; // @[Modules.scala 143:74:@53951.4]
  wire [4:0] _T_944; // @[Modules.scala 143:103:@53953.4]
  wire [3:0] _T_945; // @[Modules.scala 143:103:@53954.4]
  wire [3:0] _T_946; // @[Modules.scala 143:103:@53955.4]
  wire [4:0] _T_951; // @[Modules.scala 143:103:@53959.4]
  wire [3:0] _T_952; // @[Modules.scala 143:103:@53960.4]
  wire [3:0] _T_953; // @[Modules.scala 143:103:@53961.4]
  wire [3:0] _T_958; // @[Modules.scala 143:103:@53965.4]
  wire [2:0] _T_959; // @[Modules.scala 143:103:@53966.4]
  wire [2:0] _T_960; // @[Modules.scala 143:103:@53967.4]
  wire [3:0] _GEN_7; // @[Modules.scala 143:103:@53971.4]
  wire [4:0] _T_965; // @[Modules.scala 143:103:@53971.4]
  wire [3:0] _T_966; // @[Modules.scala 143:103:@53972.4]
  wire [3:0] _T_967; // @[Modules.scala 143:103:@53973.4]
  wire [3:0] _GEN_8; // @[Modules.scala 143:103:@53977.4]
  wire [4:0] _T_972; // @[Modules.scala 143:103:@53977.4]
  wire [3:0] _T_973; // @[Modules.scala 143:103:@53978.4]
  wire [3:0] _T_974; // @[Modules.scala 143:103:@53979.4]
  wire [5:0] buffer_2_0; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_2_1; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_975; // @[Modules.scala 166:64:@53981.4]
  wire [5:0] _T_976; // @[Modules.scala 166:64:@53982.4]
  wire [5:0] buffer_2_7; // @[Modules.scala 166:64:@53983.4]
  wire [5:0] buffer_2_2; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_2_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_978; // @[Modules.scala 166:64:@53985.4]
  wire [5:0] _T_979; // @[Modules.scala 166:64:@53986.4]
  wire [5:0] buffer_2_8; // @[Modules.scala 166:64:@53987.4]
  wire [5:0] buffer_2_4; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_2_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_981; // @[Modules.scala 166:64:@53989.4]
  wire [5:0] _T_982; // @[Modules.scala 166:64:@53990.4]
  wire [5:0] buffer_2_9; // @[Modules.scala 166:64:@53991.4]
  wire [6:0] _T_984; // @[Modules.scala 166:64:@53993.4]
  wire [5:0] _T_985; // @[Modules.scala 166:64:@53994.4]
  wire [5:0] buffer_2_10; // @[Modules.scala 166:64:@53995.4]
  wire [5:0] buffer_2_6; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_987; // @[Modules.scala 172:66:@53997.4]
  wire [5:0] _T_988; // @[Modules.scala 172:66:@53998.4]
  wire [5:0] buffer_2_11; // @[Modules.scala 172:66:@53999.4]
  wire [6:0] _T_990; // @[Modules.scala 160:64:@54001.4]
  wire [5:0] _T_991; // @[Modules.scala 160:64:@54002.4]
  wire [5:0] buffer_2_12; // @[Modules.scala 160:64:@54003.4]
  wire [3:0] _T_997; // @[Modules.scala 150:103:@54010.4]
  wire [2:0] _T_998; // @[Modules.scala 150:103:@54011.4]
  wire [2:0] _T_999; // @[Modules.scala 150:103:@54012.4]
  wire [3:0] _GEN_9; // @[Modules.scala 150:103:@54016.4]
  wire [4:0] _T_1004; // @[Modules.scala 150:103:@54016.4]
  wire [3:0] _T_1005; // @[Modules.scala 150:103:@54017.4]
  wire [3:0] _T_1006; // @[Modules.scala 150:103:@54018.4]
  wire [3:0] _T_1008; // @[Modules.scala 150:74:@54020.4]
  wire [4:0] _T_1011; // @[Modules.scala 150:103:@54022.4]
  wire [3:0] _T_1012; // @[Modules.scala 150:103:@54023.4]
  wire [3:0] _T_1013; // @[Modules.scala 150:103:@54024.4]
  wire [3:0] _T_1017; // @[Modules.scala 151:80:@54027.4]
  wire [3:0] _GEN_10; // @[Modules.scala 150:103:@54028.4]
  wire [4:0] _T_1018; // @[Modules.scala 150:103:@54028.4]
  wire [3:0] _T_1019; // @[Modules.scala 150:103:@54029.4]
  wire [3:0] _T_1020; // @[Modules.scala 150:103:@54030.4]
  wire [4:0] _T_1032; // @[Modules.scala 150:103:@54040.4]
  wire [3:0] _T_1033; // @[Modules.scala 150:103:@54041.4]
  wire [3:0] _T_1034; // @[Modules.scala 150:103:@54042.4]
  wire [2:0] _T_1038; // @[Modules.scala 151:80:@54045.4]
  wire [3:0] _T_1039; // @[Modules.scala 150:103:@54046.4]
  wire [2:0] _T_1040; // @[Modules.scala 150:103:@54047.4]
  wire [2:0] _T_1041; // @[Modules.scala 150:103:@54048.4]
  wire [5:0] buffer_3_0; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_3_1; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1044; // @[Modules.scala 160:64:@54052.4]
  wire [5:0] _T_1045; // @[Modules.scala 160:64:@54053.4]
  wire [5:0] buffer_3_8; // @[Modules.scala 160:64:@54054.4]
  wire [5:0] buffer_3_2; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_3_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1047; // @[Modules.scala 160:64:@54056.4]
  wire [5:0] _T_1048; // @[Modules.scala 160:64:@54057.4]
  wire [5:0] buffer_3_9; // @[Modules.scala 160:64:@54058.4]
  wire [5:0] buffer_3_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1050; // @[Modules.scala 160:64:@54060.4]
  wire [5:0] _T_1051; // @[Modules.scala 160:64:@54061.4]
  wire [5:0] buffer_3_10; // @[Modules.scala 160:64:@54062.4]
  wire [5:0] buffer_3_6; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_3_7; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1053; // @[Modules.scala 160:64:@54064.4]
  wire [5:0] _T_1054; // @[Modules.scala 160:64:@54065.4]
  wire [5:0] buffer_3_11; // @[Modules.scala 160:64:@54066.4]
  wire [6:0] _T_1056; // @[Modules.scala 160:64:@54068.4]
  wire [5:0] _T_1057; // @[Modules.scala 160:64:@54069.4]
  wire [5:0] buffer_3_12; // @[Modules.scala 160:64:@54070.4]
  wire [6:0] _T_1059; // @[Modules.scala 160:64:@54072.4]
  wire [5:0] _T_1060; // @[Modules.scala 160:64:@54073.4]
  wire [5:0] buffer_3_13; // @[Modules.scala 160:64:@54074.4]
  wire [6:0] _T_1062; // @[Modules.scala 160:64:@54076.4]
  wire [5:0] _T_1063; // @[Modules.scala 160:64:@54077.4]
  wire [5:0] buffer_3_14; // @[Modules.scala 160:64:@54078.4]
  wire [4:0] _T_1069; // @[Modules.scala 143:103:@54083.4]
  wire [3:0] _T_1070; // @[Modules.scala 143:103:@54084.4]
  wire [3:0] _T_1071; // @[Modules.scala 143:103:@54085.4]
  wire [3:0] _T_1076; // @[Modules.scala 143:103:@54089.4]
  wire [2:0] _T_1077; // @[Modules.scala 143:103:@54090.4]
  wire [2:0] _T_1078; // @[Modules.scala 143:103:@54091.4]
  wire [4:0] _T_1090; // @[Modules.scala 143:103:@54101.4]
  wire [3:0] _T_1091; // @[Modules.scala 143:103:@54102.4]
  wire [3:0] _T_1092; // @[Modules.scala 143:103:@54103.4]
  wire [3:0] _T_1097; // @[Modules.scala 143:103:@54107.4]
  wire [2:0] _T_1098; // @[Modules.scala 143:103:@54108.4]
  wire [2:0] _T_1099; // @[Modules.scala 143:103:@54109.4]
  wire [3:0] _GEN_13; // @[Modules.scala 143:103:@54113.4]
  wire [4:0] _T_1104; // @[Modules.scala 143:103:@54113.4]
  wire [3:0] _T_1105; // @[Modules.scala 143:103:@54114.4]
  wire [3:0] _T_1106; // @[Modules.scala 143:103:@54115.4]
  wire [4:0] _T_1111; // @[Modules.scala 143:103:@54119.4]
  wire [3:0] _T_1112; // @[Modules.scala 143:103:@54120.4]
  wire [3:0] _T_1113; // @[Modules.scala 143:103:@54121.4]
  wire [3:0] _GEN_15; // @[Modules.scala 143:103:@54125.4]
  wire [4:0] _T_1118; // @[Modules.scala 143:103:@54125.4]
  wire [3:0] _T_1119; // @[Modules.scala 143:103:@54126.4]
  wire [3:0] _T_1120; // @[Modules.scala 143:103:@54127.4]
  wire [5:0] buffer_4_0; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_4_1; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1121; // @[Modules.scala 160:64:@54129.4]
  wire [5:0] _T_1122; // @[Modules.scala 160:64:@54130.4]
  wire [5:0] buffer_4_8; // @[Modules.scala 160:64:@54131.4]
  wire [5:0] buffer_4_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1124; // @[Modules.scala 160:64:@54133.4]
  wire [5:0] _T_1125; // @[Modules.scala 160:64:@54134.4]
  wire [5:0] buffer_4_9; // @[Modules.scala 160:64:@54135.4]
  wire [5:0] buffer_4_4; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_4_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1127; // @[Modules.scala 160:64:@54137.4]
  wire [5:0] _T_1128; // @[Modules.scala 160:64:@54138.4]
  wire [5:0] buffer_4_10; // @[Modules.scala 160:64:@54139.4]
  wire [5:0] buffer_4_6; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_4_7; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1130; // @[Modules.scala 160:64:@54141.4]
  wire [5:0] _T_1131; // @[Modules.scala 160:64:@54142.4]
  wire [5:0] buffer_4_11; // @[Modules.scala 160:64:@54143.4]
  wire [6:0] _T_1133; // @[Modules.scala 160:64:@54145.4]
  wire [5:0] _T_1134; // @[Modules.scala 160:64:@54146.4]
  wire [5:0] buffer_4_12; // @[Modules.scala 160:64:@54147.4]
  wire [6:0] _T_1136; // @[Modules.scala 160:64:@54149.4]
  wire [5:0] _T_1137; // @[Modules.scala 160:64:@54150.4]
  wire [5:0] buffer_4_13; // @[Modules.scala 160:64:@54151.4]
  wire [6:0] _T_1139; // @[Modules.scala 160:64:@54153.4]
  wire [5:0] _T_1140; // @[Modules.scala 160:64:@54154.4]
  wire [5:0] buffer_4_14; // @[Modules.scala 160:64:@54155.4]
  wire [4:0] _T_1167; // @[Modules.scala 143:103:@54178.4]
  wire [3:0] _T_1168; // @[Modules.scala 143:103:@54179.4]
  wire [3:0] _T_1169; // @[Modules.scala 143:103:@54180.4]
  wire [4:0] _T_1174; // @[Modules.scala 143:103:@54184.4]
  wire [3:0] _T_1175; // @[Modules.scala 143:103:@54185.4]
  wire [3:0] _T_1176; // @[Modules.scala 143:103:@54186.4]
  wire [4:0] _T_1181; // @[Modules.scala 143:103:@54190.4]
  wire [3:0] _T_1182; // @[Modules.scala 143:103:@54191.4]
  wire [3:0] _T_1183; // @[Modules.scala 143:103:@54192.4]
  wire [6:0] _T_1191; // @[Modules.scala 166:64:@54200.4]
  wire [5:0] _T_1192; // @[Modules.scala 166:64:@54201.4]
  wire [5:0] buffer_5_7; // @[Modules.scala 166:64:@54202.4]
  wire [5:0] buffer_5_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1194; // @[Modules.scala 166:64:@54204.4]
  wire [5:0] _T_1195; // @[Modules.scala 166:64:@54205.4]
  wire [5:0] buffer_5_8; // @[Modules.scala 166:64:@54206.4]
  wire [5:0] buffer_5_4; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_5_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1197; // @[Modules.scala 166:64:@54208.4]
  wire [5:0] _T_1198; // @[Modules.scala 166:64:@54209.4]
  wire [5:0] buffer_5_9; // @[Modules.scala 166:64:@54210.4]
  wire [6:0] _T_1200; // @[Modules.scala 166:64:@54212.4]
  wire [5:0] _T_1201; // @[Modules.scala 166:64:@54213.4]
  wire [5:0] buffer_5_10; // @[Modules.scala 166:64:@54214.4]
  wire [6:0] _T_1203; // @[Modules.scala 172:66:@54216.4]
  wire [5:0] _T_1204; // @[Modules.scala 172:66:@54217.4]
  wire [5:0] buffer_5_11; // @[Modules.scala 172:66:@54218.4]
  wire [6:0] _T_1206; // @[Modules.scala 160:64:@54220.4]
  wire [5:0] _T_1207; // @[Modules.scala 160:64:@54221.4]
  wire [5:0] buffer_5_12; // @[Modules.scala 160:64:@54222.4]
  wire [4:0] _T_1220; // @[Modules.scala 143:103:@54235.4]
  wire [3:0] _T_1221; // @[Modules.scala 143:103:@54236.4]
  wire [3:0] _T_1222; // @[Modules.scala 143:103:@54237.4]
  wire [4:0] _T_1248; // @[Modules.scala 143:103:@54259.4]
  wire [3:0] _T_1249; // @[Modules.scala 143:103:@54260.4]
  wire [3:0] _T_1250; // @[Modules.scala 143:103:@54261.4]
  wire [5:0] buffer_6_1; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1251; // @[Modules.scala 160:64:@54263.4]
  wire [5:0] _T_1252; // @[Modules.scala 160:64:@54264.4]
  wire [5:0] buffer_6_6; // @[Modules.scala 160:64:@54265.4]
  wire [6:0] _T_1254; // @[Modules.scala 160:64:@54267.4]
  wire [5:0] _T_1255; // @[Modules.scala 160:64:@54268.4]
  wire [5:0] buffer_6_7; // @[Modules.scala 160:64:@54269.4]
  wire [5:0] buffer_6_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1257; // @[Modules.scala 160:64:@54271.4]
  wire [5:0] _T_1258; // @[Modules.scala 160:64:@54272.4]
  wire [5:0] buffer_6_8; // @[Modules.scala 160:64:@54273.4]
  wire [6:0] _T_1260; // @[Modules.scala 166:64:@54275.4]
  wire [5:0] _T_1261; // @[Modules.scala 166:64:@54276.4]
  wire [5:0] buffer_6_9; // @[Modules.scala 166:64:@54277.4]
  wire [6:0] _T_1263; // @[Modules.scala 172:66:@54279.4]
  wire [5:0] _T_1264; // @[Modules.scala 172:66:@54280.4]
  wire [5:0] buffer_6_10; // @[Modules.scala 172:66:@54281.4]
  wire [3:0] _T_1284; // @[Modules.scala 150:103:@54302.4]
  wire [2:0] _T_1285; // @[Modules.scala 150:103:@54303.4]
  wire [2:0] _T_1286; // @[Modules.scala 150:103:@54304.4]
  wire [3:0] _GEN_20; // @[Modules.scala 150:103:@54308.4]
  wire [4:0] _T_1291; // @[Modules.scala 150:103:@54308.4]
  wire [3:0] _T_1292; // @[Modules.scala 150:103:@54309.4]
  wire [3:0] _T_1293; // @[Modules.scala 150:103:@54310.4]
  wire [4:0] _T_1298; // @[Modules.scala 150:103:@54314.4]
  wire [3:0] _T_1299; // @[Modules.scala 150:103:@54315.4]
  wire [3:0] _T_1300; // @[Modules.scala 150:103:@54316.4]
  wire [6:0] _T_1310; // @[Modules.scala 166:64:@54326.4]
  wire [5:0] _T_1311; // @[Modules.scala 166:64:@54327.4]
  wire [5:0] buffer_7_7; // @[Modules.scala 166:64:@54328.4]
  wire [5:0] buffer_7_2; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_7_3; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1313; // @[Modules.scala 166:64:@54330.4]
  wire [5:0] _T_1314; // @[Modules.scala 166:64:@54331.4]
  wire [5:0] buffer_7_8; // @[Modules.scala 166:64:@54332.4]
  wire [5:0] buffer_7_4; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1316; // @[Modules.scala 166:64:@54334.4]
  wire [5:0] _T_1317; // @[Modules.scala 166:64:@54335.4]
  wire [5:0] buffer_7_9; // @[Modules.scala 166:64:@54336.4]
  wire [6:0] _T_1319; // @[Modules.scala 166:64:@54338.4]
  wire [5:0] _T_1320; // @[Modules.scala 166:64:@54339.4]
  wire [5:0] buffer_7_10; // @[Modules.scala 166:64:@54340.4]
  wire [5:0] buffer_7_6; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1322; // @[Modules.scala 172:66:@54342.4]
  wire [5:0] _T_1323; // @[Modules.scala 172:66:@54343.4]
  wire [5:0] buffer_7_11; // @[Modules.scala 172:66:@54344.4]
  wire [6:0] _T_1325; // @[Modules.scala 160:64:@54346.4]
  wire [5:0] _T_1326; // @[Modules.scala 160:64:@54347.4]
  wire [5:0] buffer_7_12; // @[Modules.scala 160:64:@54348.4]
  wire [3:0] _GEN_22; // @[Modules.scala 143:103:@54355.4]
  wire [4:0] _T_1332; // @[Modules.scala 143:103:@54355.4]
  wire [3:0] _T_1333; // @[Modules.scala 143:103:@54356.4]
  wire [3:0] _T_1334; // @[Modules.scala 143:103:@54357.4]
  wire [3:0] _GEN_23; // @[Modules.scala 143:103:@54367.4]
  wire [4:0] _T_1346; // @[Modules.scala 143:103:@54367.4]
  wire [3:0] _T_1347; // @[Modules.scala 143:103:@54368.4]
  wire [3:0] _T_1348; // @[Modules.scala 143:103:@54369.4]
  wire [3:0] _T_1360; // @[Modules.scala 143:103:@54379.4]
  wire [2:0] _T_1361; // @[Modules.scala 143:103:@54380.4]
  wire [2:0] _T_1362; // @[Modules.scala 143:103:@54381.4]
  wire [3:0] _T_1367; // @[Modules.scala 143:103:@54385.4]
  wire [2:0] _T_1368; // @[Modules.scala 143:103:@54386.4]
  wire [2:0] _T_1369; // @[Modules.scala 143:103:@54387.4]
  wire [5:0] buffer_8_0; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1370; // @[Modules.scala 160:64:@54389.4]
  wire [5:0] _T_1371; // @[Modules.scala 160:64:@54390.4]
  wire [5:0] buffer_8_6; // @[Modules.scala 160:64:@54391.4]
  wire [5:0] buffer_8_2; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1373; // @[Modules.scala 160:64:@54393.4]
  wire [5:0] _T_1374; // @[Modules.scala 160:64:@54394.4]
  wire [5:0] buffer_8_7; // @[Modules.scala 160:64:@54395.4]
  wire [5:0] buffer_8_4; // @[Modules.scala 112:22:@53800.4]
  wire [5:0] buffer_8_5; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1376; // @[Modules.scala 160:64:@54397.4]
  wire [5:0] _T_1377; // @[Modules.scala 160:64:@54398.4]
  wire [5:0] buffer_8_8; // @[Modules.scala 160:64:@54399.4]
  wire [6:0] _T_1379; // @[Modules.scala 166:64:@54401.4]
  wire [5:0] _T_1380; // @[Modules.scala 166:64:@54402.4]
  wire [5:0] buffer_8_9; // @[Modules.scala 166:64:@54403.4]
  wire [6:0] _T_1382; // @[Modules.scala 172:66:@54405.4]
  wire [5:0] _T_1383; // @[Modules.scala 172:66:@54406.4]
  wire [5:0] buffer_8_10; // @[Modules.scala 172:66:@54407.4]
  wire [4:0] _T_1431; // @[Modules.scala 150:103:@54452.4]
  wire [3:0] _T_1432; // @[Modules.scala 150:103:@54453.4]
  wire [3:0] _T_1433; // @[Modules.scala 150:103:@54454.4]
  wire [6:0] _T_1439; // @[Modules.scala 160:64:@54462.4]
  wire [5:0] _T_1440; // @[Modules.scala 160:64:@54463.4]
  wire [5:0] buffer_9_9; // @[Modules.scala 160:64:@54464.4]
  wire [6:0] _T_1442; // @[Modules.scala 160:64:@54466.4]
  wire [5:0] _T_1443; // @[Modules.scala 160:64:@54467.4]
  wire [5:0] buffer_9_10; // @[Modules.scala 160:64:@54468.4]
  wire [5:0] buffer_9_6; // @[Modules.scala 112:22:@53800.4]
  wire [6:0] _T_1445; // @[Modules.scala 160:64:@54470.4]
  wire [5:0] _T_1446; // @[Modules.scala 160:64:@54471.4]
  wire [5:0] buffer_9_11; // @[Modules.scala 160:64:@54472.4]
  wire [6:0] _T_1448; // @[Modules.scala 160:64:@54474.4]
  wire [5:0] _T_1449; // @[Modules.scala 160:64:@54475.4]
  wire [5:0] buffer_9_12; // @[Modules.scala 160:64:@54476.4]
  wire [6:0] _T_1451; // @[Modules.scala 160:64:@54478.4]
  wire [5:0] _T_1452; // @[Modules.scala 160:64:@54479.4]
  wire [5:0] buffer_9_13; // @[Modules.scala 160:64:@54480.4]
  wire [6:0] _T_1454; // @[Modules.scala 160:64:@54482.4]
  wire [5:0] _T_1455; // @[Modules.scala 160:64:@54483.4]
  wire [5:0] buffer_9_14; // @[Modules.scala 160:64:@54484.4]
  assign _T_793 = $signed(-2'sh1) * $signed(io_in_0); // @[Modules.scala 143:74:@53801.4]
  assign _T_795 = $signed(-2'sh1) * $signed(io_in_2); // @[Modules.scala 144:80:@53802.4]
  assign _T_796 = $signed(_T_793) + $signed(_T_795); // @[Modules.scala 143:103:@53803.4]
  assign _T_797 = _T_796[2:0]; // @[Modules.scala 143:103:@53804.4]
  assign _T_798 = $signed(_T_797); // @[Modules.scala 143:103:@53805.4]
  assign _T_800 = $signed(-2'sh1) * $signed(io_in_3); // @[Modules.scala 143:74:@53807.4]
  assign _T_802 = $signed(-2'sh1) * $signed(io_in_5); // @[Modules.scala 144:80:@53808.4]
  assign _T_803 = $signed(_T_800) + $signed(_T_802); // @[Modules.scala 143:103:@53809.4]
  assign _T_804 = _T_803[2:0]; // @[Modules.scala 143:103:@53810.4]
  assign _T_805 = $signed(_T_804); // @[Modules.scala 143:103:@53811.4]
  assign _T_807 = $signed(-2'sh1) * $signed(io_in_6); // @[Modules.scala 143:74:@53813.4]
  assign _T_809 = $signed(-2'sh1) * $signed(io_in_7); // @[Modules.scala 144:80:@53814.4]
  assign _T_810 = $signed(_T_807) + $signed(_T_809); // @[Modules.scala 143:103:@53815.4]
  assign _T_811 = _T_810[2:0]; // @[Modules.scala 143:103:@53816.4]
  assign _T_812 = $signed(_T_811); // @[Modules.scala 143:103:@53817.4]
  assign _T_814 = $signed(-2'sh1) * $signed(io_in_8); // @[Modules.scala 143:74:@53819.4]
  assign _T_816 = $signed(2'sh1) * $signed(io_in_9); // @[Modules.scala 144:80:@53820.4]
  assign _GEN_0 = {{1{_T_814[2]}},_T_814}; // @[Modules.scala 143:103:@53821.4]
  assign _T_817 = $signed(_GEN_0) + $signed(_T_816); // @[Modules.scala 143:103:@53821.4]
  assign _T_818 = _T_817[3:0]; // @[Modules.scala 143:103:@53822.4]
  assign _T_819 = $signed(_T_818); // @[Modules.scala 143:103:@53823.4]
  assign _T_821 = $signed(2'sh1) * $signed(io_in_10); // @[Modules.scala 143:74:@53825.4]
  assign _T_823 = $signed(-2'sh1) * $signed(io_in_11); // @[Modules.scala 144:80:@53826.4]
  assign _GEN_1 = {{1{_T_823[2]}},_T_823}; // @[Modules.scala 143:103:@53827.4]
  assign _T_824 = $signed(_T_821) + $signed(_GEN_1); // @[Modules.scala 143:103:@53827.4]
  assign _T_825 = _T_824[3:0]; // @[Modules.scala 143:103:@53828.4]
  assign _T_826 = $signed(_T_825); // @[Modules.scala 143:103:@53829.4]
  assign _T_828 = $signed(2'sh1) * $signed(io_in_12); // @[Modules.scala 143:74:@53831.4]
  assign _T_830 = $signed(2'sh1) * $signed(io_in_13); // @[Modules.scala 144:80:@53832.4]
  assign _T_831 = $signed(_T_828) + $signed(_T_830); // @[Modules.scala 143:103:@53833.4]
  assign _T_832 = _T_831[3:0]; // @[Modules.scala 143:103:@53834.4]
  assign _T_833 = $signed(_T_832); // @[Modules.scala 143:103:@53835.4]
  assign _T_835 = $signed(2'sh1) * $signed(io_in_14); // @[Modules.scala 143:74:@53837.4]
  assign _T_837 = $signed(2'sh1) * $signed(io_in_15); // @[Modules.scala 144:80:@53838.4]
  assign _T_838 = $signed(_T_835) + $signed(_T_837); // @[Modules.scala 143:103:@53839.4]
  assign _T_839 = _T_838[3:0]; // @[Modules.scala 143:103:@53840.4]
  assign _T_840 = $signed(_T_839); // @[Modules.scala 143:103:@53841.4]
  assign buffer_0_0 = {{3{_T_798[2]}},_T_798}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_0_1 = {{3{_T_805[2]}},_T_805}; // @[Modules.scala 112:22:@53800.4]
  assign _T_841 = $signed(buffer_0_0) + $signed(buffer_0_1); // @[Modules.scala 166:64:@53843.4]
  assign _T_842 = _T_841[5:0]; // @[Modules.scala 166:64:@53844.4]
  assign buffer_0_7 = $signed(_T_842); // @[Modules.scala 166:64:@53845.4]
  assign buffer_0_2 = {{3{_T_812[2]}},_T_812}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_0_3 = {{2{_T_819[3]}},_T_819}; // @[Modules.scala 112:22:@53800.4]
  assign _T_844 = $signed(buffer_0_2) + $signed(buffer_0_3); // @[Modules.scala 166:64:@53847.4]
  assign _T_845 = _T_844[5:0]; // @[Modules.scala 166:64:@53848.4]
  assign buffer_0_8 = $signed(_T_845); // @[Modules.scala 166:64:@53849.4]
  assign buffer_0_4 = {{2{_T_826[3]}},_T_826}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_0_5 = {{2{_T_833[3]}},_T_833}; // @[Modules.scala 112:22:@53800.4]
  assign _T_847 = $signed(buffer_0_4) + $signed(buffer_0_5); // @[Modules.scala 166:64:@53851.4]
  assign _T_848 = _T_847[5:0]; // @[Modules.scala 166:64:@53852.4]
  assign buffer_0_9 = $signed(_T_848); // @[Modules.scala 166:64:@53853.4]
  assign _T_850 = $signed(buffer_0_7) + $signed(buffer_0_8); // @[Modules.scala 166:64:@53855.4]
  assign _T_851 = _T_850[5:0]; // @[Modules.scala 166:64:@53856.4]
  assign buffer_0_10 = $signed(_T_851); // @[Modules.scala 166:64:@53857.4]
  assign buffer_0_6 = {{2{_T_840[3]}},_T_840}; // @[Modules.scala 112:22:@53800.4]
  assign _T_853 = $signed(buffer_0_9) + $signed(buffer_0_6); // @[Modules.scala 172:66:@53859.4]
  assign _T_854 = _T_853[5:0]; // @[Modules.scala 172:66:@53860.4]
  assign buffer_0_11 = $signed(_T_854); // @[Modules.scala 172:66:@53861.4]
  assign _T_856 = $signed(buffer_0_10) + $signed(buffer_0_11); // @[Modules.scala 160:64:@53863.4]
  assign _T_857 = _T_856[5:0]; // @[Modules.scala 160:64:@53864.4]
  assign buffer_0_12 = $signed(_T_857); // @[Modules.scala 160:64:@53865.4]
  assign _T_860 = $signed(2'sh1) * $signed(io_in_0); // @[Modules.scala 143:74:@53870.4]
  assign _T_862 = $signed(-2'sh1) * $signed(io_in_1); // @[Modules.scala 144:80:@53871.4]
  assign _GEN_2 = {{1{_T_862[2]}},_T_862}; // @[Modules.scala 143:103:@53872.4]
  assign _T_863 = $signed(_T_860) + $signed(_GEN_2); // @[Modules.scala 143:103:@53872.4]
  assign _T_864 = _T_863[3:0]; // @[Modules.scala 143:103:@53873.4]
  assign _T_865 = $signed(_T_864); // @[Modules.scala 143:103:@53874.4]
  assign _T_867 = $signed(2'sh1) * $signed(io_in_2); // @[Modules.scala 143:74:@53876.4]
  assign _T_869 = $signed(2'sh1) * $signed(io_in_3); // @[Modules.scala 144:80:@53877.4]
  assign _T_870 = $signed(_T_867) + $signed(_T_869); // @[Modules.scala 143:103:@53878.4]
  assign _T_871 = _T_870[3:0]; // @[Modules.scala 143:103:@53879.4]
  assign _T_872 = $signed(_T_871); // @[Modules.scala 143:103:@53880.4]
  assign _T_877 = $signed(_T_802) + $signed(_T_807); // @[Modules.scala 143:103:@53884.4]
  assign _T_878 = _T_877[2:0]; // @[Modules.scala 143:103:@53885.4]
  assign _T_879 = $signed(_T_878); // @[Modules.scala 143:103:@53886.4]
  assign _T_883 = $signed(2'sh1) * $signed(io_in_8); // @[Modules.scala 144:80:@53889.4]
  assign _GEN_3 = {{1{_T_809[2]}},_T_809}; // @[Modules.scala 143:103:@53890.4]
  assign _T_884 = $signed(_GEN_3) + $signed(_T_883); // @[Modules.scala 143:103:@53890.4]
  assign _T_885 = _T_884[3:0]; // @[Modules.scala 143:103:@53891.4]
  assign _T_886 = $signed(_T_885); // @[Modules.scala 143:103:@53892.4]
  assign _T_888 = $signed(-2'sh1) * $signed(io_in_9); // @[Modules.scala 143:74:@53894.4]
  assign _T_890 = $signed(-2'sh1) * $signed(io_in_10); // @[Modules.scala 144:80:@53895.4]
  assign _T_891 = $signed(_T_888) + $signed(_T_890); // @[Modules.scala 143:103:@53896.4]
  assign _T_892 = _T_891[2:0]; // @[Modules.scala 143:103:@53897.4]
  assign _T_893 = $signed(_T_892); // @[Modules.scala 143:103:@53898.4]
  assign _T_895 = $signed(2'sh1) * $signed(io_in_11); // @[Modules.scala 143:74:@53900.4]
  assign _T_897 = $signed(-2'sh1) * $signed(io_in_12); // @[Modules.scala 144:80:@53901.4]
  assign _GEN_4 = {{1{_T_897[2]}},_T_897}; // @[Modules.scala 143:103:@53902.4]
  assign _T_898 = $signed(_T_895) + $signed(_GEN_4); // @[Modules.scala 143:103:@53902.4]
  assign _T_899 = _T_898[3:0]; // @[Modules.scala 143:103:@53903.4]
  assign _T_900 = $signed(_T_899); // @[Modules.scala 143:103:@53904.4]
  assign _T_902 = $signed(-2'sh1) * $signed(io_in_13); // @[Modules.scala 143:74:@53906.4]
  assign _T_904 = $signed(-2'sh1) * $signed(io_in_15); // @[Modules.scala 144:80:@53907.4]
  assign _T_905 = $signed(_T_902) + $signed(_T_904); // @[Modules.scala 143:103:@53908.4]
  assign _T_906 = _T_905[2:0]; // @[Modules.scala 143:103:@53909.4]
  assign _T_907 = $signed(_T_906); // @[Modules.scala 143:103:@53910.4]
  assign buffer_1_0 = {{2{_T_865[3]}},_T_865}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_1_1 = {{2{_T_872[3]}},_T_872}; // @[Modules.scala 112:22:@53800.4]
  assign _T_908 = $signed(buffer_1_0) + $signed(buffer_1_1); // @[Modules.scala 166:64:@53912.4]
  assign _T_909 = _T_908[5:0]; // @[Modules.scala 166:64:@53913.4]
  assign buffer_1_7 = $signed(_T_909); // @[Modules.scala 166:64:@53914.4]
  assign buffer_1_2 = {{3{_T_879[2]}},_T_879}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_1_3 = {{2{_T_886[3]}},_T_886}; // @[Modules.scala 112:22:@53800.4]
  assign _T_911 = $signed(buffer_1_2) + $signed(buffer_1_3); // @[Modules.scala 166:64:@53916.4]
  assign _T_912 = _T_911[5:0]; // @[Modules.scala 166:64:@53917.4]
  assign buffer_1_8 = $signed(_T_912); // @[Modules.scala 166:64:@53918.4]
  assign buffer_1_4 = {{3{_T_893[2]}},_T_893}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_1_5 = {{2{_T_900[3]}},_T_900}; // @[Modules.scala 112:22:@53800.4]
  assign _T_914 = $signed(buffer_1_4) + $signed(buffer_1_5); // @[Modules.scala 166:64:@53920.4]
  assign _T_915 = _T_914[5:0]; // @[Modules.scala 166:64:@53921.4]
  assign buffer_1_9 = $signed(_T_915); // @[Modules.scala 166:64:@53922.4]
  assign _T_917 = $signed(buffer_1_7) + $signed(buffer_1_8); // @[Modules.scala 166:64:@53924.4]
  assign _T_918 = _T_917[5:0]; // @[Modules.scala 166:64:@53925.4]
  assign buffer_1_10 = $signed(_T_918); // @[Modules.scala 166:64:@53926.4]
  assign buffer_1_6 = {{3{_T_907[2]}},_T_907}; // @[Modules.scala 112:22:@53800.4]
  assign _T_920 = $signed(buffer_1_9) + $signed(buffer_1_6); // @[Modules.scala 172:66:@53928.4]
  assign _T_921 = _T_920[5:0]; // @[Modules.scala 172:66:@53929.4]
  assign buffer_1_11 = $signed(_T_921); // @[Modules.scala 172:66:@53930.4]
  assign _T_923 = $signed(buffer_1_10) + $signed(buffer_1_11); // @[Modules.scala 160:64:@53932.4]
  assign _T_924 = _T_923[5:0]; // @[Modules.scala 160:64:@53933.4]
  assign buffer_1_12 = $signed(_T_924); // @[Modules.scala 160:64:@53934.4]
  assign _T_927 = $signed(2'sh1) * $signed(io_in_1); // @[Modules.scala 143:74:@53939.4]
  assign _T_930 = $signed(_T_927) + $signed(_T_869); // @[Modules.scala 143:103:@53941.4]
  assign _T_931 = _T_930[3:0]; // @[Modules.scala 143:103:@53942.4]
  assign _T_932 = $signed(_T_931); // @[Modules.scala 143:103:@53943.4]
  assign _T_934 = $signed(-2'sh1) * $signed(io_in_4); // @[Modules.scala 143:74:@53945.4]
  assign _T_936 = $signed(2'sh1) * $signed(io_in_5); // @[Modules.scala 144:80:@53946.4]
  assign _GEN_5 = {{1{_T_934[2]}},_T_934}; // @[Modules.scala 143:103:@53947.4]
  assign _T_937 = $signed(_GEN_5) + $signed(_T_936); // @[Modules.scala 143:103:@53947.4]
  assign _T_938 = _T_937[3:0]; // @[Modules.scala 143:103:@53948.4]
  assign _T_939 = $signed(_T_938); // @[Modules.scala 143:103:@53949.4]
  assign _T_941 = $signed(2'sh1) * $signed(io_in_6); // @[Modules.scala 143:74:@53951.4]
  assign _T_944 = $signed(_T_941) + $signed(_GEN_3); // @[Modules.scala 143:103:@53953.4]
  assign _T_945 = _T_944[3:0]; // @[Modules.scala 143:103:@53954.4]
  assign _T_946 = $signed(_T_945); // @[Modules.scala 143:103:@53955.4]
  assign _T_951 = $signed(_T_883) + $signed(_T_816); // @[Modules.scala 143:103:@53959.4]
  assign _T_952 = _T_951[3:0]; // @[Modules.scala 143:103:@53960.4]
  assign _T_953 = $signed(_T_952); // @[Modules.scala 143:103:@53961.4]
  assign _T_958 = $signed(_T_890) + $signed(_T_823); // @[Modules.scala 143:103:@53965.4]
  assign _T_959 = _T_958[2:0]; // @[Modules.scala 143:103:@53966.4]
  assign _T_960 = $signed(_T_959); // @[Modules.scala 143:103:@53967.4]
  assign _GEN_7 = {{1{_T_902[2]}},_T_902}; // @[Modules.scala 143:103:@53971.4]
  assign _T_965 = $signed(_T_828) + $signed(_GEN_7); // @[Modules.scala 143:103:@53971.4]
  assign _T_966 = _T_965[3:0]; // @[Modules.scala 143:103:@53972.4]
  assign _T_967 = $signed(_T_966); // @[Modules.scala 143:103:@53973.4]
  assign _GEN_8 = {{1{_T_904[2]}},_T_904}; // @[Modules.scala 143:103:@53977.4]
  assign _T_972 = $signed(_T_835) + $signed(_GEN_8); // @[Modules.scala 143:103:@53977.4]
  assign _T_973 = _T_972[3:0]; // @[Modules.scala 143:103:@53978.4]
  assign _T_974 = $signed(_T_973); // @[Modules.scala 143:103:@53979.4]
  assign buffer_2_0 = {{2{_T_932[3]}},_T_932}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_2_1 = {{2{_T_939[3]}},_T_939}; // @[Modules.scala 112:22:@53800.4]
  assign _T_975 = $signed(buffer_2_0) + $signed(buffer_2_1); // @[Modules.scala 166:64:@53981.4]
  assign _T_976 = _T_975[5:0]; // @[Modules.scala 166:64:@53982.4]
  assign buffer_2_7 = $signed(_T_976); // @[Modules.scala 166:64:@53983.4]
  assign buffer_2_2 = {{2{_T_946[3]}},_T_946}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_2_3 = {{2{_T_953[3]}},_T_953}; // @[Modules.scala 112:22:@53800.4]
  assign _T_978 = $signed(buffer_2_2) + $signed(buffer_2_3); // @[Modules.scala 166:64:@53985.4]
  assign _T_979 = _T_978[5:0]; // @[Modules.scala 166:64:@53986.4]
  assign buffer_2_8 = $signed(_T_979); // @[Modules.scala 166:64:@53987.4]
  assign buffer_2_4 = {{3{_T_960[2]}},_T_960}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_2_5 = {{2{_T_967[3]}},_T_967}; // @[Modules.scala 112:22:@53800.4]
  assign _T_981 = $signed(buffer_2_4) + $signed(buffer_2_5); // @[Modules.scala 166:64:@53989.4]
  assign _T_982 = _T_981[5:0]; // @[Modules.scala 166:64:@53990.4]
  assign buffer_2_9 = $signed(_T_982); // @[Modules.scala 166:64:@53991.4]
  assign _T_984 = $signed(buffer_2_7) + $signed(buffer_2_8); // @[Modules.scala 166:64:@53993.4]
  assign _T_985 = _T_984[5:0]; // @[Modules.scala 166:64:@53994.4]
  assign buffer_2_10 = $signed(_T_985); // @[Modules.scala 166:64:@53995.4]
  assign buffer_2_6 = {{2{_T_974[3]}},_T_974}; // @[Modules.scala 112:22:@53800.4]
  assign _T_987 = $signed(buffer_2_9) + $signed(buffer_2_6); // @[Modules.scala 172:66:@53997.4]
  assign _T_988 = _T_987[5:0]; // @[Modules.scala 172:66:@53998.4]
  assign buffer_2_11 = $signed(_T_988); // @[Modules.scala 172:66:@53999.4]
  assign _T_990 = $signed(buffer_2_10) + $signed(buffer_2_11); // @[Modules.scala 160:64:@54001.4]
  assign _T_991 = _T_990[5:0]; // @[Modules.scala 160:64:@54002.4]
  assign buffer_2_12 = $signed(_T_991); // @[Modules.scala 160:64:@54003.4]
  assign _T_997 = $signed(_T_793) + $signed(_T_862); // @[Modules.scala 150:103:@54010.4]
  assign _T_998 = _T_997[2:0]; // @[Modules.scala 150:103:@54011.4]
  assign _T_999 = $signed(_T_998); // @[Modules.scala 150:103:@54012.4]
  assign _GEN_9 = {{1{_T_795[2]}},_T_795}; // @[Modules.scala 150:103:@54016.4]
  assign _T_1004 = $signed(_GEN_9) + $signed(_T_869); // @[Modules.scala 150:103:@54016.4]
  assign _T_1005 = _T_1004[3:0]; // @[Modules.scala 150:103:@54017.4]
  assign _T_1006 = $signed(_T_1005); // @[Modules.scala 150:103:@54018.4]
  assign _T_1008 = $signed(2'sh1) * $signed(io_in_4); // @[Modules.scala 150:74:@54020.4]
  assign _T_1011 = $signed(_T_1008) + $signed(_T_936); // @[Modules.scala 150:103:@54022.4]
  assign _T_1012 = _T_1011[3:0]; // @[Modules.scala 150:103:@54023.4]
  assign _T_1013 = $signed(_T_1012); // @[Modules.scala 150:103:@54024.4]
  assign _T_1017 = $signed(2'sh1) * $signed(io_in_7); // @[Modules.scala 151:80:@54027.4]
  assign _GEN_10 = {{1{_T_807[2]}},_T_807}; // @[Modules.scala 150:103:@54028.4]
  assign _T_1018 = $signed(_GEN_10) + $signed(_T_1017); // @[Modules.scala 150:103:@54028.4]
  assign _T_1019 = _T_1018[3:0]; // @[Modules.scala 150:103:@54029.4]
  assign _T_1020 = $signed(_T_1019); // @[Modules.scala 150:103:@54030.4]
  assign _T_1032 = $signed(_T_821) + $signed(_GEN_4); // @[Modules.scala 150:103:@54040.4]
  assign _T_1033 = _T_1032[3:0]; // @[Modules.scala 150:103:@54041.4]
  assign _T_1034 = $signed(_T_1033); // @[Modules.scala 150:103:@54042.4]
  assign _T_1038 = $signed(-2'sh1) * $signed(io_in_14); // @[Modules.scala 151:80:@54045.4]
  assign _T_1039 = $signed(_T_902) + $signed(_T_1038); // @[Modules.scala 150:103:@54046.4]
  assign _T_1040 = _T_1039[2:0]; // @[Modules.scala 150:103:@54047.4]
  assign _T_1041 = $signed(_T_1040); // @[Modules.scala 150:103:@54048.4]
  assign buffer_3_0 = {{3{_T_999[2]}},_T_999}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_3_1 = {{2{_T_1006[3]}},_T_1006}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1044 = $signed(buffer_3_0) + $signed(buffer_3_1); // @[Modules.scala 160:64:@54052.4]
  assign _T_1045 = _T_1044[5:0]; // @[Modules.scala 160:64:@54053.4]
  assign buffer_3_8 = $signed(_T_1045); // @[Modules.scala 160:64:@54054.4]
  assign buffer_3_2 = {{2{_T_1013[3]}},_T_1013}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_3_3 = {{2{_T_1020[3]}},_T_1020}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1047 = $signed(buffer_3_2) + $signed(buffer_3_3); // @[Modules.scala 160:64:@54056.4]
  assign _T_1048 = _T_1047[5:0]; // @[Modules.scala 160:64:@54057.4]
  assign buffer_3_9 = $signed(_T_1048); // @[Modules.scala 160:64:@54058.4]
  assign buffer_3_5 = {{2{_T_1034[3]}},_T_1034}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1050 = $signed(buffer_2_3) + $signed(buffer_3_5); // @[Modules.scala 160:64:@54060.4]
  assign _T_1051 = _T_1050[5:0]; // @[Modules.scala 160:64:@54061.4]
  assign buffer_3_10 = $signed(_T_1051); // @[Modules.scala 160:64:@54062.4]
  assign buffer_3_6 = {{3{_T_1041[2]}},_T_1041}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_3_7 = {{3{_T_904[2]}},_T_904}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1053 = $signed(buffer_3_6) + $signed(buffer_3_7); // @[Modules.scala 160:64:@54064.4]
  assign _T_1054 = _T_1053[5:0]; // @[Modules.scala 160:64:@54065.4]
  assign buffer_3_11 = $signed(_T_1054); // @[Modules.scala 160:64:@54066.4]
  assign _T_1056 = $signed(buffer_3_8) + $signed(buffer_3_9); // @[Modules.scala 160:64:@54068.4]
  assign _T_1057 = _T_1056[5:0]; // @[Modules.scala 160:64:@54069.4]
  assign buffer_3_12 = $signed(_T_1057); // @[Modules.scala 160:64:@54070.4]
  assign _T_1059 = $signed(buffer_3_10) + $signed(buffer_3_11); // @[Modules.scala 160:64:@54072.4]
  assign _T_1060 = _T_1059[5:0]; // @[Modules.scala 160:64:@54073.4]
  assign buffer_3_13 = $signed(_T_1060); // @[Modules.scala 160:64:@54074.4]
  assign _T_1062 = $signed(buffer_3_12) + $signed(buffer_3_13); // @[Modules.scala 160:64:@54076.4]
  assign _T_1063 = _T_1062[5:0]; // @[Modules.scala 160:64:@54077.4]
  assign buffer_3_14 = $signed(_T_1063); // @[Modules.scala 160:64:@54078.4]
  assign _T_1069 = $signed(_T_860) + $signed(_T_927); // @[Modules.scala 143:103:@54083.4]
  assign _T_1070 = _T_1069[3:0]; // @[Modules.scala 143:103:@54084.4]
  assign _T_1071 = $signed(_T_1070); // @[Modules.scala 143:103:@54085.4]
  assign _T_1076 = $signed(_T_795) + $signed(_T_800); // @[Modules.scala 143:103:@54089.4]
  assign _T_1077 = _T_1076[2:0]; // @[Modules.scala 143:103:@54090.4]
  assign _T_1078 = $signed(_T_1077); // @[Modules.scala 143:103:@54091.4]
  assign _T_1090 = $signed(_T_941) + $signed(_T_1017); // @[Modules.scala 143:103:@54101.4]
  assign _T_1091 = _T_1090[3:0]; // @[Modules.scala 143:103:@54102.4]
  assign _T_1092 = $signed(_T_1091); // @[Modules.scala 143:103:@54103.4]
  assign _T_1097 = $signed(_T_814) + $signed(_T_888); // @[Modules.scala 143:103:@54107.4]
  assign _T_1098 = _T_1097[2:0]; // @[Modules.scala 143:103:@54108.4]
  assign _T_1099 = $signed(_T_1098); // @[Modules.scala 143:103:@54109.4]
  assign _GEN_13 = {{1{_T_890[2]}},_T_890}; // @[Modules.scala 143:103:@54113.4]
  assign _T_1104 = $signed(_GEN_13) + $signed(_T_895); // @[Modules.scala 143:103:@54113.4]
  assign _T_1105 = _T_1104[3:0]; // @[Modules.scala 143:103:@54114.4]
  assign _T_1106 = $signed(_T_1105); // @[Modules.scala 143:103:@54115.4]
  assign _T_1111 = $signed(_GEN_4) + $signed(_T_830); // @[Modules.scala 143:103:@54119.4]
  assign _T_1112 = _T_1111[3:0]; // @[Modules.scala 143:103:@54120.4]
  assign _T_1113 = $signed(_T_1112); // @[Modules.scala 143:103:@54121.4]
  assign _GEN_15 = {{1{_T_1038[2]}},_T_1038}; // @[Modules.scala 143:103:@54125.4]
  assign _T_1118 = $signed(_GEN_15) + $signed(_T_837); // @[Modules.scala 143:103:@54125.4]
  assign _T_1119 = _T_1118[3:0]; // @[Modules.scala 143:103:@54126.4]
  assign _T_1120 = $signed(_T_1119); // @[Modules.scala 143:103:@54127.4]
  assign buffer_4_0 = {{2{_T_1071[3]}},_T_1071}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_4_1 = {{3{_T_1078[2]}},_T_1078}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1121 = $signed(buffer_4_0) + $signed(buffer_4_1); // @[Modules.scala 160:64:@54129.4]
  assign _T_1122 = _T_1121[5:0]; // @[Modules.scala 160:64:@54130.4]
  assign buffer_4_8 = $signed(_T_1122); // @[Modules.scala 160:64:@54131.4]
  assign buffer_4_3 = {{2{_T_1092[3]}},_T_1092}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1124 = $signed(buffer_2_1) + $signed(buffer_4_3); // @[Modules.scala 160:64:@54133.4]
  assign _T_1125 = _T_1124[5:0]; // @[Modules.scala 160:64:@54134.4]
  assign buffer_4_9 = $signed(_T_1125); // @[Modules.scala 160:64:@54135.4]
  assign buffer_4_4 = {{3{_T_1099[2]}},_T_1099}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_4_5 = {{2{_T_1106[3]}},_T_1106}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1127 = $signed(buffer_4_4) + $signed(buffer_4_5); // @[Modules.scala 160:64:@54137.4]
  assign _T_1128 = _T_1127[5:0]; // @[Modules.scala 160:64:@54138.4]
  assign buffer_4_10 = $signed(_T_1128); // @[Modules.scala 160:64:@54139.4]
  assign buffer_4_6 = {{2{_T_1113[3]}},_T_1113}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_4_7 = {{2{_T_1120[3]}},_T_1120}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1130 = $signed(buffer_4_6) + $signed(buffer_4_7); // @[Modules.scala 160:64:@54141.4]
  assign _T_1131 = _T_1130[5:0]; // @[Modules.scala 160:64:@54142.4]
  assign buffer_4_11 = $signed(_T_1131); // @[Modules.scala 160:64:@54143.4]
  assign _T_1133 = $signed(buffer_4_8) + $signed(buffer_4_9); // @[Modules.scala 160:64:@54145.4]
  assign _T_1134 = _T_1133[5:0]; // @[Modules.scala 160:64:@54146.4]
  assign buffer_4_12 = $signed(_T_1134); // @[Modules.scala 160:64:@54147.4]
  assign _T_1136 = $signed(buffer_4_10) + $signed(buffer_4_11); // @[Modules.scala 160:64:@54149.4]
  assign _T_1137 = _T_1136[5:0]; // @[Modules.scala 160:64:@54150.4]
  assign buffer_4_13 = $signed(_T_1137); // @[Modules.scala 160:64:@54151.4]
  assign _T_1139 = $signed(buffer_4_12) + $signed(buffer_4_13); // @[Modules.scala 160:64:@54153.4]
  assign _T_1140 = _T_1139[5:0]; // @[Modules.scala 160:64:@54154.4]
  assign buffer_4_14 = $signed(_T_1140); // @[Modules.scala 160:64:@54155.4]
  assign _T_1167 = $signed(_T_1017) + $signed(_GEN_0); // @[Modules.scala 143:103:@54178.4]
  assign _T_1168 = _T_1167[3:0]; // @[Modules.scala 143:103:@54179.4]
  assign _T_1169 = $signed(_T_1168); // @[Modules.scala 143:103:@54180.4]
  assign _T_1174 = $signed(_T_816) + $signed(_T_821); // @[Modules.scala 143:103:@54184.4]
  assign _T_1175 = _T_1174[3:0]; // @[Modules.scala 143:103:@54185.4]
  assign _T_1176 = $signed(_T_1175); // @[Modules.scala 143:103:@54186.4]
  assign _T_1181 = $signed(_T_895) + $signed(_T_830); // @[Modules.scala 143:103:@54190.4]
  assign _T_1182 = _T_1181[3:0]; // @[Modules.scala 143:103:@54191.4]
  assign _T_1183 = $signed(_T_1182); // @[Modules.scala 143:103:@54192.4]
  assign _T_1191 = $signed(buffer_3_0) + $signed(buffer_1_1); // @[Modules.scala 166:64:@54200.4]
  assign _T_1192 = _T_1191[5:0]; // @[Modules.scala 166:64:@54201.4]
  assign buffer_5_7 = $signed(_T_1192); // @[Modules.scala 166:64:@54202.4]
  assign buffer_5_3 = {{2{_T_1169[3]}},_T_1169}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1194 = $signed(buffer_1_2) + $signed(buffer_5_3); // @[Modules.scala 166:64:@54204.4]
  assign _T_1195 = _T_1194[5:0]; // @[Modules.scala 166:64:@54205.4]
  assign buffer_5_8 = $signed(_T_1195); // @[Modules.scala 166:64:@54206.4]
  assign buffer_5_4 = {{2{_T_1176[3]}},_T_1176}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_5_5 = {{2{_T_1183[3]}},_T_1183}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1197 = $signed(buffer_5_4) + $signed(buffer_5_5); // @[Modules.scala 166:64:@54208.4]
  assign _T_1198 = _T_1197[5:0]; // @[Modules.scala 166:64:@54209.4]
  assign buffer_5_9 = $signed(_T_1198); // @[Modules.scala 166:64:@54210.4]
  assign _T_1200 = $signed(buffer_5_7) + $signed(buffer_5_8); // @[Modules.scala 166:64:@54212.4]
  assign _T_1201 = _T_1200[5:0]; // @[Modules.scala 166:64:@54213.4]
  assign buffer_5_10 = $signed(_T_1201); // @[Modules.scala 166:64:@54214.4]
  assign _T_1203 = $signed(buffer_5_9) + $signed(buffer_4_7); // @[Modules.scala 172:66:@54216.4]
  assign _T_1204 = _T_1203[5:0]; // @[Modules.scala 172:66:@54217.4]
  assign buffer_5_11 = $signed(_T_1204); // @[Modules.scala 172:66:@54218.4]
  assign _T_1206 = $signed(buffer_5_10) + $signed(buffer_5_11); // @[Modules.scala 160:64:@54220.4]
  assign _T_1207 = _T_1206[5:0]; // @[Modules.scala 160:64:@54221.4]
  assign buffer_5_12 = $signed(_T_1207); // @[Modules.scala 160:64:@54222.4]
  assign _T_1220 = $signed(_T_867) + $signed(_T_936); // @[Modules.scala 143:103:@54235.4]
  assign _T_1221 = _T_1220[3:0]; // @[Modules.scala 143:103:@54236.4]
  assign _T_1222 = $signed(_T_1221); // @[Modules.scala 143:103:@54237.4]
  assign _T_1248 = $signed(_T_830) + $signed(_T_837); // @[Modules.scala 143:103:@54259.4]
  assign _T_1249 = _T_1248[3:0]; // @[Modules.scala 143:103:@54260.4]
  assign _T_1250 = $signed(_T_1249); // @[Modules.scala 143:103:@54261.4]
  assign buffer_6_1 = {{2{_T_1222[3]}},_T_1222}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1251 = $signed(buffer_4_0) + $signed(buffer_6_1); // @[Modules.scala 160:64:@54263.4]
  assign _T_1252 = _T_1251[5:0]; // @[Modules.scala 160:64:@54264.4]
  assign buffer_6_6 = $signed(_T_1252); // @[Modules.scala 160:64:@54265.4]
  assign _T_1254 = $signed(buffer_0_2) + $signed(buffer_2_3); // @[Modules.scala 160:64:@54267.4]
  assign _T_1255 = _T_1254[5:0]; // @[Modules.scala 160:64:@54268.4]
  assign buffer_6_7 = $signed(_T_1255); // @[Modules.scala 160:64:@54269.4]
  assign buffer_6_5 = {{2{_T_1250[3]}},_T_1250}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1257 = $signed(buffer_4_5) + $signed(buffer_6_5); // @[Modules.scala 160:64:@54271.4]
  assign _T_1258 = _T_1257[5:0]; // @[Modules.scala 160:64:@54272.4]
  assign buffer_6_8 = $signed(_T_1258); // @[Modules.scala 160:64:@54273.4]
  assign _T_1260 = $signed(buffer_6_6) + $signed(buffer_6_7); // @[Modules.scala 166:64:@54275.4]
  assign _T_1261 = _T_1260[5:0]; // @[Modules.scala 166:64:@54276.4]
  assign buffer_6_9 = $signed(_T_1261); // @[Modules.scala 166:64:@54277.4]
  assign _T_1263 = $signed(buffer_6_9) + $signed(buffer_6_8); // @[Modules.scala 172:66:@54279.4]
  assign _T_1264 = _T_1263[5:0]; // @[Modules.scala 172:66:@54280.4]
  assign buffer_6_10 = $signed(_T_1264); // @[Modules.scala 172:66:@54281.4]
  assign _T_1284 = $signed(_T_934) + $signed(_T_802); // @[Modules.scala 150:103:@54302.4]
  assign _T_1285 = _T_1284[2:0]; // @[Modules.scala 150:103:@54303.4]
  assign _T_1286 = $signed(_T_1285); // @[Modules.scala 150:103:@54304.4]
  assign _GEN_20 = {{1{_T_888[2]}},_T_888}; // @[Modules.scala 150:103:@54308.4]
  assign _T_1291 = $signed(_T_941) + $signed(_GEN_20); // @[Modules.scala 150:103:@54308.4]
  assign _T_1292 = _T_1291[3:0]; // @[Modules.scala 150:103:@54309.4]
  assign _T_1293 = $signed(_T_1292); // @[Modules.scala 150:103:@54310.4]
  assign _T_1298 = $signed(_T_821) + $signed(_T_895); // @[Modules.scala 150:103:@54314.4]
  assign _T_1299 = _T_1298[3:0]; // @[Modules.scala 150:103:@54315.4]
  assign _T_1300 = $signed(_T_1299); // @[Modules.scala 150:103:@54316.4]
  assign _T_1310 = $signed(buffer_1_0) + $signed(buffer_4_1); // @[Modules.scala 166:64:@54326.4]
  assign _T_1311 = _T_1310[5:0]; // @[Modules.scala 166:64:@54327.4]
  assign buffer_7_7 = $signed(_T_1311); // @[Modules.scala 166:64:@54328.4]
  assign buffer_7_2 = {{3{_T_1286[2]}},_T_1286}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_7_3 = {{2{_T_1293[3]}},_T_1293}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1313 = $signed(buffer_7_2) + $signed(buffer_7_3); // @[Modules.scala 166:64:@54330.4]
  assign _T_1314 = _T_1313[5:0]; // @[Modules.scala 166:64:@54331.4]
  assign buffer_7_8 = $signed(_T_1314); // @[Modules.scala 166:64:@54332.4]
  assign buffer_7_4 = {{2{_T_1300[3]}},_T_1300}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1316 = $signed(buffer_7_4) + $signed(buffer_2_5); // @[Modules.scala 166:64:@54334.4]
  assign _T_1317 = _T_1316[5:0]; // @[Modules.scala 166:64:@54335.4]
  assign buffer_7_9 = $signed(_T_1317); // @[Modules.scala 166:64:@54336.4]
  assign _T_1319 = $signed(buffer_7_7) + $signed(buffer_7_8); // @[Modules.scala 166:64:@54338.4]
  assign _T_1320 = _T_1319[5:0]; // @[Modules.scala 166:64:@54339.4]
  assign buffer_7_10 = $signed(_T_1320); // @[Modules.scala 166:64:@54340.4]
  assign buffer_7_6 = {{2{_T_835[3]}},_T_835}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1322 = $signed(buffer_7_9) + $signed(buffer_7_6); // @[Modules.scala 172:66:@54342.4]
  assign _T_1323 = _T_1322[5:0]; // @[Modules.scala 172:66:@54343.4]
  assign buffer_7_11 = $signed(_T_1323); // @[Modules.scala 172:66:@54344.4]
  assign _T_1325 = $signed(buffer_7_10) + $signed(buffer_7_11); // @[Modules.scala 160:64:@54346.4]
  assign _T_1326 = _T_1325[5:0]; // @[Modules.scala 160:64:@54347.4]
  assign buffer_7_12 = $signed(_T_1326); // @[Modules.scala 160:64:@54348.4]
  assign _GEN_22 = {{1{_T_793[2]}},_T_793}; // @[Modules.scala 143:103:@54355.4]
  assign _T_1332 = $signed(_GEN_22) + $signed(_T_927); // @[Modules.scala 143:103:@54355.4]
  assign _T_1333 = _T_1332[3:0]; // @[Modules.scala 143:103:@54356.4]
  assign _T_1334 = $signed(_T_1333); // @[Modules.scala 143:103:@54357.4]
  assign _GEN_23 = {{1{_T_802[2]}},_T_802}; // @[Modules.scala 143:103:@54367.4]
  assign _T_1346 = $signed(_T_1008) + $signed(_GEN_23); // @[Modules.scala 143:103:@54367.4]
  assign _T_1347 = _T_1346[3:0]; // @[Modules.scala 143:103:@54368.4]
  assign _T_1348 = $signed(_T_1347); // @[Modules.scala 143:103:@54369.4]
  assign _T_1360 = $signed(_T_814) + $signed(_T_823); // @[Modules.scala 143:103:@54379.4]
  assign _T_1361 = _T_1360[2:0]; // @[Modules.scala 143:103:@54380.4]
  assign _T_1362 = $signed(_T_1361); // @[Modules.scala 143:103:@54381.4]
  assign _T_1367 = $signed(_T_897) + $signed(_T_902); // @[Modules.scala 143:103:@54385.4]
  assign _T_1368 = _T_1367[2:0]; // @[Modules.scala 143:103:@54386.4]
  assign _T_1369 = $signed(_T_1368); // @[Modules.scala 143:103:@54387.4]
  assign buffer_8_0 = {{2{_T_1334[3]}},_T_1334}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1370 = $signed(buffer_8_0) + $signed(buffer_1_1); // @[Modules.scala 160:64:@54389.4]
  assign _T_1371 = _T_1370[5:0]; // @[Modules.scala 160:64:@54390.4]
  assign buffer_8_6 = $signed(_T_1371); // @[Modules.scala 160:64:@54391.4]
  assign buffer_8_2 = {{2{_T_1348[3]}},_T_1348}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1373 = $signed(buffer_8_2) + $signed(buffer_2_2); // @[Modules.scala 160:64:@54393.4]
  assign _T_1374 = _T_1373[5:0]; // @[Modules.scala 160:64:@54394.4]
  assign buffer_8_7 = $signed(_T_1374); // @[Modules.scala 160:64:@54395.4]
  assign buffer_8_4 = {{3{_T_1362[2]}},_T_1362}; // @[Modules.scala 112:22:@53800.4]
  assign buffer_8_5 = {{3{_T_1369[2]}},_T_1369}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1376 = $signed(buffer_8_4) + $signed(buffer_8_5); // @[Modules.scala 160:64:@54397.4]
  assign _T_1377 = _T_1376[5:0]; // @[Modules.scala 160:64:@54398.4]
  assign buffer_8_8 = $signed(_T_1377); // @[Modules.scala 160:64:@54399.4]
  assign _T_1379 = $signed(buffer_8_6) + $signed(buffer_8_7); // @[Modules.scala 166:64:@54401.4]
  assign _T_1380 = _T_1379[5:0]; // @[Modules.scala 166:64:@54402.4]
  assign buffer_8_9 = $signed(_T_1380); // @[Modules.scala 166:64:@54403.4]
  assign _T_1382 = $signed(buffer_8_9) + $signed(buffer_8_8); // @[Modules.scala 172:66:@54405.4]
  assign _T_1383 = _T_1382[5:0]; // @[Modules.scala 172:66:@54406.4]
  assign buffer_8_10 = $signed(_T_1383); // @[Modules.scala 172:66:@54407.4]
  assign _T_1431 = $signed(_T_830) + $signed(_T_835); // @[Modules.scala 150:103:@54452.4]
  assign _T_1432 = _T_1431[3:0]; // @[Modules.scala 150:103:@54453.4]
  assign _T_1433 = $signed(_T_1432); // @[Modules.scala 150:103:@54454.4]
  assign _T_1439 = $signed(buffer_8_2) + $signed(buffer_4_3); // @[Modules.scala 160:64:@54462.4]
  assign _T_1440 = _T_1439[5:0]; // @[Modules.scala 160:64:@54463.4]
  assign buffer_9_9 = $signed(_T_1440); // @[Modules.scala 160:64:@54464.4]
  assign _T_1442 = $signed(buffer_4_4) + $signed(buffer_1_5); // @[Modules.scala 160:64:@54466.4]
  assign _T_1443 = _T_1442[5:0]; // @[Modules.scala 160:64:@54467.4]
  assign buffer_9_10 = $signed(_T_1443); // @[Modules.scala 160:64:@54468.4]
  assign buffer_9_6 = {{2{_T_1433[3]}},_T_1433}; // @[Modules.scala 112:22:@53800.4]
  assign _T_1445 = $signed(buffer_9_6) + $signed(buffer_3_7); // @[Modules.scala 160:64:@54470.4]
  assign _T_1446 = _T_1445[5:0]; // @[Modules.scala 160:64:@54471.4]
  assign buffer_9_11 = $signed(_T_1446); // @[Modules.scala 160:64:@54472.4]
  assign _T_1448 = $signed(buffer_4_8) + $signed(buffer_9_9); // @[Modules.scala 160:64:@54474.4]
  assign _T_1449 = _T_1448[5:0]; // @[Modules.scala 160:64:@54475.4]
  assign buffer_9_12 = $signed(_T_1449); // @[Modules.scala 160:64:@54476.4]
  assign _T_1451 = $signed(buffer_9_10) + $signed(buffer_9_11); // @[Modules.scala 160:64:@54478.4]
  assign _T_1452 = _T_1451[5:0]; // @[Modules.scala 160:64:@54479.4]
  assign buffer_9_13 = $signed(_T_1452); // @[Modules.scala 160:64:@54480.4]
  assign _T_1454 = $signed(buffer_9_12) + $signed(buffer_9_13); // @[Modules.scala 160:64:@54482.4]
  assign _T_1455 = _T_1454[5:0]; // @[Modules.scala 160:64:@54483.4]
  assign buffer_9_14 = $signed(_T_1455); // @[Modules.scala 160:64:@54484.4]
  assign io_out_0 = buffer_0_12;
  assign io_out_1 = buffer_1_12;
  assign io_out_2 = buffer_2_12;
  assign io_out_3 = buffer_3_14;
  assign io_out_4 = buffer_4_14;
  assign io_out_5 = buffer_5_12;
  assign io_out_6 = buffer_6_10;
  assign io_out_7 = buffer_7_12;
  assign io_out_8 = buffer_8_10;
  assign io_out_9 = buffer_9_14;
endmodule
module SBN_2( // @[:@54488.2]
  input  [5:0] io_in_0, // @[:@54491.4]
  input  [5:0] io_in_1, // @[:@54491.4]
  input  [5:0] io_in_2, // @[:@54491.4]
  input  [5:0] io_in_3, // @[:@54491.4]
  input  [5:0] io_in_4, // @[:@54491.4]
  input  [5:0] io_in_5, // @[:@54491.4]
  input  [5:0] io_in_6, // @[:@54491.4]
  input  [5:0] io_in_7, // @[:@54491.4]
  input  [5:0] io_in_8, // @[:@54491.4]
  input  [5:0] io_in_9, // @[:@54491.4]
  output [5:0] io_out_0, // @[:@54491.4]
  output [5:0] io_out_1, // @[:@54491.4]
  output [5:0] io_out_2, // @[:@54491.4]
  output [5:0] io_out_3, // @[:@54491.4]
  output [5:0] io_out_4, // @[:@54491.4]
  output [5:0] io_out_5, // @[:@54491.4]
  output [5:0] io_out_6, // @[:@54491.4]
  output [5:0] io_out_7, // @[:@54491.4]
  output [5:0] io_out_8, // @[:@54491.4]
  output [5:0] io_out_9 // @[:@54491.4]
);
  wire [6:0] _T_63; // @[Modules.scala 264:28:@54495.4]
  wire [5:0] _T_64; // @[Modules.scala 264:28:@54496.4]
  wire [5:0] c_x_0; // @[Modules.scala 264:28:@54497.4]
  wire [5:0] x_hat_0; // @[Modules.scala 269:32:@54499.4]
  wire [6:0] _T_69; // @[Modules.scala 271:31:@54501.4]
  wire [5:0] _T_70; // @[Modules.scala 271:31:@54502.4]
  wire [5:0] _T_71; // @[Modules.scala 271:31:@54503.4]
  wire [6:0] _T_73; // @[Modules.scala 264:28:@54505.4]
  wire [5:0] _T_74; // @[Modules.scala 264:28:@54506.4]
  wire [5:0] c_x_1; // @[Modules.scala 264:28:@54507.4]
  wire [5:0] x_hat_1; // @[Modules.scala 269:32:@54509.4]
  wire [6:0] _T_79; // @[Modules.scala 271:31:@54511.4]
  wire [5:0] _T_80; // @[Modules.scala 271:31:@54512.4]
  wire [5:0] _T_81; // @[Modules.scala 271:31:@54513.4]
  wire [6:0] _T_83; // @[Modules.scala 264:28:@54515.4]
  wire [5:0] _T_84; // @[Modules.scala 264:28:@54516.4]
  wire [5:0] c_x_2; // @[Modules.scala 264:28:@54517.4]
  wire [5:0] x_hat_2; // @[Modules.scala 269:32:@54519.4]
  wire [6:0] _T_89; // @[Modules.scala 271:31:@54521.4]
  wire [5:0] _T_90; // @[Modules.scala 271:31:@54522.4]
  wire [5:0] _T_91; // @[Modules.scala 271:31:@54523.4]
  wire [6:0] _T_93; // @[Modules.scala 264:28:@54525.4]
  wire [5:0] _T_94; // @[Modules.scala 264:28:@54526.4]
  wire [5:0] c_x_3; // @[Modules.scala 264:28:@54527.4]
  wire [5:0] x_hat_3; // @[Modules.scala 269:32:@54529.4]
  wire [6:0] _T_99; // @[Modules.scala 271:31:@54531.4]
  wire [5:0] _T_100; // @[Modules.scala 271:31:@54532.4]
  wire [5:0] _T_101; // @[Modules.scala 271:31:@54533.4]
  wire [6:0] _T_103; // @[Modules.scala 264:28:@54535.4]
  wire [5:0] _T_104; // @[Modules.scala 264:28:@54536.4]
  wire [5:0] c_x_4; // @[Modules.scala 264:28:@54537.4]
  wire [5:0] x_hat_4; // @[Modules.scala 269:32:@54539.4]
  wire [6:0] _T_109; // @[Modules.scala 271:31:@54541.4]
  wire [5:0] _T_110; // @[Modules.scala 271:31:@54542.4]
  wire [5:0] _T_111; // @[Modules.scala 271:31:@54543.4]
  wire [6:0] _T_113; // @[Modules.scala 264:28:@54545.4]
  wire [5:0] _T_114; // @[Modules.scala 264:28:@54546.4]
  wire [5:0] c_x_5; // @[Modules.scala 264:28:@54547.4]
  wire [5:0] x_hat_5; // @[Modules.scala 269:32:@54549.4]
  wire [6:0] _T_119; // @[Modules.scala 271:31:@54551.4]
  wire [5:0] _T_120; // @[Modules.scala 271:31:@54552.4]
  wire [5:0] _T_121; // @[Modules.scala 271:31:@54553.4]
  wire [6:0] _T_123; // @[Modules.scala 264:28:@54555.4]
  wire [5:0] _T_124; // @[Modules.scala 264:28:@54556.4]
  wire [5:0] c_x_6; // @[Modules.scala 264:28:@54557.4]
  wire [5:0] x_hat_6; // @[Modules.scala 269:32:@54559.4]
  wire [6:0] _T_129; // @[Modules.scala 271:31:@54561.4]
  wire [5:0] _T_130; // @[Modules.scala 271:31:@54562.4]
  wire [5:0] _T_131; // @[Modules.scala 271:31:@54563.4]
  wire [6:0] _T_133; // @[Modules.scala 264:28:@54565.4]
  wire [5:0] _T_134; // @[Modules.scala 264:28:@54566.4]
  wire [5:0] c_x_7; // @[Modules.scala 264:28:@54567.4]
  wire [20:0] _GEN_0; // @[Modules.scala 266:32:@54569.4]
  wire [20:0] _T_137; // @[Modules.scala 266:32:@54569.4]
  wire [5:0] _GEN_1; // @[Modules.scala 262:21:@54494.4]
  wire [5:0] x_hat_7; // @[Modules.scala 262:21:@54494.4]
  wire [6:0] _T_139; // @[Modules.scala 271:31:@54571.4]
  wire [5:0] _T_140; // @[Modules.scala 271:31:@54572.4]
  wire [5:0] _T_141; // @[Modules.scala 271:31:@54573.4]
  wire [6:0] _T_143; // @[Modules.scala 264:28:@54575.4]
  wire [5:0] _T_144; // @[Modules.scala 264:28:@54576.4]
  wire [5:0] c_x_8; // @[Modules.scala 264:28:@54577.4]
  wire [5:0] x_hat_8; // @[Modules.scala 269:32:@54579.4]
  wire [6:0] _T_149; // @[Modules.scala 271:31:@54581.4]
  wire [5:0] _T_150; // @[Modules.scala 271:31:@54582.4]
  wire [5:0] _T_151; // @[Modules.scala 271:31:@54583.4]
  wire [6:0] _T_153; // @[Modules.scala 264:28:@54585.4]
  wire [5:0] _T_154; // @[Modules.scala 264:28:@54586.4]
  wire [5:0] c_x_9; // @[Modules.scala 264:28:@54587.4]
  wire [5:0] x_hat_9; // @[Modules.scala 269:32:@54589.4]
  wire [6:0] _T_159; // @[Modules.scala 271:31:@54591.4]
  wire [5:0] _T_160; // @[Modules.scala 271:31:@54592.4]
  wire [5:0] _T_161; // @[Modules.scala 271:31:@54593.4]
  assign _T_63 = $signed(io_in_0) - $signed(6'sh0); // @[Modules.scala 264:28:@54495.4]
  assign _T_64 = _T_63[5:0]; // @[Modules.scala 264:28:@54496.4]
  assign c_x_0 = $signed(_T_64); // @[Modules.scala 264:28:@54497.4]
  assign x_hat_0 = $signed(c_x_0) >>> 4'h1; // @[Modules.scala 269:32:@54499.4]
  assign _T_69 = $signed(x_hat_0) + $signed(-6'sh1); // @[Modules.scala 271:31:@54501.4]
  assign _T_70 = _T_69[5:0]; // @[Modules.scala 271:31:@54502.4]
  assign _T_71 = $signed(_T_70); // @[Modules.scala 271:31:@54503.4]
  assign _T_73 = $signed(io_in_1) - $signed(6'sh1); // @[Modules.scala 264:28:@54505.4]
  assign _T_74 = _T_73[5:0]; // @[Modules.scala 264:28:@54506.4]
  assign c_x_1 = $signed(_T_74); // @[Modules.scala 264:28:@54507.4]
  assign x_hat_1 = $signed(c_x_1) >>> 4'h1; // @[Modules.scala 269:32:@54509.4]
  assign _T_79 = $signed(x_hat_1) + $signed(6'sh0); // @[Modules.scala 271:31:@54511.4]
  assign _T_80 = _T_79[5:0]; // @[Modules.scala 271:31:@54512.4]
  assign _T_81 = $signed(_T_80); // @[Modules.scala 271:31:@54513.4]
  assign _T_83 = $signed(io_in_2) - $signed(6'sh0); // @[Modules.scala 264:28:@54515.4]
  assign _T_84 = _T_83[5:0]; // @[Modules.scala 264:28:@54516.4]
  assign c_x_2 = $signed(_T_84); // @[Modules.scala 264:28:@54517.4]
  assign x_hat_2 = $signed(c_x_2) >>> 4'h1; // @[Modules.scala 269:32:@54519.4]
  assign _T_89 = $signed(x_hat_2) + $signed(6'sh0); // @[Modules.scala 271:31:@54521.4]
  assign _T_90 = _T_89[5:0]; // @[Modules.scala 271:31:@54522.4]
  assign _T_91 = $signed(_T_90); // @[Modules.scala 271:31:@54523.4]
  assign _T_93 = $signed(io_in_3) - $signed(6'sh0); // @[Modules.scala 264:28:@54525.4]
  assign _T_94 = _T_93[5:0]; // @[Modules.scala 264:28:@54526.4]
  assign c_x_3 = $signed(_T_94); // @[Modules.scala 264:28:@54527.4]
  assign x_hat_3 = $signed(c_x_3) >>> 4'h1; // @[Modules.scala 269:32:@54529.4]
  assign _T_99 = $signed(x_hat_3) + $signed(6'sh0); // @[Modules.scala 271:31:@54531.4]
  assign _T_100 = _T_99[5:0]; // @[Modules.scala 271:31:@54532.4]
  assign _T_101 = $signed(_T_100); // @[Modules.scala 271:31:@54533.4]
  assign _T_103 = $signed(io_in_4) - $signed(6'sh1); // @[Modules.scala 264:28:@54535.4]
  assign _T_104 = _T_103[5:0]; // @[Modules.scala 264:28:@54536.4]
  assign c_x_4 = $signed(_T_104); // @[Modules.scala 264:28:@54537.4]
  assign x_hat_4 = $signed(c_x_4) >>> 4'h1; // @[Modules.scala 269:32:@54539.4]
  assign _T_109 = $signed(x_hat_4) + $signed(6'sh0); // @[Modules.scala 271:31:@54541.4]
  assign _T_110 = _T_109[5:0]; // @[Modules.scala 271:31:@54542.4]
  assign _T_111 = $signed(_T_110); // @[Modules.scala 271:31:@54543.4]
  assign _T_113 = $signed(io_in_5) - $signed(6'sh0); // @[Modules.scala 264:28:@54545.4]
  assign _T_114 = _T_113[5:0]; // @[Modules.scala 264:28:@54546.4]
  assign c_x_5 = $signed(_T_114); // @[Modules.scala 264:28:@54547.4]
  assign x_hat_5 = $signed(c_x_5) >>> 4'h1; // @[Modules.scala 269:32:@54549.4]
  assign _T_119 = $signed(x_hat_5) + $signed(6'sh0); // @[Modules.scala 271:31:@54551.4]
  assign _T_120 = _T_119[5:0]; // @[Modules.scala 271:31:@54552.4]
  assign _T_121 = $signed(_T_120); // @[Modules.scala 271:31:@54553.4]
  assign _T_123 = $signed(io_in_6) - $signed(6'sh0); // @[Modules.scala 264:28:@54555.4]
  assign _T_124 = _T_123[5:0]; // @[Modules.scala 264:28:@54556.4]
  assign c_x_6 = $signed(_T_124); // @[Modules.scala 264:28:@54557.4]
  assign x_hat_6 = $signed(c_x_6) >>> 4'h1; // @[Modules.scala 269:32:@54559.4]
  assign _T_129 = $signed(x_hat_6) + $signed(6'sh0); // @[Modules.scala 271:31:@54561.4]
  assign _T_130 = _T_129[5:0]; // @[Modules.scala 271:31:@54562.4]
  assign _T_131 = $signed(_T_130); // @[Modules.scala 271:31:@54563.4]
  assign _T_133 = $signed(io_in_7) - $signed(6'sh0); // @[Modules.scala 264:28:@54565.4]
  assign _T_134 = _T_133[5:0]; // @[Modules.scala 264:28:@54566.4]
  assign c_x_7 = $signed(_T_134); // @[Modules.scala 264:28:@54567.4]
  assign _GEN_0 = {{15{c_x_7[5]}},c_x_7}; // @[Modules.scala 266:32:@54569.4]
  assign _T_137 = $signed(_GEN_0) << 4'h0; // @[Modules.scala 266:32:@54569.4]
  assign _GEN_1 = _T_137[5:0]; // @[Modules.scala 262:21:@54494.4]
  assign x_hat_7 = $signed(_GEN_1); // @[Modules.scala 262:21:@54494.4]
  assign _T_139 = $signed(x_hat_7) + $signed(6'sh0); // @[Modules.scala 271:31:@54571.4]
  assign _T_140 = _T_139[5:0]; // @[Modules.scala 271:31:@54572.4]
  assign _T_141 = $signed(_T_140); // @[Modules.scala 271:31:@54573.4]
  assign _T_143 = $signed(io_in_8) - $signed(6'sh0); // @[Modules.scala 264:28:@54575.4]
  assign _T_144 = _T_143[5:0]; // @[Modules.scala 264:28:@54576.4]
  assign c_x_8 = $signed(_T_144); // @[Modules.scala 264:28:@54577.4]
  assign x_hat_8 = $signed(c_x_8) >>> 4'h1; // @[Modules.scala 269:32:@54579.4]
  assign _T_149 = $signed(x_hat_8) + $signed(6'sh0); // @[Modules.scala 271:31:@54581.4]
  assign _T_150 = _T_149[5:0]; // @[Modules.scala 271:31:@54582.4]
  assign _T_151 = $signed(_T_150); // @[Modules.scala 271:31:@54583.4]
  assign _T_153 = $signed(io_in_9) - $signed(6'sh1); // @[Modules.scala 264:28:@54585.4]
  assign _T_154 = _T_153[5:0]; // @[Modules.scala 264:28:@54586.4]
  assign c_x_9 = $signed(_T_154); // @[Modules.scala 264:28:@54587.4]
  assign x_hat_9 = $signed(c_x_9) >>> 4'h1; // @[Modules.scala 269:32:@54589.4]
  assign _T_159 = $signed(x_hat_9) + $signed(6'sh0); // @[Modules.scala 271:31:@54591.4]
  assign _T_160 = _T_159[5:0]; // @[Modules.scala 271:31:@54592.4]
  assign _T_161 = $signed(_T_160); // @[Modules.scala 271:31:@54593.4]
  assign io_out_0 = _T_71;
  assign io_out_1 = _T_81;
  assign io_out_2 = _T_91;
  assign io_out_3 = _T_101;
  assign io_out_4 = _T_111;
  assign io_out_5 = _T_121;
  assign io_out_6 = _T_131;
  assign io_out_7 = _T_141;
  assign io_out_8 = _T_151;
  assign io_out_9 = _T_161;
endmodule
module MLP( // @[:@54596.2]
  input        clock, // @[:@54597.4]
  input        reset, // @[:@54598.4]
  input  [3:0] io_in_0, // @[:@54599.4]
  input  [3:0] io_in_1, // @[:@54599.4]
  input  [3:0] io_in_2, // @[:@54599.4]
  input  [3:0] io_in_3, // @[:@54599.4]
  input  [3:0] io_in_4, // @[:@54599.4]
  input  [3:0] io_in_5, // @[:@54599.4]
  input  [3:0] io_in_6, // @[:@54599.4]
  input  [3:0] io_in_7, // @[:@54599.4]
  input  [3:0] io_in_8, // @[:@54599.4]
  input  [3:0] io_in_9, // @[:@54599.4]
  input  [3:0] io_in_10, // @[:@54599.4]
  input  [3:0] io_in_11, // @[:@54599.4]
  input  [3:0] io_in_12, // @[:@54599.4]
  input  [3:0] io_in_13, // @[:@54599.4]
  input  [3:0] io_in_14, // @[:@54599.4]
  input  [3:0] io_in_15, // @[:@54599.4]
  input  [3:0] io_in_16, // @[:@54599.4]
  input  [3:0] io_in_17, // @[:@54599.4]
  input  [3:0] io_in_18, // @[:@54599.4]
  input  [3:0] io_in_19, // @[:@54599.4]
  input  [3:0] io_in_20, // @[:@54599.4]
  input  [3:0] io_in_21, // @[:@54599.4]
  input  [3:0] io_in_22, // @[:@54599.4]
  input  [3:0] io_in_23, // @[:@54599.4]
  input  [3:0] io_in_24, // @[:@54599.4]
  input  [3:0] io_in_25, // @[:@54599.4]
  input  [3:0] io_in_26, // @[:@54599.4]
  input  [3:0] io_in_27, // @[:@54599.4]
  input  [3:0] io_in_28, // @[:@54599.4]
  input  [3:0] io_in_29, // @[:@54599.4]
  input  [3:0] io_in_30, // @[:@54599.4]
  input  [3:0] io_in_31, // @[:@54599.4]
  input  [3:0] io_in_32, // @[:@54599.4]
  input  [3:0] io_in_33, // @[:@54599.4]
  input  [3:0] io_in_34, // @[:@54599.4]
  input  [3:0] io_in_35, // @[:@54599.4]
  input  [3:0] io_in_36, // @[:@54599.4]
  input  [3:0] io_in_37, // @[:@54599.4]
  input  [3:0] io_in_38, // @[:@54599.4]
  input  [3:0] io_in_39, // @[:@54599.4]
  input  [3:0] io_in_40, // @[:@54599.4]
  input  [3:0] io_in_41, // @[:@54599.4]
  input  [3:0] io_in_42, // @[:@54599.4]
  input  [3:0] io_in_43, // @[:@54599.4]
  input  [3:0] io_in_44, // @[:@54599.4]
  input  [3:0] io_in_45, // @[:@54599.4]
  input  [3:0] io_in_46, // @[:@54599.4]
  input  [3:0] io_in_47, // @[:@54599.4]
  input  [3:0] io_in_48, // @[:@54599.4]
  input  [3:0] io_in_49, // @[:@54599.4]
  input  [3:0] io_in_50, // @[:@54599.4]
  input  [3:0] io_in_51, // @[:@54599.4]
  input  [3:0] io_in_52, // @[:@54599.4]
  input  [3:0] io_in_53, // @[:@54599.4]
  input  [3:0] io_in_54, // @[:@54599.4]
  input  [3:0] io_in_55, // @[:@54599.4]
  input  [3:0] io_in_56, // @[:@54599.4]
  input  [3:0] io_in_57, // @[:@54599.4]
  input  [3:0] io_in_58, // @[:@54599.4]
  input  [3:0] io_in_59, // @[:@54599.4]
  input  [3:0] io_in_60, // @[:@54599.4]
  input  [3:0] io_in_61, // @[:@54599.4]
  input  [3:0] io_in_62, // @[:@54599.4]
  input  [3:0] io_in_63, // @[:@54599.4]
  input  [3:0] io_in_64, // @[:@54599.4]
  input  [3:0] io_in_65, // @[:@54599.4]
  input  [3:0] io_in_66, // @[:@54599.4]
  input  [3:0] io_in_67, // @[:@54599.4]
  input  [3:0] io_in_68, // @[:@54599.4]
  input  [3:0] io_in_69, // @[:@54599.4]
  input  [3:0] io_in_70, // @[:@54599.4]
  input  [3:0] io_in_71, // @[:@54599.4]
  input  [3:0] io_in_72, // @[:@54599.4]
  input  [3:0] io_in_73, // @[:@54599.4]
  input  [3:0] io_in_74, // @[:@54599.4]
  input  [3:0] io_in_75, // @[:@54599.4]
  input  [3:0] io_in_76, // @[:@54599.4]
  input  [3:0] io_in_77, // @[:@54599.4]
  input  [3:0] io_in_78, // @[:@54599.4]
  input  [3:0] io_in_79, // @[:@54599.4]
  input  [3:0] io_in_80, // @[:@54599.4]
  input  [3:0] io_in_81, // @[:@54599.4]
  input  [3:0] io_in_82, // @[:@54599.4]
  input  [3:0] io_in_83, // @[:@54599.4]
  input  [3:0] io_in_84, // @[:@54599.4]
  input  [3:0] io_in_85, // @[:@54599.4]
  input  [3:0] io_in_86, // @[:@54599.4]
  input  [3:0] io_in_87, // @[:@54599.4]
  input  [3:0] io_in_88, // @[:@54599.4]
  input  [3:0] io_in_89, // @[:@54599.4]
  input  [3:0] io_in_90, // @[:@54599.4]
  input  [3:0] io_in_91, // @[:@54599.4]
  input  [3:0] io_in_92, // @[:@54599.4]
  input  [3:0] io_in_93, // @[:@54599.4]
  input  [3:0] io_in_94, // @[:@54599.4]
  input  [3:0] io_in_95, // @[:@54599.4]
  input  [3:0] io_in_96, // @[:@54599.4]
  input  [3:0] io_in_97, // @[:@54599.4]
  input  [3:0] io_in_98, // @[:@54599.4]
  input  [3:0] io_in_99, // @[:@54599.4]
  input  [3:0] io_in_100, // @[:@54599.4]
  input  [3:0] io_in_101, // @[:@54599.4]
  input  [3:0] io_in_102, // @[:@54599.4]
  input  [3:0] io_in_103, // @[:@54599.4]
  input  [3:0] io_in_104, // @[:@54599.4]
  input  [3:0] io_in_105, // @[:@54599.4]
  input  [3:0] io_in_106, // @[:@54599.4]
  input  [3:0] io_in_107, // @[:@54599.4]
  input  [3:0] io_in_108, // @[:@54599.4]
  input  [3:0] io_in_109, // @[:@54599.4]
  input  [3:0] io_in_110, // @[:@54599.4]
  input  [3:0] io_in_111, // @[:@54599.4]
  input  [3:0] io_in_112, // @[:@54599.4]
  input  [3:0] io_in_113, // @[:@54599.4]
  input  [3:0] io_in_114, // @[:@54599.4]
  input  [3:0] io_in_115, // @[:@54599.4]
  input  [3:0] io_in_116, // @[:@54599.4]
  input  [3:0] io_in_117, // @[:@54599.4]
  input  [3:0] io_in_118, // @[:@54599.4]
  input  [3:0] io_in_119, // @[:@54599.4]
  input  [3:0] io_in_120, // @[:@54599.4]
  input  [3:0] io_in_121, // @[:@54599.4]
  input  [3:0] io_in_122, // @[:@54599.4]
  input  [3:0] io_in_123, // @[:@54599.4]
  input  [3:0] io_in_124, // @[:@54599.4]
  input  [3:0] io_in_125, // @[:@54599.4]
  input  [3:0] io_in_126, // @[:@54599.4]
  input  [3:0] io_in_127, // @[:@54599.4]
  input  [3:0] io_in_128, // @[:@54599.4]
  input  [3:0] io_in_129, // @[:@54599.4]
  input  [3:0] io_in_130, // @[:@54599.4]
  input  [3:0] io_in_131, // @[:@54599.4]
  input  [3:0] io_in_132, // @[:@54599.4]
  input  [3:0] io_in_133, // @[:@54599.4]
  input  [3:0] io_in_134, // @[:@54599.4]
  input  [3:0] io_in_135, // @[:@54599.4]
  input  [3:0] io_in_136, // @[:@54599.4]
  input  [3:0] io_in_137, // @[:@54599.4]
  input  [3:0] io_in_138, // @[:@54599.4]
  input  [3:0] io_in_139, // @[:@54599.4]
  input  [3:0] io_in_140, // @[:@54599.4]
  input  [3:0] io_in_141, // @[:@54599.4]
  input  [3:0] io_in_142, // @[:@54599.4]
  input  [3:0] io_in_143, // @[:@54599.4]
  input  [3:0] io_in_144, // @[:@54599.4]
  input  [3:0] io_in_145, // @[:@54599.4]
  input  [3:0] io_in_146, // @[:@54599.4]
  input  [3:0] io_in_147, // @[:@54599.4]
  input  [3:0] io_in_148, // @[:@54599.4]
  input  [3:0] io_in_149, // @[:@54599.4]
  input  [3:0] io_in_150, // @[:@54599.4]
  input  [3:0] io_in_151, // @[:@54599.4]
  input  [3:0] io_in_152, // @[:@54599.4]
  input  [3:0] io_in_153, // @[:@54599.4]
  input  [3:0] io_in_154, // @[:@54599.4]
  input  [3:0] io_in_155, // @[:@54599.4]
  input  [3:0] io_in_156, // @[:@54599.4]
  input  [3:0] io_in_157, // @[:@54599.4]
  input  [3:0] io_in_158, // @[:@54599.4]
  input  [3:0] io_in_159, // @[:@54599.4]
  input  [3:0] io_in_160, // @[:@54599.4]
  input  [3:0] io_in_161, // @[:@54599.4]
  input  [3:0] io_in_162, // @[:@54599.4]
  input  [3:0] io_in_163, // @[:@54599.4]
  input  [3:0] io_in_164, // @[:@54599.4]
  input  [3:0] io_in_165, // @[:@54599.4]
  input  [3:0] io_in_166, // @[:@54599.4]
  input  [3:0] io_in_167, // @[:@54599.4]
  input  [3:0] io_in_168, // @[:@54599.4]
  input  [3:0] io_in_169, // @[:@54599.4]
  input  [3:0] io_in_170, // @[:@54599.4]
  input  [3:0] io_in_171, // @[:@54599.4]
  input  [3:0] io_in_172, // @[:@54599.4]
  input  [3:0] io_in_173, // @[:@54599.4]
  input  [3:0] io_in_174, // @[:@54599.4]
  input  [3:0] io_in_175, // @[:@54599.4]
  input  [3:0] io_in_176, // @[:@54599.4]
  input  [3:0] io_in_177, // @[:@54599.4]
  input  [3:0] io_in_178, // @[:@54599.4]
  input  [3:0] io_in_179, // @[:@54599.4]
  input  [3:0] io_in_180, // @[:@54599.4]
  input  [3:0] io_in_181, // @[:@54599.4]
  input  [3:0] io_in_182, // @[:@54599.4]
  input  [3:0] io_in_183, // @[:@54599.4]
  input  [3:0] io_in_184, // @[:@54599.4]
  input  [3:0] io_in_185, // @[:@54599.4]
  input  [3:0] io_in_186, // @[:@54599.4]
  input  [3:0] io_in_187, // @[:@54599.4]
  input  [3:0] io_in_188, // @[:@54599.4]
  input  [3:0] io_in_189, // @[:@54599.4]
  input  [3:0] io_in_190, // @[:@54599.4]
  input  [3:0] io_in_191, // @[:@54599.4]
  input  [3:0] io_in_192, // @[:@54599.4]
  input  [3:0] io_in_193, // @[:@54599.4]
  input  [3:0] io_in_194, // @[:@54599.4]
  input  [3:0] io_in_195, // @[:@54599.4]
  input  [3:0] io_in_196, // @[:@54599.4]
  input  [3:0] io_in_197, // @[:@54599.4]
  input  [3:0] io_in_198, // @[:@54599.4]
  input  [3:0] io_in_199, // @[:@54599.4]
  input  [3:0] io_in_200, // @[:@54599.4]
  input  [3:0] io_in_201, // @[:@54599.4]
  input  [3:0] io_in_202, // @[:@54599.4]
  input  [3:0] io_in_203, // @[:@54599.4]
  input  [3:0] io_in_204, // @[:@54599.4]
  input  [3:0] io_in_205, // @[:@54599.4]
  input  [3:0] io_in_206, // @[:@54599.4]
  input  [3:0] io_in_207, // @[:@54599.4]
  input  [3:0] io_in_208, // @[:@54599.4]
  input  [3:0] io_in_209, // @[:@54599.4]
  input  [3:0] io_in_210, // @[:@54599.4]
  input  [3:0] io_in_211, // @[:@54599.4]
  input  [3:0] io_in_212, // @[:@54599.4]
  input  [3:0] io_in_213, // @[:@54599.4]
  input  [3:0] io_in_214, // @[:@54599.4]
  input  [3:0] io_in_215, // @[:@54599.4]
  input  [3:0] io_in_216, // @[:@54599.4]
  input  [3:0] io_in_217, // @[:@54599.4]
  input  [3:0] io_in_218, // @[:@54599.4]
  input  [3:0] io_in_219, // @[:@54599.4]
  input  [3:0] io_in_220, // @[:@54599.4]
  input  [3:0] io_in_221, // @[:@54599.4]
  input  [3:0] io_in_222, // @[:@54599.4]
  input  [3:0] io_in_223, // @[:@54599.4]
  input  [3:0] io_in_224, // @[:@54599.4]
  input  [3:0] io_in_225, // @[:@54599.4]
  input  [3:0] io_in_226, // @[:@54599.4]
  input  [3:0] io_in_227, // @[:@54599.4]
  input  [3:0] io_in_228, // @[:@54599.4]
  input  [3:0] io_in_229, // @[:@54599.4]
  input  [3:0] io_in_230, // @[:@54599.4]
  input  [3:0] io_in_231, // @[:@54599.4]
  input  [3:0] io_in_232, // @[:@54599.4]
  input  [3:0] io_in_233, // @[:@54599.4]
  input  [3:0] io_in_234, // @[:@54599.4]
  input  [3:0] io_in_235, // @[:@54599.4]
  input  [3:0] io_in_236, // @[:@54599.4]
  input  [3:0] io_in_237, // @[:@54599.4]
  input  [3:0] io_in_238, // @[:@54599.4]
  input  [3:0] io_in_239, // @[:@54599.4]
  input  [3:0] io_in_240, // @[:@54599.4]
  input  [3:0] io_in_241, // @[:@54599.4]
  input  [3:0] io_in_242, // @[:@54599.4]
  input  [3:0] io_in_243, // @[:@54599.4]
  input  [3:0] io_in_244, // @[:@54599.4]
  input  [3:0] io_in_245, // @[:@54599.4]
  input  [3:0] io_in_246, // @[:@54599.4]
  input  [3:0] io_in_247, // @[:@54599.4]
  input  [3:0] io_in_248, // @[:@54599.4]
  input  [3:0] io_in_249, // @[:@54599.4]
  input  [3:0] io_in_250, // @[:@54599.4]
  input  [3:0] io_in_251, // @[:@54599.4]
  input  [3:0] io_in_252, // @[:@54599.4]
  input  [3:0] io_in_253, // @[:@54599.4]
  input  [3:0] io_in_254, // @[:@54599.4]
  input  [3:0] io_in_255, // @[:@54599.4]
  input  [3:0] io_in_256, // @[:@54599.4]
  input  [3:0] io_in_257, // @[:@54599.4]
  input  [3:0] io_in_258, // @[:@54599.4]
  input  [3:0] io_in_259, // @[:@54599.4]
  input  [3:0] io_in_260, // @[:@54599.4]
  input  [3:0] io_in_261, // @[:@54599.4]
  input  [3:0] io_in_262, // @[:@54599.4]
  input  [3:0] io_in_263, // @[:@54599.4]
  input  [3:0] io_in_264, // @[:@54599.4]
  input  [3:0] io_in_265, // @[:@54599.4]
  input  [3:0] io_in_266, // @[:@54599.4]
  input  [3:0] io_in_267, // @[:@54599.4]
  input  [3:0] io_in_268, // @[:@54599.4]
  input  [3:0] io_in_269, // @[:@54599.4]
  input  [3:0] io_in_270, // @[:@54599.4]
  input  [3:0] io_in_271, // @[:@54599.4]
  input  [3:0] io_in_272, // @[:@54599.4]
  input  [3:0] io_in_273, // @[:@54599.4]
  input  [3:0] io_in_274, // @[:@54599.4]
  input  [3:0] io_in_275, // @[:@54599.4]
  input  [3:0] io_in_276, // @[:@54599.4]
  input  [3:0] io_in_277, // @[:@54599.4]
  input  [3:0] io_in_278, // @[:@54599.4]
  input  [3:0] io_in_279, // @[:@54599.4]
  input  [3:0] io_in_280, // @[:@54599.4]
  input  [3:0] io_in_281, // @[:@54599.4]
  input  [3:0] io_in_282, // @[:@54599.4]
  input  [3:0] io_in_283, // @[:@54599.4]
  input  [3:0] io_in_284, // @[:@54599.4]
  input  [3:0] io_in_285, // @[:@54599.4]
  input  [3:0] io_in_286, // @[:@54599.4]
  input  [3:0] io_in_287, // @[:@54599.4]
  input  [3:0] io_in_288, // @[:@54599.4]
  input  [3:0] io_in_289, // @[:@54599.4]
  input  [3:0] io_in_290, // @[:@54599.4]
  input  [3:0] io_in_291, // @[:@54599.4]
  input  [3:0] io_in_292, // @[:@54599.4]
  input  [3:0] io_in_293, // @[:@54599.4]
  input  [3:0] io_in_294, // @[:@54599.4]
  input  [3:0] io_in_295, // @[:@54599.4]
  input  [3:0] io_in_296, // @[:@54599.4]
  input  [3:0] io_in_297, // @[:@54599.4]
  input  [3:0] io_in_298, // @[:@54599.4]
  input  [3:0] io_in_299, // @[:@54599.4]
  input  [3:0] io_in_300, // @[:@54599.4]
  input  [3:0] io_in_301, // @[:@54599.4]
  input  [3:0] io_in_302, // @[:@54599.4]
  input  [3:0] io_in_303, // @[:@54599.4]
  input  [3:0] io_in_304, // @[:@54599.4]
  input  [3:0] io_in_305, // @[:@54599.4]
  input  [3:0] io_in_306, // @[:@54599.4]
  input  [3:0] io_in_307, // @[:@54599.4]
  input  [3:0] io_in_308, // @[:@54599.4]
  input  [3:0] io_in_309, // @[:@54599.4]
  input  [3:0] io_in_310, // @[:@54599.4]
  input  [3:0] io_in_311, // @[:@54599.4]
  input  [3:0] io_in_312, // @[:@54599.4]
  input  [3:0] io_in_313, // @[:@54599.4]
  input  [3:0] io_in_314, // @[:@54599.4]
  input  [3:0] io_in_315, // @[:@54599.4]
  input  [3:0] io_in_316, // @[:@54599.4]
  input  [3:0] io_in_317, // @[:@54599.4]
  input  [3:0] io_in_318, // @[:@54599.4]
  input  [3:0] io_in_319, // @[:@54599.4]
  input  [3:0] io_in_320, // @[:@54599.4]
  input  [3:0] io_in_321, // @[:@54599.4]
  input  [3:0] io_in_322, // @[:@54599.4]
  input  [3:0] io_in_323, // @[:@54599.4]
  input  [3:0] io_in_324, // @[:@54599.4]
  input  [3:0] io_in_325, // @[:@54599.4]
  input  [3:0] io_in_326, // @[:@54599.4]
  input  [3:0] io_in_327, // @[:@54599.4]
  input  [3:0] io_in_328, // @[:@54599.4]
  input  [3:0] io_in_329, // @[:@54599.4]
  input  [3:0] io_in_330, // @[:@54599.4]
  input  [3:0] io_in_331, // @[:@54599.4]
  input  [3:0] io_in_332, // @[:@54599.4]
  input  [3:0] io_in_333, // @[:@54599.4]
  input  [3:0] io_in_334, // @[:@54599.4]
  input  [3:0] io_in_335, // @[:@54599.4]
  input  [3:0] io_in_336, // @[:@54599.4]
  input  [3:0] io_in_337, // @[:@54599.4]
  input  [3:0] io_in_338, // @[:@54599.4]
  input  [3:0] io_in_339, // @[:@54599.4]
  input  [3:0] io_in_340, // @[:@54599.4]
  input  [3:0] io_in_341, // @[:@54599.4]
  input  [3:0] io_in_342, // @[:@54599.4]
  input  [3:0] io_in_343, // @[:@54599.4]
  input  [3:0] io_in_344, // @[:@54599.4]
  input  [3:0] io_in_345, // @[:@54599.4]
  input  [3:0] io_in_346, // @[:@54599.4]
  input  [3:0] io_in_347, // @[:@54599.4]
  input  [3:0] io_in_348, // @[:@54599.4]
  input  [3:0] io_in_349, // @[:@54599.4]
  input  [3:0] io_in_350, // @[:@54599.4]
  input  [3:0] io_in_351, // @[:@54599.4]
  input  [3:0] io_in_352, // @[:@54599.4]
  input  [3:0] io_in_353, // @[:@54599.4]
  input  [3:0] io_in_354, // @[:@54599.4]
  input  [3:0] io_in_355, // @[:@54599.4]
  input  [3:0] io_in_356, // @[:@54599.4]
  input  [3:0] io_in_357, // @[:@54599.4]
  input  [3:0] io_in_358, // @[:@54599.4]
  input  [3:0] io_in_359, // @[:@54599.4]
  input  [3:0] io_in_360, // @[:@54599.4]
  input  [3:0] io_in_361, // @[:@54599.4]
  input  [3:0] io_in_362, // @[:@54599.4]
  input  [3:0] io_in_363, // @[:@54599.4]
  input  [3:0] io_in_364, // @[:@54599.4]
  input  [3:0] io_in_365, // @[:@54599.4]
  input  [3:0] io_in_366, // @[:@54599.4]
  input  [3:0] io_in_367, // @[:@54599.4]
  input  [3:0] io_in_368, // @[:@54599.4]
  input  [3:0] io_in_369, // @[:@54599.4]
  input  [3:0] io_in_370, // @[:@54599.4]
  input  [3:0] io_in_371, // @[:@54599.4]
  input  [3:0] io_in_372, // @[:@54599.4]
  input  [3:0] io_in_373, // @[:@54599.4]
  input  [3:0] io_in_374, // @[:@54599.4]
  input  [3:0] io_in_375, // @[:@54599.4]
  input  [3:0] io_in_376, // @[:@54599.4]
  input  [3:0] io_in_377, // @[:@54599.4]
  input  [3:0] io_in_378, // @[:@54599.4]
  input  [3:0] io_in_379, // @[:@54599.4]
  input  [3:0] io_in_380, // @[:@54599.4]
  input  [3:0] io_in_381, // @[:@54599.4]
  input  [3:0] io_in_382, // @[:@54599.4]
  input  [3:0] io_in_383, // @[:@54599.4]
  input  [3:0] io_in_384, // @[:@54599.4]
  input  [3:0] io_in_385, // @[:@54599.4]
  input  [3:0] io_in_386, // @[:@54599.4]
  input  [3:0] io_in_387, // @[:@54599.4]
  input  [3:0] io_in_388, // @[:@54599.4]
  input  [3:0] io_in_389, // @[:@54599.4]
  input  [3:0] io_in_390, // @[:@54599.4]
  input  [3:0] io_in_391, // @[:@54599.4]
  input  [3:0] io_in_392, // @[:@54599.4]
  input  [3:0] io_in_393, // @[:@54599.4]
  input  [3:0] io_in_394, // @[:@54599.4]
  input  [3:0] io_in_395, // @[:@54599.4]
  input  [3:0] io_in_396, // @[:@54599.4]
  input  [3:0] io_in_397, // @[:@54599.4]
  input  [3:0] io_in_398, // @[:@54599.4]
  input  [3:0] io_in_399, // @[:@54599.4]
  input  [3:0] io_in_400, // @[:@54599.4]
  input  [3:0] io_in_401, // @[:@54599.4]
  input  [3:0] io_in_402, // @[:@54599.4]
  input  [3:0] io_in_403, // @[:@54599.4]
  input  [3:0] io_in_404, // @[:@54599.4]
  input  [3:0] io_in_405, // @[:@54599.4]
  input  [3:0] io_in_406, // @[:@54599.4]
  input  [3:0] io_in_407, // @[:@54599.4]
  input  [3:0] io_in_408, // @[:@54599.4]
  input  [3:0] io_in_409, // @[:@54599.4]
  input  [3:0] io_in_410, // @[:@54599.4]
  input  [3:0] io_in_411, // @[:@54599.4]
  input  [3:0] io_in_412, // @[:@54599.4]
  input  [3:0] io_in_413, // @[:@54599.4]
  input  [3:0] io_in_414, // @[:@54599.4]
  input  [3:0] io_in_415, // @[:@54599.4]
  input  [3:0] io_in_416, // @[:@54599.4]
  input  [3:0] io_in_417, // @[:@54599.4]
  input  [3:0] io_in_418, // @[:@54599.4]
  input  [3:0] io_in_419, // @[:@54599.4]
  input  [3:0] io_in_420, // @[:@54599.4]
  input  [3:0] io_in_421, // @[:@54599.4]
  input  [3:0] io_in_422, // @[:@54599.4]
  input  [3:0] io_in_423, // @[:@54599.4]
  input  [3:0] io_in_424, // @[:@54599.4]
  input  [3:0] io_in_425, // @[:@54599.4]
  input  [3:0] io_in_426, // @[:@54599.4]
  input  [3:0] io_in_427, // @[:@54599.4]
  input  [3:0] io_in_428, // @[:@54599.4]
  input  [3:0] io_in_429, // @[:@54599.4]
  input  [3:0] io_in_430, // @[:@54599.4]
  input  [3:0] io_in_431, // @[:@54599.4]
  input  [3:0] io_in_432, // @[:@54599.4]
  input  [3:0] io_in_433, // @[:@54599.4]
  input  [3:0] io_in_434, // @[:@54599.4]
  input  [3:0] io_in_435, // @[:@54599.4]
  input  [3:0] io_in_436, // @[:@54599.4]
  input  [3:0] io_in_437, // @[:@54599.4]
  input  [3:0] io_in_438, // @[:@54599.4]
  input  [3:0] io_in_439, // @[:@54599.4]
  input  [3:0] io_in_440, // @[:@54599.4]
  input  [3:0] io_in_441, // @[:@54599.4]
  input  [3:0] io_in_442, // @[:@54599.4]
  input  [3:0] io_in_443, // @[:@54599.4]
  input  [3:0] io_in_444, // @[:@54599.4]
  input  [3:0] io_in_445, // @[:@54599.4]
  input  [3:0] io_in_446, // @[:@54599.4]
  input  [3:0] io_in_447, // @[:@54599.4]
  input  [3:0] io_in_448, // @[:@54599.4]
  input  [3:0] io_in_449, // @[:@54599.4]
  input  [3:0] io_in_450, // @[:@54599.4]
  input  [3:0] io_in_451, // @[:@54599.4]
  input  [3:0] io_in_452, // @[:@54599.4]
  input  [3:0] io_in_453, // @[:@54599.4]
  input  [3:0] io_in_454, // @[:@54599.4]
  input  [3:0] io_in_455, // @[:@54599.4]
  input  [3:0] io_in_456, // @[:@54599.4]
  input  [3:0] io_in_457, // @[:@54599.4]
  input  [3:0] io_in_458, // @[:@54599.4]
  input  [3:0] io_in_459, // @[:@54599.4]
  input  [3:0] io_in_460, // @[:@54599.4]
  input  [3:0] io_in_461, // @[:@54599.4]
  input  [3:0] io_in_462, // @[:@54599.4]
  input  [3:0] io_in_463, // @[:@54599.4]
  input  [3:0] io_in_464, // @[:@54599.4]
  input  [3:0] io_in_465, // @[:@54599.4]
  input  [3:0] io_in_466, // @[:@54599.4]
  input  [3:0] io_in_467, // @[:@54599.4]
  input  [3:0] io_in_468, // @[:@54599.4]
  input  [3:0] io_in_469, // @[:@54599.4]
  input  [3:0] io_in_470, // @[:@54599.4]
  input  [3:0] io_in_471, // @[:@54599.4]
  input  [3:0] io_in_472, // @[:@54599.4]
  input  [3:0] io_in_473, // @[:@54599.4]
  input  [3:0] io_in_474, // @[:@54599.4]
  input  [3:0] io_in_475, // @[:@54599.4]
  input  [3:0] io_in_476, // @[:@54599.4]
  input  [3:0] io_in_477, // @[:@54599.4]
  input  [3:0] io_in_478, // @[:@54599.4]
  input  [3:0] io_in_479, // @[:@54599.4]
  input  [3:0] io_in_480, // @[:@54599.4]
  input  [3:0] io_in_481, // @[:@54599.4]
  input  [3:0] io_in_482, // @[:@54599.4]
  input  [3:0] io_in_483, // @[:@54599.4]
  input  [3:0] io_in_484, // @[:@54599.4]
  input  [3:0] io_in_485, // @[:@54599.4]
  input  [3:0] io_in_486, // @[:@54599.4]
  input  [3:0] io_in_487, // @[:@54599.4]
  input  [3:0] io_in_488, // @[:@54599.4]
  input  [3:0] io_in_489, // @[:@54599.4]
  input  [3:0] io_in_490, // @[:@54599.4]
  input  [3:0] io_in_491, // @[:@54599.4]
  input  [3:0] io_in_492, // @[:@54599.4]
  input  [3:0] io_in_493, // @[:@54599.4]
  input  [3:0] io_in_494, // @[:@54599.4]
  input  [3:0] io_in_495, // @[:@54599.4]
  input  [3:0] io_in_496, // @[:@54599.4]
  input  [3:0] io_in_497, // @[:@54599.4]
  input  [3:0] io_in_498, // @[:@54599.4]
  input  [3:0] io_in_499, // @[:@54599.4]
  input  [3:0] io_in_500, // @[:@54599.4]
  input  [3:0] io_in_501, // @[:@54599.4]
  input  [3:0] io_in_502, // @[:@54599.4]
  input  [3:0] io_in_503, // @[:@54599.4]
  input  [3:0] io_in_504, // @[:@54599.4]
  input  [3:0] io_in_505, // @[:@54599.4]
  input  [3:0] io_in_506, // @[:@54599.4]
  input  [3:0] io_in_507, // @[:@54599.4]
  input  [3:0] io_in_508, // @[:@54599.4]
  input  [3:0] io_in_509, // @[:@54599.4]
  input  [3:0] io_in_510, // @[:@54599.4]
  input  [3:0] io_in_511, // @[:@54599.4]
  input  [3:0] io_in_512, // @[:@54599.4]
  input  [3:0] io_in_513, // @[:@54599.4]
  input  [3:0] io_in_514, // @[:@54599.4]
  input  [3:0] io_in_515, // @[:@54599.4]
  input  [3:0] io_in_516, // @[:@54599.4]
  input  [3:0] io_in_517, // @[:@54599.4]
  input  [3:0] io_in_518, // @[:@54599.4]
  input  [3:0] io_in_519, // @[:@54599.4]
  input  [3:0] io_in_520, // @[:@54599.4]
  input  [3:0] io_in_521, // @[:@54599.4]
  input  [3:0] io_in_522, // @[:@54599.4]
  input  [3:0] io_in_523, // @[:@54599.4]
  input  [3:0] io_in_524, // @[:@54599.4]
  input  [3:0] io_in_525, // @[:@54599.4]
  input  [3:0] io_in_526, // @[:@54599.4]
  input  [3:0] io_in_527, // @[:@54599.4]
  input  [3:0] io_in_528, // @[:@54599.4]
  input  [3:0] io_in_529, // @[:@54599.4]
  input  [3:0] io_in_530, // @[:@54599.4]
  input  [3:0] io_in_531, // @[:@54599.4]
  input  [3:0] io_in_532, // @[:@54599.4]
  input  [3:0] io_in_533, // @[:@54599.4]
  input  [3:0] io_in_534, // @[:@54599.4]
  input  [3:0] io_in_535, // @[:@54599.4]
  input  [3:0] io_in_536, // @[:@54599.4]
  input  [3:0] io_in_537, // @[:@54599.4]
  input  [3:0] io_in_538, // @[:@54599.4]
  input  [3:0] io_in_539, // @[:@54599.4]
  input  [3:0] io_in_540, // @[:@54599.4]
  input  [3:0] io_in_541, // @[:@54599.4]
  input  [3:0] io_in_542, // @[:@54599.4]
  input  [3:0] io_in_543, // @[:@54599.4]
  input  [3:0] io_in_544, // @[:@54599.4]
  input  [3:0] io_in_545, // @[:@54599.4]
  input  [3:0] io_in_546, // @[:@54599.4]
  input  [3:0] io_in_547, // @[:@54599.4]
  input  [3:0] io_in_548, // @[:@54599.4]
  input  [3:0] io_in_549, // @[:@54599.4]
  input  [3:0] io_in_550, // @[:@54599.4]
  input  [3:0] io_in_551, // @[:@54599.4]
  input  [3:0] io_in_552, // @[:@54599.4]
  input  [3:0] io_in_553, // @[:@54599.4]
  input  [3:0] io_in_554, // @[:@54599.4]
  input  [3:0] io_in_555, // @[:@54599.4]
  input  [3:0] io_in_556, // @[:@54599.4]
  input  [3:0] io_in_557, // @[:@54599.4]
  input  [3:0] io_in_558, // @[:@54599.4]
  input  [3:0] io_in_559, // @[:@54599.4]
  input  [3:0] io_in_560, // @[:@54599.4]
  input  [3:0] io_in_561, // @[:@54599.4]
  input  [3:0] io_in_562, // @[:@54599.4]
  input  [3:0] io_in_563, // @[:@54599.4]
  input  [3:0] io_in_564, // @[:@54599.4]
  input  [3:0] io_in_565, // @[:@54599.4]
  input  [3:0] io_in_566, // @[:@54599.4]
  input  [3:0] io_in_567, // @[:@54599.4]
  input  [3:0] io_in_568, // @[:@54599.4]
  input  [3:0] io_in_569, // @[:@54599.4]
  input  [3:0] io_in_570, // @[:@54599.4]
  input  [3:0] io_in_571, // @[:@54599.4]
  input  [3:0] io_in_572, // @[:@54599.4]
  input  [3:0] io_in_573, // @[:@54599.4]
  input  [3:0] io_in_574, // @[:@54599.4]
  input  [3:0] io_in_575, // @[:@54599.4]
  input  [3:0] io_in_576, // @[:@54599.4]
  input  [3:0] io_in_577, // @[:@54599.4]
  input  [3:0] io_in_578, // @[:@54599.4]
  input  [3:0] io_in_579, // @[:@54599.4]
  input  [3:0] io_in_580, // @[:@54599.4]
  input  [3:0] io_in_581, // @[:@54599.4]
  input  [3:0] io_in_582, // @[:@54599.4]
  input  [3:0] io_in_583, // @[:@54599.4]
  input  [3:0] io_in_584, // @[:@54599.4]
  input  [3:0] io_in_585, // @[:@54599.4]
  input  [3:0] io_in_586, // @[:@54599.4]
  input  [3:0] io_in_587, // @[:@54599.4]
  input  [3:0] io_in_588, // @[:@54599.4]
  input  [3:0] io_in_589, // @[:@54599.4]
  input  [3:0] io_in_590, // @[:@54599.4]
  input  [3:0] io_in_591, // @[:@54599.4]
  input  [3:0] io_in_592, // @[:@54599.4]
  input  [3:0] io_in_593, // @[:@54599.4]
  input  [3:0] io_in_594, // @[:@54599.4]
  input  [3:0] io_in_595, // @[:@54599.4]
  input  [3:0] io_in_596, // @[:@54599.4]
  input  [3:0] io_in_597, // @[:@54599.4]
  input  [3:0] io_in_598, // @[:@54599.4]
  input  [3:0] io_in_599, // @[:@54599.4]
  input  [3:0] io_in_600, // @[:@54599.4]
  input  [3:0] io_in_601, // @[:@54599.4]
  input  [3:0] io_in_602, // @[:@54599.4]
  input  [3:0] io_in_603, // @[:@54599.4]
  input  [3:0] io_in_604, // @[:@54599.4]
  input  [3:0] io_in_605, // @[:@54599.4]
  input  [3:0] io_in_606, // @[:@54599.4]
  input  [3:0] io_in_607, // @[:@54599.4]
  input  [3:0] io_in_608, // @[:@54599.4]
  input  [3:0] io_in_609, // @[:@54599.4]
  input  [3:0] io_in_610, // @[:@54599.4]
  input  [3:0] io_in_611, // @[:@54599.4]
  input  [3:0] io_in_612, // @[:@54599.4]
  input  [3:0] io_in_613, // @[:@54599.4]
  input  [3:0] io_in_614, // @[:@54599.4]
  input  [3:0] io_in_615, // @[:@54599.4]
  input  [3:0] io_in_616, // @[:@54599.4]
  input  [3:0] io_in_617, // @[:@54599.4]
  input  [3:0] io_in_618, // @[:@54599.4]
  input  [3:0] io_in_619, // @[:@54599.4]
  input  [3:0] io_in_620, // @[:@54599.4]
  input  [3:0] io_in_621, // @[:@54599.4]
  input  [3:0] io_in_622, // @[:@54599.4]
  input  [3:0] io_in_623, // @[:@54599.4]
  input  [3:0] io_in_624, // @[:@54599.4]
  input  [3:0] io_in_625, // @[:@54599.4]
  input  [3:0] io_in_626, // @[:@54599.4]
  input  [3:0] io_in_627, // @[:@54599.4]
  input  [3:0] io_in_628, // @[:@54599.4]
  input  [3:0] io_in_629, // @[:@54599.4]
  input  [3:0] io_in_630, // @[:@54599.4]
  input  [3:0] io_in_631, // @[:@54599.4]
  input  [3:0] io_in_632, // @[:@54599.4]
  input  [3:0] io_in_633, // @[:@54599.4]
  input  [3:0] io_in_634, // @[:@54599.4]
  input  [3:0] io_in_635, // @[:@54599.4]
  input  [3:0] io_in_636, // @[:@54599.4]
  input  [3:0] io_in_637, // @[:@54599.4]
  input  [3:0] io_in_638, // @[:@54599.4]
  input  [3:0] io_in_639, // @[:@54599.4]
  input  [3:0] io_in_640, // @[:@54599.4]
  input  [3:0] io_in_641, // @[:@54599.4]
  input  [3:0] io_in_642, // @[:@54599.4]
  input  [3:0] io_in_643, // @[:@54599.4]
  input  [3:0] io_in_644, // @[:@54599.4]
  input  [3:0] io_in_645, // @[:@54599.4]
  input  [3:0] io_in_646, // @[:@54599.4]
  input  [3:0] io_in_647, // @[:@54599.4]
  input  [3:0] io_in_648, // @[:@54599.4]
  input  [3:0] io_in_649, // @[:@54599.4]
  input  [3:0] io_in_650, // @[:@54599.4]
  input  [3:0] io_in_651, // @[:@54599.4]
  input  [3:0] io_in_652, // @[:@54599.4]
  input  [3:0] io_in_653, // @[:@54599.4]
  input  [3:0] io_in_654, // @[:@54599.4]
  input  [3:0] io_in_655, // @[:@54599.4]
  input  [3:0] io_in_656, // @[:@54599.4]
  input  [3:0] io_in_657, // @[:@54599.4]
  input  [3:0] io_in_658, // @[:@54599.4]
  input  [3:0] io_in_659, // @[:@54599.4]
  input  [3:0] io_in_660, // @[:@54599.4]
  input  [3:0] io_in_661, // @[:@54599.4]
  input  [3:0] io_in_662, // @[:@54599.4]
  input  [3:0] io_in_663, // @[:@54599.4]
  input  [3:0] io_in_664, // @[:@54599.4]
  input  [3:0] io_in_665, // @[:@54599.4]
  input  [3:0] io_in_666, // @[:@54599.4]
  input  [3:0] io_in_667, // @[:@54599.4]
  input  [3:0] io_in_668, // @[:@54599.4]
  input  [3:0] io_in_669, // @[:@54599.4]
  input  [3:0] io_in_670, // @[:@54599.4]
  input  [3:0] io_in_671, // @[:@54599.4]
  input  [3:0] io_in_672, // @[:@54599.4]
  input  [3:0] io_in_673, // @[:@54599.4]
  input  [3:0] io_in_674, // @[:@54599.4]
  input  [3:0] io_in_675, // @[:@54599.4]
  input  [3:0] io_in_676, // @[:@54599.4]
  input  [3:0] io_in_677, // @[:@54599.4]
  input  [3:0] io_in_678, // @[:@54599.4]
  input  [3:0] io_in_679, // @[:@54599.4]
  input  [3:0] io_in_680, // @[:@54599.4]
  input  [3:0] io_in_681, // @[:@54599.4]
  input  [3:0] io_in_682, // @[:@54599.4]
  input  [3:0] io_in_683, // @[:@54599.4]
  input  [3:0] io_in_684, // @[:@54599.4]
  input  [3:0] io_in_685, // @[:@54599.4]
  input  [3:0] io_in_686, // @[:@54599.4]
  input  [3:0] io_in_687, // @[:@54599.4]
  input  [3:0] io_in_688, // @[:@54599.4]
  input  [3:0] io_in_689, // @[:@54599.4]
  input  [3:0] io_in_690, // @[:@54599.4]
  input  [3:0] io_in_691, // @[:@54599.4]
  input  [3:0] io_in_692, // @[:@54599.4]
  input  [3:0] io_in_693, // @[:@54599.4]
  input  [3:0] io_in_694, // @[:@54599.4]
  input  [3:0] io_in_695, // @[:@54599.4]
  input  [3:0] io_in_696, // @[:@54599.4]
  input  [3:0] io_in_697, // @[:@54599.4]
  input  [3:0] io_in_698, // @[:@54599.4]
  input  [3:0] io_in_699, // @[:@54599.4]
  input  [3:0] io_in_700, // @[:@54599.4]
  input  [3:0] io_in_701, // @[:@54599.4]
  input  [3:0] io_in_702, // @[:@54599.4]
  input  [3:0] io_in_703, // @[:@54599.4]
  input  [3:0] io_in_704, // @[:@54599.4]
  input  [3:0] io_in_705, // @[:@54599.4]
  input  [3:0] io_in_706, // @[:@54599.4]
  input  [3:0] io_in_707, // @[:@54599.4]
  input  [3:0] io_in_708, // @[:@54599.4]
  input  [3:0] io_in_709, // @[:@54599.4]
  input  [3:0] io_in_710, // @[:@54599.4]
  input  [3:0] io_in_711, // @[:@54599.4]
  input  [3:0] io_in_712, // @[:@54599.4]
  input  [3:0] io_in_713, // @[:@54599.4]
  input  [3:0] io_in_714, // @[:@54599.4]
  input  [3:0] io_in_715, // @[:@54599.4]
  input  [3:0] io_in_716, // @[:@54599.4]
  input  [3:0] io_in_717, // @[:@54599.4]
  input  [3:0] io_in_718, // @[:@54599.4]
  input  [3:0] io_in_719, // @[:@54599.4]
  input  [3:0] io_in_720, // @[:@54599.4]
  input  [3:0] io_in_721, // @[:@54599.4]
  input  [3:0] io_in_722, // @[:@54599.4]
  input  [3:0] io_in_723, // @[:@54599.4]
  input  [3:0] io_in_724, // @[:@54599.4]
  input  [3:0] io_in_725, // @[:@54599.4]
  input  [3:0] io_in_726, // @[:@54599.4]
  input  [3:0] io_in_727, // @[:@54599.4]
  input  [3:0] io_in_728, // @[:@54599.4]
  input  [3:0] io_in_729, // @[:@54599.4]
  input  [3:0] io_in_730, // @[:@54599.4]
  input  [3:0] io_in_731, // @[:@54599.4]
  input  [3:0] io_in_732, // @[:@54599.4]
  input  [3:0] io_in_733, // @[:@54599.4]
  input  [3:0] io_in_734, // @[:@54599.4]
  input  [3:0] io_in_735, // @[:@54599.4]
  input  [3:0] io_in_736, // @[:@54599.4]
  input  [3:0] io_in_737, // @[:@54599.4]
  input  [3:0] io_in_738, // @[:@54599.4]
  input  [3:0] io_in_739, // @[:@54599.4]
  input  [3:0] io_in_740, // @[:@54599.4]
  input  [3:0] io_in_741, // @[:@54599.4]
  input  [3:0] io_in_742, // @[:@54599.4]
  input  [3:0] io_in_743, // @[:@54599.4]
  input  [3:0] io_in_744, // @[:@54599.4]
  input  [3:0] io_in_745, // @[:@54599.4]
  input  [3:0] io_in_746, // @[:@54599.4]
  input  [3:0] io_in_747, // @[:@54599.4]
  input  [3:0] io_in_748, // @[:@54599.4]
  input  [3:0] io_in_749, // @[:@54599.4]
  input  [3:0] io_in_750, // @[:@54599.4]
  input  [3:0] io_in_751, // @[:@54599.4]
  input  [3:0] io_in_752, // @[:@54599.4]
  input  [3:0] io_in_753, // @[:@54599.4]
  input  [3:0] io_in_754, // @[:@54599.4]
  input  [3:0] io_in_755, // @[:@54599.4]
  input  [3:0] io_in_756, // @[:@54599.4]
  input  [3:0] io_in_757, // @[:@54599.4]
  input  [3:0] io_in_758, // @[:@54599.4]
  input  [3:0] io_in_759, // @[:@54599.4]
  input  [3:0] io_in_760, // @[:@54599.4]
  input  [3:0] io_in_761, // @[:@54599.4]
  input  [3:0] io_in_762, // @[:@54599.4]
  input  [3:0] io_in_763, // @[:@54599.4]
  input  [3:0] io_in_764, // @[:@54599.4]
  input  [3:0] io_in_765, // @[:@54599.4]
  input  [3:0] io_in_766, // @[:@54599.4]
  input  [3:0] io_in_767, // @[:@54599.4]
  input  [3:0] io_in_768, // @[:@54599.4]
  input  [3:0] io_in_769, // @[:@54599.4]
  input  [3:0] io_in_770, // @[:@54599.4]
  input  [3:0] io_in_771, // @[:@54599.4]
  input  [3:0] io_in_772, // @[:@54599.4]
  input  [3:0] io_in_773, // @[:@54599.4]
  input  [3:0] io_in_774, // @[:@54599.4]
  input  [3:0] io_in_775, // @[:@54599.4]
  input  [3:0] io_in_776, // @[:@54599.4]
  input  [3:0] io_in_777, // @[:@54599.4]
  input  [3:0] io_in_778, // @[:@54599.4]
  input  [3:0] io_in_779, // @[:@54599.4]
  input  [3:0] io_in_780, // @[:@54599.4]
  input  [3:0] io_in_781, // @[:@54599.4]
  input  [3:0] io_in_782, // @[:@54599.4]
  input  [3:0] io_in_783, // @[:@54599.4]
  output [9:0] io_out_0, // @[:@54599.4]
  output [9:0] io_out_1, // @[:@54599.4]
  output [9:0] io_out_2, // @[:@54599.4]
  output [9:0] io_out_3, // @[:@54599.4]
  output [9:0] io_out_4, // @[:@54599.4]
  output [9:0] io_out_5, // @[:@54599.4]
  output [9:0] io_out_6, // @[:@54599.4]
  output [9:0] io_out_7, // @[:@54599.4]
  output [9:0] io_out_8, // @[:@54599.4]
  output [9:0] io_out_9 // @[:@54599.4]
);
  wire [3:0] fc1_io_in_0; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_3; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_5; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_10; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_12; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_13; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_14; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_15; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_19; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_21; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_23; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_25; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_28; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_29; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_30; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_32; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_33; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_34; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_35; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_36; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_37; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_38; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_39; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_40; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_41; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_42; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_43; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_44; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_45; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_46; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_47; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_48; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_49; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_50; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_51; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_52; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_54; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_56; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_59; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_60; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_61; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_62; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_63; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_64; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_65; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_66; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_67; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_68; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_69; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_70; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_71; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_72; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_73; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_74; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_75; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_76; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_77; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_78; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_79; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_80; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_81; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_82; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_83; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_86; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_87; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_88; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_89; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_90; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_91; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_92; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_93; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_94; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_95; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_96; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_97; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_98; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_99; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_100; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_101; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_102; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_103; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_104; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_105; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_106; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_107; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_108; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_109; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_110; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_113; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_114; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_115; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_116; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_117; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_118; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_119; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_120; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_121; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_122; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_123; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_124; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_125; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_126; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_127; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_128; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_129; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_130; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_131; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_132; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_133; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_134; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_135; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_136; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_137; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_138; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_139; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_140; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_142; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_143; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_144; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_145; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_146; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_147; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_148; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_149; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_150; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_151; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_152; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_153; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_154; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_155; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_156; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_157; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_158; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_159; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_160; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_161; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_162; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_163; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_164; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_165; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_166; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_167; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_168; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_169; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_170; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_171; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_172; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_173; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_174; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_175; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_176; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_177; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_178; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_179; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_180; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_181; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_182; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_183; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_184; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_185; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_186; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_187; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_188; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_189; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_190; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_191; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_192; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_193; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_194; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_195; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_196; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_197; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_198; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_199; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_200; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_201; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_202; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_203; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_204; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_205; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_206; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_207; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_208; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_209; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_210; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_211; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_212; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_213; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_214; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_215; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_216; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_217; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_218; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_219; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_220; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_221; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_222; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_223; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_224; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_225; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_226; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_227; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_228; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_229; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_230; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_231; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_232; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_233; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_234; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_235; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_236; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_237; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_238; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_239; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_240; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_241; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_242; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_243; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_244; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_245; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_246; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_247; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_248; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_249; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_250; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_251; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_252; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_253; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_254; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_255; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_256; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_257; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_258; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_259; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_260; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_261; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_262; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_263; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_264; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_265; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_266; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_267; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_268; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_269; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_270; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_271; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_272; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_273; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_274; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_275; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_276; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_277; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_278; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_279; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_280; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_281; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_282; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_283; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_284; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_285; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_286; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_287; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_288; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_289; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_290; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_291; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_292; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_293; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_294; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_295; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_296; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_297; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_298; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_299; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_300; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_301; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_302; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_303; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_304; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_305; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_306; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_307; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_308; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_309; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_310; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_311; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_312; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_313; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_314; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_315; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_316; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_317; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_318; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_319; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_320; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_321; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_322; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_323; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_324; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_325; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_326; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_327; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_328; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_329; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_330; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_331; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_332; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_333; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_334; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_335; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_336; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_337; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_338; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_339; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_340; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_341; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_342; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_343; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_344; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_345; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_346; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_347; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_348; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_349; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_350; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_351; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_352; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_353; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_354; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_355; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_356; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_357; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_358; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_359; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_360; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_361; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_362; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_363; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_364; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_365; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_366; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_367; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_368; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_369; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_370; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_371; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_372; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_373; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_374; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_375; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_376; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_377; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_378; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_379; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_380; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_381; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_382; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_383; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_384; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_385; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_386; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_387; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_388; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_389; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_390; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_391; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_392; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_393; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_394; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_395; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_396; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_397; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_398; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_399; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_400; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_401; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_402; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_403; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_404; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_405; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_406; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_407; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_408; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_409; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_410; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_411; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_412; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_413; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_414; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_415; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_416; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_417; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_418; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_419; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_420; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_421; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_422; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_423; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_424; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_425; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_426; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_427; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_428; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_429; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_430; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_431; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_432; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_433; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_434; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_435; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_436; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_437; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_438; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_439; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_440; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_441; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_442; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_443; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_444; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_445; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_446; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_447; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_448; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_449; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_450; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_451; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_452; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_453; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_454; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_455; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_456; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_457; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_458; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_459; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_460; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_461; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_462; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_463; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_464; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_465; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_466; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_467; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_468; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_469; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_470; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_471; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_472; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_473; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_474; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_475; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_476; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_477; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_478; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_479; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_480; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_481; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_482; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_483; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_484; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_485; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_486; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_487; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_488; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_489; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_490; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_491; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_492; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_493; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_494; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_495; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_496; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_497; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_498; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_499; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_500; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_501; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_502; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_503; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_504; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_505; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_506; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_507; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_508; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_509; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_510; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_511; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_512; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_513; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_514; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_515; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_516; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_517; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_518; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_519; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_520; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_521; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_522; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_523; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_524; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_525; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_526; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_527; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_528; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_529; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_530; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_531; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_532; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_533; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_534; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_535; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_536; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_537; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_538; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_539; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_540; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_541; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_542; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_543; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_544; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_545; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_546; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_547; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_548; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_549; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_550; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_551; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_552; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_553; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_554; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_555; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_556; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_557; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_558; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_559; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_561; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_562; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_563; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_564; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_565; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_566; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_567; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_568; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_569; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_570; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_571; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_572; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_573; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_574; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_575; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_576; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_577; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_578; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_579; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_580; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_581; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_582; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_583; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_584; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_585; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_586; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_587; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_588; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_589; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_590; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_591; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_592; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_593; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_594; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_595; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_596; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_597; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_598; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_599; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_600; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_601; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_602; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_603; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_604; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_605; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_606; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_607; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_608; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_609; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_610; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_611; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_612; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_613; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_614; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_615; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_616; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_617; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_618; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_619; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_620; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_621; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_622; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_623; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_624; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_625; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_626; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_627; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_628; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_629; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_630; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_631; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_632; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_633; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_634; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_635; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_636; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_637; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_638; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_639; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_640; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_641; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_642; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_646; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_647; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_648; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_649; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_650; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_651; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_652; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_653; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_654; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_655; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_656; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_657; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_658; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_659; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_660; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_661; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_662; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_663; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_664; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_665; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_666; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_667; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_668; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_669; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_670; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_673; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_674; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_675; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_676; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_677; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_678; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_679; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_680; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_681; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_682; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_683; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_684; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_685; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_686; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_687; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_688; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_689; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_690; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_691; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_692; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_693; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_694; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_695; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_696; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_697; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_698; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_699; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_702; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_703; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_704; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_705; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_706; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_707; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_708; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_709; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_710; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_711; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_712; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_713; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_714; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_715; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_716; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_717; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_718; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_719; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_720; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_721; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_722; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_723; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_724; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_725; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_726; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_728; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_729; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_731; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_732; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_733; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_734; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_735; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_736; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_737; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_738; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_739; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_740; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_741; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_742; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_743; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_744; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_745; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_746; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_747; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_748; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_749; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_750; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_751; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_752; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_753; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_756; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_758; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_760; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_761; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_762; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_763; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_764; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_765; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_766; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_767; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_768; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_769; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_770; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_771; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_772; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_773; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_774; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_775; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_776; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_777; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_778; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_779; // @[Models.scala 13:15:@54601.4]
  wire [3:0] fc1_io_in_780; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_0; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_1; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_2; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_3; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_4; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_5; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_6; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_7; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_8; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_9; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_10; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_11; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_12; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_13; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_14; // @[Models.scala 13:15:@54601.4]
  wire [13:0] fc1_io_out_15; // @[Models.scala 13:15:@54601.4]
  wire [13:0] bn_bi1_io_in_0; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_1; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_2; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_3; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_4; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_5; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_6; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_7; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_8; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_9; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_10; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_11; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_12; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_13; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_14; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_in_15; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_0; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_1; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_2; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_3; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_4; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_5; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_6; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_7; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_8; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_9; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_10; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_11; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_12; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_13; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_14; // @[Models.scala 22:24:@54610.4]
  wire [13:0] bn_bi1_io_out_15; // @[Models.scala 22:24:@54610.4]
  wire [1:0] fc2_io_in_0; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_1; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_2; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_3; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_4; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_5; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_6; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_7; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_8; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_9; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_10; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_11; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_12; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_13; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_14; // @[Models.scala 26:15:@54613.4]
  wire [1:0] fc2_io_in_15; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_0; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_1; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_2; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_3; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_4; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_5; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_6; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_7; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_8; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_9; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_10; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_11; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_12; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_13; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_14; // @[Models.scala 26:15:@54613.4]
  wire [5:0] fc2_io_out_15; // @[Models.scala 26:15:@54613.4]
  wire [5:0] bn_bi2_io_in_0; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_1; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_2; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_3; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_4; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_5; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_6; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_7; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_8; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_9; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_10; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_11; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_12; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_13; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_14; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_in_15; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_0; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_1; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_2; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_3; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_4; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_5; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_6; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_7; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_8; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_9; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_10; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_11; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_12; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_13; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_14; // @[Models.scala 35:24:@54622.4]
  wire [5:0] bn_bi2_io_out_15; // @[Models.scala 35:24:@54622.4]
  wire [1:0] fc3_io_in_0; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_1; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_2; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_3; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_4; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_5; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_6; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_7; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_8; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_9; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_10; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_11; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_12; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_13; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_14; // @[Models.scala 39:15:@54625.4]
  wire [1:0] fc3_io_in_15; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_0; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_1; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_2; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_3; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_4; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_5; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_6; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_7; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_8; // @[Models.scala 39:15:@54625.4]
  wire [5:0] fc3_io_out_9; // @[Models.scala 39:15:@54625.4]
  wire [5:0] bn3_io_in_0; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_1; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_2; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_3; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_4; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_5; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_6; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_7; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_8; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_in_9; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_0; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_1; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_2; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_3; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_4; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_5; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_6; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_7; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_8; // @[Models.scala 45:21:@54628.4]
  wire [5:0] bn3_io_out_9; // @[Models.scala 45:21:@54628.4]
  wire [1:0] _GEN_0;
  wire [1:0] _GEN_1;
  wire [1:0] _GEN_2;
  wire [1:0] _GEN_3;
  wire [1:0] _GEN_4;
  wire [1:0] _GEN_5;
  wire [1:0] _GEN_6;
  wire [1:0] _GEN_7;
  wire [1:0] _GEN_8;
  wire [1:0] _GEN_9;
  wire [1:0] _GEN_10;
  wire [1:0] _GEN_11;
  wire [1:0] _GEN_12;
  wire [1:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [1:0] _GEN_16;
  wire [1:0] _GEN_17;
  wire [1:0] _GEN_18;
  wire [1:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [1:0] _GEN_22;
  wire [1:0] _GEN_23;
  wire [1:0] _GEN_24;
  wire [1:0] _GEN_25;
  wire [1:0] _GEN_26;
  wire [1:0] _GEN_27;
  wire [1:0] _GEN_28;
  wire [1:0] _GEN_29;
  wire [1:0] _GEN_30;
  wire [1:0] _GEN_31;
  Linear_p fc1 ( // @[Models.scala 13:15:@54601.4]
    .io_in_0(fc1_io_in_0),
    .io_in_3(fc1_io_in_3),
    .io_in_5(fc1_io_in_5),
    .io_in_10(fc1_io_in_10),
    .io_in_12(fc1_io_in_12),
    .io_in_13(fc1_io_in_13),
    .io_in_14(fc1_io_in_14),
    .io_in_15(fc1_io_in_15),
    .io_in_19(fc1_io_in_19),
    .io_in_21(fc1_io_in_21),
    .io_in_23(fc1_io_in_23),
    .io_in_25(fc1_io_in_25),
    .io_in_28(fc1_io_in_28),
    .io_in_29(fc1_io_in_29),
    .io_in_30(fc1_io_in_30),
    .io_in_32(fc1_io_in_32),
    .io_in_33(fc1_io_in_33),
    .io_in_34(fc1_io_in_34),
    .io_in_35(fc1_io_in_35),
    .io_in_36(fc1_io_in_36),
    .io_in_37(fc1_io_in_37),
    .io_in_38(fc1_io_in_38),
    .io_in_39(fc1_io_in_39),
    .io_in_40(fc1_io_in_40),
    .io_in_41(fc1_io_in_41),
    .io_in_42(fc1_io_in_42),
    .io_in_43(fc1_io_in_43),
    .io_in_44(fc1_io_in_44),
    .io_in_45(fc1_io_in_45),
    .io_in_46(fc1_io_in_46),
    .io_in_47(fc1_io_in_47),
    .io_in_48(fc1_io_in_48),
    .io_in_49(fc1_io_in_49),
    .io_in_50(fc1_io_in_50),
    .io_in_51(fc1_io_in_51),
    .io_in_52(fc1_io_in_52),
    .io_in_54(fc1_io_in_54),
    .io_in_56(fc1_io_in_56),
    .io_in_59(fc1_io_in_59),
    .io_in_60(fc1_io_in_60),
    .io_in_61(fc1_io_in_61),
    .io_in_62(fc1_io_in_62),
    .io_in_63(fc1_io_in_63),
    .io_in_64(fc1_io_in_64),
    .io_in_65(fc1_io_in_65),
    .io_in_66(fc1_io_in_66),
    .io_in_67(fc1_io_in_67),
    .io_in_68(fc1_io_in_68),
    .io_in_69(fc1_io_in_69),
    .io_in_70(fc1_io_in_70),
    .io_in_71(fc1_io_in_71),
    .io_in_72(fc1_io_in_72),
    .io_in_73(fc1_io_in_73),
    .io_in_74(fc1_io_in_74),
    .io_in_75(fc1_io_in_75),
    .io_in_76(fc1_io_in_76),
    .io_in_77(fc1_io_in_77),
    .io_in_78(fc1_io_in_78),
    .io_in_79(fc1_io_in_79),
    .io_in_80(fc1_io_in_80),
    .io_in_81(fc1_io_in_81),
    .io_in_82(fc1_io_in_82),
    .io_in_83(fc1_io_in_83),
    .io_in_86(fc1_io_in_86),
    .io_in_87(fc1_io_in_87),
    .io_in_88(fc1_io_in_88),
    .io_in_89(fc1_io_in_89),
    .io_in_90(fc1_io_in_90),
    .io_in_91(fc1_io_in_91),
    .io_in_92(fc1_io_in_92),
    .io_in_93(fc1_io_in_93),
    .io_in_94(fc1_io_in_94),
    .io_in_95(fc1_io_in_95),
    .io_in_96(fc1_io_in_96),
    .io_in_97(fc1_io_in_97),
    .io_in_98(fc1_io_in_98),
    .io_in_99(fc1_io_in_99),
    .io_in_100(fc1_io_in_100),
    .io_in_101(fc1_io_in_101),
    .io_in_102(fc1_io_in_102),
    .io_in_103(fc1_io_in_103),
    .io_in_104(fc1_io_in_104),
    .io_in_105(fc1_io_in_105),
    .io_in_106(fc1_io_in_106),
    .io_in_107(fc1_io_in_107),
    .io_in_108(fc1_io_in_108),
    .io_in_109(fc1_io_in_109),
    .io_in_110(fc1_io_in_110),
    .io_in_113(fc1_io_in_113),
    .io_in_114(fc1_io_in_114),
    .io_in_115(fc1_io_in_115),
    .io_in_116(fc1_io_in_116),
    .io_in_117(fc1_io_in_117),
    .io_in_118(fc1_io_in_118),
    .io_in_119(fc1_io_in_119),
    .io_in_120(fc1_io_in_120),
    .io_in_121(fc1_io_in_121),
    .io_in_122(fc1_io_in_122),
    .io_in_123(fc1_io_in_123),
    .io_in_124(fc1_io_in_124),
    .io_in_125(fc1_io_in_125),
    .io_in_126(fc1_io_in_126),
    .io_in_127(fc1_io_in_127),
    .io_in_128(fc1_io_in_128),
    .io_in_129(fc1_io_in_129),
    .io_in_130(fc1_io_in_130),
    .io_in_131(fc1_io_in_131),
    .io_in_132(fc1_io_in_132),
    .io_in_133(fc1_io_in_133),
    .io_in_134(fc1_io_in_134),
    .io_in_135(fc1_io_in_135),
    .io_in_136(fc1_io_in_136),
    .io_in_137(fc1_io_in_137),
    .io_in_138(fc1_io_in_138),
    .io_in_139(fc1_io_in_139),
    .io_in_140(fc1_io_in_140),
    .io_in_142(fc1_io_in_142),
    .io_in_143(fc1_io_in_143),
    .io_in_144(fc1_io_in_144),
    .io_in_145(fc1_io_in_145),
    .io_in_146(fc1_io_in_146),
    .io_in_147(fc1_io_in_147),
    .io_in_148(fc1_io_in_148),
    .io_in_149(fc1_io_in_149),
    .io_in_150(fc1_io_in_150),
    .io_in_151(fc1_io_in_151),
    .io_in_152(fc1_io_in_152),
    .io_in_153(fc1_io_in_153),
    .io_in_154(fc1_io_in_154),
    .io_in_155(fc1_io_in_155),
    .io_in_156(fc1_io_in_156),
    .io_in_157(fc1_io_in_157),
    .io_in_158(fc1_io_in_158),
    .io_in_159(fc1_io_in_159),
    .io_in_160(fc1_io_in_160),
    .io_in_161(fc1_io_in_161),
    .io_in_162(fc1_io_in_162),
    .io_in_163(fc1_io_in_163),
    .io_in_164(fc1_io_in_164),
    .io_in_165(fc1_io_in_165),
    .io_in_166(fc1_io_in_166),
    .io_in_167(fc1_io_in_167),
    .io_in_168(fc1_io_in_168),
    .io_in_169(fc1_io_in_169),
    .io_in_170(fc1_io_in_170),
    .io_in_171(fc1_io_in_171),
    .io_in_172(fc1_io_in_172),
    .io_in_173(fc1_io_in_173),
    .io_in_174(fc1_io_in_174),
    .io_in_175(fc1_io_in_175),
    .io_in_176(fc1_io_in_176),
    .io_in_177(fc1_io_in_177),
    .io_in_178(fc1_io_in_178),
    .io_in_179(fc1_io_in_179),
    .io_in_180(fc1_io_in_180),
    .io_in_181(fc1_io_in_181),
    .io_in_182(fc1_io_in_182),
    .io_in_183(fc1_io_in_183),
    .io_in_184(fc1_io_in_184),
    .io_in_185(fc1_io_in_185),
    .io_in_186(fc1_io_in_186),
    .io_in_187(fc1_io_in_187),
    .io_in_188(fc1_io_in_188),
    .io_in_189(fc1_io_in_189),
    .io_in_190(fc1_io_in_190),
    .io_in_191(fc1_io_in_191),
    .io_in_192(fc1_io_in_192),
    .io_in_193(fc1_io_in_193),
    .io_in_194(fc1_io_in_194),
    .io_in_195(fc1_io_in_195),
    .io_in_196(fc1_io_in_196),
    .io_in_197(fc1_io_in_197),
    .io_in_198(fc1_io_in_198),
    .io_in_199(fc1_io_in_199),
    .io_in_200(fc1_io_in_200),
    .io_in_201(fc1_io_in_201),
    .io_in_202(fc1_io_in_202),
    .io_in_203(fc1_io_in_203),
    .io_in_204(fc1_io_in_204),
    .io_in_205(fc1_io_in_205),
    .io_in_206(fc1_io_in_206),
    .io_in_207(fc1_io_in_207),
    .io_in_208(fc1_io_in_208),
    .io_in_209(fc1_io_in_209),
    .io_in_210(fc1_io_in_210),
    .io_in_211(fc1_io_in_211),
    .io_in_212(fc1_io_in_212),
    .io_in_213(fc1_io_in_213),
    .io_in_214(fc1_io_in_214),
    .io_in_215(fc1_io_in_215),
    .io_in_216(fc1_io_in_216),
    .io_in_217(fc1_io_in_217),
    .io_in_218(fc1_io_in_218),
    .io_in_219(fc1_io_in_219),
    .io_in_220(fc1_io_in_220),
    .io_in_221(fc1_io_in_221),
    .io_in_222(fc1_io_in_222),
    .io_in_223(fc1_io_in_223),
    .io_in_224(fc1_io_in_224),
    .io_in_225(fc1_io_in_225),
    .io_in_226(fc1_io_in_226),
    .io_in_227(fc1_io_in_227),
    .io_in_228(fc1_io_in_228),
    .io_in_229(fc1_io_in_229),
    .io_in_230(fc1_io_in_230),
    .io_in_231(fc1_io_in_231),
    .io_in_232(fc1_io_in_232),
    .io_in_233(fc1_io_in_233),
    .io_in_234(fc1_io_in_234),
    .io_in_235(fc1_io_in_235),
    .io_in_236(fc1_io_in_236),
    .io_in_237(fc1_io_in_237),
    .io_in_238(fc1_io_in_238),
    .io_in_239(fc1_io_in_239),
    .io_in_240(fc1_io_in_240),
    .io_in_241(fc1_io_in_241),
    .io_in_242(fc1_io_in_242),
    .io_in_243(fc1_io_in_243),
    .io_in_244(fc1_io_in_244),
    .io_in_245(fc1_io_in_245),
    .io_in_246(fc1_io_in_246),
    .io_in_247(fc1_io_in_247),
    .io_in_248(fc1_io_in_248),
    .io_in_249(fc1_io_in_249),
    .io_in_250(fc1_io_in_250),
    .io_in_251(fc1_io_in_251),
    .io_in_252(fc1_io_in_252),
    .io_in_253(fc1_io_in_253),
    .io_in_254(fc1_io_in_254),
    .io_in_255(fc1_io_in_255),
    .io_in_256(fc1_io_in_256),
    .io_in_257(fc1_io_in_257),
    .io_in_258(fc1_io_in_258),
    .io_in_259(fc1_io_in_259),
    .io_in_260(fc1_io_in_260),
    .io_in_261(fc1_io_in_261),
    .io_in_262(fc1_io_in_262),
    .io_in_263(fc1_io_in_263),
    .io_in_264(fc1_io_in_264),
    .io_in_265(fc1_io_in_265),
    .io_in_266(fc1_io_in_266),
    .io_in_267(fc1_io_in_267),
    .io_in_268(fc1_io_in_268),
    .io_in_269(fc1_io_in_269),
    .io_in_270(fc1_io_in_270),
    .io_in_271(fc1_io_in_271),
    .io_in_272(fc1_io_in_272),
    .io_in_273(fc1_io_in_273),
    .io_in_274(fc1_io_in_274),
    .io_in_275(fc1_io_in_275),
    .io_in_276(fc1_io_in_276),
    .io_in_277(fc1_io_in_277),
    .io_in_278(fc1_io_in_278),
    .io_in_279(fc1_io_in_279),
    .io_in_280(fc1_io_in_280),
    .io_in_281(fc1_io_in_281),
    .io_in_282(fc1_io_in_282),
    .io_in_283(fc1_io_in_283),
    .io_in_284(fc1_io_in_284),
    .io_in_285(fc1_io_in_285),
    .io_in_286(fc1_io_in_286),
    .io_in_287(fc1_io_in_287),
    .io_in_288(fc1_io_in_288),
    .io_in_289(fc1_io_in_289),
    .io_in_290(fc1_io_in_290),
    .io_in_291(fc1_io_in_291),
    .io_in_292(fc1_io_in_292),
    .io_in_293(fc1_io_in_293),
    .io_in_294(fc1_io_in_294),
    .io_in_295(fc1_io_in_295),
    .io_in_296(fc1_io_in_296),
    .io_in_297(fc1_io_in_297),
    .io_in_298(fc1_io_in_298),
    .io_in_299(fc1_io_in_299),
    .io_in_300(fc1_io_in_300),
    .io_in_301(fc1_io_in_301),
    .io_in_302(fc1_io_in_302),
    .io_in_303(fc1_io_in_303),
    .io_in_304(fc1_io_in_304),
    .io_in_305(fc1_io_in_305),
    .io_in_306(fc1_io_in_306),
    .io_in_307(fc1_io_in_307),
    .io_in_308(fc1_io_in_308),
    .io_in_309(fc1_io_in_309),
    .io_in_310(fc1_io_in_310),
    .io_in_311(fc1_io_in_311),
    .io_in_312(fc1_io_in_312),
    .io_in_313(fc1_io_in_313),
    .io_in_314(fc1_io_in_314),
    .io_in_315(fc1_io_in_315),
    .io_in_316(fc1_io_in_316),
    .io_in_317(fc1_io_in_317),
    .io_in_318(fc1_io_in_318),
    .io_in_319(fc1_io_in_319),
    .io_in_320(fc1_io_in_320),
    .io_in_321(fc1_io_in_321),
    .io_in_322(fc1_io_in_322),
    .io_in_323(fc1_io_in_323),
    .io_in_324(fc1_io_in_324),
    .io_in_325(fc1_io_in_325),
    .io_in_326(fc1_io_in_326),
    .io_in_327(fc1_io_in_327),
    .io_in_328(fc1_io_in_328),
    .io_in_329(fc1_io_in_329),
    .io_in_330(fc1_io_in_330),
    .io_in_331(fc1_io_in_331),
    .io_in_332(fc1_io_in_332),
    .io_in_333(fc1_io_in_333),
    .io_in_334(fc1_io_in_334),
    .io_in_335(fc1_io_in_335),
    .io_in_336(fc1_io_in_336),
    .io_in_337(fc1_io_in_337),
    .io_in_338(fc1_io_in_338),
    .io_in_339(fc1_io_in_339),
    .io_in_340(fc1_io_in_340),
    .io_in_341(fc1_io_in_341),
    .io_in_342(fc1_io_in_342),
    .io_in_343(fc1_io_in_343),
    .io_in_344(fc1_io_in_344),
    .io_in_345(fc1_io_in_345),
    .io_in_346(fc1_io_in_346),
    .io_in_347(fc1_io_in_347),
    .io_in_348(fc1_io_in_348),
    .io_in_349(fc1_io_in_349),
    .io_in_350(fc1_io_in_350),
    .io_in_351(fc1_io_in_351),
    .io_in_352(fc1_io_in_352),
    .io_in_353(fc1_io_in_353),
    .io_in_354(fc1_io_in_354),
    .io_in_355(fc1_io_in_355),
    .io_in_356(fc1_io_in_356),
    .io_in_357(fc1_io_in_357),
    .io_in_358(fc1_io_in_358),
    .io_in_359(fc1_io_in_359),
    .io_in_360(fc1_io_in_360),
    .io_in_361(fc1_io_in_361),
    .io_in_362(fc1_io_in_362),
    .io_in_363(fc1_io_in_363),
    .io_in_364(fc1_io_in_364),
    .io_in_365(fc1_io_in_365),
    .io_in_366(fc1_io_in_366),
    .io_in_367(fc1_io_in_367),
    .io_in_368(fc1_io_in_368),
    .io_in_369(fc1_io_in_369),
    .io_in_370(fc1_io_in_370),
    .io_in_371(fc1_io_in_371),
    .io_in_372(fc1_io_in_372),
    .io_in_373(fc1_io_in_373),
    .io_in_374(fc1_io_in_374),
    .io_in_375(fc1_io_in_375),
    .io_in_376(fc1_io_in_376),
    .io_in_377(fc1_io_in_377),
    .io_in_378(fc1_io_in_378),
    .io_in_379(fc1_io_in_379),
    .io_in_380(fc1_io_in_380),
    .io_in_381(fc1_io_in_381),
    .io_in_382(fc1_io_in_382),
    .io_in_383(fc1_io_in_383),
    .io_in_384(fc1_io_in_384),
    .io_in_385(fc1_io_in_385),
    .io_in_386(fc1_io_in_386),
    .io_in_387(fc1_io_in_387),
    .io_in_388(fc1_io_in_388),
    .io_in_389(fc1_io_in_389),
    .io_in_390(fc1_io_in_390),
    .io_in_391(fc1_io_in_391),
    .io_in_392(fc1_io_in_392),
    .io_in_393(fc1_io_in_393),
    .io_in_394(fc1_io_in_394),
    .io_in_395(fc1_io_in_395),
    .io_in_396(fc1_io_in_396),
    .io_in_397(fc1_io_in_397),
    .io_in_398(fc1_io_in_398),
    .io_in_399(fc1_io_in_399),
    .io_in_400(fc1_io_in_400),
    .io_in_401(fc1_io_in_401),
    .io_in_402(fc1_io_in_402),
    .io_in_403(fc1_io_in_403),
    .io_in_404(fc1_io_in_404),
    .io_in_405(fc1_io_in_405),
    .io_in_406(fc1_io_in_406),
    .io_in_407(fc1_io_in_407),
    .io_in_408(fc1_io_in_408),
    .io_in_409(fc1_io_in_409),
    .io_in_410(fc1_io_in_410),
    .io_in_411(fc1_io_in_411),
    .io_in_412(fc1_io_in_412),
    .io_in_413(fc1_io_in_413),
    .io_in_414(fc1_io_in_414),
    .io_in_415(fc1_io_in_415),
    .io_in_416(fc1_io_in_416),
    .io_in_417(fc1_io_in_417),
    .io_in_418(fc1_io_in_418),
    .io_in_419(fc1_io_in_419),
    .io_in_420(fc1_io_in_420),
    .io_in_421(fc1_io_in_421),
    .io_in_422(fc1_io_in_422),
    .io_in_423(fc1_io_in_423),
    .io_in_424(fc1_io_in_424),
    .io_in_425(fc1_io_in_425),
    .io_in_426(fc1_io_in_426),
    .io_in_427(fc1_io_in_427),
    .io_in_428(fc1_io_in_428),
    .io_in_429(fc1_io_in_429),
    .io_in_430(fc1_io_in_430),
    .io_in_431(fc1_io_in_431),
    .io_in_432(fc1_io_in_432),
    .io_in_433(fc1_io_in_433),
    .io_in_434(fc1_io_in_434),
    .io_in_435(fc1_io_in_435),
    .io_in_436(fc1_io_in_436),
    .io_in_437(fc1_io_in_437),
    .io_in_438(fc1_io_in_438),
    .io_in_439(fc1_io_in_439),
    .io_in_440(fc1_io_in_440),
    .io_in_441(fc1_io_in_441),
    .io_in_442(fc1_io_in_442),
    .io_in_443(fc1_io_in_443),
    .io_in_444(fc1_io_in_444),
    .io_in_445(fc1_io_in_445),
    .io_in_446(fc1_io_in_446),
    .io_in_447(fc1_io_in_447),
    .io_in_448(fc1_io_in_448),
    .io_in_449(fc1_io_in_449),
    .io_in_450(fc1_io_in_450),
    .io_in_451(fc1_io_in_451),
    .io_in_452(fc1_io_in_452),
    .io_in_453(fc1_io_in_453),
    .io_in_454(fc1_io_in_454),
    .io_in_455(fc1_io_in_455),
    .io_in_456(fc1_io_in_456),
    .io_in_457(fc1_io_in_457),
    .io_in_458(fc1_io_in_458),
    .io_in_459(fc1_io_in_459),
    .io_in_460(fc1_io_in_460),
    .io_in_461(fc1_io_in_461),
    .io_in_462(fc1_io_in_462),
    .io_in_463(fc1_io_in_463),
    .io_in_464(fc1_io_in_464),
    .io_in_465(fc1_io_in_465),
    .io_in_466(fc1_io_in_466),
    .io_in_467(fc1_io_in_467),
    .io_in_468(fc1_io_in_468),
    .io_in_469(fc1_io_in_469),
    .io_in_470(fc1_io_in_470),
    .io_in_471(fc1_io_in_471),
    .io_in_472(fc1_io_in_472),
    .io_in_473(fc1_io_in_473),
    .io_in_474(fc1_io_in_474),
    .io_in_475(fc1_io_in_475),
    .io_in_476(fc1_io_in_476),
    .io_in_477(fc1_io_in_477),
    .io_in_478(fc1_io_in_478),
    .io_in_479(fc1_io_in_479),
    .io_in_480(fc1_io_in_480),
    .io_in_481(fc1_io_in_481),
    .io_in_482(fc1_io_in_482),
    .io_in_483(fc1_io_in_483),
    .io_in_484(fc1_io_in_484),
    .io_in_485(fc1_io_in_485),
    .io_in_486(fc1_io_in_486),
    .io_in_487(fc1_io_in_487),
    .io_in_488(fc1_io_in_488),
    .io_in_489(fc1_io_in_489),
    .io_in_490(fc1_io_in_490),
    .io_in_491(fc1_io_in_491),
    .io_in_492(fc1_io_in_492),
    .io_in_493(fc1_io_in_493),
    .io_in_494(fc1_io_in_494),
    .io_in_495(fc1_io_in_495),
    .io_in_496(fc1_io_in_496),
    .io_in_497(fc1_io_in_497),
    .io_in_498(fc1_io_in_498),
    .io_in_499(fc1_io_in_499),
    .io_in_500(fc1_io_in_500),
    .io_in_501(fc1_io_in_501),
    .io_in_502(fc1_io_in_502),
    .io_in_503(fc1_io_in_503),
    .io_in_504(fc1_io_in_504),
    .io_in_505(fc1_io_in_505),
    .io_in_506(fc1_io_in_506),
    .io_in_507(fc1_io_in_507),
    .io_in_508(fc1_io_in_508),
    .io_in_509(fc1_io_in_509),
    .io_in_510(fc1_io_in_510),
    .io_in_511(fc1_io_in_511),
    .io_in_512(fc1_io_in_512),
    .io_in_513(fc1_io_in_513),
    .io_in_514(fc1_io_in_514),
    .io_in_515(fc1_io_in_515),
    .io_in_516(fc1_io_in_516),
    .io_in_517(fc1_io_in_517),
    .io_in_518(fc1_io_in_518),
    .io_in_519(fc1_io_in_519),
    .io_in_520(fc1_io_in_520),
    .io_in_521(fc1_io_in_521),
    .io_in_522(fc1_io_in_522),
    .io_in_523(fc1_io_in_523),
    .io_in_524(fc1_io_in_524),
    .io_in_525(fc1_io_in_525),
    .io_in_526(fc1_io_in_526),
    .io_in_527(fc1_io_in_527),
    .io_in_528(fc1_io_in_528),
    .io_in_529(fc1_io_in_529),
    .io_in_530(fc1_io_in_530),
    .io_in_531(fc1_io_in_531),
    .io_in_532(fc1_io_in_532),
    .io_in_533(fc1_io_in_533),
    .io_in_534(fc1_io_in_534),
    .io_in_535(fc1_io_in_535),
    .io_in_536(fc1_io_in_536),
    .io_in_537(fc1_io_in_537),
    .io_in_538(fc1_io_in_538),
    .io_in_539(fc1_io_in_539),
    .io_in_540(fc1_io_in_540),
    .io_in_541(fc1_io_in_541),
    .io_in_542(fc1_io_in_542),
    .io_in_543(fc1_io_in_543),
    .io_in_544(fc1_io_in_544),
    .io_in_545(fc1_io_in_545),
    .io_in_546(fc1_io_in_546),
    .io_in_547(fc1_io_in_547),
    .io_in_548(fc1_io_in_548),
    .io_in_549(fc1_io_in_549),
    .io_in_550(fc1_io_in_550),
    .io_in_551(fc1_io_in_551),
    .io_in_552(fc1_io_in_552),
    .io_in_553(fc1_io_in_553),
    .io_in_554(fc1_io_in_554),
    .io_in_555(fc1_io_in_555),
    .io_in_556(fc1_io_in_556),
    .io_in_557(fc1_io_in_557),
    .io_in_558(fc1_io_in_558),
    .io_in_559(fc1_io_in_559),
    .io_in_561(fc1_io_in_561),
    .io_in_562(fc1_io_in_562),
    .io_in_563(fc1_io_in_563),
    .io_in_564(fc1_io_in_564),
    .io_in_565(fc1_io_in_565),
    .io_in_566(fc1_io_in_566),
    .io_in_567(fc1_io_in_567),
    .io_in_568(fc1_io_in_568),
    .io_in_569(fc1_io_in_569),
    .io_in_570(fc1_io_in_570),
    .io_in_571(fc1_io_in_571),
    .io_in_572(fc1_io_in_572),
    .io_in_573(fc1_io_in_573),
    .io_in_574(fc1_io_in_574),
    .io_in_575(fc1_io_in_575),
    .io_in_576(fc1_io_in_576),
    .io_in_577(fc1_io_in_577),
    .io_in_578(fc1_io_in_578),
    .io_in_579(fc1_io_in_579),
    .io_in_580(fc1_io_in_580),
    .io_in_581(fc1_io_in_581),
    .io_in_582(fc1_io_in_582),
    .io_in_583(fc1_io_in_583),
    .io_in_584(fc1_io_in_584),
    .io_in_585(fc1_io_in_585),
    .io_in_586(fc1_io_in_586),
    .io_in_587(fc1_io_in_587),
    .io_in_588(fc1_io_in_588),
    .io_in_589(fc1_io_in_589),
    .io_in_590(fc1_io_in_590),
    .io_in_591(fc1_io_in_591),
    .io_in_592(fc1_io_in_592),
    .io_in_593(fc1_io_in_593),
    .io_in_594(fc1_io_in_594),
    .io_in_595(fc1_io_in_595),
    .io_in_596(fc1_io_in_596),
    .io_in_597(fc1_io_in_597),
    .io_in_598(fc1_io_in_598),
    .io_in_599(fc1_io_in_599),
    .io_in_600(fc1_io_in_600),
    .io_in_601(fc1_io_in_601),
    .io_in_602(fc1_io_in_602),
    .io_in_603(fc1_io_in_603),
    .io_in_604(fc1_io_in_604),
    .io_in_605(fc1_io_in_605),
    .io_in_606(fc1_io_in_606),
    .io_in_607(fc1_io_in_607),
    .io_in_608(fc1_io_in_608),
    .io_in_609(fc1_io_in_609),
    .io_in_610(fc1_io_in_610),
    .io_in_611(fc1_io_in_611),
    .io_in_612(fc1_io_in_612),
    .io_in_613(fc1_io_in_613),
    .io_in_614(fc1_io_in_614),
    .io_in_615(fc1_io_in_615),
    .io_in_616(fc1_io_in_616),
    .io_in_617(fc1_io_in_617),
    .io_in_618(fc1_io_in_618),
    .io_in_619(fc1_io_in_619),
    .io_in_620(fc1_io_in_620),
    .io_in_621(fc1_io_in_621),
    .io_in_622(fc1_io_in_622),
    .io_in_623(fc1_io_in_623),
    .io_in_624(fc1_io_in_624),
    .io_in_625(fc1_io_in_625),
    .io_in_626(fc1_io_in_626),
    .io_in_627(fc1_io_in_627),
    .io_in_628(fc1_io_in_628),
    .io_in_629(fc1_io_in_629),
    .io_in_630(fc1_io_in_630),
    .io_in_631(fc1_io_in_631),
    .io_in_632(fc1_io_in_632),
    .io_in_633(fc1_io_in_633),
    .io_in_634(fc1_io_in_634),
    .io_in_635(fc1_io_in_635),
    .io_in_636(fc1_io_in_636),
    .io_in_637(fc1_io_in_637),
    .io_in_638(fc1_io_in_638),
    .io_in_639(fc1_io_in_639),
    .io_in_640(fc1_io_in_640),
    .io_in_641(fc1_io_in_641),
    .io_in_642(fc1_io_in_642),
    .io_in_646(fc1_io_in_646),
    .io_in_647(fc1_io_in_647),
    .io_in_648(fc1_io_in_648),
    .io_in_649(fc1_io_in_649),
    .io_in_650(fc1_io_in_650),
    .io_in_651(fc1_io_in_651),
    .io_in_652(fc1_io_in_652),
    .io_in_653(fc1_io_in_653),
    .io_in_654(fc1_io_in_654),
    .io_in_655(fc1_io_in_655),
    .io_in_656(fc1_io_in_656),
    .io_in_657(fc1_io_in_657),
    .io_in_658(fc1_io_in_658),
    .io_in_659(fc1_io_in_659),
    .io_in_660(fc1_io_in_660),
    .io_in_661(fc1_io_in_661),
    .io_in_662(fc1_io_in_662),
    .io_in_663(fc1_io_in_663),
    .io_in_664(fc1_io_in_664),
    .io_in_665(fc1_io_in_665),
    .io_in_666(fc1_io_in_666),
    .io_in_667(fc1_io_in_667),
    .io_in_668(fc1_io_in_668),
    .io_in_669(fc1_io_in_669),
    .io_in_670(fc1_io_in_670),
    .io_in_673(fc1_io_in_673),
    .io_in_674(fc1_io_in_674),
    .io_in_675(fc1_io_in_675),
    .io_in_676(fc1_io_in_676),
    .io_in_677(fc1_io_in_677),
    .io_in_678(fc1_io_in_678),
    .io_in_679(fc1_io_in_679),
    .io_in_680(fc1_io_in_680),
    .io_in_681(fc1_io_in_681),
    .io_in_682(fc1_io_in_682),
    .io_in_683(fc1_io_in_683),
    .io_in_684(fc1_io_in_684),
    .io_in_685(fc1_io_in_685),
    .io_in_686(fc1_io_in_686),
    .io_in_687(fc1_io_in_687),
    .io_in_688(fc1_io_in_688),
    .io_in_689(fc1_io_in_689),
    .io_in_690(fc1_io_in_690),
    .io_in_691(fc1_io_in_691),
    .io_in_692(fc1_io_in_692),
    .io_in_693(fc1_io_in_693),
    .io_in_694(fc1_io_in_694),
    .io_in_695(fc1_io_in_695),
    .io_in_696(fc1_io_in_696),
    .io_in_697(fc1_io_in_697),
    .io_in_698(fc1_io_in_698),
    .io_in_699(fc1_io_in_699),
    .io_in_702(fc1_io_in_702),
    .io_in_703(fc1_io_in_703),
    .io_in_704(fc1_io_in_704),
    .io_in_705(fc1_io_in_705),
    .io_in_706(fc1_io_in_706),
    .io_in_707(fc1_io_in_707),
    .io_in_708(fc1_io_in_708),
    .io_in_709(fc1_io_in_709),
    .io_in_710(fc1_io_in_710),
    .io_in_711(fc1_io_in_711),
    .io_in_712(fc1_io_in_712),
    .io_in_713(fc1_io_in_713),
    .io_in_714(fc1_io_in_714),
    .io_in_715(fc1_io_in_715),
    .io_in_716(fc1_io_in_716),
    .io_in_717(fc1_io_in_717),
    .io_in_718(fc1_io_in_718),
    .io_in_719(fc1_io_in_719),
    .io_in_720(fc1_io_in_720),
    .io_in_721(fc1_io_in_721),
    .io_in_722(fc1_io_in_722),
    .io_in_723(fc1_io_in_723),
    .io_in_724(fc1_io_in_724),
    .io_in_725(fc1_io_in_725),
    .io_in_726(fc1_io_in_726),
    .io_in_728(fc1_io_in_728),
    .io_in_729(fc1_io_in_729),
    .io_in_731(fc1_io_in_731),
    .io_in_732(fc1_io_in_732),
    .io_in_733(fc1_io_in_733),
    .io_in_734(fc1_io_in_734),
    .io_in_735(fc1_io_in_735),
    .io_in_736(fc1_io_in_736),
    .io_in_737(fc1_io_in_737),
    .io_in_738(fc1_io_in_738),
    .io_in_739(fc1_io_in_739),
    .io_in_740(fc1_io_in_740),
    .io_in_741(fc1_io_in_741),
    .io_in_742(fc1_io_in_742),
    .io_in_743(fc1_io_in_743),
    .io_in_744(fc1_io_in_744),
    .io_in_745(fc1_io_in_745),
    .io_in_746(fc1_io_in_746),
    .io_in_747(fc1_io_in_747),
    .io_in_748(fc1_io_in_748),
    .io_in_749(fc1_io_in_749),
    .io_in_750(fc1_io_in_750),
    .io_in_751(fc1_io_in_751),
    .io_in_752(fc1_io_in_752),
    .io_in_753(fc1_io_in_753),
    .io_in_756(fc1_io_in_756),
    .io_in_758(fc1_io_in_758),
    .io_in_760(fc1_io_in_760),
    .io_in_761(fc1_io_in_761),
    .io_in_762(fc1_io_in_762),
    .io_in_763(fc1_io_in_763),
    .io_in_764(fc1_io_in_764),
    .io_in_765(fc1_io_in_765),
    .io_in_766(fc1_io_in_766),
    .io_in_767(fc1_io_in_767),
    .io_in_768(fc1_io_in_768),
    .io_in_769(fc1_io_in_769),
    .io_in_770(fc1_io_in_770),
    .io_in_771(fc1_io_in_771),
    .io_in_772(fc1_io_in_772),
    .io_in_773(fc1_io_in_773),
    .io_in_774(fc1_io_in_774),
    .io_in_775(fc1_io_in_775),
    .io_in_776(fc1_io_in_776),
    .io_in_777(fc1_io_in_777),
    .io_in_778(fc1_io_in_778),
    .io_in_779(fc1_io_in_779),
    .io_in_780(fc1_io_in_780),
    .io_out_0(fc1_io_out_0),
    .io_out_1(fc1_io_out_1),
    .io_out_2(fc1_io_out_2),
    .io_out_3(fc1_io_out_3),
    .io_out_4(fc1_io_out_4),
    .io_out_5(fc1_io_out_5),
    .io_out_6(fc1_io_out_6),
    .io_out_7(fc1_io_out_7),
    .io_out_8(fc1_io_out_8),
    .io_out_9(fc1_io_out_9),
    .io_out_10(fc1_io_out_10),
    .io_out_11(fc1_io_out_11),
    .io_out_12(fc1_io_out_12),
    .io_out_13(fc1_io_out_13),
    .io_out_14(fc1_io_out_14),
    .io_out_15(fc1_io_out_15)
  );
  BN_BI bn_bi1 ( // @[Models.scala 22:24:@54610.4]
    .io_in_0(bn_bi1_io_in_0),
    .io_in_1(bn_bi1_io_in_1),
    .io_in_2(bn_bi1_io_in_2),
    .io_in_3(bn_bi1_io_in_3),
    .io_in_4(bn_bi1_io_in_4),
    .io_in_5(bn_bi1_io_in_5),
    .io_in_6(bn_bi1_io_in_6),
    .io_in_7(bn_bi1_io_in_7),
    .io_in_8(bn_bi1_io_in_8),
    .io_in_9(bn_bi1_io_in_9),
    .io_in_10(bn_bi1_io_in_10),
    .io_in_11(bn_bi1_io_in_11),
    .io_in_12(bn_bi1_io_in_12),
    .io_in_13(bn_bi1_io_in_13),
    .io_in_14(bn_bi1_io_in_14),
    .io_in_15(bn_bi1_io_in_15),
    .io_out_0(bn_bi1_io_out_0),
    .io_out_1(bn_bi1_io_out_1),
    .io_out_2(bn_bi1_io_out_2),
    .io_out_3(bn_bi1_io_out_3),
    .io_out_4(bn_bi1_io_out_4),
    .io_out_5(bn_bi1_io_out_5),
    .io_out_6(bn_bi1_io_out_6),
    .io_out_7(bn_bi1_io_out_7),
    .io_out_8(bn_bi1_io_out_8),
    .io_out_9(bn_bi1_io_out_9),
    .io_out_10(bn_bi1_io_out_10),
    .io_out_11(bn_bi1_io_out_11),
    .io_out_12(bn_bi1_io_out_12),
    .io_out_13(bn_bi1_io_out_13),
    .io_out_14(bn_bi1_io_out_14),
    .io_out_15(bn_bi1_io_out_15)
  );
  Linear_p_1 fc2 ( // @[Models.scala 26:15:@54613.4]
    .io_in_0(fc2_io_in_0),
    .io_in_1(fc2_io_in_1),
    .io_in_2(fc2_io_in_2),
    .io_in_3(fc2_io_in_3),
    .io_in_4(fc2_io_in_4),
    .io_in_5(fc2_io_in_5),
    .io_in_6(fc2_io_in_6),
    .io_in_7(fc2_io_in_7),
    .io_in_8(fc2_io_in_8),
    .io_in_9(fc2_io_in_9),
    .io_in_10(fc2_io_in_10),
    .io_in_11(fc2_io_in_11),
    .io_in_12(fc2_io_in_12),
    .io_in_13(fc2_io_in_13),
    .io_in_14(fc2_io_in_14),
    .io_in_15(fc2_io_in_15),
    .io_out_0(fc2_io_out_0),
    .io_out_1(fc2_io_out_1),
    .io_out_2(fc2_io_out_2),
    .io_out_3(fc2_io_out_3),
    .io_out_4(fc2_io_out_4),
    .io_out_5(fc2_io_out_5),
    .io_out_6(fc2_io_out_6),
    .io_out_7(fc2_io_out_7),
    .io_out_8(fc2_io_out_8),
    .io_out_9(fc2_io_out_9),
    .io_out_10(fc2_io_out_10),
    .io_out_11(fc2_io_out_11),
    .io_out_12(fc2_io_out_12),
    .io_out_13(fc2_io_out_13),
    .io_out_14(fc2_io_out_14),
    .io_out_15(fc2_io_out_15)
  );
  BN_BI_1 bn_bi2 ( // @[Models.scala 35:24:@54622.4]
    .io_in_0(bn_bi2_io_in_0),
    .io_in_1(bn_bi2_io_in_1),
    .io_in_2(bn_bi2_io_in_2),
    .io_in_3(bn_bi2_io_in_3),
    .io_in_4(bn_bi2_io_in_4),
    .io_in_5(bn_bi2_io_in_5),
    .io_in_6(bn_bi2_io_in_6),
    .io_in_7(bn_bi2_io_in_7),
    .io_in_8(bn_bi2_io_in_8),
    .io_in_9(bn_bi2_io_in_9),
    .io_in_10(bn_bi2_io_in_10),
    .io_in_11(bn_bi2_io_in_11),
    .io_in_12(bn_bi2_io_in_12),
    .io_in_13(bn_bi2_io_in_13),
    .io_in_14(bn_bi2_io_in_14),
    .io_in_15(bn_bi2_io_in_15),
    .io_out_0(bn_bi2_io_out_0),
    .io_out_1(bn_bi2_io_out_1),
    .io_out_2(bn_bi2_io_out_2),
    .io_out_3(bn_bi2_io_out_3),
    .io_out_4(bn_bi2_io_out_4),
    .io_out_5(bn_bi2_io_out_5),
    .io_out_6(bn_bi2_io_out_6),
    .io_out_7(bn_bi2_io_out_7),
    .io_out_8(bn_bi2_io_out_8),
    .io_out_9(bn_bi2_io_out_9),
    .io_out_10(bn_bi2_io_out_10),
    .io_out_11(bn_bi2_io_out_11),
    .io_out_12(bn_bi2_io_out_12),
    .io_out_13(bn_bi2_io_out_13),
    .io_out_14(bn_bi2_io_out_14),
    .io_out_15(bn_bi2_io_out_15)
  );
  Linear_p_2 fc3 ( // @[Models.scala 39:15:@54625.4]
    .io_in_0(fc3_io_in_0),
    .io_in_1(fc3_io_in_1),
    .io_in_2(fc3_io_in_2),
    .io_in_3(fc3_io_in_3),
    .io_in_4(fc3_io_in_4),
    .io_in_5(fc3_io_in_5),
    .io_in_6(fc3_io_in_6),
    .io_in_7(fc3_io_in_7),
    .io_in_8(fc3_io_in_8),
    .io_in_9(fc3_io_in_9),
    .io_in_10(fc3_io_in_10),
    .io_in_11(fc3_io_in_11),
    .io_in_12(fc3_io_in_12),
    .io_in_13(fc3_io_in_13),
    .io_in_14(fc3_io_in_14),
    .io_in_15(fc3_io_in_15),
    .io_out_0(fc3_io_out_0),
    .io_out_1(fc3_io_out_1),
    .io_out_2(fc3_io_out_2),
    .io_out_3(fc3_io_out_3),
    .io_out_4(fc3_io_out_4),
    .io_out_5(fc3_io_out_5),
    .io_out_6(fc3_io_out_6),
    .io_out_7(fc3_io_out_7),
    .io_out_8(fc3_io_out_8),
    .io_out_9(fc3_io_out_9)
  );
  SBN_2 bn3 ( // @[Models.scala 45:21:@54628.4]
    .io_in_0(bn3_io_in_0),
    .io_in_1(bn3_io_in_1),
    .io_in_2(bn3_io_in_2),
    .io_in_3(bn3_io_in_3),
    .io_in_4(bn3_io_in_4),
    .io_in_5(bn3_io_in_5),
    .io_in_6(bn3_io_in_6),
    .io_in_7(bn3_io_in_7),
    .io_in_8(bn3_io_in_8),
    .io_in_9(bn3_io_in_9),
    .io_out_0(bn3_io_out_0),
    .io_out_1(bn3_io_out_1),
    .io_out_2(bn3_io_out_2),
    .io_out_3(bn3_io_out_3),
    .io_out_4(bn3_io_out_4),
    .io_out_5(bn3_io_out_5),
    .io_out_6(bn3_io_out_6),
    .io_out_7(bn3_io_out_7),
    .io_out_8(bn3_io_out_8),
    .io_out_9(bn3_io_out_9)
  );
  assign io_out_0 = {{4{bn3_io_out_0[5]}},bn3_io_out_0};
  assign io_out_1 = {{4{bn3_io_out_1[5]}},bn3_io_out_1};
  assign io_out_2 = {{4{bn3_io_out_2[5]}},bn3_io_out_2};
  assign io_out_3 = {{4{bn3_io_out_3[5]}},bn3_io_out_3};
  assign io_out_4 = {{4{bn3_io_out_4[5]}},bn3_io_out_4};
  assign io_out_5 = {{4{bn3_io_out_5[5]}},bn3_io_out_5};
  assign io_out_6 = {{4{bn3_io_out_6[5]}},bn3_io_out_6};
  assign io_out_7 = {{4{bn3_io_out_7[5]}},bn3_io_out_7};
  assign io_out_8 = {{4{bn3_io_out_8[5]}},bn3_io_out_8};
  assign io_out_9 = {{4{bn3_io_out_9[5]}},bn3_io_out_9};
  assign fc1_io_in_0 = io_in_0;
  assign fc1_io_in_3 = io_in_3;
  assign fc1_io_in_5 = io_in_5;
  assign fc1_io_in_10 = io_in_10;
  assign fc1_io_in_12 = io_in_12;
  assign fc1_io_in_13 = io_in_13;
  assign fc1_io_in_14 = io_in_14;
  assign fc1_io_in_15 = io_in_15;
  assign fc1_io_in_19 = io_in_19;
  assign fc1_io_in_21 = io_in_21;
  assign fc1_io_in_23 = io_in_23;
  assign fc1_io_in_25 = io_in_25;
  assign fc1_io_in_28 = io_in_28;
  assign fc1_io_in_29 = io_in_29;
  assign fc1_io_in_30 = io_in_30;
  assign fc1_io_in_32 = io_in_32;
  assign fc1_io_in_33 = io_in_33;
  assign fc1_io_in_34 = io_in_34;
  assign fc1_io_in_35 = io_in_35;
  assign fc1_io_in_36 = io_in_36;
  assign fc1_io_in_37 = io_in_37;
  assign fc1_io_in_38 = io_in_38;
  assign fc1_io_in_39 = io_in_39;
  assign fc1_io_in_40 = io_in_40;
  assign fc1_io_in_41 = io_in_41;
  assign fc1_io_in_42 = io_in_42;
  assign fc1_io_in_43 = io_in_43;
  assign fc1_io_in_44 = io_in_44;
  assign fc1_io_in_45 = io_in_45;
  assign fc1_io_in_46 = io_in_46;
  assign fc1_io_in_47 = io_in_47;
  assign fc1_io_in_48 = io_in_48;
  assign fc1_io_in_49 = io_in_49;
  assign fc1_io_in_50 = io_in_50;
  assign fc1_io_in_51 = io_in_51;
  assign fc1_io_in_52 = io_in_52;
  assign fc1_io_in_54 = io_in_54;
  assign fc1_io_in_56 = io_in_56;
  assign fc1_io_in_59 = io_in_59;
  assign fc1_io_in_60 = io_in_60;
  assign fc1_io_in_61 = io_in_61;
  assign fc1_io_in_62 = io_in_62;
  assign fc1_io_in_63 = io_in_63;
  assign fc1_io_in_64 = io_in_64;
  assign fc1_io_in_65 = io_in_65;
  assign fc1_io_in_66 = io_in_66;
  assign fc1_io_in_67 = io_in_67;
  assign fc1_io_in_68 = io_in_68;
  assign fc1_io_in_69 = io_in_69;
  assign fc1_io_in_70 = io_in_70;
  assign fc1_io_in_71 = io_in_71;
  assign fc1_io_in_72 = io_in_72;
  assign fc1_io_in_73 = io_in_73;
  assign fc1_io_in_74 = io_in_74;
  assign fc1_io_in_75 = io_in_75;
  assign fc1_io_in_76 = io_in_76;
  assign fc1_io_in_77 = io_in_77;
  assign fc1_io_in_78 = io_in_78;
  assign fc1_io_in_79 = io_in_79;
  assign fc1_io_in_80 = io_in_80;
  assign fc1_io_in_81 = io_in_81;
  assign fc1_io_in_82 = io_in_82;
  assign fc1_io_in_83 = io_in_83;
  assign fc1_io_in_86 = io_in_86;
  assign fc1_io_in_87 = io_in_87;
  assign fc1_io_in_88 = io_in_88;
  assign fc1_io_in_89 = io_in_89;
  assign fc1_io_in_90 = io_in_90;
  assign fc1_io_in_91 = io_in_91;
  assign fc1_io_in_92 = io_in_92;
  assign fc1_io_in_93 = io_in_93;
  assign fc1_io_in_94 = io_in_94;
  assign fc1_io_in_95 = io_in_95;
  assign fc1_io_in_96 = io_in_96;
  assign fc1_io_in_97 = io_in_97;
  assign fc1_io_in_98 = io_in_98;
  assign fc1_io_in_99 = io_in_99;
  assign fc1_io_in_100 = io_in_100;
  assign fc1_io_in_101 = io_in_101;
  assign fc1_io_in_102 = io_in_102;
  assign fc1_io_in_103 = io_in_103;
  assign fc1_io_in_104 = io_in_104;
  assign fc1_io_in_105 = io_in_105;
  assign fc1_io_in_106 = io_in_106;
  assign fc1_io_in_107 = io_in_107;
  assign fc1_io_in_108 = io_in_108;
  assign fc1_io_in_109 = io_in_109;
  assign fc1_io_in_110 = io_in_110;
  assign fc1_io_in_113 = io_in_113;
  assign fc1_io_in_114 = io_in_114;
  assign fc1_io_in_115 = io_in_115;
  assign fc1_io_in_116 = io_in_116;
  assign fc1_io_in_117 = io_in_117;
  assign fc1_io_in_118 = io_in_118;
  assign fc1_io_in_119 = io_in_119;
  assign fc1_io_in_120 = io_in_120;
  assign fc1_io_in_121 = io_in_121;
  assign fc1_io_in_122 = io_in_122;
  assign fc1_io_in_123 = io_in_123;
  assign fc1_io_in_124 = io_in_124;
  assign fc1_io_in_125 = io_in_125;
  assign fc1_io_in_126 = io_in_126;
  assign fc1_io_in_127 = io_in_127;
  assign fc1_io_in_128 = io_in_128;
  assign fc1_io_in_129 = io_in_129;
  assign fc1_io_in_130 = io_in_130;
  assign fc1_io_in_131 = io_in_131;
  assign fc1_io_in_132 = io_in_132;
  assign fc1_io_in_133 = io_in_133;
  assign fc1_io_in_134 = io_in_134;
  assign fc1_io_in_135 = io_in_135;
  assign fc1_io_in_136 = io_in_136;
  assign fc1_io_in_137 = io_in_137;
  assign fc1_io_in_138 = io_in_138;
  assign fc1_io_in_139 = io_in_139;
  assign fc1_io_in_140 = io_in_140;
  assign fc1_io_in_142 = io_in_142;
  assign fc1_io_in_143 = io_in_143;
  assign fc1_io_in_144 = io_in_144;
  assign fc1_io_in_145 = io_in_145;
  assign fc1_io_in_146 = io_in_146;
  assign fc1_io_in_147 = io_in_147;
  assign fc1_io_in_148 = io_in_148;
  assign fc1_io_in_149 = io_in_149;
  assign fc1_io_in_150 = io_in_150;
  assign fc1_io_in_151 = io_in_151;
  assign fc1_io_in_152 = io_in_152;
  assign fc1_io_in_153 = io_in_153;
  assign fc1_io_in_154 = io_in_154;
  assign fc1_io_in_155 = io_in_155;
  assign fc1_io_in_156 = io_in_156;
  assign fc1_io_in_157 = io_in_157;
  assign fc1_io_in_158 = io_in_158;
  assign fc1_io_in_159 = io_in_159;
  assign fc1_io_in_160 = io_in_160;
  assign fc1_io_in_161 = io_in_161;
  assign fc1_io_in_162 = io_in_162;
  assign fc1_io_in_163 = io_in_163;
  assign fc1_io_in_164 = io_in_164;
  assign fc1_io_in_165 = io_in_165;
  assign fc1_io_in_166 = io_in_166;
  assign fc1_io_in_167 = io_in_167;
  assign fc1_io_in_168 = io_in_168;
  assign fc1_io_in_169 = io_in_169;
  assign fc1_io_in_170 = io_in_170;
  assign fc1_io_in_171 = io_in_171;
  assign fc1_io_in_172 = io_in_172;
  assign fc1_io_in_173 = io_in_173;
  assign fc1_io_in_174 = io_in_174;
  assign fc1_io_in_175 = io_in_175;
  assign fc1_io_in_176 = io_in_176;
  assign fc1_io_in_177 = io_in_177;
  assign fc1_io_in_178 = io_in_178;
  assign fc1_io_in_179 = io_in_179;
  assign fc1_io_in_180 = io_in_180;
  assign fc1_io_in_181 = io_in_181;
  assign fc1_io_in_182 = io_in_182;
  assign fc1_io_in_183 = io_in_183;
  assign fc1_io_in_184 = io_in_184;
  assign fc1_io_in_185 = io_in_185;
  assign fc1_io_in_186 = io_in_186;
  assign fc1_io_in_187 = io_in_187;
  assign fc1_io_in_188 = io_in_188;
  assign fc1_io_in_189 = io_in_189;
  assign fc1_io_in_190 = io_in_190;
  assign fc1_io_in_191 = io_in_191;
  assign fc1_io_in_192 = io_in_192;
  assign fc1_io_in_193 = io_in_193;
  assign fc1_io_in_194 = io_in_194;
  assign fc1_io_in_195 = io_in_195;
  assign fc1_io_in_196 = io_in_196;
  assign fc1_io_in_197 = io_in_197;
  assign fc1_io_in_198 = io_in_198;
  assign fc1_io_in_199 = io_in_199;
  assign fc1_io_in_200 = io_in_200;
  assign fc1_io_in_201 = io_in_201;
  assign fc1_io_in_202 = io_in_202;
  assign fc1_io_in_203 = io_in_203;
  assign fc1_io_in_204 = io_in_204;
  assign fc1_io_in_205 = io_in_205;
  assign fc1_io_in_206 = io_in_206;
  assign fc1_io_in_207 = io_in_207;
  assign fc1_io_in_208 = io_in_208;
  assign fc1_io_in_209 = io_in_209;
  assign fc1_io_in_210 = io_in_210;
  assign fc1_io_in_211 = io_in_211;
  assign fc1_io_in_212 = io_in_212;
  assign fc1_io_in_213 = io_in_213;
  assign fc1_io_in_214 = io_in_214;
  assign fc1_io_in_215 = io_in_215;
  assign fc1_io_in_216 = io_in_216;
  assign fc1_io_in_217 = io_in_217;
  assign fc1_io_in_218 = io_in_218;
  assign fc1_io_in_219 = io_in_219;
  assign fc1_io_in_220 = io_in_220;
  assign fc1_io_in_221 = io_in_221;
  assign fc1_io_in_222 = io_in_222;
  assign fc1_io_in_223 = io_in_223;
  assign fc1_io_in_224 = io_in_224;
  assign fc1_io_in_225 = io_in_225;
  assign fc1_io_in_226 = io_in_226;
  assign fc1_io_in_227 = io_in_227;
  assign fc1_io_in_228 = io_in_228;
  assign fc1_io_in_229 = io_in_229;
  assign fc1_io_in_230 = io_in_230;
  assign fc1_io_in_231 = io_in_231;
  assign fc1_io_in_232 = io_in_232;
  assign fc1_io_in_233 = io_in_233;
  assign fc1_io_in_234 = io_in_234;
  assign fc1_io_in_235 = io_in_235;
  assign fc1_io_in_236 = io_in_236;
  assign fc1_io_in_237 = io_in_237;
  assign fc1_io_in_238 = io_in_238;
  assign fc1_io_in_239 = io_in_239;
  assign fc1_io_in_240 = io_in_240;
  assign fc1_io_in_241 = io_in_241;
  assign fc1_io_in_242 = io_in_242;
  assign fc1_io_in_243 = io_in_243;
  assign fc1_io_in_244 = io_in_244;
  assign fc1_io_in_245 = io_in_245;
  assign fc1_io_in_246 = io_in_246;
  assign fc1_io_in_247 = io_in_247;
  assign fc1_io_in_248 = io_in_248;
  assign fc1_io_in_249 = io_in_249;
  assign fc1_io_in_250 = io_in_250;
  assign fc1_io_in_251 = io_in_251;
  assign fc1_io_in_252 = io_in_252;
  assign fc1_io_in_253 = io_in_253;
  assign fc1_io_in_254 = io_in_254;
  assign fc1_io_in_255 = io_in_255;
  assign fc1_io_in_256 = io_in_256;
  assign fc1_io_in_257 = io_in_257;
  assign fc1_io_in_258 = io_in_258;
  assign fc1_io_in_259 = io_in_259;
  assign fc1_io_in_260 = io_in_260;
  assign fc1_io_in_261 = io_in_261;
  assign fc1_io_in_262 = io_in_262;
  assign fc1_io_in_263 = io_in_263;
  assign fc1_io_in_264 = io_in_264;
  assign fc1_io_in_265 = io_in_265;
  assign fc1_io_in_266 = io_in_266;
  assign fc1_io_in_267 = io_in_267;
  assign fc1_io_in_268 = io_in_268;
  assign fc1_io_in_269 = io_in_269;
  assign fc1_io_in_270 = io_in_270;
  assign fc1_io_in_271 = io_in_271;
  assign fc1_io_in_272 = io_in_272;
  assign fc1_io_in_273 = io_in_273;
  assign fc1_io_in_274 = io_in_274;
  assign fc1_io_in_275 = io_in_275;
  assign fc1_io_in_276 = io_in_276;
  assign fc1_io_in_277 = io_in_277;
  assign fc1_io_in_278 = io_in_278;
  assign fc1_io_in_279 = io_in_279;
  assign fc1_io_in_280 = io_in_280;
  assign fc1_io_in_281 = io_in_281;
  assign fc1_io_in_282 = io_in_282;
  assign fc1_io_in_283 = io_in_283;
  assign fc1_io_in_284 = io_in_284;
  assign fc1_io_in_285 = io_in_285;
  assign fc1_io_in_286 = io_in_286;
  assign fc1_io_in_287 = io_in_287;
  assign fc1_io_in_288 = io_in_288;
  assign fc1_io_in_289 = io_in_289;
  assign fc1_io_in_290 = io_in_290;
  assign fc1_io_in_291 = io_in_291;
  assign fc1_io_in_292 = io_in_292;
  assign fc1_io_in_293 = io_in_293;
  assign fc1_io_in_294 = io_in_294;
  assign fc1_io_in_295 = io_in_295;
  assign fc1_io_in_296 = io_in_296;
  assign fc1_io_in_297 = io_in_297;
  assign fc1_io_in_298 = io_in_298;
  assign fc1_io_in_299 = io_in_299;
  assign fc1_io_in_300 = io_in_300;
  assign fc1_io_in_301 = io_in_301;
  assign fc1_io_in_302 = io_in_302;
  assign fc1_io_in_303 = io_in_303;
  assign fc1_io_in_304 = io_in_304;
  assign fc1_io_in_305 = io_in_305;
  assign fc1_io_in_306 = io_in_306;
  assign fc1_io_in_307 = io_in_307;
  assign fc1_io_in_308 = io_in_308;
  assign fc1_io_in_309 = io_in_309;
  assign fc1_io_in_310 = io_in_310;
  assign fc1_io_in_311 = io_in_311;
  assign fc1_io_in_312 = io_in_312;
  assign fc1_io_in_313 = io_in_313;
  assign fc1_io_in_314 = io_in_314;
  assign fc1_io_in_315 = io_in_315;
  assign fc1_io_in_316 = io_in_316;
  assign fc1_io_in_317 = io_in_317;
  assign fc1_io_in_318 = io_in_318;
  assign fc1_io_in_319 = io_in_319;
  assign fc1_io_in_320 = io_in_320;
  assign fc1_io_in_321 = io_in_321;
  assign fc1_io_in_322 = io_in_322;
  assign fc1_io_in_323 = io_in_323;
  assign fc1_io_in_324 = io_in_324;
  assign fc1_io_in_325 = io_in_325;
  assign fc1_io_in_326 = io_in_326;
  assign fc1_io_in_327 = io_in_327;
  assign fc1_io_in_328 = io_in_328;
  assign fc1_io_in_329 = io_in_329;
  assign fc1_io_in_330 = io_in_330;
  assign fc1_io_in_331 = io_in_331;
  assign fc1_io_in_332 = io_in_332;
  assign fc1_io_in_333 = io_in_333;
  assign fc1_io_in_334 = io_in_334;
  assign fc1_io_in_335 = io_in_335;
  assign fc1_io_in_336 = io_in_336;
  assign fc1_io_in_337 = io_in_337;
  assign fc1_io_in_338 = io_in_338;
  assign fc1_io_in_339 = io_in_339;
  assign fc1_io_in_340 = io_in_340;
  assign fc1_io_in_341 = io_in_341;
  assign fc1_io_in_342 = io_in_342;
  assign fc1_io_in_343 = io_in_343;
  assign fc1_io_in_344 = io_in_344;
  assign fc1_io_in_345 = io_in_345;
  assign fc1_io_in_346 = io_in_346;
  assign fc1_io_in_347 = io_in_347;
  assign fc1_io_in_348 = io_in_348;
  assign fc1_io_in_349 = io_in_349;
  assign fc1_io_in_350 = io_in_350;
  assign fc1_io_in_351 = io_in_351;
  assign fc1_io_in_352 = io_in_352;
  assign fc1_io_in_353 = io_in_353;
  assign fc1_io_in_354 = io_in_354;
  assign fc1_io_in_355 = io_in_355;
  assign fc1_io_in_356 = io_in_356;
  assign fc1_io_in_357 = io_in_357;
  assign fc1_io_in_358 = io_in_358;
  assign fc1_io_in_359 = io_in_359;
  assign fc1_io_in_360 = io_in_360;
  assign fc1_io_in_361 = io_in_361;
  assign fc1_io_in_362 = io_in_362;
  assign fc1_io_in_363 = io_in_363;
  assign fc1_io_in_364 = io_in_364;
  assign fc1_io_in_365 = io_in_365;
  assign fc1_io_in_366 = io_in_366;
  assign fc1_io_in_367 = io_in_367;
  assign fc1_io_in_368 = io_in_368;
  assign fc1_io_in_369 = io_in_369;
  assign fc1_io_in_370 = io_in_370;
  assign fc1_io_in_371 = io_in_371;
  assign fc1_io_in_372 = io_in_372;
  assign fc1_io_in_373 = io_in_373;
  assign fc1_io_in_374 = io_in_374;
  assign fc1_io_in_375 = io_in_375;
  assign fc1_io_in_376 = io_in_376;
  assign fc1_io_in_377 = io_in_377;
  assign fc1_io_in_378 = io_in_378;
  assign fc1_io_in_379 = io_in_379;
  assign fc1_io_in_380 = io_in_380;
  assign fc1_io_in_381 = io_in_381;
  assign fc1_io_in_382 = io_in_382;
  assign fc1_io_in_383 = io_in_383;
  assign fc1_io_in_384 = io_in_384;
  assign fc1_io_in_385 = io_in_385;
  assign fc1_io_in_386 = io_in_386;
  assign fc1_io_in_387 = io_in_387;
  assign fc1_io_in_388 = io_in_388;
  assign fc1_io_in_389 = io_in_389;
  assign fc1_io_in_390 = io_in_390;
  assign fc1_io_in_391 = io_in_391;
  assign fc1_io_in_392 = io_in_392;
  assign fc1_io_in_393 = io_in_393;
  assign fc1_io_in_394 = io_in_394;
  assign fc1_io_in_395 = io_in_395;
  assign fc1_io_in_396 = io_in_396;
  assign fc1_io_in_397 = io_in_397;
  assign fc1_io_in_398 = io_in_398;
  assign fc1_io_in_399 = io_in_399;
  assign fc1_io_in_400 = io_in_400;
  assign fc1_io_in_401 = io_in_401;
  assign fc1_io_in_402 = io_in_402;
  assign fc1_io_in_403 = io_in_403;
  assign fc1_io_in_404 = io_in_404;
  assign fc1_io_in_405 = io_in_405;
  assign fc1_io_in_406 = io_in_406;
  assign fc1_io_in_407 = io_in_407;
  assign fc1_io_in_408 = io_in_408;
  assign fc1_io_in_409 = io_in_409;
  assign fc1_io_in_410 = io_in_410;
  assign fc1_io_in_411 = io_in_411;
  assign fc1_io_in_412 = io_in_412;
  assign fc1_io_in_413 = io_in_413;
  assign fc1_io_in_414 = io_in_414;
  assign fc1_io_in_415 = io_in_415;
  assign fc1_io_in_416 = io_in_416;
  assign fc1_io_in_417 = io_in_417;
  assign fc1_io_in_418 = io_in_418;
  assign fc1_io_in_419 = io_in_419;
  assign fc1_io_in_420 = io_in_420;
  assign fc1_io_in_421 = io_in_421;
  assign fc1_io_in_422 = io_in_422;
  assign fc1_io_in_423 = io_in_423;
  assign fc1_io_in_424 = io_in_424;
  assign fc1_io_in_425 = io_in_425;
  assign fc1_io_in_426 = io_in_426;
  assign fc1_io_in_427 = io_in_427;
  assign fc1_io_in_428 = io_in_428;
  assign fc1_io_in_429 = io_in_429;
  assign fc1_io_in_430 = io_in_430;
  assign fc1_io_in_431 = io_in_431;
  assign fc1_io_in_432 = io_in_432;
  assign fc1_io_in_433 = io_in_433;
  assign fc1_io_in_434 = io_in_434;
  assign fc1_io_in_435 = io_in_435;
  assign fc1_io_in_436 = io_in_436;
  assign fc1_io_in_437 = io_in_437;
  assign fc1_io_in_438 = io_in_438;
  assign fc1_io_in_439 = io_in_439;
  assign fc1_io_in_440 = io_in_440;
  assign fc1_io_in_441 = io_in_441;
  assign fc1_io_in_442 = io_in_442;
  assign fc1_io_in_443 = io_in_443;
  assign fc1_io_in_444 = io_in_444;
  assign fc1_io_in_445 = io_in_445;
  assign fc1_io_in_446 = io_in_446;
  assign fc1_io_in_447 = io_in_447;
  assign fc1_io_in_448 = io_in_448;
  assign fc1_io_in_449 = io_in_449;
  assign fc1_io_in_450 = io_in_450;
  assign fc1_io_in_451 = io_in_451;
  assign fc1_io_in_452 = io_in_452;
  assign fc1_io_in_453 = io_in_453;
  assign fc1_io_in_454 = io_in_454;
  assign fc1_io_in_455 = io_in_455;
  assign fc1_io_in_456 = io_in_456;
  assign fc1_io_in_457 = io_in_457;
  assign fc1_io_in_458 = io_in_458;
  assign fc1_io_in_459 = io_in_459;
  assign fc1_io_in_460 = io_in_460;
  assign fc1_io_in_461 = io_in_461;
  assign fc1_io_in_462 = io_in_462;
  assign fc1_io_in_463 = io_in_463;
  assign fc1_io_in_464 = io_in_464;
  assign fc1_io_in_465 = io_in_465;
  assign fc1_io_in_466 = io_in_466;
  assign fc1_io_in_467 = io_in_467;
  assign fc1_io_in_468 = io_in_468;
  assign fc1_io_in_469 = io_in_469;
  assign fc1_io_in_470 = io_in_470;
  assign fc1_io_in_471 = io_in_471;
  assign fc1_io_in_472 = io_in_472;
  assign fc1_io_in_473 = io_in_473;
  assign fc1_io_in_474 = io_in_474;
  assign fc1_io_in_475 = io_in_475;
  assign fc1_io_in_476 = io_in_476;
  assign fc1_io_in_477 = io_in_477;
  assign fc1_io_in_478 = io_in_478;
  assign fc1_io_in_479 = io_in_479;
  assign fc1_io_in_480 = io_in_480;
  assign fc1_io_in_481 = io_in_481;
  assign fc1_io_in_482 = io_in_482;
  assign fc1_io_in_483 = io_in_483;
  assign fc1_io_in_484 = io_in_484;
  assign fc1_io_in_485 = io_in_485;
  assign fc1_io_in_486 = io_in_486;
  assign fc1_io_in_487 = io_in_487;
  assign fc1_io_in_488 = io_in_488;
  assign fc1_io_in_489 = io_in_489;
  assign fc1_io_in_490 = io_in_490;
  assign fc1_io_in_491 = io_in_491;
  assign fc1_io_in_492 = io_in_492;
  assign fc1_io_in_493 = io_in_493;
  assign fc1_io_in_494 = io_in_494;
  assign fc1_io_in_495 = io_in_495;
  assign fc1_io_in_496 = io_in_496;
  assign fc1_io_in_497 = io_in_497;
  assign fc1_io_in_498 = io_in_498;
  assign fc1_io_in_499 = io_in_499;
  assign fc1_io_in_500 = io_in_500;
  assign fc1_io_in_501 = io_in_501;
  assign fc1_io_in_502 = io_in_502;
  assign fc1_io_in_503 = io_in_503;
  assign fc1_io_in_504 = io_in_504;
  assign fc1_io_in_505 = io_in_505;
  assign fc1_io_in_506 = io_in_506;
  assign fc1_io_in_507 = io_in_507;
  assign fc1_io_in_508 = io_in_508;
  assign fc1_io_in_509 = io_in_509;
  assign fc1_io_in_510 = io_in_510;
  assign fc1_io_in_511 = io_in_511;
  assign fc1_io_in_512 = io_in_512;
  assign fc1_io_in_513 = io_in_513;
  assign fc1_io_in_514 = io_in_514;
  assign fc1_io_in_515 = io_in_515;
  assign fc1_io_in_516 = io_in_516;
  assign fc1_io_in_517 = io_in_517;
  assign fc1_io_in_518 = io_in_518;
  assign fc1_io_in_519 = io_in_519;
  assign fc1_io_in_520 = io_in_520;
  assign fc1_io_in_521 = io_in_521;
  assign fc1_io_in_522 = io_in_522;
  assign fc1_io_in_523 = io_in_523;
  assign fc1_io_in_524 = io_in_524;
  assign fc1_io_in_525 = io_in_525;
  assign fc1_io_in_526 = io_in_526;
  assign fc1_io_in_527 = io_in_527;
  assign fc1_io_in_528 = io_in_528;
  assign fc1_io_in_529 = io_in_529;
  assign fc1_io_in_530 = io_in_530;
  assign fc1_io_in_531 = io_in_531;
  assign fc1_io_in_532 = io_in_532;
  assign fc1_io_in_533 = io_in_533;
  assign fc1_io_in_534 = io_in_534;
  assign fc1_io_in_535 = io_in_535;
  assign fc1_io_in_536 = io_in_536;
  assign fc1_io_in_537 = io_in_537;
  assign fc1_io_in_538 = io_in_538;
  assign fc1_io_in_539 = io_in_539;
  assign fc1_io_in_540 = io_in_540;
  assign fc1_io_in_541 = io_in_541;
  assign fc1_io_in_542 = io_in_542;
  assign fc1_io_in_543 = io_in_543;
  assign fc1_io_in_544 = io_in_544;
  assign fc1_io_in_545 = io_in_545;
  assign fc1_io_in_546 = io_in_546;
  assign fc1_io_in_547 = io_in_547;
  assign fc1_io_in_548 = io_in_548;
  assign fc1_io_in_549 = io_in_549;
  assign fc1_io_in_550 = io_in_550;
  assign fc1_io_in_551 = io_in_551;
  assign fc1_io_in_552 = io_in_552;
  assign fc1_io_in_553 = io_in_553;
  assign fc1_io_in_554 = io_in_554;
  assign fc1_io_in_555 = io_in_555;
  assign fc1_io_in_556 = io_in_556;
  assign fc1_io_in_557 = io_in_557;
  assign fc1_io_in_558 = io_in_558;
  assign fc1_io_in_559 = io_in_559;
  assign fc1_io_in_561 = io_in_561;
  assign fc1_io_in_562 = io_in_562;
  assign fc1_io_in_563 = io_in_563;
  assign fc1_io_in_564 = io_in_564;
  assign fc1_io_in_565 = io_in_565;
  assign fc1_io_in_566 = io_in_566;
  assign fc1_io_in_567 = io_in_567;
  assign fc1_io_in_568 = io_in_568;
  assign fc1_io_in_569 = io_in_569;
  assign fc1_io_in_570 = io_in_570;
  assign fc1_io_in_571 = io_in_571;
  assign fc1_io_in_572 = io_in_572;
  assign fc1_io_in_573 = io_in_573;
  assign fc1_io_in_574 = io_in_574;
  assign fc1_io_in_575 = io_in_575;
  assign fc1_io_in_576 = io_in_576;
  assign fc1_io_in_577 = io_in_577;
  assign fc1_io_in_578 = io_in_578;
  assign fc1_io_in_579 = io_in_579;
  assign fc1_io_in_580 = io_in_580;
  assign fc1_io_in_581 = io_in_581;
  assign fc1_io_in_582 = io_in_582;
  assign fc1_io_in_583 = io_in_583;
  assign fc1_io_in_584 = io_in_584;
  assign fc1_io_in_585 = io_in_585;
  assign fc1_io_in_586 = io_in_586;
  assign fc1_io_in_587 = io_in_587;
  assign fc1_io_in_588 = io_in_588;
  assign fc1_io_in_589 = io_in_589;
  assign fc1_io_in_590 = io_in_590;
  assign fc1_io_in_591 = io_in_591;
  assign fc1_io_in_592 = io_in_592;
  assign fc1_io_in_593 = io_in_593;
  assign fc1_io_in_594 = io_in_594;
  assign fc1_io_in_595 = io_in_595;
  assign fc1_io_in_596 = io_in_596;
  assign fc1_io_in_597 = io_in_597;
  assign fc1_io_in_598 = io_in_598;
  assign fc1_io_in_599 = io_in_599;
  assign fc1_io_in_600 = io_in_600;
  assign fc1_io_in_601 = io_in_601;
  assign fc1_io_in_602 = io_in_602;
  assign fc1_io_in_603 = io_in_603;
  assign fc1_io_in_604 = io_in_604;
  assign fc1_io_in_605 = io_in_605;
  assign fc1_io_in_606 = io_in_606;
  assign fc1_io_in_607 = io_in_607;
  assign fc1_io_in_608 = io_in_608;
  assign fc1_io_in_609 = io_in_609;
  assign fc1_io_in_610 = io_in_610;
  assign fc1_io_in_611 = io_in_611;
  assign fc1_io_in_612 = io_in_612;
  assign fc1_io_in_613 = io_in_613;
  assign fc1_io_in_614 = io_in_614;
  assign fc1_io_in_615 = io_in_615;
  assign fc1_io_in_616 = io_in_616;
  assign fc1_io_in_617 = io_in_617;
  assign fc1_io_in_618 = io_in_618;
  assign fc1_io_in_619 = io_in_619;
  assign fc1_io_in_620 = io_in_620;
  assign fc1_io_in_621 = io_in_621;
  assign fc1_io_in_622 = io_in_622;
  assign fc1_io_in_623 = io_in_623;
  assign fc1_io_in_624 = io_in_624;
  assign fc1_io_in_625 = io_in_625;
  assign fc1_io_in_626 = io_in_626;
  assign fc1_io_in_627 = io_in_627;
  assign fc1_io_in_628 = io_in_628;
  assign fc1_io_in_629 = io_in_629;
  assign fc1_io_in_630 = io_in_630;
  assign fc1_io_in_631 = io_in_631;
  assign fc1_io_in_632 = io_in_632;
  assign fc1_io_in_633 = io_in_633;
  assign fc1_io_in_634 = io_in_634;
  assign fc1_io_in_635 = io_in_635;
  assign fc1_io_in_636 = io_in_636;
  assign fc1_io_in_637 = io_in_637;
  assign fc1_io_in_638 = io_in_638;
  assign fc1_io_in_639 = io_in_639;
  assign fc1_io_in_640 = io_in_640;
  assign fc1_io_in_641 = io_in_641;
  assign fc1_io_in_642 = io_in_642;
  assign fc1_io_in_646 = io_in_646;
  assign fc1_io_in_647 = io_in_647;
  assign fc1_io_in_648 = io_in_648;
  assign fc1_io_in_649 = io_in_649;
  assign fc1_io_in_650 = io_in_650;
  assign fc1_io_in_651 = io_in_651;
  assign fc1_io_in_652 = io_in_652;
  assign fc1_io_in_653 = io_in_653;
  assign fc1_io_in_654 = io_in_654;
  assign fc1_io_in_655 = io_in_655;
  assign fc1_io_in_656 = io_in_656;
  assign fc1_io_in_657 = io_in_657;
  assign fc1_io_in_658 = io_in_658;
  assign fc1_io_in_659 = io_in_659;
  assign fc1_io_in_660 = io_in_660;
  assign fc1_io_in_661 = io_in_661;
  assign fc1_io_in_662 = io_in_662;
  assign fc1_io_in_663 = io_in_663;
  assign fc1_io_in_664 = io_in_664;
  assign fc1_io_in_665 = io_in_665;
  assign fc1_io_in_666 = io_in_666;
  assign fc1_io_in_667 = io_in_667;
  assign fc1_io_in_668 = io_in_668;
  assign fc1_io_in_669 = io_in_669;
  assign fc1_io_in_670 = io_in_670;
  assign fc1_io_in_673 = io_in_673;
  assign fc1_io_in_674 = io_in_674;
  assign fc1_io_in_675 = io_in_675;
  assign fc1_io_in_676 = io_in_676;
  assign fc1_io_in_677 = io_in_677;
  assign fc1_io_in_678 = io_in_678;
  assign fc1_io_in_679 = io_in_679;
  assign fc1_io_in_680 = io_in_680;
  assign fc1_io_in_681 = io_in_681;
  assign fc1_io_in_682 = io_in_682;
  assign fc1_io_in_683 = io_in_683;
  assign fc1_io_in_684 = io_in_684;
  assign fc1_io_in_685 = io_in_685;
  assign fc1_io_in_686 = io_in_686;
  assign fc1_io_in_687 = io_in_687;
  assign fc1_io_in_688 = io_in_688;
  assign fc1_io_in_689 = io_in_689;
  assign fc1_io_in_690 = io_in_690;
  assign fc1_io_in_691 = io_in_691;
  assign fc1_io_in_692 = io_in_692;
  assign fc1_io_in_693 = io_in_693;
  assign fc1_io_in_694 = io_in_694;
  assign fc1_io_in_695 = io_in_695;
  assign fc1_io_in_696 = io_in_696;
  assign fc1_io_in_697 = io_in_697;
  assign fc1_io_in_698 = io_in_698;
  assign fc1_io_in_699 = io_in_699;
  assign fc1_io_in_702 = io_in_702;
  assign fc1_io_in_703 = io_in_703;
  assign fc1_io_in_704 = io_in_704;
  assign fc1_io_in_705 = io_in_705;
  assign fc1_io_in_706 = io_in_706;
  assign fc1_io_in_707 = io_in_707;
  assign fc1_io_in_708 = io_in_708;
  assign fc1_io_in_709 = io_in_709;
  assign fc1_io_in_710 = io_in_710;
  assign fc1_io_in_711 = io_in_711;
  assign fc1_io_in_712 = io_in_712;
  assign fc1_io_in_713 = io_in_713;
  assign fc1_io_in_714 = io_in_714;
  assign fc1_io_in_715 = io_in_715;
  assign fc1_io_in_716 = io_in_716;
  assign fc1_io_in_717 = io_in_717;
  assign fc1_io_in_718 = io_in_718;
  assign fc1_io_in_719 = io_in_719;
  assign fc1_io_in_720 = io_in_720;
  assign fc1_io_in_721 = io_in_721;
  assign fc1_io_in_722 = io_in_722;
  assign fc1_io_in_723 = io_in_723;
  assign fc1_io_in_724 = io_in_724;
  assign fc1_io_in_725 = io_in_725;
  assign fc1_io_in_726 = io_in_726;
  assign fc1_io_in_728 = io_in_728;
  assign fc1_io_in_729 = io_in_729;
  assign fc1_io_in_731 = io_in_731;
  assign fc1_io_in_732 = io_in_732;
  assign fc1_io_in_733 = io_in_733;
  assign fc1_io_in_734 = io_in_734;
  assign fc1_io_in_735 = io_in_735;
  assign fc1_io_in_736 = io_in_736;
  assign fc1_io_in_737 = io_in_737;
  assign fc1_io_in_738 = io_in_738;
  assign fc1_io_in_739 = io_in_739;
  assign fc1_io_in_740 = io_in_740;
  assign fc1_io_in_741 = io_in_741;
  assign fc1_io_in_742 = io_in_742;
  assign fc1_io_in_743 = io_in_743;
  assign fc1_io_in_744 = io_in_744;
  assign fc1_io_in_745 = io_in_745;
  assign fc1_io_in_746 = io_in_746;
  assign fc1_io_in_747 = io_in_747;
  assign fc1_io_in_748 = io_in_748;
  assign fc1_io_in_749 = io_in_749;
  assign fc1_io_in_750 = io_in_750;
  assign fc1_io_in_751 = io_in_751;
  assign fc1_io_in_752 = io_in_752;
  assign fc1_io_in_753 = io_in_753;
  assign fc1_io_in_756 = io_in_756;
  assign fc1_io_in_758 = io_in_758;
  assign fc1_io_in_760 = io_in_760;
  assign fc1_io_in_761 = io_in_761;
  assign fc1_io_in_762 = io_in_762;
  assign fc1_io_in_763 = io_in_763;
  assign fc1_io_in_764 = io_in_764;
  assign fc1_io_in_765 = io_in_765;
  assign fc1_io_in_766 = io_in_766;
  assign fc1_io_in_767 = io_in_767;
  assign fc1_io_in_768 = io_in_768;
  assign fc1_io_in_769 = io_in_769;
  assign fc1_io_in_770 = io_in_770;
  assign fc1_io_in_771 = io_in_771;
  assign fc1_io_in_772 = io_in_772;
  assign fc1_io_in_773 = io_in_773;
  assign fc1_io_in_774 = io_in_774;
  assign fc1_io_in_775 = io_in_775;
  assign fc1_io_in_776 = io_in_776;
  assign fc1_io_in_777 = io_in_777;
  assign fc1_io_in_778 = io_in_778;
  assign fc1_io_in_779 = io_in_779;
  assign fc1_io_in_780 = io_in_780;
  assign bn_bi1_io_in_0 = fc1_io_out_0;
  assign bn_bi1_io_in_1 = fc1_io_out_1;
  assign bn_bi1_io_in_2 = fc1_io_out_2;
  assign bn_bi1_io_in_3 = fc1_io_out_3;
  assign bn_bi1_io_in_4 = fc1_io_out_4;
  assign bn_bi1_io_in_5 = fc1_io_out_5;
  assign bn_bi1_io_in_6 = fc1_io_out_6;
  assign bn_bi1_io_in_7 = fc1_io_out_7;
  assign bn_bi1_io_in_8 = fc1_io_out_8;
  assign bn_bi1_io_in_9 = fc1_io_out_9;
  assign bn_bi1_io_in_10 = fc1_io_out_10;
  assign bn_bi1_io_in_11 = fc1_io_out_11;
  assign bn_bi1_io_in_12 = fc1_io_out_12;
  assign bn_bi1_io_in_13 = fc1_io_out_13;
  assign bn_bi1_io_in_14 = fc1_io_out_14;
  assign bn_bi1_io_in_15 = fc1_io_out_15;
  assign _GEN_0 = bn_bi1_io_out_0[1:0];
  assign fc2_io_in_0 = $signed(_GEN_0);
  assign _GEN_1 = bn_bi1_io_out_1[1:0];
  assign fc2_io_in_1 = $signed(_GEN_1);
  assign _GEN_2 = bn_bi1_io_out_2[1:0];
  assign fc2_io_in_2 = $signed(_GEN_2);
  assign _GEN_3 = bn_bi1_io_out_3[1:0];
  assign fc2_io_in_3 = $signed(_GEN_3);
  assign _GEN_4 = bn_bi1_io_out_4[1:0];
  assign fc2_io_in_4 = $signed(_GEN_4);
  assign _GEN_5 = bn_bi1_io_out_5[1:0];
  assign fc2_io_in_5 = $signed(_GEN_5);
  assign _GEN_6 = bn_bi1_io_out_6[1:0];
  assign fc2_io_in_6 = $signed(_GEN_6);
  assign _GEN_7 = bn_bi1_io_out_7[1:0];
  assign fc2_io_in_7 = $signed(_GEN_7);
  assign _GEN_8 = bn_bi1_io_out_8[1:0];
  assign fc2_io_in_8 = $signed(_GEN_8);
  assign _GEN_9 = bn_bi1_io_out_9[1:0];
  assign fc2_io_in_9 = $signed(_GEN_9);
  assign _GEN_10 = bn_bi1_io_out_10[1:0];
  assign fc2_io_in_10 = $signed(_GEN_10);
  assign _GEN_11 = bn_bi1_io_out_11[1:0];
  assign fc2_io_in_11 = $signed(_GEN_11);
  assign _GEN_12 = bn_bi1_io_out_12[1:0];
  assign fc2_io_in_12 = $signed(_GEN_12);
  assign _GEN_13 = bn_bi1_io_out_13[1:0];
  assign fc2_io_in_13 = $signed(_GEN_13);
  assign _GEN_14 = bn_bi1_io_out_14[1:0];
  assign fc2_io_in_14 = $signed(_GEN_14);
  assign _GEN_15 = bn_bi1_io_out_15[1:0];
  assign fc2_io_in_15 = $signed(_GEN_15);
  assign bn_bi2_io_in_0 = fc2_io_out_0;
  assign bn_bi2_io_in_1 = fc2_io_out_1;
  assign bn_bi2_io_in_2 = fc2_io_out_2;
  assign bn_bi2_io_in_3 = fc2_io_out_3;
  assign bn_bi2_io_in_4 = fc2_io_out_4;
  assign bn_bi2_io_in_5 = fc2_io_out_5;
  assign bn_bi2_io_in_6 = fc2_io_out_6;
  assign bn_bi2_io_in_7 = fc2_io_out_7;
  assign bn_bi2_io_in_8 = fc2_io_out_8;
  assign bn_bi2_io_in_9 = fc2_io_out_9;
  assign bn_bi2_io_in_10 = fc2_io_out_10;
  assign bn_bi2_io_in_11 = fc2_io_out_11;
  assign bn_bi2_io_in_12 = fc2_io_out_12;
  assign bn_bi2_io_in_13 = fc2_io_out_13;
  assign bn_bi2_io_in_14 = fc2_io_out_14;
  assign bn_bi2_io_in_15 = fc2_io_out_15;
  assign _GEN_16 = bn_bi2_io_out_0[1:0];
  assign fc3_io_in_0 = $signed(_GEN_16);
  assign _GEN_17 = bn_bi2_io_out_1[1:0];
  assign fc3_io_in_1 = $signed(_GEN_17);
  assign _GEN_18 = bn_bi2_io_out_2[1:0];
  assign fc3_io_in_2 = $signed(_GEN_18);
  assign _GEN_19 = bn_bi2_io_out_3[1:0];
  assign fc3_io_in_3 = $signed(_GEN_19);
  assign _GEN_20 = bn_bi2_io_out_4[1:0];
  assign fc3_io_in_4 = $signed(_GEN_20);
  assign _GEN_21 = bn_bi2_io_out_5[1:0];
  assign fc3_io_in_5 = $signed(_GEN_21);
  assign _GEN_22 = bn_bi2_io_out_6[1:0];
  assign fc3_io_in_6 = $signed(_GEN_22);
  assign _GEN_23 = bn_bi2_io_out_7[1:0];
  assign fc3_io_in_7 = $signed(_GEN_23);
  assign _GEN_24 = bn_bi2_io_out_8[1:0];
  assign fc3_io_in_8 = $signed(_GEN_24);
  assign _GEN_25 = bn_bi2_io_out_9[1:0];
  assign fc3_io_in_9 = $signed(_GEN_25);
  assign _GEN_26 = bn_bi2_io_out_10[1:0];
  assign fc3_io_in_10 = $signed(_GEN_26);
  assign _GEN_27 = bn_bi2_io_out_11[1:0];
  assign fc3_io_in_11 = $signed(_GEN_27);
  assign _GEN_28 = bn_bi2_io_out_12[1:0];
  assign fc3_io_in_12 = $signed(_GEN_28);
  assign _GEN_29 = bn_bi2_io_out_13[1:0];
  assign fc3_io_in_13 = $signed(_GEN_29);
  assign _GEN_30 = bn_bi2_io_out_14[1:0];
  assign fc3_io_in_14 = $signed(_GEN_30);
  assign _GEN_31 = bn_bi2_io_out_15[1:0];
  assign fc3_io_in_15 = $signed(_GEN_31);
  assign bn3_io_in_0 = fc3_io_out_0;
  assign bn3_io_in_1 = fc3_io_out_1;
  assign bn3_io_in_2 = fc3_io_out_2;
  assign bn3_io_in_3 = fc3_io_out_3;
  assign bn3_io_in_4 = fc3_io_out_4;
  assign bn3_io_in_5 = fc3_io_out_5;
  assign bn3_io_in_6 = fc3_io_out_6;
  assign bn3_io_in_7 = fc3_io_out_7;
  assign bn3_io_in_8 = fc3_io_out_8;
  assign bn3_io_in_9 = fc3_io_out_9;
endmodule
