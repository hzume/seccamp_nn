`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module ShifBatchNorm( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [10:0] io_in_0, // @[:@6.4]
  input  [10:0] io_in_1, // @[:@6.4]
  input  [10:0] io_in_2, // @[:@6.4]
  input  [10:0] io_in_3, // @[:@6.4]
  input  [10:0] io_in_4, // @[:@6.4]
  input  [10:0] io_in_5, // @[:@6.4]
  input  [10:0] io_in_6, // @[:@6.4]
  input  [10:0] io_in_7, // @[:@6.4]
  input  [10:0] io_in_8, // @[:@6.4]
  input  [10:0] io_in_9, // @[:@6.4]
  input  [10:0] io_in_10, // @[:@6.4]
  input  [10:0] io_in_11, // @[:@6.4]
  input  [10:0] io_in_12, // @[:@6.4]
  input  [10:0] io_in_13, // @[:@6.4]
  input  [10:0] io_in_14, // @[:@6.4]
  input  [10:0] io_in_15, // @[:@6.4]
  output [10:0] io_out_0, // @[:@6.4]
  output [10:0] io_out_1, // @[:@6.4]
  output [10:0] io_out_2, // @[:@6.4]
  output [10:0] io_out_3, // @[:@6.4]
  output [10:0] io_out_4, // @[:@6.4]
  output [10:0] io_out_5, // @[:@6.4]
  output [10:0] io_out_6, // @[:@6.4]
  output [10:0] io_out_7, // @[:@6.4]
  output [10:0] io_out_8, // @[:@6.4]
  output [10:0] io_out_9, // @[:@6.4]
  output [10:0] io_out_10, // @[:@6.4]
  output [10:0] io_out_11, // @[:@6.4]
  output [10:0] io_out_12, // @[:@6.4]
  output [10:0] io_out_13, // @[:@6.4]
  output [10:0] io_out_14, // @[:@6.4]
  output [10:0] io_out_15 // @[:@6.4]
);
  wire [11:0] _T_108; // @[Modules.scala 111:28:@11.4]
  wire [10:0] _T_109; // @[Modules.scala 111:28:@12.4]
  wire [10:0] c_x_0; // @[Modules.scala 111:28:@13.4]
  wire [25:0] _GEN_0; // @[Modules.scala 116:32:@15.4]
  wire [25:0] _T_112; // @[Modules.scala 116:32:@15.4]
  wire [10:0] _GEN_1; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_0; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_2; // @[Modules.scala 118:37:@17.4]
  wire [25:0] _T_114; // @[Modules.scala 118:37:@17.4]
  wire [10:0] _GEN_3; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_0; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_116; // @[Modules.scala 119:38:@19.4]
  wire [10:0] _T_117; // @[Modules.scala 119:38:@20.4]
  wire [10:0] _T_118; // @[Modules.scala 119:38:@21.4]
  wire [11:0] _T_120; // @[Modules.scala 111:28:@23.4]
  wire [10:0] _T_121; // @[Modules.scala 111:28:@24.4]
  wire [10:0] c_x_1; // @[Modules.scala 111:28:@25.4]
  wire [25:0] _GEN_4; // @[Modules.scala 116:32:@27.4]
  wire [25:0] _T_124; // @[Modules.scala 116:32:@27.4]
  wire [10:0] _GEN_5; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_1; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_6; // @[Modules.scala 118:37:@29.4]
  wire [25:0] _T_126; // @[Modules.scala 118:37:@29.4]
  wire [10:0] _GEN_7; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_1; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_128; // @[Modules.scala 119:38:@31.4]
  wire [10:0] _T_129; // @[Modules.scala 119:38:@32.4]
  wire [10:0] _T_130; // @[Modules.scala 119:38:@33.4]
  wire [11:0] _T_132; // @[Modules.scala 111:28:@35.4]
  wire [10:0] _T_133; // @[Modules.scala 111:28:@36.4]
  wire [10:0] c_x_2; // @[Modules.scala 111:28:@37.4]
  wire [25:0] _GEN_8; // @[Modules.scala 116:32:@39.4]
  wire [25:0] _T_136; // @[Modules.scala 116:32:@39.4]
  wire [10:0] _GEN_9; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_2; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_10; // @[Modules.scala 118:37:@41.4]
  wire [25:0] _T_138; // @[Modules.scala 118:37:@41.4]
  wire [10:0] _GEN_11; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_2; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_140; // @[Modules.scala 119:38:@43.4]
  wire [10:0] _T_141; // @[Modules.scala 119:38:@44.4]
  wire [10:0] _T_142; // @[Modules.scala 119:38:@45.4]
  wire [11:0] _T_144; // @[Modules.scala 111:28:@47.4]
  wire [10:0] _T_145; // @[Modules.scala 111:28:@48.4]
  wire [10:0] c_x_3; // @[Modules.scala 111:28:@49.4]
  wire [25:0] _GEN_12; // @[Modules.scala 116:32:@51.4]
  wire [25:0] _T_148; // @[Modules.scala 116:32:@51.4]
  wire [10:0] _GEN_13; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_3; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_14; // @[Modules.scala 118:37:@53.4]
  wire [25:0] _T_150; // @[Modules.scala 118:37:@53.4]
  wire [10:0] _GEN_15; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_3; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_152; // @[Modules.scala 119:38:@55.4]
  wire [10:0] _T_153; // @[Modules.scala 119:38:@56.4]
  wire [10:0] _T_154; // @[Modules.scala 119:38:@57.4]
  wire [11:0] _T_156; // @[Modules.scala 111:28:@59.4]
  wire [10:0] _T_157; // @[Modules.scala 111:28:@60.4]
  wire [10:0] c_x_4; // @[Modules.scala 111:28:@61.4]
  wire [25:0] _GEN_16; // @[Modules.scala 116:32:@63.4]
  wire [25:0] _T_160; // @[Modules.scala 116:32:@63.4]
  wire [10:0] _GEN_17; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_4; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_18; // @[Modules.scala 118:37:@65.4]
  wire [25:0] _T_162; // @[Modules.scala 118:37:@65.4]
  wire [10:0] _GEN_19; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_4; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_164; // @[Modules.scala 119:38:@67.4]
  wire [10:0] _T_165; // @[Modules.scala 119:38:@68.4]
  wire [10:0] _T_166; // @[Modules.scala 119:38:@69.4]
  wire [11:0] _T_168; // @[Modules.scala 111:28:@71.4]
  wire [10:0] _T_169; // @[Modules.scala 111:28:@72.4]
  wire [10:0] c_x_5; // @[Modules.scala 111:28:@73.4]
  wire [25:0] _GEN_20; // @[Modules.scala 116:32:@75.4]
  wire [25:0] _T_172; // @[Modules.scala 116:32:@75.4]
  wire [10:0] _GEN_21; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_5; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_22; // @[Modules.scala 118:37:@77.4]
  wire [25:0] _T_174; // @[Modules.scala 118:37:@77.4]
  wire [10:0] _GEN_23; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_5; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_176; // @[Modules.scala 119:38:@79.4]
  wire [10:0] _T_177; // @[Modules.scala 119:38:@80.4]
  wire [10:0] _T_178; // @[Modules.scala 119:38:@81.4]
  wire [11:0] _T_180; // @[Modules.scala 111:28:@83.4]
  wire [10:0] _T_181; // @[Modules.scala 111:28:@84.4]
  wire [10:0] c_x_6; // @[Modules.scala 111:28:@85.4]
  wire [25:0] _GEN_24; // @[Modules.scala 116:32:@87.4]
  wire [25:0] _T_184; // @[Modules.scala 116:32:@87.4]
  wire [10:0] _GEN_25; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_6; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_26; // @[Modules.scala 118:37:@89.4]
  wire [25:0] _T_186; // @[Modules.scala 118:37:@89.4]
  wire [10:0] _GEN_27; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_6; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_188; // @[Modules.scala 119:38:@91.4]
  wire [10:0] _T_189; // @[Modules.scala 119:38:@92.4]
  wire [10:0] _T_190; // @[Modules.scala 119:38:@93.4]
  wire [11:0] _T_192; // @[Modules.scala 111:28:@95.4]
  wire [10:0] _T_193; // @[Modules.scala 111:28:@96.4]
  wire [10:0] c_x_7; // @[Modules.scala 111:28:@97.4]
  wire [25:0] _GEN_28; // @[Modules.scala 116:32:@99.4]
  wire [25:0] _T_196; // @[Modules.scala 116:32:@99.4]
  wire [10:0] _GEN_29; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_7; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_30; // @[Modules.scala 118:37:@101.4]
  wire [25:0] _T_198; // @[Modules.scala 118:37:@101.4]
  wire [10:0] _GEN_31; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_7; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_200; // @[Modules.scala 119:38:@103.4]
  wire [10:0] _T_201; // @[Modules.scala 119:38:@104.4]
  wire [10:0] _T_202; // @[Modules.scala 119:38:@105.4]
  wire [11:0] _T_204; // @[Modules.scala 111:28:@107.4]
  wire [10:0] _T_205; // @[Modules.scala 111:28:@108.4]
  wire [10:0] c_x_8; // @[Modules.scala 111:28:@109.4]
  wire [25:0] _GEN_32; // @[Modules.scala 116:32:@111.4]
  wire [25:0] _T_208; // @[Modules.scala 116:32:@111.4]
  wire [10:0] _GEN_33; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_8; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_34; // @[Modules.scala 118:37:@113.4]
  wire [25:0] _T_210; // @[Modules.scala 118:37:@113.4]
  wire [10:0] _GEN_35; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_8; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_212; // @[Modules.scala 119:38:@115.4]
  wire [10:0] _T_213; // @[Modules.scala 119:38:@116.4]
  wire [10:0] _T_214; // @[Modules.scala 119:38:@117.4]
  wire [11:0] _T_216; // @[Modules.scala 111:28:@119.4]
  wire [10:0] _T_217; // @[Modules.scala 111:28:@120.4]
  wire [10:0] c_x_9; // @[Modules.scala 111:28:@121.4]
  wire [25:0] _GEN_36; // @[Modules.scala 116:32:@123.4]
  wire [25:0] _T_220; // @[Modules.scala 116:32:@123.4]
  wire [10:0] _GEN_37; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_9; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_38; // @[Modules.scala 118:37:@125.4]
  wire [25:0] _T_222; // @[Modules.scala 118:37:@125.4]
  wire [10:0] _GEN_39; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_9; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_224; // @[Modules.scala 119:38:@127.4]
  wire [10:0] _T_225; // @[Modules.scala 119:38:@128.4]
  wire [10:0] _T_226; // @[Modules.scala 119:38:@129.4]
  wire [11:0] _T_228; // @[Modules.scala 111:28:@131.4]
  wire [10:0] _T_229; // @[Modules.scala 111:28:@132.4]
  wire [10:0] c_x_10; // @[Modules.scala 111:28:@133.4]
  wire [25:0] _GEN_40; // @[Modules.scala 116:32:@135.4]
  wire [25:0] _T_232; // @[Modules.scala 116:32:@135.4]
  wire [10:0] _GEN_41; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_10; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_42; // @[Modules.scala 118:37:@137.4]
  wire [25:0] _T_234; // @[Modules.scala 118:37:@137.4]
  wire [10:0] _GEN_43; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_10; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_236; // @[Modules.scala 119:38:@139.4]
  wire [10:0] _T_237; // @[Modules.scala 119:38:@140.4]
  wire [10:0] _T_238; // @[Modules.scala 119:38:@141.4]
  wire [11:0] _T_240; // @[Modules.scala 111:28:@143.4]
  wire [10:0] _T_241; // @[Modules.scala 111:28:@144.4]
  wire [10:0] c_x_11; // @[Modules.scala 111:28:@145.4]
  wire [25:0] _GEN_44; // @[Modules.scala 116:32:@147.4]
  wire [25:0] _T_244; // @[Modules.scala 116:32:@147.4]
  wire [10:0] _GEN_45; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_11; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_46; // @[Modules.scala 118:37:@149.4]
  wire [25:0] _T_246; // @[Modules.scala 118:37:@149.4]
  wire [10:0] _GEN_47; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_11; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_248; // @[Modules.scala 119:38:@151.4]
  wire [10:0] _T_249; // @[Modules.scala 119:38:@152.4]
  wire [10:0] _T_250; // @[Modules.scala 119:38:@153.4]
  wire [11:0] _T_252; // @[Modules.scala 111:28:@155.4]
  wire [10:0] _T_253; // @[Modules.scala 111:28:@156.4]
  wire [10:0] c_x_12; // @[Modules.scala 111:28:@157.4]
  wire [25:0] _GEN_48; // @[Modules.scala 116:32:@159.4]
  wire [25:0] _T_256; // @[Modules.scala 116:32:@159.4]
  wire [10:0] _GEN_49; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_12; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_50; // @[Modules.scala 118:37:@161.4]
  wire [25:0] _T_258; // @[Modules.scala 118:37:@161.4]
  wire [10:0] _GEN_51; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_12; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_260; // @[Modules.scala 119:38:@163.4]
  wire [10:0] _T_261; // @[Modules.scala 119:38:@164.4]
  wire [10:0] _T_262; // @[Modules.scala 119:38:@165.4]
  wire [11:0] _T_264; // @[Modules.scala 111:28:@167.4]
  wire [10:0] _T_265; // @[Modules.scala 111:28:@168.4]
  wire [10:0] c_x_13; // @[Modules.scala 111:28:@169.4]
  wire [25:0] _GEN_52; // @[Modules.scala 116:32:@171.4]
  wire [25:0] _T_268; // @[Modules.scala 116:32:@171.4]
  wire [10:0] _GEN_53; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_13; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_54; // @[Modules.scala 118:37:@173.4]
  wire [25:0] _T_270; // @[Modules.scala 118:37:@173.4]
  wire [10:0] _GEN_55; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_13; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_272; // @[Modules.scala 119:38:@175.4]
  wire [10:0] _T_273; // @[Modules.scala 119:38:@176.4]
  wire [10:0] _T_274; // @[Modules.scala 119:38:@177.4]
  wire [11:0] _T_276; // @[Modules.scala 111:28:@179.4]
  wire [10:0] _T_277; // @[Modules.scala 111:28:@180.4]
  wire [10:0] c_x_14; // @[Modules.scala 111:28:@181.4]
  wire [25:0] _GEN_56; // @[Modules.scala 116:32:@183.4]
  wire [25:0] _T_280; // @[Modules.scala 116:32:@183.4]
  wire [10:0] _GEN_57; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_14; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_58; // @[Modules.scala 118:37:@185.4]
  wire [25:0] _T_282; // @[Modules.scala 118:37:@185.4]
  wire [10:0] _GEN_59; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_14; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_284; // @[Modules.scala 119:38:@187.4]
  wire [10:0] _T_285; // @[Modules.scala 119:38:@188.4]
  wire [10:0] _T_286; // @[Modules.scala 119:38:@189.4]
  wire [11:0] _T_288; // @[Modules.scala 111:28:@191.4]
  wire [10:0] _T_289; // @[Modules.scala 111:28:@192.4]
  wire [10:0] c_x_15; // @[Modules.scala 111:28:@193.4]
  wire [25:0] _GEN_60; // @[Modules.scala 116:32:@195.4]
  wire [25:0] _T_292; // @[Modules.scala 116:32:@195.4]
  wire [10:0] _GEN_61; // @[Modules.scala 108:21:@9.4]
  wire [10:0] x_hat_15; // @[Modules.scala 108:21:@9.4]
  wire [25:0] _GEN_62; // @[Modules.scala 118:37:@197.4]
  wire [25:0] _T_294; // @[Modules.scala 118:37:@197.4]
  wire [10:0] _GEN_63; // @[Modules.scala 109:28:@10.4]
  wire [10:0] normed_x_hat_15; // @[Modules.scala 109:28:@10.4]
  wire [11:0] _T_296; // @[Modules.scala 119:38:@199.4]
  wire [10:0] _T_297; // @[Modules.scala 119:38:@200.4]
  wire [10:0] _T_298; // @[Modules.scala 119:38:@201.4]
  assign _T_108 = $signed(io_in_0) - $signed(11'sh49); // @[Modules.scala 111:28:@11.4]
  assign _T_109 = _T_108[10:0]; // @[Modules.scala 111:28:@12.4]
  assign c_x_0 = $signed(_T_109); // @[Modules.scala 111:28:@13.4]
  assign _GEN_0 = {{15{c_x_0[10]}},c_x_0}; // @[Modules.scala 116:32:@15.4]
  assign _T_112 = $signed(_GEN_0) << 4'h4; // @[Modules.scala 116:32:@15.4]
  assign _GEN_1 = _T_112[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_0 = $signed(_GEN_1); // @[Modules.scala 108:21:@9.4]
  assign _GEN_2 = {{15{x_hat_0[10]}},x_hat_0}; // @[Modules.scala 118:37:@17.4]
  assign _T_114 = $signed(_GEN_2) << 4'h2; // @[Modules.scala 118:37:@17.4]
  assign _GEN_3 = _T_114[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_0 = $signed(_GEN_3); // @[Modules.scala 109:28:@10.4]
  assign _T_116 = $signed(normed_x_hat_0) + $signed(-11'shf); // @[Modules.scala 119:38:@19.4]
  assign _T_117 = _T_116[10:0]; // @[Modules.scala 119:38:@20.4]
  assign _T_118 = $signed(_T_117); // @[Modules.scala 119:38:@21.4]
  assign _T_120 = $signed(io_in_1) - $signed(-11'sh2f); // @[Modules.scala 111:28:@23.4]
  assign _T_121 = _T_120[10:0]; // @[Modules.scala 111:28:@24.4]
  assign c_x_1 = $signed(_T_121); // @[Modules.scala 111:28:@25.4]
  assign _GEN_4 = {{15{c_x_1[10]}},c_x_1}; // @[Modules.scala 116:32:@27.4]
  assign _T_124 = $signed(_GEN_4) << 4'h4; // @[Modules.scala 116:32:@27.4]
  assign _GEN_5 = _T_124[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_1 = $signed(_GEN_5); // @[Modules.scala 108:21:@9.4]
  assign _GEN_6 = {{15{x_hat_1[10]}},x_hat_1}; // @[Modules.scala 118:37:@29.4]
  assign _T_126 = $signed(_GEN_6) << 4'h2; // @[Modules.scala 118:37:@29.4]
  assign _GEN_7 = _T_126[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_1 = $signed(_GEN_7); // @[Modules.scala 109:28:@10.4]
  assign _T_128 = $signed(normed_x_hat_1) + $signed(-11'sh5); // @[Modules.scala 119:38:@31.4]
  assign _T_129 = _T_128[10:0]; // @[Modules.scala 119:38:@32.4]
  assign _T_130 = $signed(_T_129); // @[Modules.scala 119:38:@33.4]
  assign _T_132 = $signed(io_in_2) - $signed(11'sh4a); // @[Modules.scala 111:28:@35.4]
  assign _T_133 = _T_132[10:0]; // @[Modules.scala 111:28:@36.4]
  assign c_x_2 = $signed(_T_133); // @[Modules.scala 111:28:@37.4]
  assign _GEN_8 = {{15{c_x_2[10]}},c_x_2}; // @[Modules.scala 116:32:@39.4]
  assign _T_136 = $signed(_GEN_8) << 4'h4; // @[Modules.scala 116:32:@39.4]
  assign _GEN_9 = _T_136[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_2 = $signed(_GEN_9); // @[Modules.scala 108:21:@9.4]
  assign _GEN_10 = {{15{x_hat_2[10]}},x_hat_2}; // @[Modules.scala 118:37:@41.4]
  assign _T_138 = $signed(_GEN_10) << 4'h2; // @[Modules.scala 118:37:@41.4]
  assign _GEN_11 = _T_138[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_2 = $signed(_GEN_11); // @[Modules.scala 109:28:@10.4]
  assign _T_140 = $signed(normed_x_hat_2) + $signed(-11'sh2); // @[Modules.scala 119:38:@43.4]
  assign _T_141 = _T_140[10:0]; // @[Modules.scala 119:38:@44.4]
  assign _T_142 = $signed(_T_141); // @[Modules.scala 119:38:@45.4]
  assign _T_144 = $signed(io_in_3) - $signed(-11'sh90); // @[Modules.scala 111:28:@47.4]
  assign _T_145 = _T_144[10:0]; // @[Modules.scala 111:28:@48.4]
  assign c_x_3 = $signed(_T_145); // @[Modules.scala 111:28:@49.4]
  assign _GEN_12 = {{15{c_x_3[10]}},c_x_3}; // @[Modules.scala 116:32:@51.4]
  assign _T_148 = $signed(_GEN_12) << 4'h4; // @[Modules.scala 116:32:@51.4]
  assign _GEN_13 = _T_148[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_3 = $signed(_GEN_13); // @[Modules.scala 108:21:@9.4]
  assign _GEN_14 = {{15{x_hat_3[10]}},x_hat_3}; // @[Modules.scala 118:37:@53.4]
  assign _T_150 = $signed(_GEN_14) << 4'h2; // @[Modules.scala 118:37:@53.4]
  assign _GEN_15 = _T_150[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_3 = $signed(_GEN_15); // @[Modules.scala 109:28:@10.4]
  assign _T_152 = $signed(normed_x_hat_3) + $signed(11'sh0); // @[Modules.scala 119:38:@55.4]
  assign _T_153 = _T_152[10:0]; // @[Modules.scala 119:38:@56.4]
  assign _T_154 = $signed(_T_153); // @[Modules.scala 119:38:@57.4]
  assign _T_156 = $signed(io_in_4) - $signed(-11'shc); // @[Modules.scala 111:28:@59.4]
  assign _T_157 = _T_156[10:0]; // @[Modules.scala 111:28:@60.4]
  assign c_x_4 = $signed(_T_157); // @[Modules.scala 111:28:@61.4]
  assign _GEN_16 = {{15{c_x_4[10]}},c_x_4}; // @[Modules.scala 116:32:@63.4]
  assign _T_160 = $signed(_GEN_16) << 4'h4; // @[Modules.scala 116:32:@63.4]
  assign _GEN_17 = _T_160[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_4 = $signed(_GEN_17); // @[Modules.scala 108:21:@9.4]
  assign _GEN_18 = {{15{x_hat_4[10]}},x_hat_4}; // @[Modules.scala 118:37:@65.4]
  assign _T_162 = $signed(_GEN_18) << 4'h2; // @[Modules.scala 118:37:@65.4]
  assign _GEN_19 = _T_162[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_4 = $signed(_GEN_19); // @[Modules.scala 109:28:@10.4]
  assign _T_164 = $signed(normed_x_hat_4) + $signed(11'sh11); // @[Modules.scala 119:38:@67.4]
  assign _T_165 = _T_164[10:0]; // @[Modules.scala 119:38:@68.4]
  assign _T_166 = $signed(_T_165); // @[Modules.scala 119:38:@69.4]
  assign _T_168 = $signed(io_in_5) - $signed(11'shc); // @[Modules.scala 111:28:@71.4]
  assign _T_169 = _T_168[10:0]; // @[Modules.scala 111:28:@72.4]
  assign c_x_5 = $signed(_T_169); // @[Modules.scala 111:28:@73.4]
  assign _GEN_20 = {{15{c_x_5[10]}},c_x_5}; // @[Modules.scala 116:32:@75.4]
  assign _T_172 = $signed(_GEN_20) << 4'h4; // @[Modules.scala 116:32:@75.4]
  assign _GEN_21 = _T_172[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_5 = $signed(_GEN_21); // @[Modules.scala 108:21:@9.4]
  assign _GEN_22 = {{15{x_hat_5[10]}},x_hat_5}; // @[Modules.scala 118:37:@77.4]
  assign _T_174 = $signed(_GEN_22) << 4'h2; // @[Modules.scala 118:37:@77.4]
  assign _GEN_23 = _T_174[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_5 = $signed(_GEN_23); // @[Modules.scala 109:28:@10.4]
  assign _T_176 = $signed(normed_x_hat_5) + $signed(11'sh3); // @[Modules.scala 119:38:@79.4]
  assign _T_177 = _T_176[10:0]; // @[Modules.scala 119:38:@80.4]
  assign _T_178 = $signed(_T_177); // @[Modules.scala 119:38:@81.4]
  assign _T_180 = $signed(io_in_6) - $signed(11'sh7d); // @[Modules.scala 111:28:@83.4]
  assign _T_181 = _T_180[10:0]; // @[Modules.scala 111:28:@84.4]
  assign c_x_6 = $signed(_T_181); // @[Modules.scala 111:28:@85.4]
  assign _GEN_24 = {{15{c_x_6[10]}},c_x_6}; // @[Modules.scala 116:32:@87.4]
  assign _T_184 = $signed(_GEN_24) << 4'h4; // @[Modules.scala 116:32:@87.4]
  assign _GEN_25 = _T_184[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_6 = $signed(_GEN_25); // @[Modules.scala 108:21:@9.4]
  assign _GEN_26 = {{15{x_hat_6[10]}},x_hat_6}; // @[Modules.scala 118:37:@89.4]
  assign _T_186 = $signed(_GEN_26) << 4'h2; // @[Modules.scala 118:37:@89.4]
  assign _GEN_27 = _T_186[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_6 = $signed(_GEN_27); // @[Modules.scala 109:28:@10.4]
  assign _T_188 = $signed(normed_x_hat_6) + $signed(-11'sh11); // @[Modules.scala 119:38:@91.4]
  assign _T_189 = _T_188[10:0]; // @[Modules.scala 119:38:@92.4]
  assign _T_190 = $signed(_T_189); // @[Modules.scala 119:38:@93.4]
  assign _T_192 = $signed(io_in_7) - $signed(11'sh3); // @[Modules.scala 111:28:@95.4]
  assign _T_193 = _T_192[10:0]; // @[Modules.scala 111:28:@96.4]
  assign c_x_7 = $signed(_T_193); // @[Modules.scala 111:28:@97.4]
  assign _GEN_28 = {{15{c_x_7[10]}},c_x_7}; // @[Modules.scala 116:32:@99.4]
  assign _T_196 = $signed(_GEN_28) << 4'h4; // @[Modules.scala 116:32:@99.4]
  assign _GEN_29 = _T_196[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_7 = $signed(_GEN_29); // @[Modules.scala 108:21:@9.4]
  assign _GEN_30 = {{15{x_hat_7[10]}},x_hat_7}; // @[Modules.scala 118:37:@101.4]
  assign _T_198 = $signed(_GEN_30) << 4'h1; // @[Modules.scala 118:37:@101.4]
  assign _GEN_31 = _T_198[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_7 = $signed(_GEN_31); // @[Modules.scala 109:28:@10.4]
  assign _T_200 = $signed(normed_x_hat_7) + $signed(11'sh1); // @[Modules.scala 119:38:@103.4]
  assign _T_201 = _T_200[10:0]; // @[Modules.scala 119:38:@104.4]
  assign _T_202 = $signed(_T_201); // @[Modules.scala 119:38:@105.4]
  assign _T_204 = $signed(io_in_8) - $signed(-11'sh5); // @[Modules.scala 111:28:@107.4]
  assign _T_205 = _T_204[10:0]; // @[Modules.scala 111:28:@108.4]
  assign c_x_8 = $signed(_T_205); // @[Modules.scala 111:28:@109.4]
  assign _GEN_32 = {{15{c_x_8[10]}},c_x_8}; // @[Modules.scala 116:32:@111.4]
  assign _T_208 = $signed(_GEN_32) << 4'h4; // @[Modules.scala 116:32:@111.4]
  assign _GEN_33 = _T_208[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_8 = $signed(_GEN_33); // @[Modules.scala 108:21:@9.4]
  assign _GEN_34 = {{15{x_hat_8[10]}},x_hat_8}; // @[Modules.scala 118:37:@113.4]
  assign _T_210 = $signed(_GEN_34) << 4'h2; // @[Modules.scala 118:37:@113.4]
  assign _GEN_35 = _T_210[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_8 = $signed(_GEN_35); // @[Modules.scala 109:28:@10.4]
  assign _T_212 = $signed(normed_x_hat_8) + $signed(-11'sh6); // @[Modules.scala 119:38:@115.4]
  assign _T_213 = _T_212[10:0]; // @[Modules.scala 119:38:@116.4]
  assign _T_214 = $signed(_T_213); // @[Modules.scala 119:38:@117.4]
  assign _T_216 = $signed(io_in_9) - $signed(-11'sh3d); // @[Modules.scala 111:28:@119.4]
  assign _T_217 = _T_216[10:0]; // @[Modules.scala 111:28:@120.4]
  assign c_x_9 = $signed(_T_217); // @[Modules.scala 111:28:@121.4]
  assign _GEN_36 = {{15{c_x_9[10]}},c_x_9}; // @[Modules.scala 116:32:@123.4]
  assign _T_220 = $signed(_GEN_36) << 4'h4; // @[Modules.scala 116:32:@123.4]
  assign _GEN_37 = _T_220[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_9 = $signed(_GEN_37); // @[Modules.scala 108:21:@9.4]
  assign _GEN_38 = {{15{x_hat_9[10]}},x_hat_9}; // @[Modules.scala 118:37:@125.4]
  assign _T_222 = $signed(_GEN_38) << 4'h1; // @[Modules.scala 118:37:@125.4]
  assign _GEN_39 = _T_222[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_9 = $signed(_GEN_39); // @[Modules.scala 109:28:@10.4]
  assign _T_224 = $signed(normed_x_hat_9) + $signed(11'sh1); // @[Modules.scala 119:38:@127.4]
  assign _T_225 = _T_224[10:0]; // @[Modules.scala 119:38:@128.4]
  assign _T_226 = $signed(_T_225); // @[Modules.scala 119:38:@129.4]
  assign _T_228 = $signed(io_in_10) - $signed(-11'shaf); // @[Modules.scala 111:28:@131.4]
  assign _T_229 = _T_228[10:0]; // @[Modules.scala 111:28:@132.4]
  assign c_x_10 = $signed(_T_229); // @[Modules.scala 111:28:@133.4]
  assign _GEN_40 = {{15{c_x_10[10]}},c_x_10}; // @[Modules.scala 116:32:@135.4]
  assign _T_232 = $signed(_GEN_40) << 4'h4; // @[Modules.scala 116:32:@135.4]
  assign _GEN_41 = _T_232[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_10 = $signed(_GEN_41); // @[Modules.scala 108:21:@9.4]
  assign _GEN_42 = {{15{x_hat_10[10]}},x_hat_10}; // @[Modules.scala 118:37:@137.4]
  assign _T_234 = $signed(_GEN_42) << 4'h2; // @[Modules.scala 118:37:@137.4]
  assign _GEN_43 = _T_234[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_10 = $signed(_GEN_43); // @[Modules.scala 109:28:@10.4]
  assign _T_236 = $signed(normed_x_hat_10) + $signed(-11'sh6); // @[Modules.scala 119:38:@139.4]
  assign _T_237 = _T_236[10:0]; // @[Modules.scala 119:38:@140.4]
  assign _T_238 = $signed(_T_237); // @[Modules.scala 119:38:@141.4]
  assign _T_240 = $signed(io_in_11) - $signed(11'sh75); // @[Modules.scala 111:28:@143.4]
  assign _T_241 = _T_240[10:0]; // @[Modules.scala 111:28:@144.4]
  assign c_x_11 = $signed(_T_241); // @[Modules.scala 111:28:@145.4]
  assign _GEN_44 = {{15{c_x_11[10]}},c_x_11}; // @[Modules.scala 116:32:@147.4]
  assign _T_244 = $signed(_GEN_44) << 4'h4; // @[Modules.scala 116:32:@147.4]
  assign _GEN_45 = _T_244[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_11 = $signed(_GEN_45); // @[Modules.scala 108:21:@9.4]
  assign _GEN_46 = {{15{x_hat_11[10]}},x_hat_11}; // @[Modules.scala 118:37:@149.4]
  assign _T_246 = $signed(_GEN_46) << 4'h1; // @[Modules.scala 118:37:@149.4]
  assign _GEN_47 = _T_246[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_11 = $signed(_GEN_47); // @[Modules.scala 109:28:@10.4]
  assign _T_248 = $signed(normed_x_hat_11) + $signed(-11'sh9); // @[Modules.scala 119:38:@151.4]
  assign _T_249 = _T_248[10:0]; // @[Modules.scala 119:38:@152.4]
  assign _T_250 = $signed(_T_249); // @[Modules.scala 119:38:@153.4]
  assign _T_252 = $signed(io_in_12) - $signed(-11'sh32); // @[Modules.scala 111:28:@155.4]
  assign _T_253 = _T_252[10:0]; // @[Modules.scala 111:28:@156.4]
  assign c_x_12 = $signed(_T_253); // @[Modules.scala 111:28:@157.4]
  assign _GEN_48 = {{15{c_x_12[10]}},c_x_12}; // @[Modules.scala 116:32:@159.4]
  assign _T_256 = $signed(_GEN_48) << 4'h4; // @[Modules.scala 116:32:@159.4]
  assign _GEN_49 = _T_256[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_12 = $signed(_GEN_49); // @[Modules.scala 108:21:@9.4]
  assign _GEN_50 = {{15{x_hat_12[10]}},x_hat_12}; // @[Modules.scala 118:37:@161.4]
  assign _T_258 = $signed(_GEN_50) << 4'h2; // @[Modules.scala 118:37:@161.4]
  assign _GEN_51 = _T_258[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_12 = $signed(_GEN_51); // @[Modules.scala 109:28:@10.4]
  assign _T_260 = $signed(normed_x_hat_12) + $signed(-11'sh9); // @[Modules.scala 119:38:@163.4]
  assign _T_261 = _T_260[10:0]; // @[Modules.scala 119:38:@164.4]
  assign _T_262 = $signed(_T_261); // @[Modules.scala 119:38:@165.4]
  assign _T_264 = $signed(io_in_13) - $signed(11'sh77); // @[Modules.scala 111:28:@167.4]
  assign _T_265 = _T_264[10:0]; // @[Modules.scala 111:28:@168.4]
  assign c_x_13 = $signed(_T_265); // @[Modules.scala 111:28:@169.4]
  assign _GEN_52 = {{15{c_x_13[10]}},c_x_13}; // @[Modules.scala 116:32:@171.4]
  assign _T_268 = $signed(_GEN_52) << 4'h4; // @[Modules.scala 116:32:@171.4]
  assign _GEN_53 = _T_268[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_13 = $signed(_GEN_53); // @[Modules.scala 108:21:@9.4]
  assign _GEN_54 = {{15{x_hat_13[10]}},x_hat_13}; // @[Modules.scala 118:37:@173.4]
  assign _T_270 = $signed(_GEN_54) << 4'h1; // @[Modules.scala 118:37:@173.4]
  assign _GEN_55 = _T_270[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_13 = $signed(_GEN_55); // @[Modules.scala 109:28:@10.4]
  assign _T_272 = $signed(normed_x_hat_13) + $signed(11'sh5); // @[Modules.scala 119:38:@175.4]
  assign _T_273 = _T_272[10:0]; // @[Modules.scala 119:38:@176.4]
  assign _T_274 = $signed(_T_273); // @[Modules.scala 119:38:@177.4]
  assign _T_276 = $signed(io_in_14) - $signed(11'sh19); // @[Modules.scala 111:28:@179.4]
  assign _T_277 = _T_276[10:0]; // @[Modules.scala 111:28:@180.4]
  assign c_x_14 = $signed(_T_277); // @[Modules.scala 111:28:@181.4]
  assign _GEN_56 = {{15{c_x_14[10]}},c_x_14}; // @[Modules.scala 116:32:@183.4]
  assign _T_280 = $signed(_GEN_56) << 4'h4; // @[Modules.scala 116:32:@183.4]
  assign _GEN_57 = _T_280[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_14 = $signed(_GEN_57); // @[Modules.scala 108:21:@9.4]
  assign _GEN_58 = {{15{x_hat_14[10]}},x_hat_14}; // @[Modules.scala 118:37:@185.4]
  assign _T_282 = $signed(_GEN_58) << 4'h2; // @[Modules.scala 118:37:@185.4]
  assign _GEN_59 = _T_282[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_14 = $signed(_GEN_59); // @[Modules.scala 109:28:@10.4]
  assign _T_284 = $signed(normed_x_hat_14) + $signed(11'sh7); // @[Modules.scala 119:38:@187.4]
  assign _T_285 = _T_284[10:0]; // @[Modules.scala 119:38:@188.4]
  assign _T_286 = $signed(_T_285); // @[Modules.scala 119:38:@189.4]
  assign _T_288 = $signed(io_in_15) - $signed(-11'sh64); // @[Modules.scala 111:28:@191.4]
  assign _T_289 = _T_288[10:0]; // @[Modules.scala 111:28:@192.4]
  assign c_x_15 = $signed(_T_289); // @[Modules.scala 111:28:@193.4]
  assign _GEN_60 = {{15{c_x_15[10]}},c_x_15}; // @[Modules.scala 116:32:@195.4]
  assign _T_292 = $signed(_GEN_60) << 4'h4; // @[Modules.scala 116:32:@195.4]
  assign _GEN_61 = _T_292[10:0]; // @[Modules.scala 108:21:@9.4]
  assign x_hat_15 = $signed(_GEN_61); // @[Modules.scala 108:21:@9.4]
  assign _GEN_62 = {{15{x_hat_15[10]}},x_hat_15}; // @[Modules.scala 118:37:@197.4]
  assign _T_294 = $signed(_GEN_62) << 4'h1; // @[Modules.scala 118:37:@197.4]
  assign _GEN_63 = _T_294[10:0]; // @[Modules.scala 109:28:@10.4]
  assign normed_x_hat_15 = $signed(_GEN_63); // @[Modules.scala 109:28:@10.4]
  assign _T_296 = $signed(normed_x_hat_15) + $signed(11'sh4); // @[Modules.scala 119:38:@199.4]
  assign _T_297 = _T_296[10:0]; // @[Modules.scala 119:38:@200.4]
  assign _T_298 = $signed(_T_297); // @[Modules.scala 119:38:@201.4]
  assign io_out_0 = _T_118;
  assign io_out_1 = _T_130;
  assign io_out_2 = _T_142;
  assign io_out_3 = _T_154;
  assign io_out_4 = _T_166;
  assign io_out_5 = _T_178;
  assign io_out_6 = _T_190;
  assign io_out_7 = _T_202;
  assign io_out_8 = _T_214;
  assign io_out_9 = _T_226;
  assign io_out_10 = _T_238;
  assign io_out_11 = _T_250;
  assign io_out_12 = _T_262;
  assign io_out_13 = _T_274;
  assign io_out_14 = _T_286;
  assign io_out_15 = _T_298;
endmodule
