`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Linear_p( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [4:0]  io_in_0, // @[:@6.4]
  input  [4:0]  io_in_1, // @[:@6.4]
  input  [4:0]  io_in_2, // @[:@6.4]
  input  [4:0]  io_in_3, // @[:@6.4]
  input  [4:0]  io_in_4, // @[:@6.4]
  input  [4:0]  io_in_5, // @[:@6.4]
  input  [4:0]  io_in_6, // @[:@6.4]
  input  [4:0]  io_in_7, // @[:@6.4]
  input  [4:0]  io_in_8, // @[:@6.4]
  input  [4:0]  io_in_9, // @[:@6.4]
  input  [4:0]  io_in_10, // @[:@6.4]
  input  [4:0]  io_in_11, // @[:@6.4]
  input  [4:0]  io_in_12, // @[:@6.4]
  input  [4:0]  io_in_13, // @[:@6.4]
  input  [4:0]  io_in_14, // @[:@6.4]
  input  [4:0]  io_in_15, // @[:@6.4]
  input  [4:0]  io_in_16, // @[:@6.4]
  input  [4:0]  io_in_17, // @[:@6.4]
  input  [4:0]  io_in_18, // @[:@6.4]
  input  [4:0]  io_in_19, // @[:@6.4]
  input  [4:0]  io_in_20, // @[:@6.4]
  input  [4:0]  io_in_21, // @[:@6.4]
  input  [4:0]  io_in_22, // @[:@6.4]
  input  [4:0]  io_in_23, // @[:@6.4]
  input  [4:0]  io_in_24, // @[:@6.4]
  input  [4:0]  io_in_25, // @[:@6.4]
  input  [4:0]  io_in_26, // @[:@6.4]
  input  [4:0]  io_in_27, // @[:@6.4]
  input  [4:0]  io_in_28, // @[:@6.4]
  input  [4:0]  io_in_29, // @[:@6.4]
  input  [4:0]  io_in_30, // @[:@6.4]
  input  [4:0]  io_in_31, // @[:@6.4]
  input  [4:0]  io_in_32, // @[:@6.4]
  input  [4:0]  io_in_33, // @[:@6.4]
  input  [4:0]  io_in_34, // @[:@6.4]
  input  [4:0]  io_in_35, // @[:@6.4]
  input  [4:0]  io_in_36, // @[:@6.4]
  input  [4:0]  io_in_37, // @[:@6.4]
  input  [4:0]  io_in_38, // @[:@6.4]
  input  [4:0]  io_in_39, // @[:@6.4]
  input  [4:0]  io_in_40, // @[:@6.4]
  input  [4:0]  io_in_41, // @[:@6.4]
  input  [4:0]  io_in_42, // @[:@6.4]
  input  [4:0]  io_in_43, // @[:@6.4]
  input  [4:0]  io_in_44, // @[:@6.4]
  input  [4:0]  io_in_45, // @[:@6.4]
  input  [4:0]  io_in_46, // @[:@6.4]
  input  [4:0]  io_in_47, // @[:@6.4]
  input  [4:0]  io_in_48, // @[:@6.4]
  input  [4:0]  io_in_49, // @[:@6.4]
  input  [4:0]  io_in_50, // @[:@6.4]
  input  [4:0]  io_in_51, // @[:@6.4]
  input  [4:0]  io_in_52, // @[:@6.4]
  input  [4:0]  io_in_53, // @[:@6.4]
  input  [4:0]  io_in_54, // @[:@6.4]
  input  [4:0]  io_in_55, // @[:@6.4]
  input  [4:0]  io_in_56, // @[:@6.4]
  input  [4:0]  io_in_57, // @[:@6.4]
  input  [4:0]  io_in_58, // @[:@6.4]
  input  [4:0]  io_in_59, // @[:@6.4]
  input  [4:0]  io_in_60, // @[:@6.4]
  input  [4:0]  io_in_61, // @[:@6.4]
  input  [4:0]  io_in_62, // @[:@6.4]
  input  [4:0]  io_in_63, // @[:@6.4]
  input  [4:0]  io_in_64, // @[:@6.4]
  input  [4:0]  io_in_65, // @[:@6.4]
  input  [4:0]  io_in_66, // @[:@6.4]
  input  [4:0]  io_in_67, // @[:@6.4]
  input  [4:0]  io_in_68, // @[:@6.4]
  input  [4:0]  io_in_69, // @[:@6.4]
  input  [4:0]  io_in_70, // @[:@6.4]
  input  [4:0]  io_in_71, // @[:@6.4]
  input  [4:0]  io_in_72, // @[:@6.4]
  input  [4:0]  io_in_73, // @[:@6.4]
  input  [4:0]  io_in_74, // @[:@6.4]
  input  [4:0]  io_in_75, // @[:@6.4]
  input  [4:0]  io_in_76, // @[:@6.4]
  input  [4:0]  io_in_77, // @[:@6.4]
  input  [4:0]  io_in_78, // @[:@6.4]
  input  [4:0]  io_in_79, // @[:@6.4]
  input  [4:0]  io_in_80, // @[:@6.4]
  input  [4:0]  io_in_81, // @[:@6.4]
  input  [4:0]  io_in_82, // @[:@6.4]
  input  [4:0]  io_in_83, // @[:@6.4]
  input  [4:0]  io_in_84, // @[:@6.4]
  input  [4:0]  io_in_85, // @[:@6.4]
  input  [4:0]  io_in_86, // @[:@6.4]
  input  [4:0]  io_in_87, // @[:@6.4]
  input  [4:0]  io_in_88, // @[:@6.4]
  input  [4:0]  io_in_89, // @[:@6.4]
  input  [4:0]  io_in_90, // @[:@6.4]
  input  [4:0]  io_in_91, // @[:@6.4]
  input  [4:0]  io_in_92, // @[:@6.4]
  input  [4:0]  io_in_93, // @[:@6.4]
  input  [4:0]  io_in_94, // @[:@6.4]
  input  [4:0]  io_in_95, // @[:@6.4]
  input  [4:0]  io_in_96, // @[:@6.4]
  input  [4:0]  io_in_97, // @[:@6.4]
  input  [4:0]  io_in_98, // @[:@6.4]
  input  [4:0]  io_in_99, // @[:@6.4]
  input  [4:0]  io_in_100, // @[:@6.4]
  input  [4:0]  io_in_101, // @[:@6.4]
  input  [4:0]  io_in_102, // @[:@6.4]
  input  [4:0]  io_in_103, // @[:@6.4]
  input  [4:0]  io_in_104, // @[:@6.4]
  input  [4:0]  io_in_105, // @[:@6.4]
  input  [4:0]  io_in_106, // @[:@6.4]
  input  [4:0]  io_in_107, // @[:@6.4]
  input  [4:0]  io_in_108, // @[:@6.4]
  input  [4:0]  io_in_109, // @[:@6.4]
  input  [4:0]  io_in_110, // @[:@6.4]
  input  [4:0]  io_in_111, // @[:@6.4]
  input  [4:0]  io_in_112, // @[:@6.4]
  input  [4:0]  io_in_113, // @[:@6.4]
  input  [4:0]  io_in_114, // @[:@6.4]
  input  [4:0]  io_in_115, // @[:@6.4]
  input  [4:0]  io_in_116, // @[:@6.4]
  input  [4:0]  io_in_117, // @[:@6.4]
  input  [4:0]  io_in_118, // @[:@6.4]
  input  [4:0]  io_in_119, // @[:@6.4]
  input  [4:0]  io_in_120, // @[:@6.4]
  input  [4:0]  io_in_121, // @[:@6.4]
  input  [4:0]  io_in_122, // @[:@6.4]
  input  [4:0]  io_in_123, // @[:@6.4]
  input  [4:0]  io_in_124, // @[:@6.4]
  input  [4:0]  io_in_125, // @[:@6.4]
  input  [4:0]  io_in_126, // @[:@6.4]
  input  [4:0]  io_in_127, // @[:@6.4]
  input  [4:0]  io_in_128, // @[:@6.4]
  input  [4:0]  io_in_129, // @[:@6.4]
  input  [4:0]  io_in_130, // @[:@6.4]
  input  [4:0]  io_in_131, // @[:@6.4]
  input  [4:0]  io_in_132, // @[:@6.4]
  input  [4:0]  io_in_133, // @[:@6.4]
  input  [4:0]  io_in_134, // @[:@6.4]
  input  [4:0]  io_in_135, // @[:@6.4]
  input  [4:0]  io_in_136, // @[:@6.4]
  input  [4:0]  io_in_137, // @[:@6.4]
  input  [4:0]  io_in_138, // @[:@6.4]
  input  [4:0]  io_in_139, // @[:@6.4]
  input  [4:0]  io_in_140, // @[:@6.4]
  input  [4:0]  io_in_141, // @[:@6.4]
  input  [4:0]  io_in_142, // @[:@6.4]
  input  [4:0]  io_in_143, // @[:@6.4]
  input  [4:0]  io_in_144, // @[:@6.4]
  input  [4:0]  io_in_145, // @[:@6.4]
  input  [4:0]  io_in_146, // @[:@6.4]
  input  [4:0]  io_in_147, // @[:@6.4]
  input  [4:0]  io_in_148, // @[:@6.4]
  input  [4:0]  io_in_149, // @[:@6.4]
  input  [4:0]  io_in_150, // @[:@6.4]
  input  [4:0]  io_in_151, // @[:@6.4]
  input  [4:0]  io_in_152, // @[:@6.4]
  input  [4:0]  io_in_153, // @[:@6.4]
  input  [4:0]  io_in_154, // @[:@6.4]
  input  [4:0]  io_in_155, // @[:@6.4]
  input  [4:0]  io_in_156, // @[:@6.4]
  input  [4:0]  io_in_157, // @[:@6.4]
  input  [4:0]  io_in_158, // @[:@6.4]
  input  [4:0]  io_in_159, // @[:@6.4]
  input  [4:0]  io_in_160, // @[:@6.4]
  input  [4:0]  io_in_161, // @[:@6.4]
  input  [4:0]  io_in_162, // @[:@6.4]
  input  [4:0]  io_in_163, // @[:@6.4]
  input  [4:0]  io_in_164, // @[:@6.4]
  input  [4:0]  io_in_165, // @[:@6.4]
  input  [4:0]  io_in_166, // @[:@6.4]
  input  [4:0]  io_in_167, // @[:@6.4]
  input  [4:0]  io_in_168, // @[:@6.4]
  input  [4:0]  io_in_169, // @[:@6.4]
  input  [4:0]  io_in_170, // @[:@6.4]
  input  [4:0]  io_in_171, // @[:@6.4]
  input  [4:0]  io_in_172, // @[:@6.4]
  input  [4:0]  io_in_173, // @[:@6.4]
  input  [4:0]  io_in_174, // @[:@6.4]
  input  [4:0]  io_in_175, // @[:@6.4]
  input  [4:0]  io_in_176, // @[:@6.4]
  input  [4:0]  io_in_177, // @[:@6.4]
  input  [4:0]  io_in_178, // @[:@6.4]
  input  [4:0]  io_in_179, // @[:@6.4]
  input  [4:0]  io_in_180, // @[:@6.4]
  input  [4:0]  io_in_181, // @[:@6.4]
  input  [4:0]  io_in_182, // @[:@6.4]
  input  [4:0]  io_in_183, // @[:@6.4]
  input  [4:0]  io_in_184, // @[:@6.4]
  input  [4:0]  io_in_185, // @[:@6.4]
  input  [4:0]  io_in_186, // @[:@6.4]
  input  [4:0]  io_in_187, // @[:@6.4]
  input  [4:0]  io_in_188, // @[:@6.4]
  input  [4:0]  io_in_189, // @[:@6.4]
  input  [4:0]  io_in_190, // @[:@6.4]
  input  [4:0]  io_in_191, // @[:@6.4]
  input  [4:0]  io_in_192, // @[:@6.4]
  input  [4:0]  io_in_193, // @[:@6.4]
  input  [4:0]  io_in_194, // @[:@6.4]
  input  [4:0]  io_in_195, // @[:@6.4]
  input  [4:0]  io_in_196, // @[:@6.4]
  input  [4:0]  io_in_197, // @[:@6.4]
  input  [4:0]  io_in_198, // @[:@6.4]
  input  [4:0]  io_in_199, // @[:@6.4]
  input  [4:0]  io_in_200, // @[:@6.4]
  input  [4:0]  io_in_201, // @[:@6.4]
  input  [4:0]  io_in_202, // @[:@6.4]
  input  [4:0]  io_in_203, // @[:@6.4]
  input  [4:0]  io_in_204, // @[:@6.4]
  input  [4:0]  io_in_205, // @[:@6.4]
  input  [4:0]  io_in_206, // @[:@6.4]
  input  [4:0]  io_in_207, // @[:@6.4]
  input  [4:0]  io_in_208, // @[:@6.4]
  input  [4:0]  io_in_209, // @[:@6.4]
  input  [4:0]  io_in_210, // @[:@6.4]
  input  [4:0]  io_in_211, // @[:@6.4]
  input  [4:0]  io_in_212, // @[:@6.4]
  input  [4:0]  io_in_213, // @[:@6.4]
  input  [4:0]  io_in_214, // @[:@6.4]
  input  [4:0]  io_in_215, // @[:@6.4]
  input  [4:0]  io_in_216, // @[:@6.4]
  input  [4:0]  io_in_217, // @[:@6.4]
  input  [4:0]  io_in_218, // @[:@6.4]
  input  [4:0]  io_in_219, // @[:@6.4]
  input  [4:0]  io_in_220, // @[:@6.4]
  input  [4:0]  io_in_221, // @[:@6.4]
  input  [4:0]  io_in_222, // @[:@6.4]
  input  [4:0]  io_in_223, // @[:@6.4]
  input  [4:0]  io_in_224, // @[:@6.4]
  input  [4:0]  io_in_225, // @[:@6.4]
  input  [4:0]  io_in_226, // @[:@6.4]
  input  [4:0]  io_in_227, // @[:@6.4]
  input  [4:0]  io_in_228, // @[:@6.4]
  input  [4:0]  io_in_229, // @[:@6.4]
  input  [4:0]  io_in_230, // @[:@6.4]
  input  [4:0]  io_in_231, // @[:@6.4]
  input  [4:0]  io_in_232, // @[:@6.4]
  input  [4:0]  io_in_233, // @[:@6.4]
  input  [4:0]  io_in_234, // @[:@6.4]
  input  [4:0]  io_in_235, // @[:@6.4]
  input  [4:0]  io_in_236, // @[:@6.4]
  input  [4:0]  io_in_237, // @[:@6.4]
  input  [4:0]  io_in_238, // @[:@6.4]
  input  [4:0]  io_in_239, // @[:@6.4]
  input  [4:0]  io_in_240, // @[:@6.4]
  input  [4:0]  io_in_241, // @[:@6.4]
  input  [4:0]  io_in_242, // @[:@6.4]
  input  [4:0]  io_in_243, // @[:@6.4]
  input  [4:0]  io_in_244, // @[:@6.4]
  input  [4:0]  io_in_245, // @[:@6.4]
  input  [4:0]  io_in_246, // @[:@6.4]
  input  [4:0]  io_in_247, // @[:@6.4]
  input  [4:0]  io_in_248, // @[:@6.4]
  input  [4:0]  io_in_249, // @[:@6.4]
  input  [4:0]  io_in_250, // @[:@6.4]
  input  [4:0]  io_in_251, // @[:@6.4]
  input  [4:0]  io_in_252, // @[:@6.4]
  input  [4:0]  io_in_253, // @[:@6.4]
  input  [4:0]  io_in_254, // @[:@6.4]
  input  [4:0]  io_in_255, // @[:@6.4]
  input  [4:0]  io_in_256, // @[:@6.4]
  input  [4:0]  io_in_257, // @[:@6.4]
  input  [4:0]  io_in_258, // @[:@6.4]
  input  [4:0]  io_in_259, // @[:@6.4]
  input  [4:0]  io_in_260, // @[:@6.4]
  input  [4:0]  io_in_261, // @[:@6.4]
  input  [4:0]  io_in_262, // @[:@6.4]
  input  [4:0]  io_in_263, // @[:@6.4]
  input  [4:0]  io_in_264, // @[:@6.4]
  input  [4:0]  io_in_265, // @[:@6.4]
  input  [4:0]  io_in_266, // @[:@6.4]
  input  [4:0]  io_in_267, // @[:@6.4]
  input  [4:0]  io_in_268, // @[:@6.4]
  input  [4:0]  io_in_269, // @[:@6.4]
  input  [4:0]  io_in_270, // @[:@6.4]
  input  [4:0]  io_in_271, // @[:@6.4]
  input  [4:0]  io_in_272, // @[:@6.4]
  input  [4:0]  io_in_273, // @[:@6.4]
  input  [4:0]  io_in_274, // @[:@6.4]
  input  [4:0]  io_in_275, // @[:@6.4]
  input  [4:0]  io_in_276, // @[:@6.4]
  input  [4:0]  io_in_277, // @[:@6.4]
  input  [4:0]  io_in_278, // @[:@6.4]
  input  [4:0]  io_in_279, // @[:@6.4]
  input  [4:0]  io_in_280, // @[:@6.4]
  input  [4:0]  io_in_281, // @[:@6.4]
  input  [4:0]  io_in_282, // @[:@6.4]
  input  [4:0]  io_in_283, // @[:@6.4]
  input  [4:0]  io_in_284, // @[:@6.4]
  input  [4:0]  io_in_285, // @[:@6.4]
  input  [4:0]  io_in_286, // @[:@6.4]
  input  [4:0]  io_in_287, // @[:@6.4]
  input  [4:0]  io_in_288, // @[:@6.4]
  input  [4:0]  io_in_289, // @[:@6.4]
  input  [4:0]  io_in_290, // @[:@6.4]
  input  [4:0]  io_in_291, // @[:@6.4]
  input  [4:0]  io_in_292, // @[:@6.4]
  input  [4:0]  io_in_293, // @[:@6.4]
  input  [4:0]  io_in_294, // @[:@6.4]
  input  [4:0]  io_in_295, // @[:@6.4]
  input  [4:0]  io_in_296, // @[:@6.4]
  input  [4:0]  io_in_297, // @[:@6.4]
  input  [4:0]  io_in_298, // @[:@6.4]
  input  [4:0]  io_in_299, // @[:@6.4]
  input  [4:0]  io_in_300, // @[:@6.4]
  input  [4:0]  io_in_301, // @[:@6.4]
  input  [4:0]  io_in_302, // @[:@6.4]
  input  [4:0]  io_in_303, // @[:@6.4]
  input  [4:0]  io_in_304, // @[:@6.4]
  input  [4:0]  io_in_305, // @[:@6.4]
  input  [4:0]  io_in_306, // @[:@6.4]
  input  [4:0]  io_in_307, // @[:@6.4]
  input  [4:0]  io_in_308, // @[:@6.4]
  input  [4:0]  io_in_309, // @[:@6.4]
  input  [4:0]  io_in_310, // @[:@6.4]
  input  [4:0]  io_in_311, // @[:@6.4]
  input  [4:0]  io_in_312, // @[:@6.4]
  input  [4:0]  io_in_313, // @[:@6.4]
  input  [4:0]  io_in_314, // @[:@6.4]
  input  [4:0]  io_in_315, // @[:@6.4]
  input  [4:0]  io_in_316, // @[:@6.4]
  input  [4:0]  io_in_317, // @[:@6.4]
  input  [4:0]  io_in_318, // @[:@6.4]
  input  [4:0]  io_in_319, // @[:@6.4]
  input  [4:0]  io_in_320, // @[:@6.4]
  input  [4:0]  io_in_321, // @[:@6.4]
  input  [4:0]  io_in_322, // @[:@6.4]
  input  [4:0]  io_in_323, // @[:@6.4]
  input  [4:0]  io_in_324, // @[:@6.4]
  input  [4:0]  io_in_325, // @[:@6.4]
  input  [4:0]  io_in_326, // @[:@6.4]
  input  [4:0]  io_in_327, // @[:@6.4]
  input  [4:0]  io_in_328, // @[:@6.4]
  input  [4:0]  io_in_329, // @[:@6.4]
  input  [4:0]  io_in_330, // @[:@6.4]
  input  [4:0]  io_in_331, // @[:@6.4]
  input  [4:0]  io_in_332, // @[:@6.4]
  input  [4:0]  io_in_333, // @[:@6.4]
  input  [4:0]  io_in_334, // @[:@6.4]
  input  [4:0]  io_in_335, // @[:@6.4]
  input  [4:0]  io_in_336, // @[:@6.4]
  input  [4:0]  io_in_337, // @[:@6.4]
  input  [4:0]  io_in_338, // @[:@6.4]
  input  [4:0]  io_in_339, // @[:@6.4]
  input  [4:0]  io_in_340, // @[:@6.4]
  input  [4:0]  io_in_341, // @[:@6.4]
  input  [4:0]  io_in_342, // @[:@6.4]
  input  [4:0]  io_in_343, // @[:@6.4]
  input  [4:0]  io_in_344, // @[:@6.4]
  input  [4:0]  io_in_345, // @[:@6.4]
  input  [4:0]  io_in_346, // @[:@6.4]
  input  [4:0]  io_in_347, // @[:@6.4]
  input  [4:0]  io_in_348, // @[:@6.4]
  input  [4:0]  io_in_349, // @[:@6.4]
  input  [4:0]  io_in_350, // @[:@6.4]
  input  [4:0]  io_in_351, // @[:@6.4]
  input  [4:0]  io_in_352, // @[:@6.4]
  input  [4:0]  io_in_353, // @[:@6.4]
  input  [4:0]  io_in_354, // @[:@6.4]
  input  [4:0]  io_in_355, // @[:@6.4]
  input  [4:0]  io_in_356, // @[:@6.4]
  input  [4:0]  io_in_357, // @[:@6.4]
  input  [4:0]  io_in_358, // @[:@6.4]
  input  [4:0]  io_in_359, // @[:@6.4]
  input  [4:0]  io_in_360, // @[:@6.4]
  input  [4:0]  io_in_361, // @[:@6.4]
  input  [4:0]  io_in_362, // @[:@6.4]
  input  [4:0]  io_in_363, // @[:@6.4]
  input  [4:0]  io_in_364, // @[:@6.4]
  input  [4:0]  io_in_365, // @[:@6.4]
  input  [4:0]  io_in_366, // @[:@6.4]
  input  [4:0]  io_in_367, // @[:@6.4]
  input  [4:0]  io_in_368, // @[:@6.4]
  input  [4:0]  io_in_369, // @[:@6.4]
  input  [4:0]  io_in_370, // @[:@6.4]
  input  [4:0]  io_in_371, // @[:@6.4]
  input  [4:0]  io_in_372, // @[:@6.4]
  input  [4:0]  io_in_373, // @[:@6.4]
  input  [4:0]  io_in_374, // @[:@6.4]
  input  [4:0]  io_in_375, // @[:@6.4]
  input  [4:0]  io_in_376, // @[:@6.4]
  input  [4:0]  io_in_377, // @[:@6.4]
  input  [4:0]  io_in_378, // @[:@6.4]
  input  [4:0]  io_in_379, // @[:@6.4]
  input  [4:0]  io_in_380, // @[:@6.4]
  input  [4:0]  io_in_381, // @[:@6.4]
  input  [4:0]  io_in_382, // @[:@6.4]
  input  [4:0]  io_in_383, // @[:@6.4]
  input  [4:0]  io_in_384, // @[:@6.4]
  input  [4:0]  io_in_385, // @[:@6.4]
  input  [4:0]  io_in_386, // @[:@6.4]
  input  [4:0]  io_in_387, // @[:@6.4]
  input  [4:0]  io_in_388, // @[:@6.4]
  input  [4:0]  io_in_389, // @[:@6.4]
  input  [4:0]  io_in_390, // @[:@6.4]
  input  [4:0]  io_in_391, // @[:@6.4]
  input  [4:0]  io_in_392, // @[:@6.4]
  input  [4:0]  io_in_393, // @[:@6.4]
  input  [4:0]  io_in_394, // @[:@6.4]
  input  [4:0]  io_in_395, // @[:@6.4]
  input  [4:0]  io_in_396, // @[:@6.4]
  input  [4:0]  io_in_397, // @[:@6.4]
  input  [4:0]  io_in_398, // @[:@6.4]
  input  [4:0]  io_in_399, // @[:@6.4]
  input  [4:0]  io_in_400, // @[:@6.4]
  input  [4:0]  io_in_401, // @[:@6.4]
  input  [4:0]  io_in_402, // @[:@6.4]
  input  [4:0]  io_in_403, // @[:@6.4]
  input  [4:0]  io_in_404, // @[:@6.4]
  input  [4:0]  io_in_405, // @[:@6.4]
  input  [4:0]  io_in_406, // @[:@6.4]
  input  [4:0]  io_in_407, // @[:@6.4]
  input  [4:0]  io_in_408, // @[:@6.4]
  input  [4:0]  io_in_409, // @[:@6.4]
  input  [4:0]  io_in_410, // @[:@6.4]
  input  [4:0]  io_in_411, // @[:@6.4]
  input  [4:0]  io_in_412, // @[:@6.4]
  input  [4:0]  io_in_413, // @[:@6.4]
  input  [4:0]  io_in_414, // @[:@6.4]
  input  [4:0]  io_in_415, // @[:@6.4]
  input  [4:0]  io_in_416, // @[:@6.4]
  input  [4:0]  io_in_417, // @[:@6.4]
  input  [4:0]  io_in_418, // @[:@6.4]
  input  [4:0]  io_in_419, // @[:@6.4]
  input  [4:0]  io_in_420, // @[:@6.4]
  input  [4:0]  io_in_421, // @[:@6.4]
  input  [4:0]  io_in_422, // @[:@6.4]
  input  [4:0]  io_in_423, // @[:@6.4]
  input  [4:0]  io_in_424, // @[:@6.4]
  input  [4:0]  io_in_425, // @[:@6.4]
  input  [4:0]  io_in_426, // @[:@6.4]
  input  [4:0]  io_in_427, // @[:@6.4]
  input  [4:0]  io_in_428, // @[:@6.4]
  input  [4:0]  io_in_429, // @[:@6.4]
  input  [4:0]  io_in_430, // @[:@6.4]
  input  [4:0]  io_in_431, // @[:@6.4]
  input  [4:0]  io_in_432, // @[:@6.4]
  input  [4:0]  io_in_433, // @[:@6.4]
  input  [4:0]  io_in_434, // @[:@6.4]
  input  [4:0]  io_in_435, // @[:@6.4]
  input  [4:0]  io_in_436, // @[:@6.4]
  input  [4:0]  io_in_437, // @[:@6.4]
  input  [4:0]  io_in_438, // @[:@6.4]
  input  [4:0]  io_in_439, // @[:@6.4]
  input  [4:0]  io_in_440, // @[:@6.4]
  input  [4:0]  io_in_441, // @[:@6.4]
  input  [4:0]  io_in_442, // @[:@6.4]
  input  [4:0]  io_in_443, // @[:@6.4]
  input  [4:0]  io_in_444, // @[:@6.4]
  input  [4:0]  io_in_445, // @[:@6.4]
  input  [4:0]  io_in_446, // @[:@6.4]
  input  [4:0]  io_in_447, // @[:@6.4]
  input  [4:0]  io_in_448, // @[:@6.4]
  input  [4:0]  io_in_449, // @[:@6.4]
  input  [4:0]  io_in_450, // @[:@6.4]
  input  [4:0]  io_in_451, // @[:@6.4]
  input  [4:0]  io_in_452, // @[:@6.4]
  input  [4:0]  io_in_453, // @[:@6.4]
  input  [4:0]  io_in_454, // @[:@6.4]
  input  [4:0]  io_in_455, // @[:@6.4]
  input  [4:0]  io_in_456, // @[:@6.4]
  input  [4:0]  io_in_457, // @[:@6.4]
  input  [4:0]  io_in_458, // @[:@6.4]
  input  [4:0]  io_in_459, // @[:@6.4]
  input  [4:0]  io_in_460, // @[:@6.4]
  input  [4:0]  io_in_461, // @[:@6.4]
  input  [4:0]  io_in_462, // @[:@6.4]
  input  [4:0]  io_in_463, // @[:@6.4]
  input  [4:0]  io_in_464, // @[:@6.4]
  input  [4:0]  io_in_465, // @[:@6.4]
  input  [4:0]  io_in_466, // @[:@6.4]
  input  [4:0]  io_in_467, // @[:@6.4]
  input  [4:0]  io_in_468, // @[:@6.4]
  input  [4:0]  io_in_469, // @[:@6.4]
  input  [4:0]  io_in_470, // @[:@6.4]
  input  [4:0]  io_in_471, // @[:@6.4]
  input  [4:0]  io_in_472, // @[:@6.4]
  input  [4:0]  io_in_473, // @[:@6.4]
  input  [4:0]  io_in_474, // @[:@6.4]
  input  [4:0]  io_in_475, // @[:@6.4]
  input  [4:0]  io_in_476, // @[:@6.4]
  input  [4:0]  io_in_477, // @[:@6.4]
  input  [4:0]  io_in_478, // @[:@6.4]
  input  [4:0]  io_in_479, // @[:@6.4]
  input  [4:0]  io_in_480, // @[:@6.4]
  input  [4:0]  io_in_481, // @[:@6.4]
  input  [4:0]  io_in_482, // @[:@6.4]
  input  [4:0]  io_in_483, // @[:@6.4]
  input  [4:0]  io_in_484, // @[:@6.4]
  input  [4:0]  io_in_485, // @[:@6.4]
  input  [4:0]  io_in_486, // @[:@6.4]
  input  [4:0]  io_in_487, // @[:@6.4]
  input  [4:0]  io_in_488, // @[:@6.4]
  input  [4:0]  io_in_489, // @[:@6.4]
  input  [4:0]  io_in_490, // @[:@6.4]
  input  [4:0]  io_in_491, // @[:@6.4]
  input  [4:0]  io_in_492, // @[:@6.4]
  input  [4:0]  io_in_493, // @[:@6.4]
  input  [4:0]  io_in_494, // @[:@6.4]
  input  [4:0]  io_in_495, // @[:@6.4]
  input  [4:0]  io_in_496, // @[:@6.4]
  input  [4:0]  io_in_497, // @[:@6.4]
  input  [4:0]  io_in_498, // @[:@6.4]
  input  [4:0]  io_in_499, // @[:@6.4]
  input  [4:0]  io_in_500, // @[:@6.4]
  input  [4:0]  io_in_501, // @[:@6.4]
  input  [4:0]  io_in_502, // @[:@6.4]
  input  [4:0]  io_in_503, // @[:@6.4]
  input  [4:0]  io_in_504, // @[:@6.4]
  input  [4:0]  io_in_505, // @[:@6.4]
  input  [4:0]  io_in_506, // @[:@6.4]
  input  [4:0]  io_in_507, // @[:@6.4]
  input  [4:0]  io_in_508, // @[:@6.4]
  input  [4:0]  io_in_509, // @[:@6.4]
  input  [4:0]  io_in_510, // @[:@6.4]
  input  [4:0]  io_in_511, // @[:@6.4]
  input  [4:0]  io_in_512, // @[:@6.4]
  input  [4:0]  io_in_513, // @[:@6.4]
  input  [4:0]  io_in_514, // @[:@6.4]
  input  [4:0]  io_in_515, // @[:@6.4]
  input  [4:0]  io_in_516, // @[:@6.4]
  input  [4:0]  io_in_517, // @[:@6.4]
  input  [4:0]  io_in_518, // @[:@6.4]
  input  [4:0]  io_in_519, // @[:@6.4]
  input  [4:0]  io_in_520, // @[:@6.4]
  input  [4:0]  io_in_521, // @[:@6.4]
  input  [4:0]  io_in_522, // @[:@6.4]
  input  [4:0]  io_in_523, // @[:@6.4]
  input  [4:0]  io_in_524, // @[:@6.4]
  input  [4:0]  io_in_525, // @[:@6.4]
  input  [4:0]  io_in_526, // @[:@6.4]
  input  [4:0]  io_in_527, // @[:@6.4]
  input  [4:0]  io_in_528, // @[:@6.4]
  input  [4:0]  io_in_529, // @[:@6.4]
  input  [4:0]  io_in_530, // @[:@6.4]
  input  [4:0]  io_in_531, // @[:@6.4]
  input  [4:0]  io_in_532, // @[:@6.4]
  input  [4:0]  io_in_533, // @[:@6.4]
  input  [4:0]  io_in_534, // @[:@6.4]
  input  [4:0]  io_in_535, // @[:@6.4]
  input  [4:0]  io_in_536, // @[:@6.4]
  input  [4:0]  io_in_537, // @[:@6.4]
  input  [4:0]  io_in_538, // @[:@6.4]
  input  [4:0]  io_in_539, // @[:@6.4]
  input  [4:0]  io_in_540, // @[:@6.4]
  input  [4:0]  io_in_541, // @[:@6.4]
  input  [4:0]  io_in_542, // @[:@6.4]
  input  [4:0]  io_in_543, // @[:@6.4]
  input  [4:0]  io_in_544, // @[:@6.4]
  input  [4:0]  io_in_545, // @[:@6.4]
  input  [4:0]  io_in_546, // @[:@6.4]
  input  [4:0]  io_in_547, // @[:@6.4]
  input  [4:0]  io_in_548, // @[:@6.4]
  input  [4:0]  io_in_549, // @[:@6.4]
  input  [4:0]  io_in_550, // @[:@6.4]
  input  [4:0]  io_in_551, // @[:@6.4]
  input  [4:0]  io_in_552, // @[:@6.4]
  input  [4:0]  io_in_553, // @[:@6.4]
  input  [4:0]  io_in_554, // @[:@6.4]
  input  [4:0]  io_in_555, // @[:@6.4]
  input  [4:0]  io_in_556, // @[:@6.4]
  input  [4:0]  io_in_557, // @[:@6.4]
  input  [4:0]  io_in_558, // @[:@6.4]
  input  [4:0]  io_in_559, // @[:@6.4]
  input  [4:0]  io_in_560, // @[:@6.4]
  input  [4:0]  io_in_561, // @[:@6.4]
  input  [4:0]  io_in_562, // @[:@6.4]
  input  [4:0]  io_in_563, // @[:@6.4]
  input  [4:0]  io_in_564, // @[:@6.4]
  input  [4:0]  io_in_565, // @[:@6.4]
  input  [4:0]  io_in_566, // @[:@6.4]
  input  [4:0]  io_in_567, // @[:@6.4]
  input  [4:0]  io_in_568, // @[:@6.4]
  input  [4:0]  io_in_569, // @[:@6.4]
  input  [4:0]  io_in_570, // @[:@6.4]
  input  [4:0]  io_in_571, // @[:@6.4]
  input  [4:0]  io_in_572, // @[:@6.4]
  input  [4:0]  io_in_573, // @[:@6.4]
  input  [4:0]  io_in_574, // @[:@6.4]
  input  [4:0]  io_in_575, // @[:@6.4]
  input  [4:0]  io_in_576, // @[:@6.4]
  input  [4:0]  io_in_577, // @[:@6.4]
  input  [4:0]  io_in_578, // @[:@6.4]
  input  [4:0]  io_in_579, // @[:@6.4]
  input  [4:0]  io_in_580, // @[:@6.4]
  input  [4:0]  io_in_581, // @[:@6.4]
  input  [4:0]  io_in_582, // @[:@6.4]
  input  [4:0]  io_in_583, // @[:@6.4]
  input  [4:0]  io_in_584, // @[:@6.4]
  input  [4:0]  io_in_585, // @[:@6.4]
  input  [4:0]  io_in_586, // @[:@6.4]
  input  [4:0]  io_in_587, // @[:@6.4]
  input  [4:0]  io_in_588, // @[:@6.4]
  input  [4:0]  io_in_589, // @[:@6.4]
  input  [4:0]  io_in_590, // @[:@6.4]
  input  [4:0]  io_in_591, // @[:@6.4]
  input  [4:0]  io_in_592, // @[:@6.4]
  input  [4:0]  io_in_593, // @[:@6.4]
  input  [4:0]  io_in_594, // @[:@6.4]
  input  [4:0]  io_in_595, // @[:@6.4]
  input  [4:0]  io_in_596, // @[:@6.4]
  input  [4:0]  io_in_597, // @[:@6.4]
  input  [4:0]  io_in_598, // @[:@6.4]
  input  [4:0]  io_in_599, // @[:@6.4]
  input  [4:0]  io_in_600, // @[:@6.4]
  input  [4:0]  io_in_601, // @[:@6.4]
  input  [4:0]  io_in_602, // @[:@6.4]
  input  [4:0]  io_in_603, // @[:@6.4]
  input  [4:0]  io_in_604, // @[:@6.4]
  input  [4:0]  io_in_605, // @[:@6.4]
  input  [4:0]  io_in_606, // @[:@6.4]
  input  [4:0]  io_in_607, // @[:@6.4]
  input  [4:0]  io_in_608, // @[:@6.4]
  input  [4:0]  io_in_609, // @[:@6.4]
  input  [4:0]  io_in_610, // @[:@6.4]
  input  [4:0]  io_in_611, // @[:@6.4]
  input  [4:0]  io_in_612, // @[:@6.4]
  input  [4:0]  io_in_613, // @[:@6.4]
  input  [4:0]  io_in_614, // @[:@6.4]
  input  [4:0]  io_in_615, // @[:@6.4]
  input  [4:0]  io_in_616, // @[:@6.4]
  input  [4:0]  io_in_617, // @[:@6.4]
  input  [4:0]  io_in_618, // @[:@6.4]
  input  [4:0]  io_in_619, // @[:@6.4]
  input  [4:0]  io_in_620, // @[:@6.4]
  input  [4:0]  io_in_621, // @[:@6.4]
  input  [4:0]  io_in_622, // @[:@6.4]
  input  [4:0]  io_in_623, // @[:@6.4]
  input  [4:0]  io_in_624, // @[:@6.4]
  input  [4:0]  io_in_625, // @[:@6.4]
  input  [4:0]  io_in_626, // @[:@6.4]
  input  [4:0]  io_in_627, // @[:@6.4]
  input  [4:0]  io_in_628, // @[:@6.4]
  input  [4:0]  io_in_629, // @[:@6.4]
  input  [4:0]  io_in_630, // @[:@6.4]
  input  [4:0]  io_in_631, // @[:@6.4]
  input  [4:0]  io_in_632, // @[:@6.4]
  input  [4:0]  io_in_633, // @[:@6.4]
  input  [4:0]  io_in_634, // @[:@6.4]
  input  [4:0]  io_in_635, // @[:@6.4]
  input  [4:0]  io_in_636, // @[:@6.4]
  input  [4:0]  io_in_637, // @[:@6.4]
  input  [4:0]  io_in_638, // @[:@6.4]
  input  [4:0]  io_in_639, // @[:@6.4]
  input  [4:0]  io_in_640, // @[:@6.4]
  input  [4:0]  io_in_641, // @[:@6.4]
  input  [4:0]  io_in_642, // @[:@6.4]
  input  [4:0]  io_in_643, // @[:@6.4]
  input  [4:0]  io_in_644, // @[:@6.4]
  input  [4:0]  io_in_645, // @[:@6.4]
  input  [4:0]  io_in_646, // @[:@6.4]
  input  [4:0]  io_in_647, // @[:@6.4]
  input  [4:0]  io_in_648, // @[:@6.4]
  input  [4:0]  io_in_649, // @[:@6.4]
  input  [4:0]  io_in_650, // @[:@6.4]
  input  [4:0]  io_in_651, // @[:@6.4]
  input  [4:0]  io_in_652, // @[:@6.4]
  input  [4:0]  io_in_653, // @[:@6.4]
  input  [4:0]  io_in_654, // @[:@6.4]
  input  [4:0]  io_in_655, // @[:@6.4]
  input  [4:0]  io_in_656, // @[:@6.4]
  input  [4:0]  io_in_657, // @[:@6.4]
  input  [4:0]  io_in_658, // @[:@6.4]
  input  [4:0]  io_in_659, // @[:@6.4]
  input  [4:0]  io_in_660, // @[:@6.4]
  input  [4:0]  io_in_661, // @[:@6.4]
  input  [4:0]  io_in_662, // @[:@6.4]
  input  [4:0]  io_in_663, // @[:@6.4]
  input  [4:0]  io_in_664, // @[:@6.4]
  input  [4:0]  io_in_665, // @[:@6.4]
  input  [4:0]  io_in_666, // @[:@6.4]
  input  [4:0]  io_in_667, // @[:@6.4]
  input  [4:0]  io_in_668, // @[:@6.4]
  input  [4:0]  io_in_669, // @[:@6.4]
  input  [4:0]  io_in_670, // @[:@6.4]
  input  [4:0]  io_in_671, // @[:@6.4]
  input  [4:0]  io_in_672, // @[:@6.4]
  input  [4:0]  io_in_673, // @[:@6.4]
  input  [4:0]  io_in_674, // @[:@6.4]
  input  [4:0]  io_in_675, // @[:@6.4]
  input  [4:0]  io_in_676, // @[:@6.4]
  input  [4:0]  io_in_677, // @[:@6.4]
  input  [4:0]  io_in_678, // @[:@6.4]
  input  [4:0]  io_in_679, // @[:@6.4]
  input  [4:0]  io_in_680, // @[:@6.4]
  input  [4:0]  io_in_681, // @[:@6.4]
  input  [4:0]  io_in_682, // @[:@6.4]
  input  [4:0]  io_in_683, // @[:@6.4]
  input  [4:0]  io_in_684, // @[:@6.4]
  input  [4:0]  io_in_685, // @[:@6.4]
  input  [4:0]  io_in_686, // @[:@6.4]
  input  [4:0]  io_in_687, // @[:@6.4]
  input  [4:0]  io_in_688, // @[:@6.4]
  input  [4:0]  io_in_689, // @[:@6.4]
  input  [4:0]  io_in_690, // @[:@6.4]
  input  [4:0]  io_in_691, // @[:@6.4]
  input  [4:0]  io_in_692, // @[:@6.4]
  input  [4:0]  io_in_693, // @[:@6.4]
  input  [4:0]  io_in_694, // @[:@6.4]
  input  [4:0]  io_in_695, // @[:@6.4]
  input  [4:0]  io_in_696, // @[:@6.4]
  input  [4:0]  io_in_697, // @[:@6.4]
  input  [4:0]  io_in_698, // @[:@6.4]
  input  [4:0]  io_in_699, // @[:@6.4]
  input  [4:0]  io_in_700, // @[:@6.4]
  input  [4:0]  io_in_701, // @[:@6.4]
  input  [4:0]  io_in_702, // @[:@6.4]
  input  [4:0]  io_in_703, // @[:@6.4]
  input  [4:0]  io_in_704, // @[:@6.4]
  input  [4:0]  io_in_705, // @[:@6.4]
  input  [4:0]  io_in_706, // @[:@6.4]
  input  [4:0]  io_in_707, // @[:@6.4]
  input  [4:0]  io_in_708, // @[:@6.4]
  input  [4:0]  io_in_709, // @[:@6.4]
  input  [4:0]  io_in_710, // @[:@6.4]
  input  [4:0]  io_in_711, // @[:@6.4]
  input  [4:0]  io_in_712, // @[:@6.4]
  input  [4:0]  io_in_713, // @[:@6.4]
  input  [4:0]  io_in_714, // @[:@6.4]
  input  [4:0]  io_in_715, // @[:@6.4]
  input  [4:0]  io_in_716, // @[:@6.4]
  input  [4:0]  io_in_717, // @[:@6.4]
  input  [4:0]  io_in_718, // @[:@6.4]
  input  [4:0]  io_in_719, // @[:@6.4]
  input  [4:0]  io_in_720, // @[:@6.4]
  input  [4:0]  io_in_721, // @[:@6.4]
  input  [4:0]  io_in_722, // @[:@6.4]
  input  [4:0]  io_in_723, // @[:@6.4]
  input  [4:0]  io_in_724, // @[:@6.4]
  input  [4:0]  io_in_725, // @[:@6.4]
  input  [4:0]  io_in_726, // @[:@6.4]
  input  [4:0]  io_in_727, // @[:@6.4]
  input  [4:0]  io_in_728, // @[:@6.4]
  input  [4:0]  io_in_729, // @[:@6.4]
  input  [4:0]  io_in_730, // @[:@6.4]
  input  [4:0]  io_in_731, // @[:@6.4]
  input  [4:0]  io_in_732, // @[:@6.4]
  input  [4:0]  io_in_733, // @[:@6.4]
  input  [4:0]  io_in_734, // @[:@6.4]
  input  [4:0]  io_in_735, // @[:@6.4]
  input  [4:0]  io_in_736, // @[:@6.4]
  input  [4:0]  io_in_737, // @[:@6.4]
  input  [4:0]  io_in_738, // @[:@6.4]
  input  [4:0]  io_in_739, // @[:@6.4]
  input  [4:0]  io_in_740, // @[:@6.4]
  input  [4:0]  io_in_741, // @[:@6.4]
  input  [4:0]  io_in_742, // @[:@6.4]
  input  [4:0]  io_in_743, // @[:@6.4]
  input  [4:0]  io_in_744, // @[:@6.4]
  input  [4:0]  io_in_745, // @[:@6.4]
  input  [4:0]  io_in_746, // @[:@6.4]
  input  [4:0]  io_in_747, // @[:@6.4]
  input  [4:0]  io_in_748, // @[:@6.4]
  input  [4:0]  io_in_749, // @[:@6.4]
  input  [4:0]  io_in_750, // @[:@6.4]
  input  [4:0]  io_in_751, // @[:@6.4]
  input  [4:0]  io_in_752, // @[:@6.4]
  input  [4:0]  io_in_753, // @[:@6.4]
  input  [4:0]  io_in_754, // @[:@6.4]
  input  [4:0]  io_in_755, // @[:@6.4]
  input  [4:0]  io_in_756, // @[:@6.4]
  input  [4:0]  io_in_757, // @[:@6.4]
  input  [4:0]  io_in_758, // @[:@6.4]
  input  [4:0]  io_in_759, // @[:@6.4]
  input  [4:0]  io_in_760, // @[:@6.4]
  input  [4:0]  io_in_761, // @[:@6.4]
  input  [4:0]  io_in_762, // @[:@6.4]
  input  [4:0]  io_in_763, // @[:@6.4]
  input  [4:0]  io_in_764, // @[:@6.4]
  input  [4:0]  io_in_765, // @[:@6.4]
  input  [4:0]  io_in_766, // @[:@6.4]
  input  [4:0]  io_in_767, // @[:@6.4]
  input  [4:0]  io_in_768, // @[:@6.4]
  input  [4:0]  io_in_769, // @[:@6.4]
  input  [4:0]  io_in_770, // @[:@6.4]
  input  [4:0]  io_in_771, // @[:@6.4]
  input  [4:0]  io_in_772, // @[:@6.4]
  input  [4:0]  io_in_773, // @[:@6.4]
  input  [4:0]  io_in_774, // @[:@6.4]
  input  [4:0]  io_in_775, // @[:@6.4]
  input  [4:0]  io_in_776, // @[:@6.4]
  input  [4:0]  io_in_777, // @[:@6.4]
  input  [4:0]  io_in_778, // @[:@6.4]
  input  [4:0]  io_in_779, // @[:@6.4]
  input  [4:0]  io_in_780, // @[:@6.4]
  input  [4:0]  io_in_781, // @[:@6.4]
  input  [4:0]  io_in_782, // @[:@6.4]
  input  [4:0]  io_in_783, // @[:@6.4]
  output [10:0] io_out_0, // @[:@6.4]
  output [10:0] io_out_1, // @[:@6.4]
  output [10:0] io_out_2, // @[:@6.4]
  output [10:0] io_out_3, // @[:@6.4]
  output [10:0] io_out_4, // @[:@6.4]
  output [10:0] io_out_5, // @[:@6.4]
  output [10:0] io_out_6, // @[:@6.4]
  output [10:0] io_out_7, // @[:@6.4]
  output [10:0] io_out_8, // @[:@6.4]
  output [10:0] io_out_9, // @[:@6.4]
  output [10:0] io_out_10, // @[:@6.4]
  output [10:0] io_out_11, // @[:@6.4]
  output [10:0] io_out_12, // @[:@6.4]
  output [10:0] io_out_13, // @[:@6.4]
  output [10:0] io_out_14, // @[:@6.4]
  output [10:0] io_out_15 // @[:@6.4]
);
  wire [5:0] _T_54267; // @[Modules.scala 43:37:@9.4]
  wire [4:0] _T_54268; // @[Modules.scala 43:37:@10.4]
  wire [4:0] _T_54269; // @[Modules.scala 43:37:@11.4]
  wire [5:0] _T_54270; // @[Modules.scala 43:47:@12.4]
  wire [4:0] _T_54271; // @[Modules.scala 43:47:@13.4]
  wire [4:0] _T_54272; // @[Modules.scala 43:47:@14.4]
  wire [5:0] _T_54274; // @[Modules.scala 46:37:@16.4]
  wire [4:0] _T_54275; // @[Modules.scala 46:37:@17.4]
  wire [4:0] _T_54276; // @[Modules.scala 46:37:@18.4]
  wire [5:0] _T_54277; // @[Modules.scala 46:47:@19.4]
  wire [4:0] _T_54278; // @[Modules.scala 46:47:@20.4]
  wire [4:0] _T_54279; // @[Modules.scala 46:47:@21.4]
  wire [5:0] _T_54281; // @[Modules.scala 43:37:@23.4]
  wire [4:0] _T_54282; // @[Modules.scala 43:37:@24.4]
  wire [4:0] _T_54283; // @[Modules.scala 43:37:@25.4]
  wire [5:0] _T_54284; // @[Modules.scala 43:47:@26.4]
  wire [4:0] _T_54285; // @[Modules.scala 43:47:@27.4]
  wire [4:0] _T_54286; // @[Modules.scala 43:47:@28.4]
  wire [5:0] _T_54288; // @[Modules.scala 43:37:@30.4]
  wire [4:0] _T_54289; // @[Modules.scala 43:37:@31.4]
  wire [4:0] _T_54290; // @[Modules.scala 43:37:@32.4]
  wire [5:0] _T_54291; // @[Modules.scala 43:47:@33.4]
  wire [4:0] _T_54292; // @[Modules.scala 43:47:@34.4]
  wire [4:0] _T_54293; // @[Modules.scala 43:47:@35.4]
  wire [5:0] _T_54295; // @[Modules.scala 43:37:@37.4]
  wire [4:0] _T_54296; // @[Modules.scala 43:37:@38.4]
  wire [4:0] _T_54297; // @[Modules.scala 43:37:@39.4]
  wire [5:0] _T_54298; // @[Modules.scala 43:47:@40.4]
  wire [4:0] _T_54299; // @[Modules.scala 43:47:@41.4]
  wire [4:0] _T_54300; // @[Modules.scala 43:47:@42.4]
  wire [5:0] _T_54302; // @[Modules.scala 46:37:@44.4]
  wire [4:0] _T_54303; // @[Modules.scala 46:37:@45.4]
  wire [4:0] _T_54304; // @[Modules.scala 46:37:@46.4]
  wire [5:0] _T_54305; // @[Modules.scala 46:47:@47.4]
  wire [4:0] _T_54306; // @[Modules.scala 46:47:@48.4]
  wire [4:0] _T_54307; // @[Modules.scala 46:47:@49.4]
  wire [5:0] _T_54309; // @[Modules.scala 46:37:@51.4]
  wire [4:0] _T_54310; // @[Modules.scala 46:37:@52.4]
  wire [4:0] _T_54311; // @[Modules.scala 46:37:@53.4]
  wire [5:0] _T_54312; // @[Modules.scala 46:47:@54.4]
  wire [4:0] _T_54313; // @[Modules.scala 46:47:@55.4]
  wire [4:0] _T_54314; // @[Modules.scala 46:47:@56.4]
  wire [5:0] _T_54316; // @[Modules.scala 46:37:@58.4]
  wire [4:0] _T_54317; // @[Modules.scala 46:37:@59.4]
  wire [4:0] _T_54318; // @[Modules.scala 46:37:@60.4]
  wire [5:0] _T_54319; // @[Modules.scala 46:47:@61.4]
  wire [4:0] _T_54320; // @[Modules.scala 46:47:@62.4]
  wire [4:0] _T_54321; // @[Modules.scala 46:47:@63.4]
  wire [5:0] _T_54322; // @[Modules.scala 37:46:@65.4]
  wire [4:0] _T_54323; // @[Modules.scala 37:46:@66.4]
  wire [4:0] _T_54324; // @[Modules.scala 37:46:@67.4]
  wire [5:0] _T_54326; // @[Modules.scala 46:37:@69.4]
  wire [4:0] _T_54327; // @[Modules.scala 46:37:@70.4]
  wire [4:0] _T_54328; // @[Modules.scala 46:37:@71.4]
  wire [5:0] _T_54329; // @[Modules.scala 46:47:@72.4]
  wire [4:0] _T_54330; // @[Modules.scala 46:47:@73.4]
  wire [4:0] _T_54331; // @[Modules.scala 46:47:@74.4]
  wire [5:0] _T_54332; // @[Modules.scala 37:46:@76.4]
  wire [4:0] _T_54333; // @[Modules.scala 37:46:@77.4]
  wire [4:0] _T_54334; // @[Modules.scala 37:46:@78.4]
  wire [5:0] _T_54336; // @[Modules.scala 43:37:@80.4]
  wire [4:0] _T_54337; // @[Modules.scala 43:37:@81.4]
  wire [4:0] _T_54338; // @[Modules.scala 43:37:@82.4]
  wire [5:0] _T_54339; // @[Modules.scala 43:47:@83.4]
  wire [4:0] _T_54340; // @[Modules.scala 43:47:@84.4]
  wire [4:0] _T_54341; // @[Modules.scala 43:47:@85.4]
  wire [5:0] _T_54343; // @[Modules.scala 43:37:@87.4]
  wire [4:0] _T_54344; // @[Modules.scala 43:37:@88.4]
  wire [4:0] _T_54345; // @[Modules.scala 43:37:@89.4]
  wire [5:0] _T_54346; // @[Modules.scala 43:47:@90.4]
  wire [4:0] _T_54347; // @[Modules.scala 43:47:@91.4]
  wire [4:0] _T_54348; // @[Modules.scala 43:47:@92.4]
  wire [5:0] _T_54349; // @[Modules.scala 40:46:@94.4]
  wire [4:0] _T_54350; // @[Modules.scala 40:46:@95.4]
  wire [4:0] _T_54351; // @[Modules.scala 40:46:@96.4]
  wire [5:0] _T_54353; // @[Modules.scala 46:37:@98.4]
  wire [4:0] _T_54354; // @[Modules.scala 46:37:@99.4]
  wire [4:0] _T_54355; // @[Modules.scala 46:37:@100.4]
  wire [5:0] _T_54356; // @[Modules.scala 46:47:@101.4]
  wire [4:0] _T_54357; // @[Modules.scala 46:47:@102.4]
  wire [4:0] _T_54358; // @[Modules.scala 46:47:@103.4]
  wire [5:0] _T_54360; // @[Modules.scala 43:37:@105.4]
  wire [4:0] _T_54361; // @[Modules.scala 43:37:@106.4]
  wire [4:0] _T_54362; // @[Modules.scala 43:37:@107.4]
  wire [5:0] _T_54363; // @[Modules.scala 43:47:@108.4]
  wire [4:0] _T_54364; // @[Modules.scala 43:47:@109.4]
  wire [4:0] _T_54365; // @[Modules.scala 43:47:@110.4]
  wire [5:0] _T_54366; // @[Modules.scala 37:46:@112.4]
  wire [4:0] _T_54367; // @[Modules.scala 37:46:@113.4]
  wire [4:0] _T_54368; // @[Modules.scala 37:46:@114.4]
  wire [5:0] _T_54370; // @[Modules.scala 46:37:@116.4]
  wire [4:0] _T_54371; // @[Modules.scala 46:37:@117.4]
  wire [4:0] _T_54372; // @[Modules.scala 46:37:@118.4]
  wire [5:0] _T_54373; // @[Modules.scala 46:47:@119.4]
  wire [4:0] _T_54374; // @[Modules.scala 46:47:@120.4]
  wire [4:0] _T_54375; // @[Modules.scala 46:47:@121.4]
  wire [5:0] _T_54377; // @[Modules.scala 46:37:@123.4]
  wire [4:0] _T_54378; // @[Modules.scala 46:37:@124.4]
  wire [4:0] _T_54379; // @[Modules.scala 46:37:@125.4]
  wire [5:0] _T_54380; // @[Modules.scala 46:47:@126.4]
  wire [4:0] _T_54381; // @[Modules.scala 46:47:@127.4]
  wire [4:0] _T_54382; // @[Modules.scala 46:47:@128.4]
  wire [5:0] _T_54384; // @[Modules.scala 46:37:@130.4]
  wire [4:0] _T_54385; // @[Modules.scala 46:37:@131.4]
  wire [4:0] _T_54386; // @[Modules.scala 46:37:@132.4]
  wire [5:0] _T_54387; // @[Modules.scala 46:47:@133.4]
  wire [4:0] _T_54388; // @[Modules.scala 46:47:@134.4]
  wire [4:0] _T_54389; // @[Modules.scala 46:47:@135.4]
  wire [5:0] _T_54391; // @[Modules.scala 46:37:@137.4]
  wire [4:0] _T_54392; // @[Modules.scala 46:37:@138.4]
  wire [4:0] _T_54393; // @[Modules.scala 46:37:@139.4]
  wire [5:0] _T_54394; // @[Modules.scala 46:47:@140.4]
  wire [4:0] _T_54395; // @[Modules.scala 46:47:@141.4]
  wire [4:0] _T_54396; // @[Modules.scala 46:47:@142.4]
  wire [5:0] _T_54398; // @[Modules.scala 46:37:@144.4]
  wire [4:0] _T_54399; // @[Modules.scala 46:37:@145.4]
  wire [4:0] _T_54400; // @[Modules.scala 46:37:@146.4]
  wire [5:0] _T_54401; // @[Modules.scala 46:47:@147.4]
  wire [4:0] _T_54402; // @[Modules.scala 46:47:@148.4]
  wire [4:0] _T_54403; // @[Modules.scala 46:47:@149.4]
  wire [5:0] _T_54405; // @[Modules.scala 46:37:@151.4]
  wire [4:0] _T_54406; // @[Modules.scala 46:37:@152.4]
  wire [4:0] _T_54407; // @[Modules.scala 46:37:@153.4]
  wire [5:0] _T_54408; // @[Modules.scala 46:47:@154.4]
  wire [4:0] _T_54409; // @[Modules.scala 46:47:@155.4]
  wire [4:0] _T_54410; // @[Modules.scala 46:47:@156.4]
  wire [5:0] _T_54412; // @[Modules.scala 46:37:@158.4]
  wire [4:0] _T_54413; // @[Modules.scala 46:37:@159.4]
  wire [4:0] _T_54414; // @[Modules.scala 46:37:@160.4]
  wire [5:0] _T_54415; // @[Modules.scala 46:47:@161.4]
  wire [4:0] _T_54416; // @[Modules.scala 46:47:@162.4]
  wire [4:0] _T_54417; // @[Modules.scala 46:47:@163.4]
  wire [5:0] _T_54419; // @[Modules.scala 46:37:@165.4]
  wire [4:0] _T_54420; // @[Modules.scala 46:37:@166.4]
  wire [4:0] _T_54421; // @[Modules.scala 46:37:@167.4]
  wire [5:0] _T_54422; // @[Modules.scala 46:47:@168.4]
  wire [4:0] _T_54423; // @[Modules.scala 46:47:@169.4]
  wire [4:0] _T_54424; // @[Modules.scala 46:47:@170.4]
  wire [5:0] _T_54426; // @[Modules.scala 46:37:@172.4]
  wire [4:0] _T_54427; // @[Modules.scala 46:37:@173.4]
  wire [4:0] _T_54428; // @[Modules.scala 46:37:@174.4]
  wire [5:0] _T_54429; // @[Modules.scala 46:47:@175.4]
  wire [4:0] _T_54430; // @[Modules.scala 46:47:@176.4]
  wire [4:0] _T_54431; // @[Modules.scala 46:47:@177.4]
  wire [5:0] _T_54432; // @[Modules.scala 37:46:@179.4]
  wire [4:0] _T_54433; // @[Modules.scala 37:46:@180.4]
  wire [4:0] _T_54434; // @[Modules.scala 37:46:@181.4]
  wire [5:0] _T_54435; // @[Modules.scala 40:46:@183.4]
  wire [4:0] _T_54436; // @[Modules.scala 40:46:@184.4]
  wire [4:0] _T_54437; // @[Modules.scala 40:46:@185.4]
  wire [5:0] _T_54438; // @[Modules.scala 40:46:@187.4]
  wire [4:0] _T_54439; // @[Modules.scala 40:46:@188.4]
  wire [4:0] _T_54440; // @[Modules.scala 40:46:@189.4]
  wire [5:0] _T_54442; // @[Modules.scala 46:37:@191.4]
  wire [4:0] _T_54443; // @[Modules.scala 46:37:@192.4]
  wire [4:0] _T_54444; // @[Modules.scala 46:37:@193.4]
  wire [5:0] _T_54445; // @[Modules.scala 46:47:@194.4]
  wire [4:0] _T_54446; // @[Modules.scala 46:47:@195.4]
  wire [4:0] _T_54447; // @[Modules.scala 46:47:@196.4]
  wire [5:0] _T_54449; // @[Modules.scala 46:37:@198.4]
  wire [4:0] _T_54450; // @[Modules.scala 46:37:@199.4]
  wire [4:0] _T_54451; // @[Modules.scala 46:37:@200.4]
  wire [5:0] _T_54452; // @[Modules.scala 46:47:@201.4]
  wire [4:0] _T_54453; // @[Modules.scala 46:47:@202.4]
  wire [4:0] _T_54454; // @[Modules.scala 46:47:@203.4]
  wire [5:0] _T_54456; // @[Modules.scala 46:37:@205.4]
  wire [4:0] _T_54457; // @[Modules.scala 46:37:@206.4]
  wire [4:0] _T_54458; // @[Modules.scala 46:37:@207.4]
  wire [5:0] _T_54459; // @[Modules.scala 46:47:@208.4]
  wire [4:0] _T_54460; // @[Modules.scala 46:47:@209.4]
  wire [4:0] _T_54461; // @[Modules.scala 46:47:@210.4]
  wire [5:0] _T_54463; // @[Modules.scala 43:37:@212.4]
  wire [4:0] _T_54464; // @[Modules.scala 43:37:@213.4]
  wire [4:0] _T_54465; // @[Modules.scala 43:37:@214.4]
  wire [5:0] _T_54466; // @[Modules.scala 43:47:@215.4]
  wire [4:0] _T_54467; // @[Modules.scala 43:47:@216.4]
  wire [4:0] _T_54468; // @[Modules.scala 43:47:@217.4]
  wire [5:0] _T_54470; // @[Modules.scala 46:37:@219.4]
  wire [4:0] _T_54471; // @[Modules.scala 46:37:@220.4]
  wire [4:0] _T_54472; // @[Modules.scala 46:37:@221.4]
  wire [5:0] _T_54473; // @[Modules.scala 46:47:@222.4]
  wire [4:0] _T_54474; // @[Modules.scala 46:47:@223.4]
  wire [4:0] _T_54475; // @[Modules.scala 46:47:@224.4]
  wire [5:0] _T_54477; // @[Modules.scala 46:37:@226.4]
  wire [4:0] _T_54478; // @[Modules.scala 46:37:@227.4]
  wire [4:0] _T_54479; // @[Modules.scala 46:37:@228.4]
  wire [5:0] _T_54480; // @[Modules.scala 46:47:@229.4]
  wire [4:0] _T_54481; // @[Modules.scala 46:47:@230.4]
  wire [4:0] _T_54482; // @[Modules.scala 46:47:@231.4]
  wire [5:0] _T_54484; // @[Modules.scala 46:37:@233.4]
  wire [4:0] _T_54485; // @[Modules.scala 46:37:@234.4]
  wire [4:0] _T_54486; // @[Modules.scala 46:37:@235.4]
  wire [5:0] _T_54487; // @[Modules.scala 46:47:@236.4]
  wire [4:0] _T_54488; // @[Modules.scala 46:47:@237.4]
  wire [4:0] _T_54489; // @[Modules.scala 46:47:@238.4]
  wire [5:0] _T_54491; // @[Modules.scala 46:37:@240.4]
  wire [4:0] _T_54492; // @[Modules.scala 46:37:@241.4]
  wire [4:0] _T_54493; // @[Modules.scala 46:37:@242.4]
  wire [5:0] _T_54494; // @[Modules.scala 46:47:@243.4]
  wire [4:0] _T_54495; // @[Modules.scala 46:47:@244.4]
  wire [4:0] _T_54496; // @[Modules.scala 46:47:@245.4]
  wire [5:0] _T_54498; // @[Modules.scala 43:37:@247.4]
  wire [4:0] _T_54499; // @[Modules.scala 43:37:@248.4]
  wire [4:0] _T_54500; // @[Modules.scala 43:37:@249.4]
  wire [5:0] _T_54501; // @[Modules.scala 43:47:@250.4]
  wire [4:0] _T_54502; // @[Modules.scala 43:47:@251.4]
  wire [4:0] _T_54503; // @[Modules.scala 43:47:@252.4]
  wire [5:0] _T_54504; // @[Modules.scala 40:46:@254.4]
  wire [4:0] _T_54505; // @[Modules.scala 40:46:@255.4]
  wire [4:0] _T_54506; // @[Modules.scala 40:46:@256.4]
  wire [5:0] _T_54507; // @[Modules.scala 37:46:@258.4]
  wire [4:0] _T_54508; // @[Modules.scala 37:46:@259.4]
  wire [4:0] _T_54509; // @[Modules.scala 37:46:@260.4]
  wire [5:0] _T_54511; // @[Modules.scala 46:37:@262.4]
  wire [4:0] _T_54512; // @[Modules.scala 46:37:@263.4]
  wire [4:0] _T_54513; // @[Modules.scala 46:37:@264.4]
  wire [5:0] _T_54514; // @[Modules.scala 46:47:@265.4]
  wire [4:0] _T_54515; // @[Modules.scala 46:47:@266.4]
  wire [4:0] _T_54516; // @[Modules.scala 46:47:@267.4]
  wire [5:0] _T_54517; // @[Modules.scala 40:46:@269.4]
  wire [4:0] _T_54518; // @[Modules.scala 40:46:@270.4]
  wire [4:0] _T_54519; // @[Modules.scala 40:46:@271.4]
  wire [5:0] _T_54520; // @[Modules.scala 40:46:@273.4]
  wire [4:0] _T_54521; // @[Modules.scala 40:46:@274.4]
  wire [4:0] _T_54522; // @[Modules.scala 40:46:@275.4]
  wire [5:0] _T_54524; // @[Modules.scala 46:37:@277.4]
  wire [4:0] _T_54525; // @[Modules.scala 46:37:@278.4]
  wire [4:0] _T_54526; // @[Modules.scala 46:37:@279.4]
  wire [5:0] _T_54527; // @[Modules.scala 46:47:@280.4]
  wire [4:0] _T_54528; // @[Modules.scala 46:47:@281.4]
  wire [4:0] _T_54529; // @[Modules.scala 46:47:@282.4]
  wire [5:0] _T_54530; // @[Modules.scala 37:46:@284.4]
  wire [4:0] _T_54531; // @[Modules.scala 37:46:@285.4]
  wire [4:0] _T_54532; // @[Modules.scala 37:46:@286.4]
  wire [5:0] _T_54533; // @[Modules.scala 37:46:@288.4]
  wire [4:0] _T_54534; // @[Modules.scala 37:46:@289.4]
  wire [4:0] _T_54535; // @[Modules.scala 37:46:@290.4]
  wire [5:0] _T_54537; // @[Modules.scala 43:37:@292.4]
  wire [4:0] _T_54538; // @[Modules.scala 43:37:@293.4]
  wire [4:0] _T_54539; // @[Modules.scala 43:37:@294.4]
  wire [5:0] _T_54540; // @[Modules.scala 43:47:@295.4]
  wire [4:0] _T_54541; // @[Modules.scala 43:47:@296.4]
  wire [4:0] _T_54542; // @[Modules.scala 43:47:@297.4]
  wire [5:0] _T_54543; // @[Modules.scala 37:46:@299.4]
  wire [4:0] _T_54544; // @[Modules.scala 37:46:@300.4]
  wire [4:0] _T_54545; // @[Modules.scala 37:46:@301.4]
  wire [5:0] _T_54547; // @[Modules.scala 43:37:@303.4]
  wire [4:0] _T_54548; // @[Modules.scala 43:37:@304.4]
  wire [4:0] _T_54549; // @[Modules.scala 43:37:@305.4]
  wire [5:0] _T_54550; // @[Modules.scala 43:47:@306.4]
  wire [4:0] _T_54551; // @[Modules.scala 43:47:@307.4]
  wire [4:0] _T_54552; // @[Modules.scala 43:47:@308.4]
  wire [5:0] _T_54553; // @[Modules.scala 37:46:@310.4]
  wire [4:0] _T_54554; // @[Modules.scala 37:46:@311.4]
  wire [4:0] _T_54555; // @[Modules.scala 37:46:@312.4]
  wire [5:0] _T_54556; // @[Modules.scala 37:46:@314.4]
  wire [4:0] _T_54557; // @[Modules.scala 37:46:@315.4]
  wire [4:0] _T_54558; // @[Modules.scala 37:46:@316.4]
  wire [5:0] _T_54559; // @[Modules.scala 37:46:@318.4]
  wire [4:0] _T_54560; // @[Modules.scala 37:46:@319.4]
  wire [4:0] _T_54561; // @[Modules.scala 37:46:@320.4]
  wire [5:0] _T_54562; // @[Modules.scala 37:46:@322.4]
  wire [4:0] _T_54563; // @[Modules.scala 37:46:@323.4]
  wire [4:0] _T_54564; // @[Modules.scala 37:46:@324.4]
  wire [5:0] _T_54565; // @[Modules.scala 37:46:@326.4]
  wire [4:0] _T_54566; // @[Modules.scala 37:46:@327.4]
  wire [4:0] _T_54567; // @[Modules.scala 37:46:@328.4]
  wire [5:0] _T_54568; // @[Modules.scala 40:46:@330.4]
  wire [4:0] _T_54569; // @[Modules.scala 40:46:@331.4]
  wire [4:0] _T_54570; // @[Modules.scala 40:46:@332.4]
  wire [5:0] _T_54571; // @[Modules.scala 37:46:@334.4]
  wire [4:0] _T_54572; // @[Modules.scala 37:46:@335.4]
  wire [4:0] _T_54573; // @[Modules.scala 37:46:@336.4]
  wire [5:0] _T_54575; // @[Modules.scala 43:37:@338.4]
  wire [4:0] _T_54576; // @[Modules.scala 43:37:@339.4]
  wire [4:0] _T_54577; // @[Modules.scala 43:37:@340.4]
  wire [5:0] _T_54578; // @[Modules.scala 43:47:@341.4]
  wire [4:0] _T_54579; // @[Modules.scala 43:47:@342.4]
  wire [4:0] _T_54580; // @[Modules.scala 43:47:@343.4]
  wire [5:0] _T_54582; // @[Modules.scala 46:37:@345.4]
  wire [4:0] _T_54583; // @[Modules.scala 46:37:@346.4]
  wire [4:0] _T_54584; // @[Modules.scala 46:37:@347.4]
  wire [5:0] _T_54585; // @[Modules.scala 46:47:@348.4]
  wire [4:0] _T_54586; // @[Modules.scala 46:47:@349.4]
  wire [4:0] _T_54587; // @[Modules.scala 46:47:@350.4]
  wire [5:0] _T_54588; // @[Modules.scala 40:46:@352.4]
  wire [4:0] _T_54589; // @[Modules.scala 40:46:@353.4]
  wire [4:0] _T_54590; // @[Modules.scala 40:46:@354.4]
  wire [5:0] _T_54591; // @[Modules.scala 37:46:@356.4]
  wire [4:0] _T_54592; // @[Modules.scala 37:46:@357.4]
  wire [4:0] _T_54593; // @[Modules.scala 37:46:@358.4]
  wire [5:0] _T_54595; // @[Modules.scala 46:37:@360.4]
  wire [4:0] _T_54596; // @[Modules.scala 46:37:@361.4]
  wire [4:0] _T_54597; // @[Modules.scala 46:37:@362.4]
  wire [5:0] _T_54598; // @[Modules.scala 46:47:@363.4]
  wire [4:0] _T_54599; // @[Modules.scala 46:47:@364.4]
  wire [4:0] _T_54600; // @[Modules.scala 46:47:@365.4]
  wire [5:0] _T_54602; // @[Modules.scala 46:37:@367.4]
  wire [4:0] _T_54603; // @[Modules.scala 46:37:@368.4]
  wire [4:0] _T_54604; // @[Modules.scala 46:37:@369.4]
  wire [5:0] _T_54605; // @[Modules.scala 46:47:@370.4]
  wire [4:0] _T_54606; // @[Modules.scala 46:47:@371.4]
  wire [4:0] _T_54607; // @[Modules.scala 46:47:@372.4]
  wire [5:0] _T_54609; // @[Modules.scala 46:37:@374.4]
  wire [4:0] _T_54610; // @[Modules.scala 46:37:@375.4]
  wire [4:0] _T_54611; // @[Modules.scala 46:37:@376.4]
  wire [5:0] _T_54612; // @[Modules.scala 46:47:@377.4]
  wire [4:0] _T_54613; // @[Modules.scala 46:47:@378.4]
  wire [4:0] _T_54614; // @[Modules.scala 46:47:@379.4]
  wire [5:0] _T_54616; // @[Modules.scala 46:37:@381.4]
  wire [4:0] _T_54617; // @[Modules.scala 46:37:@382.4]
  wire [4:0] _T_54618; // @[Modules.scala 46:37:@383.4]
  wire [5:0] _T_54619; // @[Modules.scala 46:47:@384.4]
  wire [4:0] _T_54620; // @[Modules.scala 46:47:@385.4]
  wire [4:0] _T_54621; // @[Modules.scala 46:47:@386.4]
  wire [5:0] _T_54623; // @[Modules.scala 43:37:@388.4]
  wire [4:0] _T_54624; // @[Modules.scala 43:37:@389.4]
  wire [4:0] _T_54625; // @[Modules.scala 43:37:@390.4]
  wire [5:0] _T_54626; // @[Modules.scala 43:47:@391.4]
  wire [4:0] _T_54627; // @[Modules.scala 43:47:@392.4]
  wire [4:0] _T_54628; // @[Modules.scala 43:47:@393.4]
  wire [5:0] _T_54630; // @[Modules.scala 43:37:@395.4]
  wire [4:0] _T_54631; // @[Modules.scala 43:37:@396.4]
  wire [4:0] _T_54632; // @[Modules.scala 43:37:@397.4]
  wire [5:0] _T_54633; // @[Modules.scala 43:47:@398.4]
  wire [4:0] _T_54634; // @[Modules.scala 43:47:@399.4]
  wire [4:0] _T_54635; // @[Modules.scala 43:47:@400.4]
  wire [5:0] _T_54636; // @[Modules.scala 37:46:@402.4]
  wire [4:0] _T_54637; // @[Modules.scala 37:46:@403.4]
  wire [4:0] _T_54638; // @[Modules.scala 37:46:@404.4]
  wire [5:0] _T_54639; // @[Modules.scala 37:46:@406.4]
  wire [4:0] _T_54640; // @[Modules.scala 37:46:@407.4]
  wire [4:0] _T_54641; // @[Modules.scala 37:46:@408.4]
  wire [5:0] _T_54642; // @[Modules.scala 40:46:@410.4]
  wire [4:0] _T_54643; // @[Modules.scala 40:46:@411.4]
  wire [4:0] _T_54644; // @[Modules.scala 40:46:@412.4]
  wire [5:0] _T_54646; // @[Modules.scala 46:37:@414.4]
  wire [4:0] _T_54647; // @[Modules.scala 46:37:@415.4]
  wire [4:0] _T_54648; // @[Modules.scala 46:37:@416.4]
  wire [5:0] _T_54649; // @[Modules.scala 46:47:@417.4]
  wire [4:0] _T_54650; // @[Modules.scala 46:47:@418.4]
  wire [4:0] _T_54651; // @[Modules.scala 46:47:@419.4]
  wire [5:0] _T_54652; // @[Modules.scala 37:46:@421.4]
  wire [4:0] _T_54653; // @[Modules.scala 37:46:@422.4]
  wire [4:0] _T_54654; // @[Modules.scala 37:46:@423.4]
  wire [5:0] _T_54656; // @[Modules.scala 46:37:@425.4]
  wire [4:0] _T_54657; // @[Modules.scala 46:37:@426.4]
  wire [4:0] _T_54658; // @[Modules.scala 46:37:@427.4]
  wire [5:0] _T_54659; // @[Modules.scala 46:47:@428.4]
  wire [4:0] _T_54660; // @[Modules.scala 46:47:@429.4]
  wire [4:0] _T_54661; // @[Modules.scala 46:47:@430.4]
  wire [5:0] _T_54662; // @[Modules.scala 40:46:@432.4]
  wire [4:0] _T_54663; // @[Modules.scala 40:46:@433.4]
  wire [4:0] _T_54664; // @[Modules.scala 40:46:@434.4]
  wire [5:0] _T_54665; // @[Modules.scala 37:46:@436.4]
  wire [4:0] _T_54666; // @[Modules.scala 37:46:@437.4]
  wire [4:0] _T_54667; // @[Modules.scala 37:46:@438.4]
  wire [5:0] _T_54668; // @[Modules.scala 37:46:@440.4]
  wire [4:0] _T_54669; // @[Modules.scala 37:46:@441.4]
  wire [4:0] _T_54670; // @[Modules.scala 37:46:@442.4]
  wire [5:0] _T_54672; // @[Modules.scala 46:37:@444.4]
  wire [4:0] _T_54673; // @[Modules.scala 46:37:@445.4]
  wire [4:0] _T_54674; // @[Modules.scala 46:37:@446.4]
  wire [5:0] _T_54675; // @[Modules.scala 46:47:@447.4]
  wire [4:0] _T_54676; // @[Modules.scala 46:47:@448.4]
  wire [4:0] _T_54677; // @[Modules.scala 46:47:@449.4]
  wire [5:0] _T_54679; // @[Modules.scala 46:37:@451.4]
  wire [4:0] _T_54680; // @[Modules.scala 46:37:@452.4]
  wire [4:0] _T_54681; // @[Modules.scala 46:37:@453.4]
  wire [5:0] _T_54682; // @[Modules.scala 46:47:@454.4]
  wire [4:0] _T_54683; // @[Modules.scala 46:47:@455.4]
  wire [4:0] _T_54684; // @[Modules.scala 46:47:@456.4]
  wire [5:0] _T_54686; // @[Modules.scala 46:37:@458.4]
  wire [4:0] _T_54687; // @[Modules.scala 46:37:@459.4]
  wire [4:0] _T_54688; // @[Modules.scala 46:37:@460.4]
  wire [5:0] _T_54689; // @[Modules.scala 46:47:@461.4]
  wire [4:0] _T_54690; // @[Modules.scala 46:47:@462.4]
  wire [4:0] _T_54691; // @[Modules.scala 46:47:@463.4]
  wire [5:0] _T_54693; // @[Modules.scala 46:37:@465.4]
  wire [4:0] _T_54694; // @[Modules.scala 46:37:@466.4]
  wire [4:0] _T_54695; // @[Modules.scala 46:37:@467.4]
  wire [5:0] _T_54696; // @[Modules.scala 46:47:@468.4]
  wire [4:0] _T_54697; // @[Modules.scala 46:47:@469.4]
  wire [4:0] _T_54698; // @[Modules.scala 46:47:@470.4]
  wire [5:0] _T_54700; // @[Modules.scala 46:37:@472.4]
  wire [4:0] _T_54701; // @[Modules.scala 46:37:@473.4]
  wire [4:0] _T_54702; // @[Modules.scala 46:37:@474.4]
  wire [5:0] _T_54703; // @[Modules.scala 46:47:@475.4]
  wire [4:0] _T_54704; // @[Modules.scala 46:47:@476.4]
  wire [4:0] _T_54705; // @[Modules.scala 46:47:@477.4]
  wire [5:0] _T_54707; // @[Modules.scala 46:37:@479.4]
  wire [4:0] _T_54708; // @[Modules.scala 46:37:@480.4]
  wire [4:0] _T_54709; // @[Modules.scala 46:37:@481.4]
  wire [5:0] _T_54710; // @[Modules.scala 46:47:@482.4]
  wire [4:0] _T_54711; // @[Modules.scala 46:47:@483.4]
  wire [4:0] _T_54712; // @[Modules.scala 46:47:@484.4]
  wire [5:0] _T_54713; // @[Modules.scala 37:46:@486.4]
  wire [4:0] _T_54714; // @[Modules.scala 37:46:@487.4]
  wire [4:0] _T_54715; // @[Modules.scala 37:46:@488.4]
  wire [5:0] _T_54716; // @[Modules.scala 40:46:@490.4]
  wire [4:0] _T_54717; // @[Modules.scala 40:46:@491.4]
  wire [4:0] _T_54718; // @[Modules.scala 40:46:@492.4]
  wire [5:0] _T_54720; // @[Modules.scala 43:37:@494.4]
  wire [4:0] _T_54721; // @[Modules.scala 43:37:@495.4]
  wire [4:0] _T_54722; // @[Modules.scala 43:37:@496.4]
  wire [5:0] _T_54723; // @[Modules.scala 43:47:@497.4]
  wire [4:0] _T_54724; // @[Modules.scala 43:47:@498.4]
  wire [4:0] _T_54725; // @[Modules.scala 43:47:@499.4]
  wire [5:0] _T_54727; // @[Modules.scala 46:37:@501.4]
  wire [4:0] _T_54728; // @[Modules.scala 46:37:@502.4]
  wire [4:0] _T_54729; // @[Modules.scala 46:37:@503.4]
  wire [5:0] _T_54730; // @[Modules.scala 46:47:@504.4]
  wire [4:0] _T_54731; // @[Modules.scala 46:47:@505.4]
  wire [4:0] _T_54732; // @[Modules.scala 46:47:@506.4]
  wire [5:0] _T_54734; // @[Modules.scala 46:37:@508.4]
  wire [4:0] _T_54735; // @[Modules.scala 46:37:@509.4]
  wire [4:0] _T_54736; // @[Modules.scala 46:37:@510.4]
  wire [5:0] _T_54737; // @[Modules.scala 46:47:@511.4]
  wire [4:0] _T_54738; // @[Modules.scala 46:47:@512.4]
  wire [4:0] _T_54739; // @[Modules.scala 46:47:@513.4]
  wire [5:0] _T_54740; // @[Modules.scala 40:46:@515.4]
  wire [4:0] _T_54741; // @[Modules.scala 40:46:@516.4]
  wire [4:0] _T_54742; // @[Modules.scala 40:46:@517.4]
  wire [5:0] _T_54744; // @[Modules.scala 46:37:@519.4]
  wire [4:0] _T_54745; // @[Modules.scala 46:37:@520.4]
  wire [4:0] _T_54746; // @[Modules.scala 46:37:@521.4]
  wire [5:0] _T_54747; // @[Modules.scala 46:47:@522.4]
  wire [4:0] _T_54748; // @[Modules.scala 46:47:@523.4]
  wire [4:0] _T_54749; // @[Modules.scala 46:47:@524.4]
  wire [5:0] _T_54751; // @[Modules.scala 46:37:@526.4]
  wire [4:0] _T_54752; // @[Modules.scala 46:37:@527.4]
  wire [4:0] _T_54753; // @[Modules.scala 46:37:@528.4]
  wire [5:0] _T_54754; // @[Modules.scala 46:47:@529.4]
  wire [4:0] _T_54755; // @[Modules.scala 46:47:@530.4]
  wire [4:0] _T_54756; // @[Modules.scala 46:47:@531.4]
  wire [5:0] _T_54758; // @[Modules.scala 46:37:@533.4]
  wire [4:0] _T_54759; // @[Modules.scala 46:37:@534.4]
  wire [4:0] _T_54760; // @[Modules.scala 46:37:@535.4]
  wire [5:0] _T_54761; // @[Modules.scala 46:47:@536.4]
  wire [4:0] _T_54762; // @[Modules.scala 46:47:@537.4]
  wire [4:0] _T_54763; // @[Modules.scala 46:47:@538.4]
  wire [5:0] _T_54765; // @[Modules.scala 46:37:@540.4]
  wire [4:0] _T_54766; // @[Modules.scala 46:37:@541.4]
  wire [4:0] _T_54767; // @[Modules.scala 46:37:@542.4]
  wire [5:0] _T_54768; // @[Modules.scala 46:47:@543.4]
  wire [4:0] _T_54769; // @[Modules.scala 46:47:@544.4]
  wire [4:0] _T_54770; // @[Modules.scala 46:47:@545.4]
  wire [5:0] _T_54772; // @[Modules.scala 46:37:@547.4]
  wire [4:0] _T_54773; // @[Modules.scala 46:37:@548.4]
  wire [4:0] _T_54774; // @[Modules.scala 46:37:@549.4]
  wire [5:0] _T_54775; // @[Modules.scala 46:47:@550.4]
  wire [4:0] _T_54776; // @[Modules.scala 46:47:@551.4]
  wire [4:0] _T_54777; // @[Modules.scala 46:47:@552.4]
  wire [5:0] _T_54779; // @[Modules.scala 46:37:@554.4]
  wire [4:0] _T_54780; // @[Modules.scala 46:37:@555.4]
  wire [4:0] _T_54781; // @[Modules.scala 46:37:@556.4]
  wire [5:0] _T_54782; // @[Modules.scala 46:47:@557.4]
  wire [4:0] _T_54783; // @[Modules.scala 46:47:@558.4]
  wire [4:0] _T_54784; // @[Modules.scala 46:47:@559.4]
  wire [5:0] _T_54785; // @[Modules.scala 37:46:@561.4]
  wire [4:0] _T_54786; // @[Modules.scala 37:46:@562.4]
  wire [4:0] _T_54787; // @[Modules.scala 37:46:@563.4]
  wire [5:0] _T_54789; // @[Modules.scala 46:37:@565.4]
  wire [4:0] _T_54790; // @[Modules.scala 46:37:@566.4]
  wire [4:0] _T_54791; // @[Modules.scala 46:37:@567.4]
  wire [5:0] _T_54792; // @[Modules.scala 46:47:@568.4]
  wire [4:0] _T_54793; // @[Modules.scala 46:47:@569.4]
  wire [4:0] _T_54794; // @[Modules.scala 46:47:@570.4]
  wire [5:0] _T_54795; // @[Modules.scala 40:46:@572.4]
  wire [4:0] _T_54796; // @[Modules.scala 40:46:@573.4]
  wire [4:0] _T_54797; // @[Modules.scala 40:46:@574.4]
  wire [5:0] _T_54799; // @[Modules.scala 46:37:@576.4]
  wire [4:0] _T_54800; // @[Modules.scala 46:37:@577.4]
  wire [4:0] _T_54801; // @[Modules.scala 46:37:@578.4]
  wire [5:0] _T_54802; // @[Modules.scala 46:47:@579.4]
  wire [4:0] _T_54803; // @[Modules.scala 46:47:@580.4]
  wire [4:0] _T_54804; // @[Modules.scala 46:47:@581.4]
  wire [5:0] _T_54806; // @[Modules.scala 46:37:@583.4]
  wire [4:0] _T_54807; // @[Modules.scala 46:37:@584.4]
  wire [4:0] _T_54808; // @[Modules.scala 46:37:@585.4]
  wire [5:0] _T_54809; // @[Modules.scala 46:47:@586.4]
  wire [4:0] _T_54810; // @[Modules.scala 46:47:@587.4]
  wire [4:0] _T_54811; // @[Modules.scala 46:47:@588.4]
  wire [5:0] _T_54812; // @[Modules.scala 40:46:@590.4]
  wire [4:0] _T_54813; // @[Modules.scala 40:46:@591.4]
  wire [4:0] _T_54814; // @[Modules.scala 40:46:@592.4]
  wire [5:0] _T_54815; // @[Modules.scala 40:46:@594.4]
  wire [4:0] _T_54816; // @[Modules.scala 40:46:@595.4]
  wire [4:0] _T_54817; // @[Modules.scala 40:46:@596.4]
  wire [5:0] _T_54819; // @[Modules.scala 46:37:@598.4]
  wire [4:0] _T_54820; // @[Modules.scala 46:37:@599.4]
  wire [4:0] _T_54821; // @[Modules.scala 46:37:@600.4]
  wire [5:0] _T_54822; // @[Modules.scala 46:47:@601.4]
  wire [4:0] _T_54823; // @[Modules.scala 46:47:@602.4]
  wire [4:0] _T_54824; // @[Modules.scala 46:47:@603.4]
  wire [5:0] _T_54826; // @[Modules.scala 46:37:@605.4]
  wire [4:0] _T_54827; // @[Modules.scala 46:37:@606.4]
  wire [4:0] _T_54828; // @[Modules.scala 46:37:@607.4]
  wire [5:0] _T_54829; // @[Modules.scala 46:47:@608.4]
  wire [4:0] _T_54830; // @[Modules.scala 46:47:@609.4]
  wire [4:0] _T_54831; // @[Modules.scala 46:47:@610.4]
  wire [5:0] _T_54833; // @[Modules.scala 46:37:@612.4]
  wire [4:0] _T_54834; // @[Modules.scala 46:37:@613.4]
  wire [4:0] _T_54835; // @[Modules.scala 46:37:@614.4]
  wire [5:0] _T_54836; // @[Modules.scala 46:47:@615.4]
  wire [4:0] _T_54837; // @[Modules.scala 46:47:@616.4]
  wire [4:0] _T_54838; // @[Modules.scala 46:47:@617.4]
  wire [5:0] _T_54840; // @[Modules.scala 43:37:@619.4]
  wire [4:0] _T_54841; // @[Modules.scala 43:37:@620.4]
  wire [4:0] _T_54842; // @[Modules.scala 43:37:@621.4]
  wire [5:0] _T_54843; // @[Modules.scala 43:47:@622.4]
  wire [4:0] _T_54844; // @[Modules.scala 43:47:@623.4]
  wire [4:0] _T_54845; // @[Modules.scala 43:47:@624.4]
  wire [5:0] _T_54847; // @[Modules.scala 43:37:@626.4]
  wire [4:0] _T_54848; // @[Modules.scala 43:37:@627.4]
  wire [4:0] _T_54849; // @[Modules.scala 43:37:@628.4]
  wire [5:0] _T_54850; // @[Modules.scala 43:47:@629.4]
  wire [4:0] _T_54851; // @[Modules.scala 43:47:@630.4]
  wire [4:0] _T_54852; // @[Modules.scala 43:47:@631.4]
  wire [5:0] _T_54853; // @[Modules.scala 37:46:@633.4]
  wire [4:0] _T_54854; // @[Modules.scala 37:46:@634.4]
  wire [4:0] _T_54855; // @[Modules.scala 37:46:@635.4]
  wire [5:0] _T_54856; // @[Modules.scala 40:46:@637.4]
  wire [4:0] _T_54857; // @[Modules.scala 40:46:@638.4]
  wire [4:0] _T_54858; // @[Modules.scala 40:46:@639.4]
  wire [5:0] _T_54860; // @[Modules.scala 46:37:@641.4]
  wire [4:0] _T_54861; // @[Modules.scala 46:37:@642.4]
  wire [4:0] _T_54862; // @[Modules.scala 46:37:@643.4]
  wire [5:0] _T_54863; // @[Modules.scala 46:47:@644.4]
  wire [4:0] _T_54864; // @[Modules.scala 46:47:@645.4]
  wire [4:0] _T_54865; // @[Modules.scala 46:47:@646.4]
  wire [5:0] _T_54867; // @[Modules.scala 46:37:@648.4]
  wire [4:0] _T_54868; // @[Modules.scala 46:37:@649.4]
  wire [4:0] _T_54869; // @[Modules.scala 46:37:@650.4]
  wire [5:0] _T_54870; // @[Modules.scala 46:47:@651.4]
  wire [4:0] _T_54871; // @[Modules.scala 46:47:@652.4]
  wire [4:0] _T_54872; // @[Modules.scala 46:47:@653.4]
  wire [5:0] _T_54874; // @[Modules.scala 46:37:@655.4]
  wire [4:0] _T_54875; // @[Modules.scala 46:37:@656.4]
  wire [4:0] _T_54876; // @[Modules.scala 46:37:@657.4]
  wire [5:0] _T_54877; // @[Modules.scala 46:47:@658.4]
  wire [4:0] _T_54878; // @[Modules.scala 46:47:@659.4]
  wire [4:0] _T_54879; // @[Modules.scala 46:47:@660.4]
  wire [5:0] _T_54881; // @[Modules.scala 46:37:@662.4]
  wire [4:0] _T_54882; // @[Modules.scala 46:37:@663.4]
  wire [4:0] _T_54883; // @[Modules.scala 46:37:@664.4]
  wire [5:0] _T_54884; // @[Modules.scala 46:47:@665.4]
  wire [4:0] _T_54885; // @[Modules.scala 46:47:@666.4]
  wire [4:0] _T_54886; // @[Modules.scala 46:47:@667.4]
  wire [5:0] _T_54888; // @[Modules.scala 46:37:@669.4]
  wire [4:0] _T_54889; // @[Modules.scala 46:37:@670.4]
  wire [4:0] _T_54890; // @[Modules.scala 46:37:@671.4]
  wire [5:0] _T_54891; // @[Modules.scala 46:47:@672.4]
  wire [4:0] _T_54892; // @[Modules.scala 46:47:@673.4]
  wire [4:0] _T_54893; // @[Modules.scala 46:47:@674.4]
  wire [5:0] _T_54895; // @[Modules.scala 46:37:@676.4]
  wire [4:0] _T_54896; // @[Modules.scala 46:37:@677.4]
  wire [4:0] _T_54897; // @[Modules.scala 46:37:@678.4]
  wire [5:0] _T_54898; // @[Modules.scala 46:47:@679.4]
  wire [4:0] _T_54899; // @[Modules.scala 46:47:@680.4]
  wire [4:0] _T_54900; // @[Modules.scala 46:47:@681.4]
  wire [5:0] _T_54902; // @[Modules.scala 46:37:@683.4]
  wire [4:0] _T_54903; // @[Modules.scala 46:37:@684.4]
  wire [4:0] _T_54904; // @[Modules.scala 46:37:@685.4]
  wire [5:0] _T_54905; // @[Modules.scala 46:47:@686.4]
  wire [4:0] _T_54906; // @[Modules.scala 46:47:@687.4]
  wire [4:0] _T_54907; // @[Modules.scala 46:47:@688.4]
  wire [5:0] _T_54909; // @[Modules.scala 46:37:@690.4]
  wire [4:0] _T_54910; // @[Modules.scala 46:37:@691.4]
  wire [4:0] _T_54911; // @[Modules.scala 46:37:@692.4]
  wire [5:0] _T_54912; // @[Modules.scala 46:47:@693.4]
  wire [4:0] _T_54913; // @[Modules.scala 46:47:@694.4]
  wire [4:0] _T_54914; // @[Modules.scala 46:47:@695.4]
  wire [5:0] _T_54916; // @[Modules.scala 46:37:@697.4]
  wire [4:0] _T_54917; // @[Modules.scala 46:37:@698.4]
  wire [4:0] _T_54918; // @[Modules.scala 46:37:@699.4]
  wire [5:0] _T_54919; // @[Modules.scala 46:47:@700.4]
  wire [4:0] _T_54920; // @[Modules.scala 46:47:@701.4]
  wire [4:0] _T_54921; // @[Modules.scala 46:47:@702.4]
  wire [5:0] _T_54923; // @[Modules.scala 46:37:@704.4]
  wire [4:0] _T_54924; // @[Modules.scala 46:37:@705.4]
  wire [4:0] _T_54925; // @[Modules.scala 46:37:@706.4]
  wire [5:0] _T_54926; // @[Modules.scala 46:47:@707.4]
  wire [4:0] _T_54927; // @[Modules.scala 46:47:@708.4]
  wire [4:0] _T_54928; // @[Modules.scala 46:47:@709.4]
  wire [5:0] _T_54930; // @[Modules.scala 46:37:@711.4]
  wire [4:0] _T_54931; // @[Modules.scala 46:37:@712.4]
  wire [4:0] _T_54932; // @[Modules.scala 46:37:@713.4]
  wire [5:0] _T_54933; // @[Modules.scala 46:47:@714.4]
  wire [4:0] _T_54934; // @[Modules.scala 46:47:@715.4]
  wire [4:0] _T_54935; // @[Modules.scala 46:47:@716.4]
  wire [5:0] _T_54937; // @[Modules.scala 43:37:@718.4]
  wire [4:0] _T_54938; // @[Modules.scala 43:37:@719.4]
  wire [4:0] _T_54939; // @[Modules.scala 43:37:@720.4]
  wire [5:0] _T_54940; // @[Modules.scala 43:47:@721.4]
  wire [4:0] _T_54941; // @[Modules.scala 43:47:@722.4]
  wire [4:0] _T_54942; // @[Modules.scala 43:47:@723.4]
  wire [5:0] _T_54944; // @[Modules.scala 46:37:@725.4]
  wire [4:0] _T_54945; // @[Modules.scala 46:37:@726.4]
  wire [4:0] _T_54946; // @[Modules.scala 46:37:@727.4]
  wire [5:0] _T_54947; // @[Modules.scala 46:47:@728.4]
  wire [4:0] _T_54948; // @[Modules.scala 46:47:@729.4]
  wire [4:0] _T_54949; // @[Modules.scala 46:47:@730.4]
  wire [5:0] _T_54951; // @[Modules.scala 46:37:@732.4]
  wire [4:0] _T_54952; // @[Modules.scala 46:37:@733.4]
  wire [4:0] _T_54953; // @[Modules.scala 46:37:@734.4]
  wire [5:0] _T_54954; // @[Modules.scala 46:47:@735.4]
  wire [4:0] _T_54955; // @[Modules.scala 46:47:@736.4]
  wire [4:0] _T_54956; // @[Modules.scala 46:47:@737.4]
  wire [5:0] _T_54958; // @[Modules.scala 46:37:@739.4]
  wire [4:0] _T_54959; // @[Modules.scala 46:37:@740.4]
  wire [4:0] _T_54960; // @[Modules.scala 46:37:@741.4]
  wire [5:0] _T_54961; // @[Modules.scala 46:47:@742.4]
  wire [4:0] _T_54962; // @[Modules.scala 46:47:@743.4]
  wire [4:0] _T_54963; // @[Modules.scala 46:47:@744.4]
  wire [5:0] _T_54965; // @[Modules.scala 46:37:@746.4]
  wire [4:0] _T_54966; // @[Modules.scala 46:37:@747.4]
  wire [4:0] _T_54967; // @[Modules.scala 46:37:@748.4]
  wire [5:0] _T_54968; // @[Modules.scala 46:47:@749.4]
  wire [4:0] _T_54969; // @[Modules.scala 46:47:@750.4]
  wire [4:0] _T_54970; // @[Modules.scala 46:47:@751.4]
  wire [5:0] _T_54972; // @[Modules.scala 46:37:@753.4]
  wire [4:0] _T_54973; // @[Modules.scala 46:37:@754.4]
  wire [4:0] _T_54974; // @[Modules.scala 46:37:@755.4]
  wire [5:0] _T_54975; // @[Modules.scala 46:47:@756.4]
  wire [4:0] _T_54976; // @[Modules.scala 46:47:@757.4]
  wire [4:0] _T_54977; // @[Modules.scala 46:47:@758.4]
  wire [5:0] _T_54979; // @[Modules.scala 46:37:@760.4]
  wire [4:0] _T_54980; // @[Modules.scala 46:37:@761.4]
  wire [4:0] _T_54981; // @[Modules.scala 46:37:@762.4]
  wire [5:0] _T_54982; // @[Modules.scala 46:47:@763.4]
  wire [4:0] _T_54983; // @[Modules.scala 46:47:@764.4]
  wire [4:0] _T_54984; // @[Modules.scala 46:47:@765.4]
  wire [5:0] _T_54986; // @[Modules.scala 46:37:@767.4]
  wire [4:0] _T_54987; // @[Modules.scala 46:37:@768.4]
  wire [4:0] _T_54988; // @[Modules.scala 46:37:@769.4]
  wire [5:0] _T_54989; // @[Modules.scala 46:47:@770.4]
  wire [4:0] _T_54990; // @[Modules.scala 46:47:@771.4]
  wire [4:0] _T_54991; // @[Modules.scala 46:47:@772.4]
  wire [5:0] _T_54993; // @[Modules.scala 46:37:@774.4]
  wire [4:0] _T_54994; // @[Modules.scala 46:37:@775.4]
  wire [4:0] _T_54995; // @[Modules.scala 46:37:@776.4]
  wire [5:0] _T_54996; // @[Modules.scala 46:47:@777.4]
  wire [4:0] _T_54997; // @[Modules.scala 46:47:@778.4]
  wire [4:0] _T_54998; // @[Modules.scala 46:47:@779.4]
  wire [5:0] _T_55000; // @[Modules.scala 46:37:@781.4]
  wire [4:0] _T_55001; // @[Modules.scala 46:37:@782.4]
  wire [4:0] _T_55002; // @[Modules.scala 46:37:@783.4]
  wire [5:0] _T_55003; // @[Modules.scala 46:47:@784.4]
  wire [4:0] _T_55004; // @[Modules.scala 46:47:@785.4]
  wire [4:0] _T_55005; // @[Modules.scala 46:47:@786.4]
  wire [5:0] _T_55007; // @[Modules.scala 46:37:@788.4]
  wire [4:0] _T_55008; // @[Modules.scala 46:37:@789.4]
  wire [4:0] _T_55009; // @[Modules.scala 46:37:@790.4]
  wire [5:0] _T_55010; // @[Modules.scala 46:47:@791.4]
  wire [4:0] _T_55011; // @[Modules.scala 46:47:@792.4]
  wire [4:0] _T_55012; // @[Modules.scala 46:47:@793.4]
  wire [5:0] _T_55014; // @[Modules.scala 46:37:@795.4]
  wire [4:0] _T_55015; // @[Modules.scala 46:37:@796.4]
  wire [4:0] _T_55016; // @[Modules.scala 46:37:@797.4]
  wire [5:0] _T_55017; // @[Modules.scala 46:47:@798.4]
  wire [4:0] _T_55018; // @[Modules.scala 46:47:@799.4]
  wire [4:0] _T_55019; // @[Modules.scala 46:47:@800.4]
  wire [5:0] _T_55021; // @[Modules.scala 46:37:@802.4]
  wire [4:0] _T_55022; // @[Modules.scala 46:37:@803.4]
  wire [4:0] _T_55023; // @[Modules.scala 46:37:@804.4]
  wire [5:0] _T_55024; // @[Modules.scala 46:47:@805.4]
  wire [4:0] _T_55025; // @[Modules.scala 46:47:@806.4]
  wire [4:0] _T_55026; // @[Modules.scala 46:47:@807.4]
  wire [5:0] _T_55027; // @[Modules.scala 40:46:@809.4]
  wire [4:0] _T_55028; // @[Modules.scala 40:46:@810.4]
  wire [4:0] _T_55029; // @[Modules.scala 40:46:@811.4]
  wire [5:0] _T_55031; // @[Modules.scala 46:37:@813.4]
  wire [4:0] _T_55032; // @[Modules.scala 46:37:@814.4]
  wire [4:0] _T_55033; // @[Modules.scala 46:37:@815.4]
  wire [5:0] _T_55034; // @[Modules.scala 46:47:@816.4]
  wire [4:0] _T_55035; // @[Modules.scala 46:47:@817.4]
  wire [4:0] _T_55036; // @[Modules.scala 46:47:@818.4]
  wire [5:0] _T_55038; // @[Modules.scala 46:37:@820.4]
  wire [4:0] _T_55039; // @[Modules.scala 46:37:@821.4]
  wire [4:0] _T_55040; // @[Modules.scala 46:37:@822.4]
  wire [5:0] _T_55041; // @[Modules.scala 46:47:@823.4]
  wire [4:0] _T_55042; // @[Modules.scala 46:47:@824.4]
  wire [4:0] _T_55043; // @[Modules.scala 46:47:@825.4]
  wire [5:0] _T_55045; // @[Modules.scala 46:37:@827.4]
  wire [4:0] _T_55046; // @[Modules.scala 46:37:@828.4]
  wire [4:0] _T_55047; // @[Modules.scala 46:37:@829.4]
  wire [5:0] _T_55048; // @[Modules.scala 46:47:@830.4]
  wire [4:0] _T_55049; // @[Modules.scala 46:47:@831.4]
  wire [4:0] _T_55050; // @[Modules.scala 46:47:@832.4]
  wire [5:0] _T_55052; // @[Modules.scala 46:37:@834.4]
  wire [4:0] _T_55053; // @[Modules.scala 46:37:@835.4]
  wire [4:0] _T_55054; // @[Modules.scala 46:37:@836.4]
  wire [5:0] _T_55055; // @[Modules.scala 46:47:@837.4]
  wire [4:0] _T_55056; // @[Modules.scala 46:47:@838.4]
  wire [4:0] _T_55057; // @[Modules.scala 46:47:@839.4]
  wire [5:0] _T_55059; // @[Modules.scala 46:37:@841.4]
  wire [4:0] _T_55060; // @[Modules.scala 46:37:@842.4]
  wire [4:0] _T_55061; // @[Modules.scala 46:37:@843.4]
  wire [5:0] _T_55062; // @[Modules.scala 46:47:@844.4]
  wire [4:0] _T_55063; // @[Modules.scala 46:47:@845.4]
  wire [4:0] _T_55064; // @[Modules.scala 46:47:@846.4]
  wire [5:0] _T_55066; // @[Modules.scala 46:37:@848.4]
  wire [4:0] _T_55067; // @[Modules.scala 46:37:@849.4]
  wire [4:0] _T_55068; // @[Modules.scala 46:37:@850.4]
  wire [5:0] _T_55069; // @[Modules.scala 46:47:@851.4]
  wire [4:0] _T_55070; // @[Modules.scala 46:47:@852.4]
  wire [4:0] _T_55071; // @[Modules.scala 46:47:@853.4]
  wire [5:0] _T_55073; // @[Modules.scala 46:37:@855.4]
  wire [4:0] _T_55074; // @[Modules.scala 46:37:@856.4]
  wire [4:0] _T_55075; // @[Modules.scala 46:37:@857.4]
  wire [5:0] _T_55076; // @[Modules.scala 46:47:@858.4]
  wire [4:0] _T_55077; // @[Modules.scala 46:47:@859.4]
  wire [4:0] _T_55078; // @[Modules.scala 46:47:@860.4]
  wire [5:0] _T_55080; // @[Modules.scala 46:37:@862.4]
  wire [4:0] _T_55081; // @[Modules.scala 46:37:@863.4]
  wire [4:0] _T_55082; // @[Modules.scala 46:37:@864.4]
  wire [5:0] _T_55083; // @[Modules.scala 46:47:@865.4]
  wire [4:0] _T_55084; // @[Modules.scala 46:47:@866.4]
  wire [4:0] _T_55085; // @[Modules.scala 46:47:@867.4]
  wire [5:0] _T_55087; // @[Modules.scala 46:37:@869.4]
  wire [4:0] _T_55088; // @[Modules.scala 46:37:@870.4]
  wire [4:0] _T_55089; // @[Modules.scala 46:37:@871.4]
  wire [5:0] _T_55090; // @[Modules.scala 46:47:@872.4]
  wire [4:0] _T_55091; // @[Modules.scala 46:47:@873.4]
  wire [4:0] _T_55092; // @[Modules.scala 46:47:@874.4]
  wire [5:0] _T_55094; // @[Modules.scala 46:37:@876.4]
  wire [4:0] _T_55095; // @[Modules.scala 46:37:@877.4]
  wire [4:0] _T_55096; // @[Modules.scala 46:37:@878.4]
  wire [5:0] _T_55097; // @[Modules.scala 46:47:@879.4]
  wire [4:0] _T_55098; // @[Modules.scala 46:47:@880.4]
  wire [4:0] _T_55099; // @[Modules.scala 46:47:@881.4]
  wire [5:0] _T_55101; // @[Modules.scala 46:37:@883.4]
  wire [4:0] _T_55102; // @[Modules.scala 46:37:@884.4]
  wire [4:0] _T_55103; // @[Modules.scala 46:37:@885.4]
  wire [5:0] _T_55104; // @[Modules.scala 46:47:@886.4]
  wire [4:0] _T_55105; // @[Modules.scala 46:47:@887.4]
  wire [4:0] _T_55106; // @[Modules.scala 46:47:@888.4]
  wire [5:0] _T_55108; // @[Modules.scala 46:37:@890.4]
  wire [4:0] _T_55109; // @[Modules.scala 46:37:@891.4]
  wire [4:0] _T_55110; // @[Modules.scala 46:37:@892.4]
  wire [5:0] _T_55111; // @[Modules.scala 46:47:@893.4]
  wire [4:0] _T_55112; // @[Modules.scala 46:47:@894.4]
  wire [4:0] _T_55113; // @[Modules.scala 46:47:@895.4]
  wire [5:0] _T_55115; // @[Modules.scala 43:37:@897.4]
  wire [4:0] _T_55116; // @[Modules.scala 43:37:@898.4]
  wire [4:0] _T_55117; // @[Modules.scala 43:37:@899.4]
  wire [5:0] _T_55118; // @[Modules.scala 43:47:@900.4]
  wire [4:0] _T_55119; // @[Modules.scala 43:47:@901.4]
  wire [4:0] _T_55120; // @[Modules.scala 43:47:@902.4]
  wire [5:0] _T_55122; // @[Modules.scala 46:37:@904.4]
  wire [4:0] _T_55123; // @[Modules.scala 46:37:@905.4]
  wire [4:0] _T_55124; // @[Modules.scala 46:37:@906.4]
  wire [5:0] _T_55125; // @[Modules.scala 46:47:@907.4]
  wire [4:0] _T_55126; // @[Modules.scala 46:47:@908.4]
  wire [4:0] _T_55127; // @[Modules.scala 46:47:@909.4]
  wire [5:0] _T_55129; // @[Modules.scala 46:37:@911.4]
  wire [4:0] _T_55130; // @[Modules.scala 46:37:@912.4]
  wire [4:0] _T_55131; // @[Modules.scala 46:37:@913.4]
  wire [5:0] _T_55132; // @[Modules.scala 46:47:@914.4]
  wire [4:0] _T_55133; // @[Modules.scala 46:47:@915.4]
  wire [4:0] _T_55134; // @[Modules.scala 46:47:@916.4]
  wire [5:0] _T_55136; // @[Modules.scala 46:37:@918.4]
  wire [4:0] _T_55137; // @[Modules.scala 46:37:@919.4]
  wire [4:0] _T_55138; // @[Modules.scala 46:37:@920.4]
  wire [5:0] _T_55139; // @[Modules.scala 46:47:@921.4]
  wire [4:0] _T_55140; // @[Modules.scala 46:47:@922.4]
  wire [4:0] _T_55141; // @[Modules.scala 46:47:@923.4]
  wire [5:0] _T_55143; // @[Modules.scala 46:37:@925.4]
  wire [4:0] _T_55144; // @[Modules.scala 46:37:@926.4]
  wire [4:0] _T_55145; // @[Modules.scala 46:37:@927.4]
  wire [5:0] _T_55146; // @[Modules.scala 46:47:@928.4]
  wire [4:0] _T_55147; // @[Modules.scala 46:47:@929.4]
  wire [4:0] _T_55148; // @[Modules.scala 46:47:@930.4]
  wire [5:0] _T_55150; // @[Modules.scala 46:37:@932.4]
  wire [4:0] _T_55151; // @[Modules.scala 46:37:@933.4]
  wire [4:0] _T_55152; // @[Modules.scala 46:37:@934.4]
  wire [5:0] _T_55153; // @[Modules.scala 46:47:@935.4]
  wire [4:0] _T_55154; // @[Modules.scala 46:47:@936.4]
  wire [4:0] _T_55155; // @[Modules.scala 46:47:@937.4]
  wire [5:0] _T_55157; // @[Modules.scala 46:37:@939.4]
  wire [4:0] _T_55158; // @[Modules.scala 46:37:@940.4]
  wire [4:0] _T_55159; // @[Modules.scala 46:37:@941.4]
  wire [5:0] _T_55160; // @[Modules.scala 46:47:@942.4]
  wire [4:0] _T_55161; // @[Modules.scala 46:47:@943.4]
  wire [4:0] _T_55162; // @[Modules.scala 46:47:@944.4]
  wire [5:0] _T_55164; // @[Modules.scala 46:37:@946.4]
  wire [4:0] _T_55165; // @[Modules.scala 46:37:@947.4]
  wire [4:0] _T_55166; // @[Modules.scala 46:37:@948.4]
  wire [5:0] _T_55167; // @[Modules.scala 46:47:@949.4]
  wire [4:0] _T_55168; // @[Modules.scala 46:47:@950.4]
  wire [4:0] _T_55169; // @[Modules.scala 46:47:@951.4]
  wire [5:0] _T_55171; // @[Modules.scala 46:37:@953.4]
  wire [4:0] _T_55172; // @[Modules.scala 46:37:@954.4]
  wire [4:0] _T_55173; // @[Modules.scala 46:37:@955.4]
  wire [5:0] _T_55174; // @[Modules.scala 46:47:@956.4]
  wire [4:0] _T_55175; // @[Modules.scala 46:47:@957.4]
  wire [4:0] _T_55176; // @[Modules.scala 46:47:@958.4]
  wire [5:0] _T_55178; // @[Modules.scala 46:37:@960.4]
  wire [4:0] _T_55179; // @[Modules.scala 46:37:@961.4]
  wire [4:0] _T_55180; // @[Modules.scala 46:37:@962.4]
  wire [5:0] _T_55181; // @[Modules.scala 46:47:@963.4]
  wire [4:0] _T_55182; // @[Modules.scala 46:47:@964.4]
  wire [4:0] _T_55183; // @[Modules.scala 46:47:@965.4]
  wire [5:0] _T_55185; // @[Modules.scala 46:37:@967.4]
  wire [4:0] _T_55186; // @[Modules.scala 46:37:@968.4]
  wire [4:0] _T_55187; // @[Modules.scala 46:37:@969.4]
  wire [5:0] _T_55188; // @[Modules.scala 46:47:@970.4]
  wire [4:0] _T_55189; // @[Modules.scala 46:47:@971.4]
  wire [4:0] _T_55190; // @[Modules.scala 46:47:@972.4]
  wire [5:0] _T_55192; // @[Modules.scala 46:37:@974.4]
  wire [4:0] _T_55193; // @[Modules.scala 46:37:@975.4]
  wire [4:0] _T_55194; // @[Modules.scala 46:37:@976.4]
  wire [5:0] _T_55195; // @[Modules.scala 46:47:@977.4]
  wire [4:0] _T_55196; // @[Modules.scala 46:47:@978.4]
  wire [4:0] _T_55197; // @[Modules.scala 46:47:@979.4]
  wire [5:0] _T_55199; // @[Modules.scala 46:37:@981.4]
  wire [4:0] _T_55200; // @[Modules.scala 46:37:@982.4]
  wire [4:0] _T_55201; // @[Modules.scala 46:37:@983.4]
  wire [5:0] _T_55202; // @[Modules.scala 46:47:@984.4]
  wire [4:0] _T_55203; // @[Modules.scala 46:47:@985.4]
  wire [4:0] _T_55204; // @[Modules.scala 46:47:@986.4]
  wire [5:0] _T_55206; // @[Modules.scala 43:37:@988.4]
  wire [4:0] _T_55207; // @[Modules.scala 43:37:@989.4]
  wire [4:0] _T_55208; // @[Modules.scala 43:37:@990.4]
  wire [5:0] _T_55209; // @[Modules.scala 43:47:@991.4]
  wire [4:0] _T_55210; // @[Modules.scala 43:47:@992.4]
  wire [4:0] _T_55211; // @[Modules.scala 43:47:@993.4]
  wire [5:0] _T_55212; // @[Modules.scala 37:46:@995.4]
  wire [4:0] _T_55213; // @[Modules.scala 37:46:@996.4]
  wire [4:0] _T_55214; // @[Modules.scala 37:46:@997.4]
  wire [5:0] _T_55215; // @[Modules.scala 37:46:@999.4]
  wire [4:0] _T_55216; // @[Modules.scala 37:46:@1000.4]
  wire [4:0] _T_55217; // @[Modules.scala 37:46:@1001.4]
  wire [5:0] _T_55219; // @[Modules.scala 46:37:@1003.4]
  wire [4:0] _T_55220; // @[Modules.scala 46:37:@1004.4]
  wire [4:0] _T_55221; // @[Modules.scala 46:37:@1005.4]
  wire [5:0] _T_55222; // @[Modules.scala 46:47:@1006.4]
  wire [4:0] _T_55223; // @[Modules.scala 46:47:@1007.4]
  wire [4:0] _T_55224; // @[Modules.scala 46:47:@1008.4]
  wire [5:0] _T_55226; // @[Modules.scala 46:37:@1010.4]
  wire [4:0] _T_55227; // @[Modules.scala 46:37:@1011.4]
  wire [4:0] _T_55228; // @[Modules.scala 46:37:@1012.4]
  wire [5:0] _T_55229; // @[Modules.scala 46:47:@1013.4]
  wire [4:0] _T_55230; // @[Modules.scala 46:47:@1014.4]
  wire [4:0] _T_55231; // @[Modules.scala 46:47:@1015.4]
  wire [5:0] _T_55233; // @[Modules.scala 43:37:@1017.4]
  wire [4:0] _T_55234; // @[Modules.scala 43:37:@1018.4]
  wire [4:0] _T_55235; // @[Modules.scala 43:37:@1019.4]
  wire [5:0] _T_55236; // @[Modules.scala 43:47:@1020.4]
  wire [4:0] _T_55237; // @[Modules.scala 43:47:@1021.4]
  wire [4:0] _T_55238; // @[Modules.scala 43:47:@1022.4]
  wire [5:0] _T_55240; // @[Modules.scala 46:37:@1024.4]
  wire [4:0] _T_55241; // @[Modules.scala 46:37:@1025.4]
  wire [4:0] _T_55242; // @[Modules.scala 46:37:@1026.4]
  wire [5:0] _T_55243; // @[Modules.scala 46:47:@1027.4]
  wire [4:0] _T_55244; // @[Modules.scala 46:47:@1028.4]
  wire [4:0] _T_55245; // @[Modules.scala 46:47:@1029.4]
  wire [5:0] _T_55246; // @[Modules.scala 37:46:@1031.4]
  wire [4:0] _T_55247; // @[Modules.scala 37:46:@1032.4]
  wire [4:0] _T_55248; // @[Modules.scala 37:46:@1033.4]
  wire [5:0] _T_55250; // @[Modules.scala 46:37:@1035.4]
  wire [4:0] _T_55251; // @[Modules.scala 46:37:@1036.4]
  wire [4:0] _T_55252; // @[Modules.scala 46:37:@1037.4]
  wire [5:0] _T_55253; // @[Modules.scala 46:47:@1038.4]
  wire [4:0] _T_55254; // @[Modules.scala 46:47:@1039.4]
  wire [4:0] _T_55255; // @[Modules.scala 46:47:@1040.4]
  wire [5:0] _T_55257; // @[Modules.scala 46:37:@1042.4]
  wire [4:0] _T_55258; // @[Modules.scala 46:37:@1043.4]
  wire [4:0] _T_55259; // @[Modules.scala 46:37:@1044.4]
  wire [5:0] _T_55260; // @[Modules.scala 46:47:@1045.4]
  wire [4:0] _T_55261; // @[Modules.scala 46:47:@1046.4]
  wire [4:0] _T_55262; // @[Modules.scala 46:47:@1047.4]
  wire [5:0] _T_55264; // @[Modules.scala 43:37:@1049.4]
  wire [4:0] _T_55265; // @[Modules.scala 43:37:@1050.4]
  wire [4:0] _T_55266; // @[Modules.scala 43:37:@1051.4]
  wire [5:0] _T_55267; // @[Modules.scala 43:47:@1052.4]
  wire [4:0] _T_55268; // @[Modules.scala 43:47:@1053.4]
  wire [4:0] _T_55269; // @[Modules.scala 43:47:@1054.4]
  wire [5:0] _T_55270; // @[Modules.scala 40:46:@1056.4]
  wire [4:0] _T_55271; // @[Modules.scala 40:46:@1057.4]
  wire [4:0] _T_55272; // @[Modules.scala 40:46:@1058.4]
  wire [5:0] _T_55274; // @[Modules.scala 46:37:@1060.4]
  wire [4:0] _T_55275; // @[Modules.scala 46:37:@1061.4]
  wire [4:0] _T_55276; // @[Modules.scala 46:37:@1062.4]
  wire [5:0] _T_55277; // @[Modules.scala 46:47:@1063.4]
  wire [4:0] _T_55278; // @[Modules.scala 46:47:@1064.4]
  wire [4:0] _T_55279; // @[Modules.scala 46:47:@1065.4]
  wire [5:0] _T_55281; // @[Modules.scala 43:37:@1067.4]
  wire [4:0] _T_55282; // @[Modules.scala 43:37:@1068.4]
  wire [4:0] _T_55283; // @[Modules.scala 43:37:@1069.4]
  wire [5:0] _T_55284; // @[Modules.scala 43:47:@1070.4]
  wire [4:0] _T_55285; // @[Modules.scala 43:47:@1071.4]
  wire [4:0] _T_55286; // @[Modules.scala 43:47:@1072.4]
  wire [5:0] _T_55287; // @[Modules.scala 37:46:@1074.4]
  wire [4:0] _T_55288; // @[Modules.scala 37:46:@1075.4]
  wire [4:0] _T_55289; // @[Modules.scala 37:46:@1076.4]
  wire [5:0] _T_55290; // @[Modules.scala 37:46:@1078.4]
  wire [4:0] _T_55291; // @[Modules.scala 37:46:@1079.4]
  wire [4:0] _T_55292; // @[Modules.scala 37:46:@1080.4]
  wire [5:0] _T_55293; // @[Modules.scala 37:46:@1082.4]
  wire [4:0] _T_55294; // @[Modules.scala 37:46:@1083.4]
  wire [4:0] _T_55295; // @[Modules.scala 37:46:@1084.4]
  wire [5:0] _T_55296; // @[Modules.scala 37:46:@1086.4]
  wire [4:0] _T_55297; // @[Modules.scala 37:46:@1087.4]
  wire [4:0] _T_55298; // @[Modules.scala 37:46:@1088.4]
  wire [5:0] _T_55299; // @[Modules.scala 37:46:@1090.4]
  wire [4:0] _T_55300; // @[Modules.scala 37:46:@1091.4]
  wire [4:0] _T_55301; // @[Modules.scala 37:46:@1092.4]
  wire [5:0] _T_55302; // @[Modules.scala 37:46:@1094.4]
  wire [4:0] _T_55303; // @[Modules.scala 37:46:@1095.4]
  wire [4:0] _T_55304; // @[Modules.scala 37:46:@1096.4]
  wire [5:0] _T_55305; // @[Modules.scala 37:46:@1098.4]
  wire [4:0] _T_55306; // @[Modules.scala 37:46:@1099.4]
  wire [4:0] _T_55307; // @[Modules.scala 37:46:@1100.4]
  wire [5:0] _T_55308; // @[Modules.scala 37:46:@1102.4]
  wire [4:0] _T_55309; // @[Modules.scala 37:46:@1103.4]
  wire [4:0] _T_55310; // @[Modules.scala 37:46:@1104.4]
  wire [5:0] _T_55311; // @[Modules.scala 37:46:@1106.4]
  wire [4:0] _T_55312; // @[Modules.scala 37:46:@1107.4]
  wire [4:0] _T_55313; // @[Modules.scala 37:46:@1108.4]
  wire [5:0] _T_55315; // @[Modules.scala 46:37:@1110.4]
  wire [4:0] _T_55316; // @[Modules.scala 46:37:@1111.4]
  wire [4:0] _T_55317; // @[Modules.scala 46:37:@1112.4]
  wire [5:0] _T_55318; // @[Modules.scala 46:47:@1113.4]
  wire [4:0] _T_55319; // @[Modules.scala 46:47:@1114.4]
  wire [4:0] _T_55320; // @[Modules.scala 46:47:@1115.4]
  wire [5:0] _T_55322; // @[Modules.scala 43:37:@1117.4]
  wire [4:0] _T_55323; // @[Modules.scala 43:37:@1118.4]
  wire [4:0] _T_55324; // @[Modules.scala 43:37:@1119.4]
  wire [5:0] _T_55325; // @[Modules.scala 43:47:@1120.4]
  wire [4:0] _T_55326; // @[Modules.scala 43:47:@1121.4]
  wire [4:0] _T_55327; // @[Modules.scala 43:47:@1122.4]
  wire [5:0] _T_55329; // @[Modules.scala 46:37:@1124.4]
  wire [4:0] _T_55330; // @[Modules.scala 46:37:@1125.4]
  wire [4:0] _T_55331; // @[Modules.scala 46:37:@1126.4]
  wire [5:0] _T_55332; // @[Modules.scala 46:47:@1127.4]
  wire [4:0] _T_55333; // @[Modules.scala 46:47:@1128.4]
  wire [4:0] _T_55334; // @[Modules.scala 46:47:@1129.4]
  wire [5:0] _T_55336; // @[Modules.scala 46:37:@1131.4]
  wire [4:0] _T_55337; // @[Modules.scala 46:37:@1132.4]
  wire [4:0] _T_55338; // @[Modules.scala 46:37:@1133.4]
  wire [5:0] _T_55339; // @[Modules.scala 46:47:@1134.4]
  wire [4:0] _T_55340; // @[Modules.scala 46:47:@1135.4]
  wire [4:0] _T_55341; // @[Modules.scala 46:47:@1136.4]
  wire [5:0] _T_55342; // @[Modules.scala 37:46:@1138.4]
  wire [4:0] _T_55343; // @[Modules.scala 37:46:@1139.4]
  wire [4:0] _T_55344; // @[Modules.scala 37:46:@1140.4]
  wire [5:0] _T_55345; // @[Modules.scala 37:46:@1142.4]
  wire [4:0] _T_55346; // @[Modules.scala 37:46:@1143.4]
  wire [4:0] _T_55347; // @[Modules.scala 37:46:@1144.4]
  wire [5:0] _T_55348; // @[Modules.scala 37:46:@1146.4]
  wire [4:0] _T_55349; // @[Modules.scala 37:46:@1147.4]
  wire [4:0] _T_55350; // @[Modules.scala 37:46:@1148.4]
  wire [5:0] _T_55351; // @[Modules.scala 37:46:@1150.4]
  wire [4:0] _T_55352; // @[Modules.scala 37:46:@1151.4]
  wire [4:0] _T_55353; // @[Modules.scala 37:46:@1152.4]
  wire [5:0] _T_55354; // @[Modules.scala 37:46:@1154.4]
  wire [4:0] _T_55355; // @[Modules.scala 37:46:@1155.4]
  wire [4:0] _T_55356; // @[Modules.scala 37:46:@1156.4]
  wire [5:0] _T_55357; // @[Modules.scala 37:46:@1158.4]
  wire [4:0] _T_55358; // @[Modules.scala 37:46:@1159.4]
  wire [4:0] _T_55359; // @[Modules.scala 37:46:@1160.4]
  wire [5:0] _T_55360; // @[Modules.scala 37:46:@1162.4]
  wire [4:0] _T_55361; // @[Modules.scala 37:46:@1163.4]
  wire [4:0] _T_55362; // @[Modules.scala 37:46:@1164.4]
  wire [5:0] _T_55363; // @[Modules.scala 37:46:@1166.4]
  wire [4:0] _T_55364; // @[Modules.scala 37:46:@1167.4]
  wire [4:0] _T_55365; // @[Modules.scala 37:46:@1168.4]
  wire [5:0] _T_55367; // @[Modules.scala 43:37:@1170.4]
  wire [4:0] _T_55368; // @[Modules.scala 43:37:@1171.4]
  wire [4:0] _T_55369; // @[Modules.scala 43:37:@1172.4]
  wire [5:0] _T_55370; // @[Modules.scala 43:47:@1173.4]
  wire [4:0] _T_55371; // @[Modules.scala 43:47:@1174.4]
  wire [4:0] _T_55372; // @[Modules.scala 43:47:@1175.4]
  wire [5:0] _T_55373; // @[Modules.scala 37:46:@1177.4]
  wire [4:0] _T_55374; // @[Modules.scala 37:46:@1178.4]
  wire [4:0] _T_55375; // @[Modules.scala 37:46:@1179.4]
  wire [5:0] _T_55376; // @[Modules.scala 40:46:@1181.4]
  wire [4:0] _T_55377; // @[Modules.scala 40:46:@1182.4]
  wire [4:0] _T_55378; // @[Modules.scala 40:46:@1183.4]
  wire [5:0] _T_55380; // @[Modules.scala 43:37:@1185.4]
  wire [4:0] _T_55381; // @[Modules.scala 43:37:@1186.4]
  wire [4:0] _T_55382; // @[Modules.scala 43:37:@1187.4]
  wire [5:0] _T_55383; // @[Modules.scala 43:47:@1188.4]
  wire [4:0] _T_55384; // @[Modules.scala 43:47:@1189.4]
  wire [4:0] _T_55385; // @[Modules.scala 43:47:@1190.4]
  wire [5:0] _T_55387; // @[Modules.scala 46:37:@1192.4]
  wire [4:0] _T_55388; // @[Modules.scala 46:37:@1193.4]
  wire [4:0] _T_55389; // @[Modules.scala 46:37:@1194.4]
  wire [5:0] _T_55390; // @[Modules.scala 46:47:@1195.4]
  wire [4:0] _T_55391; // @[Modules.scala 46:47:@1196.4]
  wire [4:0] _T_55392; // @[Modules.scala 46:47:@1197.4]
  wire [5:0] _T_55394; // @[Modules.scala 46:37:@1199.4]
  wire [4:0] _T_55395; // @[Modules.scala 46:37:@1200.4]
  wire [4:0] _T_55396; // @[Modules.scala 46:37:@1201.4]
  wire [5:0] _T_55397; // @[Modules.scala 46:47:@1202.4]
  wire [4:0] _T_55398; // @[Modules.scala 46:47:@1203.4]
  wire [4:0] _T_55399; // @[Modules.scala 46:47:@1204.4]
  wire [5:0] _T_55400; // @[Modules.scala 37:46:@1206.4]
  wire [4:0] _T_55401; // @[Modules.scala 37:46:@1207.4]
  wire [4:0] _T_55402; // @[Modules.scala 37:46:@1208.4]
  wire [5:0] _T_55403; // @[Modules.scala 37:46:@1210.4]
  wire [4:0] _T_55404; // @[Modules.scala 37:46:@1211.4]
  wire [4:0] _T_55405; // @[Modules.scala 37:46:@1212.4]
  wire [5:0] _T_55406; // @[Modules.scala 37:46:@1214.4]
  wire [4:0] _T_55407; // @[Modules.scala 37:46:@1215.4]
  wire [4:0] _T_55408; // @[Modules.scala 37:46:@1216.4]
  wire [5:0] _T_55409; // @[Modules.scala 37:46:@1218.4]
  wire [4:0] _T_55410; // @[Modules.scala 37:46:@1219.4]
  wire [4:0] _T_55411; // @[Modules.scala 37:46:@1220.4]
  wire [5:0] _T_55412; // @[Modules.scala 37:46:@1222.4]
  wire [4:0] _T_55413; // @[Modules.scala 37:46:@1223.4]
  wire [4:0] _T_55414; // @[Modules.scala 37:46:@1224.4]
  wire [5:0] _T_55415; // @[Modules.scala 37:46:@1226.4]
  wire [4:0] _T_55416; // @[Modules.scala 37:46:@1227.4]
  wire [4:0] _T_55417; // @[Modules.scala 37:46:@1228.4]
  wire [5:0] _T_55418; // @[Modules.scala 37:46:@1230.4]
  wire [4:0] _T_55419; // @[Modules.scala 37:46:@1231.4]
  wire [4:0] _T_55420; // @[Modules.scala 37:46:@1232.4]
  wire [5:0] _T_55421; // @[Modules.scala 37:46:@1234.4]
  wire [4:0] _T_55422; // @[Modules.scala 37:46:@1235.4]
  wire [4:0] _T_55423; // @[Modules.scala 37:46:@1236.4]
  wire [5:0] _T_55424; // @[Modules.scala 37:46:@1238.4]
  wire [4:0] _T_55425; // @[Modules.scala 37:46:@1239.4]
  wire [4:0] _T_55426; // @[Modules.scala 37:46:@1240.4]
  wire [5:0] _T_55427; // @[Modules.scala 37:46:@1242.4]
  wire [4:0] _T_55428; // @[Modules.scala 37:46:@1243.4]
  wire [4:0] _T_55429; // @[Modules.scala 37:46:@1244.4]
  wire [5:0] _T_55430; // @[Modules.scala 40:46:@1246.4]
  wire [4:0] _T_55431; // @[Modules.scala 40:46:@1247.4]
  wire [4:0] _T_55432; // @[Modules.scala 40:46:@1248.4]
  wire [5:0] _T_55434; // @[Modules.scala 43:37:@1250.4]
  wire [4:0] _T_55435; // @[Modules.scala 43:37:@1251.4]
  wire [4:0] _T_55436; // @[Modules.scala 43:37:@1252.4]
  wire [5:0] _T_55437; // @[Modules.scala 43:47:@1253.4]
  wire [4:0] _T_55438; // @[Modules.scala 43:47:@1254.4]
  wire [4:0] _T_55439; // @[Modules.scala 43:47:@1255.4]
  wire [5:0] _T_55441; // @[Modules.scala 43:37:@1257.4]
  wire [4:0] _T_55442; // @[Modules.scala 43:37:@1258.4]
  wire [4:0] _T_55443; // @[Modules.scala 43:37:@1259.4]
  wire [5:0] _T_55444; // @[Modules.scala 43:47:@1260.4]
  wire [4:0] _T_55445; // @[Modules.scala 43:47:@1261.4]
  wire [4:0] _T_55446; // @[Modules.scala 43:47:@1262.4]
  wire [5:0] _T_55448; // @[Modules.scala 46:37:@1264.4]
  wire [4:0] _T_55449; // @[Modules.scala 46:37:@1265.4]
  wire [4:0] _T_55450; // @[Modules.scala 46:37:@1266.4]
  wire [5:0] _T_55451; // @[Modules.scala 46:47:@1267.4]
  wire [4:0] _T_55452; // @[Modules.scala 46:47:@1268.4]
  wire [4:0] _T_55453; // @[Modules.scala 46:47:@1269.4]
  wire [5:0] _T_55455; // @[Modules.scala 43:37:@1271.4]
  wire [4:0] _T_55456; // @[Modules.scala 43:37:@1272.4]
  wire [4:0] _T_55457; // @[Modules.scala 43:37:@1273.4]
  wire [5:0] _T_55458; // @[Modules.scala 43:47:@1274.4]
  wire [4:0] _T_55459; // @[Modules.scala 43:47:@1275.4]
  wire [4:0] _T_55460; // @[Modules.scala 43:47:@1276.4]
  wire [5:0] _T_55461; // @[Modules.scala 37:46:@1278.4]
  wire [4:0] _T_55462; // @[Modules.scala 37:46:@1279.4]
  wire [4:0] _T_55463; // @[Modules.scala 37:46:@1280.4]
  wire [5:0] _T_55464; // @[Modules.scala 37:46:@1282.4]
  wire [4:0] _T_55465; // @[Modules.scala 37:46:@1283.4]
  wire [4:0] _T_55466; // @[Modules.scala 37:46:@1284.4]
  wire [5:0] _T_55467; // @[Modules.scala 37:46:@1286.4]
  wire [4:0] _T_55468; // @[Modules.scala 37:46:@1287.4]
  wire [4:0] _T_55469; // @[Modules.scala 37:46:@1288.4]
  wire [5:0] _T_55470; // @[Modules.scala 37:46:@1290.4]
  wire [4:0] _T_55471; // @[Modules.scala 37:46:@1291.4]
  wire [4:0] _T_55472; // @[Modules.scala 37:46:@1292.4]
  wire [5:0] _T_55473; // @[Modules.scala 37:46:@1294.4]
  wire [4:0] _T_55474; // @[Modules.scala 37:46:@1295.4]
  wire [4:0] _T_55475; // @[Modules.scala 37:46:@1296.4]
  wire [5:0] _T_55476; // @[Modules.scala 37:46:@1298.4]
  wire [4:0] _T_55477; // @[Modules.scala 37:46:@1299.4]
  wire [4:0] _T_55478; // @[Modules.scala 37:46:@1300.4]
  wire [5:0] _T_55479; // @[Modules.scala 40:46:@1302.4]
  wire [4:0] _T_55480; // @[Modules.scala 40:46:@1303.4]
  wire [4:0] _T_55481; // @[Modules.scala 40:46:@1304.4]
  wire [5:0] _T_55482; // @[Modules.scala 40:46:@1306.4]
  wire [4:0] _T_55483; // @[Modules.scala 40:46:@1307.4]
  wire [4:0] _T_55484; // @[Modules.scala 40:46:@1308.4]
  wire [5:0] _T_55486; // @[Modules.scala 43:37:@1310.4]
  wire [4:0] _T_55487; // @[Modules.scala 43:37:@1311.4]
  wire [4:0] _T_55488; // @[Modules.scala 43:37:@1312.4]
  wire [5:0] _T_55489; // @[Modules.scala 43:47:@1313.4]
  wire [4:0] _T_55490; // @[Modules.scala 43:47:@1314.4]
  wire [4:0] _T_55491; // @[Modules.scala 43:47:@1315.4]
  wire [5:0] _T_55493; // @[Modules.scala 46:37:@1317.4]
  wire [4:0] _T_55494; // @[Modules.scala 46:37:@1318.4]
  wire [4:0] _T_55495; // @[Modules.scala 46:37:@1319.4]
  wire [5:0] _T_55496; // @[Modules.scala 46:47:@1320.4]
  wire [4:0] _T_55497; // @[Modules.scala 46:47:@1321.4]
  wire [4:0] _T_55498; // @[Modules.scala 46:47:@1322.4]
  wire [5:0] _T_55500; // @[Modules.scala 46:37:@1324.4]
  wire [4:0] _T_55501; // @[Modules.scala 46:37:@1325.4]
  wire [4:0] _T_55502; // @[Modules.scala 46:37:@1326.4]
  wire [5:0] _T_55503; // @[Modules.scala 46:47:@1327.4]
  wire [4:0] _T_55504; // @[Modules.scala 46:47:@1328.4]
  wire [4:0] _T_55505; // @[Modules.scala 46:47:@1329.4]
  wire [5:0] _T_55506; // @[Modules.scala 37:46:@1331.4]
  wire [4:0] _T_55507; // @[Modules.scala 37:46:@1332.4]
  wire [4:0] _T_55508; // @[Modules.scala 37:46:@1333.4]
  wire [5:0] _T_55510; // @[Modules.scala 46:37:@1335.4]
  wire [4:0] _T_55511; // @[Modules.scala 46:37:@1336.4]
  wire [4:0] _T_55512; // @[Modules.scala 46:37:@1337.4]
  wire [5:0] _T_55513; // @[Modules.scala 46:47:@1338.4]
  wire [4:0] _T_55514; // @[Modules.scala 46:47:@1339.4]
  wire [4:0] _T_55515; // @[Modules.scala 46:47:@1340.4]
  wire [5:0] _T_55517; // @[Modules.scala 43:37:@1342.4]
  wire [4:0] _T_55518; // @[Modules.scala 43:37:@1343.4]
  wire [4:0] _T_55519; // @[Modules.scala 43:37:@1344.4]
  wire [5:0] _T_55520; // @[Modules.scala 43:47:@1345.4]
  wire [4:0] _T_55521; // @[Modules.scala 43:47:@1346.4]
  wire [4:0] _T_55522; // @[Modules.scala 43:47:@1347.4]
  wire [5:0] _T_55523; // @[Modules.scala 37:46:@1349.4]
  wire [4:0] _T_55524; // @[Modules.scala 37:46:@1350.4]
  wire [4:0] _T_55525; // @[Modules.scala 37:46:@1351.4]
  wire [5:0] _T_55526; // @[Modules.scala 37:46:@1353.4]
  wire [4:0] _T_55527; // @[Modules.scala 37:46:@1354.4]
  wire [4:0] _T_55528; // @[Modules.scala 37:46:@1355.4]
  wire [5:0] _T_55529; // @[Modules.scala 37:46:@1357.4]
  wire [4:0] _T_55530; // @[Modules.scala 37:46:@1358.4]
  wire [4:0] _T_55531; // @[Modules.scala 37:46:@1359.4]
  wire [5:0] _T_55532; // @[Modules.scala 40:46:@1361.4]
  wire [4:0] _T_55533; // @[Modules.scala 40:46:@1362.4]
  wire [4:0] _T_55534; // @[Modules.scala 40:46:@1363.4]
  wire [5:0] _T_55535; // @[Modules.scala 37:46:@1365.4]
  wire [4:0] _T_55536; // @[Modules.scala 37:46:@1366.4]
  wire [4:0] _T_55537; // @[Modules.scala 37:46:@1367.4]
  wire [5:0] _T_55538; // @[Modules.scala 37:46:@1369.4]
  wire [4:0] _T_55539; // @[Modules.scala 37:46:@1370.4]
  wire [4:0] _T_55540; // @[Modules.scala 37:46:@1371.4]
  wire [5:0] _T_55541; // @[Modules.scala 37:46:@1373.4]
  wire [4:0] _T_55542; // @[Modules.scala 37:46:@1374.4]
  wire [4:0] _T_55543; // @[Modules.scala 37:46:@1375.4]
  wire [5:0] _T_55544; // @[Modules.scala 40:46:@1377.4]
  wire [4:0] _T_55545; // @[Modules.scala 40:46:@1378.4]
  wire [4:0] _T_55546; // @[Modules.scala 40:46:@1379.4]
  wire [5:0] _T_55548; // @[Modules.scala 46:37:@1381.4]
  wire [4:0] _T_55549; // @[Modules.scala 46:37:@1382.4]
  wire [4:0] _T_55550; // @[Modules.scala 46:37:@1383.4]
  wire [5:0] _T_55551; // @[Modules.scala 46:47:@1384.4]
  wire [4:0] _T_55552; // @[Modules.scala 46:47:@1385.4]
  wire [4:0] _T_55553; // @[Modules.scala 46:47:@1386.4]
  wire [5:0] _T_55555; // @[Modules.scala 46:37:@1388.4]
  wire [4:0] _T_55556; // @[Modules.scala 46:37:@1389.4]
  wire [4:0] _T_55557; // @[Modules.scala 46:37:@1390.4]
  wire [5:0] _T_55558; // @[Modules.scala 46:47:@1391.4]
  wire [4:0] _T_55559; // @[Modules.scala 46:47:@1392.4]
  wire [4:0] _T_55560; // @[Modules.scala 46:47:@1393.4]
  wire [5:0] _T_55562; // @[Modules.scala 46:37:@1395.4]
  wire [4:0] _T_55563; // @[Modules.scala 46:37:@1396.4]
  wire [4:0] _T_55564; // @[Modules.scala 46:37:@1397.4]
  wire [5:0] _T_55565; // @[Modules.scala 46:47:@1398.4]
  wire [4:0] _T_55566; // @[Modules.scala 46:47:@1399.4]
  wire [4:0] _T_55567; // @[Modules.scala 46:47:@1400.4]
  wire [5:0] _T_55569; // @[Modules.scala 46:37:@1402.4]
  wire [4:0] _T_55570; // @[Modules.scala 46:37:@1403.4]
  wire [4:0] _T_55571; // @[Modules.scala 46:37:@1404.4]
  wire [5:0] _T_55572; // @[Modules.scala 46:47:@1405.4]
  wire [4:0] _T_55573; // @[Modules.scala 46:47:@1406.4]
  wire [4:0] _T_55574; // @[Modules.scala 46:47:@1407.4]
  wire [5:0] _T_55575; // @[Modules.scala 40:46:@1409.4]
  wire [4:0] _T_55576; // @[Modules.scala 40:46:@1410.4]
  wire [4:0] _T_55577; // @[Modules.scala 40:46:@1411.4]
  wire [5:0] _T_55579; // @[Modules.scala 46:37:@1413.4]
  wire [4:0] _T_55580; // @[Modules.scala 46:37:@1414.4]
  wire [4:0] _T_55581; // @[Modules.scala 46:37:@1415.4]
  wire [5:0] _T_55582; // @[Modules.scala 46:47:@1416.4]
  wire [4:0] _T_55583; // @[Modules.scala 46:47:@1417.4]
  wire [4:0] _T_55584; // @[Modules.scala 46:47:@1418.4]
  wire [5:0] _T_55585; // @[Modules.scala 37:46:@1420.4]
  wire [4:0] _T_55586; // @[Modules.scala 37:46:@1421.4]
  wire [4:0] _T_55587; // @[Modules.scala 37:46:@1422.4]
  wire [5:0] _T_55588; // @[Modules.scala 37:46:@1424.4]
  wire [4:0] _T_55589; // @[Modules.scala 37:46:@1425.4]
  wire [4:0] _T_55590; // @[Modules.scala 37:46:@1426.4]
  wire [5:0] _T_55591; // @[Modules.scala 37:46:@1428.4]
  wire [4:0] _T_55592; // @[Modules.scala 37:46:@1429.4]
  wire [4:0] _T_55593; // @[Modules.scala 37:46:@1430.4]
  wire [5:0] _T_55595; // @[Modules.scala 43:37:@1432.4]
  wire [4:0] _T_55596; // @[Modules.scala 43:37:@1433.4]
  wire [4:0] _T_55597; // @[Modules.scala 43:37:@1434.4]
  wire [5:0] _T_55598; // @[Modules.scala 43:47:@1435.4]
  wire [4:0] _T_55599; // @[Modules.scala 43:47:@1436.4]
  wire [4:0] _T_55600; // @[Modules.scala 43:47:@1437.4]
  wire [5:0] _T_55601; // @[Modules.scala 37:46:@1439.4]
  wire [4:0] _T_55602; // @[Modules.scala 37:46:@1440.4]
  wire [4:0] _T_55603; // @[Modules.scala 37:46:@1441.4]
  wire [5:0] _T_55604; // @[Modules.scala 40:46:@1443.4]
  wire [4:0] _T_55605; // @[Modules.scala 40:46:@1444.4]
  wire [4:0] _T_55606; // @[Modules.scala 40:46:@1445.4]
  wire [5:0] _T_55607; // @[Modules.scala 40:46:@1447.4]
  wire [4:0] _T_55608; // @[Modules.scala 40:46:@1448.4]
  wire [4:0] _T_55609; // @[Modules.scala 40:46:@1449.4]
  wire [5:0] _T_55611; // @[Modules.scala 46:37:@1451.4]
  wire [4:0] _T_55612; // @[Modules.scala 46:37:@1452.4]
  wire [4:0] _T_55613; // @[Modules.scala 46:37:@1453.4]
  wire [5:0] _T_55614; // @[Modules.scala 46:47:@1454.4]
  wire [4:0] _T_55615; // @[Modules.scala 46:47:@1455.4]
  wire [4:0] _T_55616; // @[Modules.scala 46:47:@1456.4]
  wire [5:0] _T_55617; // @[Modules.scala 37:46:@1458.4]
  wire [4:0] _T_55618; // @[Modules.scala 37:46:@1459.4]
  wire [4:0] _T_55619; // @[Modules.scala 37:46:@1460.4]
  wire [5:0] _T_55621; // @[Modules.scala 46:37:@1462.4]
  wire [4:0] _T_55622; // @[Modules.scala 46:37:@1463.4]
  wire [4:0] _T_55623; // @[Modules.scala 46:37:@1464.4]
  wire [5:0] _T_55624; // @[Modules.scala 46:47:@1465.4]
  wire [4:0] _T_55625; // @[Modules.scala 46:47:@1466.4]
  wire [4:0] _T_55626; // @[Modules.scala 46:47:@1467.4]
  wire [5:0] _T_55628; // @[Modules.scala 46:37:@1469.4]
  wire [4:0] _T_55629; // @[Modules.scala 46:37:@1470.4]
  wire [4:0] _T_55630; // @[Modules.scala 46:37:@1471.4]
  wire [5:0] _T_55631; // @[Modules.scala 46:47:@1472.4]
  wire [4:0] _T_55632; // @[Modules.scala 46:47:@1473.4]
  wire [4:0] _T_55633; // @[Modules.scala 46:47:@1474.4]
  wire [5:0] _T_55635; // @[Modules.scala 46:37:@1476.4]
  wire [4:0] _T_55636; // @[Modules.scala 46:37:@1477.4]
  wire [4:0] _T_55637; // @[Modules.scala 46:37:@1478.4]
  wire [5:0] _T_55638; // @[Modules.scala 46:47:@1479.4]
  wire [4:0] _T_55639; // @[Modules.scala 46:47:@1480.4]
  wire [4:0] _T_55640; // @[Modules.scala 46:47:@1481.4]
  wire [5:0] _T_55642; // @[Modules.scala 43:37:@1483.4]
  wire [4:0] _T_55643; // @[Modules.scala 43:37:@1484.4]
  wire [4:0] _T_55644; // @[Modules.scala 43:37:@1485.4]
  wire [5:0] _T_55645; // @[Modules.scala 43:47:@1486.4]
  wire [4:0] _T_55646; // @[Modules.scala 43:47:@1487.4]
  wire [4:0] _T_55647; // @[Modules.scala 43:47:@1488.4]
  wire [5:0] _T_55649; // @[Modules.scala 46:37:@1490.4]
  wire [4:0] _T_55650; // @[Modules.scala 46:37:@1491.4]
  wire [4:0] _T_55651; // @[Modules.scala 46:37:@1492.4]
  wire [5:0] _T_55652; // @[Modules.scala 46:47:@1493.4]
  wire [4:0] _T_55653; // @[Modules.scala 46:47:@1494.4]
  wire [4:0] _T_55654; // @[Modules.scala 46:47:@1495.4]
  wire [5:0] _T_55656; // @[Modules.scala 46:37:@1497.4]
  wire [4:0] _T_55657; // @[Modules.scala 46:37:@1498.4]
  wire [4:0] _T_55658; // @[Modules.scala 46:37:@1499.4]
  wire [5:0] _T_55659; // @[Modules.scala 46:47:@1500.4]
  wire [4:0] _T_55660; // @[Modules.scala 46:47:@1501.4]
  wire [4:0] _T_55661; // @[Modules.scala 46:47:@1502.4]
  wire [5:0] _T_55662; // @[Modules.scala 37:46:@1504.4]
  wire [4:0] _T_55663; // @[Modules.scala 37:46:@1505.4]
  wire [4:0] _T_55664; // @[Modules.scala 37:46:@1506.4]
  wire [5:0] _T_55665; // @[Modules.scala 37:46:@1508.4]
  wire [4:0] _T_55666; // @[Modules.scala 37:46:@1509.4]
  wire [4:0] _T_55667; // @[Modules.scala 37:46:@1510.4]
  wire [5:0] _T_55668; // @[Modules.scala 40:46:@1512.4]
  wire [4:0] _T_55669; // @[Modules.scala 40:46:@1513.4]
  wire [4:0] _T_55670; // @[Modules.scala 40:46:@1514.4]
  wire [5:0] _T_55671; // @[Modules.scala 37:46:@1516.4]
  wire [4:0] _T_55672; // @[Modules.scala 37:46:@1517.4]
  wire [4:0] _T_55673; // @[Modules.scala 37:46:@1518.4]
  wire [5:0] _T_55675; // @[Modules.scala 43:37:@1520.4]
  wire [4:0] _T_55676; // @[Modules.scala 43:37:@1521.4]
  wire [4:0] _T_55677; // @[Modules.scala 43:37:@1522.4]
  wire [5:0] _T_55678; // @[Modules.scala 43:47:@1523.4]
  wire [4:0] _T_55679; // @[Modules.scala 43:47:@1524.4]
  wire [4:0] _T_55680; // @[Modules.scala 43:47:@1525.4]
  wire [5:0] _T_55682; // @[Modules.scala 43:37:@1527.4]
  wire [4:0] _T_55683; // @[Modules.scala 43:37:@1528.4]
  wire [4:0] _T_55684; // @[Modules.scala 43:37:@1529.4]
  wire [5:0] _T_55685; // @[Modules.scala 43:47:@1530.4]
  wire [4:0] _T_55686; // @[Modules.scala 43:47:@1531.4]
  wire [4:0] _T_55687; // @[Modules.scala 43:47:@1532.4]
  wire [5:0] _T_55689; // @[Modules.scala 43:37:@1534.4]
  wire [4:0] _T_55690; // @[Modules.scala 43:37:@1535.4]
  wire [4:0] _T_55691; // @[Modules.scala 43:37:@1536.4]
  wire [5:0] _T_55692; // @[Modules.scala 43:47:@1537.4]
  wire [4:0] _T_55693; // @[Modules.scala 43:47:@1538.4]
  wire [4:0] _T_55694; // @[Modules.scala 43:47:@1539.4]
  wire [5:0] _T_55695; // @[Modules.scala 37:46:@1541.4]
  wire [4:0] _T_55696; // @[Modules.scala 37:46:@1542.4]
  wire [4:0] _T_55697; // @[Modules.scala 37:46:@1543.4]
  wire [5:0] _T_55698; // @[Modules.scala 37:46:@1545.4]
  wire [4:0] _T_55699; // @[Modules.scala 37:46:@1546.4]
  wire [4:0] _T_55700; // @[Modules.scala 37:46:@1547.4]
  wire [5:0] _T_55702; // @[Modules.scala 46:37:@1549.4]
  wire [4:0] _T_55703; // @[Modules.scala 46:37:@1550.4]
  wire [4:0] _T_55704; // @[Modules.scala 46:37:@1551.4]
  wire [5:0] _T_55705; // @[Modules.scala 46:47:@1552.4]
  wire [4:0] _T_55706; // @[Modules.scala 46:47:@1553.4]
  wire [4:0] _T_55707; // @[Modules.scala 46:47:@1554.4]
  wire [5:0] _T_55708; // @[Modules.scala 40:46:@1556.4]
  wire [4:0] _T_55709; // @[Modules.scala 40:46:@1557.4]
  wire [4:0] _T_55710; // @[Modules.scala 40:46:@1558.4]
  wire [5:0] _T_55712; // @[Modules.scala 43:37:@1560.4]
  wire [4:0] _T_55713; // @[Modules.scala 43:37:@1561.4]
  wire [4:0] _T_55714; // @[Modules.scala 43:37:@1562.4]
  wire [5:0] _T_55715; // @[Modules.scala 43:47:@1563.4]
  wire [4:0] _T_55716; // @[Modules.scala 43:47:@1564.4]
  wire [4:0] _T_55717; // @[Modules.scala 43:47:@1565.4]
  wire [5:0] _T_55719; // @[Modules.scala 46:37:@1567.4]
  wire [4:0] _T_55720; // @[Modules.scala 46:37:@1568.4]
  wire [4:0] _T_55721; // @[Modules.scala 46:37:@1569.4]
  wire [5:0] _T_55722; // @[Modules.scala 46:47:@1570.4]
  wire [4:0] _T_55723; // @[Modules.scala 46:47:@1571.4]
  wire [4:0] _T_55724; // @[Modules.scala 46:47:@1572.4]
  wire [5:0] _T_55726; // @[Modules.scala 46:37:@1574.4]
  wire [4:0] _T_55727; // @[Modules.scala 46:37:@1575.4]
  wire [4:0] _T_55728; // @[Modules.scala 46:37:@1576.4]
  wire [5:0] _T_55729; // @[Modules.scala 46:47:@1577.4]
  wire [4:0] _T_55730; // @[Modules.scala 46:47:@1578.4]
  wire [4:0] _T_55731; // @[Modules.scala 46:47:@1579.4]
  wire [5:0] _T_55733; // @[Modules.scala 46:37:@1581.4]
  wire [4:0] _T_55734; // @[Modules.scala 46:37:@1582.4]
  wire [4:0] _T_55735; // @[Modules.scala 46:37:@1583.4]
  wire [5:0] _T_55736; // @[Modules.scala 46:47:@1584.4]
  wire [4:0] _T_55737; // @[Modules.scala 46:47:@1585.4]
  wire [4:0] _T_55738; // @[Modules.scala 46:47:@1586.4]
  wire [5:0] _T_55740; // @[Modules.scala 43:37:@1588.4]
  wire [4:0] _T_55741; // @[Modules.scala 43:37:@1589.4]
  wire [4:0] _T_55742; // @[Modules.scala 43:37:@1590.4]
  wire [5:0] _T_55743; // @[Modules.scala 43:47:@1591.4]
  wire [4:0] _T_55744; // @[Modules.scala 43:47:@1592.4]
  wire [4:0] _T_55745; // @[Modules.scala 43:47:@1593.4]
  wire [5:0] _T_55747; // @[Modules.scala 46:37:@1595.4]
  wire [4:0] _T_55748; // @[Modules.scala 46:37:@1596.4]
  wire [4:0] _T_55749; // @[Modules.scala 46:37:@1597.4]
  wire [5:0] _T_55750; // @[Modules.scala 46:47:@1598.4]
  wire [4:0] _T_55751; // @[Modules.scala 46:47:@1599.4]
  wire [4:0] _T_55752; // @[Modules.scala 46:47:@1600.4]
  wire [5:0] _T_55754; // @[Modules.scala 46:37:@1602.4]
  wire [4:0] _T_55755; // @[Modules.scala 46:37:@1603.4]
  wire [4:0] _T_55756; // @[Modules.scala 46:37:@1604.4]
  wire [5:0] _T_55757; // @[Modules.scala 46:47:@1605.4]
  wire [4:0] _T_55758; // @[Modules.scala 46:47:@1606.4]
  wire [4:0] _T_55759; // @[Modules.scala 46:47:@1607.4]
  wire [5:0] _T_55761; // @[Modules.scala 46:37:@1609.4]
  wire [4:0] _T_55762; // @[Modules.scala 46:37:@1610.4]
  wire [4:0] _T_55763; // @[Modules.scala 46:37:@1611.4]
  wire [5:0] _T_55764; // @[Modules.scala 46:47:@1612.4]
  wire [4:0] _T_55765; // @[Modules.scala 46:47:@1613.4]
  wire [4:0] _T_55766; // @[Modules.scala 46:47:@1614.4]
  wire [5:0] _T_55767; // @[Modules.scala 40:46:@1616.4]
  wire [4:0] _T_55768; // @[Modules.scala 40:46:@1617.4]
  wire [4:0] _T_55769; // @[Modules.scala 40:46:@1618.4]
  wire [5:0] _T_55770; // @[Modules.scala 40:46:@1620.4]
  wire [4:0] _T_55771; // @[Modules.scala 40:46:@1621.4]
  wire [4:0] _T_55772; // @[Modules.scala 40:46:@1622.4]
  wire [5:0] _T_55774; // @[Modules.scala 46:37:@1624.4]
  wire [4:0] _T_55775; // @[Modules.scala 46:37:@1625.4]
  wire [4:0] _T_55776; // @[Modules.scala 46:37:@1626.4]
  wire [5:0] _T_55777; // @[Modules.scala 46:47:@1627.4]
  wire [4:0] _T_55778; // @[Modules.scala 46:47:@1628.4]
  wire [4:0] _T_55779; // @[Modules.scala 46:47:@1629.4]
  wire [5:0] _T_55780; // @[Modules.scala 40:46:@1631.4]
  wire [4:0] _T_55781; // @[Modules.scala 40:46:@1632.4]
  wire [4:0] _T_55782; // @[Modules.scala 40:46:@1633.4]
  wire [5:0] _T_55784; // @[Modules.scala 43:37:@1635.4]
  wire [4:0] _T_55785; // @[Modules.scala 43:37:@1636.4]
  wire [4:0] _T_55786; // @[Modules.scala 43:37:@1637.4]
  wire [5:0] _T_55787; // @[Modules.scala 43:47:@1638.4]
  wire [4:0] _T_55788; // @[Modules.scala 43:47:@1639.4]
  wire [4:0] _T_55789; // @[Modules.scala 43:47:@1640.4]
  wire [5:0] _T_55791; // @[Modules.scala 46:37:@1642.4]
  wire [4:0] _T_55792; // @[Modules.scala 46:37:@1643.4]
  wire [4:0] _T_55793; // @[Modules.scala 46:37:@1644.4]
  wire [5:0] _T_55794; // @[Modules.scala 46:47:@1645.4]
  wire [4:0] _T_55795; // @[Modules.scala 46:47:@1646.4]
  wire [4:0] _T_55796; // @[Modules.scala 46:47:@1647.4]
  wire [5:0] _T_55798; // @[Modules.scala 46:37:@1649.4]
  wire [4:0] _T_55799; // @[Modules.scala 46:37:@1650.4]
  wire [4:0] _T_55800; // @[Modules.scala 46:37:@1651.4]
  wire [5:0] _T_55801; // @[Modules.scala 46:47:@1652.4]
  wire [4:0] _T_55802; // @[Modules.scala 46:47:@1653.4]
  wire [4:0] _T_55803; // @[Modules.scala 46:47:@1654.4]
  wire [5:0] _T_55805; // @[Modules.scala 46:37:@1656.4]
  wire [4:0] _T_55806; // @[Modules.scala 46:37:@1657.4]
  wire [4:0] _T_55807; // @[Modules.scala 46:37:@1658.4]
  wire [5:0] _T_55808; // @[Modules.scala 46:47:@1659.4]
  wire [4:0] _T_55809; // @[Modules.scala 46:47:@1660.4]
  wire [4:0] _T_55810; // @[Modules.scala 46:47:@1661.4]
  wire [5:0] _T_55812; // @[Modules.scala 46:37:@1663.4]
  wire [4:0] _T_55813; // @[Modules.scala 46:37:@1664.4]
  wire [4:0] _T_55814; // @[Modules.scala 46:37:@1665.4]
  wire [5:0] _T_55815; // @[Modules.scala 46:47:@1666.4]
  wire [4:0] _T_55816; // @[Modules.scala 46:47:@1667.4]
  wire [4:0] _T_55817; // @[Modules.scala 46:47:@1668.4]
  wire [5:0] _T_55819; // @[Modules.scala 46:37:@1670.4]
  wire [4:0] _T_55820; // @[Modules.scala 46:37:@1671.4]
  wire [4:0] _T_55821; // @[Modules.scala 46:37:@1672.4]
  wire [5:0] _T_55822; // @[Modules.scala 46:47:@1673.4]
  wire [4:0] _T_55823; // @[Modules.scala 46:47:@1674.4]
  wire [4:0] _T_55824; // @[Modules.scala 46:47:@1675.4]
  wire [5:0] _T_55826; // @[Modules.scala 43:37:@1677.4]
  wire [4:0] _T_55827; // @[Modules.scala 43:37:@1678.4]
  wire [4:0] _T_55828; // @[Modules.scala 43:37:@1679.4]
  wire [5:0] _T_55829; // @[Modules.scala 43:47:@1680.4]
  wire [4:0] _T_55830; // @[Modules.scala 43:47:@1681.4]
  wire [4:0] _T_55831; // @[Modules.scala 43:47:@1682.4]
  wire [5:0] _T_55833; // @[Modules.scala 43:37:@1684.4]
  wire [4:0] _T_55834; // @[Modules.scala 43:37:@1685.4]
  wire [4:0] _T_55835; // @[Modules.scala 43:37:@1686.4]
  wire [5:0] _T_55836; // @[Modules.scala 43:47:@1687.4]
  wire [4:0] _T_55837; // @[Modules.scala 43:47:@1688.4]
  wire [4:0] _T_55838; // @[Modules.scala 43:47:@1689.4]
  wire [5:0] _T_55840; // @[Modules.scala 43:37:@1691.4]
  wire [4:0] _T_55841; // @[Modules.scala 43:37:@1692.4]
  wire [4:0] _T_55842; // @[Modules.scala 43:37:@1693.4]
  wire [5:0] _T_55843; // @[Modules.scala 43:47:@1694.4]
  wire [4:0] _T_55844; // @[Modules.scala 43:47:@1695.4]
  wire [4:0] _T_55845; // @[Modules.scala 43:47:@1696.4]
  wire [5:0] _T_55846; // @[Modules.scala 37:46:@1698.4]
  wire [4:0] _T_55847; // @[Modules.scala 37:46:@1699.4]
  wire [4:0] _T_55848; // @[Modules.scala 37:46:@1700.4]
  wire [5:0] _T_55849; // @[Modules.scala 40:46:@1702.4]
  wire [4:0] _T_55850; // @[Modules.scala 40:46:@1703.4]
  wire [4:0] _T_55851; // @[Modules.scala 40:46:@1704.4]
  wire [5:0] _T_55852; // @[Modules.scala 40:46:@1706.4]
  wire [4:0] _T_55853; // @[Modules.scala 40:46:@1707.4]
  wire [4:0] _T_55854; // @[Modules.scala 40:46:@1708.4]
  wire [5:0] _T_55856; // @[Modules.scala 46:37:@1710.4]
  wire [4:0] _T_55857; // @[Modules.scala 46:37:@1711.4]
  wire [4:0] _T_55858; // @[Modules.scala 46:37:@1712.4]
  wire [5:0] _T_55859; // @[Modules.scala 46:47:@1713.4]
  wire [4:0] _T_55860; // @[Modules.scala 46:47:@1714.4]
  wire [4:0] _T_55861; // @[Modules.scala 46:47:@1715.4]
  wire [5:0] _T_55862; // @[Modules.scala 37:46:@1717.4]
  wire [4:0] _T_55863; // @[Modules.scala 37:46:@1718.4]
  wire [4:0] _T_55864; // @[Modules.scala 37:46:@1719.4]
  wire [5:0] _T_55866; // @[Modules.scala 43:37:@1721.4]
  wire [4:0] _T_55867; // @[Modules.scala 43:37:@1722.4]
  wire [4:0] _T_55868; // @[Modules.scala 43:37:@1723.4]
  wire [5:0] _T_55869; // @[Modules.scala 43:47:@1724.4]
  wire [4:0] _T_55870; // @[Modules.scala 43:47:@1725.4]
  wire [4:0] _T_55871; // @[Modules.scala 43:47:@1726.4]
  wire [5:0] _T_55873; // @[Modules.scala 43:37:@1728.4]
  wire [4:0] _T_55874; // @[Modules.scala 43:37:@1729.4]
  wire [4:0] _T_55875; // @[Modules.scala 43:37:@1730.4]
  wire [5:0] _T_55876; // @[Modules.scala 43:47:@1731.4]
  wire [4:0] _T_55877; // @[Modules.scala 43:47:@1732.4]
  wire [4:0] _T_55878; // @[Modules.scala 43:47:@1733.4]
  wire [5:0] _T_55880; // @[Modules.scala 46:37:@1735.4]
  wire [4:0] _T_55881; // @[Modules.scala 46:37:@1736.4]
  wire [4:0] _T_55882; // @[Modules.scala 46:37:@1737.4]
  wire [5:0] _T_55883; // @[Modules.scala 46:47:@1738.4]
  wire [4:0] _T_55884; // @[Modules.scala 46:47:@1739.4]
  wire [4:0] _T_55885; // @[Modules.scala 46:47:@1740.4]
  wire [5:0] _T_55887; // @[Modules.scala 46:37:@1742.4]
  wire [4:0] _T_55888; // @[Modules.scala 46:37:@1743.4]
  wire [4:0] _T_55889; // @[Modules.scala 46:37:@1744.4]
  wire [5:0] _T_55890; // @[Modules.scala 46:47:@1745.4]
  wire [4:0] _T_55891; // @[Modules.scala 46:47:@1746.4]
  wire [4:0] _T_55892; // @[Modules.scala 46:47:@1747.4]
  wire [5:0] _T_55894; // @[Modules.scala 46:37:@1749.4]
  wire [4:0] _T_55895; // @[Modules.scala 46:37:@1750.4]
  wire [4:0] _T_55896; // @[Modules.scala 46:37:@1751.4]
  wire [5:0] _T_55897; // @[Modules.scala 46:47:@1752.4]
  wire [4:0] _T_55898; // @[Modules.scala 46:47:@1753.4]
  wire [4:0] _T_55899; // @[Modules.scala 46:47:@1754.4]
  wire [5:0] _T_55901; // @[Modules.scala 46:37:@1756.4]
  wire [4:0] _T_55902; // @[Modules.scala 46:37:@1757.4]
  wire [4:0] _T_55903; // @[Modules.scala 46:37:@1758.4]
  wire [5:0] _T_55904; // @[Modules.scala 46:47:@1759.4]
  wire [4:0] _T_55905; // @[Modules.scala 46:47:@1760.4]
  wire [4:0] _T_55906; // @[Modules.scala 46:47:@1761.4]
  wire [5:0] _T_55908; // @[Modules.scala 46:37:@1763.4]
  wire [4:0] _T_55909; // @[Modules.scala 46:37:@1764.4]
  wire [4:0] _T_55910; // @[Modules.scala 46:37:@1765.4]
  wire [5:0] _T_55911; // @[Modules.scala 46:47:@1766.4]
  wire [4:0] _T_55912; // @[Modules.scala 46:47:@1767.4]
  wire [4:0] _T_55913; // @[Modules.scala 46:47:@1768.4]
  wire [5:0] _T_55914; // @[Modules.scala 37:46:@1770.4]
  wire [4:0] _T_55915; // @[Modules.scala 37:46:@1771.4]
  wire [4:0] _T_55916; // @[Modules.scala 37:46:@1772.4]
  wire [5:0] _T_55917; // @[Modules.scala 40:46:@1774.4]
  wire [4:0] _T_55918; // @[Modules.scala 40:46:@1775.4]
  wire [4:0] _T_55919; // @[Modules.scala 40:46:@1776.4]
  wire [5:0] _T_55920; // @[Modules.scala 37:46:@1778.4]
  wire [4:0] _T_55921; // @[Modules.scala 37:46:@1779.4]
  wire [4:0] _T_55922; // @[Modules.scala 37:46:@1780.4]
  wire [5:0] _T_55923; // @[Modules.scala 37:46:@1782.4]
  wire [4:0] _T_55924; // @[Modules.scala 37:46:@1783.4]
  wire [4:0] _T_55925; // @[Modules.scala 37:46:@1784.4]
  wire [5:0] _T_55927; // @[Modules.scala 46:37:@1786.4]
  wire [4:0] _T_55928; // @[Modules.scala 46:37:@1787.4]
  wire [4:0] _T_55929; // @[Modules.scala 46:37:@1788.4]
  wire [5:0] _T_55930; // @[Modules.scala 46:47:@1789.4]
  wire [4:0] _T_55931; // @[Modules.scala 46:47:@1790.4]
  wire [4:0] _T_55932; // @[Modules.scala 46:47:@1791.4]
  wire [5:0] _T_55934; // @[Modules.scala 46:37:@1793.4]
  wire [4:0] _T_55935; // @[Modules.scala 46:37:@1794.4]
  wire [4:0] _T_55936; // @[Modules.scala 46:37:@1795.4]
  wire [5:0] _T_55937; // @[Modules.scala 46:47:@1796.4]
  wire [4:0] _T_55938; // @[Modules.scala 46:47:@1797.4]
  wire [4:0] _T_55939; // @[Modules.scala 46:47:@1798.4]
  wire [5:0] _T_55940; // @[Modules.scala 37:46:@1800.4]
  wire [4:0] _T_55941; // @[Modules.scala 37:46:@1801.4]
  wire [4:0] _T_55942; // @[Modules.scala 37:46:@1802.4]
  wire [5:0] _T_55944; // @[Modules.scala 43:37:@1804.4]
  wire [4:0] _T_55945; // @[Modules.scala 43:37:@1805.4]
  wire [4:0] _T_55946; // @[Modules.scala 43:37:@1806.4]
  wire [5:0] _T_55947; // @[Modules.scala 43:47:@1807.4]
  wire [4:0] _T_55948; // @[Modules.scala 43:47:@1808.4]
  wire [4:0] _T_55949; // @[Modules.scala 43:47:@1809.4]
  wire [5:0] _T_55951; // @[Modules.scala 43:37:@1811.4]
  wire [4:0] _T_55952; // @[Modules.scala 43:37:@1812.4]
  wire [4:0] _T_55953; // @[Modules.scala 43:37:@1813.4]
  wire [5:0] _T_55954; // @[Modules.scala 43:47:@1814.4]
  wire [4:0] _T_55955; // @[Modules.scala 43:47:@1815.4]
  wire [4:0] _T_55956; // @[Modules.scala 43:47:@1816.4]
  wire [5:0] _T_55957; // @[Modules.scala 37:46:@1818.4]
  wire [4:0] _T_55958; // @[Modules.scala 37:46:@1819.4]
  wire [4:0] _T_55959; // @[Modules.scala 37:46:@1820.4]
  wire [5:0] _T_55961; // @[Modules.scala 46:37:@1822.4]
  wire [4:0] _T_55962; // @[Modules.scala 46:37:@1823.4]
  wire [4:0] _T_55963; // @[Modules.scala 46:37:@1824.4]
  wire [5:0] _T_55964; // @[Modules.scala 46:47:@1825.4]
  wire [4:0] _T_55965; // @[Modules.scala 46:47:@1826.4]
  wire [4:0] _T_55966; // @[Modules.scala 46:47:@1827.4]
  wire [5:0] _T_55968; // @[Modules.scala 46:37:@1829.4]
  wire [4:0] _T_55969; // @[Modules.scala 46:37:@1830.4]
  wire [4:0] _T_55970; // @[Modules.scala 46:37:@1831.4]
  wire [5:0] _T_55971; // @[Modules.scala 46:47:@1832.4]
  wire [4:0] _T_55972; // @[Modules.scala 46:47:@1833.4]
  wire [4:0] _T_55973; // @[Modules.scala 46:47:@1834.4]
  wire [5:0] _T_55975; // @[Modules.scala 46:37:@1836.4]
  wire [4:0] _T_55976; // @[Modules.scala 46:37:@1837.4]
  wire [4:0] _T_55977; // @[Modules.scala 46:37:@1838.4]
  wire [5:0] _T_55978; // @[Modules.scala 46:47:@1839.4]
  wire [4:0] _T_55979; // @[Modules.scala 46:47:@1840.4]
  wire [4:0] _T_55980; // @[Modules.scala 46:47:@1841.4]
  wire [5:0] _T_55982; // @[Modules.scala 46:37:@1843.4]
  wire [4:0] _T_55983; // @[Modules.scala 46:37:@1844.4]
  wire [4:0] _T_55984; // @[Modules.scala 46:37:@1845.4]
  wire [5:0] _T_55985; // @[Modules.scala 46:47:@1846.4]
  wire [4:0] _T_55986; // @[Modules.scala 46:47:@1847.4]
  wire [4:0] _T_55987; // @[Modules.scala 46:47:@1848.4]
  wire [5:0] _T_55989; // @[Modules.scala 46:37:@1850.4]
  wire [4:0] _T_55990; // @[Modules.scala 46:37:@1851.4]
  wire [4:0] _T_55991; // @[Modules.scala 46:37:@1852.4]
  wire [5:0] _T_55992; // @[Modules.scala 46:47:@1853.4]
  wire [4:0] _T_55993; // @[Modules.scala 46:47:@1854.4]
  wire [4:0] _T_55994; // @[Modules.scala 46:47:@1855.4]
  wire [5:0] _T_55996; // @[Modules.scala 46:37:@1857.4]
  wire [4:0] _T_55997; // @[Modules.scala 46:37:@1858.4]
  wire [4:0] _T_55998; // @[Modules.scala 46:37:@1859.4]
  wire [5:0] _T_55999; // @[Modules.scala 46:47:@1860.4]
  wire [4:0] _T_56000; // @[Modules.scala 46:47:@1861.4]
  wire [4:0] _T_56001; // @[Modules.scala 46:47:@1862.4]
  wire [5:0] _T_56003; // @[Modules.scala 46:37:@1864.4]
  wire [4:0] _T_56004; // @[Modules.scala 46:37:@1865.4]
  wire [4:0] _T_56005; // @[Modules.scala 46:37:@1866.4]
  wire [5:0] _T_56006; // @[Modules.scala 46:47:@1867.4]
  wire [4:0] _T_56007; // @[Modules.scala 46:47:@1868.4]
  wire [4:0] _T_56008; // @[Modules.scala 46:47:@1869.4]
  wire [5:0] _T_56010; // @[Modules.scala 46:37:@1871.4]
  wire [4:0] _T_56011; // @[Modules.scala 46:37:@1872.4]
  wire [4:0] _T_56012; // @[Modules.scala 46:37:@1873.4]
  wire [5:0] _T_56013; // @[Modules.scala 46:47:@1874.4]
  wire [4:0] _T_56014; // @[Modules.scala 46:47:@1875.4]
  wire [4:0] _T_56015; // @[Modules.scala 46:47:@1876.4]
  wire [5:0] _T_56017; // @[Modules.scala 46:37:@1878.4]
  wire [4:0] _T_56018; // @[Modules.scala 46:37:@1879.4]
  wire [4:0] _T_56019; // @[Modules.scala 46:37:@1880.4]
  wire [5:0] _T_56020; // @[Modules.scala 46:47:@1881.4]
  wire [4:0] _T_56021; // @[Modules.scala 46:47:@1882.4]
  wire [4:0] _T_56022; // @[Modules.scala 46:47:@1883.4]
  wire [5:0] _T_56024; // @[Modules.scala 43:37:@1885.4]
  wire [4:0] _T_56025; // @[Modules.scala 43:37:@1886.4]
  wire [4:0] _T_56026; // @[Modules.scala 43:37:@1887.4]
  wire [5:0] _T_56027; // @[Modules.scala 43:47:@1888.4]
  wire [4:0] _T_56028; // @[Modules.scala 43:47:@1889.4]
  wire [4:0] _T_56029; // @[Modules.scala 43:47:@1890.4]
  wire [5:0] _T_56030; // @[Modules.scala 37:46:@1892.4]
  wire [4:0] _T_56031; // @[Modules.scala 37:46:@1893.4]
  wire [4:0] _T_56032; // @[Modules.scala 37:46:@1894.4]
  wire [5:0] _T_56034; // @[Modules.scala 43:37:@1896.4]
  wire [4:0] _T_56035; // @[Modules.scala 43:37:@1897.4]
  wire [4:0] _T_56036; // @[Modules.scala 43:37:@1898.4]
  wire [5:0] _T_56037; // @[Modules.scala 43:47:@1899.4]
  wire [4:0] _T_56038; // @[Modules.scala 43:47:@1900.4]
  wire [4:0] _T_56039; // @[Modules.scala 43:47:@1901.4]
  wire [5:0] _T_56041; // @[Modules.scala 43:37:@1903.4]
  wire [4:0] _T_56042; // @[Modules.scala 43:37:@1904.4]
  wire [4:0] _T_56043; // @[Modules.scala 43:37:@1905.4]
  wire [5:0] _T_56044; // @[Modules.scala 43:47:@1906.4]
  wire [4:0] _T_56045; // @[Modules.scala 43:47:@1907.4]
  wire [4:0] _T_56046; // @[Modules.scala 43:47:@1908.4]
  wire [5:0] _T_56047; // @[Modules.scala 37:46:@1910.4]
  wire [4:0] _T_56048; // @[Modules.scala 37:46:@1911.4]
  wire [4:0] _T_56049; // @[Modules.scala 37:46:@1912.4]
  wire [5:0] _T_56051; // @[Modules.scala 46:37:@1914.4]
  wire [4:0] _T_56052; // @[Modules.scala 46:37:@1915.4]
  wire [4:0] _T_56053; // @[Modules.scala 46:37:@1916.4]
  wire [5:0] _T_56054; // @[Modules.scala 46:47:@1917.4]
  wire [4:0] _T_56055; // @[Modules.scala 46:47:@1918.4]
  wire [4:0] _T_56056; // @[Modules.scala 46:47:@1919.4]
  wire [5:0] _T_56058; // @[Modules.scala 46:37:@1921.4]
  wire [4:0] _T_56059; // @[Modules.scala 46:37:@1922.4]
  wire [4:0] _T_56060; // @[Modules.scala 46:37:@1923.4]
  wire [5:0] _T_56061; // @[Modules.scala 46:47:@1924.4]
  wire [4:0] _T_56062; // @[Modules.scala 46:47:@1925.4]
  wire [4:0] _T_56063; // @[Modules.scala 46:47:@1926.4]
  wire [5:0] _T_56065; // @[Modules.scala 46:37:@1928.4]
  wire [4:0] _T_56066; // @[Modules.scala 46:37:@1929.4]
  wire [4:0] _T_56067; // @[Modules.scala 46:37:@1930.4]
  wire [5:0] _T_56068; // @[Modules.scala 46:47:@1931.4]
  wire [4:0] _T_56069; // @[Modules.scala 46:47:@1932.4]
  wire [4:0] _T_56070; // @[Modules.scala 46:47:@1933.4]
  wire [5:0] _T_56072; // @[Modules.scala 46:37:@1935.4]
  wire [4:0] _T_56073; // @[Modules.scala 46:37:@1936.4]
  wire [4:0] _T_56074; // @[Modules.scala 46:37:@1937.4]
  wire [5:0] _T_56075; // @[Modules.scala 46:47:@1938.4]
  wire [4:0] _T_56076; // @[Modules.scala 46:47:@1939.4]
  wire [4:0] _T_56077; // @[Modules.scala 46:47:@1940.4]
  wire [5:0] _T_56079; // @[Modules.scala 46:37:@1942.4]
  wire [4:0] _T_56080; // @[Modules.scala 46:37:@1943.4]
  wire [4:0] _T_56081; // @[Modules.scala 46:37:@1944.4]
  wire [5:0] _T_56082; // @[Modules.scala 46:47:@1945.4]
  wire [4:0] _T_56083; // @[Modules.scala 46:47:@1946.4]
  wire [4:0] _T_56084; // @[Modules.scala 46:47:@1947.4]
  wire [5:0] _T_56086; // @[Modules.scala 46:37:@1949.4]
  wire [4:0] _T_56087; // @[Modules.scala 46:37:@1950.4]
  wire [4:0] _T_56088; // @[Modules.scala 46:37:@1951.4]
  wire [5:0] _T_56089; // @[Modules.scala 46:47:@1952.4]
  wire [4:0] _T_56090; // @[Modules.scala 46:47:@1953.4]
  wire [4:0] _T_56091; // @[Modules.scala 46:47:@1954.4]
  wire [5:0] _T_56093; // @[Modules.scala 46:37:@1956.4]
  wire [4:0] _T_56094; // @[Modules.scala 46:37:@1957.4]
  wire [4:0] _T_56095; // @[Modules.scala 46:37:@1958.4]
  wire [5:0] _T_56096; // @[Modules.scala 46:47:@1959.4]
  wire [4:0] _T_56097; // @[Modules.scala 46:47:@1960.4]
  wire [4:0] _T_56098; // @[Modules.scala 46:47:@1961.4]
  wire [5:0] _T_56100; // @[Modules.scala 43:37:@1963.4]
  wire [4:0] _T_56101; // @[Modules.scala 43:37:@1964.4]
  wire [4:0] _T_56102; // @[Modules.scala 43:37:@1965.4]
  wire [5:0] _T_56103; // @[Modules.scala 43:47:@1966.4]
  wire [4:0] _T_56104; // @[Modules.scala 43:47:@1967.4]
  wire [4:0] _T_56105; // @[Modules.scala 43:47:@1968.4]
  wire [5:0] _T_56106; // @[Modules.scala 37:46:@1970.4]
  wire [4:0] _T_56107; // @[Modules.scala 37:46:@1971.4]
  wire [4:0] _T_56108; // @[Modules.scala 37:46:@1972.4]
  wire [5:0] _T_56109; // @[Modules.scala 37:46:@1974.4]
  wire [4:0] _T_56110; // @[Modules.scala 37:46:@1975.4]
  wire [4:0] _T_56111; // @[Modules.scala 37:46:@1976.4]
  wire [5:0] _T_56112; // @[Modules.scala 37:46:@1978.4]
  wire [4:0] _T_56113; // @[Modules.scala 37:46:@1979.4]
  wire [4:0] _T_56114; // @[Modules.scala 37:46:@1980.4]
  wire [5:0] _T_56116; // @[Modules.scala 46:37:@1982.4]
  wire [4:0] _T_56117; // @[Modules.scala 46:37:@1983.4]
  wire [4:0] _T_56118; // @[Modules.scala 46:37:@1984.4]
  wire [5:0] _T_56119; // @[Modules.scala 46:47:@1985.4]
  wire [4:0] _T_56120; // @[Modules.scala 46:47:@1986.4]
  wire [4:0] _T_56121; // @[Modules.scala 46:47:@1987.4]
  wire [5:0] _T_56123; // @[Modules.scala 43:37:@1989.4]
  wire [4:0] _T_56124; // @[Modules.scala 43:37:@1990.4]
  wire [4:0] _T_56125; // @[Modules.scala 43:37:@1991.4]
  wire [5:0] _T_56126; // @[Modules.scala 43:47:@1992.4]
  wire [4:0] _T_56127; // @[Modules.scala 43:47:@1993.4]
  wire [4:0] _T_56128; // @[Modules.scala 43:47:@1994.4]
  wire [5:0] _T_56129; // @[Modules.scala 40:46:@1996.4]
  wire [4:0] _T_56130; // @[Modules.scala 40:46:@1997.4]
  wire [4:0] _T_56131; // @[Modules.scala 40:46:@1998.4]
  wire [5:0] _T_56132; // @[Modules.scala 37:46:@2000.4]
  wire [4:0] _T_56133; // @[Modules.scala 37:46:@2001.4]
  wire [4:0] _T_56134; // @[Modules.scala 37:46:@2002.4]
  wire [5:0] _T_56135; // @[Modules.scala 37:46:@2004.4]
  wire [4:0] _T_56136; // @[Modules.scala 37:46:@2005.4]
  wire [4:0] _T_56137; // @[Modules.scala 37:46:@2006.4]
  wire [5:0] _T_56138; // @[Modules.scala 37:46:@2008.4]
  wire [4:0] _T_56139; // @[Modules.scala 37:46:@2009.4]
  wire [4:0] _T_56140; // @[Modules.scala 37:46:@2010.4]
  wire [5:0] _T_56141; // @[Modules.scala 40:46:@2012.4]
  wire [4:0] _T_56142; // @[Modules.scala 40:46:@2013.4]
  wire [4:0] _T_56143; // @[Modules.scala 40:46:@2014.4]
  wire [5:0] _T_56145; // @[Modules.scala 46:37:@2016.4]
  wire [4:0] _T_56146; // @[Modules.scala 46:37:@2017.4]
  wire [4:0] _T_56147; // @[Modules.scala 46:37:@2018.4]
  wire [5:0] _T_56148; // @[Modules.scala 46:47:@2019.4]
  wire [4:0] _T_56149; // @[Modules.scala 46:47:@2020.4]
  wire [4:0] _T_56150; // @[Modules.scala 46:47:@2021.4]
  wire [5:0] _T_56152; // @[Modules.scala 46:37:@2023.4]
  wire [4:0] _T_56153; // @[Modules.scala 46:37:@2024.4]
  wire [4:0] _T_56154; // @[Modules.scala 46:37:@2025.4]
  wire [5:0] _T_56155; // @[Modules.scala 46:47:@2026.4]
  wire [4:0] _T_56156; // @[Modules.scala 46:47:@2027.4]
  wire [4:0] _T_56157; // @[Modules.scala 46:47:@2028.4]
  wire [5:0] _T_56158; // @[Modules.scala 37:46:@2030.4]
  wire [4:0] _T_56159; // @[Modules.scala 37:46:@2031.4]
  wire [4:0] _T_56160; // @[Modules.scala 37:46:@2032.4]
  wire [5:0] _T_56161; // @[Modules.scala 37:46:@2034.4]
  wire [4:0] _T_56162; // @[Modules.scala 37:46:@2035.4]
  wire [4:0] _T_56163; // @[Modules.scala 37:46:@2036.4]
  wire [5:0] _T_56164; // @[Modules.scala 37:46:@2038.4]
  wire [4:0] _T_56165; // @[Modules.scala 37:46:@2039.4]
  wire [4:0] _T_56166; // @[Modules.scala 37:46:@2040.4]
  wire [5:0] _T_56167; // @[Modules.scala 37:46:@2042.4]
  wire [4:0] _T_56168; // @[Modules.scala 37:46:@2043.4]
  wire [4:0] _T_56169; // @[Modules.scala 37:46:@2044.4]
  wire [5:0] _T_56170; // @[Modules.scala 37:46:@2046.4]
  wire [4:0] _T_56171; // @[Modules.scala 37:46:@2047.4]
  wire [4:0] _T_56172; // @[Modules.scala 37:46:@2048.4]
  wire [5:0] _T_56174; // @[Modules.scala 43:37:@2050.4]
  wire [4:0] _T_56175; // @[Modules.scala 43:37:@2051.4]
  wire [4:0] _T_56176; // @[Modules.scala 43:37:@2052.4]
  wire [5:0] _T_56177; // @[Modules.scala 43:47:@2053.4]
  wire [4:0] _T_56178; // @[Modules.scala 43:47:@2054.4]
  wire [4:0] _T_56179; // @[Modules.scala 43:47:@2055.4]
  wire [5:0] _T_56181; // @[Modules.scala 43:37:@2057.4]
  wire [4:0] _T_56182; // @[Modules.scala 43:37:@2058.4]
  wire [4:0] _T_56183; // @[Modules.scala 43:37:@2059.4]
  wire [5:0] _T_56184; // @[Modules.scala 43:47:@2060.4]
  wire [4:0] _T_56185; // @[Modules.scala 43:47:@2061.4]
  wire [4:0] _T_56186; // @[Modules.scala 43:47:@2062.4]
  wire [5:0] _T_56187; // @[Modules.scala 40:46:@2064.4]
  wire [4:0] _T_56188; // @[Modules.scala 40:46:@2065.4]
  wire [4:0] _T_56189; // @[Modules.scala 40:46:@2066.4]
  wire [5:0] _T_56190; // @[Modules.scala 37:46:@2068.4]
  wire [4:0] _T_56191; // @[Modules.scala 37:46:@2069.4]
  wire [4:0] _T_56192; // @[Modules.scala 37:46:@2070.4]
  wire [5:0] _T_56193; // @[Modules.scala 37:46:@2072.4]
  wire [4:0] _T_56194; // @[Modules.scala 37:46:@2073.4]
  wire [4:0] _T_56195; // @[Modules.scala 37:46:@2074.4]
  wire [5:0] _T_56196; // @[Modules.scala 37:46:@2076.4]
  wire [4:0] _T_56197; // @[Modules.scala 37:46:@2077.4]
  wire [4:0] _T_56198; // @[Modules.scala 37:46:@2078.4]
  wire [5:0] _T_56199; // @[Modules.scala 40:46:@2080.4]
  wire [4:0] _T_56200; // @[Modules.scala 40:46:@2081.4]
  wire [4:0] _T_56201; // @[Modules.scala 40:46:@2082.4]
  wire [5:0] _T_56202; // @[Modules.scala 37:46:@2084.4]
  wire [4:0] _T_56203; // @[Modules.scala 37:46:@2085.4]
  wire [4:0] _T_56204; // @[Modules.scala 37:46:@2086.4]
  wire [5:0] _T_56205; // @[Modules.scala 37:46:@2088.4]
  wire [4:0] _T_56206; // @[Modules.scala 37:46:@2089.4]
  wire [4:0] _T_56207; // @[Modules.scala 37:46:@2090.4]
  wire [5:0] _T_56208; // @[Modules.scala 37:46:@2092.4]
  wire [4:0] _T_56209; // @[Modules.scala 37:46:@2093.4]
  wire [4:0] _T_56210; // @[Modules.scala 37:46:@2094.4]
  wire [5:0] _T_56211; // @[Modules.scala 37:46:@2096.4]
  wire [4:0] _T_56212; // @[Modules.scala 37:46:@2097.4]
  wire [4:0] _T_56213; // @[Modules.scala 37:46:@2098.4]
  wire [5:0] _T_56214; // @[Modules.scala 37:46:@2100.4]
  wire [4:0] _T_56215; // @[Modules.scala 37:46:@2101.4]
  wire [4:0] _T_56216; // @[Modules.scala 37:46:@2102.4]
  wire [5:0] _T_56217; // @[Modules.scala 37:46:@2104.4]
  wire [4:0] _T_56218; // @[Modules.scala 37:46:@2105.4]
  wire [4:0] _T_56219; // @[Modules.scala 37:46:@2106.4]
  wire [5:0] _T_56220; // @[Modules.scala 40:46:@2108.4]
  wire [4:0] _T_56221; // @[Modules.scala 40:46:@2109.4]
  wire [4:0] _T_56222; // @[Modules.scala 40:46:@2110.4]
  wire [5:0] _T_56224; // @[Modules.scala 46:37:@2112.4]
  wire [4:0] _T_56225; // @[Modules.scala 46:37:@2113.4]
  wire [4:0] _T_56226; // @[Modules.scala 46:37:@2114.4]
  wire [5:0] _T_56227; // @[Modules.scala 46:47:@2115.4]
  wire [4:0] _T_56228; // @[Modules.scala 46:47:@2116.4]
  wire [4:0] _T_56229; // @[Modules.scala 46:47:@2117.4]
  wire [5:0] _T_56230; // @[Modules.scala 40:46:@2119.4]
  wire [4:0] _T_56231; // @[Modules.scala 40:46:@2120.4]
  wire [4:0] _T_56232; // @[Modules.scala 40:46:@2121.4]
  wire [5:0] _T_56234; // @[Modules.scala 43:37:@2123.4]
  wire [4:0] _T_56235; // @[Modules.scala 43:37:@2124.4]
  wire [4:0] _T_56236; // @[Modules.scala 43:37:@2125.4]
  wire [5:0] _T_56237; // @[Modules.scala 43:47:@2126.4]
  wire [4:0] _T_56238; // @[Modules.scala 43:47:@2127.4]
  wire [4:0] _T_56239; // @[Modules.scala 43:47:@2128.4]
  wire [5:0] _T_56240; // @[Modules.scala 37:46:@2130.4]
  wire [4:0] _T_56241; // @[Modules.scala 37:46:@2131.4]
  wire [4:0] _T_56242; // @[Modules.scala 37:46:@2132.4]
  wire [5:0] _T_56243; // @[Modules.scala 37:46:@2134.4]
  wire [4:0] _T_56244; // @[Modules.scala 37:46:@2135.4]
  wire [4:0] _T_56245; // @[Modules.scala 37:46:@2136.4]
  wire [5:0] _T_56247; // @[Modules.scala 46:37:@2138.4]
  wire [4:0] _T_56248; // @[Modules.scala 46:37:@2139.4]
  wire [4:0] _T_56249; // @[Modules.scala 46:37:@2140.4]
  wire [5:0] _T_56250; // @[Modules.scala 46:47:@2141.4]
  wire [4:0] _T_56251; // @[Modules.scala 46:47:@2142.4]
  wire [4:0] _T_56252; // @[Modules.scala 46:47:@2143.4]
  wire [5:0] _T_56254; // @[Modules.scala 46:37:@2145.4]
  wire [4:0] _T_56255; // @[Modules.scala 46:37:@2146.4]
  wire [4:0] _T_56256; // @[Modules.scala 46:37:@2147.4]
  wire [5:0] _T_56257; // @[Modules.scala 46:47:@2148.4]
  wire [4:0] _T_56258; // @[Modules.scala 46:47:@2149.4]
  wire [4:0] _T_56259; // @[Modules.scala 46:47:@2150.4]
  wire [5:0] _T_56260; // @[Modules.scala 40:46:@2152.4]
  wire [4:0] _T_56261; // @[Modules.scala 40:46:@2153.4]
  wire [4:0] _T_56262; // @[Modules.scala 40:46:@2154.4]
  wire [5:0] _T_56263; // @[Modules.scala 40:46:@2156.4]
  wire [4:0] _T_56264; // @[Modules.scala 40:46:@2157.4]
  wire [4:0] _T_56265; // @[Modules.scala 40:46:@2158.4]
  wire [5:0] _T_56267; // @[Modules.scala 46:37:@2160.4]
  wire [4:0] _T_56268; // @[Modules.scala 46:37:@2161.4]
  wire [4:0] _T_56269; // @[Modules.scala 46:37:@2162.4]
  wire [5:0] _T_56270; // @[Modules.scala 46:47:@2163.4]
  wire [4:0] _T_56271; // @[Modules.scala 46:47:@2164.4]
  wire [4:0] _T_56272; // @[Modules.scala 46:47:@2165.4]
  wire [5:0] _T_56274; // @[Modules.scala 46:37:@2167.4]
  wire [4:0] _T_56275; // @[Modules.scala 46:37:@2168.4]
  wire [4:0] _T_56276; // @[Modules.scala 46:37:@2169.4]
  wire [5:0] _T_56277; // @[Modules.scala 46:47:@2170.4]
  wire [4:0] _T_56278; // @[Modules.scala 46:47:@2171.4]
  wire [4:0] _T_56279; // @[Modules.scala 46:47:@2172.4]
  wire [5:0] _T_56280; // @[Modules.scala 37:46:@2174.4]
  wire [4:0] _T_56281; // @[Modules.scala 37:46:@2175.4]
  wire [4:0] _T_56282; // @[Modules.scala 37:46:@2176.4]
  wire [5:0] _T_56283; // @[Modules.scala 40:46:@2178.4]
  wire [4:0] _T_56284; // @[Modules.scala 40:46:@2179.4]
  wire [4:0] _T_56285; // @[Modules.scala 40:46:@2180.4]
  wire [5:0] _T_56286; // @[Modules.scala 37:46:@2182.4]
  wire [4:0] _T_56287; // @[Modules.scala 37:46:@2183.4]
  wire [4:0] _T_56288; // @[Modules.scala 37:46:@2184.4]
  wire [5:0] _T_56289; // @[Modules.scala 37:46:@2186.4]
  wire [4:0] _T_56290; // @[Modules.scala 37:46:@2187.4]
  wire [4:0] _T_56291; // @[Modules.scala 37:46:@2188.4]
  wire [5:0] _T_56293; // @[Modules.scala 43:37:@2190.4]
  wire [4:0] _T_56294; // @[Modules.scala 43:37:@2191.4]
  wire [4:0] _T_56295; // @[Modules.scala 43:37:@2192.4]
  wire [5:0] _T_56296; // @[Modules.scala 43:47:@2193.4]
  wire [4:0] _T_56297; // @[Modules.scala 43:47:@2194.4]
  wire [4:0] _T_56298; // @[Modules.scala 43:47:@2195.4]
  wire [5:0] _T_56300; // @[Modules.scala 46:37:@2197.4]
  wire [4:0] _T_56301; // @[Modules.scala 46:37:@2198.4]
  wire [4:0] _T_56302; // @[Modules.scala 46:37:@2199.4]
  wire [5:0] _T_56303; // @[Modules.scala 46:47:@2200.4]
  wire [4:0] _T_56304; // @[Modules.scala 46:47:@2201.4]
  wire [4:0] _T_56305; // @[Modules.scala 46:47:@2202.4]
  wire [5:0] _T_56306; // @[Modules.scala 40:46:@2204.4]
  wire [4:0] _T_56307; // @[Modules.scala 40:46:@2205.4]
  wire [4:0] _T_56308; // @[Modules.scala 40:46:@2206.4]
  wire [5:0] _T_56310; // @[Modules.scala 46:37:@2208.4]
  wire [4:0] _T_56311; // @[Modules.scala 46:37:@2209.4]
  wire [4:0] _T_56312; // @[Modules.scala 46:37:@2210.4]
  wire [5:0] _T_56313; // @[Modules.scala 46:47:@2211.4]
  wire [4:0] _T_56314; // @[Modules.scala 46:47:@2212.4]
  wire [4:0] _T_56315; // @[Modules.scala 46:47:@2213.4]
  wire [5:0] _T_56317; // @[Modules.scala 46:37:@2215.4]
  wire [4:0] _T_56318; // @[Modules.scala 46:37:@2216.4]
  wire [4:0] _T_56319; // @[Modules.scala 46:37:@2217.4]
  wire [5:0] _T_56320; // @[Modules.scala 46:47:@2218.4]
  wire [4:0] _T_56321; // @[Modules.scala 46:47:@2219.4]
  wire [4:0] _T_56322; // @[Modules.scala 46:47:@2220.4]
  wire [5:0] _T_56324; // @[Modules.scala 46:37:@2222.4]
  wire [4:0] _T_56325; // @[Modules.scala 46:37:@2223.4]
  wire [4:0] _T_56326; // @[Modules.scala 46:37:@2224.4]
  wire [5:0] _T_56327; // @[Modules.scala 46:47:@2225.4]
  wire [4:0] _T_56328; // @[Modules.scala 46:47:@2226.4]
  wire [4:0] _T_56329; // @[Modules.scala 46:47:@2227.4]
  wire [5:0] _T_56330; // @[Modules.scala 40:46:@2229.4]
  wire [4:0] _T_56331; // @[Modules.scala 40:46:@2230.4]
  wire [4:0] _T_56332; // @[Modules.scala 40:46:@2231.4]
  wire [5:0] _T_56334; // @[Modules.scala 43:37:@2233.4]
  wire [4:0] _T_56335; // @[Modules.scala 43:37:@2234.4]
  wire [4:0] _T_56336; // @[Modules.scala 43:37:@2235.4]
  wire [5:0] _T_56337; // @[Modules.scala 43:47:@2236.4]
  wire [4:0] _T_56338; // @[Modules.scala 43:47:@2237.4]
  wire [4:0] _T_56339; // @[Modules.scala 43:47:@2238.4]
  wire [5:0] _T_56341; // @[Modules.scala 46:37:@2240.4]
  wire [4:0] _T_56342; // @[Modules.scala 46:37:@2241.4]
  wire [4:0] _T_56343; // @[Modules.scala 46:37:@2242.4]
  wire [5:0] _T_56344; // @[Modules.scala 46:47:@2243.4]
  wire [4:0] _T_56345; // @[Modules.scala 46:47:@2244.4]
  wire [4:0] _T_56346; // @[Modules.scala 46:47:@2245.4]
  wire [5:0] _T_56348; // @[Modules.scala 46:37:@2247.4]
  wire [4:0] _T_56349; // @[Modules.scala 46:37:@2248.4]
  wire [4:0] _T_56350; // @[Modules.scala 46:37:@2249.4]
  wire [5:0] _T_56351; // @[Modules.scala 46:47:@2250.4]
  wire [4:0] _T_56352; // @[Modules.scala 46:47:@2251.4]
  wire [4:0] _T_56353; // @[Modules.scala 46:47:@2252.4]
  wire [5:0] _T_56354; // @[Modules.scala 37:46:@2254.4]
  wire [4:0] _T_56355; // @[Modules.scala 37:46:@2255.4]
  wire [4:0] _T_56356; // @[Modules.scala 37:46:@2256.4]
  wire [5:0] _T_56358; // @[Modules.scala 46:37:@2258.4]
  wire [4:0] _T_56359; // @[Modules.scala 46:37:@2259.4]
  wire [4:0] _T_56360; // @[Modules.scala 46:37:@2260.4]
  wire [5:0] _T_56361; // @[Modules.scala 46:47:@2261.4]
  wire [4:0] _T_56362; // @[Modules.scala 46:47:@2262.4]
  wire [4:0] _T_56363; // @[Modules.scala 46:47:@2263.4]
  wire [5:0] _T_56365; // @[Modules.scala 43:37:@2265.4]
  wire [4:0] _T_56366; // @[Modules.scala 43:37:@2266.4]
  wire [4:0] _T_56367; // @[Modules.scala 43:37:@2267.4]
  wire [5:0] _T_56368; // @[Modules.scala 43:47:@2268.4]
  wire [4:0] _T_56369; // @[Modules.scala 43:47:@2269.4]
  wire [4:0] _T_56370; // @[Modules.scala 43:47:@2270.4]
  wire [5:0] _T_56371; // @[Modules.scala 37:46:@2272.4]
  wire [4:0] _T_56372; // @[Modules.scala 37:46:@2273.4]
  wire [4:0] _T_56373; // @[Modules.scala 37:46:@2274.4]
  wire [10:0] buffer_0_0; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56374; // @[Modules.scala 50:57:@2276.4]
  wire [10:0] _T_56375; // @[Modules.scala 50:57:@2277.4]
  wire [10:0] buffer_0_392; // @[Modules.scala 50:57:@2278.4]
  wire [10:0] buffer_0_2; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_3; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56377; // @[Modules.scala 50:57:@2280.4]
  wire [10:0] _T_56378; // @[Modules.scala 50:57:@2281.4]
  wire [10:0] buffer_0_393; // @[Modules.scala 50:57:@2282.4]
  wire [10:0] buffer_0_4; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56380; // @[Modules.scala 50:57:@2284.4]
  wire [10:0] _T_56381; // @[Modules.scala 50:57:@2285.4]
  wire [10:0] buffer_0_394; // @[Modules.scala 50:57:@2286.4]
  wire [10:0] buffer_0_6; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_7; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56383; // @[Modules.scala 50:57:@2288.4]
  wire [10:0] _T_56384; // @[Modules.scala 50:57:@2289.4]
  wire [10:0] buffer_0_395; // @[Modules.scala 50:57:@2290.4]
  wire [10:0] buffer_0_8; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56386; // @[Modules.scala 50:57:@2292.4]
  wire [10:0] _T_56387; // @[Modules.scala 50:57:@2293.4]
  wire [10:0] buffer_0_396; // @[Modules.scala 50:57:@2294.4]
  wire [10:0] buffer_0_10; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56389; // @[Modules.scala 50:57:@2296.4]
  wire [10:0] _T_56390; // @[Modules.scala 50:57:@2297.4]
  wire [10:0] buffer_0_397; // @[Modules.scala 50:57:@2298.4]
  wire [10:0] buffer_0_12; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56392; // @[Modules.scala 50:57:@2300.4]
  wire [10:0] _T_56393; // @[Modules.scala 50:57:@2301.4]
  wire [10:0] buffer_0_398; // @[Modules.scala 50:57:@2302.4]
  wire [10:0] buffer_0_14; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56395; // @[Modules.scala 50:57:@2304.4]
  wire [10:0] _T_56396; // @[Modules.scala 50:57:@2305.4]
  wire [10:0] buffer_0_399; // @[Modules.scala 50:57:@2306.4]
  wire [10:0] buffer_0_16; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_17; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56398; // @[Modules.scala 50:57:@2308.4]
  wire [10:0] _T_56399; // @[Modules.scala 50:57:@2309.4]
  wire [10:0] buffer_0_400; // @[Modules.scala 50:57:@2310.4]
  wire [10:0] buffer_0_18; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_19; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56401; // @[Modules.scala 50:57:@2312.4]
  wire [10:0] _T_56402; // @[Modules.scala 50:57:@2313.4]
  wire [10:0] buffer_0_401; // @[Modules.scala 50:57:@2314.4]
  wire [10:0] buffer_0_20; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_21; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56404; // @[Modules.scala 50:57:@2316.4]
  wire [10:0] _T_56405; // @[Modules.scala 50:57:@2317.4]
  wire [10:0] buffer_0_402; // @[Modules.scala 50:57:@2318.4]
  wire [10:0] buffer_0_22; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_23; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56407; // @[Modules.scala 50:57:@2320.4]
  wire [10:0] _T_56408; // @[Modules.scala 50:57:@2321.4]
  wire [10:0] buffer_0_403; // @[Modules.scala 50:57:@2322.4]
  wire [10:0] buffer_0_24; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_25; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56410; // @[Modules.scala 50:57:@2324.4]
  wire [10:0] _T_56411; // @[Modules.scala 50:57:@2325.4]
  wire [10:0] buffer_0_404; // @[Modules.scala 50:57:@2326.4]
  wire [10:0] buffer_0_26; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56413; // @[Modules.scala 50:57:@2328.4]
  wire [10:0] _T_56414; // @[Modules.scala 50:57:@2329.4]
  wire [10:0] buffer_0_405; // @[Modules.scala 50:57:@2330.4]
  wire [10:0] buffer_0_28; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56416; // @[Modules.scala 50:57:@2332.4]
  wire [10:0] _T_56417; // @[Modules.scala 50:57:@2333.4]
  wire [10:0] buffer_0_406; // @[Modules.scala 50:57:@2334.4]
  wire [10:0] buffer_0_30; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_31; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56419; // @[Modules.scala 50:57:@2336.4]
  wire [10:0] _T_56420; // @[Modules.scala 50:57:@2337.4]
  wire [10:0] buffer_0_407; // @[Modules.scala 50:57:@2338.4]
  wire [10:0] buffer_0_32; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_33; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56422; // @[Modules.scala 50:57:@2340.4]
  wire [10:0] _T_56423; // @[Modules.scala 50:57:@2341.4]
  wire [10:0] buffer_0_408; // @[Modules.scala 50:57:@2342.4]
  wire [10:0] buffer_0_34; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56425; // @[Modules.scala 50:57:@2344.4]
  wire [10:0] _T_56426; // @[Modules.scala 50:57:@2345.4]
  wire [10:0] buffer_0_409; // @[Modules.scala 50:57:@2346.4]
  wire [10:0] buffer_0_36; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_37; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56428; // @[Modules.scala 50:57:@2348.4]
  wire [10:0] _T_56429; // @[Modules.scala 50:57:@2349.4]
  wire [10:0] buffer_0_410; // @[Modules.scala 50:57:@2350.4]
  wire [10:0] buffer_0_38; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_39; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56431; // @[Modules.scala 50:57:@2352.4]
  wire [10:0] _T_56432; // @[Modules.scala 50:57:@2353.4]
  wire [10:0] buffer_0_411; // @[Modules.scala 50:57:@2354.4]
  wire [10:0] buffer_0_40; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56434; // @[Modules.scala 50:57:@2356.4]
  wire [10:0] _T_56435; // @[Modules.scala 50:57:@2357.4]
  wire [10:0] buffer_0_412; // @[Modules.scala 50:57:@2358.4]
  wire [10:0] buffer_0_42; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56437; // @[Modules.scala 50:57:@2360.4]
  wire [10:0] _T_56438; // @[Modules.scala 50:57:@2361.4]
  wire [10:0] buffer_0_413; // @[Modules.scala 50:57:@2362.4]
  wire [10:0] buffer_0_44; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_45; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56440; // @[Modules.scala 50:57:@2364.4]
  wire [10:0] _T_56441; // @[Modules.scala 50:57:@2365.4]
  wire [10:0] buffer_0_414; // @[Modules.scala 50:57:@2366.4]
  wire [10:0] buffer_0_46; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_47; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56443; // @[Modules.scala 50:57:@2368.4]
  wire [10:0] _T_56444; // @[Modules.scala 50:57:@2369.4]
  wire [10:0] buffer_0_415; // @[Modules.scala 50:57:@2370.4]
  wire [10:0] buffer_0_48; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_49; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56446; // @[Modules.scala 50:57:@2372.4]
  wire [10:0] _T_56447; // @[Modules.scala 50:57:@2373.4]
  wire [10:0] buffer_0_416; // @[Modules.scala 50:57:@2374.4]
  wire [10:0] buffer_0_50; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_51; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56449; // @[Modules.scala 50:57:@2376.4]
  wire [10:0] _T_56450; // @[Modules.scala 50:57:@2377.4]
  wire [10:0] buffer_0_417; // @[Modules.scala 50:57:@2378.4]
  wire [10:0] buffer_0_52; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_53; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56452; // @[Modules.scala 50:57:@2380.4]
  wire [10:0] _T_56453; // @[Modules.scala 50:57:@2381.4]
  wire [10:0] buffer_0_418; // @[Modules.scala 50:57:@2382.4]
  wire [10:0] buffer_0_54; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56455; // @[Modules.scala 50:57:@2384.4]
  wire [10:0] _T_56456; // @[Modules.scala 50:57:@2385.4]
  wire [10:0] buffer_0_419; // @[Modules.scala 50:57:@2386.4]
  wire [10:0] buffer_0_56; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56458; // @[Modules.scala 50:57:@2388.4]
  wire [10:0] _T_56459; // @[Modules.scala 50:57:@2389.4]
  wire [10:0] buffer_0_420; // @[Modules.scala 50:57:@2390.4]
  wire [10:0] buffer_0_58; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_59; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56461; // @[Modules.scala 50:57:@2392.4]
  wire [10:0] _T_56462; // @[Modules.scala 50:57:@2393.4]
  wire [10:0] buffer_0_421; // @[Modules.scala 50:57:@2394.4]
  wire [10:0] buffer_0_60; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56464; // @[Modules.scala 50:57:@2396.4]
  wire [10:0] _T_56465; // @[Modules.scala 50:57:@2397.4]
  wire [10:0] buffer_0_422; // @[Modules.scala 50:57:@2398.4]
  wire [10:0] buffer_0_62; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56467; // @[Modules.scala 50:57:@2400.4]
  wire [10:0] _T_56468; // @[Modules.scala 50:57:@2401.4]
  wire [10:0] buffer_0_423; // @[Modules.scala 50:57:@2402.4]
  wire [10:0] buffer_0_64; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_65; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56470; // @[Modules.scala 50:57:@2404.4]
  wire [10:0] _T_56471; // @[Modules.scala 50:57:@2405.4]
  wire [10:0] buffer_0_424; // @[Modules.scala 50:57:@2406.4]
  wire [10:0] buffer_0_66; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_67; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56473; // @[Modules.scala 50:57:@2408.4]
  wire [10:0] _T_56474; // @[Modules.scala 50:57:@2409.4]
  wire [10:0] buffer_0_425; // @[Modules.scala 50:57:@2410.4]
  wire [10:0] buffer_0_68; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56476; // @[Modules.scala 50:57:@2412.4]
  wire [10:0] _T_56477; // @[Modules.scala 50:57:@2413.4]
  wire [10:0] buffer_0_426; // @[Modules.scala 50:57:@2414.4]
  wire [10:0] buffer_0_70; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56479; // @[Modules.scala 50:57:@2416.4]
  wire [10:0] _T_56480; // @[Modules.scala 50:57:@2417.4]
  wire [10:0] buffer_0_427; // @[Modules.scala 50:57:@2418.4]
  wire [10:0] buffer_0_72; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56482; // @[Modules.scala 50:57:@2420.4]
  wire [10:0] _T_56483; // @[Modules.scala 50:57:@2421.4]
  wire [10:0] buffer_0_428; // @[Modules.scala 50:57:@2422.4]
  wire [10:0] buffer_0_74; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56485; // @[Modules.scala 50:57:@2424.4]
  wire [10:0] _T_56486; // @[Modules.scala 50:57:@2425.4]
  wire [10:0] buffer_0_429; // @[Modules.scala 50:57:@2426.4]
  wire [10:0] buffer_0_76; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_77; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56488; // @[Modules.scala 50:57:@2428.4]
  wire [10:0] _T_56489; // @[Modules.scala 50:57:@2429.4]
  wire [10:0] buffer_0_430; // @[Modules.scala 50:57:@2430.4]
  wire [10:0] buffer_0_78; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56491; // @[Modules.scala 50:57:@2432.4]
  wire [10:0] _T_56492; // @[Modules.scala 50:57:@2433.4]
  wire [10:0] buffer_0_431; // @[Modules.scala 50:57:@2434.4]
  wire [10:0] buffer_0_80; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_81; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56494; // @[Modules.scala 50:57:@2436.4]
  wire [10:0] _T_56495; // @[Modules.scala 50:57:@2437.4]
  wire [10:0] buffer_0_432; // @[Modules.scala 50:57:@2438.4]
  wire [10:0] buffer_0_82; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56497; // @[Modules.scala 50:57:@2440.4]
  wire [10:0] _T_56498; // @[Modules.scala 50:57:@2441.4]
  wire [10:0] buffer_0_433; // @[Modules.scala 50:57:@2442.4]
  wire [10:0] buffer_0_84; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56500; // @[Modules.scala 50:57:@2444.4]
  wire [10:0] _T_56501; // @[Modules.scala 50:57:@2445.4]
  wire [10:0] buffer_0_434; // @[Modules.scala 50:57:@2446.4]
  wire [10:0] buffer_0_86; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56503; // @[Modules.scala 50:57:@2448.4]
  wire [10:0] _T_56504; // @[Modules.scala 50:57:@2449.4]
  wire [10:0] buffer_0_435; // @[Modules.scala 50:57:@2450.4]
  wire [10:0] buffer_0_88; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56506; // @[Modules.scala 50:57:@2452.4]
  wire [10:0] _T_56507; // @[Modules.scala 50:57:@2453.4]
  wire [10:0] buffer_0_436; // @[Modules.scala 50:57:@2454.4]
  wire [10:0] buffer_0_90; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56509; // @[Modules.scala 50:57:@2456.4]
  wire [10:0] _T_56510; // @[Modules.scala 50:57:@2457.4]
  wire [10:0] buffer_0_437; // @[Modules.scala 50:57:@2458.4]
  wire [10:0] buffer_0_92; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56512; // @[Modules.scala 50:57:@2460.4]
  wire [10:0] _T_56513; // @[Modules.scala 50:57:@2461.4]
  wire [10:0] buffer_0_438; // @[Modules.scala 50:57:@2462.4]
  wire [10:0] buffer_0_94; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56515; // @[Modules.scala 50:57:@2464.4]
  wire [10:0] _T_56516; // @[Modules.scala 50:57:@2465.4]
  wire [10:0] buffer_0_439; // @[Modules.scala 50:57:@2466.4]
  wire [10:0] buffer_0_96; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56518; // @[Modules.scala 50:57:@2468.4]
  wire [10:0] _T_56519; // @[Modules.scala 50:57:@2469.4]
  wire [10:0] buffer_0_440; // @[Modules.scala 50:57:@2470.4]
  wire [10:0] buffer_0_98; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56521; // @[Modules.scala 50:57:@2472.4]
  wire [10:0] _T_56522; // @[Modules.scala 50:57:@2473.4]
  wire [10:0] buffer_0_441; // @[Modules.scala 50:57:@2474.4]
  wire [10:0] buffer_0_100; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56524; // @[Modules.scala 50:57:@2476.4]
  wire [10:0] _T_56525; // @[Modules.scala 50:57:@2477.4]
  wire [10:0] buffer_0_442; // @[Modules.scala 50:57:@2478.4]
  wire [10:0] buffer_0_102; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56527; // @[Modules.scala 50:57:@2480.4]
  wire [10:0] _T_56528; // @[Modules.scala 50:57:@2481.4]
  wire [10:0] buffer_0_443; // @[Modules.scala 50:57:@2482.4]
  wire [10:0] buffer_0_104; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56530; // @[Modules.scala 50:57:@2484.4]
  wire [10:0] _T_56531; // @[Modules.scala 50:57:@2485.4]
  wire [10:0] buffer_0_444; // @[Modules.scala 50:57:@2486.4]
  wire [10:0] buffer_0_106; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56533; // @[Modules.scala 50:57:@2488.4]
  wire [10:0] _T_56534; // @[Modules.scala 50:57:@2489.4]
  wire [10:0] buffer_0_445; // @[Modules.scala 50:57:@2490.4]
  wire [10:0] buffer_0_108; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56536; // @[Modules.scala 50:57:@2492.4]
  wire [10:0] _T_56537; // @[Modules.scala 50:57:@2493.4]
  wire [10:0] buffer_0_446; // @[Modules.scala 50:57:@2494.4]
  wire [10:0] buffer_0_110; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56539; // @[Modules.scala 50:57:@2496.4]
  wire [10:0] _T_56540; // @[Modules.scala 50:57:@2497.4]
  wire [10:0] buffer_0_447; // @[Modules.scala 50:57:@2498.4]
  wire [10:0] buffer_0_112; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56542; // @[Modules.scala 50:57:@2500.4]
  wire [10:0] _T_56543; // @[Modules.scala 50:57:@2501.4]
  wire [10:0] buffer_0_448; // @[Modules.scala 50:57:@2502.4]
  wire [10:0] buffer_0_114; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56545; // @[Modules.scala 50:57:@2504.4]
  wire [10:0] _T_56546; // @[Modules.scala 50:57:@2505.4]
  wire [10:0] buffer_0_449; // @[Modules.scala 50:57:@2506.4]
  wire [10:0] buffer_0_116; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56548; // @[Modules.scala 50:57:@2508.4]
  wire [10:0] _T_56549; // @[Modules.scala 50:57:@2509.4]
  wire [10:0] buffer_0_450; // @[Modules.scala 50:57:@2510.4]
  wire [10:0] buffer_0_118; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56551; // @[Modules.scala 50:57:@2512.4]
  wire [10:0] _T_56552; // @[Modules.scala 50:57:@2513.4]
  wire [10:0] buffer_0_451; // @[Modules.scala 50:57:@2514.4]
  wire [10:0] buffer_0_120; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56554; // @[Modules.scala 50:57:@2516.4]
  wire [10:0] _T_56555; // @[Modules.scala 50:57:@2517.4]
  wire [10:0] buffer_0_452; // @[Modules.scala 50:57:@2518.4]
  wire [10:0] buffer_0_122; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56557; // @[Modules.scala 50:57:@2520.4]
  wire [10:0] _T_56558; // @[Modules.scala 50:57:@2521.4]
  wire [10:0] buffer_0_453; // @[Modules.scala 50:57:@2522.4]
  wire [10:0] buffer_0_124; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_125; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56560; // @[Modules.scala 50:57:@2524.4]
  wire [10:0] _T_56561; // @[Modules.scala 50:57:@2525.4]
  wire [10:0] buffer_0_454; // @[Modules.scala 50:57:@2526.4]
  wire [10:0] buffer_0_126; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_127; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56563; // @[Modules.scala 50:57:@2528.4]
  wire [10:0] _T_56564; // @[Modules.scala 50:57:@2529.4]
  wire [10:0] buffer_0_455; // @[Modules.scala 50:57:@2530.4]
  wire [10:0] buffer_0_128; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56566; // @[Modules.scala 50:57:@2532.4]
  wire [10:0] _T_56567; // @[Modules.scala 50:57:@2533.4]
  wire [10:0] buffer_0_456; // @[Modules.scala 50:57:@2534.4]
  wire [10:0] buffer_0_130; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56569; // @[Modules.scala 50:57:@2536.4]
  wire [10:0] _T_56570; // @[Modules.scala 50:57:@2537.4]
  wire [10:0] buffer_0_457; // @[Modules.scala 50:57:@2538.4]
  wire [10:0] buffer_0_132; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_133; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56572; // @[Modules.scala 50:57:@2540.4]
  wire [10:0] _T_56573; // @[Modules.scala 50:57:@2541.4]
  wire [10:0] buffer_0_458; // @[Modules.scala 50:57:@2542.4]
  wire [10:0] buffer_0_134; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56575; // @[Modules.scala 50:57:@2544.4]
  wire [10:0] _T_56576; // @[Modules.scala 50:57:@2545.4]
  wire [10:0] buffer_0_459; // @[Modules.scala 50:57:@2546.4]
  wire [10:0] buffer_0_136; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56578; // @[Modules.scala 50:57:@2548.4]
  wire [10:0] _T_56579; // @[Modules.scala 50:57:@2549.4]
  wire [10:0] buffer_0_460; // @[Modules.scala 50:57:@2550.4]
  wire [10:0] buffer_0_138; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_139; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56581; // @[Modules.scala 50:57:@2552.4]
  wire [10:0] _T_56582; // @[Modules.scala 50:57:@2553.4]
  wire [10:0] buffer_0_461; // @[Modules.scala 50:57:@2554.4]
  wire [10:0] buffer_0_140; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56584; // @[Modules.scala 50:57:@2556.4]
  wire [10:0] _T_56585; // @[Modules.scala 50:57:@2557.4]
  wire [10:0] buffer_0_462; // @[Modules.scala 50:57:@2558.4]
  wire [10:0] buffer_0_142; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56587; // @[Modules.scala 50:57:@2560.4]
  wire [10:0] _T_56588; // @[Modules.scala 50:57:@2561.4]
  wire [10:0] buffer_0_463; // @[Modules.scala 50:57:@2562.4]
  wire [10:0] buffer_0_144; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56590; // @[Modules.scala 50:57:@2564.4]
  wire [10:0] _T_56591; // @[Modules.scala 50:57:@2565.4]
  wire [10:0] buffer_0_464; // @[Modules.scala 50:57:@2566.4]
  wire [10:0] buffer_0_146; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56593; // @[Modules.scala 50:57:@2568.4]
  wire [10:0] _T_56594; // @[Modules.scala 50:57:@2569.4]
  wire [10:0] buffer_0_465; // @[Modules.scala 50:57:@2570.4]
  wire [10:0] buffer_0_148; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_149; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56596; // @[Modules.scala 50:57:@2572.4]
  wire [10:0] _T_56597; // @[Modules.scala 50:57:@2573.4]
  wire [10:0] buffer_0_466; // @[Modules.scala 50:57:@2574.4]
  wire [10:0] buffer_0_150; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56599; // @[Modules.scala 50:57:@2576.4]
  wire [10:0] _T_56600; // @[Modules.scala 50:57:@2577.4]
  wire [10:0] buffer_0_467; // @[Modules.scala 50:57:@2578.4]
  wire [10:0] buffer_0_152; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_153; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56602; // @[Modules.scala 50:57:@2580.4]
  wire [10:0] _T_56603; // @[Modules.scala 50:57:@2581.4]
  wire [10:0] buffer_0_468; // @[Modules.scala 50:57:@2582.4]
  wire [10:0] buffer_0_154; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56605; // @[Modules.scala 50:57:@2584.4]
  wire [10:0] _T_56606; // @[Modules.scala 50:57:@2585.4]
  wire [10:0] buffer_0_469; // @[Modules.scala 50:57:@2586.4]
  wire [10:0] buffer_0_156; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56608; // @[Modules.scala 50:57:@2588.4]
  wire [10:0] _T_56609; // @[Modules.scala 50:57:@2589.4]
  wire [10:0] buffer_0_470; // @[Modules.scala 50:57:@2590.4]
  wire [10:0] buffer_0_158; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_159; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56611; // @[Modules.scala 50:57:@2592.4]
  wire [10:0] _T_56612; // @[Modules.scala 50:57:@2593.4]
  wire [10:0] buffer_0_471; // @[Modules.scala 50:57:@2594.4]
  wire [10:0] buffer_0_160; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56614; // @[Modules.scala 50:57:@2596.4]
  wire [10:0] _T_56615; // @[Modules.scala 50:57:@2597.4]
  wire [10:0] buffer_0_472; // @[Modules.scala 50:57:@2598.4]
  wire [10:0] buffer_0_162; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_163; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56617; // @[Modules.scala 50:57:@2600.4]
  wire [10:0] _T_56618; // @[Modules.scala 50:57:@2601.4]
  wire [10:0] buffer_0_473; // @[Modules.scala 50:57:@2602.4]
  wire [10:0] buffer_0_164; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_165; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56620; // @[Modules.scala 50:57:@2604.4]
  wire [10:0] _T_56621; // @[Modules.scala 50:57:@2605.4]
  wire [10:0] buffer_0_474; // @[Modules.scala 50:57:@2606.4]
  wire [10:0] buffer_0_166; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56623; // @[Modules.scala 50:57:@2608.4]
  wire [10:0] _T_56624; // @[Modules.scala 50:57:@2609.4]
  wire [10:0] buffer_0_475; // @[Modules.scala 50:57:@2610.4]
  wire [10:0] buffer_0_168; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56626; // @[Modules.scala 50:57:@2612.4]
  wire [10:0] _T_56627; // @[Modules.scala 50:57:@2613.4]
  wire [10:0] buffer_0_476; // @[Modules.scala 50:57:@2614.4]
  wire [10:0] buffer_0_170; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56629; // @[Modules.scala 50:57:@2616.4]
  wire [10:0] _T_56630; // @[Modules.scala 50:57:@2617.4]
  wire [10:0] buffer_0_477; // @[Modules.scala 50:57:@2618.4]
  wire [10:0] buffer_0_172; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56632; // @[Modules.scala 50:57:@2620.4]
  wire [10:0] _T_56633; // @[Modules.scala 50:57:@2621.4]
  wire [10:0] buffer_0_478; // @[Modules.scala 50:57:@2622.4]
  wire [10:0] buffer_0_174; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_175; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56635; // @[Modules.scala 50:57:@2624.4]
  wire [10:0] _T_56636; // @[Modules.scala 50:57:@2625.4]
  wire [10:0] buffer_0_479; // @[Modules.scala 50:57:@2626.4]
  wire [10:0] buffer_0_176; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56638; // @[Modules.scala 50:57:@2628.4]
  wire [10:0] _T_56639; // @[Modules.scala 50:57:@2629.4]
  wire [10:0] buffer_0_480; // @[Modules.scala 50:57:@2630.4]
  wire [10:0] buffer_0_178; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56641; // @[Modules.scala 50:57:@2632.4]
  wire [10:0] _T_56642; // @[Modules.scala 50:57:@2633.4]
  wire [10:0] buffer_0_481; // @[Modules.scala 50:57:@2634.4]
  wire [10:0] buffer_0_180; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56644; // @[Modules.scala 50:57:@2636.4]
  wire [10:0] _T_56645; // @[Modules.scala 50:57:@2637.4]
  wire [10:0] buffer_0_482; // @[Modules.scala 50:57:@2638.4]
  wire [10:0] buffer_0_182; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56647; // @[Modules.scala 50:57:@2640.4]
  wire [10:0] _T_56648; // @[Modules.scala 50:57:@2641.4]
  wire [10:0] buffer_0_483; // @[Modules.scala 50:57:@2642.4]
  wire [10:0] buffer_0_184; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56650; // @[Modules.scala 50:57:@2644.4]
  wire [10:0] _T_56651; // @[Modules.scala 50:57:@2645.4]
  wire [10:0] buffer_0_484; // @[Modules.scala 50:57:@2646.4]
  wire [10:0] buffer_0_186; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_187; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56653; // @[Modules.scala 50:57:@2648.4]
  wire [10:0] _T_56654; // @[Modules.scala 50:57:@2649.4]
  wire [10:0] buffer_0_485; // @[Modules.scala 50:57:@2650.4]
  wire [10:0] buffer_0_188; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56656; // @[Modules.scala 50:57:@2652.4]
  wire [10:0] _T_56657; // @[Modules.scala 50:57:@2653.4]
  wire [10:0] buffer_0_486; // @[Modules.scala 50:57:@2654.4]
  wire [10:0] buffer_0_190; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56659; // @[Modules.scala 50:57:@2656.4]
  wire [10:0] _T_56660; // @[Modules.scala 50:57:@2657.4]
  wire [10:0] buffer_0_487; // @[Modules.scala 50:57:@2658.4]
  wire [10:0] buffer_0_192; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_193; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56662; // @[Modules.scala 50:57:@2660.4]
  wire [10:0] _T_56663; // @[Modules.scala 50:57:@2661.4]
  wire [10:0] buffer_0_488; // @[Modules.scala 50:57:@2662.4]
  wire [10:0] buffer_0_194; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56665; // @[Modules.scala 50:57:@2664.4]
  wire [10:0] _T_56666; // @[Modules.scala 50:57:@2665.4]
  wire [10:0] buffer_0_489; // @[Modules.scala 50:57:@2666.4]
  wire [10:0] buffer_0_196; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56668; // @[Modules.scala 50:57:@2668.4]
  wire [10:0] _T_56669; // @[Modules.scala 50:57:@2669.4]
  wire [10:0] buffer_0_490; // @[Modules.scala 50:57:@2670.4]
  wire [10:0] buffer_0_198; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56671; // @[Modules.scala 50:57:@2672.4]
  wire [10:0] _T_56672; // @[Modules.scala 50:57:@2673.4]
  wire [10:0] buffer_0_491; // @[Modules.scala 50:57:@2674.4]
  wire [10:0] buffer_0_200; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_201; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56674; // @[Modules.scala 50:57:@2676.4]
  wire [10:0] _T_56675; // @[Modules.scala 50:57:@2677.4]
  wire [10:0] buffer_0_492; // @[Modules.scala 50:57:@2678.4]
  wire [10:0] buffer_0_202; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56677; // @[Modules.scala 50:57:@2680.4]
  wire [10:0] _T_56678; // @[Modules.scala 50:57:@2681.4]
  wire [10:0] buffer_0_493; // @[Modules.scala 50:57:@2682.4]
  wire [10:0] buffer_0_204; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56680; // @[Modules.scala 50:57:@2684.4]
  wire [10:0] _T_56681; // @[Modules.scala 50:57:@2685.4]
  wire [10:0] buffer_0_494; // @[Modules.scala 50:57:@2686.4]
  wire [10:0] buffer_0_206; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_207; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56683; // @[Modules.scala 50:57:@2688.4]
  wire [10:0] _T_56684; // @[Modules.scala 50:57:@2689.4]
  wire [10:0] buffer_0_495; // @[Modules.scala 50:57:@2690.4]
  wire [10:0] buffer_0_208; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56686; // @[Modules.scala 50:57:@2692.4]
  wire [10:0] _T_56687; // @[Modules.scala 50:57:@2693.4]
  wire [10:0] buffer_0_496; // @[Modules.scala 50:57:@2694.4]
  wire [10:0] buffer_0_210; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56689; // @[Modules.scala 50:57:@2696.4]
  wire [10:0] _T_56690; // @[Modules.scala 50:57:@2697.4]
  wire [10:0] buffer_0_497; // @[Modules.scala 50:57:@2698.4]
  wire [10:0] buffer_0_212; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56692; // @[Modules.scala 50:57:@2700.4]
  wire [10:0] _T_56693; // @[Modules.scala 50:57:@2701.4]
  wire [10:0] buffer_0_498; // @[Modules.scala 50:57:@2702.4]
  wire [10:0] buffer_0_214; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56695; // @[Modules.scala 50:57:@2704.4]
  wire [10:0] _T_56696; // @[Modules.scala 50:57:@2705.4]
  wire [10:0] buffer_0_499; // @[Modules.scala 50:57:@2706.4]
  wire [10:0] buffer_0_216; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56698; // @[Modules.scala 50:57:@2708.4]
  wire [10:0] _T_56699; // @[Modules.scala 50:57:@2709.4]
  wire [10:0] buffer_0_500; // @[Modules.scala 50:57:@2710.4]
  wire [10:0] buffer_0_218; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56701; // @[Modules.scala 50:57:@2712.4]
  wire [10:0] _T_56702; // @[Modules.scala 50:57:@2713.4]
  wire [10:0] buffer_0_501; // @[Modules.scala 50:57:@2714.4]
  wire [10:0] buffer_0_220; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56704; // @[Modules.scala 50:57:@2716.4]
  wire [10:0] _T_56705; // @[Modules.scala 50:57:@2717.4]
  wire [10:0] buffer_0_502; // @[Modules.scala 50:57:@2718.4]
  wire [10:0] buffer_0_222; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_223; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56707; // @[Modules.scala 50:57:@2720.4]
  wire [10:0] _T_56708; // @[Modules.scala 50:57:@2721.4]
  wire [10:0] buffer_0_503; // @[Modules.scala 50:57:@2722.4]
  wire [10:0] buffer_0_224; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56710; // @[Modules.scala 50:57:@2724.4]
  wire [10:0] _T_56711; // @[Modules.scala 50:57:@2725.4]
  wire [10:0] buffer_0_504; // @[Modules.scala 50:57:@2726.4]
  wire [10:0] buffer_0_226; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56713; // @[Modules.scala 50:57:@2728.4]
  wire [10:0] _T_56714; // @[Modules.scala 50:57:@2729.4]
  wire [10:0] buffer_0_505; // @[Modules.scala 50:57:@2730.4]
  wire [10:0] buffer_0_228; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56716; // @[Modules.scala 50:57:@2732.4]
  wire [10:0] _T_56717; // @[Modules.scala 50:57:@2733.4]
  wire [10:0] buffer_0_506; // @[Modules.scala 50:57:@2734.4]
  wire [10:0] buffer_0_230; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56719; // @[Modules.scala 50:57:@2736.4]
  wire [10:0] _T_56720; // @[Modules.scala 50:57:@2737.4]
  wire [10:0] buffer_0_507; // @[Modules.scala 50:57:@2738.4]
  wire [10:0] buffer_0_232; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56722; // @[Modules.scala 50:57:@2740.4]
  wire [10:0] _T_56723; // @[Modules.scala 50:57:@2741.4]
  wire [10:0] buffer_0_508; // @[Modules.scala 50:57:@2742.4]
  wire [10:0] buffer_0_234; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56725; // @[Modules.scala 50:57:@2744.4]
  wire [10:0] _T_56726; // @[Modules.scala 50:57:@2745.4]
  wire [10:0] buffer_0_509; // @[Modules.scala 50:57:@2746.4]
  wire [10:0] buffer_0_236; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_237; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56728; // @[Modules.scala 50:57:@2748.4]
  wire [10:0] _T_56729; // @[Modules.scala 50:57:@2749.4]
  wire [10:0] buffer_0_510; // @[Modules.scala 50:57:@2750.4]
  wire [10:0] buffer_0_238; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56731; // @[Modules.scala 50:57:@2752.4]
  wire [10:0] _T_56732; // @[Modules.scala 50:57:@2753.4]
  wire [10:0] buffer_0_511; // @[Modules.scala 50:57:@2754.4]
  wire [10:0] buffer_0_240; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56734; // @[Modules.scala 50:57:@2756.4]
  wire [10:0] _T_56735; // @[Modules.scala 50:57:@2757.4]
  wire [10:0] buffer_0_512; // @[Modules.scala 50:57:@2758.4]
  wire [10:0] buffer_0_242; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_243; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56737; // @[Modules.scala 50:57:@2760.4]
  wire [10:0] _T_56738; // @[Modules.scala 50:57:@2761.4]
  wire [10:0] buffer_0_513; // @[Modules.scala 50:57:@2762.4]
  wire [10:0] buffer_0_244; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56740; // @[Modules.scala 50:57:@2764.4]
  wire [10:0] _T_56741; // @[Modules.scala 50:57:@2765.4]
  wire [10:0] buffer_0_514; // @[Modules.scala 50:57:@2766.4]
  wire [10:0] buffer_0_246; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56743; // @[Modules.scala 50:57:@2768.4]
  wire [10:0] _T_56744; // @[Modules.scala 50:57:@2769.4]
  wire [10:0] buffer_0_515; // @[Modules.scala 50:57:@2770.4]
  wire [10:0] buffer_0_248; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56746; // @[Modules.scala 50:57:@2772.4]
  wire [10:0] _T_56747; // @[Modules.scala 50:57:@2773.4]
  wire [10:0] buffer_0_516; // @[Modules.scala 50:57:@2774.4]
  wire [10:0] buffer_0_250; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_251; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56749; // @[Modules.scala 50:57:@2776.4]
  wire [10:0] _T_56750; // @[Modules.scala 50:57:@2777.4]
  wire [10:0] buffer_0_517; // @[Modules.scala 50:57:@2778.4]
  wire [10:0] buffer_0_252; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56752; // @[Modules.scala 50:57:@2780.4]
  wire [10:0] _T_56753; // @[Modules.scala 50:57:@2781.4]
  wire [10:0] buffer_0_518; // @[Modules.scala 50:57:@2782.4]
  wire [10:0] buffer_0_254; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56755; // @[Modules.scala 50:57:@2784.4]
  wire [10:0] _T_56756; // @[Modules.scala 50:57:@2785.4]
  wire [10:0] buffer_0_519; // @[Modules.scala 50:57:@2786.4]
  wire [10:0] buffer_0_256; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_257; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56758; // @[Modules.scala 50:57:@2788.4]
  wire [10:0] _T_56759; // @[Modules.scala 50:57:@2789.4]
  wire [10:0] buffer_0_520; // @[Modules.scala 50:57:@2790.4]
  wire [10:0] buffer_0_258; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56761; // @[Modules.scala 50:57:@2792.4]
  wire [10:0] _T_56762; // @[Modules.scala 50:57:@2793.4]
  wire [10:0] buffer_0_521; // @[Modules.scala 50:57:@2794.4]
  wire [10:0] buffer_0_260; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_261; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56764; // @[Modules.scala 50:57:@2796.4]
  wire [10:0] _T_56765; // @[Modules.scala 50:57:@2797.4]
  wire [10:0] buffer_0_522; // @[Modules.scala 50:57:@2798.4]
  wire [10:0] buffer_0_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56767; // @[Modules.scala 50:57:@2800.4]
  wire [10:0] _T_56768; // @[Modules.scala 50:57:@2801.4]
  wire [10:0] buffer_0_523; // @[Modules.scala 50:57:@2802.4]
  wire [10:0] buffer_0_264; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_265; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56770; // @[Modules.scala 50:57:@2804.4]
  wire [10:0] _T_56771; // @[Modules.scala 50:57:@2805.4]
  wire [10:0] buffer_0_524; // @[Modules.scala 50:57:@2806.4]
  wire [10:0] buffer_0_266; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_267; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56773; // @[Modules.scala 50:57:@2808.4]
  wire [10:0] _T_56774; // @[Modules.scala 50:57:@2809.4]
  wire [10:0] buffer_0_525; // @[Modules.scala 50:57:@2810.4]
  wire [10:0] buffer_0_268; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56776; // @[Modules.scala 50:57:@2812.4]
  wire [10:0] _T_56777; // @[Modules.scala 50:57:@2813.4]
  wire [10:0] buffer_0_526; // @[Modules.scala 50:57:@2814.4]
  wire [10:0] buffer_0_270; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_271; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56779; // @[Modules.scala 50:57:@2816.4]
  wire [10:0] _T_56780; // @[Modules.scala 50:57:@2817.4]
  wire [10:0] buffer_0_527; // @[Modules.scala 50:57:@2818.4]
  wire [10:0] buffer_0_272; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56782; // @[Modules.scala 50:57:@2820.4]
  wire [10:0] _T_56783; // @[Modules.scala 50:57:@2821.4]
  wire [10:0] buffer_0_528; // @[Modules.scala 50:57:@2822.4]
  wire [10:0] buffer_0_274; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56785; // @[Modules.scala 50:57:@2824.4]
  wire [10:0] _T_56786; // @[Modules.scala 50:57:@2825.4]
  wire [10:0] buffer_0_529; // @[Modules.scala 50:57:@2826.4]
  wire [10:0] buffer_0_276; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56788; // @[Modules.scala 50:57:@2828.4]
  wire [10:0] _T_56789; // @[Modules.scala 50:57:@2829.4]
  wire [10:0] buffer_0_530; // @[Modules.scala 50:57:@2830.4]
  wire [10:0] buffer_0_278; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56791; // @[Modules.scala 50:57:@2832.4]
  wire [10:0] _T_56792; // @[Modules.scala 50:57:@2833.4]
  wire [10:0] buffer_0_531; // @[Modules.scala 50:57:@2834.4]
  wire [10:0] buffer_0_280; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56794; // @[Modules.scala 50:57:@2836.4]
  wire [10:0] _T_56795; // @[Modules.scala 50:57:@2837.4]
  wire [10:0] buffer_0_532; // @[Modules.scala 50:57:@2838.4]
  wire [10:0] buffer_0_282; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56797; // @[Modules.scala 50:57:@2840.4]
  wire [10:0] _T_56798; // @[Modules.scala 50:57:@2841.4]
  wire [10:0] buffer_0_533; // @[Modules.scala 50:57:@2842.4]
  wire [10:0] buffer_0_284; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_285; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56800; // @[Modules.scala 50:57:@2844.4]
  wire [10:0] _T_56801; // @[Modules.scala 50:57:@2845.4]
  wire [10:0] buffer_0_534; // @[Modules.scala 50:57:@2846.4]
  wire [10:0] buffer_0_286; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56803; // @[Modules.scala 50:57:@2848.4]
  wire [10:0] _T_56804; // @[Modules.scala 50:57:@2849.4]
  wire [10:0] buffer_0_535; // @[Modules.scala 50:57:@2850.4]
  wire [10:0] buffer_0_288; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56806; // @[Modules.scala 50:57:@2852.4]
  wire [10:0] _T_56807; // @[Modules.scala 50:57:@2853.4]
  wire [10:0] buffer_0_536; // @[Modules.scala 50:57:@2854.4]
  wire [10:0] buffer_0_290; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56809; // @[Modules.scala 50:57:@2856.4]
  wire [10:0] _T_56810; // @[Modules.scala 50:57:@2857.4]
  wire [10:0] buffer_0_537; // @[Modules.scala 50:57:@2858.4]
  wire [10:0] buffer_0_292; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56812; // @[Modules.scala 50:57:@2860.4]
  wire [10:0] _T_56813; // @[Modules.scala 50:57:@2861.4]
  wire [10:0] buffer_0_538; // @[Modules.scala 50:57:@2862.4]
  wire [10:0] buffer_0_294; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_295; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56815; // @[Modules.scala 50:57:@2864.4]
  wire [10:0] _T_56816; // @[Modules.scala 50:57:@2865.4]
  wire [10:0] buffer_0_539; // @[Modules.scala 50:57:@2866.4]
  wire [10:0] buffer_0_296; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56818; // @[Modules.scala 50:57:@2868.4]
  wire [10:0] _T_56819; // @[Modules.scala 50:57:@2869.4]
  wire [10:0] buffer_0_540; // @[Modules.scala 50:57:@2870.4]
  wire [10:0] buffer_0_298; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56821; // @[Modules.scala 50:57:@2872.4]
  wire [10:0] _T_56822; // @[Modules.scala 50:57:@2873.4]
  wire [10:0] buffer_0_541; // @[Modules.scala 50:57:@2874.4]
  wire [10:0] buffer_0_300; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56824; // @[Modules.scala 50:57:@2876.4]
  wire [10:0] _T_56825; // @[Modules.scala 50:57:@2877.4]
  wire [10:0] buffer_0_542; // @[Modules.scala 50:57:@2878.4]
  wire [10:0] buffer_0_302; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_303; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56827; // @[Modules.scala 50:57:@2880.4]
  wire [10:0] _T_56828; // @[Modules.scala 50:57:@2881.4]
  wire [10:0] buffer_0_543; // @[Modules.scala 50:57:@2882.4]
  wire [10:0] buffer_0_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56830; // @[Modules.scala 50:57:@2884.4]
  wire [10:0] _T_56831; // @[Modules.scala 50:57:@2885.4]
  wire [10:0] buffer_0_544; // @[Modules.scala 50:57:@2886.4]
  wire [10:0] buffer_0_306; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56833; // @[Modules.scala 50:57:@2888.4]
  wire [10:0] _T_56834; // @[Modules.scala 50:57:@2889.4]
  wire [10:0] buffer_0_545; // @[Modules.scala 50:57:@2890.4]
  wire [10:0] buffer_0_308; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56836; // @[Modules.scala 50:57:@2892.4]
  wire [10:0] _T_56837; // @[Modules.scala 50:57:@2893.4]
  wire [10:0] buffer_0_546; // @[Modules.scala 50:57:@2894.4]
  wire [10:0] buffer_0_310; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56839; // @[Modules.scala 50:57:@2896.4]
  wire [10:0] _T_56840; // @[Modules.scala 50:57:@2897.4]
  wire [10:0] buffer_0_547; // @[Modules.scala 50:57:@2898.4]
  wire [10:0] buffer_0_312; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56842; // @[Modules.scala 50:57:@2900.4]
  wire [10:0] _T_56843; // @[Modules.scala 50:57:@2901.4]
  wire [10:0] buffer_0_548; // @[Modules.scala 50:57:@2902.4]
  wire [10:0] buffer_0_314; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56845; // @[Modules.scala 50:57:@2904.4]
  wire [10:0] _T_56846; // @[Modules.scala 50:57:@2905.4]
  wire [10:0] buffer_0_549; // @[Modules.scala 50:57:@2906.4]
  wire [10:0] buffer_0_316; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56848; // @[Modules.scala 50:57:@2908.4]
  wire [10:0] _T_56849; // @[Modules.scala 50:57:@2909.4]
  wire [10:0] buffer_0_550; // @[Modules.scala 50:57:@2910.4]
  wire [10:0] buffer_0_318; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56851; // @[Modules.scala 50:57:@2912.4]
  wire [10:0] _T_56852; // @[Modules.scala 50:57:@2913.4]
  wire [10:0] buffer_0_551; // @[Modules.scala 50:57:@2914.4]
  wire [10:0] buffer_0_320; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56854; // @[Modules.scala 50:57:@2916.4]
  wire [10:0] _T_56855; // @[Modules.scala 50:57:@2917.4]
  wire [10:0] buffer_0_552; // @[Modules.scala 50:57:@2918.4]
  wire [10:0] buffer_0_322; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_323; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56857; // @[Modules.scala 50:57:@2920.4]
  wire [10:0] _T_56858; // @[Modules.scala 50:57:@2921.4]
  wire [10:0] buffer_0_553; // @[Modules.scala 50:57:@2922.4]
  wire [10:0] buffer_0_324; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56860; // @[Modules.scala 50:57:@2924.4]
  wire [10:0] _T_56861; // @[Modules.scala 50:57:@2925.4]
  wire [10:0] buffer_0_554; // @[Modules.scala 50:57:@2926.4]
  wire [10:0] buffer_0_326; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56863; // @[Modules.scala 50:57:@2928.4]
  wire [10:0] _T_56864; // @[Modules.scala 50:57:@2929.4]
  wire [10:0] buffer_0_555; // @[Modules.scala 50:57:@2930.4]
  wire [10:0] buffer_0_328; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56866; // @[Modules.scala 50:57:@2932.4]
  wire [10:0] _T_56867; // @[Modules.scala 50:57:@2933.4]
  wire [10:0] buffer_0_556; // @[Modules.scala 50:57:@2934.4]
  wire [10:0] buffer_0_330; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_331; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56869; // @[Modules.scala 50:57:@2936.4]
  wire [10:0] _T_56870; // @[Modules.scala 50:57:@2937.4]
  wire [10:0] buffer_0_557; // @[Modules.scala 50:57:@2938.4]
  wire [10:0] buffer_0_332; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_333; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56872; // @[Modules.scala 50:57:@2940.4]
  wire [10:0] _T_56873; // @[Modules.scala 50:57:@2941.4]
  wire [10:0] buffer_0_558; // @[Modules.scala 50:57:@2942.4]
  wire [10:0] buffer_0_334; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56875; // @[Modules.scala 50:57:@2944.4]
  wire [10:0] _T_56876; // @[Modules.scala 50:57:@2945.4]
  wire [10:0] buffer_0_559; // @[Modules.scala 50:57:@2946.4]
  wire [10:0] buffer_0_336; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56878; // @[Modules.scala 50:57:@2948.4]
  wire [10:0] _T_56879; // @[Modules.scala 50:57:@2949.4]
  wire [10:0] buffer_0_560; // @[Modules.scala 50:57:@2950.4]
  wire [10:0] buffer_0_338; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56881; // @[Modules.scala 50:57:@2952.4]
  wire [10:0] _T_56882; // @[Modules.scala 50:57:@2953.4]
  wire [10:0] buffer_0_561; // @[Modules.scala 50:57:@2954.4]
  wire [10:0] buffer_0_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56884; // @[Modules.scala 50:57:@2956.4]
  wire [10:0] _T_56885; // @[Modules.scala 50:57:@2957.4]
  wire [10:0] buffer_0_562; // @[Modules.scala 50:57:@2958.4]
  wire [10:0] buffer_0_342; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56887; // @[Modules.scala 50:57:@2960.4]
  wire [10:0] _T_56888; // @[Modules.scala 50:57:@2961.4]
  wire [10:0] buffer_0_563; // @[Modules.scala 50:57:@2962.4]
  wire [10:0] buffer_0_344; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56890; // @[Modules.scala 50:57:@2964.4]
  wire [10:0] _T_56891; // @[Modules.scala 50:57:@2965.4]
  wire [10:0] buffer_0_564; // @[Modules.scala 50:57:@2966.4]
  wire [10:0] buffer_0_346; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56893; // @[Modules.scala 50:57:@2968.4]
  wire [10:0] _T_56894; // @[Modules.scala 50:57:@2969.4]
  wire [10:0] buffer_0_565; // @[Modules.scala 50:57:@2970.4]
  wire [10:0] buffer_0_348; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56896; // @[Modules.scala 50:57:@2972.4]
  wire [10:0] _T_56897; // @[Modules.scala 50:57:@2973.4]
  wire [10:0] buffer_0_566; // @[Modules.scala 50:57:@2974.4]
  wire [10:0] buffer_0_350; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56899; // @[Modules.scala 50:57:@2976.4]
  wire [10:0] _T_56900; // @[Modules.scala 50:57:@2977.4]
  wire [10:0] buffer_0_567; // @[Modules.scala 50:57:@2978.4]
  wire [10:0] buffer_0_352; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_353; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56902; // @[Modules.scala 50:57:@2980.4]
  wire [10:0] _T_56903; // @[Modules.scala 50:57:@2981.4]
  wire [10:0] buffer_0_568; // @[Modules.scala 50:57:@2982.4]
  wire [10:0] buffer_0_354; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56905; // @[Modules.scala 50:57:@2984.4]
  wire [10:0] _T_56906; // @[Modules.scala 50:57:@2985.4]
  wire [10:0] buffer_0_569; // @[Modules.scala 50:57:@2986.4]
  wire [10:0] buffer_0_356; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56908; // @[Modules.scala 50:57:@2988.4]
  wire [10:0] _T_56909; // @[Modules.scala 50:57:@2989.4]
  wire [10:0] buffer_0_570; // @[Modules.scala 50:57:@2990.4]
  wire [10:0] buffer_0_358; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_359; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56911; // @[Modules.scala 50:57:@2992.4]
  wire [10:0] _T_56912; // @[Modules.scala 50:57:@2993.4]
  wire [10:0] buffer_0_571; // @[Modules.scala 50:57:@2994.4]
  wire [10:0] buffer_0_360; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56914; // @[Modules.scala 50:57:@2996.4]
  wire [10:0] _T_56915; // @[Modules.scala 50:57:@2997.4]
  wire [10:0] buffer_0_572; // @[Modules.scala 50:57:@2998.4]
  wire [10:0] buffer_0_362; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56917; // @[Modules.scala 50:57:@3000.4]
  wire [10:0] _T_56918; // @[Modules.scala 50:57:@3001.4]
  wire [10:0] buffer_0_573; // @[Modules.scala 50:57:@3002.4]
  wire [10:0] buffer_0_364; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56920; // @[Modules.scala 50:57:@3004.4]
  wire [10:0] _T_56921; // @[Modules.scala 50:57:@3005.4]
  wire [10:0] buffer_0_574; // @[Modules.scala 50:57:@3006.4]
  wire [10:0] buffer_0_366; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56923; // @[Modules.scala 50:57:@3008.4]
  wire [10:0] _T_56924; // @[Modules.scala 50:57:@3009.4]
  wire [10:0] buffer_0_575; // @[Modules.scala 50:57:@3010.4]
  wire [10:0] buffer_0_368; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_369; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56926; // @[Modules.scala 50:57:@3012.4]
  wire [10:0] _T_56927; // @[Modules.scala 50:57:@3013.4]
  wire [10:0] buffer_0_576; // @[Modules.scala 50:57:@3014.4]
  wire [10:0] buffer_0_370; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56929; // @[Modules.scala 50:57:@3016.4]
  wire [10:0] _T_56930; // @[Modules.scala 50:57:@3017.4]
  wire [10:0] buffer_0_577; // @[Modules.scala 50:57:@3018.4]
  wire [10:0] buffer_0_372; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_373; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56932; // @[Modules.scala 50:57:@3020.4]
  wire [10:0] _T_56933; // @[Modules.scala 50:57:@3021.4]
  wire [10:0] buffer_0_578; // @[Modules.scala 50:57:@3022.4]
  wire [10:0] buffer_0_374; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56935; // @[Modules.scala 50:57:@3024.4]
  wire [10:0] _T_56936; // @[Modules.scala 50:57:@3025.4]
  wire [10:0] buffer_0_579; // @[Modules.scala 50:57:@3026.4]
  wire [10:0] buffer_0_376; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56938; // @[Modules.scala 50:57:@3028.4]
  wire [10:0] _T_56939; // @[Modules.scala 50:57:@3029.4]
  wire [10:0] buffer_0_580; // @[Modules.scala 50:57:@3030.4]
  wire [10:0] buffer_0_378; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56941; // @[Modules.scala 50:57:@3032.4]
  wire [10:0] _T_56942; // @[Modules.scala 50:57:@3033.4]
  wire [10:0] buffer_0_581; // @[Modules.scala 50:57:@3034.4]
  wire [10:0] buffer_0_380; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_381; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56944; // @[Modules.scala 50:57:@3036.4]
  wire [10:0] _T_56945; // @[Modules.scala 50:57:@3037.4]
  wire [10:0] buffer_0_582; // @[Modules.scala 50:57:@3038.4]
  wire [10:0] buffer_0_382; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56947; // @[Modules.scala 50:57:@3040.4]
  wire [10:0] _T_56948; // @[Modules.scala 50:57:@3041.4]
  wire [10:0] buffer_0_583; // @[Modules.scala 50:57:@3042.4]
  wire [10:0] buffer_0_384; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_385; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56950; // @[Modules.scala 50:57:@3044.4]
  wire [10:0] _T_56951; // @[Modules.scala 50:57:@3045.4]
  wire [10:0] buffer_0_584; // @[Modules.scala 50:57:@3046.4]
  wire [10:0] buffer_0_386; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_387; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56953; // @[Modules.scala 50:57:@3048.4]
  wire [10:0] _T_56954; // @[Modules.scala 50:57:@3049.4]
  wire [10:0] buffer_0_585; // @[Modules.scala 50:57:@3050.4]
  wire [10:0] buffer_0_388; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56956; // @[Modules.scala 50:57:@3052.4]
  wire [10:0] _T_56957; // @[Modules.scala 50:57:@3053.4]
  wire [10:0] buffer_0_586; // @[Modules.scala 50:57:@3054.4]
  wire [10:0] buffer_0_390; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56959; // @[Modules.scala 50:57:@3056.4]
  wire [10:0] _T_56960; // @[Modules.scala 50:57:@3057.4]
  wire [10:0] buffer_0_587; // @[Modules.scala 50:57:@3058.4]
  wire [11:0] _T_56962; // @[Modules.scala 53:83:@3060.4]
  wire [10:0] _T_56963; // @[Modules.scala 53:83:@3061.4]
  wire [10:0] buffer_0_588; // @[Modules.scala 53:83:@3062.4]
  wire [11:0] _T_56965; // @[Modules.scala 53:83:@3064.4]
  wire [10:0] _T_56966; // @[Modules.scala 53:83:@3065.4]
  wire [10:0] buffer_0_589; // @[Modules.scala 53:83:@3066.4]
  wire [11:0] _T_56968; // @[Modules.scala 53:83:@3068.4]
  wire [10:0] _T_56969; // @[Modules.scala 53:83:@3069.4]
  wire [10:0] buffer_0_590; // @[Modules.scala 53:83:@3070.4]
  wire [11:0] _T_56971; // @[Modules.scala 53:83:@3072.4]
  wire [10:0] _T_56972; // @[Modules.scala 53:83:@3073.4]
  wire [10:0] buffer_0_591; // @[Modules.scala 53:83:@3074.4]
  wire [11:0] _T_56974; // @[Modules.scala 53:83:@3076.4]
  wire [10:0] _T_56975; // @[Modules.scala 53:83:@3077.4]
  wire [10:0] buffer_0_592; // @[Modules.scala 53:83:@3078.4]
  wire [11:0] _T_56977; // @[Modules.scala 53:83:@3080.4]
  wire [10:0] _T_56978; // @[Modules.scala 53:83:@3081.4]
  wire [10:0] buffer_0_593; // @[Modules.scala 53:83:@3082.4]
  wire [11:0] _T_56980; // @[Modules.scala 53:83:@3084.4]
  wire [10:0] _T_56981; // @[Modules.scala 53:83:@3085.4]
  wire [10:0] buffer_0_594; // @[Modules.scala 53:83:@3086.4]
  wire [11:0] _T_56983; // @[Modules.scala 53:83:@3088.4]
  wire [10:0] _T_56984; // @[Modules.scala 53:83:@3089.4]
  wire [10:0] buffer_0_595; // @[Modules.scala 53:83:@3090.4]
  wire [11:0] _T_56986; // @[Modules.scala 53:83:@3092.4]
  wire [10:0] _T_56987; // @[Modules.scala 53:83:@3093.4]
  wire [10:0] buffer_0_596; // @[Modules.scala 53:83:@3094.4]
  wire [11:0] _T_56989; // @[Modules.scala 53:83:@3096.4]
  wire [10:0] _T_56990; // @[Modules.scala 53:83:@3097.4]
  wire [10:0] buffer_0_597; // @[Modules.scala 53:83:@3098.4]
  wire [11:0] _T_56992; // @[Modules.scala 53:83:@3100.4]
  wire [10:0] _T_56993; // @[Modules.scala 53:83:@3101.4]
  wire [10:0] buffer_0_598; // @[Modules.scala 53:83:@3102.4]
  wire [11:0] _T_56995; // @[Modules.scala 53:83:@3104.4]
  wire [10:0] _T_56996; // @[Modules.scala 53:83:@3105.4]
  wire [10:0] buffer_0_599; // @[Modules.scala 53:83:@3106.4]
  wire [11:0] _T_56998; // @[Modules.scala 53:83:@3108.4]
  wire [10:0] _T_56999; // @[Modules.scala 53:83:@3109.4]
  wire [10:0] buffer_0_600; // @[Modules.scala 53:83:@3110.4]
  wire [11:0] _T_57001; // @[Modules.scala 53:83:@3112.4]
  wire [10:0] _T_57002; // @[Modules.scala 53:83:@3113.4]
  wire [10:0] buffer_0_601; // @[Modules.scala 53:83:@3114.4]
  wire [11:0] _T_57004; // @[Modules.scala 53:83:@3116.4]
  wire [10:0] _T_57005; // @[Modules.scala 53:83:@3117.4]
  wire [10:0] buffer_0_602; // @[Modules.scala 53:83:@3118.4]
  wire [11:0] _T_57007; // @[Modules.scala 53:83:@3120.4]
  wire [10:0] _T_57008; // @[Modules.scala 53:83:@3121.4]
  wire [10:0] buffer_0_603; // @[Modules.scala 53:83:@3122.4]
  wire [11:0] _T_57010; // @[Modules.scala 53:83:@3124.4]
  wire [10:0] _T_57011; // @[Modules.scala 53:83:@3125.4]
  wire [10:0] buffer_0_604; // @[Modules.scala 53:83:@3126.4]
  wire [11:0] _T_57013; // @[Modules.scala 53:83:@3128.4]
  wire [10:0] _T_57014; // @[Modules.scala 53:83:@3129.4]
  wire [10:0] buffer_0_605; // @[Modules.scala 53:83:@3130.4]
  wire [11:0] _T_57016; // @[Modules.scala 53:83:@3132.4]
  wire [10:0] _T_57017; // @[Modules.scala 53:83:@3133.4]
  wire [10:0] buffer_0_606; // @[Modules.scala 53:83:@3134.4]
  wire [11:0] _T_57019; // @[Modules.scala 53:83:@3136.4]
  wire [10:0] _T_57020; // @[Modules.scala 53:83:@3137.4]
  wire [10:0] buffer_0_607; // @[Modules.scala 53:83:@3138.4]
  wire [11:0] _T_57022; // @[Modules.scala 53:83:@3140.4]
  wire [10:0] _T_57023; // @[Modules.scala 53:83:@3141.4]
  wire [10:0] buffer_0_608; // @[Modules.scala 53:83:@3142.4]
  wire [11:0] _T_57025; // @[Modules.scala 53:83:@3144.4]
  wire [10:0] _T_57026; // @[Modules.scala 53:83:@3145.4]
  wire [10:0] buffer_0_609; // @[Modules.scala 53:83:@3146.4]
  wire [11:0] _T_57028; // @[Modules.scala 53:83:@3148.4]
  wire [10:0] _T_57029; // @[Modules.scala 53:83:@3149.4]
  wire [10:0] buffer_0_610; // @[Modules.scala 53:83:@3150.4]
  wire [11:0] _T_57031; // @[Modules.scala 53:83:@3152.4]
  wire [10:0] _T_57032; // @[Modules.scala 53:83:@3153.4]
  wire [10:0] buffer_0_611; // @[Modules.scala 53:83:@3154.4]
  wire [11:0] _T_57034; // @[Modules.scala 53:83:@3156.4]
  wire [10:0] _T_57035; // @[Modules.scala 53:83:@3157.4]
  wire [10:0] buffer_0_612; // @[Modules.scala 53:83:@3158.4]
  wire [11:0] _T_57037; // @[Modules.scala 53:83:@3160.4]
  wire [10:0] _T_57038; // @[Modules.scala 53:83:@3161.4]
  wire [10:0] buffer_0_613; // @[Modules.scala 53:83:@3162.4]
  wire [11:0] _T_57040; // @[Modules.scala 53:83:@3164.4]
  wire [10:0] _T_57041; // @[Modules.scala 53:83:@3165.4]
  wire [10:0] buffer_0_614; // @[Modules.scala 53:83:@3166.4]
  wire [11:0] _T_57043; // @[Modules.scala 53:83:@3168.4]
  wire [10:0] _T_57044; // @[Modules.scala 53:83:@3169.4]
  wire [10:0] buffer_0_615; // @[Modules.scala 53:83:@3170.4]
  wire [11:0] _T_57046; // @[Modules.scala 53:83:@3172.4]
  wire [10:0] _T_57047; // @[Modules.scala 53:83:@3173.4]
  wire [10:0] buffer_0_616; // @[Modules.scala 53:83:@3174.4]
  wire [11:0] _T_57049; // @[Modules.scala 53:83:@3176.4]
  wire [10:0] _T_57050; // @[Modules.scala 53:83:@3177.4]
  wire [10:0] buffer_0_617; // @[Modules.scala 53:83:@3178.4]
  wire [11:0] _T_57052; // @[Modules.scala 53:83:@3180.4]
  wire [10:0] _T_57053; // @[Modules.scala 53:83:@3181.4]
  wire [10:0] buffer_0_618; // @[Modules.scala 53:83:@3182.4]
  wire [11:0] _T_57055; // @[Modules.scala 53:83:@3184.4]
  wire [10:0] _T_57056; // @[Modules.scala 53:83:@3185.4]
  wire [10:0] buffer_0_619; // @[Modules.scala 53:83:@3186.4]
  wire [11:0] _T_57058; // @[Modules.scala 53:83:@3188.4]
  wire [10:0] _T_57059; // @[Modules.scala 53:83:@3189.4]
  wire [10:0] buffer_0_620; // @[Modules.scala 53:83:@3190.4]
  wire [11:0] _T_57061; // @[Modules.scala 53:83:@3192.4]
  wire [10:0] _T_57062; // @[Modules.scala 53:83:@3193.4]
  wire [10:0] buffer_0_621; // @[Modules.scala 53:83:@3194.4]
  wire [11:0] _T_57064; // @[Modules.scala 53:83:@3196.4]
  wire [10:0] _T_57065; // @[Modules.scala 53:83:@3197.4]
  wire [10:0] buffer_0_622; // @[Modules.scala 53:83:@3198.4]
  wire [11:0] _T_57067; // @[Modules.scala 53:83:@3200.4]
  wire [10:0] _T_57068; // @[Modules.scala 53:83:@3201.4]
  wire [10:0] buffer_0_623; // @[Modules.scala 53:83:@3202.4]
  wire [11:0] _T_57070; // @[Modules.scala 53:83:@3204.4]
  wire [10:0] _T_57071; // @[Modules.scala 53:83:@3205.4]
  wire [10:0] buffer_0_624; // @[Modules.scala 53:83:@3206.4]
  wire [11:0] _T_57073; // @[Modules.scala 53:83:@3208.4]
  wire [10:0] _T_57074; // @[Modules.scala 53:83:@3209.4]
  wire [10:0] buffer_0_625; // @[Modules.scala 53:83:@3210.4]
  wire [11:0] _T_57076; // @[Modules.scala 53:83:@3212.4]
  wire [10:0] _T_57077; // @[Modules.scala 53:83:@3213.4]
  wire [10:0] buffer_0_626; // @[Modules.scala 53:83:@3214.4]
  wire [11:0] _T_57079; // @[Modules.scala 53:83:@3216.4]
  wire [10:0] _T_57080; // @[Modules.scala 53:83:@3217.4]
  wire [10:0] buffer_0_627; // @[Modules.scala 53:83:@3218.4]
  wire [11:0] _T_57082; // @[Modules.scala 53:83:@3220.4]
  wire [10:0] _T_57083; // @[Modules.scala 53:83:@3221.4]
  wire [10:0] buffer_0_628; // @[Modules.scala 53:83:@3222.4]
  wire [11:0] _T_57085; // @[Modules.scala 53:83:@3224.4]
  wire [10:0] _T_57086; // @[Modules.scala 53:83:@3225.4]
  wire [10:0] buffer_0_629; // @[Modules.scala 53:83:@3226.4]
  wire [11:0] _T_57088; // @[Modules.scala 53:83:@3228.4]
  wire [10:0] _T_57089; // @[Modules.scala 53:83:@3229.4]
  wire [10:0] buffer_0_630; // @[Modules.scala 53:83:@3230.4]
  wire [11:0] _T_57091; // @[Modules.scala 53:83:@3232.4]
  wire [10:0] _T_57092; // @[Modules.scala 53:83:@3233.4]
  wire [10:0] buffer_0_631; // @[Modules.scala 53:83:@3234.4]
  wire [11:0] _T_57094; // @[Modules.scala 53:83:@3236.4]
  wire [10:0] _T_57095; // @[Modules.scala 53:83:@3237.4]
  wire [10:0] buffer_0_632; // @[Modules.scala 53:83:@3238.4]
  wire [11:0] _T_57097; // @[Modules.scala 53:83:@3240.4]
  wire [10:0] _T_57098; // @[Modules.scala 53:83:@3241.4]
  wire [10:0] buffer_0_633; // @[Modules.scala 53:83:@3242.4]
  wire [11:0] _T_57100; // @[Modules.scala 53:83:@3244.4]
  wire [10:0] _T_57101; // @[Modules.scala 53:83:@3245.4]
  wire [10:0] buffer_0_634; // @[Modules.scala 53:83:@3246.4]
  wire [11:0] _T_57103; // @[Modules.scala 53:83:@3248.4]
  wire [10:0] _T_57104; // @[Modules.scala 53:83:@3249.4]
  wire [10:0] buffer_0_635; // @[Modules.scala 53:83:@3250.4]
  wire [11:0] _T_57106; // @[Modules.scala 53:83:@3252.4]
  wire [10:0] _T_57107; // @[Modules.scala 53:83:@3253.4]
  wire [10:0] buffer_0_636; // @[Modules.scala 53:83:@3254.4]
  wire [11:0] _T_57109; // @[Modules.scala 53:83:@3256.4]
  wire [10:0] _T_57110; // @[Modules.scala 53:83:@3257.4]
  wire [10:0] buffer_0_637; // @[Modules.scala 53:83:@3258.4]
  wire [11:0] _T_57112; // @[Modules.scala 53:83:@3260.4]
  wire [10:0] _T_57113; // @[Modules.scala 53:83:@3261.4]
  wire [10:0] buffer_0_638; // @[Modules.scala 53:83:@3262.4]
  wire [11:0] _T_57115; // @[Modules.scala 53:83:@3264.4]
  wire [10:0] _T_57116; // @[Modules.scala 53:83:@3265.4]
  wire [10:0] buffer_0_639; // @[Modules.scala 53:83:@3266.4]
  wire [11:0] _T_57118; // @[Modules.scala 53:83:@3268.4]
  wire [10:0] _T_57119; // @[Modules.scala 53:83:@3269.4]
  wire [10:0] buffer_0_640; // @[Modules.scala 53:83:@3270.4]
  wire [11:0] _T_57121; // @[Modules.scala 53:83:@3272.4]
  wire [10:0] _T_57122; // @[Modules.scala 53:83:@3273.4]
  wire [10:0] buffer_0_641; // @[Modules.scala 53:83:@3274.4]
  wire [11:0] _T_57124; // @[Modules.scala 53:83:@3276.4]
  wire [10:0] _T_57125; // @[Modules.scala 53:83:@3277.4]
  wire [10:0] buffer_0_642; // @[Modules.scala 53:83:@3278.4]
  wire [11:0] _T_57127; // @[Modules.scala 53:83:@3280.4]
  wire [10:0] _T_57128; // @[Modules.scala 53:83:@3281.4]
  wire [10:0] buffer_0_643; // @[Modules.scala 53:83:@3282.4]
  wire [11:0] _T_57130; // @[Modules.scala 53:83:@3284.4]
  wire [10:0] _T_57131; // @[Modules.scala 53:83:@3285.4]
  wire [10:0] buffer_0_644; // @[Modules.scala 53:83:@3286.4]
  wire [11:0] _T_57133; // @[Modules.scala 53:83:@3288.4]
  wire [10:0] _T_57134; // @[Modules.scala 53:83:@3289.4]
  wire [10:0] buffer_0_645; // @[Modules.scala 53:83:@3290.4]
  wire [11:0] _T_57136; // @[Modules.scala 53:83:@3292.4]
  wire [10:0] _T_57137; // @[Modules.scala 53:83:@3293.4]
  wire [10:0] buffer_0_646; // @[Modules.scala 53:83:@3294.4]
  wire [11:0] _T_57139; // @[Modules.scala 53:83:@3296.4]
  wire [10:0] _T_57140; // @[Modules.scala 53:83:@3297.4]
  wire [10:0] buffer_0_647; // @[Modules.scala 53:83:@3298.4]
  wire [11:0] _T_57142; // @[Modules.scala 53:83:@3300.4]
  wire [10:0] _T_57143; // @[Modules.scala 53:83:@3301.4]
  wire [10:0] buffer_0_648; // @[Modules.scala 53:83:@3302.4]
  wire [11:0] _T_57145; // @[Modules.scala 53:83:@3304.4]
  wire [10:0] _T_57146; // @[Modules.scala 53:83:@3305.4]
  wire [10:0] buffer_0_649; // @[Modules.scala 53:83:@3306.4]
  wire [11:0] _T_57148; // @[Modules.scala 53:83:@3308.4]
  wire [10:0] _T_57149; // @[Modules.scala 53:83:@3309.4]
  wire [10:0] buffer_0_650; // @[Modules.scala 53:83:@3310.4]
  wire [11:0] _T_57151; // @[Modules.scala 53:83:@3312.4]
  wire [10:0] _T_57152; // @[Modules.scala 53:83:@3313.4]
  wire [10:0] buffer_0_651; // @[Modules.scala 53:83:@3314.4]
  wire [11:0] _T_57154; // @[Modules.scala 53:83:@3316.4]
  wire [10:0] _T_57155; // @[Modules.scala 53:83:@3317.4]
  wire [10:0] buffer_0_652; // @[Modules.scala 53:83:@3318.4]
  wire [11:0] _T_57157; // @[Modules.scala 53:83:@3320.4]
  wire [10:0] _T_57158; // @[Modules.scala 53:83:@3321.4]
  wire [10:0] buffer_0_653; // @[Modules.scala 53:83:@3322.4]
  wire [11:0] _T_57160; // @[Modules.scala 53:83:@3324.4]
  wire [10:0] _T_57161; // @[Modules.scala 53:83:@3325.4]
  wire [10:0] buffer_0_654; // @[Modules.scala 53:83:@3326.4]
  wire [11:0] _T_57163; // @[Modules.scala 53:83:@3328.4]
  wire [10:0] _T_57164; // @[Modules.scala 53:83:@3329.4]
  wire [10:0] buffer_0_655; // @[Modules.scala 53:83:@3330.4]
  wire [11:0] _T_57166; // @[Modules.scala 53:83:@3332.4]
  wire [10:0] _T_57167; // @[Modules.scala 53:83:@3333.4]
  wire [10:0] buffer_0_656; // @[Modules.scala 53:83:@3334.4]
  wire [11:0] _T_57169; // @[Modules.scala 53:83:@3336.4]
  wire [10:0] _T_57170; // @[Modules.scala 53:83:@3337.4]
  wire [10:0] buffer_0_657; // @[Modules.scala 53:83:@3338.4]
  wire [11:0] _T_57172; // @[Modules.scala 53:83:@3340.4]
  wire [10:0] _T_57173; // @[Modules.scala 53:83:@3341.4]
  wire [10:0] buffer_0_658; // @[Modules.scala 53:83:@3342.4]
  wire [11:0] _T_57175; // @[Modules.scala 53:83:@3344.4]
  wire [10:0] _T_57176; // @[Modules.scala 53:83:@3345.4]
  wire [10:0] buffer_0_659; // @[Modules.scala 53:83:@3346.4]
  wire [11:0] _T_57178; // @[Modules.scala 53:83:@3348.4]
  wire [10:0] _T_57179; // @[Modules.scala 53:83:@3349.4]
  wire [10:0] buffer_0_660; // @[Modules.scala 53:83:@3350.4]
  wire [11:0] _T_57181; // @[Modules.scala 53:83:@3352.4]
  wire [10:0] _T_57182; // @[Modules.scala 53:83:@3353.4]
  wire [10:0] buffer_0_661; // @[Modules.scala 53:83:@3354.4]
  wire [11:0] _T_57184; // @[Modules.scala 53:83:@3356.4]
  wire [10:0] _T_57185; // @[Modules.scala 53:83:@3357.4]
  wire [10:0] buffer_0_662; // @[Modules.scala 53:83:@3358.4]
  wire [11:0] _T_57187; // @[Modules.scala 53:83:@3360.4]
  wire [10:0] _T_57188; // @[Modules.scala 53:83:@3361.4]
  wire [10:0] buffer_0_663; // @[Modules.scala 53:83:@3362.4]
  wire [11:0] _T_57190; // @[Modules.scala 53:83:@3364.4]
  wire [10:0] _T_57191; // @[Modules.scala 53:83:@3365.4]
  wire [10:0] buffer_0_664; // @[Modules.scala 53:83:@3366.4]
  wire [11:0] _T_57193; // @[Modules.scala 53:83:@3368.4]
  wire [10:0] _T_57194; // @[Modules.scala 53:83:@3369.4]
  wire [10:0] buffer_0_665; // @[Modules.scala 53:83:@3370.4]
  wire [11:0] _T_57196; // @[Modules.scala 53:83:@3372.4]
  wire [10:0] _T_57197; // @[Modules.scala 53:83:@3373.4]
  wire [10:0] buffer_0_666; // @[Modules.scala 53:83:@3374.4]
  wire [11:0] _T_57199; // @[Modules.scala 53:83:@3376.4]
  wire [10:0] _T_57200; // @[Modules.scala 53:83:@3377.4]
  wire [10:0] buffer_0_667; // @[Modules.scala 53:83:@3378.4]
  wire [11:0] _T_57202; // @[Modules.scala 53:83:@3380.4]
  wire [10:0] _T_57203; // @[Modules.scala 53:83:@3381.4]
  wire [10:0] buffer_0_668; // @[Modules.scala 53:83:@3382.4]
  wire [11:0] _T_57205; // @[Modules.scala 53:83:@3384.4]
  wire [10:0] _T_57206; // @[Modules.scala 53:83:@3385.4]
  wire [10:0] buffer_0_669; // @[Modules.scala 53:83:@3386.4]
  wire [11:0] _T_57208; // @[Modules.scala 53:83:@3388.4]
  wire [10:0] _T_57209; // @[Modules.scala 53:83:@3389.4]
  wire [10:0] buffer_0_670; // @[Modules.scala 53:83:@3390.4]
  wire [11:0] _T_57211; // @[Modules.scala 53:83:@3392.4]
  wire [10:0] _T_57212; // @[Modules.scala 53:83:@3393.4]
  wire [10:0] buffer_0_671; // @[Modules.scala 53:83:@3394.4]
  wire [11:0] _T_57214; // @[Modules.scala 53:83:@3396.4]
  wire [10:0] _T_57215; // @[Modules.scala 53:83:@3397.4]
  wire [10:0] buffer_0_672; // @[Modules.scala 53:83:@3398.4]
  wire [11:0] _T_57217; // @[Modules.scala 53:83:@3400.4]
  wire [10:0] _T_57218; // @[Modules.scala 53:83:@3401.4]
  wire [10:0] buffer_0_673; // @[Modules.scala 53:83:@3402.4]
  wire [11:0] _T_57220; // @[Modules.scala 53:83:@3404.4]
  wire [10:0] _T_57221; // @[Modules.scala 53:83:@3405.4]
  wire [10:0] buffer_0_674; // @[Modules.scala 53:83:@3406.4]
  wire [11:0] _T_57223; // @[Modules.scala 53:83:@3408.4]
  wire [10:0] _T_57224; // @[Modules.scala 53:83:@3409.4]
  wire [10:0] buffer_0_675; // @[Modules.scala 53:83:@3410.4]
  wire [11:0] _T_57226; // @[Modules.scala 53:83:@3412.4]
  wire [10:0] _T_57227; // @[Modules.scala 53:83:@3413.4]
  wire [10:0] buffer_0_676; // @[Modules.scala 53:83:@3414.4]
  wire [11:0] _T_57229; // @[Modules.scala 53:83:@3416.4]
  wire [10:0] _T_57230; // @[Modules.scala 53:83:@3417.4]
  wire [10:0] buffer_0_677; // @[Modules.scala 53:83:@3418.4]
  wire [11:0] _T_57232; // @[Modules.scala 53:83:@3420.4]
  wire [10:0] _T_57233; // @[Modules.scala 53:83:@3421.4]
  wire [10:0] buffer_0_678; // @[Modules.scala 53:83:@3422.4]
  wire [11:0] _T_57235; // @[Modules.scala 53:83:@3424.4]
  wire [10:0] _T_57236; // @[Modules.scala 53:83:@3425.4]
  wire [10:0] buffer_0_679; // @[Modules.scala 53:83:@3426.4]
  wire [11:0] _T_57238; // @[Modules.scala 53:83:@3428.4]
  wire [10:0] _T_57239; // @[Modules.scala 53:83:@3429.4]
  wire [10:0] buffer_0_680; // @[Modules.scala 53:83:@3430.4]
  wire [11:0] _T_57241; // @[Modules.scala 53:83:@3432.4]
  wire [10:0] _T_57242; // @[Modules.scala 53:83:@3433.4]
  wire [10:0] buffer_0_681; // @[Modules.scala 53:83:@3434.4]
  wire [11:0] _T_57244; // @[Modules.scala 53:83:@3436.4]
  wire [10:0] _T_57245; // @[Modules.scala 53:83:@3437.4]
  wire [10:0] buffer_0_682; // @[Modules.scala 53:83:@3438.4]
  wire [11:0] _T_57247; // @[Modules.scala 53:83:@3440.4]
  wire [10:0] _T_57248; // @[Modules.scala 53:83:@3441.4]
  wire [10:0] buffer_0_683; // @[Modules.scala 53:83:@3442.4]
  wire [11:0] _T_57250; // @[Modules.scala 53:83:@3444.4]
  wire [10:0] _T_57251; // @[Modules.scala 53:83:@3445.4]
  wire [10:0] buffer_0_684; // @[Modules.scala 53:83:@3446.4]
  wire [11:0] _T_57253; // @[Modules.scala 53:83:@3448.4]
  wire [10:0] _T_57254; // @[Modules.scala 53:83:@3449.4]
  wire [10:0] buffer_0_685; // @[Modules.scala 53:83:@3450.4]
  wire [11:0] _T_57256; // @[Modules.scala 56:109:@3452.4]
  wire [10:0] _T_57257; // @[Modules.scala 56:109:@3453.4]
  wire [10:0] buffer_0_686; // @[Modules.scala 56:109:@3454.4]
  wire [11:0] _T_57259; // @[Modules.scala 56:109:@3456.4]
  wire [10:0] _T_57260; // @[Modules.scala 56:109:@3457.4]
  wire [10:0] buffer_0_687; // @[Modules.scala 56:109:@3458.4]
  wire [11:0] _T_57262; // @[Modules.scala 56:109:@3460.4]
  wire [10:0] _T_57263; // @[Modules.scala 56:109:@3461.4]
  wire [10:0] buffer_0_688; // @[Modules.scala 56:109:@3462.4]
  wire [11:0] _T_57265; // @[Modules.scala 56:109:@3464.4]
  wire [10:0] _T_57266; // @[Modules.scala 56:109:@3465.4]
  wire [10:0] buffer_0_689; // @[Modules.scala 56:109:@3466.4]
  wire [11:0] _T_57268; // @[Modules.scala 56:109:@3468.4]
  wire [10:0] _T_57269; // @[Modules.scala 56:109:@3469.4]
  wire [10:0] buffer_0_690; // @[Modules.scala 56:109:@3470.4]
  wire [11:0] _T_57271; // @[Modules.scala 56:109:@3472.4]
  wire [10:0] _T_57272; // @[Modules.scala 56:109:@3473.4]
  wire [10:0] buffer_0_691; // @[Modules.scala 56:109:@3474.4]
  wire [11:0] _T_57274; // @[Modules.scala 56:109:@3476.4]
  wire [10:0] _T_57275; // @[Modules.scala 56:109:@3477.4]
  wire [10:0] buffer_0_692; // @[Modules.scala 56:109:@3478.4]
  wire [11:0] _T_57277; // @[Modules.scala 56:109:@3480.4]
  wire [10:0] _T_57278; // @[Modules.scala 56:109:@3481.4]
  wire [10:0] buffer_0_693; // @[Modules.scala 56:109:@3482.4]
  wire [11:0] _T_57280; // @[Modules.scala 56:109:@3484.4]
  wire [10:0] _T_57281; // @[Modules.scala 56:109:@3485.4]
  wire [10:0] buffer_0_694; // @[Modules.scala 56:109:@3486.4]
  wire [11:0] _T_57283; // @[Modules.scala 56:109:@3488.4]
  wire [10:0] _T_57284; // @[Modules.scala 56:109:@3489.4]
  wire [10:0] buffer_0_695; // @[Modules.scala 56:109:@3490.4]
  wire [11:0] _T_57286; // @[Modules.scala 56:109:@3492.4]
  wire [10:0] _T_57287; // @[Modules.scala 56:109:@3493.4]
  wire [10:0] buffer_0_696; // @[Modules.scala 56:109:@3494.4]
  wire [11:0] _T_57289; // @[Modules.scala 56:109:@3496.4]
  wire [10:0] _T_57290; // @[Modules.scala 56:109:@3497.4]
  wire [10:0] buffer_0_697; // @[Modules.scala 56:109:@3498.4]
  wire [11:0] _T_57292; // @[Modules.scala 56:109:@3500.4]
  wire [10:0] _T_57293; // @[Modules.scala 56:109:@3501.4]
  wire [10:0] buffer_0_698; // @[Modules.scala 56:109:@3502.4]
  wire [11:0] _T_57295; // @[Modules.scala 56:109:@3504.4]
  wire [10:0] _T_57296; // @[Modules.scala 56:109:@3505.4]
  wire [10:0] buffer_0_699; // @[Modules.scala 56:109:@3506.4]
  wire [11:0] _T_57298; // @[Modules.scala 56:109:@3508.4]
  wire [10:0] _T_57299; // @[Modules.scala 56:109:@3509.4]
  wire [10:0] buffer_0_700; // @[Modules.scala 56:109:@3510.4]
  wire [11:0] _T_57301; // @[Modules.scala 56:109:@3512.4]
  wire [10:0] _T_57302; // @[Modules.scala 56:109:@3513.4]
  wire [10:0] buffer_0_701; // @[Modules.scala 56:109:@3514.4]
  wire [11:0] _T_57304; // @[Modules.scala 56:109:@3516.4]
  wire [10:0] _T_57305; // @[Modules.scala 56:109:@3517.4]
  wire [10:0] buffer_0_702; // @[Modules.scala 56:109:@3518.4]
  wire [11:0] _T_57307; // @[Modules.scala 56:109:@3520.4]
  wire [10:0] _T_57308; // @[Modules.scala 56:109:@3521.4]
  wire [10:0] buffer_0_703; // @[Modules.scala 56:109:@3522.4]
  wire [11:0] _T_57310; // @[Modules.scala 56:109:@3524.4]
  wire [10:0] _T_57311; // @[Modules.scala 56:109:@3525.4]
  wire [10:0] buffer_0_704; // @[Modules.scala 56:109:@3526.4]
  wire [11:0] _T_57313; // @[Modules.scala 56:109:@3528.4]
  wire [10:0] _T_57314; // @[Modules.scala 56:109:@3529.4]
  wire [10:0] buffer_0_705; // @[Modules.scala 56:109:@3530.4]
  wire [11:0] _T_57316; // @[Modules.scala 56:109:@3532.4]
  wire [10:0] _T_57317; // @[Modules.scala 56:109:@3533.4]
  wire [10:0] buffer_0_706; // @[Modules.scala 56:109:@3534.4]
  wire [11:0] _T_57319; // @[Modules.scala 56:109:@3536.4]
  wire [10:0] _T_57320; // @[Modules.scala 56:109:@3537.4]
  wire [10:0] buffer_0_707; // @[Modules.scala 56:109:@3538.4]
  wire [11:0] _T_57322; // @[Modules.scala 56:109:@3540.4]
  wire [10:0] _T_57323; // @[Modules.scala 56:109:@3541.4]
  wire [10:0] buffer_0_708; // @[Modules.scala 56:109:@3542.4]
  wire [11:0] _T_57325; // @[Modules.scala 56:109:@3544.4]
  wire [10:0] _T_57326; // @[Modules.scala 56:109:@3545.4]
  wire [10:0] buffer_0_709; // @[Modules.scala 56:109:@3546.4]
  wire [11:0] _T_57328; // @[Modules.scala 56:109:@3548.4]
  wire [10:0] _T_57329; // @[Modules.scala 56:109:@3549.4]
  wire [10:0] buffer_0_710; // @[Modules.scala 56:109:@3550.4]
  wire [11:0] _T_57331; // @[Modules.scala 56:109:@3552.4]
  wire [10:0] _T_57332; // @[Modules.scala 56:109:@3553.4]
  wire [10:0] buffer_0_711; // @[Modules.scala 56:109:@3554.4]
  wire [11:0] _T_57334; // @[Modules.scala 56:109:@3556.4]
  wire [10:0] _T_57335; // @[Modules.scala 56:109:@3557.4]
  wire [10:0] buffer_0_712; // @[Modules.scala 56:109:@3558.4]
  wire [11:0] _T_57337; // @[Modules.scala 56:109:@3560.4]
  wire [10:0] _T_57338; // @[Modules.scala 56:109:@3561.4]
  wire [10:0] buffer_0_713; // @[Modules.scala 56:109:@3562.4]
  wire [11:0] _T_57340; // @[Modules.scala 56:109:@3564.4]
  wire [10:0] _T_57341; // @[Modules.scala 56:109:@3565.4]
  wire [10:0] buffer_0_714; // @[Modules.scala 56:109:@3566.4]
  wire [11:0] _T_57343; // @[Modules.scala 56:109:@3568.4]
  wire [10:0] _T_57344; // @[Modules.scala 56:109:@3569.4]
  wire [10:0] buffer_0_715; // @[Modules.scala 56:109:@3570.4]
  wire [11:0] _T_57346; // @[Modules.scala 56:109:@3572.4]
  wire [10:0] _T_57347; // @[Modules.scala 56:109:@3573.4]
  wire [10:0] buffer_0_716; // @[Modules.scala 56:109:@3574.4]
  wire [11:0] _T_57349; // @[Modules.scala 56:109:@3576.4]
  wire [10:0] _T_57350; // @[Modules.scala 56:109:@3577.4]
  wire [10:0] buffer_0_717; // @[Modules.scala 56:109:@3578.4]
  wire [11:0] _T_57352; // @[Modules.scala 56:109:@3580.4]
  wire [10:0] _T_57353; // @[Modules.scala 56:109:@3581.4]
  wire [10:0] buffer_0_718; // @[Modules.scala 56:109:@3582.4]
  wire [11:0] _T_57355; // @[Modules.scala 56:109:@3584.4]
  wire [10:0] _T_57356; // @[Modules.scala 56:109:@3585.4]
  wire [10:0] buffer_0_719; // @[Modules.scala 56:109:@3586.4]
  wire [11:0] _T_57358; // @[Modules.scala 56:109:@3588.4]
  wire [10:0] _T_57359; // @[Modules.scala 56:109:@3589.4]
  wire [10:0] buffer_0_720; // @[Modules.scala 56:109:@3590.4]
  wire [11:0] _T_57361; // @[Modules.scala 56:109:@3592.4]
  wire [10:0] _T_57362; // @[Modules.scala 56:109:@3593.4]
  wire [10:0] buffer_0_721; // @[Modules.scala 56:109:@3594.4]
  wire [11:0] _T_57364; // @[Modules.scala 56:109:@3596.4]
  wire [10:0] _T_57365; // @[Modules.scala 56:109:@3597.4]
  wire [10:0] buffer_0_722; // @[Modules.scala 56:109:@3598.4]
  wire [11:0] _T_57367; // @[Modules.scala 56:109:@3600.4]
  wire [10:0] _T_57368; // @[Modules.scala 56:109:@3601.4]
  wire [10:0] buffer_0_723; // @[Modules.scala 56:109:@3602.4]
  wire [11:0] _T_57370; // @[Modules.scala 56:109:@3604.4]
  wire [10:0] _T_57371; // @[Modules.scala 56:109:@3605.4]
  wire [10:0] buffer_0_724; // @[Modules.scala 56:109:@3606.4]
  wire [11:0] _T_57373; // @[Modules.scala 56:109:@3608.4]
  wire [10:0] _T_57374; // @[Modules.scala 56:109:@3609.4]
  wire [10:0] buffer_0_725; // @[Modules.scala 56:109:@3610.4]
  wire [11:0] _T_57376; // @[Modules.scala 56:109:@3612.4]
  wire [10:0] _T_57377; // @[Modules.scala 56:109:@3613.4]
  wire [10:0] buffer_0_726; // @[Modules.scala 56:109:@3614.4]
  wire [11:0] _T_57379; // @[Modules.scala 56:109:@3616.4]
  wire [10:0] _T_57380; // @[Modules.scala 56:109:@3617.4]
  wire [10:0] buffer_0_727; // @[Modules.scala 56:109:@3618.4]
  wire [11:0] _T_57382; // @[Modules.scala 56:109:@3620.4]
  wire [10:0] _T_57383; // @[Modules.scala 56:109:@3621.4]
  wire [10:0] buffer_0_728; // @[Modules.scala 56:109:@3622.4]
  wire [11:0] _T_57385; // @[Modules.scala 56:109:@3624.4]
  wire [10:0] _T_57386; // @[Modules.scala 56:109:@3625.4]
  wire [10:0] buffer_0_729; // @[Modules.scala 56:109:@3626.4]
  wire [11:0] _T_57388; // @[Modules.scala 56:109:@3628.4]
  wire [10:0] _T_57389; // @[Modules.scala 56:109:@3629.4]
  wire [10:0] buffer_0_730; // @[Modules.scala 56:109:@3630.4]
  wire [11:0] _T_57391; // @[Modules.scala 56:109:@3632.4]
  wire [10:0] _T_57392; // @[Modules.scala 56:109:@3633.4]
  wire [10:0] buffer_0_731; // @[Modules.scala 56:109:@3634.4]
  wire [11:0] _T_57394; // @[Modules.scala 56:109:@3636.4]
  wire [10:0] _T_57395; // @[Modules.scala 56:109:@3637.4]
  wire [10:0] buffer_0_732; // @[Modules.scala 56:109:@3638.4]
  wire [11:0] _T_57397; // @[Modules.scala 56:109:@3640.4]
  wire [10:0] _T_57398; // @[Modules.scala 56:109:@3641.4]
  wire [10:0] buffer_0_733; // @[Modules.scala 56:109:@3642.4]
  wire [11:0] _T_57400; // @[Modules.scala 56:109:@3644.4]
  wire [10:0] _T_57401; // @[Modules.scala 56:109:@3645.4]
  wire [10:0] buffer_0_734; // @[Modules.scala 56:109:@3646.4]
  wire [11:0] _T_57403; // @[Modules.scala 63:156:@3649.4]
  wire [10:0] _T_57404; // @[Modules.scala 63:156:@3650.4]
  wire [10:0] buffer_0_736; // @[Modules.scala 63:156:@3651.4]
  wire [11:0] _T_57406; // @[Modules.scala 63:156:@3653.4]
  wire [10:0] _T_57407; // @[Modules.scala 63:156:@3654.4]
  wire [10:0] buffer_0_737; // @[Modules.scala 63:156:@3655.4]
  wire [11:0] _T_57409; // @[Modules.scala 63:156:@3657.4]
  wire [10:0] _T_57410; // @[Modules.scala 63:156:@3658.4]
  wire [10:0] buffer_0_738; // @[Modules.scala 63:156:@3659.4]
  wire [11:0] _T_57412; // @[Modules.scala 63:156:@3661.4]
  wire [10:0] _T_57413; // @[Modules.scala 63:156:@3662.4]
  wire [10:0] buffer_0_739; // @[Modules.scala 63:156:@3663.4]
  wire [11:0] _T_57415; // @[Modules.scala 63:156:@3665.4]
  wire [10:0] _T_57416; // @[Modules.scala 63:156:@3666.4]
  wire [10:0] buffer_0_740; // @[Modules.scala 63:156:@3667.4]
  wire [11:0] _T_57418; // @[Modules.scala 63:156:@3669.4]
  wire [10:0] _T_57419; // @[Modules.scala 63:156:@3670.4]
  wire [10:0] buffer_0_741; // @[Modules.scala 63:156:@3671.4]
  wire [11:0] _T_57421; // @[Modules.scala 63:156:@3673.4]
  wire [10:0] _T_57422; // @[Modules.scala 63:156:@3674.4]
  wire [10:0] buffer_0_742; // @[Modules.scala 63:156:@3675.4]
  wire [11:0] _T_57424; // @[Modules.scala 63:156:@3677.4]
  wire [10:0] _T_57425; // @[Modules.scala 63:156:@3678.4]
  wire [10:0] buffer_0_743; // @[Modules.scala 63:156:@3679.4]
  wire [11:0] _T_57427; // @[Modules.scala 63:156:@3681.4]
  wire [10:0] _T_57428; // @[Modules.scala 63:156:@3682.4]
  wire [10:0] buffer_0_744; // @[Modules.scala 63:156:@3683.4]
  wire [11:0] _T_57430; // @[Modules.scala 63:156:@3685.4]
  wire [10:0] _T_57431; // @[Modules.scala 63:156:@3686.4]
  wire [10:0] buffer_0_745; // @[Modules.scala 63:156:@3687.4]
  wire [11:0] _T_57433; // @[Modules.scala 63:156:@3689.4]
  wire [10:0] _T_57434; // @[Modules.scala 63:156:@3690.4]
  wire [10:0] buffer_0_746; // @[Modules.scala 63:156:@3691.4]
  wire [11:0] _T_57436; // @[Modules.scala 63:156:@3693.4]
  wire [10:0] _T_57437; // @[Modules.scala 63:156:@3694.4]
  wire [10:0] buffer_0_747; // @[Modules.scala 63:156:@3695.4]
  wire [11:0] _T_57439; // @[Modules.scala 63:156:@3697.4]
  wire [10:0] _T_57440; // @[Modules.scala 63:156:@3698.4]
  wire [10:0] buffer_0_748; // @[Modules.scala 63:156:@3699.4]
  wire [11:0] _T_57442; // @[Modules.scala 63:156:@3701.4]
  wire [10:0] _T_57443; // @[Modules.scala 63:156:@3702.4]
  wire [10:0] buffer_0_749; // @[Modules.scala 63:156:@3703.4]
  wire [11:0] _T_57445; // @[Modules.scala 63:156:@3705.4]
  wire [10:0] _T_57446; // @[Modules.scala 63:156:@3706.4]
  wire [10:0] buffer_0_750; // @[Modules.scala 63:156:@3707.4]
  wire [11:0] _T_57448; // @[Modules.scala 63:156:@3709.4]
  wire [10:0] _T_57449; // @[Modules.scala 63:156:@3710.4]
  wire [10:0] buffer_0_751; // @[Modules.scala 63:156:@3711.4]
  wire [11:0] _T_57451; // @[Modules.scala 63:156:@3713.4]
  wire [10:0] _T_57452; // @[Modules.scala 63:156:@3714.4]
  wire [10:0] buffer_0_752; // @[Modules.scala 63:156:@3715.4]
  wire [11:0] _T_57454; // @[Modules.scala 63:156:@3717.4]
  wire [10:0] _T_57455; // @[Modules.scala 63:156:@3718.4]
  wire [10:0] buffer_0_753; // @[Modules.scala 63:156:@3719.4]
  wire [11:0] _T_57457; // @[Modules.scala 63:156:@3721.4]
  wire [10:0] _T_57458; // @[Modules.scala 63:156:@3722.4]
  wire [10:0] buffer_0_754; // @[Modules.scala 63:156:@3723.4]
  wire [11:0] _T_57460; // @[Modules.scala 63:156:@3725.4]
  wire [10:0] _T_57461; // @[Modules.scala 63:156:@3726.4]
  wire [10:0] buffer_0_755; // @[Modules.scala 63:156:@3727.4]
  wire [11:0] _T_57463; // @[Modules.scala 63:156:@3729.4]
  wire [10:0] _T_57464; // @[Modules.scala 63:156:@3730.4]
  wire [10:0] buffer_0_756; // @[Modules.scala 63:156:@3731.4]
  wire [11:0] _T_57466; // @[Modules.scala 63:156:@3733.4]
  wire [10:0] _T_57467; // @[Modules.scala 63:156:@3734.4]
  wire [10:0] buffer_0_757; // @[Modules.scala 63:156:@3735.4]
  wire [11:0] _T_57469; // @[Modules.scala 63:156:@3737.4]
  wire [10:0] _T_57470; // @[Modules.scala 63:156:@3738.4]
  wire [10:0] buffer_0_758; // @[Modules.scala 63:156:@3739.4]
  wire [11:0] _T_57472; // @[Modules.scala 63:156:@3741.4]
  wire [10:0] _T_57473; // @[Modules.scala 63:156:@3742.4]
  wire [10:0] buffer_0_759; // @[Modules.scala 63:156:@3743.4]
  wire [11:0] _T_57475; // @[Modules.scala 63:156:@3745.4]
  wire [10:0] _T_57476; // @[Modules.scala 63:156:@3746.4]
  wire [10:0] buffer_0_760; // @[Modules.scala 63:156:@3747.4]
  wire [11:0] _T_57478; // @[Modules.scala 63:156:@3749.4]
  wire [10:0] _T_57479; // @[Modules.scala 63:156:@3750.4]
  wire [10:0] buffer_0_761; // @[Modules.scala 63:156:@3751.4]
  wire [11:0] _T_57481; // @[Modules.scala 63:156:@3753.4]
  wire [10:0] _T_57482; // @[Modules.scala 63:156:@3754.4]
  wire [10:0] buffer_0_762; // @[Modules.scala 63:156:@3755.4]
  wire [11:0] _T_57484; // @[Modules.scala 63:156:@3757.4]
  wire [10:0] _T_57485; // @[Modules.scala 63:156:@3758.4]
  wire [10:0] buffer_0_763; // @[Modules.scala 63:156:@3759.4]
  wire [11:0] _T_57487; // @[Modules.scala 63:156:@3761.4]
  wire [10:0] _T_57488; // @[Modules.scala 63:156:@3762.4]
  wire [10:0] buffer_0_764; // @[Modules.scala 63:156:@3763.4]
  wire [11:0] _T_57490; // @[Modules.scala 63:156:@3765.4]
  wire [10:0] _T_57491; // @[Modules.scala 63:156:@3766.4]
  wire [10:0] buffer_0_765; // @[Modules.scala 63:156:@3767.4]
  wire [11:0] _T_57493; // @[Modules.scala 63:156:@3769.4]
  wire [10:0] _T_57494; // @[Modules.scala 63:156:@3770.4]
  wire [10:0] buffer_0_766; // @[Modules.scala 63:156:@3771.4]
  wire [11:0] _T_57496; // @[Modules.scala 63:156:@3773.4]
  wire [10:0] _T_57497; // @[Modules.scala 63:156:@3774.4]
  wire [10:0] buffer_0_767; // @[Modules.scala 63:156:@3775.4]
  wire [11:0] _T_57499; // @[Modules.scala 63:156:@3777.4]
  wire [10:0] _T_57500; // @[Modules.scala 63:156:@3778.4]
  wire [10:0] buffer_0_768; // @[Modules.scala 63:156:@3779.4]
  wire [11:0] _T_57502; // @[Modules.scala 63:156:@3781.4]
  wire [10:0] _T_57503; // @[Modules.scala 63:156:@3782.4]
  wire [10:0] buffer_0_769; // @[Modules.scala 63:156:@3783.4]
  wire [11:0] _T_57505; // @[Modules.scala 63:156:@3785.4]
  wire [10:0] _T_57506; // @[Modules.scala 63:156:@3786.4]
  wire [10:0] buffer_0_770; // @[Modules.scala 63:156:@3787.4]
  wire [11:0] _T_57508; // @[Modules.scala 63:156:@3789.4]
  wire [10:0] _T_57509; // @[Modules.scala 63:156:@3790.4]
  wire [10:0] buffer_0_771; // @[Modules.scala 63:156:@3791.4]
  wire [11:0] _T_57511; // @[Modules.scala 63:156:@3793.4]
  wire [10:0] _T_57512; // @[Modules.scala 63:156:@3794.4]
  wire [10:0] buffer_0_772; // @[Modules.scala 63:156:@3795.4]
  wire [11:0] _T_57514; // @[Modules.scala 63:156:@3797.4]
  wire [10:0] _T_57515; // @[Modules.scala 63:156:@3798.4]
  wire [10:0] buffer_0_773; // @[Modules.scala 63:156:@3799.4]
  wire [11:0] _T_57517; // @[Modules.scala 63:156:@3801.4]
  wire [10:0] _T_57518; // @[Modules.scala 63:156:@3802.4]
  wire [10:0] buffer_0_774; // @[Modules.scala 63:156:@3803.4]
  wire [11:0] _T_57520; // @[Modules.scala 63:156:@3805.4]
  wire [10:0] _T_57521; // @[Modules.scala 63:156:@3806.4]
  wire [10:0] buffer_0_775; // @[Modules.scala 63:156:@3807.4]
  wire [11:0] _T_57523; // @[Modules.scala 63:156:@3809.4]
  wire [10:0] _T_57524; // @[Modules.scala 63:156:@3810.4]
  wire [10:0] buffer_0_776; // @[Modules.scala 63:156:@3811.4]
  wire [11:0] _T_57526; // @[Modules.scala 63:156:@3813.4]
  wire [10:0] _T_57527; // @[Modules.scala 63:156:@3814.4]
  wire [10:0] buffer_0_777; // @[Modules.scala 63:156:@3815.4]
  wire [11:0] _T_57529; // @[Modules.scala 63:156:@3817.4]
  wire [10:0] _T_57530; // @[Modules.scala 63:156:@3818.4]
  wire [10:0] buffer_0_778; // @[Modules.scala 63:156:@3819.4]
  wire [11:0] _T_57532; // @[Modules.scala 63:156:@3821.4]
  wire [10:0] _T_57533; // @[Modules.scala 63:156:@3822.4]
  wire [10:0] buffer_0_779; // @[Modules.scala 63:156:@3823.4]
  wire [11:0] _T_57535; // @[Modules.scala 63:156:@3825.4]
  wire [10:0] _T_57536; // @[Modules.scala 63:156:@3826.4]
  wire [10:0] buffer_0_780; // @[Modules.scala 63:156:@3827.4]
  wire [11:0] _T_57538; // @[Modules.scala 63:156:@3829.4]
  wire [10:0] _T_57539; // @[Modules.scala 63:156:@3830.4]
  wire [10:0] buffer_0_781; // @[Modules.scala 63:156:@3831.4]
  wire [11:0] _T_57541; // @[Modules.scala 63:156:@3833.4]
  wire [10:0] _T_57542; // @[Modules.scala 63:156:@3834.4]
  wire [10:0] buffer_0_782; // @[Modules.scala 63:156:@3835.4]
  wire [11:0] _T_57544; // @[Modules.scala 63:156:@3837.4]
  wire [10:0] _T_57545; // @[Modules.scala 63:156:@3838.4]
  wire [10:0] buffer_0_783; // @[Modules.scala 63:156:@3839.4]
  wire [5:0] _T_57551; // @[Modules.scala 46:47:@3845.4]
  wire [4:0] _T_57552; // @[Modules.scala 46:47:@3846.4]
  wire [4:0] _T_57553; // @[Modules.scala 46:47:@3847.4]
  wire [5:0] _T_57561; // @[Modules.scala 37:46:@3856.4]
  wire [4:0] _T_57562; // @[Modules.scala 37:46:@3857.4]
  wire [4:0] _T_57563; // @[Modules.scala 37:46:@3858.4]
  wire [5:0] _T_57564; // @[Modules.scala 37:46:@3860.4]
  wire [4:0] _T_57565; // @[Modules.scala 37:46:@3861.4]
  wire [4:0] _T_57566; // @[Modules.scala 37:46:@3862.4]
  wire [5:0] _T_57567; // @[Modules.scala 37:46:@3864.4]
  wire [4:0] _T_57568; // @[Modules.scala 37:46:@3865.4]
  wire [4:0] _T_57569; // @[Modules.scala 37:46:@3866.4]
  wire [5:0] _T_57577; // @[Modules.scala 37:46:@3875.4]
  wire [4:0] _T_57578; // @[Modules.scala 37:46:@3876.4]
  wire [4:0] _T_57579; // @[Modules.scala 37:46:@3877.4]
  wire [5:0] _T_57580; // @[Modules.scala 37:46:@3879.4]
  wire [4:0] _T_57581; // @[Modules.scala 37:46:@3880.4]
  wire [4:0] _T_57582; // @[Modules.scala 37:46:@3881.4]
  wire [5:0] _T_57583; // @[Modules.scala 40:46:@3883.4]
  wire [4:0] _T_57584; // @[Modules.scala 40:46:@3884.4]
  wire [4:0] _T_57585; // @[Modules.scala 40:46:@3885.4]
  wire [5:0] _T_57586; // @[Modules.scala 40:46:@3887.4]
  wire [4:0] _T_57587; // @[Modules.scala 40:46:@3888.4]
  wire [4:0] _T_57588; // @[Modules.scala 40:46:@3889.4]
  wire [5:0] _T_57592; // @[Modules.scala 40:46:@3895.4]
  wire [4:0] _T_57593; // @[Modules.scala 40:46:@3896.4]
  wire [4:0] _T_57594; // @[Modules.scala 40:46:@3897.4]
  wire [5:0] _T_57595; // @[Modules.scala 37:46:@3899.4]
  wire [4:0] _T_57596; // @[Modules.scala 37:46:@3900.4]
  wire [4:0] _T_57597; // @[Modules.scala 37:46:@3901.4]
  wire [5:0] _T_57599; // @[Modules.scala 46:37:@3903.4]
  wire [4:0] _T_57600; // @[Modules.scala 46:37:@3904.4]
  wire [4:0] _T_57601; // @[Modules.scala 46:37:@3905.4]
  wire [5:0] _T_57602; // @[Modules.scala 46:47:@3906.4]
  wire [4:0] _T_57603; // @[Modules.scala 46:47:@3907.4]
  wire [4:0] _T_57604; // @[Modules.scala 46:47:@3908.4]
  wire [5:0] _T_57605; // @[Modules.scala 40:46:@3910.4]
  wire [4:0] _T_57606; // @[Modules.scala 40:46:@3911.4]
  wire [4:0] _T_57607; // @[Modules.scala 40:46:@3912.4]
  wire [5:0] _T_57608; // @[Modules.scala 37:46:@3914.4]
  wire [4:0] _T_57609; // @[Modules.scala 37:46:@3915.4]
  wire [4:0] _T_57610; // @[Modules.scala 37:46:@3916.4]
  wire [5:0] _T_57614; // @[Modules.scala 37:46:@3922.4]
  wire [4:0] _T_57615; // @[Modules.scala 37:46:@3923.4]
  wire [4:0] _T_57616; // @[Modules.scala 37:46:@3924.4]
  wire [5:0] _T_57617; // @[Modules.scala 37:46:@3926.4]
  wire [4:0] _T_57618; // @[Modules.scala 37:46:@3927.4]
  wire [4:0] _T_57619; // @[Modules.scala 37:46:@3928.4]
  wire [5:0] _T_57620; // @[Modules.scala 37:46:@3930.4]
  wire [4:0] _T_57621; // @[Modules.scala 37:46:@3931.4]
  wire [4:0] _T_57622; // @[Modules.scala 37:46:@3932.4]
  wire [5:0] _T_57623; // @[Modules.scala 37:46:@3934.4]
  wire [4:0] _T_57624; // @[Modules.scala 37:46:@3935.4]
  wire [4:0] _T_57625; // @[Modules.scala 37:46:@3936.4]
  wire [5:0] _T_57626; // @[Modules.scala 37:46:@3938.4]
  wire [4:0] _T_57627; // @[Modules.scala 37:46:@3939.4]
  wire [4:0] _T_57628; // @[Modules.scala 37:46:@3940.4]
  wire [5:0] _T_57633; // @[Modules.scala 43:47:@3945.4]
  wire [4:0] _T_57634; // @[Modules.scala 43:47:@3946.4]
  wire [4:0] _T_57635; // @[Modules.scala 43:47:@3947.4]
  wire [5:0] _T_57636; // @[Modules.scala 37:46:@3949.4]
  wire [4:0] _T_57637; // @[Modules.scala 37:46:@3950.4]
  wire [4:0] _T_57638; // @[Modules.scala 37:46:@3951.4]
  wire [5:0] _T_57639; // @[Modules.scala 37:46:@3953.4]
  wire [4:0] _T_57640; // @[Modules.scala 37:46:@3954.4]
  wire [4:0] _T_57641; // @[Modules.scala 37:46:@3955.4]
  wire [5:0] _T_57642; // @[Modules.scala 37:46:@3957.4]
  wire [4:0] _T_57643; // @[Modules.scala 37:46:@3958.4]
  wire [4:0] _T_57644; // @[Modules.scala 37:46:@3959.4]
  wire [5:0] _T_57645; // @[Modules.scala 40:46:@3961.4]
  wire [4:0] _T_57646; // @[Modules.scala 40:46:@3962.4]
  wire [4:0] _T_57647; // @[Modules.scala 40:46:@3963.4]
  wire [5:0] _T_57649; // @[Modules.scala 43:37:@3965.4]
  wire [4:0] _T_57650; // @[Modules.scala 43:37:@3966.4]
  wire [4:0] _T_57651; // @[Modules.scala 43:37:@3967.4]
  wire [5:0] _T_57652; // @[Modules.scala 43:47:@3968.4]
  wire [4:0] _T_57653; // @[Modules.scala 43:47:@3969.4]
  wire [4:0] _T_57654; // @[Modules.scala 43:47:@3970.4]
  wire [5:0] _T_57656; // @[Modules.scala 43:37:@3972.4]
  wire [4:0] _T_57657; // @[Modules.scala 43:37:@3973.4]
  wire [4:0] _T_57658; // @[Modules.scala 43:37:@3974.4]
  wire [5:0] _T_57659; // @[Modules.scala 43:47:@3975.4]
  wire [4:0] _T_57660; // @[Modules.scala 43:47:@3976.4]
  wire [4:0] _T_57661; // @[Modules.scala 43:47:@3977.4]
  wire [5:0] _T_57662; // @[Modules.scala 37:46:@3979.4]
  wire [4:0] _T_57663; // @[Modules.scala 37:46:@3980.4]
  wire [4:0] _T_57664; // @[Modules.scala 37:46:@3981.4]
  wire [5:0] _T_57665; // @[Modules.scala 37:46:@3983.4]
  wire [4:0] _T_57666; // @[Modules.scala 37:46:@3984.4]
  wire [4:0] _T_57667; // @[Modules.scala 37:46:@3985.4]
  wire [5:0] _T_57668; // @[Modules.scala 37:46:@3987.4]
  wire [4:0] _T_57669; // @[Modules.scala 37:46:@3988.4]
  wire [4:0] _T_57670; // @[Modules.scala 37:46:@3989.4]
  wire [5:0] _T_57671; // @[Modules.scala 37:46:@3991.4]
  wire [4:0] _T_57672; // @[Modules.scala 37:46:@3992.4]
  wire [4:0] _T_57673; // @[Modules.scala 37:46:@3993.4]
  wire [5:0] _T_57674; // @[Modules.scala 37:46:@3995.4]
  wire [4:0] _T_57675; // @[Modules.scala 37:46:@3996.4]
  wire [4:0] _T_57676; // @[Modules.scala 37:46:@3997.4]
  wire [5:0] _T_57677; // @[Modules.scala 37:46:@3999.4]
  wire [4:0] _T_57678; // @[Modules.scala 37:46:@4000.4]
  wire [4:0] _T_57679; // @[Modules.scala 37:46:@4001.4]
  wire [5:0] _T_57680; // @[Modules.scala 37:46:@4003.4]
  wire [4:0] _T_57681; // @[Modules.scala 37:46:@4004.4]
  wire [4:0] _T_57682; // @[Modules.scala 37:46:@4005.4]
  wire [5:0] _T_57683; // @[Modules.scala 37:46:@4007.4]
  wire [4:0] _T_57684; // @[Modules.scala 37:46:@4008.4]
  wire [4:0] _T_57685; // @[Modules.scala 37:46:@4009.4]
  wire [5:0] _T_57686; // @[Modules.scala 37:46:@4011.4]
  wire [4:0] _T_57687; // @[Modules.scala 37:46:@4012.4]
  wire [4:0] _T_57688; // @[Modules.scala 37:46:@4013.4]
  wire [5:0] _T_57689; // @[Modules.scala 37:46:@4015.4]
  wire [4:0] _T_57690; // @[Modules.scala 37:46:@4016.4]
  wire [4:0] _T_57691; // @[Modules.scala 37:46:@4017.4]
  wire [5:0] _T_57695; // @[Modules.scala 37:46:@4023.4]
  wire [4:0] _T_57696; // @[Modules.scala 37:46:@4024.4]
  wire [4:0] _T_57697; // @[Modules.scala 37:46:@4025.4]
  wire [5:0] _T_57699; // @[Modules.scala 46:37:@4027.4]
  wire [4:0] _T_57700; // @[Modules.scala 46:37:@4028.4]
  wire [4:0] _T_57701; // @[Modules.scala 46:37:@4029.4]
  wire [5:0] _T_57702; // @[Modules.scala 46:47:@4030.4]
  wire [4:0] _T_57703; // @[Modules.scala 46:47:@4031.4]
  wire [4:0] _T_57704; // @[Modules.scala 46:47:@4032.4]
  wire [5:0] _T_57706; // @[Modules.scala 43:37:@4034.4]
  wire [4:0] _T_57707; // @[Modules.scala 43:37:@4035.4]
  wire [4:0] _T_57708; // @[Modules.scala 43:37:@4036.4]
  wire [5:0] _T_57709; // @[Modules.scala 43:47:@4037.4]
  wire [4:0] _T_57710; // @[Modules.scala 43:47:@4038.4]
  wire [4:0] _T_57711; // @[Modules.scala 43:47:@4039.4]
  wire [5:0] _T_57716; // @[Modules.scala 43:47:@4044.4]
  wire [4:0] _T_57717; // @[Modules.scala 43:47:@4045.4]
  wire [4:0] _T_57718; // @[Modules.scala 43:47:@4046.4]
  wire [5:0] _T_57725; // @[Modules.scala 37:46:@4056.4]
  wire [4:0] _T_57726; // @[Modules.scala 37:46:@4057.4]
  wire [4:0] _T_57727; // @[Modules.scala 37:46:@4058.4]
  wire [5:0] _T_57731; // @[Modules.scala 37:46:@4064.4]
  wire [4:0] _T_57732; // @[Modules.scala 37:46:@4065.4]
  wire [4:0] _T_57733; // @[Modules.scala 37:46:@4066.4]
  wire [5:0] _T_57749; // @[Modules.scala 37:46:@4088.4]
  wire [4:0] _T_57750; // @[Modules.scala 37:46:@4089.4]
  wire [4:0] _T_57751; // @[Modules.scala 37:46:@4090.4]
  wire [5:0] _T_57759; // @[Modules.scala 46:47:@4099.4]
  wire [4:0] _T_57760; // @[Modules.scala 46:47:@4100.4]
  wire [4:0] _T_57761; // @[Modules.scala 46:47:@4101.4]
  wire [5:0] _T_57766; // @[Modules.scala 43:47:@4106.4]
  wire [4:0] _T_57767; // @[Modules.scala 43:47:@4107.4]
  wire [4:0] _T_57768; // @[Modules.scala 43:47:@4108.4]
  wire [5:0] _T_57773; // @[Modules.scala 46:37:@4114.4]
  wire [4:0] _T_57774; // @[Modules.scala 46:37:@4115.4]
  wire [4:0] _T_57775; // @[Modules.scala 46:37:@4116.4]
  wire [5:0] _T_57776; // @[Modules.scala 46:47:@4117.4]
  wire [4:0] _T_57777; // @[Modules.scala 46:47:@4118.4]
  wire [4:0] _T_57778; // @[Modules.scala 46:47:@4119.4]
  wire [5:0] _T_57804; // @[Modules.scala 43:47:@4145.4]
  wire [4:0] _T_57805; // @[Modules.scala 43:47:@4146.4]
  wire [4:0] _T_57806; // @[Modules.scala 43:47:@4147.4]
  wire [5:0] _T_57807; // @[Modules.scala 37:46:@4149.4]
  wire [4:0] _T_57808; // @[Modules.scala 37:46:@4150.4]
  wire [4:0] _T_57809; // @[Modules.scala 37:46:@4151.4]
  wire [5:0] _T_57810; // @[Modules.scala 37:46:@4153.4]
  wire [4:0] _T_57811; // @[Modules.scala 37:46:@4154.4]
  wire [4:0] _T_57812; // @[Modules.scala 37:46:@4155.4]
  wire [5:0] _T_57814; // @[Modules.scala 43:37:@4157.4]
  wire [4:0] _T_57815; // @[Modules.scala 43:37:@4158.4]
  wire [4:0] _T_57816; // @[Modules.scala 43:37:@4159.4]
  wire [5:0] _T_57817; // @[Modules.scala 43:47:@4160.4]
  wire [4:0] _T_57818; // @[Modules.scala 43:47:@4161.4]
  wire [4:0] _T_57819; // @[Modules.scala 43:47:@4162.4]
  wire [5:0] _T_57823; // @[Modules.scala 37:46:@4168.4]
  wire [4:0] _T_57824; // @[Modules.scala 37:46:@4169.4]
  wire [4:0] _T_57825; // @[Modules.scala 37:46:@4170.4]
  wire [5:0] _T_57830; // @[Modules.scala 43:47:@4175.4]
  wire [4:0] _T_57831; // @[Modules.scala 43:47:@4176.4]
  wire [4:0] _T_57832; // @[Modules.scala 43:47:@4177.4]
  wire [5:0] _T_57833; // @[Modules.scala 40:46:@4179.4]
  wire [4:0] _T_57834; // @[Modules.scala 40:46:@4180.4]
  wire [4:0] _T_57835; // @[Modules.scala 40:46:@4181.4]
  wire [5:0] _T_57840; // @[Modules.scala 43:47:@4186.4]
  wire [4:0] _T_57841; // @[Modules.scala 43:47:@4187.4]
  wire [4:0] _T_57842; // @[Modules.scala 43:47:@4188.4]
  wire [5:0] _T_57844; // @[Modules.scala 46:37:@4190.4]
  wire [4:0] _T_57845; // @[Modules.scala 46:37:@4191.4]
  wire [4:0] _T_57846; // @[Modules.scala 46:37:@4192.4]
  wire [5:0] _T_57847; // @[Modules.scala 46:47:@4193.4]
  wire [4:0] _T_57848; // @[Modules.scala 46:47:@4194.4]
  wire [4:0] _T_57849; // @[Modules.scala 46:47:@4195.4]
  wire [5:0] _T_57851; // @[Modules.scala 46:37:@4197.4]
  wire [4:0] _T_57852; // @[Modules.scala 46:37:@4198.4]
  wire [4:0] _T_57853; // @[Modules.scala 46:37:@4199.4]
  wire [5:0] _T_57854; // @[Modules.scala 46:47:@4200.4]
  wire [4:0] _T_57855; // @[Modules.scala 46:47:@4201.4]
  wire [4:0] _T_57856; // @[Modules.scala 46:47:@4202.4]
  wire [5:0] _T_57857; // @[Modules.scala 40:46:@4204.4]
  wire [4:0] _T_57858; // @[Modules.scala 40:46:@4205.4]
  wire [4:0] _T_57859; // @[Modules.scala 40:46:@4206.4]
  wire [5:0] _T_57860; // @[Modules.scala 40:46:@4208.4]
  wire [4:0] _T_57861; // @[Modules.scala 40:46:@4209.4]
  wire [4:0] _T_57862; // @[Modules.scala 40:46:@4210.4]
  wire [5:0] _T_57877; // @[Modules.scala 40:46:@4226.4]
  wire [4:0] _T_57878; // @[Modules.scala 40:46:@4227.4]
  wire [4:0] _T_57879; // @[Modules.scala 40:46:@4228.4]
  wire [5:0] _T_57895; // @[Modules.scala 43:37:@4244.4]
  wire [4:0] _T_57896; // @[Modules.scala 43:37:@4245.4]
  wire [4:0] _T_57897; // @[Modules.scala 43:37:@4246.4]
  wire [5:0] _T_57898; // @[Modules.scala 43:47:@4247.4]
  wire [4:0] _T_57899; // @[Modules.scala 43:47:@4248.4]
  wire [4:0] _T_57900; // @[Modules.scala 43:47:@4249.4]
  wire [5:0] _T_57902; // @[Modules.scala 46:37:@4251.4]
  wire [4:0] _T_57903; // @[Modules.scala 46:37:@4252.4]
  wire [4:0] _T_57904; // @[Modules.scala 46:37:@4253.4]
  wire [5:0] _T_57905; // @[Modules.scala 46:47:@4254.4]
  wire [4:0] _T_57906; // @[Modules.scala 46:47:@4255.4]
  wire [4:0] _T_57907; // @[Modules.scala 46:47:@4256.4]
  wire [5:0] _T_57908; // @[Modules.scala 37:46:@4258.4]
  wire [4:0] _T_57909; // @[Modules.scala 37:46:@4259.4]
  wire [4:0] _T_57910; // @[Modules.scala 37:46:@4260.4]
  wire [5:0] _T_57915; // @[Modules.scala 43:47:@4265.4]
  wire [4:0] _T_57916; // @[Modules.scala 43:47:@4266.4]
  wire [4:0] _T_57917; // @[Modules.scala 43:47:@4267.4]
  wire [5:0] _T_57918; // @[Modules.scala 37:46:@4269.4]
  wire [4:0] _T_57919; // @[Modules.scala 37:46:@4270.4]
  wire [4:0] _T_57920; // @[Modules.scala 37:46:@4271.4]
  wire [5:0] _T_57924; // @[Modules.scala 37:46:@4277.4]
  wire [4:0] _T_57925; // @[Modules.scala 37:46:@4278.4]
  wire [4:0] _T_57926; // @[Modules.scala 37:46:@4279.4]
  wire [5:0] _T_57927; // @[Modules.scala 37:46:@4281.4]
  wire [4:0] _T_57928; // @[Modules.scala 37:46:@4282.4]
  wire [4:0] _T_57929; // @[Modules.scala 37:46:@4283.4]
  wire [5:0] _T_57930; // @[Modules.scala 40:46:@4285.4]
  wire [4:0] _T_57931; // @[Modules.scala 40:46:@4286.4]
  wire [4:0] _T_57932; // @[Modules.scala 40:46:@4287.4]
  wire [5:0] _T_57940; // @[Modules.scala 40:46:@4296.4]
  wire [4:0] _T_57941; // @[Modules.scala 40:46:@4297.4]
  wire [4:0] _T_57942; // @[Modules.scala 40:46:@4298.4]
  wire [5:0] _T_57953; // @[Modules.scala 40:46:@4311.4]
  wire [4:0] _T_57954; // @[Modules.scala 40:46:@4312.4]
  wire [4:0] _T_57955; // @[Modules.scala 40:46:@4313.4]
  wire [5:0] _T_57957; // @[Modules.scala 43:37:@4315.4]
  wire [4:0] _T_57958; // @[Modules.scala 43:37:@4316.4]
  wire [4:0] _T_57959; // @[Modules.scala 43:37:@4317.4]
  wire [5:0] _T_57960; // @[Modules.scala 43:47:@4318.4]
  wire [4:0] _T_57961; // @[Modules.scala 43:47:@4319.4]
  wire [4:0] _T_57962; // @[Modules.scala 43:47:@4320.4]
  wire [5:0] _T_57967; // @[Modules.scala 43:47:@4325.4]
  wire [4:0] _T_57968; // @[Modules.scala 43:47:@4326.4]
  wire [4:0] _T_57969; // @[Modules.scala 43:47:@4327.4]
  wire [5:0] _T_57974; // @[Modules.scala 43:47:@4332.4]
  wire [4:0] _T_57975; // @[Modules.scala 43:47:@4333.4]
  wire [4:0] _T_57976; // @[Modules.scala 43:47:@4334.4]
  wire [5:0] _T_57977; // @[Modules.scala 37:46:@4336.4]
  wire [4:0] _T_57978; // @[Modules.scala 37:46:@4337.4]
  wire [4:0] _T_57979; // @[Modules.scala 37:46:@4338.4]
  wire [5:0] _T_57981; // @[Modules.scala 43:37:@4340.4]
  wire [4:0] _T_57982; // @[Modules.scala 43:37:@4341.4]
  wire [4:0] _T_57983; // @[Modules.scala 43:37:@4342.4]
  wire [5:0] _T_57984; // @[Modules.scala 43:47:@4343.4]
  wire [4:0] _T_57985; // @[Modules.scala 43:47:@4344.4]
  wire [4:0] _T_57986; // @[Modules.scala 43:47:@4345.4]
  wire [5:0] _T_57991; // @[Modules.scala 43:47:@4350.4]
  wire [4:0] _T_57992; // @[Modules.scala 43:47:@4351.4]
  wire [4:0] _T_57993; // @[Modules.scala 43:47:@4352.4]
  wire [5:0] _T_57994; // @[Modules.scala 37:46:@4354.4]
  wire [4:0] _T_57995; // @[Modules.scala 37:46:@4355.4]
  wire [4:0] _T_57996; // @[Modules.scala 37:46:@4356.4]
  wire [5:0] _T_58001; // @[Modules.scala 43:47:@4361.4]
  wire [4:0] _T_58002; // @[Modules.scala 43:47:@4362.4]
  wire [4:0] _T_58003; // @[Modules.scala 43:47:@4363.4]
  wire [5:0] _T_58004; // @[Modules.scala 40:46:@4365.4]
  wire [4:0] _T_58005; // @[Modules.scala 40:46:@4366.4]
  wire [4:0] _T_58006; // @[Modules.scala 40:46:@4367.4]
  wire [5:0] _T_58007; // @[Modules.scala 40:46:@4369.4]
  wire [4:0] _T_58008; // @[Modules.scala 40:46:@4370.4]
  wire [4:0] _T_58009; // @[Modules.scala 40:46:@4371.4]
  wire [5:0] _T_58014; // @[Modules.scala 43:37:@4377.4]
  wire [4:0] _T_58015; // @[Modules.scala 43:37:@4378.4]
  wire [4:0] _T_58016; // @[Modules.scala 43:37:@4379.4]
  wire [5:0] _T_58017; // @[Modules.scala 43:47:@4380.4]
  wire [4:0] _T_58018; // @[Modules.scala 43:47:@4381.4]
  wire [4:0] _T_58019; // @[Modules.scala 43:47:@4382.4]
  wire [5:0] _T_58024; // @[Modules.scala 43:47:@4387.4]
  wire [4:0] _T_58025; // @[Modules.scala 43:47:@4388.4]
  wire [4:0] _T_58026; // @[Modules.scala 43:47:@4389.4]
  wire [5:0] _T_58031; // @[Modules.scala 43:47:@4394.4]
  wire [4:0] _T_58032; // @[Modules.scala 43:47:@4395.4]
  wire [4:0] _T_58033; // @[Modules.scala 43:47:@4396.4]
  wire [5:0] _T_58038; // @[Modules.scala 43:47:@4401.4]
  wire [4:0] _T_58039; // @[Modules.scala 43:47:@4402.4]
  wire [4:0] _T_58040; // @[Modules.scala 43:47:@4403.4]
  wire [5:0] _T_58041; // @[Modules.scala 37:46:@4405.4]
  wire [4:0] _T_58042; // @[Modules.scala 37:46:@4406.4]
  wire [4:0] _T_58043; // @[Modules.scala 37:46:@4407.4]
  wire [5:0] _T_58048; // @[Modules.scala 43:47:@4412.4]
  wire [4:0] _T_58049; // @[Modules.scala 43:47:@4413.4]
  wire [4:0] _T_58050; // @[Modules.scala 43:47:@4414.4]
  wire [5:0] _T_58051; // @[Modules.scala 37:46:@4416.4]
  wire [4:0] _T_58052; // @[Modules.scala 37:46:@4417.4]
  wire [4:0] _T_58053; // @[Modules.scala 37:46:@4418.4]
  wire [5:0] _T_58093; // @[Modules.scala 46:47:@4458.4]
  wire [4:0] _T_58094; // @[Modules.scala 46:47:@4459.4]
  wire [4:0] _T_58095; // @[Modules.scala 46:47:@4460.4]
  wire [5:0] _T_58103; // @[Modules.scala 37:46:@4469.4]
  wire [4:0] _T_58104; // @[Modules.scala 37:46:@4470.4]
  wire [4:0] _T_58105; // @[Modules.scala 37:46:@4471.4]
  wire [5:0] _T_58124; // @[Modules.scala 43:47:@4490.4]
  wire [4:0] _T_58125; // @[Modules.scala 43:47:@4491.4]
  wire [4:0] _T_58126; // @[Modules.scala 43:47:@4492.4]
  wire [5:0] _T_58127; // @[Modules.scala 37:46:@4494.4]
  wire [4:0] _T_58128; // @[Modules.scala 37:46:@4495.4]
  wire [4:0] _T_58129; // @[Modules.scala 37:46:@4496.4]
  wire [5:0] _T_58130; // @[Modules.scala 37:46:@4498.4]
  wire [4:0] _T_58131; // @[Modules.scala 37:46:@4499.4]
  wire [4:0] _T_58132; // @[Modules.scala 37:46:@4500.4]
  wire [5:0] _T_58137; // @[Modules.scala 43:47:@4505.4]
  wire [4:0] _T_58138; // @[Modules.scala 43:47:@4506.4]
  wire [4:0] _T_58139; // @[Modules.scala 43:47:@4507.4]
  wire [5:0] _T_58161; // @[Modules.scala 40:46:@4530.4]
  wire [4:0] _T_58162; // @[Modules.scala 40:46:@4531.4]
  wire [4:0] _T_58163; // @[Modules.scala 40:46:@4532.4]
  wire [5:0] _T_58165; // @[Modules.scala 46:37:@4534.4]
  wire [4:0] _T_58166; // @[Modules.scala 46:37:@4535.4]
  wire [4:0] _T_58167; // @[Modules.scala 46:37:@4536.4]
  wire [5:0] _T_58168; // @[Modules.scala 46:47:@4537.4]
  wire [4:0] _T_58169; // @[Modules.scala 46:47:@4538.4]
  wire [4:0] _T_58170; // @[Modules.scala 46:47:@4539.4]
  wire [5:0] _T_58178; // @[Modules.scala 37:46:@4548.4]
  wire [4:0] _T_58179; // @[Modules.scala 37:46:@4549.4]
  wire [4:0] _T_58180; // @[Modules.scala 37:46:@4550.4]
  wire [5:0] _T_58206; // @[Modules.scala 43:47:@4576.4]
  wire [4:0] _T_58207; // @[Modules.scala 43:47:@4577.4]
  wire [4:0] _T_58208; // @[Modules.scala 43:47:@4578.4]
  wire [5:0] _T_58209; // @[Modules.scala 37:46:@4580.4]
  wire [4:0] _T_58210; // @[Modules.scala 37:46:@4581.4]
  wire [4:0] _T_58211; // @[Modules.scala 37:46:@4582.4]
  wire [5:0] _T_58212; // @[Modules.scala 37:46:@4584.4]
  wire [4:0] _T_58213; // @[Modules.scala 37:46:@4585.4]
  wire [4:0] _T_58214; // @[Modules.scala 37:46:@4586.4]
  wire [5:0] _T_58219; // @[Modules.scala 43:47:@4591.4]
  wire [4:0] _T_58220; // @[Modules.scala 43:47:@4592.4]
  wire [4:0] _T_58221; // @[Modules.scala 43:47:@4593.4]
  wire [5:0] _T_58226; // @[Modules.scala 43:47:@4598.4]
  wire [4:0] _T_58227; // @[Modules.scala 43:47:@4599.4]
  wire [4:0] _T_58228; // @[Modules.scala 43:47:@4600.4]
  wire [5:0] _T_58257; // @[Modules.scala 37:46:@4630.4]
  wire [4:0] _T_58258; // @[Modules.scala 37:46:@4631.4]
  wire [4:0] _T_58259; // @[Modules.scala 37:46:@4632.4]
  wire [5:0] _T_58260; // @[Modules.scala 40:46:@4634.4]
  wire [4:0] _T_58261; // @[Modules.scala 40:46:@4635.4]
  wire [4:0] _T_58262; // @[Modules.scala 40:46:@4636.4]
  wire [5:0] _T_58288; // @[Modules.scala 43:47:@4662.4]
  wire [4:0] _T_58289; // @[Modules.scala 43:47:@4663.4]
  wire [4:0] _T_58290; // @[Modules.scala 43:47:@4664.4]
  wire [5:0] _T_58291; // @[Modules.scala 37:46:@4666.4]
  wire [4:0] _T_58292; // @[Modules.scala 37:46:@4667.4]
  wire [4:0] _T_58293; // @[Modules.scala 37:46:@4668.4]
  wire [5:0] _T_58294; // @[Modules.scala 37:46:@4670.4]
  wire [4:0] _T_58295; // @[Modules.scala 37:46:@4671.4]
  wire [4:0] _T_58296; // @[Modules.scala 37:46:@4672.4]
  wire [5:0] _T_58318; // @[Modules.scala 40:46:@4695.4]
  wire [4:0] _T_58319; // @[Modules.scala 40:46:@4696.4]
  wire [4:0] _T_58320; // @[Modules.scala 40:46:@4697.4]
  wire [5:0] _T_58322; // @[Modules.scala 46:37:@4699.4]
  wire [4:0] _T_58323; // @[Modules.scala 46:37:@4700.4]
  wire [4:0] _T_58324; // @[Modules.scala 46:37:@4701.4]
  wire [5:0] _T_58325; // @[Modules.scala 46:47:@4702.4]
  wire [4:0] _T_58326; // @[Modules.scala 46:47:@4703.4]
  wire [4:0] _T_58327; // @[Modules.scala 46:47:@4704.4]
  wire [5:0] _T_58331; // @[Modules.scala 37:46:@4710.4]
  wire [4:0] _T_58332; // @[Modules.scala 37:46:@4711.4]
  wire [4:0] _T_58333; // @[Modules.scala 37:46:@4712.4]
  wire [5:0] _T_58334; // @[Modules.scala 40:46:@4714.4]
  wire [4:0] _T_58335; // @[Modules.scala 40:46:@4715.4]
  wire [4:0] _T_58336; // @[Modules.scala 40:46:@4716.4]
  wire [5:0] _T_58341; // @[Modules.scala 46:47:@4721.4]
  wire [4:0] _T_58342; // @[Modules.scala 46:47:@4722.4]
  wire [4:0] _T_58343; // @[Modules.scala 46:47:@4723.4]
  wire [5:0] _T_58352; // @[Modules.scala 46:37:@4732.4]
  wire [4:0] _T_58353; // @[Modules.scala 46:37:@4733.4]
  wire [4:0] _T_58354; // @[Modules.scala 46:37:@4734.4]
  wire [5:0] _T_58355; // @[Modules.scala 46:47:@4735.4]
  wire [4:0] _T_58356; // @[Modules.scala 46:47:@4736.4]
  wire [4:0] _T_58357; // @[Modules.scala 46:47:@4737.4]
  wire [5:0] _T_58362; // @[Modules.scala 43:47:@4742.4]
  wire [4:0] _T_58363; // @[Modules.scala 43:47:@4743.4]
  wire [4:0] _T_58364; // @[Modules.scala 43:47:@4744.4]
  wire [5:0] _T_58365; // @[Modules.scala 37:46:@4746.4]
  wire [4:0] _T_58366; // @[Modules.scala 37:46:@4747.4]
  wire [4:0] _T_58367; // @[Modules.scala 37:46:@4748.4]
  wire [5:0] _T_58368; // @[Modules.scala 37:46:@4750.4]
  wire [4:0] _T_58369; // @[Modules.scala 37:46:@4751.4]
  wire [4:0] _T_58370; // @[Modules.scala 37:46:@4752.4]
  wire [5:0] _T_58401; // @[Modules.scala 46:37:@4788.4]
  wire [4:0] _T_58402; // @[Modules.scala 46:37:@4789.4]
  wire [4:0] _T_58403; // @[Modules.scala 46:37:@4790.4]
  wire [5:0] _T_58404; // @[Modules.scala 46:47:@4791.4]
  wire [4:0] _T_58405; // @[Modules.scala 46:47:@4792.4]
  wire [4:0] _T_58406; // @[Modules.scala 46:47:@4793.4]
  wire [5:0] _T_58408; // @[Modules.scala 46:37:@4795.4]
  wire [4:0] _T_58409; // @[Modules.scala 46:37:@4796.4]
  wire [4:0] _T_58410; // @[Modules.scala 46:37:@4797.4]
  wire [5:0] _T_58411; // @[Modules.scala 46:47:@4798.4]
  wire [4:0] _T_58412; // @[Modules.scala 46:47:@4799.4]
  wire [4:0] _T_58413; // @[Modules.scala 46:47:@4800.4]
  wire [5:0] _T_58415; // @[Modules.scala 46:37:@4802.4]
  wire [4:0] _T_58416; // @[Modules.scala 46:37:@4803.4]
  wire [4:0] _T_58417; // @[Modules.scala 46:37:@4804.4]
  wire [5:0] _T_58418; // @[Modules.scala 46:47:@4805.4]
  wire [4:0] _T_58419; // @[Modules.scala 46:47:@4806.4]
  wire [4:0] _T_58420; // @[Modules.scala 46:47:@4807.4]
  wire [5:0] _T_58422; // @[Modules.scala 46:37:@4809.4]
  wire [4:0] _T_58423; // @[Modules.scala 46:37:@4810.4]
  wire [4:0] _T_58424; // @[Modules.scala 46:37:@4811.4]
  wire [5:0] _T_58425; // @[Modules.scala 46:47:@4812.4]
  wire [4:0] _T_58426; // @[Modules.scala 46:47:@4813.4]
  wire [4:0] _T_58427; // @[Modules.scala 46:47:@4814.4]
  wire [5:0] _T_58429; // @[Modules.scala 43:37:@4816.4]
  wire [4:0] _T_58430; // @[Modules.scala 43:37:@4817.4]
  wire [4:0] _T_58431; // @[Modules.scala 43:37:@4818.4]
  wire [5:0] _T_58432; // @[Modules.scala 43:47:@4819.4]
  wire [4:0] _T_58433; // @[Modules.scala 43:47:@4820.4]
  wire [4:0] _T_58434; // @[Modules.scala 43:47:@4821.4]
  wire [5:0] _T_58435; // @[Modules.scala 37:46:@4823.4]
  wire [4:0] _T_58436; // @[Modules.scala 37:46:@4824.4]
  wire [4:0] _T_58437; // @[Modules.scala 37:46:@4825.4]
  wire [5:0] _T_58442; // @[Modules.scala 46:47:@4830.4]
  wire [4:0] _T_58443; // @[Modules.scala 46:47:@4831.4]
  wire [4:0] _T_58444; // @[Modules.scala 46:47:@4832.4]
  wire [5:0] _T_58460; // @[Modules.scala 43:37:@4848.4]
  wire [4:0] _T_58461; // @[Modules.scala 43:37:@4849.4]
  wire [4:0] _T_58462; // @[Modules.scala 43:37:@4850.4]
  wire [5:0] _T_58463; // @[Modules.scala 43:47:@4851.4]
  wire [4:0] _T_58464; // @[Modules.scala 43:47:@4852.4]
  wire [4:0] _T_58465; // @[Modules.scala 43:47:@4853.4]
  wire [5:0] _T_58479; // @[Modules.scala 46:37:@4871.4]
  wire [4:0] _T_58480; // @[Modules.scala 46:37:@4872.4]
  wire [4:0] _T_58481; // @[Modules.scala 46:37:@4873.4]
  wire [5:0] _T_58482; // @[Modules.scala 46:47:@4874.4]
  wire [4:0] _T_58483; // @[Modules.scala 46:47:@4875.4]
  wire [4:0] _T_58484; // @[Modules.scala 46:47:@4876.4]
  wire [5:0] _T_58486; // @[Modules.scala 46:37:@4878.4]
  wire [4:0] _T_58487; // @[Modules.scala 46:37:@4879.4]
  wire [4:0] _T_58488; // @[Modules.scala 46:37:@4880.4]
  wire [5:0] _T_58489; // @[Modules.scala 46:47:@4881.4]
  wire [4:0] _T_58490; // @[Modules.scala 46:47:@4882.4]
  wire [4:0] _T_58491; // @[Modules.scala 46:47:@4883.4]
  wire [5:0] _T_58493; // @[Modules.scala 46:37:@4885.4]
  wire [4:0] _T_58494; // @[Modules.scala 46:37:@4886.4]
  wire [4:0] _T_58495; // @[Modules.scala 46:37:@4887.4]
  wire [5:0] _T_58496; // @[Modules.scala 46:47:@4888.4]
  wire [4:0] _T_58497; // @[Modules.scala 46:47:@4889.4]
  wire [4:0] _T_58498; // @[Modules.scala 46:47:@4890.4]
  wire [5:0] _T_58516; // @[Modules.scala 46:47:@4910.4]
  wire [4:0] _T_58517; // @[Modules.scala 46:47:@4911.4]
  wire [4:0] _T_58518; // @[Modules.scala 46:47:@4912.4]
  wire [5:0] _T_58519; // @[Modules.scala 37:46:@4914.4]
  wire [4:0] _T_58520; // @[Modules.scala 37:46:@4915.4]
  wire [4:0] _T_58521; // @[Modules.scala 37:46:@4916.4]
  wire [5:0] _T_58530; // @[Modules.scala 43:37:@4925.4]
  wire [4:0] _T_58531; // @[Modules.scala 43:37:@4926.4]
  wire [4:0] _T_58532; // @[Modules.scala 43:37:@4927.4]
  wire [5:0] _T_58533; // @[Modules.scala 43:47:@4928.4]
  wire [4:0] _T_58534; // @[Modules.scala 43:47:@4929.4]
  wire [4:0] _T_58535; // @[Modules.scala 43:47:@4930.4]
  wire [5:0] _T_58545; // @[Modules.scala 40:46:@4944.4]
  wire [4:0] _T_58546; // @[Modules.scala 40:46:@4945.4]
  wire [4:0] _T_58547; // @[Modules.scala 40:46:@4946.4]
  wire [5:0] _T_58549; // @[Modules.scala 46:37:@4948.4]
  wire [4:0] _T_58550; // @[Modules.scala 46:37:@4949.4]
  wire [4:0] _T_58551; // @[Modules.scala 46:37:@4950.4]
  wire [5:0] _T_58552; // @[Modules.scala 46:47:@4951.4]
  wire [4:0] _T_58553; // @[Modules.scala 46:47:@4952.4]
  wire [4:0] _T_58554; // @[Modules.scala 46:47:@4953.4]
  wire [5:0] _T_58555; // @[Modules.scala 40:46:@4955.4]
  wire [4:0] _T_58556; // @[Modules.scala 40:46:@4956.4]
  wire [4:0] _T_58557; // @[Modules.scala 40:46:@4957.4]
  wire [5:0] _T_58559; // @[Modules.scala 46:37:@4959.4]
  wire [4:0] _T_58560; // @[Modules.scala 46:37:@4960.4]
  wire [4:0] _T_58561; // @[Modules.scala 46:37:@4961.4]
  wire [5:0] _T_58562; // @[Modules.scala 46:47:@4962.4]
  wire [4:0] _T_58563; // @[Modules.scala 46:47:@4963.4]
  wire [4:0] _T_58564; // @[Modules.scala 46:47:@4964.4]
  wire [5:0] _T_58578; // @[Modules.scala 46:47:@4981.4]
  wire [4:0] _T_58579; // @[Modules.scala 46:47:@4982.4]
  wire [4:0] _T_58580; // @[Modules.scala 46:47:@4983.4]
  wire [5:0] _T_58588; // @[Modules.scala 40:46:@4992.4]
  wire [4:0] _T_58589; // @[Modules.scala 40:46:@4993.4]
  wire [4:0] _T_58590; // @[Modules.scala 40:46:@4994.4]
  wire [5:0] _T_58599; // @[Modules.scala 46:37:@5003.4]
  wire [4:0] _T_58600; // @[Modules.scala 46:37:@5004.4]
  wire [4:0] _T_58601; // @[Modules.scala 46:37:@5005.4]
  wire [5:0] _T_58602; // @[Modules.scala 46:47:@5006.4]
  wire [4:0] _T_58603; // @[Modules.scala 46:47:@5007.4]
  wire [4:0] _T_58604; // @[Modules.scala 46:47:@5008.4]
  wire [5:0] _T_58612; // @[Modules.scala 46:37:@5018.4]
  wire [4:0] _T_58613; // @[Modules.scala 46:37:@5019.4]
  wire [4:0] _T_58614; // @[Modules.scala 46:37:@5020.4]
  wire [5:0] _T_58615; // @[Modules.scala 46:47:@5021.4]
  wire [4:0] _T_58616; // @[Modules.scala 46:47:@5022.4]
  wire [4:0] _T_58617; // @[Modules.scala 46:47:@5023.4]
  wire [5:0] _T_58619; // @[Modules.scala 46:37:@5025.4]
  wire [4:0] _T_58620; // @[Modules.scala 46:37:@5026.4]
  wire [4:0] _T_58621; // @[Modules.scala 46:37:@5027.4]
  wire [5:0] _T_58622; // @[Modules.scala 46:47:@5028.4]
  wire [4:0] _T_58623; // @[Modules.scala 46:47:@5029.4]
  wire [4:0] _T_58624; // @[Modules.scala 46:47:@5030.4]
  wire [5:0] _T_58626; // @[Modules.scala 46:37:@5032.4]
  wire [4:0] _T_58627; // @[Modules.scala 46:37:@5033.4]
  wire [4:0] _T_58628; // @[Modules.scala 46:37:@5034.4]
  wire [5:0] _T_58629; // @[Modules.scala 46:47:@5035.4]
  wire [4:0] _T_58630; // @[Modules.scala 46:47:@5036.4]
  wire [4:0] _T_58631; // @[Modules.scala 46:47:@5037.4]
  wire [5:0] _T_58633; // @[Modules.scala 43:37:@5039.4]
  wire [4:0] _T_58634; // @[Modules.scala 43:37:@5040.4]
  wire [4:0] _T_58635; // @[Modules.scala 43:37:@5041.4]
  wire [5:0] _T_58636; // @[Modules.scala 43:47:@5042.4]
  wire [4:0] _T_58637; // @[Modules.scala 43:47:@5043.4]
  wire [4:0] _T_58638; // @[Modules.scala 43:47:@5044.4]
  wire [5:0] _T_58639; // @[Modules.scala 37:46:@5046.4]
  wire [4:0] _T_58640; // @[Modules.scala 37:46:@5047.4]
  wire [4:0] _T_58641; // @[Modules.scala 37:46:@5048.4]
  wire [5:0] _T_58642; // @[Modules.scala 37:46:@5050.4]
  wire [4:0] _T_58643; // @[Modules.scala 37:46:@5051.4]
  wire [4:0] _T_58644; // @[Modules.scala 37:46:@5052.4]
  wire [5:0] _T_58645; // @[Modules.scala 40:46:@5054.4]
  wire [4:0] _T_58646; // @[Modules.scala 40:46:@5055.4]
  wire [4:0] _T_58647; // @[Modules.scala 40:46:@5056.4]
  wire [5:0] _T_58656; // @[Modules.scala 43:37:@5065.4]
  wire [4:0] _T_58657; // @[Modules.scala 43:37:@5066.4]
  wire [4:0] _T_58658; // @[Modules.scala 43:37:@5067.4]
  wire [5:0] _T_58659; // @[Modules.scala 43:47:@5068.4]
  wire [4:0] _T_58660; // @[Modules.scala 43:47:@5069.4]
  wire [4:0] _T_58661; // @[Modules.scala 43:47:@5070.4]
  wire [5:0] _T_58662; // @[Modules.scala 37:46:@5072.4]
  wire [4:0] _T_58663; // @[Modules.scala 37:46:@5073.4]
  wire [4:0] _T_58664; // @[Modules.scala 37:46:@5074.4]
  wire [5:0] _T_58669; // @[Modules.scala 46:47:@5079.4]
  wire [4:0] _T_58670; // @[Modules.scala 46:47:@5080.4]
  wire [4:0] _T_58671; // @[Modules.scala 46:47:@5081.4]
  wire [5:0] _T_58673; // @[Modules.scala 46:37:@5083.4]
  wire [4:0] _T_58674; // @[Modules.scala 46:37:@5084.4]
  wire [4:0] _T_58675; // @[Modules.scala 46:37:@5085.4]
  wire [5:0] _T_58676; // @[Modules.scala 46:47:@5086.4]
  wire [4:0] _T_58677; // @[Modules.scala 46:47:@5087.4]
  wire [4:0] _T_58678; // @[Modules.scala 46:47:@5088.4]
  wire [5:0] _T_58680; // @[Modules.scala 43:37:@5090.4]
  wire [4:0] _T_58681; // @[Modules.scala 43:37:@5091.4]
  wire [4:0] _T_58682; // @[Modules.scala 43:37:@5092.4]
  wire [5:0] _T_58683; // @[Modules.scala 43:47:@5093.4]
  wire [4:0] _T_58684; // @[Modules.scala 43:47:@5094.4]
  wire [4:0] _T_58685; // @[Modules.scala 43:47:@5095.4]
  wire [5:0] _T_58686; // @[Modules.scala 40:46:@5097.4]
  wire [4:0] _T_58687; // @[Modules.scala 40:46:@5098.4]
  wire [4:0] _T_58688; // @[Modules.scala 40:46:@5099.4]
  wire [5:0] _T_58690; // @[Modules.scala 46:37:@5101.4]
  wire [4:0] _T_58691; // @[Modules.scala 46:37:@5102.4]
  wire [4:0] _T_58692; // @[Modules.scala 46:37:@5103.4]
  wire [5:0] _T_58693; // @[Modules.scala 46:47:@5104.4]
  wire [4:0] _T_58694; // @[Modules.scala 46:47:@5105.4]
  wire [4:0] _T_58695; // @[Modules.scala 46:47:@5106.4]
  wire [5:0] _T_58697; // @[Modules.scala 46:37:@5108.4]
  wire [4:0] _T_58698; // @[Modules.scala 46:37:@5109.4]
  wire [4:0] _T_58699; // @[Modules.scala 46:37:@5110.4]
  wire [5:0] _T_58700; // @[Modules.scala 46:47:@5111.4]
  wire [4:0] _T_58701; // @[Modules.scala 46:47:@5112.4]
  wire [4:0] _T_58702; // @[Modules.scala 46:47:@5113.4]
  wire [5:0] _T_58704; // @[Modules.scala 46:37:@5115.4]
  wire [4:0] _T_58705; // @[Modules.scala 46:37:@5116.4]
  wire [4:0] _T_58706; // @[Modules.scala 46:37:@5117.4]
  wire [5:0] _T_58707; // @[Modules.scala 46:47:@5118.4]
  wire [4:0] _T_58708; // @[Modules.scala 46:47:@5119.4]
  wire [4:0] _T_58709; // @[Modules.scala 46:47:@5120.4]
  wire [5:0] _T_58711; // @[Modules.scala 43:37:@5122.4]
  wire [4:0] _T_58712; // @[Modules.scala 43:37:@5123.4]
  wire [4:0] _T_58713; // @[Modules.scala 43:37:@5124.4]
  wire [5:0] _T_58714; // @[Modules.scala 43:47:@5125.4]
  wire [4:0] _T_58715; // @[Modules.scala 43:47:@5126.4]
  wire [4:0] _T_58716; // @[Modules.scala 43:47:@5127.4]
  wire [5:0] _T_58717; // @[Modules.scala 37:46:@5129.4]
  wire [4:0] _T_58718; // @[Modules.scala 37:46:@5130.4]
  wire [4:0] _T_58719; // @[Modules.scala 37:46:@5131.4]
  wire [5:0] _T_58720; // @[Modules.scala 37:46:@5133.4]
  wire [4:0] _T_58721; // @[Modules.scala 37:46:@5134.4]
  wire [4:0] _T_58722; // @[Modules.scala 37:46:@5135.4]
  wire [5:0] _T_58723; // @[Modules.scala 40:46:@5137.4]
  wire [4:0] _T_58724; // @[Modules.scala 40:46:@5138.4]
  wire [4:0] _T_58725; // @[Modules.scala 40:46:@5139.4]
  wire [5:0] _T_58737; // @[Modules.scala 43:47:@5151.4]
  wire [4:0] _T_58738; // @[Modules.scala 43:47:@5152.4]
  wire [4:0] _T_58739; // @[Modules.scala 43:47:@5153.4]
  wire [5:0] _T_58740; // @[Modules.scala 37:46:@5155.4]
  wire [4:0] _T_58741; // @[Modules.scala 37:46:@5156.4]
  wire [4:0] _T_58742; // @[Modules.scala 37:46:@5157.4]
  wire [5:0] _T_58754; // @[Modules.scala 46:37:@5170.4]
  wire [4:0] _T_58755; // @[Modules.scala 46:37:@5171.4]
  wire [4:0] _T_58756; // @[Modules.scala 46:37:@5172.4]
  wire [5:0] _T_58757; // @[Modules.scala 46:47:@5173.4]
  wire [4:0] _T_58758; // @[Modules.scala 46:47:@5174.4]
  wire [4:0] _T_58759; // @[Modules.scala 46:47:@5175.4]
  wire [5:0] _T_58761; // @[Modules.scala 46:37:@5177.4]
  wire [4:0] _T_58762; // @[Modules.scala 46:37:@5178.4]
  wire [4:0] _T_58763; // @[Modules.scala 46:37:@5179.4]
  wire [5:0] _T_58764; // @[Modules.scala 46:47:@5180.4]
  wire [4:0] _T_58765; // @[Modules.scala 46:47:@5181.4]
  wire [4:0] _T_58766; // @[Modules.scala 46:47:@5182.4]
  wire [5:0] _T_58771; // @[Modules.scala 46:47:@5187.4]
  wire [4:0] _T_58772; // @[Modules.scala 46:47:@5188.4]
  wire [4:0] _T_58773; // @[Modules.scala 46:47:@5189.4]
  wire [5:0] _T_58775; // @[Modules.scala 46:37:@5191.4]
  wire [4:0] _T_58776; // @[Modules.scala 46:37:@5192.4]
  wire [4:0] _T_58777; // @[Modules.scala 46:37:@5193.4]
  wire [5:0] _T_58778; // @[Modules.scala 46:47:@5194.4]
  wire [4:0] _T_58779; // @[Modules.scala 46:47:@5195.4]
  wire [4:0] _T_58780; // @[Modules.scala 46:47:@5196.4]
  wire [5:0] _T_58782; // @[Modules.scala 46:37:@5198.4]
  wire [4:0] _T_58783; // @[Modules.scala 46:37:@5199.4]
  wire [4:0] _T_58784; // @[Modules.scala 46:37:@5200.4]
  wire [5:0] _T_58785; // @[Modules.scala 46:47:@5201.4]
  wire [4:0] _T_58786; // @[Modules.scala 46:47:@5202.4]
  wire [4:0] _T_58787; // @[Modules.scala 46:47:@5203.4]
  wire [5:0] _T_58788; // @[Modules.scala 37:46:@5205.4]
  wire [4:0] _T_58789; // @[Modules.scala 37:46:@5206.4]
  wire [4:0] _T_58790; // @[Modules.scala 37:46:@5207.4]
  wire [5:0] _T_58791; // @[Modules.scala 37:46:@5209.4]
  wire [4:0] _T_58792; // @[Modules.scala 37:46:@5210.4]
  wire [4:0] _T_58793; // @[Modules.scala 37:46:@5211.4]
  wire [5:0] _T_58815; // @[Modules.scala 43:47:@5234.4]
  wire [4:0] _T_58816; // @[Modules.scala 43:47:@5235.4]
  wire [4:0] _T_58817; // @[Modules.scala 43:47:@5236.4]
  wire [5:0] _T_58818; // @[Modules.scala 37:46:@5238.4]
  wire [4:0] _T_58819; // @[Modules.scala 37:46:@5239.4]
  wire [4:0] _T_58820; // @[Modules.scala 37:46:@5240.4]
  wire [5:0] _T_58821; // @[Modules.scala 40:46:@5242.4]
  wire [4:0] _T_58822; // @[Modules.scala 40:46:@5243.4]
  wire [4:0] _T_58823; // @[Modules.scala 40:46:@5244.4]
  wire [5:0] _T_58824; // @[Modules.scala 37:46:@5246.4]
  wire [4:0] _T_58825; // @[Modules.scala 37:46:@5247.4]
  wire [4:0] _T_58826; // @[Modules.scala 37:46:@5248.4]
  wire [5:0] _T_58828; // @[Modules.scala 46:37:@5250.4]
  wire [4:0] _T_58829; // @[Modules.scala 46:37:@5251.4]
  wire [4:0] _T_58830; // @[Modules.scala 46:37:@5252.4]
  wire [5:0] _T_58831; // @[Modules.scala 46:47:@5253.4]
  wire [4:0] _T_58832; // @[Modules.scala 46:47:@5254.4]
  wire [4:0] _T_58833; // @[Modules.scala 46:47:@5255.4]
  wire [5:0] _T_58838; // @[Modules.scala 46:37:@5261.4]
  wire [4:0] _T_58839; // @[Modules.scala 46:37:@5262.4]
  wire [4:0] _T_58840; // @[Modules.scala 46:37:@5263.4]
  wire [5:0] _T_58841; // @[Modules.scala 46:47:@5264.4]
  wire [4:0] _T_58842; // @[Modules.scala 46:47:@5265.4]
  wire [4:0] _T_58843; // @[Modules.scala 46:47:@5266.4]
  wire [5:0] _T_58845; // @[Modules.scala 46:37:@5268.4]
  wire [4:0] _T_58846; // @[Modules.scala 46:37:@5269.4]
  wire [4:0] _T_58847; // @[Modules.scala 46:37:@5270.4]
  wire [5:0] _T_58848; // @[Modules.scala 46:47:@5271.4]
  wire [4:0] _T_58849; // @[Modules.scala 46:47:@5272.4]
  wire [4:0] _T_58850; // @[Modules.scala 46:47:@5273.4]
  wire [5:0] _T_58851; // @[Modules.scala 37:46:@5275.4]
  wire [4:0] _T_58852; // @[Modules.scala 37:46:@5276.4]
  wire [4:0] _T_58853; // @[Modules.scala 37:46:@5277.4]
  wire [5:0] _T_58854; // @[Modules.scala 37:46:@5279.4]
  wire [4:0] _T_58855; // @[Modules.scala 37:46:@5280.4]
  wire [4:0] _T_58856; // @[Modules.scala 37:46:@5281.4]
  wire [5:0] _T_58857; // @[Modules.scala 37:46:@5283.4]
  wire [4:0] _T_58858; // @[Modules.scala 37:46:@5284.4]
  wire [4:0] _T_58859; // @[Modules.scala 37:46:@5285.4]
  wire [5:0] _T_58860; // @[Modules.scala 40:46:@5287.4]
  wire [4:0] _T_58861; // @[Modules.scala 40:46:@5288.4]
  wire [4:0] _T_58862; // @[Modules.scala 40:46:@5289.4]
  wire [5:0] _T_58864; // @[Modules.scala 46:37:@5291.4]
  wire [4:0] _T_58865; // @[Modules.scala 46:37:@5292.4]
  wire [4:0] _T_58866; // @[Modules.scala 46:37:@5293.4]
  wire [5:0] _T_58867; // @[Modules.scala 46:47:@5294.4]
  wire [4:0] _T_58868; // @[Modules.scala 46:47:@5295.4]
  wire [4:0] _T_58869; // @[Modules.scala 46:47:@5296.4]
  wire [5:0] _T_58877; // @[Modules.scala 37:46:@5305.4]
  wire [4:0] _T_58878; // @[Modules.scala 37:46:@5306.4]
  wire [4:0] _T_58879; // @[Modules.scala 37:46:@5307.4]
  wire [5:0] _T_58880; // @[Modules.scala 37:46:@5309.4]
  wire [4:0] _T_58881; // @[Modules.scala 37:46:@5310.4]
  wire [4:0] _T_58882; // @[Modules.scala 37:46:@5311.4]
  wire [5:0] _T_58883; // @[Modules.scala 37:46:@5313.4]
  wire [4:0] _T_58884; // @[Modules.scala 37:46:@5314.4]
  wire [4:0] _T_58885; // @[Modules.scala 37:46:@5315.4]
  wire [5:0] _T_58886; // @[Modules.scala 37:46:@5317.4]
  wire [4:0] _T_58887; // @[Modules.scala 37:46:@5318.4]
  wire [4:0] _T_58888; // @[Modules.scala 37:46:@5319.4]
  wire [5:0] _T_58889; // @[Modules.scala 37:46:@5321.4]
  wire [4:0] _T_58890; // @[Modules.scala 37:46:@5322.4]
  wire [4:0] _T_58891; // @[Modules.scala 37:46:@5323.4]
  wire [5:0] _T_58892; // @[Modules.scala 37:46:@5325.4]
  wire [4:0] _T_58893; // @[Modules.scala 37:46:@5326.4]
  wire [4:0] _T_58894; // @[Modules.scala 37:46:@5327.4]
  wire [5:0] _T_58895; // @[Modules.scala 37:46:@5329.4]
  wire [4:0] _T_58896; // @[Modules.scala 37:46:@5330.4]
  wire [4:0] _T_58897; // @[Modules.scala 37:46:@5331.4]
  wire [5:0] _T_58902; // @[Modules.scala 43:47:@5336.4]
  wire [4:0] _T_58903; // @[Modules.scala 43:47:@5337.4]
  wire [4:0] _T_58904; // @[Modules.scala 43:47:@5338.4]
  wire [5:0] _T_58905; // @[Modules.scala 37:46:@5340.4]
  wire [4:0] _T_58906; // @[Modules.scala 37:46:@5341.4]
  wire [4:0] _T_58907; // @[Modules.scala 37:46:@5342.4]
  wire [5:0] _T_58908; // @[Modules.scala 37:46:@5344.4]
  wire [4:0] _T_58909; // @[Modules.scala 37:46:@5345.4]
  wire [4:0] _T_58910; // @[Modules.scala 37:46:@5346.4]
  wire [5:0] _T_58914; // @[Modules.scala 40:46:@5352.4]
  wire [4:0] _T_58915; // @[Modules.scala 40:46:@5353.4]
  wire [4:0] _T_58916; // @[Modules.scala 40:46:@5354.4]
  wire [5:0] _T_58918; // @[Modules.scala 46:37:@5356.4]
  wire [4:0] _T_58919; // @[Modules.scala 46:37:@5357.4]
  wire [4:0] _T_58920; // @[Modules.scala 46:37:@5358.4]
  wire [5:0] _T_58921; // @[Modules.scala 46:47:@5359.4]
  wire [4:0] _T_58922; // @[Modules.scala 46:47:@5360.4]
  wire [4:0] _T_58923; // @[Modules.scala 46:47:@5361.4]
  wire [5:0] _T_58928; // @[Modules.scala 46:47:@5366.4]
  wire [4:0] _T_58929; // @[Modules.scala 46:47:@5367.4]
  wire [4:0] _T_58930; // @[Modules.scala 46:47:@5368.4]
  wire [5:0] _T_58935; // @[Modules.scala 43:47:@5373.4]
  wire [4:0] _T_58936; // @[Modules.scala 43:47:@5374.4]
  wire [4:0] _T_58937; // @[Modules.scala 43:47:@5375.4]
  wire [5:0] _T_58938; // @[Modules.scala 37:46:@5377.4]
  wire [4:0] _T_58939; // @[Modules.scala 37:46:@5378.4]
  wire [4:0] _T_58940; // @[Modules.scala 37:46:@5379.4]
  wire [5:0] _T_58941; // @[Modules.scala 37:46:@5381.4]
  wire [4:0] _T_58942; // @[Modules.scala 37:46:@5382.4]
  wire [4:0] _T_58943; // @[Modules.scala 37:46:@5383.4]
  wire [5:0] _T_58944; // @[Modules.scala 40:46:@5385.4]
  wire [4:0] _T_58945; // @[Modules.scala 40:46:@5386.4]
  wire [4:0] _T_58946; // @[Modules.scala 40:46:@5387.4]
  wire [5:0] _T_58947; // @[Modules.scala 37:46:@5389.4]
  wire [4:0] _T_58948; // @[Modules.scala 37:46:@5390.4]
  wire [4:0] _T_58949; // @[Modules.scala 37:46:@5391.4]
  wire [5:0] _T_58950; // @[Modules.scala 37:46:@5393.4]
  wire [4:0] _T_58951; // @[Modules.scala 37:46:@5394.4]
  wire [4:0] _T_58952; // @[Modules.scala 37:46:@5395.4]
  wire [5:0] _T_58953; // @[Modules.scala 37:46:@5397.4]
  wire [4:0] _T_58954; // @[Modules.scala 37:46:@5398.4]
  wire [4:0] _T_58955; // @[Modules.scala 37:46:@5399.4]
  wire [5:0] _T_58956; // @[Modules.scala 37:46:@5401.4]
  wire [4:0] _T_58957; // @[Modules.scala 37:46:@5402.4]
  wire [4:0] _T_58958; // @[Modules.scala 37:46:@5403.4]
  wire [5:0] _T_58959; // @[Modules.scala 40:46:@5405.4]
  wire [4:0] _T_58960; // @[Modules.scala 40:46:@5406.4]
  wire [4:0] _T_58961; // @[Modules.scala 40:46:@5407.4]
  wire [5:0] _T_58962; // @[Modules.scala 37:46:@5409.4]
  wire [4:0] _T_58963; // @[Modules.scala 37:46:@5410.4]
  wire [4:0] _T_58964; // @[Modules.scala 37:46:@5411.4]
  wire [5:0] _T_58968; // @[Modules.scala 40:46:@5417.4]
  wire [4:0] _T_58969; // @[Modules.scala 40:46:@5418.4]
  wire [4:0] _T_58970; // @[Modules.scala 40:46:@5419.4]
  wire [5:0] _T_58972; // @[Modules.scala 46:37:@5421.4]
  wire [4:0] _T_58973; // @[Modules.scala 46:37:@5422.4]
  wire [4:0] _T_58974; // @[Modules.scala 46:37:@5423.4]
  wire [5:0] _T_58975; // @[Modules.scala 46:47:@5424.4]
  wire [4:0] _T_58976; // @[Modules.scala 46:47:@5425.4]
  wire [4:0] _T_58977; // @[Modules.scala 46:47:@5426.4]
  wire [5:0] _T_58989; // @[Modules.scala 46:47:@5438.4]
  wire [4:0] _T_58990; // @[Modules.scala 46:47:@5439.4]
  wire [4:0] _T_58991; // @[Modules.scala 46:47:@5440.4]
  wire [5:0] _T_58992; // @[Modules.scala 37:46:@5442.4]
  wire [4:0] _T_58993; // @[Modules.scala 37:46:@5443.4]
  wire [4:0] _T_58994; // @[Modules.scala 37:46:@5444.4]
  wire [5:0] _T_58995; // @[Modules.scala 37:46:@5446.4]
  wire [4:0] _T_58996; // @[Modules.scala 37:46:@5447.4]
  wire [4:0] _T_58997; // @[Modules.scala 37:46:@5448.4]
  wire [5:0] _T_58998; // @[Modules.scala 40:46:@5450.4]
  wire [4:0] _T_58999; // @[Modules.scala 40:46:@5451.4]
  wire [4:0] _T_59000; // @[Modules.scala 40:46:@5452.4]
  wire [5:0] _T_59001; // @[Modules.scala 40:46:@5454.4]
  wire [4:0] _T_59002; // @[Modules.scala 40:46:@5455.4]
  wire [4:0] _T_59003; // @[Modules.scala 40:46:@5456.4]
  wire [5:0] _T_59004; // @[Modules.scala 37:46:@5458.4]
  wire [4:0] _T_59005; // @[Modules.scala 37:46:@5459.4]
  wire [4:0] _T_59006; // @[Modules.scala 37:46:@5460.4]
  wire [5:0] _T_59010; // @[Modules.scala 37:46:@5466.4]
  wire [4:0] _T_59011; // @[Modules.scala 37:46:@5467.4]
  wire [4:0] _T_59012; // @[Modules.scala 37:46:@5468.4]
  wire [5:0] _T_59034; // @[Modules.scala 46:37:@5492.4]
  wire [4:0] _T_59035; // @[Modules.scala 46:37:@5493.4]
  wire [4:0] _T_59036; // @[Modules.scala 46:37:@5494.4]
  wire [5:0] _T_59037; // @[Modules.scala 46:47:@5495.4]
  wire [4:0] _T_59038; // @[Modules.scala 46:47:@5496.4]
  wire [4:0] _T_59039; // @[Modules.scala 46:47:@5497.4]
  wire [5:0] _T_59051; // @[Modules.scala 46:47:@5509.4]
  wire [4:0] _T_59052; // @[Modules.scala 46:47:@5510.4]
  wire [4:0] _T_59053; // @[Modules.scala 46:47:@5511.4]
  wire [5:0] _T_59057; // @[Modules.scala 40:46:@5517.4]
  wire [4:0] _T_59058; // @[Modules.scala 40:46:@5518.4]
  wire [4:0] _T_59059; // @[Modules.scala 40:46:@5519.4]
  wire [5:0] _T_59067; // @[Modules.scala 37:46:@5528.4]
  wire [4:0] _T_59068; // @[Modules.scala 37:46:@5529.4]
  wire [4:0] _T_59069; // @[Modules.scala 37:46:@5530.4]
  wire [5:0] _T_59070; // @[Modules.scala 37:46:@5532.4]
  wire [4:0] _T_59071; // @[Modules.scala 37:46:@5533.4]
  wire [4:0] _T_59072; // @[Modules.scala 37:46:@5534.4]
  wire [5:0] _T_59073; // @[Modules.scala 37:46:@5536.4]
  wire [4:0] _T_59074; // @[Modules.scala 37:46:@5537.4]
  wire [4:0] _T_59075; // @[Modules.scala 37:46:@5538.4]
  wire [5:0] _T_59076; // @[Modules.scala 37:46:@5540.4]
  wire [4:0] _T_59077; // @[Modules.scala 37:46:@5541.4]
  wire [4:0] _T_59078; // @[Modules.scala 37:46:@5542.4]
  wire [5:0] _T_59079; // @[Modules.scala 37:46:@5544.4]
  wire [4:0] _T_59080; // @[Modules.scala 37:46:@5545.4]
  wire [4:0] _T_59081; // @[Modules.scala 37:46:@5546.4]
  wire [5:0] _T_59082; // @[Modules.scala 40:46:@5548.4]
  wire [4:0] _T_59083; // @[Modules.scala 40:46:@5549.4]
  wire [4:0] _T_59084; // @[Modules.scala 40:46:@5550.4]
  wire [5:0] _T_59085; // @[Modules.scala 37:46:@5552.4]
  wire [4:0] _T_59086; // @[Modules.scala 37:46:@5553.4]
  wire [4:0] _T_59087; // @[Modules.scala 37:46:@5554.4]
  wire [5:0] _T_59088; // @[Modules.scala 40:46:@5556.4]
  wire [4:0] _T_59089; // @[Modules.scala 40:46:@5557.4]
  wire [4:0] _T_59090; // @[Modules.scala 40:46:@5558.4]
  wire [5:0] _T_59092; // @[Modules.scala 46:37:@5560.4]
  wire [4:0] _T_59093; // @[Modules.scala 46:37:@5561.4]
  wire [4:0] _T_59094; // @[Modules.scala 46:37:@5562.4]
  wire [5:0] _T_59095; // @[Modules.scala 46:47:@5563.4]
  wire [4:0] _T_59096; // @[Modules.scala 46:47:@5564.4]
  wire [4:0] _T_59097; // @[Modules.scala 46:47:@5565.4]
  wire [5:0] _T_59098; // @[Modules.scala 37:46:@5567.4]
  wire [4:0] _T_59099; // @[Modules.scala 37:46:@5568.4]
  wire [4:0] _T_59100; // @[Modules.scala 37:46:@5569.4]
  wire [5:0] _T_59105; // @[Modules.scala 46:47:@5574.4]
  wire [4:0] _T_59106; // @[Modules.scala 46:47:@5575.4]
  wire [4:0] _T_59107; // @[Modules.scala 46:47:@5576.4]
  wire [5:0] _T_59111; // @[Modules.scala 37:46:@5582.4]
  wire [4:0] _T_59112; // @[Modules.scala 37:46:@5583.4]
  wire [4:0] _T_59113; // @[Modules.scala 37:46:@5584.4]
  wire [5:0] _T_59114; // @[Modules.scala 37:46:@5586.4]
  wire [4:0] _T_59115; // @[Modules.scala 37:46:@5587.4]
  wire [4:0] _T_59116; // @[Modules.scala 37:46:@5588.4]
  wire [5:0] _T_59117; // @[Modules.scala 37:46:@5590.4]
  wire [4:0] _T_59118; // @[Modules.scala 37:46:@5591.4]
  wire [4:0] _T_59119; // @[Modules.scala 37:46:@5592.4]
  wire [5:0] _T_59120; // @[Modules.scala 37:46:@5594.4]
  wire [4:0] _T_59121; // @[Modules.scala 37:46:@5595.4]
  wire [4:0] _T_59122; // @[Modules.scala 37:46:@5596.4]
  wire [5:0] _T_59123; // @[Modules.scala 37:46:@5598.4]
  wire [4:0] _T_59124; // @[Modules.scala 37:46:@5599.4]
  wire [4:0] _T_59125; // @[Modules.scala 37:46:@5600.4]
  wire [5:0] _T_59126; // @[Modules.scala 37:46:@5602.4]
  wire [4:0] _T_59127; // @[Modules.scala 37:46:@5603.4]
  wire [4:0] _T_59128; // @[Modules.scala 37:46:@5604.4]
  wire [5:0] _T_59136; // @[Modules.scala 37:46:@5613.4]
  wire [4:0] _T_59137; // @[Modules.scala 37:46:@5614.4]
  wire [4:0] _T_59138; // @[Modules.scala 37:46:@5615.4]
  wire [5:0] _T_59140; // @[Modules.scala 46:37:@5617.4]
  wire [4:0] _T_59141; // @[Modules.scala 46:37:@5618.4]
  wire [4:0] _T_59142; // @[Modules.scala 46:37:@5619.4]
  wire [5:0] _T_59143; // @[Modules.scala 46:47:@5620.4]
  wire [4:0] _T_59144; // @[Modules.scala 46:47:@5621.4]
  wire [4:0] _T_59145; // @[Modules.scala 46:47:@5622.4]
  wire [5:0] _T_59147; // @[Modules.scala 46:37:@5624.4]
  wire [4:0] _T_59148; // @[Modules.scala 46:37:@5625.4]
  wire [4:0] _T_59149; // @[Modules.scala 46:37:@5626.4]
  wire [5:0] _T_59150; // @[Modules.scala 46:47:@5627.4]
  wire [4:0] _T_59151; // @[Modules.scala 46:47:@5628.4]
  wire [4:0] _T_59152; // @[Modules.scala 46:47:@5629.4]
  wire [5:0] _T_59154; // @[Modules.scala 46:37:@5631.4]
  wire [4:0] _T_59155; // @[Modules.scala 46:37:@5632.4]
  wire [4:0] _T_59156; // @[Modules.scala 46:37:@5633.4]
  wire [5:0] _T_59157; // @[Modules.scala 46:47:@5634.4]
  wire [4:0] _T_59158; // @[Modules.scala 46:47:@5635.4]
  wire [4:0] _T_59159; // @[Modules.scala 46:47:@5636.4]
  wire [5:0] _T_59171; // @[Modules.scala 46:47:@5648.4]
  wire [4:0] _T_59172; // @[Modules.scala 46:47:@5649.4]
  wire [4:0] _T_59173; // @[Modules.scala 46:47:@5650.4]
  wire [5:0] _T_59174; // @[Modules.scala 37:46:@5652.4]
  wire [4:0] _T_59175; // @[Modules.scala 37:46:@5653.4]
  wire [4:0] _T_59176; // @[Modules.scala 37:46:@5654.4]
  wire [5:0] _T_59184; // @[Modules.scala 43:37:@5664.4]
  wire [4:0] _T_59185; // @[Modules.scala 43:37:@5665.4]
  wire [4:0] _T_59186; // @[Modules.scala 43:37:@5666.4]
  wire [5:0] _T_59187; // @[Modules.scala 43:47:@5667.4]
  wire [4:0] _T_59188; // @[Modules.scala 43:47:@5668.4]
  wire [4:0] _T_59189; // @[Modules.scala 43:47:@5669.4]
  wire [5:0] _T_59190; // @[Modules.scala 37:46:@5671.4]
  wire [4:0] _T_59191; // @[Modules.scala 37:46:@5672.4]
  wire [4:0] _T_59192; // @[Modules.scala 37:46:@5673.4]
  wire [5:0] _T_59193; // @[Modules.scala 37:46:@5675.4]
  wire [4:0] _T_59194; // @[Modules.scala 37:46:@5676.4]
  wire [4:0] _T_59195; // @[Modules.scala 37:46:@5677.4]
  wire [5:0] _T_59196; // @[Modules.scala 40:46:@5679.4]
  wire [4:0] _T_59197; // @[Modules.scala 40:46:@5680.4]
  wire [4:0] _T_59198; // @[Modules.scala 40:46:@5681.4]
  wire [5:0] _T_59199; // @[Modules.scala 40:46:@5683.4]
  wire [4:0] _T_59200; // @[Modules.scala 40:46:@5684.4]
  wire [4:0] _T_59201; // @[Modules.scala 40:46:@5685.4]
  wire [5:0] _T_59202; // @[Modules.scala 40:46:@5687.4]
  wire [4:0] _T_59203; // @[Modules.scala 40:46:@5688.4]
  wire [4:0] _T_59204; // @[Modules.scala 40:46:@5689.4]
  wire [5:0] _T_59206; // @[Modules.scala 46:37:@5691.4]
  wire [4:0] _T_59207; // @[Modules.scala 46:37:@5692.4]
  wire [4:0] _T_59208; // @[Modules.scala 46:37:@5693.4]
  wire [5:0] _T_59209; // @[Modules.scala 46:47:@5694.4]
  wire [4:0] _T_59210; // @[Modules.scala 46:47:@5695.4]
  wire [4:0] _T_59211; // @[Modules.scala 46:47:@5696.4]
  wire [5:0] _T_59213; // @[Modules.scala 43:37:@5698.4]
  wire [4:0] _T_59214; // @[Modules.scala 43:37:@5699.4]
  wire [4:0] _T_59215; // @[Modules.scala 43:37:@5700.4]
  wire [5:0] _T_59216; // @[Modules.scala 43:47:@5701.4]
  wire [4:0] _T_59217; // @[Modules.scala 43:47:@5702.4]
  wire [4:0] _T_59218; // @[Modules.scala 43:47:@5703.4]
  wire [5:0] _T_59219; // @[Modules.scala 40:46:@5705.4]
  wire [4:0] _T_59220; // @[Modules.scala 40:46:@5706.4]
  wire [4:0] _T_59221; // @[Modules.scala 40:46:@5707.4]
  wire [5:0] _T_59226; // @[Modules.scala 46:47:@5712.4]
  wire [4:0] _T_59227; // @[Modules.scala 46:47:@5713.4]
  wire [4:0] _T_59228; // @[Modules.scala 46:47:@5714.4]
  wire [5:0] _T_59229; // @[Modules.scala 37:46:@5716.4]
  wire [4:0] _T_59230; // @[Modules.scala 37:46:@5717.4]
  wire [4:0] _T_59231; // @[Modules.scala 37:46:@5718.4]
  wire [5:0] _T_59232; // @[Modules.scala 37:46:@5720.4]
  wire [4:0] _T_59233; // @[Modules.scala 37:46:@5721.4]
  wire [4:0] _T_59234; // @[Modules.scala 37:46:@5722.4]
  wire [5:0] _T_59242; // @[Modules.scala 46:37:@5732.4]
  wire [4:0] _T_59243; // @[Modules.scala 46:37:@5733.4]
  wire [4:0] _T_59244; // @[Modules.scala 46:37:@5734.4]
  wire [5:0] _T_59245; // @[Modules.scala 46:47:@5735.4]
  wire [4:0] _T_59246; // @[Modules.scala 46:47:@5736.4]
  wire [4:0] _T_59247; // @[Modules.scala 46:47:@5737.4]
  wire [5:0] _T_59249; // @[Modules.scala 43:37:@5739.4]
  wire [4:0] _T_59250; // @[Modules.scala 43:37:@5740.4]
  wire [4:0] _T_59251; // @[Modules.scala 43:37:@5741.4]
  wire [5:0] _T_59252; // @[Modules.scala 43:47:@5742.4]
  wire [4:0] _T_59253; // @[Modules.scala 43:47:@5743.4]
  wire [4:0] _T_59254; // @[Modules.scala 43:47:@5744.4]
  wire [5:0] _T_59256; // @[Modules.scala 46:37:@5746.4]
  wire [4:0] _T_59257; // @[Modules.scala 46:37:@5747.4]
  wire [4:0] _T_59258; // @[Modules.scala 46:37:@5748.4]
  wire [5:0] _T_59259; // @[Modules.scala 46:47:@5749.4]
  wire [4:0] _T_59260; // @[Modules.scala 46:47:@5750.4]
  wire [4:0] _T_59261; // @[Modules.scala 46:47:@5751.4]
  wire [5:0] _T_59263; // @[Modules.scala 43:37:@5753.4]
  wire [4:0] _T_59264; // @[Modules.scala 43:37:@5754.4]
  wire [4:0] _T_59265; // @[Modules.scala 43:37:@5755.4]
  wire [5:0] _T_59266; // @[Modules.scala 43:47:@5756.4]
  wire [4:0] _T_59267; // @[Modules.scala 43:47:@5757.4]
  wire [4:0] _T_59268; // @[Modules.scala 43:47:@5758.4]
  wire [5:0] _T_59269; // @[Modules.scala 40:46:@5760.4]
  wire [4:0] _T_59270; // @[Modules.scala 40:46:@5761.4]
  wire [4:0] _T_59271; // @[Modules.scala 40:46:@5762.4]
  wire [5:0] _T_59273; // @[Modules.scala 46:37:@5764.4]
  wire [4:0] _T_59274; // @[Modules.scala 46:37:@5765.4]
  wire [4:0] _T_59275; // @[Modules.scala 46:37:@5766.4]
  wire [5:0] _T_59276; // @[Modules.scala 46:47:@5767.4]
  wire [4:0] _T_59277; // @[Modules.scala 46:47:@5768.4]
  wire [4:0] _T_59278; // @[Modules.scala 46:47:@5769.4]
  wire [5:0] _T_59280; // @[Modules.scala 46:37:@5771.4]
  wire [4:0] _T_59281; // @[Modules.scala 46:37:@5772.4]
  wire [4:0] _T_59282; // @[Modules.scala 46:37:@5773.4]
  wire [5:0] _T_59283; // @[Modules.scala 46:47:@5774.4]
  wire [4:0] _T_59284; // @[Modules.scala 46:47:@5775.4]
  wire [4:0] _T_59285; // @[Modules.scala 46:47:@5776.4]
  wire [5:0] _T_59289; // @[Modules.scala 37:46:@5782.4]
  wire [4:0] _T_59290; // @[Modules.scala 37:46:@5783.4]
  wire [4:0] _T_59291; // @[Modules.scala 37:46:@5784.4]
  wire [5:0] _T_59292; // @[Modules.scala 40:46:@5786.4]
  wire [4:0] _T_59293; // @[Modules.scala 40:46:@5787.4]
  wire [4:0] _T_59294; // @[Modules.scala 40:46:@5788.4]
  wire [5:0] _T_59296; // @[Modules.scala 46:37:@5790.4]
  wire [4:0] _T_59297; // @[Modules.scala 46:37:@5791.4]
  wire [4:0] _T_59298; // @[Modules.scala 46:37:@5792.4]
  wire [5:0] _T_59299; // @[Modules.scala 46:47:@5793.4]
  wire [4:0] _T_59300; // @[Modules.scala 46:47:@5794.4]
  wire [4:0] _T_59301; // @[Modules.scala 46:47:@5795.4]
  wire [5:0] _T_59306; // @[Modules.scala 46:47:@5800.4]
  wire [4:0] _T_59307; // @[Modules.scala 46:47:@5801.4]
  wire [4:0] _T_59308; // @[Modules.scala 46:47:@5802.4]
  wire [5:0] _T_59310; // @[Modules.scala 46:37:@5804.4]
  wire [4:0] _T_59311; // @[Modules.scala 46:37:@5805.4]
  wire [4:0] _T_59312; // @[Modules.scala 46:37:@5806.4]
  wire [5:0] _T_59313; // @[Modules.scala 46:47:@5807.4]
  wire [4:0] _T_59314; // @[Modules.scala 46:47:@5808.4]
  wire [4:0] _T_59315; // @[Modules.scala 46:47:@5809.4]
  wire [5:0] _T_59317; // @[Modules.scala 46:37:@5811.4]
  wire [4:0] _T_59318; // @[Modules.scala 46:37:@5812.4]
  wire [4:0] _T_59319; // @[Modules.scala 46:37:@5813.4]
  wire [5:0] _T_59320; // @[Modules.scala 46:47:@5814.4]
  wire [4:0] _T_59321; // @[Modules.scala 46:47:@5815.4]
  wire [4:0] _T_59322; // @[Modules.scala 46:47:@5816.4]
  wire [5:0] _T_59338; // @[Modules.scala 46:37:@5832.4]
  wire [4:0] _T_59339; // @[Modules.scala 46:37:@5833.4]
  wire [4:0] _T_59340; // @[Modules.scala 46:37:@5834.4]
  wire [5:0] _T_59341; // @[Modules.scala 46:47:@5835.4]
  wire [4:0] _T_59342; // @[Modules.scala 46:47:@5836.4]
  wire [4:0] _T_59343; // @[Modules.scala 46:47:@5837.4]
  wire [5:0] _T_59345; // @[Modules.scala 46:37:@5839.4]
  wire [4:0] _T_59346; // @[Modules.scala 46:37:@5840.4]
  wire [4:0] _T_59347; // @[Modules.scala 46:37:@5841.4]
  wire [5:0] _T_59348; // @[Modules.scala 46:47:@5842.4]
  wire [4:0] _T_59349; // @[Modules.scala 46:47:@5843.4]
  wire [4:0] _T_59350; // @[Modules.scala 46:47:@5844.4]
  wire [5:0] _T_59377; // @[Modules.scala 40:46:@5876.4]
  wire [4:0] _T_59378; // @[Modules.scala 40:46:@5877.4]
  wire [4:0] _T_59379; // @[Modules.scala 40:46:@5878.4]
  wire [5:0] _T_59380; // @[Modules.scala 37:46:@5880.4]
  wire [4:0] _T_59381; // @[Modules.scala 37:46:@5881.4]
  wire [4:0] _T_59382; // @[Modules.scala 37:46:@5882.4]
  wire [5:0] _T_59383; // @[Modules.scala 37:46:@5884.4]
  wire [4:0] _T_59384; // @[Modules.scala 37:46:@5885.4]
  wire [4:0] _T_59385; // @[Modules.scala 37:46:@5886.4]
  wire [5:0] _T_59386; // @[Modules.scala 37:46:@5888.4]
  wire [4:0] _T_59387; // @[Modules.scala 37:46:@5889.4]
  wire [4:0] _T_59388; // @[Modules.scala 37:46:@5890.4]
  wire [5:0] _T_59396; // @[Modules.scala 37:46:@5899.4]
  wire [4:0] _T_59397; // @[Modules.scala 37:46:@5900.4]
  wire [4:0] _T_59398; // @[Modules.scala 37:46:@5901.4]
  wire [5:0] _T_59400; // @[Modules.scala 46:37:@5903.4]
  wire [4:0] _T_59401; // @[Modules.scala 46:37:@5904.4]
  wire [4:0] _T_59402; // @[Modules.scala 46:37:@5905.4]
  wire [5:0] _T_59403; // @[Modules.scala 46:47:@5906.4]
  wire [4:0] _T_59404; // @[Modules.scala 46:47:@5907.4]
  wire [4:0] _T_59405; // @[Modules.scala 46:47:@5908.4]
  wire [5:0] _T_59410; // @[Modules.scala 46:47:@5913.4]
  wire [4:0] _T_59411; // @[Modules.scala 46:47:@5914.4]
  wire [4:0] _T_59412; // @[Modules.scala 46:47:@5915.4]
  wire [5:0] _T_59428; // @[Modules.scala 46:37:@5931.4]
  wire [4:0] _T_59429; // @[Modules.scala 46:37:@5932.4]
  wire [4:0] _T_59430; // @[Modules.scala 46:37:@5933.4]
  wire [5:0] _T_59431; // @[Modules.scala 46:47:@5934.4]
  wire [4:0] _T_59432; // @[Modules.scala 46:47:@5935.4]
  wire [4:0] _T_59433; // @[Modules.scala 46:47:@5936.4]
  wire [5:0] _T_59441; // @[Modules.scala 40:46:@5945.4]
  wire [4:0] _T_59442; // @[Modules.scala 40:46:@5946.4]
  wire [4:0] _T_59443; // @[Modules.scala 40:46:@5947.4]
  wire [5:0] _T_59445; // @[Modules.scala 46:37:@5949.4]
  wire [4:0] _T_59446; // @[Modules.scala 46:37:@5950.4]
  wire [4:0] _T_59447; // @[Modules.scala 46:37:@5951.4]
  wire [5:0] _T_59448; // @[Modules.scala 46:47:@5952.4]
  wire [4:0] _T_59449; // @[Modules.scala 46:47:@5953.4]
  wire [4:0] _T_59450; // @[Modules.scala 46:47:@5954.4]
  wire [10:0] buffer_1_0; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59451; // @[Modules.scala 50:57:@5956.4]
  wire [10:0] _T_59452; // @[Modules.scala 50:57:@5957.4]
  wire [10:0] buffer_1_392; // @[Modules.scala 50:57:@5958.4]
  wire [10:0] buffer_1_2; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_3; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59454; // @[Modules.scala 50:57:@5960.4]
  wire [10:0] _T_59455; // @[Modules.scala 50:57:@5961.4]
  wire [10:0] buffer_1_393; // @[Modules.scala 50:57:@5962.4]
  wire [10:0] buffer_1_4; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59457; // @[Modules.scala 50:57:@5964.4]
  wire [10:0] _T_59458; // @[Modules.scala 50:57:@5965.4]
  wire [10:0] buffer_1_394; // @[Modules.scala 50:57:@5966.4]
  wire [10:0] buffer_1_6; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_7; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59460; // @[Modules.scala 50:57:@5968.4]
  wire [10:0] _T_59461; // @[Modules.scala 50:57:@5969.4]
  wire [10:0] buffer_1_395; // @[Modules.scala 50:57:@5970.4]
  wire [10:0] buffer_1_8; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59463; // @[Modules.scala 50:57:@5972.4]
  wire [10:0] _T_59464; // @[Modules.scala 50:57:@5973.4]
  wire [10:0] buffer_1_396; // @[Modules.scala 50:57:@5974.4]
  wire [10:0] buffer_1_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59466; // @[Modules.scala 50:57:@5976.4]
  wire [10:0] _T_59467; // @[Modules.scala 50:57:@5977.4]
  wire [10:0] buffer_1_397; // @[Modules.scala 50:57:@5978.4]
  wire [10:0] buffer_1_12; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59469; // @[Modules.scala 50:57:@5980.4]
  wire [10:0] _T_59470; // @[Modules.scala 50:57:@5981.4]
  wire [10:0] buffer_1_398; // @[Modules.scala 50:57:@5982.4]
  wire [10:0] buffer_1_14; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59472; // @[Modules.scala 50:57:@5984.4]
  wire [10:0] _T_59473; // @[Modules.scala 50:57:@5985.4]
  wire [10:0] buffer_1_399; // @[Modules.scala 50:57:@5986.4]
  wire [10:0] buffer_1_17; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59475; // @[Modules.scala 50:57:@5988.4]
  wire [10:0] _T_59476; // @[Modules.scala 50:57:@5989.4]
  wire [10:0] buffer_1_400; // @[Modules.scala 50:57:@5990.4]
  wire [10:0] buffer_1_18; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_19; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59478; // @[Modules.scala 50:57:@5992.4]
  wire [10:0] _T_59479; // @[Modules.scala 50:57:@5993.4]
  wire [10:0] buffer_1_401; // @[Modules.scala 50:57:@5994.4]
  wire [10:0] buffer_1_20; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_21; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59481; // @[Modules.scala 50:57:@5996.4]
  wire [10:0] _T_59482; // @[Modules.scala 50:57:@5997.4]
  wire [10:0] buffer_1_402; // @[Modules.scala 50:57:@5998.4]
  wire [10:0] buffer_1_22; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_23; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59484; // @[Modules.scala 50:57:@6000.4]
  wire [10:0] _T_59485; // @[Modules.scala 50:57:@6001.4]
  wire [10:0] buffer_1_403; // @[Modules.scala 50:57:@6002.4]
  wire [10:0] buffer_1_24; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_25; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59487; // @[Modules.scala 50:57:@6004.4]
  wire [10:0] _T_59488; // @[Modules.scala 50:57:@6005.4]
  wire [10:0] buffer_1_404; // @[Modules.scala 50:57:@6006.4]
  wire [10:0] buffer_1_26; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59490; // @[Modules.scala 50:57:@6008.4]
  wire [10:0] _T_59491; // @[Modules.scala 50:57:@6009.4]
  wire [10:0] buffer_1_405; // @[Modules.scala 50:57:@6010.4]
  wire [10:0] buffer_1_28; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59493; // @[Modules.scala 50:57:@6012.4]
  wire [10:0] _T_59494; // @[Modules.scala 50:57:@6013.4]
  wire [10:0] buffer_1_406; // @[Modules.scala 50:57:@6014.4]
  wire [10:0] buffer_1_30; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_31; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59496; // @[Modules.scala 50:57:@6016.4]
  wire [10:0] _T_59497; // @[Modules.scala 50:57:@6017.4]
  wire [10:0] buffer_1_407; // @[Modules.scala 50:57:@6018.4]
  wire [10:0] buffer_1_32; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_33; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59499; // @[Modules.scala 50:57:@6020.4]
  wire [10:0] _T_59500; // @[Modules.scala 50:57:@6021.4]
  wire [10:0] buffer_1_408; // @[Modules.scala 50:57:@6022.4]
  wire [10:0] buffer_1_34; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59502; // @[Modules.scala 50:57:@6024.4]
  wire [10:0] _T_59503; // @[Modules.scala 50:57:@6025.4]
  wire [10:0] buffer_1_409; // @[Modules.scala 50:57:@6026.4]
  wire [10:0] buffer_1_36; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_37; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59505; // @[Modules.scala 50:57:@6028.4]
  wire [10:0] _T_59506; // @[Modules.scala 50:57:@6029.4]
  wire [10:0] buffer_1_410; // @[Modules.scala 50:57:@6030.4]
  wire [10:0] buffer_1_38; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59508; // @[Modules.scala 50:57:@6032.4]
  wire [10:0] _T_59509; // @[Modules.scala 50:57:@6033.4]
  wire [10:0] buffer_1_411; // @[Modules.scala 50:57:@6034.4]
  wire [10:0] buffer_1_40; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59511; // @[Modules.scala 50:57:@6036.4]
  wire [10:0] _T_59512; // @[Modules.scala 50:57:@6037.4]
  wire [10:0] buffer_1_412; // @[Modules.scala 50:57:@6038.4]
  wire [10:0] buffer_1_42; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59514; // @[Modules.scala 50:57:@6040.4]
  wire [10:0] _T_59515; // @[Modules.scala 50:57:@6041.4]
  wire [10:0] buffer_1_413; // @[Modules.scala 50:57:@6042.4]
  wire [10:0] buffer_1_46; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59520; // @[Modules.scala 50:57:@6048.4]
  wire [10:0] _T_59521; // @[Modules.scala 50:57:@6049.4]
  wire [10:0] buffer_1_415; // @[Modules.scala 50:57:@6050.4]
  wire [10:0] buffer_1_48; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59523; // @[Modules.scala 50:57:@6052.4]
  wire [10:0] _T_59524; // @[Modules.scala 50:57:@6053.4]
  wire [10:0] buffer_1_416; // @[Modules.scala 50:57:@6054.4]
  wire [10:0] buffer_1_54; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59532; // @[Modules.scala 50:57:@6064.4]
  wire [10:0] _T_59533; // @[Modules.scala 50:57:@6065.4]
  wire [10:0] buffer_1_419; // @[Modules.scala 50:57:@6066.4]
  wire [10:0] buffer_1_56; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59535; // @[Modules.scala 50:57:@6068.4]
  wire [10:0] _T_59536; // @[Modules.scala 50:57:@6069.4]
  wire [10:0] buffer_1_420; // @[Modules.scala 50:57:@6070.4]
  wire [10:0] buffer_1_59; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59538; // @[Modules.scala 50:57:@6072.4]
  wire [10:0] _T_59539; // @[Modules.scala 50:57:@6073.4]
  wire [10:0] buffer_1_421; // @[Modules.scala 50:57:@6074.4]
  wire [10:0] buffer_1_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59544; // @[Modules.scala 50:57:@6080.4]
  wire [10:0] _T_59545; // @[Modules.scala 50:57:@6081.4]
  wire [10:0] buffer_1_423; // @[Modules.scala 50:57:@6082.4]
  wire [10:0] buffer_1_64; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_65; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59547; // @[Modules.scala 50:57:@6084.4]
  wire [10:0] _T_59548; // @[Modules.scala 50:57:@6085.4]
  wire [10:0] buffer_1_424; // @[Modules.scala 50:57:@6086.4]
  wire [10:0] buffer_1_66; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59550; // @[Modules.scala 50:57:@6088.4]
  wire [10:0] _T_59551; // @[Modules.scala 50:57:@6089.4]
  wire [10:0] buffer_1_425; // @[Modules.scala 50:57:@6090.4]
  wire [10:0] buffer_1_68; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59553; // @[Modules.scala 50:57:@6092.4]
  wire [10:0] _T_59554; // @[Modules.scala 50:57:@6093.4]
  wire [10:0] buffer_1_426; // @[Modules.scala 50:57:@6094.4]
  wire [10:0] buffer_1_70; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59556; // @[Modules.scala 50:57:@6096.4]
  wire [10:0] _T_59557; // @[Modules.scala 50:57:@6097.4]
  wire [10:0] buffer_1_427; // @[Modules.scala 50:57:@6098.4]
  wire [10:0] buffer_1_72; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59559; // @[Modules.scala 50:57:@6100.4]
  wire [10:0] _T_59560; // @[Modules.scala 50:57:@6101.4]
  wire [10:0] buffer_1_428; // @[Modules.scala 50:57:@6102.4]
  wire [10:0] buffer_1_74; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59562; // @[Modules.scala 50:57:@6104.4]
  wire [10:0] _T_59563; // @[Modules.scala 50:57:@6105.4]
  wire [10:0] buffer_1_429; // @[Modules.scala 50:57:@6106.4]
  wire [10:0] buffer_1_78; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59568; // @[Modules.scala 50:57:@6112.4]
  wire [10:0] _T_59569; // @[Modules.scala 50:57:@6113.4]
  wire [10:0] buffer_1_431; // @[Modules.scala 50:57:@6114.4]
  wire [10:0] buffer_1_81; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59571; // @[Modules.scala 50:57:@6116.4]
  wire [10:0] _T_59572; // @[Modules.scala 50:57:@6117.4]
  wire [10:0] buffer_1_432; // @[Modules.scala 50:57:@6118.4]
  wire [10:0] buffer_1_82; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59574; // @[Modules.scala 50:57:@6120.4]
  wire [10:0] _T_59575; // @[Modules.scala 50:57:@6121.4]
  wire [10:0] buffer_1_433; // @[Modules.scala 50:57:@6122.4]
  wire [10:0] buffer_1_84; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59577; // @[Modules.scala 50:57:@6124.4]
  wire [10:0] _T_59578; // @[Modules.scala 50:57:@6125.4]
  wire [10:0] buffer_1_434; // @[Modules.scala 50:57:@6126.4]
  wire [10:0] buffer_1_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59580; // @[Modules.scala 50:57:@6128.4]
  wire [10:0] _T_59581; // @[Modules.scala 50:57:@6129.4]
  wire [10:0] buffer_1_435; // @[Modules.scala 50:57:@6130.4]
  wire [10:0] buffer_1_88; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59583; // @[Modules.scala 50:57:@6132.4]
  wire [10:0] _T_59584; // @[Modules.scala 50:57:@6133.4]
  wire [10:0] buffer_1_436; // @[Modules.scala 50:57:@6134.4]
  wire [10:0] buffer_1_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59586; // @[Modules.scala 50:57:@6136.4]
  wire [10:0] _T_59587; // @[Modules.scala 50:57:@6137.4]
  wire [10:0] buffer_1_437; // @[Modules.scala 50:57:@6138.4]
  wire [10:0] buffer_1_94; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59592; // @[Modules.scala 50:57:@6144.4]
  wire [10:0] _T_59593; // @[Modules.scala 50:57:@6145.4]
  wire [10:0] buffer_1_439; // @[Modules.scala 50:57:@6146.4]
  wire [10:0] buffer_1_96; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59595; // @[Modules.scala 50:57:@6148.4]
  wire [10:0] _T_59596; // @[Modules.scala 50:57:@6149.4]
  wire [10:0] buffer_1_440; // @[Modules.scala 50:57:@6150.4]
  wire [10:0] buffer_1_98; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59598; // @[Modules.scala 50:57:@6152.4]
  wire [10:0] _T_59599; // @[Modules.scala 50:57:@6153.4]
  wire [10:0] buffer_1_441; // @[Modules.scala 50:57:@6154.4]
  wire [10:0] buffer_1_100; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59601; // @[Modules.scala 50:57:@6156.4]
  wire [10:0] _T_59602; // @[Modules.scala 50:57:@6157.4]
  wire [10:0] buffer_1_442; // @[Modules.scala 50:57:@6158.4]
  wire [10:0] buffer_1_102; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59604; // @[Modules.scala 50:57:@6160.4]
  wire [10:0] _T_59605; // @[Modules.scala 50:57:@6161.4]
  wire [10:0] buffer_1_443; // @[Modules.scala 50:57:@6162.4]
  wire [10:0] buffer_1_104; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59607; // @[Modules.scala 50:57:@6164.4]
  wire [10:0] _T_59608; // @[Modules.scala 50:57:@6165.4]
  wire [10:0] buffer_1_444; // @[Modules.scala 50:57:@6166.4]
  wire [10:0] buffer_1_106; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59610; // @[Modules.scala 50:57:@6168.4]
  wire [10:0] _T_59611; // @[Modules.scala 50:57:@6169.4]
  wire [10:0] buffer_1_445; // @[Modules.scala 50:57:@6170.4]
  wire [10:0] buffer_1_108; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59613; // @[Modules.scala 50:57:@6172.4]
  wire [10:0] _T_59614; // @[Modules.scala 50:57:@6173.4]
  wire [10:0] buffer_1_446; // @[Modules.scala 50:57:@6174.4]
  wire [10:0] buffer_1_110; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59616; // @[Modules.scala 50:57:@6176.4]
  wire [10:0] _T_59617; // @[Modules.scala 50:57:@6177.4]
  wire [10:0] buffer_1_447; // @[Modules.scala 50:57:@6178.4]
  wire [10:0] buffer_1_112; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59619; // @[Modules.scala 50:57:@6180.4]
  wire [10:0] _T_59620; // @[Modules.scala 50:57:@6181.4]
  wire [10:0] buffer_1_448; // @[Modules.scala 50:57:@6182.4]
  wire [10:0] buffer_1_118; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59628; // @[Modules.scala 50:57:@6192.4]
  wire [10:0] _T_59629; // @[Modules.scala 50:57:@6193.4]
  wire [10:0] buffer_1_451; // @[Modules.scala 50:57:@6194.4]
  wire [10:0] buffer_1_120; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59631; // @[Modules.scala 50:57:@6196.4]
  wire [10:0] _T_59632; // @[Modules.scala 50:57:@6197.4]
  wire [10:0] buffer_1_452; // @[Modules.scala 50:57:@6198.4]
  wire [10:0] buffer_1_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59634; // @[Modules.scala 50:57:@6200.4]
  wire [10:0] _T_59635; // @[Modules.scala 50:57:@6201.4]
  wire [10:0] buffer_1_453; // @[Modules.scala 50:57:@6202.4]
  wire [10:0] buffer_1_124; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_125; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59637; // @[Modules.scala 50:57:@6204.4]
  wire [10:0] _T_59638; // @[Modules.scala 50:57:@6205.4]
  wire [10:0] buffer_1_454; // @[Modules.scala 50:57:@6206.4]
  wire [10:0] buffer_1_126; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59640; // @[Modules.scala 50:57:@6208.4]
  wire [10:0] _T_59641; // @[Modules.scala 50:57:@6209.4]
  wire [10:0] buffer_1_455; // @[Modules.scala 50:57:@6210.4]
  wire [10:0] buffer_1_130; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59646; // @[Modules.scala 50:57:@6216.4]
  wire [10:0] _T_59647; // @[Modules.scala 50:57:@6217.4]
  wire [10:0] buffer_1_457; // @[Modules.scala 50:57:@6218.4]
  wire [10:0] buffer_1_133; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59649; // @[Modules.scala 50:57:@6220.4]
  wire [10:0] _T_59650; // @[Modules.scala 50:57:@6221.4]
  wire [10:0] buffer_1_458; // @[Modules.scala 50:57:@6222.4]
  wire [10:0] buffer_1_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59655; // @[Modules.scala 50:57:@6228.4]
  wire [10:0] _T_59656; // @[Modules.scala 50:57:@6229.4]
  wire [10:0] buffer_1_460; // @[Modules.scala 50:57:@6230.4]
  wire [10:0] buffer_1_138; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_139; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59658; // @[Modules.scala 50:57:@6232.4]
  wire [10:0] _T_59659; // @[Modules.scala 50:57:@6233.4]
  wire [10:0] buffer_1_461; // @[Modules.scala 50:57:@6234.4]
  wire [10:0] buffer_1_140; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59661; // @[Modules.scala 50:57:@6236.4]
  wire [10:0] _T_59662; // @[Modules.scala 50:57:@6237.4]
  wire [10:0] buffer_1_462; // @[Modules.scala 50:57:@6238.4]
  wire [10:0] buffer_1_146; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59670; // @[Modules.scala 50:57:@6248.4]
  wire [10:0] _T_59671; // @[Modules.scala 50:57:@6249.4]
  wire [10:0] buffer_1_465; // @[Modules.scala 50:57:@6250.4]
  wire [10:0] buffer_1_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59676; // @[Modules.scala 50:57:@6256.4]
  wire [10:0] _T_59677; // @[Modules.scala 50:57:@6257.4]
  wire [10:0] buffer_1_467; // @[Modules.scala 50:57:@6258.4]
  wire [10:0] buffer_1_152; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_153; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59679; // @[Modules.scala 50:57:@6260.4]
  wire [10:0] _T_59680; // @[Modules.scala 50:57:@6261.4]
  wire [10:0] buffer_1_468; // @[Modules.scala 50:57:@6262.4]
  wire [10:0] buffer_1_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59685; // @[Modules.scala 50:57:@6268.4]
  wire [10:0] _T_59686; // @[Modules.scala 50:57:@6269.4]
  wire [10:0] buffer_1_470; // @[Modules.scala 50:57:@6270.4]
  wire [10:0] buffer_1_158; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59688; // @[Modules.scala 50:57:@6272.4]
  wire [10:0] _T_59689; // @[Modules.scala 50:57:@6273.4]
  wire [10:0] buffer_1_471; // @[Modules.scala 50:57:@6274.4]
  wire [10:0] buffer_1_160; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59691; // @[Modules.scala 50:57:@6276.4]
  wire [10:0] _T_59692; // @[Modules.scala 50:57:@6277.4]
  wire [10:0] buffer_1_472; // @[Modules.scala 50:57:@6278.4]
  wire [10:0] buffer_1_162; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59694; // @[Modules.scala 50:57:@6280.4]
  wire [10:0] _T_59695; // @[Modules.scala 50:57:@6281.4]
  wire [10:0] buffer_1_473; // @[Modules.scala 50:57:@6282.4]
  wire [10:0] buffer_1_164; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_165; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59697; // @[Modules.scala 50:57:@6284.4]
  wire [10:0] _T_59698; // @[Modules.scala 50:57:@6285.4]
  wire [10:0] buffer_1_474; // @[Modules.scala 50:57:@6286.4]
  wire [10:0] buffer_1_166; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59700; // @[Modules.scala 50:57:@6288.4]
  wire [10:0] _T_59701; // @[Modules.scala 50:57:@6289.4]
  wire [10:0] buffer_1_475; // @[Modules.scala 50:57:@6290.4]
  wire [10:0] buffer_1_175; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59712; // @[Modules.scala 50:57:@6304.4]
  wire [10:0] _T_59713; // @[Modules.scala 50:57:@6305.4]
  wire [10:0] buffer_1_479; // @[Modules.scala 50:57:@6306.4]
  wire [10:0] buffer_1_176; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59715; // @[Modules.scala 50:57:@6308.4]
  wire [10:0] _T_59716; // @[Modules.scala 50:57:@6309.4]
  wire [10:0] buffer_1_480; // @[Modules.scala 50:57:@6310.4]
  wire [10:0] buffer_1_178; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59718; // @[Modules.scala 50:57:@6312.4]
  wire [10:0] _T_59719; // @[Modules.scala 50:57:@6313.4]
  wire [10:0] buffer_1_481; // @[Modules.scala 50:57:@6314.4]
  wire [10:0] buffer_1_180; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59721; // @[Modules.scala 50:57:@6316.4]
  wire [10:0] _T_59722; // @[Modules.scala 50:57:@6317.4]
  wire [10:0] buffer_1_482; // @[Modules.scala 50:57:@6318.4]
  wire [10:0] buffer_1_184; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59727; // @[Modules.scala 50:57:@6324.4]
  wire [10:0] _T_59728; // @[Modules.scala 50:57:@6325.4]
  wire [10:0] buffer_1_484; // @[Modules.scala 50:57:@6326.4]
  wire [10:0] buffer_1_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59733; // @[Modules.scala 50:57:@6332.4]
  wire [10:0] _T_59734; // @[Modules.scala 50:57:@6333.4]
  wire [10:0] buffer_1_486; // @[Modules.scala 50:57:@6334.4]
  wire [10:0] buffer_1_190; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59736; // @[Modules.scala 50:57:@6336.4]
  wire [10:0] _T_59737; // @[Modules.scala 50:57:@6337.4]
  wire [10:0] buffer_1_487; // @[Modules.scala 50:57:@6338.4]
  wire [10:0] buffer_1_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59742; // @[Modules.scala 50:57:@6344.4]
  wire [10:0] _T_59743; // @[Modules.scala 50:57:@6345.4]
  wire [10:0] buffer_1_489; // @[Modules.scala 50:57:@6346.4]
  wire [10:0] buffer_1_196; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59745; // @[Modules.scala 50:57:@6348.4]
  wire [10:0] _T_59746; // @[Modules.scala 50:57:@6349.4]
  wire [10:0] buffer_1_490; // @[Modules.scala 50:57:@6350.4]
  wire [10:0] buffer_1_198; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59748; // @[Modules.scala 50:57:@6352.4]
  wire [10:0] _T_59749; // @[Modules.scala 50:57:@6353.4]
  wire [10:0] buffer_1_491; // @[Modules.scala 50:57:@6354.4]
  wire [10:0] buffer_1_202; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59754; // @[Modules.scala 50:57:@6360.4]
  wire [10:0] _T_59755; // @[Modules.scala 50:57:@6361.4]
  wire [10:0] buffer_1_493; // @[Modules.scala 50:57:@6362.4]
  wire [10:0] buffer_1_204; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59757; // @[Modules.scala 50:57:@6364.4]
  wire [10:0] _T_59758; // @[Modules.scala 50:57:@6365.4]
  wire [10:0] buffer_1_494; // @[Modules.scala 50:57:@6366.4]
  wire [10:0] buffer_1_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59763; // @[Modules.scala 50:57:@6372.4]
  wire [10:0] _T_59764; // @[Modules.scala 50:57:@6373.4]
  wire [10:0] buffer_1_496; // @[Modules.scala 50:57:@6374.4]
  wire [10:0] buffer_1_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59766; // @[Modules.scala 50:57:@6376.4]
  wire [10:0] _T_59767; // @[Modules.scala 50:57:@6377.4]
  wire [10:0] buffer_1_497; // @[Modules.scala 50:57:@6378.4]
  wire [10:0] buffer_1_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59769; // @[Modules.scala 50:57:@6380.4]
  wire [10:0] _T_59770; // @[Modules.scala 50:57:@6381.4]
  wire [10:0] buffer_1_498; // @[Modules.scala 50:57:@6382.4]
  wire [10:0] buffer_1_216; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59775; // @[Modules.scala 50:57:@6388.4]
  wire [10:0] _T_59776; // @[Modules.scala 50:57:@6389.4]
  wire [10:0] buffer_1_500; // @[Modules.scala 50:57:@6390.4]
  wire [10:0] buffer_1_218; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59778; // @[Modules.scala 50:57:@6392.4]
  wire [10:0] _T_59779; // @[Modules.scala 50:57:@6393.4]
  wire [10:0] buffer_1_501; // @[Modules.scala 50:57:@6394.4]
  wire [10:0] buffer_1_220; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59781; // @[Modules.scala 50:57:@6396.4]
  wire [10:0] _T_59782; // @[Modules.scala 50:57:@6397.4]
  wire [10:0] buffer_1_502; // @[Modules.scala 50:57:@6398.4]
  wire [10:0] buffer_1_222; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59784; // @[Modules.scala 50:57:@6400.4]
  wire [10:0] _T_59785; // @[Modules.scala 50:57:@6401.4]
  wire [10:0] buffer_1_503; // @[Modules.scala 50:57:@6402.4]
  wire [10:0] buffer_1_224; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59787; // @[Modules.scala 50:57:@6404.4]
  wire [10:0] _T_59788; // @[Modules.scala 50:57:@6405.4]
  wire [10:0] buffer_1_504; // @[Modules.scala 50:57:@6406.4]
  wire [10:0] buffer_1_226; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59790; // @[Modules.scala 50:57:@6408.4]
  wire [10:0] _T_59791; // @[Modules.scala 50:57:@6409.4]
  wire [10:0] buffer_1_505; // @[Modules.scala 50:57:@6410.4]
  wire [10:0] buffer_1_228; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59793; // @[Modules.scala 50:57:@6412.4]
  wire [10:0] _T_59794; // @[Modules.scala 50:57:@6413.4]
  wire [10:0] buffer_1_506; // @[Modules.scala 50:57:@6414.4]
  wire [10:0] buffer_1_230; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59796; // @[Modules.scala 50:57:@6416.4]
  wire [10:0] _T_59797; // @[Modules.scala 50:57:@6417.4]
  wire [10:0] buffer_1_507; // @[Modules.scala 50:57:@6418.4]
  wire [10:0] buffer_1_232; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59799; // @[Modules.scala 50:57:@6420.4]
  wire [10:0] _T_59800; // @[Modules.scala 50:57:@6421.4]
  wire [10:0] buffer_1_508; // @[Modules.scala 50:57:@6422.4]
  wire [10:0] buffer_1_234; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59802; // @[Modules.scala 50:57:@6424.4]
  wire [10:0] _T_59803; // @[Modules.scala 50:57:@6425.4]
  wire [10:0] buffer_1_509; // @[Modules.scala 50:57:@6426.4]
  wire [10:0] buffer_1_236; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59805; // @[Modules.scala 50:57:@6428.4]
  wire [10:0] _T_59806; // @[Modules.scala 50:57:@6429.4]
  wire [10:0] buffer_1_510; // @[Modules.scala 50:57:@6430.4]
  wire [10:0] buffer_1_238; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59808; // @[Modules.scala 50:57:@6432.4]
  wire [10:0] _T_59809; // @[Modules.scala 50:57:@6433.4]
  wire [10:0] buffer_1_511; // @[Modules.scala 50:57:@6434.4]
  wire [10:0] buffer_1_242; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_243; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59814; // @[Modules.scala 50:57:@6440.4]
  wire [10:0] _T_59815; // @[Modules.scala 50:57:@6441.4]
  wire [10:0] buffer_1_513; // @[Modules.scala 50:57:@6442.4]
  wire [10:0] buffer_1_244; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59817; // @[Modules.scala 50:57:@6444.4]
  wire [10:0] _T_59818; // @[Modules.scala 50:57:@6445.4]
  wire [10:0] buffer_1_514; // @[Modules.scala 50:57:@6446.4]
  wire [10:0] buffer_1_246; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59820; // @[Modules.scala 50:57:@6448.4]
  wire [10:0] _T_59821; // @[Modules.scala 50:57:@6449.4]
  wire [10:0] buffer_1_515; // @[Modules.scala 50:57:@6450.4]
  wire [10:0] buffer_1_248; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59823; // @[Modules.scala 50:57:@6452.4]
  wire [10:0] _T_59824; // @[Modules.scala 50:57:@6453.4]
  wire [10:0] buffer_1_516; // @[Modules.scala 50:57:@6454.4]
  wire [10:0] buffer_1_252; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59829; // @[Modules.scala 50:57:@6460.4]
  wire [10:0] _T_59830; // @[Modules.scala 50:57:@6461.4]
  wire [10:0] buffer_1_518; // @[Modules.scala 50:57:@6462.4]
  wire [10:0] buffer_1_254; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59832; // @[Modules.scala 50:57:@6464.4]
  wire [10:0] _T_59833; // @[Modules.scala 50:57:@6465.4]
  wire [10:0] buffer_1_519; // @[Modules.scala 50:57:@6466.4]
  wire [10:0] buffer_1_256; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59835; // @[Modules.scala 50:57:@6468.4]
  wire [10:0] _T_59836; // @[Modules.scala 50:57:@6469.4]
  wire [10:0] buffer_1_520; // @[Modules.scala 50:57:@6470.4]
  wire [10:0] buffer_1_258; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59838; // @[Modules.scala 50:57:@6472.4]
  wire [10:0] _T_59839; // @[Modules.scala 50:57:@6473.4]
  wire [10:0] buffer_1_521; // @[Modules.scala 50:57:@6474.4]
  wire [10:0] buffer_1_260; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_261; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59841; // @[Modules.scala 50:57:@6476.4]
  wire [10:0] _T_59842; // @[Modules.scala 50:57:@6477.4]
  wire [10:0] buffer_1_522; // @[Modules.scala 50:57:@6478.4]
  wire [10:0] buffer_1_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59844; // @[Modules.scala 50:57:@6480.4]
  wire [10:0] _T_59845; // @[Modules.scala 50:57:@6481.4]
  wire [10:0] buffer_1_523; // @[Modules.scala 50:57:@6482.4]
  wire [10:0] buffer_1_264; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59847; // @[Modules.scala 50:57:@6484.4]
  wire [10:0] _T_59848; // @[Modules.scala 50:57:@6485.4]
  wire [10:0] buffer_1_524; // @[Modules.scala 50:57:@6486.4]
  wire [10:0] buffer_1_266; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_267; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59850; // @[Modules.scala 50:57:@6488.4]
  wire [10:0] _T_59851; // @[Modules.scala 50:57:@6489.4]
  wire [10:0] buffer_1_525; // @[Modules.scala 50:57:@6490.4]
  wire [10:0] buffer_1_268; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59853; // @[Modules.scala 50:57:@6492.4]
  wire [10:0] _T_59854; // @[Modules.scala 50:57:@6493.4]
  wire [10:0] buffer_1_526; // @[Modules.scala 50:57:@6494.4]
  wire [10:0] buffer_1_270; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_271; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59856; // @[Modules.scala 50:57:@6496.4]
  wire [10:0] _T_59857; // @[Modules.scala 50:57:@6497.4]
  wire [10:0] buffer_1_527; // @[Modules.scala 50:57:@6498.4]
  wire [10:0] buffer_1_272; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59859; // @[Modules.scala 50:57:@6500.4]
  wire [10:0] _T_59860; // @[Modules.scala 50:57:@6501.4]
  wire [10:0] buffer_1_528; // @[Modules.scala 50:57:@6502.4]
  wire [10:0] buffer_1_274; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59862; // @[Modules.scala 50:57:@6504.4]
  wire [10:0] _T_59863; // @[Modules.scala 50:57:@6505.4]
  wire [10:0] buffer_1_529; // @[Modules.scala 50:57:@6506.4]
  wire [10:0] buffer_1_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59865; // @[Modules.scala 50:57:@6508.4]
  wire [10:0] _T_59866; // @[Modules.scala 50:57:@6509.4]
  wire [10:0] buffer_1_530; // @[Modules.scala 50:57:@6510.4]
  wire [10:0] buffer_1_278; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59868; // @[Modules.scala 50:57:@6512.4]
  wire [10:0] _T_59869; // @[Modules.scala 50:57:@6513.4]
  wire [10:0] buffer_1_531; // @[Modules.scala 50:57:@6514.4]
  wire [10:0] buffer_1_280; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59871; // @[Modules.scala 50:57:@6516.4]
  wire [10:0] _T_59872; // @[Modules.scala 50:57:@6517.4]
  wire [10:0] buffer_1_532; // @[Modules.scala 50:57:@6518.4]
  wire [10:0] buffer_1_282; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59874; // @[Modules.scala 50:57:@6520.4]
  wire [10:0] _T_59875; // @[Modules.scala 50:57:@6521.4]
  wire [10:0] buffer_1_533; // @[Modules.scala 50:57:@6522.4]
  wire [10:0] buffer_1_284; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_285; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59877; // @[Modules.scala 50:57:@6524.4]
  wire [10:0] _T_59878; // @[Modules.scala 50:57:@6525.4]
  wire [10:0] buffer_1_534; // @[Modules.scala 50:57:@6526.4]
  wire [10:0] buffer_1_286; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59880; // @[Modules.scala 50:57:@6528.4]
  wire [10:0] _T_59881; // @[Modules.scala 50:57:@6529.4]
  wire [10:0] buffer_1_535; // @[Modules.scala 50:57:@6530.4]
  wire [10:0] buffer_1_288; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59883; // @[Modules.scala 50:57:@6532.4]
  wire [10:0] _T_59884; // @[Modules.scala 50:57:@6533.4]
  wire [10:0] buffer_1_536; // @[Modules.scala 50:57:@6534.4]
  wire [10:0] buffer_1_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59886; // @[Modules.scala 50:57:@6536.4]
  wire [10:0] _T_59887; // @[Modules.scala 50:57:@6537.4]
  wire [10:0] buffer_1_537; // @[Modules.scala 50:57:@6538.4]
  wire [10:0] buffer_1_292; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59889; // @[Modules.scala 50:57:@6540.4]
  wire [10:0] _T_59890; // @[Modules.scala 50:57:@6541.4]
  wire [10:0] buffer_1_538; // @[Modules.scala 50:57:@6542.4]
  wire [10:0] buffer_1_294; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_295; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59892; // @[Modules.scala 50:57:@6544.4]
  wire [10:0] _T_59893; // @[Modules.scala 50:57:@6545.4]
  wire [10:0] buffer_1_539; // @[Modules.scala 50:57:@6546.4]
  wire [10:0] buffer_1_296; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59895; // @[Modules.scala 50:57:@6548.4]
  wire [10:0] _T_59896; // @[Modules.scala 50:57:@6549.4]
  wire [10:0] buffer_1_540; // @[Modules.scala 50:57:@6550.4]
  wire [10:0] buffer_1_298; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59898; // @[Modules.scala 50:57:@6552.4]
  wire [10:0] _T_59899; // @[Modules.scala 50:57:@6553.4]
  wire [10:0] buffer_1_541; // @[Modules.scala 50:57:@6554.4]
  wire [10:0] buffer_1_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59901; // @[Modules.scala 50:57:@6556.4]
  wire [10:0] _T_59902; // @[Modules.scala 50:57:@6557.4]
  wire [10:0] buffer_1_542; // @[Modules.scala 50:57:@6558.4]
  wire [10:0] buffer_1_306; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59910; // @[Modules.scala 50:57:@6568.4]
  wire [10:0] _T_59911; // @[Modules.scala 50:57:@6569.4]
  wire [10:0] buffer_1_545; // @[Modules.scala 50:57:@6570.4]
  wire [10:0] buffer_1_308; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59913; // @[Modules.scala 50:57:@6572.4]
  wire [10:0] _T_59914; // @[Modules.scala 50:57:@6573.4]
  wire [10:0] buffer_1_546; // @[Modules.scala 50:57:@6574.4]
  wire [10:0] buffer_1_310; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59916; // @[Modules.scala 50:57:@6576.4]
  wire [10:0] _T_59917; // @[Modules.scala 50:57:@6577.4]
  wire [10:0] buffer_1_547; // @[Modules.scala 50:57:@6578.4]
  wire [10:0] buffer_1_312; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59919; // @[Modules.scala 50:57:@6580.4]
  wire [10:0] _T_59920; // @[Modules.scala 50:57:@6581.4]
  wire [10:0] buffer_1_548; // @[Modules.scala 50:57:@6582.4]
  wire [10:0] buffer_1_314; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59922; // @[Modules.scala 50:57:@6584.4]
  wire [10:0] _T_59923; // @[Modules.scala 50:57:@6585.4]
  wire [10:0] buffer_1_549; // @[Modules.scala 50:57:@6586.4]
  wire [10:0] buffer_1_316; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59925; // @[Modules.scala 50:57:@6588.4]
  wire [10:0] _T_59926; // @[Modules.scala 50:57:@6589.4]
  wire [10:0] buffer_1_550; // @[Modules.scala 50:57:@6590.4]
  wire [10:0] buffer_1_318; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59928; // @[Modules.scala 50:57:@6592.4]
  wire [10:0] _T_59929; // @[Modules.scala 50:57:@6593.4]
  wire [10:0] buffer_1_551; // @[Modules.scala 50:57:@6594.4]
  wire [10:0] buffer_1_320; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59931; // @[Modules.scala 50:57:@6596.4]
  wire [10:0] _T_59932; // @[Modules.scala 50:57:@6597.4]
  wire [10:0] buffer_1_552; // @[Modules.scala 50:57:@6598.4]
  wire [10:0] buffer_1_322; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59934; // @[Modules.scala 50:57:@6600.4]
  wire [10:0] _T_59935; // @[Modules.scala 50:57:@6601.4]
  wire [10:0] buffer_1_553; // @[Modules.scala 50:57:@6602.4]
  wire [10:0] buffer_1_324; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59937; // @[Modules.scala 50:57:@6604.4]
  wire [10:0] _T_59938; // @[Modules.scala 50:57:@6605.4]
  wire [10:0] buffer_1_554; // @[Modules.scala 50:57:@6606.4]
  wire [10:0] buffer_1_326; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59940; // @[Modules.scala 50:57:@6608.4]
  wire [10:0] _T_59941; // @[Modules.scala 50:57:@6609.4]
  wire [10:0] buffer_1_555; // @[Modules.scala 50:57:@6610.4]
  wire [10:0] buffer_1_328; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59943; // @[Modules.scala 50:57:@6612.4]
  wire [10:0] _T_59944; // @[Modules.scala 50:57:@6613.4]
  wire [10:0] buffer_1_556; // @[Modules.scala 50:57:@6614.4]
  wire [10:0] buffer_1_331; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59946; // @[Modules.scala 50:57:@6616.4]
  wire [10:0] _T_59947; // @[Modules.scala 50:57:@6617.4]
  wire [10:0] buffer_1_557; // @[Modules.scala 50:57:@6618.4]
  wire [10:0] buffer_1_332; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_333; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59949; // @[Modules.scala 50:57:@6620.4]
  wire [10:0] _T_59950; // @[Modules.scala 50:57:@6621.4]
  wire [10:0] buffer_1_558; // @[Modules.scala 50:57:@6622.4]
  wire [10:0] buffer_1_334; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59952; // @[Modules.scala 50:57:@6624.4]
  wire [10:0] _T_59953; // @[Modules.scala 50:57:@6625.4]
  wire [10:0] buffer_1_559; // @[Modules.scala 50:57:@6626.4]
  wire [10:0] buffer_1_336; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59955; // @[Modules.scala 50:57:@6628.4]
  wire [10:0] _T_59956; // @[Modules.scala 50:57:@6629.4]
  wire [10:0] buffer_1_560; // @[Modules.scala 50:57:@6630.4]
  wire [10:0] buffer_1_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59961; // @[Modules.scala 50:57:@6636.4]
  wire [10:0] _T_59962; // @[Modules.scala 50:57:@6637.4]
  wire [10:0] buffer_1_562; // @[Modules.scala 50:57:@6638.4]
  wire [10:0] buffer_1_342; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59964; // @[Modules.scala 50:57:@6640.4]
  wire [10:0] _T_59965; // @[Modules.scala 50:57:@6641.4]
  wire [10:0] buffer_1_563; // @[Modules.scala 50:57:@6642.4]
  wire [10:0] buffer_1_344; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59967; // @[Modules.scala 50:57:@6644.4]
  wire [10:0] _T_59968; // @[Modules.scala 50:57:@6645.4]
  wire [10:0] buffer_1_564; // @[Modules.scala 50:57:@6646.4]
  wire [10:0] buffer_1_346; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59970; // @[Modules.scala 50:57:@6648.4]
  wire [10:0] _T_59971; // @[Modules.scala 50:57:@6649.4]
  wire [10:0] buffer_1_565; // @[Modules.scala 50:57:@6650.4]
  wire [10:0] buffer_1_348; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59973; // @[Modules.scala 50:57:@6652.4]
  wire [10:0] _T_59974; // @[Modules.scala 50:57:@6653.4]
  wire [10:0] buffer_1_566; // @[Modules.scala 50:57:@6654.4]
  wire [10:0] buffer_1_350; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59976; // @[Modules.scala 50:57:@6656.4]
  wire [10:0] _T_59977; // @[Modules.scala 50:57:@6657.4]
  wire [10:0] buffer_1_567; // @[Modules.scala 50:57:@6658.4]
  wire [10:0] buffer_1_354; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59982; // @[Modules.scala 50:57:@6664.4]
  wire [10:0] _T_59983; // @[Modules.scala 50:57:@6665.4]
  wire [10:0] buffer_1_569; // @[Modules.scala 50:57:@6666.4]
  wire [10:0] buffer_1_356; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59985; // @[Modules.scala 50:57:@6668.4]
  wire [10:0] _T_59986; // @[Modules.scala 50:57:@6669.4]
  wire [10:0] buffer_1_570; // @[Modules.scala 50:57:@6670.4]
  wire [10:0] buffer_1_358; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_359; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59988; // @[Modules.scala 50:57:@6672.4]
  wire [10:0] _T_59989; // @[Modules.scala 50:57:@6673.4]
  wire [10:0] buffer_1_571; // @[Modules.scala 50:57:@6674.4]
  wire [10:0] buffer_1_360; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59991; // @[Modules.scala 50:57:@6676.4]
  wire [10:0] _T_59992; // @[Modules.scala 50:57:@6677.4]
  wire [10:0] buffer_1_572; // @[Modules.scala 50:57:@6678.4]
  wire [10:0] buffer_1_362; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59994; // @[Modules.scala 50:57:@6680.4]
  wire [10:0] _T_59995; // @[Modules.scala 50:57:@6681.4]
  wire [10:0] buffer_1_573; // @[Modules.scala 50:57:@6682.4]
  wire [10:0] buffer_1_364; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_59997; // @[Modules.scala 50:57:@6684.4]
  wire [10:0] _T_59998; // @[Modules.scala 50:57:@6685.4]
  wire [10:0] buffer_1_574; // @[Modules.scala 50:57:@6686.4]
  wire [10:0] buffer_1_366; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60000; // @[Modules.scala 50:57:@6688.4]
  wire [10:0] _T_60001; // @[Modules.scala 50:57:@6689.4]
  wire [10:0] buffer_1_575; // @[Modules.scala 50:57:@6690.4]
  wire [10:0] buffer_1_370; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60006; // @[Modules.scala 50:57:@6696.4]
  wire [10:0] _T_60007; // @[Modules.scala 50:57:@6697.4]
  wire [10:0] buffer_1_577; // @[Modules.scala 50:57:@6698.4]
  wire [10:0] buffer_1_378; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60018; // @[Modules.scala 50:57:@6712.4]
  wire [10:0] _T_60019; // @[Modules.scala 50:57:@6713.4]
  wire [10:0] buffer_1_581; // @[Modules.scala 50:57:@6714.4]
  wire [10:0] buffer_1_380; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_381; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60021; // @[Modules.scala 50:57:@6716.4]
  wire [10:0] _T_60022; // @[Modules.scala 50:57:@6717.4]
  wire [10:0] buffer_1_582; // @[Modules.scala 50:57:@6718.4]
  wire [10:0] buffer_1_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60024; // @[Modules.scala 50:57:@6720.4]
  wire [10:0] _T_60025; // @[Modules.scala 50:57:@6721.4]
  wire [10:0] buffer_1_583; // @[Modules.scala 50:57:@6722.4]
  wire [10:0] buffer_1_384; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_385; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60027; // @[Modules.scala 50:57:@6724.4]
  wire [10:0] _T_60028; // @[Modules.scala 50:57:@6725.4]
  wire [10:0] buffer_1_584; // @[Modules.scala 50:57:@6726.4]
  wire [10:0] buffer_1_388; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60033; // @[Modules.scala 50:57:@6732.4]
  wire [10:0] _T_60034; // @[Modules.scala 50:57:@6733.4]
  wire [10:0] buffer_1_586; // @[Modules.scala 50:57:@6734.4]
  wire [10:0] buffer_1_390; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60036; // @[Modules.scala 50:57:@6736.4]
  wire [10:0] _T_60037; // @[Modules.scala 50:57:@6737.4]
  wire [10:0] buffer_1_587; // @[Modules.scala 50:57:@6738.4]
  wire [11:0] _T_60039; // @[Modules.scala 53:83:@6740.4]
  wire [10:0] _T_60040; // @[Modules.scala 53:83:@6741.4]
  wire [10:0] buffer_1_588; // @[Modules.scala 53:83:@6742.4]
  wire [11:0] _T_60042; // @[Modules.scala 53:83:@6744.4]
  wire [10:0] _T_60043; // @[Modules.scala 53:83:@6745.4]
  wire [10:0] buffer_1_589; // @[Modules.scala 53:83:@6746.4]
  wire [11:0] _T_60045; // @[Modules.scala 53:83:@6748.4]
  wire [10:0] _T_60046; // @[Modules.scala 53:83:@6749.4]
  wire [10:0] buffer_1_590; // @[Modules.scala 53:83:@6750.4]
  wire [11:0] _T_60048; // @[Modules.scala 53:83:@6752.4]
  wire [10:0] _T_60049; // @[Modules.scala 53:83:@6753.4]
  wire [10:0] buffer_1_591; // @[Modules.scala 53:83:@6754.4]
  wire [11:0] _T_60051; // @[Modules.scala 53:83:@6756.4]
  wire [10:0] _T_60052; // @[Modules.scala 53:83:@6757.4]
  wire [10:0] buffer_1_592; // @[Modules.scala 53:83:@6758.4]
  wire [11:0] _T_60054; // @[Modules.scala 53:83:@6760.4]
  wire [10:0] _T_60055; // @[Modules.scala 53:83:@6761.4]
  wire [10:0] buffer_1_593; // @[Modules.scala 53:83:@6762.4]
  wire [11:0] _T_60057; // @[Modules.scala 53:83:@6764.4]
  wire [10:0] _T_60058; // @[Modules.scala 53:83:@6765.4]
  wire [10:0] buffer_1_594; // @[Modules.scala 53:83:@6766.4]
  wire [11:0] _T_60060; // @[Modules.scala 53:83:@6768.4]
  wire [10:0] _T_60061; // @[Modules.scala 53:83:@6769.4]
  wire [10:0] buffer_1_595; // @[Modules.scala 53:83:@6770.4]
  wire [11:0] _T_60063; // @[Modules.scala 53:83:@6772.4]
  wire [10:0] _T_60064; // @[Modules.scala 53:83:@6773.4]
  wire [10:0] buffer_1_596; // @[Modules.scala 53:83:@6774.4]
  wire [11:0] _T_60066; // @[Modules.scala 53:83:@6776.4]
  wire [10:0] _T_60067; // @[Modules.scala 53:83:@6777.4]
  wire [10:0] buffer_1_597; // @[Modules.scala 53:83:@6778.4]
  wire [11:0] _T_60069; // @[Modules.scala 53:83:@6780.4]
  wire [10:0] _T_60070; // @[Modules.scala 53:83:@6781.4]
  wire [10:0] buffer_1_598; // @[Modules.scala 53:83:@6782.4]
  wire [11:0] _T_60072; // @[Modules.scala 53:83:@6784.4]
  wire [10:0] _T_60073; // @[Modules.scala 53:83:@6785.4]
  wire [10:0] buffer_1_599; // @[Modules.scala 53:83:@6786.4]
  wire [11:0] _T_60075; // @[Modules.scala 53:83:@6788.4]
  wire [10:0] _T_60076; // @[Modules.scala 53:83:@6789.4]
  wire [10:0] buffer_1_600; // @[Modules.scala 53:83:@6790.4]
  wire [11:0] _T_60078; // @[Modules.scala 53:83:@6792.4]
  wire [10:0] _T_60079; // @[Modules.scala 53:83:@6793.4]
  wire [10:0] buffer_1_601; // @[Modules.scala 53:83:@6794.4]
  wire [11:0] _T_60081; // @[Modules.scala 53:83:@6796.4]
  wire [10:0] _T_60082; // @[Modules.scala 53:83:@6797.4]
  wire [10:0] buffer_1_602; // @[Modules.scala 53:83:@6798.4]
  wire [11:0] _T_60084; // @[Modules.scala 53:83:@6800.4]
  wire [10:0] _T_60085; // @[Modules.scala 53:83:@6801.4]
  wire [10:0] buffer_1_603; // @[Modules.scala 53:83:@6802.4]
  wire [11:0] _T_60087; // @[Modules.scala 53:83:@6804.4]
  wire [10:0] _T_60088; // @[Modules.scala 53:83:@6805.4]
  wire [10:0] buffer_1_604; // @[Modules.scala 53:83:@6806.4]
  wire [11:0] _T_60090; // @[Modules.scala 53:83:@6808.4]
  wire [10:0] _T_60091; // @[Modules.scala 53:83:@6809.4]
  wire [10:0] buffer_1_605; // @[Modules.scala 53:83:@6810.4]
  wire [11:0] _T_60093; // @[Modules.scala 53:83:@6812.4]
  wire [10:0] _T_60094; // @[Modules.scala 53:83:@6813.4]
  wire [10:0] buffer_1_606; // @[Modules.scala 53:83:@6814.4]
  wire [11:0] _T_60096; // @[Modules.scala 53:83:@6816.4]
  wire [10:0] _T_60097; // @[Modules.scala 53:83:@6817.4]
  wire [10:0] buffer_1_607; // @[Modules.scala 53:83:@6818.4]
  wire [11:0] _T_60099; // @[Modules.scala 53:83:@6820.4]
  wire [10:0] _T_60100; // @[Modules.scala 53:83:@6821.4]
  wire [10:0] buffer_1_608; // @[Modules.scala 53:83:@6822.4]
  wire [11:0] _T_60102; // @[Modules.scala 53:83:@6824.4]
  wire [10:0] _T_60103; // @[Modules.scala 53:83:@6825.4]
  wire [10:0] buffer_1_609; // @[Modules.scala 53:83:@6826.4]
  wire [11:0] _T_60105; // @[Modules.scala 53:83:@6828.4]
  wire [10:0] _T_60106; // @[Modules.scala 53:83:@6829.4]
  wire [10:0] buffer_1_610; // @[Modules.scala 53:83:@6830.4]
  wire [11:0] _T_60108; // @[Modules.scala 53:83:@6832.4]
  wire [10:0] _T_60109; // @[Modules.scala 53:83:@6833.4]
  wire [10:0] buffer_1_611; // @[Modules.scala 53:83:@6834.4]
  wire [11:0] _T_60111; // @[Modules.scala 53:83:@6836.4]
  wire [10:0] _T_60112; // @[Modules.scala 53:83:@6837.4]
  wire [10:0] buffer_1_612; // @[Modules.scala 53:83:@6838.4]
  wire [11:0] _T_60114; // @[Modules.scala 53:83:@6840.4]
  wire [10:0] _T_60115; // @[Modules.scala 53:83:@6841.4]
  wire [10:0] buffer_1_613; // @[Modules.scala 53:83:@6842.4]
  wire [11:0] _T_60117; // @[Modules.scala 53:83:@6844.4]
  wire [10:0] _T_60118; // @[Modules.scala 53:83:@6845.4]
  wire [10:0] buffer_1_614; // @[Modules.scala 53:83:@6846.4]
  wire [11:0] _T_60120; // @[Modules.scala 53:83:@6848.4]
  wire [10:0] _T_60121; // @[Modules.scala 53:83:@6849.4]
  wire [10:0] buffer_1_615; // @[Modules.scala 53:83:@6850.4]
  wire [11:0] _T_60123; // @[Modules.scala 53:83:@6852.4]
  wire [10:0] _T_60124; // @[Modules.scala 53:83:@6853.4]
  wire [10:0] buffer_1_616; // @[Modules.scala 53:83:@6854.4]
  wire [11:0] _T_60126; // @[Modules.scala 53:83:@6856.4]
  wire [10:0] _T_60127; // @[Modules.scala 53:83:@6857.4]
  wire [10:0] buffer_1_617; // @[Modules.scala 53:83:@6858.4]
  wire [11:0] _T_60129; // @[Modules.scala 53:83:@6860.4]
  wire [10:0] _T_60130; // @[Modules.scala 53:83:@6861.4]
  wire [10:0] buffer_1_618; // @[Modules.scala 53:83:@6862.4]
  wire [11:0] _T_60132; // @[Modules.scala 53:83:@6864.4]
  wire [10:0] _T_60133; // @[Modules.scala 53:83:@6865.4]
  wire [10:0] buffer_1_619; // @[Modules.scala 53:83:@6866.4]
  wire [11:0] _T_60135; // @[Modules.scala 53:83:@6868.4]
  wire [10:0] _T_60136; // @[Modules.scala 53:83:@6869.4]
  wire [10:0] buffer_1_620; // @[Modules.scala 53:83:@6870.4]
  wire [11:0] _T_60138; // @[Modules.scala 53:83:@6872.4]
  wire [10:0] _T_60139; // @[Modules.scala 53:83:@6873.4]
  wire [10:0] buffer_1_621; // @[Modules.scala 53:83:@6874.4]
  wire [11:0] _T_60141; // @[Modules.scala 53:83:@6876.4]
  wire [10:0] _T_60142; // @[Modules.scala 53:83:@6877.4]
  wire [10:0] buffer_1_622; // @[Modules.scala 53:83:@6878.4]
  wire [11:0] _T_60144; // @[Modules.scala 53:83:@6880.4]
  wire [10:0] _T_60145; // @[Modules.scala 53:83:@6881.4]
  wire [10:0] buffer_1_623; // @[Modules.scala 53:83:@6882.4]
  wire [11:0] _T_60147; // @[Modules.scala 53:83:@6884.4]
  wire [10:0] _T_60148; // @[Modules.scala 53:83:@6885.4]
  wire [10:0] buffer_1_624; // @[Modules.scala 53:83:@6886.4]
  wire [11:0] _T_60150; // @[Modules.scala 53:83:@6888.4]
  wire [10:0] _T_60151; // @[Modules.scala 53:83:@6889.4]
  wire [10:0] buffer_1_625; // @[Modules.scala 53:83:@6890.4]
  wire [11:0] _T_60153; // @[Modules.scala 53:83:@6892.4]
  wire [10:0] _T_60154; // @[Modules.scala 53:83:@6893.4]
  wire [10:0] buffer_1_626; // @[Modules.scala 53:83:@6894.4]
  wire [11:0] _T_60156; // @[Modules.scala 53:83:@6896.4]
  wire [10:0] _T_60157; // @[Modules.scala 53:83:@6897.4]
  wire [10:0] buffer_1_627; // @[Modules.scala 53:83:@6898.4]
  wire [11:0] _T_60159; // @[Modules.scala 53:83:@6900.4]
  wire [10:0] _T_60160; // @[Modules.scala 53:83:@6901.4]
  wire [10:0] buffer_1_628; // @[Modules.scala 53:83:@6902.4]
  wire [11:0] _T_60162; // @[Modules.scala 53:83:@6904.4]
  wire [10:0] _T_60163; // @[Modules.scala 53:83:@6905.4]
  wire [10:0] buffer_1_629; // @[Modules.scala 53:83:@6906.4]
  wire [11:0] _T_60168; // @[Modules.scala 53:83:@6912.4]
  wire [10:0] _T_60169; // @[Modules.scala 53:83:@6913.4]
  wire [10:0] buffer_1_631; // @[Modules.scala 53:83:@6914.4]
  wire [11:0] _T_60171; // @[Modules.scala 53:83:@6916.4]
  wire [10:0] _T_60172; // @[Modules.scala 53:83:@6917.4]
  wire [10:0] buffer_1_632; // @[Modules.scala 53:83:@6918.4]
  wire [11:0] _T_60174; // @[Modules.scala 53:83:@6920.4]
  wire [10:0] _T_60175; // @[Modules.scala 53:83:@6921.4]
  wire [10:0] buffer_1_633; // @[Modules.scala 53:83:@6922.4]
  wire [11:0] _T_60177; // @[Modules.scala 53:83:@6924.4]
  wire [10:0] _T_60178; // @[Modules.scala 53:83:@6925.4]
  wire [10:0] buffer_1_634; // @[Modules.scala 53:83:@6926.4]
  wire [11:0] _T_60180; // @[Modules.scala 53:83:@6928.4]
  wire [10:0] _T_60181; // @[Modules.scala 53:83:@6929.4]
  wire [10:0] buffer_1_635; // @[Modules.scala 53:83:@6930.4]
  wire [11:0] _T_60183; // @[Modules.scala 53:83:@6932.4]
  wire [10:0] _T_60184; // @[Modules.scala 53:83:@6933.4]
  wire [10:0] buffer_1_636; // @[Modules.scala 53:83:@6934.4]
  wire [11:0] _T_60186; // @[Modules.scala 53:83:@6936.4]
  wire [10:0] _T_60187; // @[Modules.scala 53:83:@6937.4]
  wire [10:0] buffer_1_637; // @[Modules.scala 53:83:@6938.4]
  wire [11:0] _T_60189; // @[Modules.scala 53:83:@6940.4]
  wire [10:0] _T_60190; // @[Modules.scala 53:83:@6941.4]
  wire [10:0] buffer_1_638; // @[Modules.scala 53:83:@6942.4]
  wire [11:0] _T_60192; // @[Modules.scala 53:83:@6944.4]
  wire [10:0] _T_60193; // @[Modules.scala 53:83:@6945.4]
  wire [10:0] buffer_1_639; // @[Modules.scala 53:83:@6946.4]
  wire [11:0] _T_60195; // @[Modules.scala 53:83:@6948.4]
  wire [10:0] _T_60196; // @[Modules.scala 53:83:@6949.4]
  wire [10:0] buffer_1_640; // @[Modules.scala 53:83:@6950.4]
  wire [11:0] _T_60198; // @[Modules.scala 53:83:@6952.4]
  wire [10:0] _T_60199; // @[Modules.scala 53:83:@6953.4]
  wire [10:0] buffer_1_641; // @[Modules.scala 53:83:@6954.4]
  wire [11:0] _T_60201; // @[Modules.scala 53:83:@6956.4]
  wire [10:0] _T_60202; // @[Modules.scala 53:83:@6957.4]
  wire [10:0] buffer_1_642; // @[Modules.scala 53:83:@6958.4]
  wire [11:0] _T_60204; // @[Modules.scala 53:83:@6960.4]
  wire [10:0] _T_60205; // @[Modules.scala 53:83:@6961.4]
  wire [10:0] buffer_1_643; // @[Modules.scala 53:83:@6962.4]
  wire [11:0] _T_60207; // @[Modules.scala 53:83:@6964.4]
  wire [10:0] _T_60208; // @[Modules.scala 53:83:@6965.4]
  wire [10:0] buffer_1_644; // @[Modules.scala 53:83:@6966.4]
  wire [11:0] _T_60210; // @[Modules.scala 53:83:@6968.4]
  wire [10:0] _T_60211; // @[Modules.scala 53:83:@6969.4]
  wire [10:0] buffer_1_645; // @[Modules.scala 53:83:@6970.4]
  wire [11:0] _T_60213; // @[Modules.scala 53:83:@6972.4]
  wire [10:0] _T_60214; // @[Modules.scala 53:83:@6973.4]
  wire [10:0] buffer_1_646; // @[Modules.scala 53:83:@6974.4]
  wire [11:0] _T_60216; // @[Modules.scala 53:83:@6976.4]
  wire [10:0] _T_60217; // @[Modules.scala 53:83:@6977.4]
  wire [10:0] buffer_1_647; // @[Modules.scala 53:83:@6978.4]
  wire [11:0] _T_60219; // @[Modules.scala 53:83:@6980.4]
  wire [10:0] _T_60220; // @[Modules.scala 53:83:@6981.4]
  wire [10:0] buffer_1_648; // @[Modules.scala 53:83:@6982.4]
  wire [11:0] _T_60222; // @[Modules.scala 53:83:@6984.4]
  wire [10:0] _T_60223; // @[Modules.scala 53:83:@6985.4]
  wire [10:0] buffer_1_649; // @[Modules.scala 53:83:@6986.4]
  wire [11:0] _T_60225; // @[Modules.scala 53:83:@6988.4]
  wire [10:0] _T_60226; // @[Modules.scala 53:83:@6989.4]
  wire [10:0] buffer_1_650; // @[Modules.scala 53:83:@6990.4]
  wire [11:0] _T_60228; // @[Modules.scala 53:83:@6992.4]
  wire [10:0] _T_60229; // @[Modules.scala 53:83:@6993.4]
  wire [10:0] buffer_1_651; // @[Modules.scala 53:83:@6994.4]
  wire [11:0] _T_60231; // @[Modules.scala 53:83:@6996.4]
  wire [10:0] _T_60232; // @[Modules.scala 53:83:@6997.4]
  wire [10:0] buffer_1_652; // @[Modules.scala 53:83:@6998.4]
  wire [11:0] _T_60234; // @[Modules.scala 53:83:@7000.4]
  wire [10:0] _T_60235; // @[Modules.scala 53:83:@7001.4]
  wire [10:0] buffer_1_653; // @[Modules.scala 53:83:@7002.4]
  wire [11:0] _T_60237; // @[Modules.scala 53:83:@7004.4]
  wire [10:0] _T_60238; // @[Modules.scala 53:83:@7005.4]
  wire [10:0] buffer_1_654; // @[Modules.scala 53:83:@7006.4]
  wire [11:0] _T_60240; // @[Modules.scala 53:83:@7008.4]
  wire [10:0] _T_60241; // @[Modules.scala 53:83:@7009.4]
  wire [10:0] buffer_1_655; // @[Modules.scala 53:83:@7010.4]
  wire [11:0] _T_60243; // @[Modules.scala 53:83:@7012.4]
  wire [10:0] _T_60244; // @[Modules.scala 53:83:@7013.4]
  wire [10:0] buffer_1_656; // @[Modules.scala 53:83:@7014.4]
  wire [11:0] _T_60246; // @[Modules.scala 53:83:@7016.4]
  wire [10:0] _T_60247; // @[Modules.scala 53:83:@7017.4]
  wire [10:0] buffer_1_657; // @[Modules.scala 53:83:@7018.4]
  wire [11:0] _T_60249; // @[Modules.scala 53:83:@7020.4]
  wire [10:0] _T_60250; // @[Modules.scala 53:83:@7021.4]
  wire [10:0] buffer_1_658; // @[Modules.scala 53:83:@7022.4]
  wire [11:0] _T_60252; // @[Modules.scala 53:83:@7024.4]
  wire [10:0] _T_60253; // @[Modules.scala 53:83:@7025.4]
  wire [10:0] buffer_1_659; // @[Modules.scala 53:83:@7026.4]
  wire [11:0] _T_60255; // @[Modules.scala 53:83:@7028.4]
  wire [10:0] _T_60256; // @[Modules.scala 53:83:@7029.4]
  wire [10:0] buffer_1_660; // @[Modules.scala 53:83:@7030.4]
  wire [11:0] _T_60258; // @[Modules.scala 53:83:@7032.4]
  wire [10:0] _T_60259; // @[Modules.scala 53:83:@7033.4]
  wire [10:0] buffer_1_661; // @[Modules.scala 53:83:@7034.4]
  wire [11:0] _T_60261; // @[Modules.scala 53:83:@7036.4]
  wire [10:0] _T_60262; // @[Modules.scala 53:83:@7037.4]
  wire [10:0] buffer_1_662; // @[Modules.scala 53:83:@7038.4]
  wire [11:0] _T_60264; // @[Modules.scala 53:83:@7040.4]
  wire [10:0] _T_60265; // @[Modules.scala 53:83:@7041.4]
  wire [10:0] buffer_1_663; // @[Modules.scala 53:83:@7042.4]
  wire [11:0] _T_60267; // @[Modules.scala 53:83:@7044.4]
  wire [10:0] _T_60268; // @[Modules.scala 53:83:@7045.4]
  wire [10:0] buffer_1_664; // @[Modules.scala 53:83:@7046.4]
  wire [11:0] _T_60270; // @[Modules.scala 53:83:@7048.4]
  wire [10:0] _T_60271; // @[Modules.scala 53:83:@7049.4]
  wire [10:0] buffer_1_665; // @[Modules.scala 53:83:@7050.4]
  wire [11:0] _T_60273; // @[Modules.scala 53:83:@7052.4]
  wire [10:0] _T_60274; // @[Modules.scala 53:83:@7053.4]
  wire [10:0] buffer_1_666; // @[Modules.scala 53:83:@7054.4]
  wire [11:0] _T_60276; // @[Modules.scala 53:83:@7056.4]
  wire [10:0] _T_60277; // @[Modules.scala 53:83:@7057.4]
  wire [10:0] buffer_1_667; // @[Modules.scala 53:83:@7058.4]
  wire [11:0] _T_60279; // @[Modules.scala 53:83:@7060.4]
  wire [10:0] _T_60280; // @[Modules.scala 53:83:@7061.4]
  wire [10:0] buffer_1_668; // @[Modules.scala 53:83:@7062.4]
  wire [11:0] _T_60282; // @[Modules.scala 53:83:@7064.4]
  wire [10:0] _T_60283; // @[Modules.scala 53:83:@7065.4]
  wire [10:0] buffer_1_669; // @[Modules.scala 53:83:@7066.4]
  wire [11:0] _T_60285; // @[Modules.scala 53:83:@7068.4]
  wire [10:0] _T_60286; // @[Modules.scala 53:83:@7069.4]
  wire [10:0] buffer_1_670; // @[Modules.scala 53:83:@7070.4]
  wire [11:0] _T_60288; // @[Modules.scala 53:83:@7072.4]
  wire [10:0] _T_60289; // @[Modules.scala 53:83:@7073.4]
  wire [10:0] buffer_1_671; // @[Modules.scala 53:83:@7074.4]
  wire [11:0] _T_60291; // @[Modules.scala 53:83:@7076.4]
  wire [10:0] _T_60292; // @[Modules.scala 53:83:@7077.4]
  wire [10:0] buffer_1_672; // @[Modules.scala 53:83:@7078.4]
  wire [11:0] _T_60294; // @[Modules.scala 53:83:@7080.4]
  wire [10:0] _T_60295; // @[Modules.scala 53:83:@7081.4]
  wire [10:0] buffer_1_673; // @[Modules.scala 53:83:@7082.4]
  wire [11:0] _T_60297; // @[Modules.scala 53:83:@7084.4]
  wire [10:0] _T_60298; // @[Modules.scala 53:83:@7085.4]
  wire [10:0] buffer_1_674; // @[Modules.scala 53:83:@7086.4]
  wire [11:0] _T_60300; // @[Modules.scala 53:83:@7088.4]
  wire [10:0] _T_60301; // @[Modules.scala 53:83:@7089.4]
  wire [10:0] buffer_1_675; // @[Modules.scala 53:83:@7090.4]
  wire [11:0] _T_60303; // @[Modules.scala 53:83:@7092.4]
  wire [10:0] _T_60304; // @[Modules.scala 53:83:@7093.4]
  wire [10:0] buffer_1_676; // @[Modules.scala 53:83:@7094.4]
  wire [11:0] _T_60306; // @[Modules.scala 53:83:@7096.4]
  wire [10:0] _T_60307; // @[Modules.scala 53:83:@7097.4]
  wire [10:0] buffer_1_677; // @[Modules.scala 53:83:@7098.4]
  wire [11:0] _T_60309; // @[Modules.scala 53:83:@7100.4]
  wire [10:0] _T_60310; // @[Modules.scala 53:83:@7101.4]
  wire [10:0] buffer_1_678; // @[Modules.scala 53:83:@7102.4]
  wire [11:0] _T_60312; // @[Modules.scala 53:83:@7104.4]
  wire [10:0] _T_60313; // @[Modules.scala 53:83:@7105.4]
  wire [10:0] buffer_1_679; // @[Modules.scala 53:83:@7106.4]
  wire [11:0] _T_60315; // @[Modules.scala 53:83:@7108.4]
  wire [10:0] _T_60316; // @[Modules.scala 53:83:@7109.4]
  wire [10:0] buffer_1_680; // @[Modules.scala 53:83:@7110.4]
  wire [11:0] _T_60321; // @[Modules.scala 53:83:@7116.4]
  wire [10:0] _T_60322; // @[Modules.scala 53:83:@7117.4]
  wire [10:0] buffer_1_682; // @[Modules.scala 53:83:@7118.4]
  wire [11:0] _T_60324; // @[Modules.scala 53:83:@7120.4]
  wire [10:0] _T_60325; // @[Modules.scala 53:83:@7121.4]
  wire [10:0] buffer_1_683; // @[Modules.scala 53:83:@7122.4]
  wire [11:0] _T_60327; // @[Modules.scala 53:83:@7124.4]
  wire [10:0] _T_60328; // @[Modules.scala 53:83:@7125.4]
  wire [10:0] buffer_1_684; // @[Modules.scala 53:83:@7126.4]
  wire [11:0] _T_60330; // @[Modules.scala 53:83:@7128.4]
  wire [10:0] _T_60331; // @[Modules.scala 53:83:@7129.4]
  wire [10:0] buffer_1_685; // @[Modules.scala 53:83:@7130.4]
  wire [11:0] _T_60333; // @[Modules.scala 56:109:@7132.4]
  wire [10:0] _T_60334; // @[Modules.scala 56:109:@7133.4]
  wire [10:0] buffer_1_686; // @[Modules.scala 56:109:@7134.4]
  wire [11:0] _T_60336; // @[Modules.scala 56:109:@7136.4]
  wire [10:0] _T_60337; // @[Modules.scala 56:109:@7137.4]
  wire [10:0] buffer_1_687; // @[Modules.scala 56:109:@7138.4]
  wire [11:0] _T_60339; // @[Modules.scala 56:109:@7140.4]
  wire [10:0] _T_60340; // @[Modules.scala 56:109:@7141.4]
  wire [10:0] buffer_1_688; // @[Modules.scala 56:109:@7142.4]
  wire [11:0] _T_60342; // @[Modules.scala 56:109:@7144.4]
  wire [10:0] _T_60343; // @[Modules.scala 56:109:@7145.4]
  wire [10:0] buffer_1_689; // @[Modules.scala 56:109:@7146.4]
  wire [11:0] _T_60345; // @[Modules.scala 56:109:@7148.4]
  wire [10:0] _T_60346; // @[Modules.scala 56:109:@7149.4]
  wire [10:0] buffer_1_690; // @[Modules.scala 56:109:@7150.4]
  wire [11:0] _T_60348; // @[Modules.scala 56:109:@7152.4]
  wire [10:0] _T_60349; // @[Modules.scala 56:109:@7153.4]
  wire [10:0] buffer_1_691; // @[Modules.scala 56:109:@7154.4]
  wire [11:0] _T_60351; // @[Modules.scala 56:109:@7156.4]
  wire [10:0] _T_60352; // @[Modules.scala 56:109:@7157.4]
  wire [10:0] buffer_1_692; // @[Modules.scala 56:109:@7158.4]
  wire [11:0] _T_60354; // @[Modules.scala 56:109:@7160.4]
  wire [10:0] _T_60355; // @[Modules.scala 56:109:@7161.4]
  wire [10:0] buffer_1_693; // @[Modules.scala 56:109:@7162.4]
  wire [11:0] _T_60357; // @[Modules.scala 56:109:@7164.4]
  wire [10:0] _T_60358; // @[Modules.scala 56:109:@7165.4]
  wire [10:0] buffer_1_694; // @[Modules.scala 56:109:@7166.4]
  wire [11:0] _T_60360; // @[Modules.scala 56:109:@7168.4]
  wire [10:0] _T_60361; // @[Modules.scala 56:109:@7169.4]
  wire [10:0] buffer_1_695; // @[Modules.scala 56:109:@7170.4]
  wire [11:0] _T_60363; // @[Modules.scala 56:109:@7172.4]
  wire [10:0] _T_60364; // @[Modules.scala 56:109:@7173.4]
  wire [10:0] buffer_1_696; // @[Modules.scala 56:109:@7174.4]
  wire [11:0] _T_60366; // @[Modules.scala 56:109:@7176.4]
  wire [10:0] _T_60367; // @[Modules.scala 56:109:@7177.4]
  wire [10:0] buffer_1_697; // @[Modules.scala 56:109:@7178.4]
  wire [11:0] _T_60369; // @[Modules.scala 56:109:@7180.4]
  wire [10:0] _T_60370; // @[Modules.scala 56:109:@7181.4]
  wire [10:0] buffer_1_698; // @[Modules.scala 56:109:@7182.4]
  wire [11:0] _T_60372; // @[Modules.scala 56:109:@7184.4]
  wire [10:0] _T_60373; // @[Modules.scala 56:109:@7185.4]
  wire [10:0] buffer_1_699; // @[Modules.scala 56:109:@7186.4]
  wire [11:0] _T_60375; // @[Modules.scala 56:109:@7188.4]
  wire [10:0] _T_60376; // @[Modules.scala 56:109:@7189.4]
  wire [10:0] buffer_1_700; // @[Modules.scala 56:109:@7190.4]
  wire [11:0] _T_60378; // @[Modules.scala 56:109:@7192.4]
  wire [10:0] _T_60379; // @[Modules.scala 56:109:@7193.4]
  wire [10:0] buffer_1_701; // @[Modules.scala 56:109:@7194.4]
  wire [11:0] _T_60381; // @[Modules.scala 56:109:@7196.4]
  wire [10:0] _T_60382; // @[Modules.scala 56:109:@7197.4]
  wire [10:0] buffer_1_702; // @[Modules.scala 56:109:@7198.4]
  wire [11:0] _T_60384; // @[Modules.scala 56:109:@7200.4]
  wire [10:0] _T_60385; // @[Modules.scala 56:109:@7201.4]
  wire [10:0] buffer_1_703; // @[Modules.scala 56:109:@7202.4]
  wire [11:0] _T_60387; // @[Modules.scala 56:109:@7204.4]
  wire [10:0] _T_60388; // @[Modules.scala 56:109:@7205.4]
  wire [10:0] buffer_1_704; // @[Modules.scala 56:109:@7206.4]
  wire [11:0] _T_60390; // @[Modules.scala 56:109:@7208.4]
  wire [10:0] _T_60391; // @[Modules.scala 56:109:@7209.4]
  wire [10:0] buffer_1_705; // @[Modules.scala 56:109:@7210.4]
  wire [11:0] _T_60393; // @[Modules.scala 56:109:@7212.4]
  wire [10:0] _T_60394; // @[Modules.scala 56:109:@7213.4]
  wire [10:0] buffer_1_706; // @[Modules.scala 56:109:@7214.4]
  wire [11:0] _T_60396; // @[Modules.scala 56:109:@7216.4]
  wire [10:0] _T_60397; // @[Modules.scala 56:109:@7217.4]
  wire [10:0] buffer_1_707; // @[Modules.scala 56:109:@7218.4]
  wire [11:0] _T_60399; // @[Modules.scala 56:109:@7220.4]
  wire [10:0] _T_60400; // @[Modules.scala 56:109:@7221.4]
  wire [10:0] buffer_1_708; // @[Modules.scala 56:109:@7222.4]
  wire [11:0] _T_60402; // @[Modules.scala 56:109:@7224.4]
  wire [10:0] _T_60403; // @[Modules.scala 56:109:@7225.4]
  wire [10:0] buffer_1_709; // @[Modules.scala 56:109:@7226.4]
  wire [11:0] _T_60405; // @[Modules.scala 56:109:@7228.4]
  wire [10:0] _T_60406; // @[Modules.scala 56:109:@7229.4]
  wire [10:0] buffer_1_710; // @[Modules.scala 56:109:@7230.4]
  wire [11:0] _T_60408; // @[Modules.scala 56:109:@7232.4]
  wire [10:0] _T_60409; // @[Modules.scala 56:109:@7233.4]
  wire [10:0] buffer_1_711; // @[Modules.scala 56:109:@7234.4]
  wire [11:0] _T_60411; // @[Modules.scala 56:109:@7236.4]
  wire [10:0] _T_60412; // @[Modules.scala 56:109:@7237.4]
  wire [10:0] buffer_1_712; // @[Modules.scala 56:109:@7238.4]
  wire [11:0] _T_60414; // @[Modules.scala 56:109:@7240.4]
  wire [10:0] _T_60415; // @[Modules.scala 56:109:@7241.4]
  wire [10:0] buffer_1_713; // @[Modules.scala 56:109:@7242.4]
  wire [11:0] _T_60417; // @[Modules.scala 56:109:@7244.4]
  wire [10:0] _T_60418; // @[Modules.scala 56:109:@7245.4]
  wire [10:0] buffer_1_714; // @[Modules.scala 56:109:@7246.4]
  wire [11:0] _T_60420; // @[Modules.scala 56:109:@7248.4]
  wire [10:0] _T_60421; // @[Modules.scala 56:109:@7249.4]
  wire [10:0] buffer_1_715; // @[Modules.scala 56:109:@7250.4]
  wire [11:0] _T_60423; // @[Modules.scala 56:109:@7252.4]
  wire [10:0] _T_60424; // @[Modules.scala 56:109:@7253.4]
  wire [10:0] buffer_1_716; // @[Modules.scala 56:109:@7254.4]
  wire [11:0] _T_60426; // @[Modules.scala 56:109:@7256.4]
  wire [10:0] _T_60427; // @[Modules.scala 56:109:@7257.4]
  wire [10:0] buffer_1_717; // @[Modules.scala 56:109:@7258.4]
  wire [11:0] _T_60429; // @[Modules.scala 56:109:@7260.4]
  wire [10:0] _T_60430; // @[Modules.scala 56:109:@7261.4]
  wire [10:0] buffer_1_718; // @[Modules.scala 56:109:@7262.4]
  wire [11:0] _T_60432; // @[Modules.scala 56:109:@7264.4]
  wire [10:0] _T_60433; // @[Modules.scala 56:109:@7265.4]
  wire [10:0] buffer_1_719; // @[Modules.scala 56:109:@7266.4]
  wire [11:0] _T_60435; // @[Modules.scala 56:109:@7268.4]
  wire [10:0] _T_60436; // @[Modules.scala 56:109:@7269.4]
  wire [10:0] buffer_1_720; // @[Modules.scala 56:109:@7270.4]
  wire [11:0] _T_60438; // @[Modules.scala 56:109:@7272.4]
  wire [10:0] _T_60439; // @[Modules.scala 56:109:@7273.4]
  wire [10:0] buffer_1_721; // @[Modules.scala 56:109:@7274.4]
  wire [11:0] _T_60441; // @[Modules.scala 56:109:@7276.4]
  wire [10:0] _T_60442; // @[Modules.scala 56:109:@7277.4]
  wire [10:0] buffer_1_722; // @[Modules.scala 56:109:@7278.4]
  wire [11:0] _T_60444; // @[Modules.scala 56:109:@7280.4]
  wire [10:0] _T_60445; // @[Modules.scala 56:109:@7281.4]
  wire [10:0] buffer_1_723; // @[Modules.scala 56:109:@7282.4]
  wire [11:0] _T_60447; // @[Modules.scala 56:109:@7284.4]
  wire [10:0] _T_60448; // @[Modules.scala 56:109:@7285.4]
  wire [10:0] buffer_1_724; // @[Modules.scala 56:109:@7286.4]
  wire [11:0] _T_60450; // @[Modules.scala 56:109:@7288.4]
  wire [10:0] _T_60451; // @[Modules.scala 56:109:@7289.4]
  wire [10:0] buffer_1_725; // @[Modules.scala 56:109:@7290.4]
  wire [11:0] _T_60453; // @[Modules.scala 56:109:@7292.4]
  wire [10:0] _T_60454; // @[Modules.scala 56:109:@7293.4]
  wire [10:0] buffer_1_726; // @[Modules.scala 56:109:@7294.4]
  wire [11:0] _T_60456; // @[Modules.scala 56:109:@7296.4]
  wire [10:0] _T_60457; // @[Modules.scala 56:109:@7297.4]
  wire [10:0] buffer_1_727; // @[Modules.scala 56:109:@7298.4]
  wire [11:0] _T_60459; // @[Modules.scala 56:109:@7300.4]
  wire [10:0] _T_60460; // @[Modules.scala 56:109:@7301.4]
  wire [10:0] buffer_1_728; // @[Modules.scala 56:109:@7302.4]
  wire [11:0] _T_60462; // @[Modules.scala 56:109:@7304.4]
  wire [10:0] _T_60463; // @[Modules.scala 56:109:@7305.4]
  wire [10:0] buffer_1_729; // @[Modules.scala 56:109:@7306.4]
  wire [11:0] _T_60465; // @[Modules.scala 56:109:@7308.4]
  wire [10:0] _T_60466; // @[Modules.scala 56:109:@7309.4]
  wire [10:0] buffer_1_730; // @[Modules.scala 56:109:@7310.4]
  wire [11:0] _T_60468; // @[Modules.scala 56:109:@7312.4]
  wire [10:0] _T_60469; // @[Modules.scala 56:109:@7313.4]
  wire [10:0] buffer_1_731; // @[Modules.scala 56:109:@7314.4]
  wire [11:0] _T_60471; // @[Modules.scala 56:109:@7316.4]
  wire [10:0] _T_60472; // @[Modules.scala 56:109:@7317.4]
  wire [10:0] buffer_1_732; // @[Modules.scala 56:109:@7318.4]
  wire [11:0] _T_60474; // @[Modules.scala 56:109:@7320.4]
  wire [10:0] _T_60475; // @[Modules.scala 56:109:@7321.4]
  wire [10:0] buffer_1_733; // @[Modules.scala 56:109:@7322.4]
  wire [11:0] _T_60477; // @[Modules.scala 56:109:@7324.4]
  wire [10:0] _T_60478; // @[Modules.scala 56:109:@7325.4]
  wire [10:0] buffer_1_734; // @[Modules.scala 56:109:@7326.4]
  wire [11:0] _T_60480; // @[Modules.scala 63:156:@7329.4]
  wire [10:0] _T_60481; // @[Modules.scala 63:156:@7330.4]
  wire [10:0] buffer_1_736; // @[Modules.scala 63:156:@7331.4]
  wire [11:0] _T_60483; // @[Modules.scala 63:156:@7333.4]
  wire [10:0] _T_60484; // @[Modules.scala 63:156:@7334.4]
  wire [10:0] buffer_1_737; // @[Modules.scala 63:156:@7335.4]
  wire [11:0] _T_60486; // @[Modules.scala 63:156:@7337.4]
  wire [10:0] _T_60487; // @[Modules.scala 63:156:@7338.4]
  wire [10:0] buffer_1_738; // @[Modules.scala 63:156:@7339.4]
  wire [11:0] _T_60489; // @[Modules.scala 63:156:@7341.4]
  wire [10:0] _T_60490; // @[Modules.scala 63:156:@7342.4]
  wire [10:0] buffer_1_739; // @[Modules.scala 63:156:@7343.4]
  wire [11:0] _T_60492; // @[Modules.scala 63:156:@7345.4]
  wire [10:0] _T_60493; // @[Modules.scala 63:156:@7346.4]
  wire [10:0] buffer_1_740; // @[Modules.scala 63:156:@7347.4]
  wire [11:0] _T_60495; // @[Modules.scala 63:156:@7349.4]
  wire [10:0] _T_60496; // @[Modules.scala 63:156:@7350.4]
  wire [10:0] buffer_1_741; // @[Modules.scala 63:156:@7351.4]
  wire [11:0] _T_60498; // @[Modules.scala 63:156:@7353.4]
  wire [10:0] _T_60499; // @[Modules.scala 63:156:@7354.4]
  wire [10:0] buffer_1_742; // @[Modules.scala 63:156:@7355.4]
  wire [11:0] _T_60501; // @[Modules.scala 63:156:@7357.4]
  wire [10:0] _T_60502; // @[Modules.scala 63:156:@7358.4]
  wire [10:0] buffer_1_743; // @[Modules.scala 63:156:@7359.4]
  wire [11:0] _T_60504; // @[Modules.scala 63:156:@7361.4]
  wire [10:0] _T_60505; // @[Modules.scala 63:156:@7362.4]
  wire [10:0] buffer_1_744; // @[Modules.scala 63:156:@7363.4]
  wire [11:0] _T_60507; // @[Modules.scala 63:156:@7365.4]
  wire [10:0] _T_60508; // @[Modules.scala 63:156:@7366.4]
  wire [10:0] buffer_1_745; // @[Modules.scala 63:156:@7367.4]
  wire [11:0] _T_60510; // @[Modules.scala 63:156:@7369.4]
  wire [10:0] _T_60511; // @[Modules.scala 63:156:@7370.4]
  wire [10:0] buffer_1_746; // @[Modules.scala 63:156:@7371.4]
  wire [11:0] _T_60513; // @[Modules.scala 63:156:@7373.4]
  wire [10:0] _T_60514; // @[Modules.scala 63:156:@7374.4]
  wire [10:0] buffer_1_747; // @[Modules.scala 63:156:@7375.4]
  wire [11:0] _T_60516; // @[Modules.scala 63:156:@7377.4]
  wire [10:0] _T_60517; // @[Modules.scala 63:156:@7378.4]
  wire [10:0] buffer_1_748; // @[Modules.scala 63:156:@7379.4]
  wire [11:0] _T_60519; // @[Modules.scala 63:156:@7381.4]
  wire [10:0] _T_60520; // @[Modules.scala 63:156:@7382.4]
  wire [10:0] buffer_1_749; // @[Modules.scala 63:156:@7383.4]
  wire [11:0] _T_60522; // @[Modules.scala 63:156:@7385.4]
  wire [10:0] _T_60523; // @[Modules.scala 63:156:@7386.4]
  wire [10:0] buffer_1_750; // @[Modules.scala 63:156:@7387.4]
  wire [11:0] _T_60525; // @[Modules.scala 63:156:@7389.4]
  wire [10:0] _T_60526; // @[Modules.scala 63:156:@7390.4]
  wire [10:0] buffer_1_751; // @[Modules.scala 63:156:@7391.4]
  wire [11:0] _T_60528; // @[Modules.scala 63:156:@7393.4]
  wire [10:0] _T_60529; // @[Modules.scala 63:156:@7394.4]
  wire [10:0] buffer_1_752; // @[Modules.scala 63:156:@7395.4]
  wire [11:0] _T_60531; // @[Modules.scala 63:156:@7397.4]
  wire [10:0] _T_60532; // @[Modules.scala 63:156:@7398.4]
  wire [10:0] buffer_1_753; // @[Modules.scala 63:156:@7399.4]
  wire [11:0] _T_60534; // @[Modules.scala 63:156:@7401.4]
  wire [10:0] _T_60535; // @[Modules.scala 63:156:@7402.4]
  wire [10:0] buffer_1_754; // @[Modules.scala 63:156:@7403.4]
  wire [11:0] _T_60537; // @[Modules.scala 63:156:@7405.4]
  wire [10:0] _T_60538; // @[Modules.scala 63:156:@7406.4]
  wire [10:0] buffer_1_755; // @[Modules.scala 63:156:@7407.4]
  wire [11:0] _T_60540; // @[Modules.scala 63:156:@7409.4]
  wire [10:0] _T_60541; // @[Modules.scala 63:156:@7410.4]
  wire [10:0] buffer_1_756; // @[Modules.scala 63:156:@7411.4]
  wire [11:0] _T_60543; // @[Modules.scala 63:156:@7413.4]
  wire [10:0] _T_60544; // @[Modules.scala 63:156:@7414.4]
  wire [10:0] buffer_1_757; // @[Modules.scala 63:156:@7415.4]
  wire [11:0] _T_60546; // @[Modules.scala 63:156:@7417.4]
  wire [10:0] _T_60547; // @[Modules.scala 63:156:@7418.4]
  wire [10:0] buffer_1_758; // @[Modules.scala 63:156:@7419.4]
  wire [11:0] _T_60549; // @[Modules.scala 63:156:@7421.4]
  wire [10:0] _T_60550; // @[Modules.scala 63:156:@7422.4]
  wire [10:0] buffer_1_759; // @[Modules.scala 63:156:@7423.4]
  wire [11:0] _T_60552; // @[Modules.scala 63:156:@7425.4]
  wire [10:0] _T_60553; // @[Modules.scala 63:156:@7426.4]
  wire [10:0] buffer_1_760; // @[Modules.scala 63:156:@7427.4]
  wire [11:0] _T_60555; // @[Modules.scala 63:156:@7429.4]
  wire [10:0] _T_60556; // @[Modules.scala 63:156:@7430.4]
  wire [10:0] buffer_1_761; // @[Modules.scala 63:156:@7431.4]
  wire [11:0] _T_60558; // @[Modules.scala 63:156:@7433.4]
  wire [10:0] _T_60559; // @[Modules.scala 63:156:@7434.4]
  wire [10:0] buffer_1_762; // @[Modules.scala 63:156:@7435.4]
  wire [11:0] _T_60561; // @[Modules.scala 63:156:@7437.4]
  wire [10:0] _T_60562; // @[Modules.scala 63:156:@7438.4]
  wire [10:0] buffer_1_763; // @[Modules.scala 63:156:@7439.4]
  wire [11:0] _T_60564; // @[Modules.scala 63:156:@7441.4]
  wire [10:0] _T_60565; // @[Modules.scala 63:156:@7442.4]
  wire [10:0] buffer_1_764; // @[Modules.scala 63:156:@7443.4]
  wire [11:0] _T_60567; // @[Modules.scala 63:156:@7445.4]
  wire [10:0] _T_60568; // @[Modules.scala 63:156:@7446.4]
  wire [10:0] buffer_1_765; // @[Modules.scala 63:156:@7447.4]
  wire [11:0] _T_60570; // @[Modules.scala 63:156:@7449.4]
  wire [10:0] _T_60571; // @[Modules.scala 63:156:@7450.4]
  wire [10:0] buffer_1_766; // @[Modules.scala 63:156:@7451.4]
  wire [11:0] _T_60573; // @[Modules.scala 63:156:@7453.4]
  wire [10:0] _T_60574; // @[Modules.scala 63:156:@7454.4]
  wire [10:0] buffer_1_767; // @[Modules.scala 63:156:@7455.4]
  wire [11:0] _T_60576; // @[Modules.scala 63:156:@7457.4]
  wire [10:0] _T_60577; // @[Modules.scala 63:156:@7458.4]
  wire [10:0] buffer_1_768; // @[Modules.scala 63:156:@7459.4]
  wire [11:0] _T_60579; // @[Modules.scala 63:156:@7461.4]
  wire [10:0] _T_60580; // @[Modules.scala 63:156:@7462.4]
  wire [10:0] buffer_1_769; // @[Modules.scala 63:156:@7463.4]
  wire [11:0] _T_60582; // @[Modules.scala 63:156:@7465.4]
  wire [10:0] _T_60583; // @[Modules.scala 63:156:@7466.4]
  wire [10:0] buffer_1_770; // @[Modules.scala 63:156:@7467.4]
  wire [11:0] _T_60585; // @[Modules.scala 63:156:@7469.4]
  wire [10:0] _T_60586; // @[Modules.scala 63:156:@7470.4]
  wire [10:0] buffer_1_771; // @[Modules.scala 63:156:@7471.4]
  wire [11:0] _T_60588; // @[Modules.scala 63:156:@7473.4]
  wire [10:0] _T_60589; // @[Modules.scala 63:156:@7474.4]
  wire [10:0] buffer_1_772; // @[Modules.scala 63:156:@7475.4]
  wire [11:0] _T_60591; // @[Modules.scala 63:156:@7477.4]
  wire [10:0] _T_60592; // @[Modules.scala 63:156:@7478.4]
  wire [10:0] buffer_1_773; // @[Modules.scala 63:156:@7479.4]
  wire [11:0] _T_60594; // @[Modules.scala 63:156:@7481.4]
  wire [10:0] _T_60595; // @[Modules.scala 63:156:@7482.4]
  wire [10:0] buffer_1_774; // @[Modules.scala 63:156:@7483.4]
  wire [11:0] _T_60597; // @[Modules.scala 63:156:@7485.4]
  wire [10:0] _T_60598; // @[Modules.scala 63:156:@7486.4]
  wire [10:0] buffer_1_775; // @[Modules.scala 63:156:@7487.4]
  wire [11:0] _T_60600; // @[Modules.scala 63:156:@7489.4]
  wire [10:0] _T_60601; // @[Modules.scala 63:156:@7490.4]
  wire [10:0] buffer_1_776; // @[Modules.scala 63:156:@7491.4]
  wire [11:0] _T_60603; // @[Modules.scala 63:156:@7493.4]
  wire [10:0] _T_60604; // @[Modules.scala 63:156:@7494.4]
  wire [10:0] buffer_1_777; // @[Modules.scala 63:156:@7495.4]
  wire [11:0] _T_60606; // @[Modules.scala 63:156:@7497.4]
  wire [10:0] _T_60607; // @[Modules.scala 63:156:@7498.4]
  wire [10:0] buffer_1_778; // @[Modules.scala 63:156:@7499.4]
  wire [11:0] _T_60609; // @[Modules.scala 63:156:@7501.4]
  wire [10:0] _T_60610; // @[Modules.scala 63:156:@7502.4]
  wire [10:0] buffer_1_779; // @[Modules.scala 63:156:@7503.4]
  wire [11:0] _T_60612; // @[Modules.scala 63:156:@7505.4]
  wire [10:0] _T_60613; // @[Modules.scala 63:156:@7506.4]
  wire [10:0] buffer_1_780; // @[Modules.scala 63:156:@7507.4]
  wire [11:0] _T_60615; // @[Modules.scala 63:156:@7509.4]
  wire [10:0] _T_60616; // @[Modules.scala 63:156:@7510.4]
  wire [10:0] buffer_1_781; // @[Modules.scala 63:156:@7511.4]
  wire [11:0] _T_60618; // @[Modules.scala 63:156:@7513.4]
  wire [10:0] _T_60619; // @[Modules.scala 63:156:@7514.4]
  wire [10:0] buffer_1_782; // @[Modules.scala 63:156:@7515.4]
  wire [11:0] _T_60621; // @[Modules.scala 63:156:@7517.4]
  wire [10:0] _T_60622; // @[Modules.scala 63:156:@7518.4]
  wire [10:0] buffer_1_783; // @[Modules.scala 63:156:@7519.4]
  wire [5:0] _T_60638; // @[Modules.scala 40:46:@7536.4]
  wire [4:0] _T_60639; // @[Modules.scala 40:46:@7537.4]
  wire [4:0] _T_60640; // @[Modules.scala 40:46:@7538.4]
  wire [5:0] _T_60645; // @[Modules.scala 46:47:@7543.4]
  wire [4:0] _T_60646; // @[Modules.scala 46:47:@7544.4]
  wire [4:0] _T_60647; // @[Modules.scala 46:47:@7545.4]
  wire [5:0] _T_60648; // @[Modules.scala 40:46:@7547.4]
  wire [4:0] _T_60649; // @[Modules.scala 40:46:@7548.4]
  wire [4:0] _T_60650; // @[Modules.scala 40:46:@7549.4]
  wire [5:0] _T_60651; // @[Modules.scala 37:46:@7551.4]
  wire [4:0] _T_60652; // @[Modules.scala 37:46:@7552.4]
  wire [4:0] _T_60653; // @[Modules.scala 37:46:@7553.4]
  wire [5:0] _T_60675; // @[Modules.scala 43:47:@7576.4]
  wire [4:0] _T_60676; // @[Modules.scala 43:47:@7577.4]
  wire [4:0] _T_60677; // @[Modules.scala 43:47:@7578.4]
  wire [5:0] _T_60678; // @[Modules.scala 40:46:@7580.4]
  wire [4:0] _T_60679; // @[Modules.scala 40:46:@7581.4]
  wire [4:0] _T_60680; // @[Modules.scala 40:46:@7582.4]
  wire [5:0] _T_60681; // @[Modules.scala 37:46:@7584.4]
  wire [4:0] _T_60682; // @[Modules.scala 37:46:@7585.4]
  wire [4:0] _T_60683; // @[Modules.scala 37:46:@7586.4]
  wire [5:0] _T_60688; // @[Modules.scala 46:47:@7591.4]
  wire [4:0] _T_60689; // @[Modules.scala 46:47:@7592.4]
  wire [4:0] _T_60690; // @[Modules.scala 46:47:@7593.4]
  wire [5:0] _T_60701; // @[Modules.scala 40:46:@7606.4]
  wire [4:0] _T_60702; // @[Modules.scala 40:46:@7607.4]
  wire [4:0] _T_60703; // @[Modules.scala 40:46:@7608.4]
  wire [5:0] _T_60705; // @[Modules.scala 46:37:@7610.4]
  wire [4:0] _T_60706; // @[Modules.scala 46:37:@7611.4]
  wire [4:0] _T_60707; // @[Modules.scala 46:37:@7612.4]
  wire [5:0] _T_60708; // @[Modules.scala 46:47:@7613.4]
  wire [4:0] _T_60709; // @[Modules.scala 46:47:@7614.4]
  wire [4:0] _T_60710; // @[Modules.scala 46:47:@7615.4]
  wire [5:0] _T_60720; // @[Modules.scala 40:46:@7629.4]
  wire [4:0] _T_60721; // @[Modules.scala 40:46:@7630.4]
  wire [4:0] _T_60722; // @[Modules.scala 40:46:@7631.4]
  wire [5:0] _T_60743; // @[Modules.scala 46:37:@7656.4]
  wire [4:0] _T_60744; // @[Modules.scala 46:37:@7657.4]
  wire [4:0] _T_60745; // @[Modules.scala 46:37:@7658.4]
  wire [5:0] _T_60746; // @[Modules.scala 46:47:@7659.4]
  wire [4:0] _T_60747; // @[Modules.scala 46:47:@7660.4]
  wire [4:0] _T_60748; // @[Modules.scala 46:47:@7661.4]
  wire [5:0] _T_60756; // @[Modules.scala 37:46:@7670.4]
  wire [4:0] _T_60757; // @[Modules.scala 37:46:@7671.4]
  wire [4:0] _T_60758; // @[Modules.scala 37:46:@7672.4]
  wire [5:0] _T_60763; // @[Modules.scala 43:47:@7677.4]
  wire [4:0] _T_60764; // @[Modules.scala 43:47:@7678.4]
  wire [4:0] _T_60765; // @[Modules.scala 43:47:@7679.4]
  wire [5:0] _T_60777; // @[Modules.scala 43:47:@7691.4]
  wire [4:0] _T_60778; // @[Modules.scala 43:47:@7692.4]
  wire [4:0] _T_60779; // @[Modules.scala 43:47:@7693.4]
  wire [5:0] _T_60793; // @[Modules.scala 43:47:@7710.4]
  wire [4:0] _T_60794; // @[Modules.scala 43:47:@7711.4]
  wire [4:0] _T_60795; // @[Modules.scala 43:47:@7712.4]
  wire [5:0] _T_60805; // @[Modules.scala 40:46:@7726.4]
  wire [4:0] _T_60806; // @[Modules.scala 40:46:@7727.4]
  wire [4:0] _T_60807; // @[Modules.scala 40:46:@7728.4]
  wire [5:0] _T_60815; // @[Modules.scala 37:46:@7737.4]
  wire [4:0] _T_60816; // @[Modules.scala 37:46:@7738.4]
  wire [4:0] _T_60817; // @[Modules.scala 37:46:@7739.4]
  wire [5:0] _T_60822; // @[Modules.scala 46:47:@7744.4]
  wire [4:0] _T_60823; // @[Modules.scala 46:47:@7745.4]
  wire [4:0] _T_60824; // @[Modules.scala 46:47:@7746.4]
  wire [5:0] _T_60832; // @[Modules.scala 40:46:@7755.4]
  wire [4:0] _T_60833; // @[Modules.scala 40:46:@7756.4]
  wire [4:0] _T_60834; // @[Modules.scala 40:46:@7757.4]
  wire [5:0] _T_60842; // @[Modules.scala 46:37:@7767.4]
  wire [4:0] _T_60843; // @[Modules.scala 46:37:@7768.4]
  wire [4:0] _T_60844; // @[Modules.scala 46:37:@7769.4]
  wire [5:0] _T_60845; // @[Modules.scala 46:47:@7770.4]
  wire [4:0] _T_60846; // @[Modules.scala 46:47:@7771.4]
  wire [4:0] _T_60847; // @[Modules.scala 46:47:@7772.4]
  wire [5:0] _T_60852; // @[Modules.scala 46:47:@7777.4]
  wire [4:0] _T_60853; // @[Modules.scala 46:47:@7778.4]
  wire [4:0] _T_60854; // @[Modules.scala 46:47:@7779.4]
  wire [5:0] _T_60856; // @[Modules.scala 46:37:@7781.4]
  wire [4:0] _T_60857; // @[Modules.scala 46:37:@7782.4]
  wire [4:0] _T_60858; // @[Modules.scala 46:37:@7783.4]
  wire [5:0] _T_60859; // @[Modules.scala 46:47:@7784.4]
  wire [4:0] _T_60860; // @[Modules.scala 46:47:@7785.4]
  wire [4:0] _T_60861; // @[Modules.scala 46:47:@7786.4]
  wire [5:0] _T_60862; // @[Modules.scala 40:46:@7788.4]
  wire [4:0] _T_60863; // @[Modules.scala 40:46:@7789.4]
  wire [4:0] _T_60864; // @[Modules.scala 40:46:@7790.4]
  wire [5:0] _T_60875; // @[Modules.scala 46:37:@7804.4]
  wire [4:0] _T_60876; // @[Modules.scala 46:37:@7805.4]
  wire [4:0] _T_60877; // @[Modules.scala 46:37:@7806.4]
  wire [5:0] _T_60878; // @[Modules.scala 46:47:@7807.4]
  wire [4:0] _T_60879; // @[Modules.scala 46:47:@7808.4]
  wire [4:0] _T_60880; // @[Modules.scala 46:47:@7809.4]
  wire [5:0] _T_60882; // @[Modules.scala 46:37:@7811.4]
  wire [4:0] _T_60883; // @[Modules.scala 46:37:@7812.4]
  wire [4:0] _T_60884; // @[Modules.scala 46:37:@7813.4]
  wire [5:0] _T_60885; // @[Modules.scala 46:47:@7814.4]
  wire [4:0] _T_60886; // @[Modules.scala 46:47:@7815.4]
  wire [4:0] _T_60887; // @[Modules.scala 46:47:@7816.4]
  wire [5:0] _T_60903; // @[Modules.scala 46:37:@7832.4]
  wire [4:0] _T_60904; // @[Modules.scala 46:37:@7833.4]
  wire [4:0] _T_60905; // @[Modules.scala 46:37:@7834.4]
  wire [5:0] _T_60906; // @[Modules.scala 46:47:@7835.4]
  wire [4:0] _T_60907; // @[Modules.scala 46:47:@7836.4]
  wire [4:0] _T_60908; // @[Modules.scala 46:47:@7837.4]
  wire [5:0] _T_60955; // @[Modules.scala 46:47:@7884.4]
  wire [4:0] _T_60956; // @[Modules.scala 46:47:@7885.4]
  wire [4:0] _T_60957; // @[Modules.scala 46:47:@7886.4]
  wire [5:0] _T_60979; // @[Modules.scala 43:37:@7910.4]
  wire [4:0] _T_60980; // @[Modules.scala 43:37:@7911.4]
  wire [4:0] _T_60981; // @[Modules.scala 43:37:@7912.4]
  wire [5:0] _T_60982; // @[Modules.scala 43:47:@7913.4]
  wire [4:0] _T_60983; // @[Modules.scala 43:47:@7914.4]
  wire [4:0] _T_60984; // @[Modules.scala 43:47:@7915.4]
  wire [5:0] _T_60985; // @[Modules.scala 40:46:@7917.4]
  wire [4:0] _T_60986; // @[Modules.scala 40:46:@7918.4]
  wire [4:0] _T_60987; // @[Modules.scala 40:46:@7919.4]
  wire [5:0] _T_61003; // @[Modules.scala 46:37:@7935.4]
  wire [4:0] _T_61004; // @[Modules.scala 46:37:@7936.4]
  wire [4:0] _T_61005; // @[Modules.scala 46:37:@7937.4]
  wire [5:0] _T_61006; // @[Modules.scala 46:47:@7938.4]
  wire [4:0] _T_61007; // @[Modules.scala 46:47:@7939.4]
  wire [4:0] _T_61008; // @[Modules.scala 46:47:@7940.4]
  wire [5:0] _T_61041; // @[Modules.scala 43:47:@7973.4]
  wire [4:0] _T_61042; // @[Modules.scala 43:47:@7974.4]
  wire [4:0] _T_61043; // @[Modules.scala 43:47:@7975.4]
  wire [5:0] _T_61044; // @[Modules.scala 37:46:@7977.4]
  wire [4:0] _T_61045; // @[Modules.scala 37:46:@7978.4]
  wire [4:0] _T_61046; // @[Modules.scala 37:46:@7979.4]
  wire [5:0] _T_61050; // @[Modules.scala 37:46:@7985.4]
  wire [4:0] _T_61051; // @[Modules.scala 37:46:@7986.4]
  wire [4:0] _T_61052; // @[Modules.scala 37:46:@7987.4]
  wire [5:0] _T_61056; // @[Modules.scala 40:46:@7993.4]
  wire [4:0] _T_61057; // @[Modules.scala 40:46:@7994.4]
  wire [4:0] _T_61058; // @[Modules.scala 40:46:@7995.4]
  wire [5:0] _T_61067; // @[Modules.scala 46:37:@8004.4]
  wire [4:0] _T_61068; // @[Modules.scala 46:37:@8005.4]
  wire [4:0] _T_61069; // @[Modules.scala 46:37:@8006.4]
  wire [5:0] _T_61070; // @[Modules.scala 46:47:@8007.4]
  wire [4:0] _T_61071; // @[Modules.scala 46:47:@8008.4]
  wire [4:0] _T_61072; // @[Modules.scala 46:47:@8009.4]
  wire [5:0] _T_61116; // @[Modules.scala 46:37:@8053.4]
  wire [4:0] _T_61117; // @[Modules.scala 46:37:@8054.4]
  wire [4:0] _T_61118; // @[Modules.scala 46:37:@8055.4]
  wire [5:0] _T_61119; // @[Modules.scala 46:47:@8056.4]
  wire [4:0] _T_61120; // @[Modules.scala 46:47:@8057.4]
  wire [4:0] _T_61121; // @[Modules.scala 46:47:@8058.4]
  wire [5:0] _T_61129; // @[Modules.scala 37:46:@8067.4]
  wire [4:0] _T_61130; // @[Modules.scala 37:46:@8068.4]
  wire [4:0] _T_61131; // @[Modules.scala 37:46:@8069.4]
  wire [5:0] _T_61132; // @[Modules.scala 37:46:@8071.4]
  wire [4:0] _T_61133; // @[Modules.scala 37:46:@8072.4]
  wire [4:0] _T_61134; // @[Modules.scala 37:46:@8073.4]
  wire [5:0] _T_61135; // @[Modules.scala 37:46:@8075.4]
  wire [4:0] _T_61136; // @[Modules.scala 37:46:@8076.4]
  wire [4:0] _T_61137; // @[Modules.scala 37:46:@8077.4]
  wire [5:0] _T_61145; // @[Modules.scala 46:47:@8086.4]
  wire [4:0] _T_61146; // @[Modules.scala 46:47:@8087.4]
  wire [4:0] _T_61147; // @[Modules.scala 46:47:@8088.4]
  wire [5:0] _T_61173; // @[Modules.scala 46:47:@8114.4]
  wire [4:0] _T_61174; // @[Modules.scala 46:47:@8115.4]
  wire [4:0] _T_61175; // @[Modules.scala 46:47:@8116.4]
  wire [5:0] _T_61180; // @[Modules.scala 46:47:@8121.4]
  wire [4:0] _T_61181; // @[Modules.scala 46:47:@8122.4]
  wire [4:0] _T_61182; // @[Modules.scala 46:47:@8123.4]
  wire [5:0] _T_61189; // @[Modules.scala 37:46:@8133.4]
  wire [4:0] _T_61190; // @[Modules.scala 37:46:@8134.4]
  wire [4:0] _T_61191; // @[Modules.scala 37:46:@8135.4]
  wire [5:0] _T_61199; // @[Modules.scala 37:46:@8144.4]
  wire [4:0] _T_61200; // @[Modules.scala 37:46:@8145.4]
  wire [4:0] _T_61201; // @[Modules.scala 37:46:@8146.4]
  wire [5:0] _T_61205; // @[Modules.scala 37:46:@8152.4]
  wire [4:0] _T_61206; // @[Modules.scala 37:46:@8153.4]
  wire [4:0] _T_61207; // @[Modules.scala 37:46:@8154.4]
  wire [5:0] _T_61247; // @[Modules.scala 43:47:@8194.4]
  wire [4:0] _T_61248; // @[Modules.scala 43:47:@8195.4]
  wire [4:0] _T_61249; // @[Modules.scala 43:47:@8196.4]
  wire [5:0] _T_61330; // @[Modules.scala 43:47:@8279.4]
  wire [4:0] _T_61331; // @[Modules.scala 43:47:@8280.4]
  wire [4:0] _T_61332; // @[Modules.scala 43:47:@8281.4]
  wire [5:0] _T_61337; // @[Modules.scala 43:47:@8286.4]
  wire [4:0] _T_61338; // @[Modules.scala 43:47:@8287.4]
  wire [4:0] _T_61339; // @[Modules.scala 43:47:@8288.4]
  wire [5:0] _T_61413; // @[Modules.scala 43:47:@8364.4]
  wire [4:0] _T_61414; // @[Modules.scala 43:47:@8365.4]
  wire [4:0] _T_61415; // @[Modules.scala 43:47:@8366.4]
  wire [5:0] _T_61416; // @[Modules.scala 37:46:@8368.4]
  wire [4:0] _T_61417; // @[Modules.scala 37:46:@8369.4]
  wire [4:0] _T_61418; // @[Modules.scala 37:46:@8370.4]
  wire [5:0] _T_61419; // @[Modules.scala 37:46:@8372.4]
  wire [4:0] _T_61420; // @[Modules.scala 37:46:@8373.4]
  wire [4:0] _T_61421; // @[Modules.scala 37:46:@8374.4]
  wire [5:0] _T_61468; // @[Modules.scala 43:47:@8421.4]
  wire [4:0] _T_61469; // @[Modules.scala 43:47:@8422.4]
  wire [4:0] _T_61470; // @[Modules.scala 43:47:@8423.4]
  wire [5:0] _T_61495; // @[Modules.scala 37:46:@8450.4]
  wire [4:0] _T_61496; // @[Modules.scala 37:46:@8451.4]
  wire [4:0] _T_61497; // @[Modules.scala 37:46:@8452.4]
  wire [5:0] _T_61504; // @[Modules.scala 40:46:@8462.4]
  wire [4:0] _T_61505; // @[Modules.scala 40:46:@8463.4]
  wire [4:0] _T_61506; // @[Modules.scala 40:46:@8464.4]
  wire [5:0] _T_61542; // @[Modules.scala 43:47:@8501.4]
  wire [4:0] _T_61543; // @[Modules.scala 43:47:@8502.4]
  wire [4:0] _T_61544; // @[Modules.scala 43:47:@8503.4]
  wire [5:0] _T_61587; // @[Modules.scala 40:46:@8554.4]
  wire [4:0] _T_61588; // @[Modules.scala 40:46:@8555.4]
  wire [4:0] _T_61589; // @[Modules.scala 40:46:@8556.4]
  wire [5:0] _T_61601; // @[Modules.scala 46:47:@8568.4]
  wire [4:0] _T_61602; // @[Modules.scala 46:47:@8569.4]
  wire [4:0] _T_61603; // @[Modules.scala 46:47:@8570.4]
  wire [5:0] _T_61608; // @[Modules.scala 43:47:@8575.4]
  wire [4:0] _T_61609; // @[Modules.scala 43:47:@8576.4]
  wire [4:0] _T_61610; // @[Modules.scala 43:47:@8577.4]
  wire [5:0] _T_61611; // @[Modules.scala 40:46:@8579.4]
  wire [4:0] _T_61612; // @[Modules.scala 40:46:@8580.4]
  wire [4:0] _T_61613; // @[Modules.scala 40:46:@8581.4]
  wire [5:0] _T_61656; // @[Modules.scala 37:46:@8632.4]
  wire [4:0] _T_61657; // @[Modules.scala 37:46:@8633.4]
  wire [4:0] _T_61658; // @[Modules.scala 37:46:@8634.4]
  wire [5:0] _T_61660; // @[Modules.scala 46:37:@8636.4]
  wire [4:0] _T_61661; // @[Modules.scala 46:37:@8637.4]
  wire [4:0] _T_61662; // @[Modules.scala 46:37:@8638.4]
  wire [5:0] _T_61663; // @[Modules.scala 46:47:@8639.4]
  wire [4:0] _T_61664; // @[Modules.scala 46:47:@8640.4]
  wire [4:0] _T_61665; // @[Modules.scala 46:47:@8641.4]
  wire [5:0] _T_61667; // @[Modules.scala 46:37:@8643.4]
  wire [4:0] _T_61668; // @[Modules.scala 46:37:@8644.4]
  wire [4:0] _T_61669; // @[Modules.scala 46:37:@8645.4]
  wire [5:0] _T_61670; // @[Modules.scala 46:47:@8646.4]
  wire [4:0] _T_61671; // @[Modules.scala 46:47:@8647.4]
  wire [4:0] _T_61672; // @[Modules.scala 46:47:@8648.4]
  wire [5:0] _T_61715; // @[Modules.scala 43:47:@8699.4]
  wire [4:0] _T_61716; // @[Modules.scala 43:47:@8700.4]
  wire [4:0] _T_61717; // @[Modules.scala 43:47:@8701.4]
  wire [5:0] _T_61725; // @[Modules.scala 46:37:@8711.4]
  wire [4:0] _T_61726; // @[Modules.scala 46:37:@8712.4]
  wire [4:0] _T_61727; // @[Modules.scala 46:37:@8713.4]
  wire [5:0] _T_61728; // @[Modules.scala 46:47:@8714.4]
  wire [4:0] _T_61729; // @[Modules.scala 46:47:@8715.4]
  wire [4:0] _T_61730; // @[Modules.scala 46:47:@8716.4]
  wire [5:0] _T_61745; // @[Modules.scala 37:46:@8732.4]
  wire [4:0] _T_61746; // @[Modules.scala 37:46:@8733.4]
  wire [4:0] _T_61747; // @[Modules.scala 37:46:@8734.4]
  wire [5:0] _T_61752; // @[Modules.scala 46:47:@8739.4]
  wire [4:0] _T_61753; // @[Modules.scala 46:47:@8740.4]
  wire [4:0] _T_61754; // @[Modules.scala 46:47:@8741.4]
  wire [5:0] _T_61762; // @[Modules.scala 46:37:@8751.4]
  wire [4:0] _T_61763; // @[Modules.scala 46:37:@8752.4]
  wire [4:0] _T_61764; // @[Modules.scala 46:37:@8753.4]
  wire [5:0] _T_61765; // @[Modules.scala 46:47:@8754.4]
  wire [4:0] _T_61766; // @[Modules.scala 46:47:@8755.4]
  wire [4:0] _T_61767; // @[Modules.scala 46:47:@8756.4]
  wire [5:0] _T_61785; // @[Modules.scala 46:47:@8776.4]
  wire [4:0] _T_61786; // @[Modules.scala 46:47:@8777.4]
  wire [4:0] _T_61787; // @[Modules.scala 46:47:@8778.4]
  wire [5:0] _T_61789; // @[Modules.scala 46:37:@8780.4]
  wire [4:0] _T_61790; // @[Modules.scala 46:37:@8781.4]
  wire [4:0] _T_61791; // @[Modules.scala 46:37:@8782.4]
  wire [5:0] _T_61792; // @[Modules.scala 46:47:@8783.4]
  wire [4:0] _T_61793; // @[Modules.scala 46:47:@8784.4]
  wire [4:0] _T_61794; // @[Modules.scala 46:47:@8785.4]
  wire [5:0] _T_61837; // @[Modules.scala 43:47:@8829.4]
  wire [4:0] _T_61838; // @[Modules.scala 43:47:@8830.4]
  wire [4:0] _T_61839; // @[Modules.scala 43:47:@8831.4]
  wire [5:0] _T_61840; // @[Modules.scala 40:46:@8833.4]
  wire [4:0] _T_61841; // @[Modules.scala 40:46:@8834.4]
  wire [4:0] _T_61842; // @[Modules.scala 40:46:@8835.4]
  wire [5:0] _T_61844; // @[Modules.scala 46:37:@8837.4]
  wire [4:0] _T_61845; // @[Modules.scala 46:37:@8838.4]
  wire [4:0] _T_61846; // @[Modules.scala 46:37:@8839.4]
  wire [5:0] _T_61847; // @[Modules.scala 46:47:@8840.4]
  wire [4:0] _T_61848; // @[Modules.scala 46:47:@8841.4]
  wire [4:0] _T_61849; // @[Modules.scala 46:47:@8842.4]
  wire [5:0] _T_61850; // @[Modules.scala 37:46:@8844.4]
  wire [4:0] _T_61851; // @[Modules.scala 37:46:@8845.4]
  wire [4:0] _T_61852; // @[Modules.scala 37:46:@8846.4]
  wire [5:0] _T_61860; // @[Modules.scala 43:47:@8855.4]
  wire [4:0] _T_61861; // @[Modules.scala 43:47:@8856.4]
  wire [4:0] _T_61862; // @[Modules.scala 43:47:@8857.4]
  wire [5:0] _T_61867; // @[Modules.scala 46:37:@8863.4]
  wire [4:0] _T_61868; // @[Modules.scala 46:37:@8864.4]
  wire [4:0] _T_61869; // @[Modules.scala 46:37:@8865.4]
  wire [5:0] _T_61870; // @[Modules.scala 46:47:@8866.4]
  wire [4:0] _T_61871; // @[Modules.scala 46:47:@8867.4]
  wire [4:0] _T_61872; // @[Modules.scala 46:47:@8868.4]
  wire [5:0] _T_61890; // @[Modules.scala 37:46:@8888.4]
  wire [4:0] _T_61891; // @[Modules.scala 37:46:@8889.4]
  wire [4:0] _T_61892; // @[Modules.scala 37:46:@8890.4]
  wire [5:0] _T_61904; // @[Modules.scala 46:37:@8903.4]
  wire [4:0] _T_61905; // @[Modules.scala 46:37:@8904.4]
  wire [4:0] _T_61906; // @[Modules.scala 46:37:@8905.4]
  wire [5:0] _T_61907; // @[Modules.scala 46:47:@8906.4]
  wire [4:0] _T_61908; // @[Modules.scala 46:47:@8907.4]
  wire [4:0] _T_61909; // @[Modules.scala 46:47:@8908.4]
  wire [5:0] _T_61914; // @[Modules.scala 43:47:@8913.4]
  wire [4:0] _T_61915; // @[Modules.scala 43:47:@8914.4]
  wire [4:0] _T_61916; // @[Modules.scala 43:47:@8915.4]
  wire [5:0] _T_61920; // @[Modules.scala 37:46:@8921.4]
  wire [4:0] _T_61921; // @[Modules.scala 37:46:@8922.4]
  wire [4:0] _T_61922; // @[Modules.scala 37:46:@8923.4]
  wire [5:0] _T_61940; // @[Modules.scala 46:37:@8944.4]
  wire [4:0] _T_61941; // @[Modules.scala 46:37:@8945.4]
  wire [4:0] _T_61942; // @[Modules.scala 46:37:@8946.4]
  wire [5:0] _T_61943; // @[Modules.scala 46:47:@8947.4]
  wire [4:0] _T_61944; // @[Modules.scala 46:47:@8948.4]
  wire [4:0] _T_61945; // @[Modules.scala 46:47:@8949.4]
  wire [5:0] _T_61971; // @[Modules.scala 46:47:@8975.4]
  wire [4:0] _T_61972; // @[Modules.scala 46:47:@8976.4]
  wire [4:0] _T_61973; // @[Modules.scala 46:47:@8977.4]
  wire [5:0] _T_61998; // @[Modules.scala 37:46:@9004.4]
  wire [4:0] _T_61999; // @[Modules.scala 37:46:@9005.4]
  wire [4:0] _T_62000; // @[Modules.scala 37:46:@9006.4]
  wire [5:0] _T_62001; // @[Modules.scala 40:46:@9008.4]
  wire [4:0] _T_62002; // @[Modules.scala 40:46:@9009.4]
  wire [4:0] _T_62003; // @[Modules.scala 40:46:@9010.4]
  wire [5:0] _T_62008; // @[Modules.scala 46:47:@9015.4]
  wire [4:0] _T_62009; // @[Modules.scala 46:47:@9016.4]
  wire [4:0] _T_62010; // @[Modules.scala 46:47:@9017.4]
  wire [5:0] _T_62022; // @[Modules.scala 46:47:@9029.4]
  wire [4:0] _T_62023; // @[Modules.scala 46:47:@9030.4]
  wire [4:0] _T_62024; // @[Modules.scala 46:47:@9031.4]
  wire [5:0] _T_62026; // @[Modules.scala 46:37:@9033.4]
  wire [4:0] _T_62027; // @[Modules.scala 46:37:@9034.4]
  wire [4:0] _T_62028; // @[Modules.scala 46:37:@9035.4]
  wire [5:0] _T_62029; // @[Modules.scala 46:47:@9036.4]
  wire [4:0] _T_62030; // @[Modules.scala 46:47:@9037.4]
  wire [4:0] _T_62031; // @[Modules.scala 46:47:@9038.4]
  wire [5:0] _T_62047; // @[Modules.scala 46:37:@9054.4]
  wire [4:0] _T_62048; // @[Modules.scala 46:37:@9055.4]
  wire [4:0] _T_62049; // @[Modules.scala 46:37:@9056.4]
  wire [5:0] _T_62050; // @[Modules.scala 46:47:@9057.4]
  wire [4:0] _T_62051; // @[Modules.scala 46:47:@9058.4]
  wire [4:0] _T_62052; // @[Modules.scala 46:47:@9059.4]
  wire [5:0] _T_62057; // @[Modules.scala 46:47:@9064.4]
  wire [4:0] _T_62058; // @[Modules.scala 46:47:@9065.4]
  wire [4:0] _T_62059; // @[Modules.scala 46:47:@9066.4]
  wire [5:0] _T_62092; // @[Modules.scala 43:47:@9099.4]
  wire [4:0] _T_62093; // @[Modules.scala 43:47:@9100.4]
  wire [4:0] _T_62094; // @[Modules.scala 43:47:@9101.4]
  wire [5:0] _T_62106; // @[Modules.scala 43:47:@9113.4]
  wire [4:0] _T_62107; // @[Modules.scala 43:47:@9114.4]
  wire [4:0] _T_62108; // @[Modules.scala 43:47:@9115.4]
  wire [5:0] _T_62110; // @[Modules.scala 43:37:@9117.4]
  wire [4:0] _T_62111; // @[Modules.scala 43:37:@9118.4]
  wire [4:0] _T_62112; // @[Modules.scala 43:37:@9119.4]
  wire [5:0] _T_62113; // @[Modules.scala 43:47:@9120.4]
  wire [4:0] _T_62114; // @[Modules.scala 43:47:@9121.4]
  wire [4:0] _T_62115; // @[Modules.scala 43:47:@9122.4]
  wire [5:0] _T_62116; // @[Modules.scala 37:46:@9124.4]
  wire [4:0] _T_62117; // @[Modules.scala 37:46:@9125.4]
  wire [4:0] _T_62118; // @[Modules.scala 37:46:@9126.4]
  wire [5:0] _T_62140; // @[Modules.scala 40:46:@9149.4]
  wire [4:0] _T_62141; // @[Modules.scala 40:46:@9150.4]
  wire [4:0] _T_62142; // @[Modules.scala 40:46:@9151.4]
  wire [5:0] _T_62182; // @[Modules.scala 46:47:@9191.4]
  wire [4:0] _T_62183; // @[Modules.scala 46:47:@9192.4]
  wire [4:0] _T_62184; // @[Modules.scala 46:47:@9193.4]
  wire [5:0] _T_62195; // @[Modules.scala 46:37:@9207.4]
  wire [4:0] _T_62196; // @[Modules.scala 46:37:@9208.4]
  wire [4:0] _T_62197; // @[Modules.scala 46:37:@9209.4]
  wire [5:0] _T_62198; // @[Modules.scala 46:47:@9210.4]
  wire [4:0] _T_62199; // @[Modules.scala 46:47:@9211.4]
  wire [4:0] _T_62200; // @[Modules.scala 46:47:@9212.4]
  wire [5:0] _T_62222; // @[Modules.scala 40:46:@9235.4]
  wire [4:0] _T_62223; // @[Modules.scala 40:46:@9236.4]
  wire [4:0] _T_62224; // @[Modules.scala 40:46:@9237.4]
  wire [5:0] _T_62225; // @[Modules.scala 40:46:@9239.4]
  wire [4:0] _T_62226; // @[Modules.scala 40:46:@9240.4]
  wire [4:0] _T_62227; // @[Modules.scala 40:46:@9241.4]
  wire [5:0] _T_62239; // @[Modules.scala 43:47:@9253.4]
  wire [4:0] _T_62240; // @[Modules.scala 43:47:@9254.4]
  wire [4:0] _T_62241; // @[Modules.scala 43:47:@9255.4]
  wire [5:0] _T_62242; // @[Modules.scala 37:46:@9257.4]
  wire [4:0] _T_62243; // @[Modules.scala 37:46:@9258.4]
  wire [4:0] _T_62244; // @[Modules.scala 37:46:@9259.4]
  wire [5:0] _T_62245; // @[Modules.scala 40:46:@9261.4]
  wire [4:0] _T_62246; // @[Modules.scala 40:46:@9262.4]
  wire [4:0] _T_62247; // @[Modules.scala 40:46:@9263.4]
  wire [5:0] _T_62249; // @[Modules.scala 43:37:@9265.4]
  wire [4:0] _T_62250; // @[Modules.scala 43:37:@9266.4]
  wire [4:0] _T_62251; // @[Modules.scala 43:37:@9267.4]
  wire [5:0] _T_62252; // @[Modules.scala 43:47:@9268.4]
  wire [4:0] _T_62253; // @[Modules.scala 43:47:@9269.4]
  wire [4:0] _T_62254; // @[Modules.scala 43:47:@9270.4]
  wire [5:0] _T_62259; // @[Modules.scala 43:37:@9276.4]
  wire [4:0] _T_62260; // @[Modules.scala 43:37:@9277.4]
  wire [4:0] _T_62261; // @[Modules.scala 43:37:@9278.4]
  wire [5:0] _T_62262; // @[Modules.scala 43:47:@9279.4]
  wire [4:0] _T_62263; // @[Modules.scala 43:47:@9280.4]
  wire [4:0] _T_62264; // @[Modules.scala 43:47:@9281.4]
  wire [5:0] _T_62266; // @[Modules.scala 46:37:@9283.4]
  wire [4:0] _T_62267; // @[Modules.scala 46:37:@9284.4]
  wire [4:0] _T_62268; // @[Modules.scala 46:37:@9285.4]
  wire [5:0] _T_62269; // @[Modules.scala 46:47:@9286.4]
  wire [4:0] _T_62270; // @[Modules.scala 46:47:@9287.4]
  wire [4:0] _T_62271; // @[Modules.scala 46:47:@9288.4]
  wire [5:0] _T_62272; // @[Modules.scala 37:46:@9290.4]
  wire [4:0] _T_62273; // @[Modules.scala 37:46:@9291.4]
  wire [4:0] _T_62274; // @[Modules.scala 37:46:@9292.4]
  wire [5:0] _T_62275; // @[Modules.scala 40:46:@9294.4]
  wire [4:0] _T_62276; // @[Modules.scala 40:46:@9295.4]
  wire [4:0] _T_62277; // @[Modules.scala 40:46:@9296.4]
  wire [5:0] _T_62292; // @[Modules.scala 37:46:@9312.4]
  wire [4:0] _T_62293; // @[Modules.scala 37:46:@9313.4]
  wire [4:0] _T_62294; // @[Modules.scala 37:46:@9314.4]
  wire [5:0] _T_62296; // @[Modules.scala 46:37:@9316.4]
  wire [4:0] _T_62297; // @[Modules.scala 46:37:@9317.4]
  wire [4:0] _T_62298; // @[Modules.scala 46:37:@9318.4]
  wire [5:0] _T_62299; // @[Modules.scala 46:47:@9319.4]
  wire [4:0] _T_62300; // @[Modules.scala 46:47:@9320.4]
  wire [4:0] _T_62301; // @[Modules.scala 46:47:@9321.4]
  wire [5:0] _T_62316; // @[Modules.scala 40:46:@9337.4]
  wire [4:0] _T_62317; // @[Modules.scala 40:46:@9338.4]
  wire [4:0] _T_62318; // @[Modules.scala 40:46:@9339.4]
  wire [5:0] _T_62343; // @[Modules.scala 37:46:@9366.4]
  wire [4:0] _T_62344; // @[Modules.scala 37:46:@9367.4]
  wire [4:0] _T_62345; // @[Modules.scala 37:46:@9368.4]
  wire [5:0] _T_62362; // @[Modules.scala 40:46:@9389.4]
  wire [4:0] _T_62363; // @[Modules.scala 40:46:@9390.4]
  wire [4:0] _T_62364; // @[Modules.scala 40:46:@9391.4]
  wire [5:0] _T_62365; // @[Modules.scala 40:46:@9393.4]
  wire [4:0] _T_62366; // @[Modules.scala 40:46:@9394.4]
  wire [4:0] _T_62367; // @[Modules.scala 40:46:@9395.4]
  wire [5:0] _T_62372; // @[Modules.scala 43:47:@9400.4]
  wire [4:0] _T_62373; // @[Modules.scala 43:47:@9401.4]
  wire [4:0] _T_62374; // @[Modules.scala 43:47:@9402.4]
  wire [5:0] _T_62375; // @[Modules.scala 40:46:@9404.4]
  wire [4:0] _T_62376; // @[Modules.scala 40:46:@9405.4]
  wire [4:0] _T_62377; // @[Modules.scala 40:46:@9406.4]
  wire [5:0] _T_62388; // @[Modules.scala 40:46:@9419.4]
  wire [4:0] _T_62389; // @[Modules.scala 40:46:@9420.4]
  wire [4:0] _T_62390; // @[Modules.scala 40:46:@9421.4]
  wire [5:0] _T_62394; // @[Modules.scala 37:46:@9427.4]
  wire [4:0] _T_62395; // @[Modules.scala 37:46:@9428.4]
  wire [4:0] _T_62396; // @[Modules.scala 37:46:@9429.4]
  wire [5:0] _T_62413; // @[Modules.scala 37:46:@9450.4]
  wire [4:0] _T_62414; // @[Modules.scala 37:46:@9451.4]
  wire [4:0] _T_62415; // @[Modules.scala 37:46:@9452.4]
  wire [5:0] _T_62427; // @[Modules.scala 46:37:@9465.4]
  wire [4:0] _T_62428; // @[Modules.scala 46:37:@9466.4]
  wire [4:0] _T_62429; // @[Modules.scala 46:37:@9467.4]
  wire [5:0] _T_62430; // @[Modules.scala 46:47:@9468.4]
  wire [4:0] _T_62431; // @[Modules.scala 46:47:@9469.4]
  wire [4:0] _T_62432; // @[Modules.scala 46:47:@9470.4]
  wire [5:0] _T_62434; // @[Modules.scala 46:37:@9472.4]
  wire [4:0] _T_62435; // @[Modules.scala 46:37:@9473.4]
  wire [4:0] _T_62436; // @[Modules.scala 46:37:@9474.4]
  wire [5:0] _T_62437; // @[Modules.scala 46:47:@9475.4]
  wire [4:0] _T_62438; // @[Modules.scala 46:47:@9476.4]
  wire [4:0] _T_62439; // @[Modules.scala 46:47:@9477.4]
  wire [5:0] _T_62444; // @[Modules.scala 46:47:@9482.4]
  wire [4:0] _T_62445; // @[Modules.scala 46:47:@9483.4]
  wire [4:0] _T_62446; // @[Modules.scala 46:47:@9484.4]
  wire [5:0] _T_62448; // @[Modules.scala 46:37:@9486.4]
  wire [4:0] _T_62449; // @[Modules.scala 46:37:@9487.4]
  wire [4:0] _T_62450; // @[Modules.scala 46:37:@9488.4]
  wire [5:0] _T_62451; // @[Modules.scala 46:47:@9489.4]
  wire [4:0] _T_62452; // @[Modules.scala 46:47:@9490.4]
  wire [4:0] _T_62453; // @[Modules.scala 46:47:@9491.4]
  wire [5:0] _T_62454; // @[Modules.scala 40:46:@9493.4]
  wire [4:0] _T_62455; // @[Modules.scala 40:46:@9494.4]
  wire [4:0] _T_62456; // @[Modules.scala 40:46:@9495.4]
  wire [5:0] _T_62465; // @[Modules.scala 43:37:@9504.4]
  wire [4:0] _T_62466; // @[Modules.scala 43:37:@9505.4]
  wire [4:0] _T_62467; // @[Modules.scala 43:37:@9506.4]
  wire [5:0] _T_62468; // @[Modules.scala 43:47:@9507.4]
  wire [4:0] _T_62469; // @[Modules.scala 43:47:@9508.4]
  wire [4:0] _T_62470; // @[Modules.scala 43:47:@9509.4]
  wire [5:0] _T_62481; // @[Modules.scala 46:37:@9523.4]
  wire [4:0] _T_62482; // @[Modules.scala 46:37:@9524.4]
  wire [4:0] _T_62483; // @[Modules.scala 46:37:@9525.4]
  wire [5:0] _T_62484; // @[Modules.scala 46:47:@9526.4]
  wire [4:0] _T_62485; // @[Modules.scala 46:47:@9527.4]
  wire [4:0] _T_62486; // @[Modules.scala 46:47:@9528.4]
  wire [5:0] _T_62498; // @[Modules.scala 46:47:@9540.4]
  wire [4:0] _T_62499; // @[Modules.scala 46:47:@9541.4]
  wire [4:0] _T_62500; // @[Modules.scala 46:47:@9542.4]
  wire [5:0] _T_62505; // @[Modules.scala 46:37:@9548.4]
  wire [4:0] _T_62506; // @[Modules.scala 46:37:@9549.4]
  wire [4:0] _T_62507; // @[Modules.scala 46:37:@9550.4]
  wire [5:0] _T_62508; // @[Modules.scala 46:47:@9551.4]
  wire [4:0] _T_62509; // @[Modules.scala 46:47:@9552.4]
  wire [4:0] _T_62510; // @[Modules.scala 46:47:@9553.4]
  wire [5:0] _T_62512; // @[Modules.scala 46:37:@9555.4]
  wire [4:0] _T_62513; // @[Modules.scala 46:37:@9556.4]
  wire [4:0] _T_62514; // @[Modules.scala 46:37:@9557.4]
  wire [5:0] _T_62515; // @[Modules.scala 46:47:@9558.4]
  wire [4:0] _T_62516; // @[Modules.scala 46:47:@9559.4]
  wire [4:0] _T_62517; // @[Modules.scala 46:47:@9560.4]
  wire [5:0] _T_62529; // @[Modules.scala 46:47:@9572.4]
  wire [4:0] _T_62530; // @[Modules.scala 46:47:@9573.4]
  wire [4:0] _T_62531; // @[Modules.scala 46:47:@9574.4]
  wire [5:0] _T_62543; // @[Modules.scala 46:47:@9586.4]
  wire [4:0] _T_62544; // @[Modules.scala 46:47:@9587.4]
  wire [4:0] _T_62545; // @[Modules.scala 46:47:@9588.4]
  wire [5:0] _T_62547; // @[Modules.scala 46:37:@9590.4]
  wire [4:0] _T_62548; // @[Modules.scala 46:37:@9591.4]
  wire [4:0] _T_62549; // @[Modules.scala 46:37:@9592.4]
  wire [5:0] _T_62550; // @[Modules.scala 46:47:@9593.4]
  wire [4:0] _T_62551; // @[Modules.scala 46:47:@9594.4]
  wire [4:0] _T_62552; // @[Modules.scala 46:47:@9595.4]
  wire [5:0] _T_62576; // @[Modules.scala 37:46:@9623.4]
  wire [4:0] _T_62577; // @[Modules.scala 37:46:@9624.4]
  wire [4:0] _T_62578; // @[Modules.scala 37:46:@9625.4]
  wire [5:0] _T_62579; // @[Modules.scala 37:46:@9627.4]
  wire [4:0] _T_62580; // @[Modules.scala 37:46:@9628.4]
  wire [4:0] _T_62581; // @[Modules.scala 37:46:@9629.4]
  wire [5:0] _T_62582; // @[Modules.scala 40:46:@9631.4]
  wire [4:0] _T_62583; // @[Modules.scala 40:46:@9632.4]
  wire [4:0] _T_62584; // @[Modules.scala 40:46:@9633.4]
  wire [5:0] _T_62634; // @[Modules.scala 40:46:@9684.4]
  wire [4:0] _T_62635; // @[Modules.scala 40:46:@9685.4]
  wire [4:0] _T_62636; // @[Modules.scala 40:46:@9686.4]
  wire [5:0] _T_62638; // @[Modules.scala 43:37:@9688.4]
  wire [4:0] _T_62639; // @[Modules.scala 43:37:@9689.4]
  wire [4:0] _T_62640; // @[Modules.scala 43:37:@9690.4]
  wire [5:0] _T_62641; // @[Modules.scala 43:47:@9691.4]
  wire [4:0] _T_62642; // @[Modules.scala 43:47:@9692.4]
  wire [4:0] _T_62643; // @[Modules.scala 43:47:@9693.4]
  wire [5:0] _T_62647; // @[Modules.scala 40:46:@9699.4]
  wire [4:0] _T_62648; // @[Modules.scala 40:46:@9700.4]
  wire [4:0] _T_62649; // @[Modules.scala 40:46:@9701.4]
  wire [5:0] _T_62654; // @[Modules.scala 46:47:@9706.4]
  wire [4:0] _T_62655; // @[Modules.scala 46:47:@9707.4]
  wire [4:0] _T_62656; // @[Modules.scala 46:47:@9708.4]
  wire [5:0] _T_62733; // @[Modules.scala 43:47:@9788.4]
  wire [4:0] _T_62734; // @[Modules.scala 43:47:@9789.4]
  wire [4:0] _T_62735; // @[Modules.scala 43:47:@9790.4]
  wire [10:0] buffer_2_2; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_3; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62739; // @[Modules.scala 50:57:@9796.4]
  wire [10:0] _T_62740; // @[Modules.scala 50:57:@9797.4]
  wire [10:0] buffer_2_393; // @[Modules.scala 50:57:@9798.4]
  wire [10:0] buffer_2_4; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62742; // @[Modules.scala 50:57:@9800.4]
  wire [10:0] _T_62743; // @[Modules.scala 50:57:@9801.4]
  wire [10:0] buffer_2_394; // @[Modules.scala 50:57:@9802.4]
  wire [10:0] buffer_2_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62748; // @[Modules.scala 50:57:@9808.4]
  wire [10:0] _T_62749; // @[Modules.scala 50:57:@9809.4]
  wire [10:0] buffer_2_396; // @[Modules.scala 50:57:@9810.4]
  wire [10:0] buffer_2_10; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62751; // @[Modules.scala 50:57:@9812.4]
  wire [10:0] _T_62752; // @[Modules.scala 50:57:@9813.4]
  wire [10:0] buffer_2_397; // @[Modules.scala 50:57:@9814.4]
  wire [10:0] buffer_2_12; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62754; // @[Modules.scala 50:57:@9816.4]
  wire [10:0] _T_62755; // @[Modules.scala 50:57:@9817.4]
  wire [10:0] buffer_2_398; // @[Modules.scala 50:57:@9818.4]
  wire [10:0] buffer_2_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62757; // @[Modules.scala 50:57:@9820.4]
  wire [10:0] _T_62758; // @[Modules.scala 50:57:@9821.4]
  wire [10:0] buffer_2_399; // @[Modules.scala 50:57:@9822.4]
  wire [10:0] buffer_2_16; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62760; // @[Modules.scala 50:57:@9824.4]
  wire [10:0] _T_62761; // @[Modules.scala 50:57:@9825.4]
  wire [10:0] buffer_2_400; // @[Modules.scala 50:57:@9826.4]
  wire [10:0] buffer_2_20; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62766; // @[Modules.scala 50:57:@9832.4]
  wire [10:0] _T_62767; // @[Modules.scala 50:57:@9833.4]
  wire [10:0] buffer_2_402; // @[Modules.scala 50:57:@9834.4]
  wire [11:0] _T_62769; // @[Modules.scala 50:57:@9836.4]
  wire [10:0] _T_62770; // @[Modules.scala 50:57:@9837.4]
  wire [10:0] buffer_2_403; // @[Modules.scala 50:57:@9838.4]
  wire [10:0] buffer_2_26; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62775; // @[Modules.scala 50:57:@9844.4]
  wire [10:0] _T_62776; // @[Modules.scala 50:57:@9845.4]
  wire [10:0] buffer_2_405; // @[Modules.scala 50:57:@9846.4]
  wire [10:0] buffer_2_28; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62778; // @[Modules.scala 50:57:@9848.4]
  wire [10:0] _T_62779; // @[Modules.scala 50:57:@9849.4]
  wire [10:0] buffer_2_406; // @[Modules.scala 50:57:@9850.4]
  wire [10:0] buffer_2_31; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62781; // @[Modules.scala 50:57:@9852.4]
  wire [10:0] _T_62782; // @[Modules.scala 50:57:@9853.4]
  wire [10:0] buffer_2_407; // @[Modules.scala 50:57:@9854.4]
  wire [10:0] buffer_2_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62787; // @[Modules.scala 50:57:@9860.4]
  wire [10:0] _T_62788; // @[Modules.scala 50:57:@9861.4]
  wire [10:0] buffer_2_409; // @[Modules.scala 50:57:@9862.4]
  wire [10:0] buffer_2_39; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62793; // @[Modules.scala 50:57:@9868.4]
  wire [10:0] _T_62794; // @[Modules.scala 50:57:@9869.4]
  wire [10:0] buffer_2_411; // @[Modules.scala 50:57:@9870.4]
  wire [10:0] buffer_2_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62796; // @[Modules.scala 50:57:@9872.4]
  wire [10:0] _T_62797; // @[Modules.scala 50:57:@9873.4]
  wire [10:0] buffer_2_412; // @[Modules.scala 50:57:@9874.4]
  wire [10:0] buffer_2_42; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62799; // @[Modules.scala 50:57:@9876.4]
  wire [10:0] _T_62800; // @[Modules.scala 50:57:@9877.4]
  wire [10:0] buffer_2_413; // @[Modules.scala 50:57:@9878.4]
  wire [10:0] buffer_2_44; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62802; // @[Modules.scala 50:57:@9880.4]
  wire [10:0] _T_62803; // @[Modules.scala 50:57:@9881.4]
  wire [10:0] buffer_2_414; // @[Modules.scala 50:57:@9882.4]
  wire [10:0] buffer_2_47; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62805; // @[Modules.scala 50:57:@9884.4]
  wire [10:0] _T_62806; // @[Modules.scala 50:57:@9885.4]
  wire [10:0] buffer_2_415; // @[Modules.scala 50:57:@9886.4]
  wire [10:0] buffer_2_48; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_49; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62808; // @[Modules.scala 50:57:@9888.4]
  wire [10:0] _T_62809; // @[Modules.scala 50:57:@9889.4]
  wire [10:0] buffer_2_416; // @[Modules.scala 50:57:@9890.4]
  wire [10:0] buffer_2_50; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62811; // @[Modules.scala 50:57:@9892.4]
  wire [10:0] _T_62812; // @[Modules.scala 50:57:@9893.4]
  wire [10:0] buffer_2_417; // @[Modules.scala 50:57:@9894.4]
  wire [10:0] buffer_2_54; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62817; // @[Modules.scala 50:57:@9900.4]
  wire [10:0] _T_62818; // @[Modules.scala 50:57:@9901.4]
  wire [10:0] buffer_2_419; // @[Modules.scala 50:57:@9902.4]
  wire [10:0] buffer_2_58; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62823; // @[Modules.scala 50:57:@9908.4]
  wire [10:0] _T_62824; // @[Modules.scala 50:57:@9909.4]
  wire [10:0] buffer_2_421; // @[Modules.scala 50:57:@9910.4]
  wire [10:0] buffer_2_65; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62832; // @[Modules.scala 50:57:@9920.4]
  wire [10:0] _T_62833; // @[Modules.scala 50:57:@9921.4]
  wire [10:0] buffer_2_424; // @[Modules.scala 50:57:@9922.4]
  wire [10:0] buffer_2_70; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62841; // @[Modules.scala 50:57:@9932.4]
  wire [10:0] _T_62842; // @[Modules.scala 50:57:@9933.4]
  wire [10:0] buffer_2_427; // @[Modules.scala 50:57:@9934.4]
  wire [10:0] buffer_2_74; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62847; // @[Modules.scala 50:57:@9940.4]
  wire [10:0] _T_62848; // @[Modules.scala 50:57:@9941.4]
  wire [10:0] buffer_2_429; // @[Modules.scala 50:57:@9942.4]
  wire [10:0] buffer_2_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62853; // @[Modules.scala 50:57:@9948.4]
  wire [10:0] _T_62854; // @[Modules.scala 50:57:@9949.4]
  wire [10:0] buffer_2_431; // @[Modules.scala 50:57:@9950.4]
  wire [10:0] buffer_2_80; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62856; // @[Modules.scala 50:57:@9952.4]
  wire [10:0] _T_62857; // @[Modules.scala 50:57:@9953.4]
  wire [10:0] buffer_2_432; // @[Modules.scala 50:57:@9954.4]
  wire [10:0] buffer_2_82; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62859; // @[Modules.scala 50:57:@9956.4]
  wire [10:0] _T_62860; // @[Modules.scala 50:57:@9957.4]
  wire [10:0] buffer_2_433; // @[Modules.scala 50:57:@9958.4]
  wire [10:0] buffer_2_84; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62862; // @[Modules.scala 50:57:@9960.4]
  wire [10:0] _T_62863; // @[Modules.scala 50:57:@9961.4]
  wire [10:0] buffer_2_434; // @[Modules.scala 50:57:@9962.4]
  wire [10:0] buffer_2_86; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62865; // @[Modules.scala 50:57:@9964.4]
  wire [10:0] _T_62866; // @[Modules.scala 50:57:@9965.4]
  wire [10:0] buffer_2_435; // @[Modules.scala 50:57:@9966.4]
  wire [10:0] buffer_2_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62874; // @[Modules.scala 50:57:@9976.4]
  wire [10:0] _T_62875; // @[Modules.scala 50:57:@9977.4]
  wire [10:0] buffer_2_438; // @[Modules.scala 50:57:@9978.4]
  wire [10:0] buffer_2_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62877; // @[Modules.scala 50:57:@9980.4]
  wire [10:0] _T_62878; // @[Modules.scala 50:57:@9981.4]
  wire [10:0] buffer_2_439; // @[Modules.scala 50:57:@9982.4]
  wire [10:0] buffer_2_96; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62880; // @[Modules.scala 50:57:@9984.4]
  wire [10:0] _T_62881; // @[Modules.scala 50:57:@9985.4]
  wire [10:0] buffer_2_440; // @[Modules.scala 50:57:@9986.4]
  wire [10:0] buffer_2_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62883; // @[Modules.scala 50:57:@9988.4]
  wire [10:0] _T_62884; // @[Modules.scala 50:57:@9989.4]
  wire [10:0] buffer_2_441; // @[Modules.scala 50:57:@9990.4]
  wire [10:0] buffer_2_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62889; // @[Modules.scala 50:57:@9996.4]
  wire [10:0] _T_62890; // @[Modules.scala 50:57:@9997.4]
  wire [10:0] buffer_2_443; // @[Modules.scala 50:57:@9998.4]
  wire [10:0] buffer_2_104; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62892; // @[Modules.scala 50:57:@10000.4]
  wire [10:0] _T_62893; // @[Modules.scala 50:57:@10001.4]
  wire [10:0] buffer_2_444; // @[Modules.scala 50:57:@10002.4]
  wire [10:0] buffer_2_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62895; // @[Modules.scala 50:57:@10004.4]
  wire [10:0] _T_62896; // @[Modules.scala 50:57:@10005.4]
  wire [10:0] buffer_2_445; // @[Modules.scala 50:57:@10006.4]
  wire [10:0] buffer_2_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62898; // @[Modules.scala 50:57:@10008.4]
  wire [10:0] _T_62899; // @[Modules.scala 50:57:@10009.4]
  wire [10:0] buffer_2_446; // @[Modules.scala 50:57:@10010.4]
  wire [10:0] buffer_2_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62901; // @[Modules.scala 50:57:@10012.4]
  wire [10:0] _T_62902; // @[Modules.scala 50:57:@10013.4]
  wire [10:0] buffer_2_447; // @[Modules.scala 50:57:@10014.4]
  wire [10:0] buffer_2_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62910; // @[Modules.scala 50:57:@10024.4]
  wire [10:0] _T_62911; // @[Modules.scala 50:57:@10025.4]
  wire [10:0] buffer_2_450; // @[Modules.scala 50:57:@10026.4]
  wire [10:0] buffer_2_130; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62931; // @[Modules.scala 50:57:@10052.4]
  wire [10:0] _T_62932; // @[Modules.scala 50:57:@10053.4]
  wire [10:0] buffer_2_457; // @[Modules.scala 50:57:@10054.4]
  wire [10:0] buffer_2_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62949; // @[Modules.scala 50:57:@10076.4]
  wire [10:0] _T_62950; // @[Modules.scala 50:57:@10077.4]
  wire [10:0] buffer_2_463; // @[Modules.scala 50:57:@10078.4]
  wire [10:0] buffer_2_144; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62952; // @[Modules.scala 50:57:@10080.4]
  wire [10:0] _T_62953; // @[Modules.scala 50:57:@10081.4]
  wire [10:0] buffer_2_464; // @[Modules.scala 50:57:@10082.4]
  wire [10:0] buffer_2_152; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62964; // @[Modules.scala 50:57:@10096.4]
  wire [10:0] _T_62965; // @[Modules.scala 50:57:@10097.4]
  wire [10:0] buffer_2_468; // @[Modules.scala 50:57:@10098.4]
  wire [10:0] buffer_2_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62970; // @[Modules.scala 50:57:@10104.4]
  wire [10:0] _T_62971; // @[Modules.scala 50:57:@10105.4]
  wire [10:0] buffer_2_470; // @[Modules.scala 50:57:@10106.4]
  wire [10:0] buffer_2_160; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62976; // @[Modules.scala 50:57:@10112.4]
  wire [10:0] _T_62977; // @[Modules.scala 50:57:@10113.4]
  wire [10:0] buffer_2_472; // @[Modules.scala 50:57:@10114.4]
  wire [11:0] _T_62982; // @[Modules.scala 50:57:@10120.4]
  wire [10:0] _T_62983; // @[Modules.scala 50:57:@10121.4]
  wire [10:0] buffer_2_474; // @[Modules.scala 50:57:@10122.4]
  wire [10:0] buffer_2_166; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62985; // @[Modules.scala 50:57:@10124.4]
  wire [10:0] _T_62986; // @[Modules.scala 50:57:@10125.4]
  wire [10:0] buffer_2_475; // @[Modules.scala 50:57:@10126.4]
  wire [10:0] buffer_2_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63000; // @[Modules.scala 50:57:@10144.4]
  wire [10:0] _T_63001; // @[Modules.scala 50:57:@10145.4]
  wire [10:0] buffer_2_480; // @[Modules.scala 50:57:@10146.4]
  wire [10:0] buffer_2_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63003; // @[Modules.scala 50:57:@10148.4]
  wire [10:0] _T_63004; // @[Modules.scala 50:57:@10149.4]
  wire [10:0] buffer_2_481; // @[Modules.scala 50:57:@10150.4]
  wire [10:0] buffer_2_180; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63006; // @[Modules.scala 50:57:@10152.4]
  wire [10:0] _T_63007; // @[Modules.scala 50:57:@10153.4]
  wire [10:0] buffer_2_482; // @[Modules.scala 50:57:@10154.4]
  wire [10:0] buffer_2_192; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_193; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63024; // @[Modules.scala 50:57:@10176.4]
  wire [10:0] _T_63025; // @[Modules.scala 50:57:@10177.4]
  wire [10:0] buffer_2_488; // @[Modules.scala 50:57:@10178.4]
  wire [10:0] buffer_2_194; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63027; // @[Modules.scala 50:57:@10180.4]
  wire [10:0] _T_63028; // @[Modules.scala 50:57:@10181.4]
  wire [10:0] buffer_2_489; // @[Modules.scala 50:57:@10182.4]
  wire [10:0] buffer_2_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63042; // @[Modules.scala 50:57:@10200.4]
  wire [10:0] _T_63043; // @[Modules.scala 50:57:@10201.4]
  wire [10:0] buffer_2_494; // @[Modules.scala 50:57:@10202.4]
  wire [10:0] buffer_2_208; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63048; // @[Modules.scala 50:57:@10208.4]
  wire [10:0] _T_63049; // @[Modules.scala 50:57:@10209.4]
  wire [10:0] buffer_2_496; // @[Modules.scala 50:57:@10210.4]
  wire [10:0] buffer_2_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63051; // @[Modules.scala 50:57:@10212.4]
  wire [10:0] _T_63052; // @[Modules.scala 50:57:@10213.4]
  wire [10:0] buffer_2_497; // @[Modules.scala 50:57:@10214.4]
  wire [10:0] buffer_2_212; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63054; // @[Modules.scala 50:57:@10216.4]
  wire [10:0] _T_63055; // @[Modules.scala 50:57:@10217.4]
  wire [10:0] buffer_2_498; // @[Modules.scala 50:57:@10218.4]
  wire [10:0] buffer_2_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63057; // @[Modules.scala 50:57:@10220.4]
  wire [10:0] _T_63058; // @[Modules.scala 50:57:@10221.4]
  wire [10:0] buffer_2_499; // @[Modules.scala 50:57:@10222.4]
  wire [10:0] buffer_2_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63063; // @[Modules.scala 50:57:@10228.4]
  wire [10:0] _T_63064; // @[Modules.scala 50:57:@10229.4]
  wire [10:0] buffer_2_501; // @[Modules.scala 50:57:@10230.4]
  wire [10:0] buffer_2_220; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63066; // @[Modules.scala 50:57:@10232.4]
  wire [10:0] _T_63067; // @[Modules.scala 50:57:@10233.4]
  wire [10:0] buffer_2_502; // @[Modules.scala 50:57:@10234.4]
  wire [11:0] _T_63072; // @[Modules.scala 50:57:@10240.4]
  wire [10:0] _T_63073; // @[Modules.scala 50:57:@10241.4]
  wire [10:0] buffer_2_504; // @[Modules.scala 50:57:@10242.4]
  wire [10:0] buffer_2_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63075; // @[Modules.scala 50:57:@10244.4]
  wire [10:0] _T_63076; // @[Modules.scala 50:57:@10245.4]
  wire [10:0] buffer_2_505; // @[Modules.scala 50:57:@10246.4]
  wire [10:0] buffer_2_228; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63078; // @[Modules.scala 50:57:@10248.4]
  wire [10:0] _T_63079; // @[Modules.scala 50:57:@10249.4]
  wire [10:0] buffer_2_506; // @[Modules.scala 50:57:@10250.4]
  wire [10:0] buffer_2_230; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63081; // @[Modules.scala 50:57:@10252.4]
  wire [10:0] _T_63082; // @[Modules.scala 50:57:@10253.4]
  wire [10:0] buffer_2_507; // @[Modules.scala 50:57:@10254.4]
  wire [10:0] buffer_2_232; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63084; // @[Modules.scala 50:57:@10256.4]
  wire [10:0] _T_63085; // @[Modules.scala 50:57:@10257.4]
  wire [10:0] buffer_2_508; // @[Modules.scala 50:57:@10258.4]
  wire [10:0] buffer_2_234; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63087; // @[Modules.scala 50:57:@10260.4]
  wire [10:0] _T_63088; // @[Modules.scala 50:57:@10261.4]
  wire [10:0] buffer_2_509; // @[Modules.scala 50:57:@10262.4]
  wire [10:0] buffer_2_238; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63093; // @[Modules.scala 50:57:@10268.4]
  wire [10:0] _T_63094; // @[Modules.scala 50:57:@10269.4]
  wire [10:0] buffer_2_511; // @[Modules.scala 50:57:@10270.4]
  wire [10:0] buffer_2_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63096; // @[Modules.scala 50:57:@10272.4]
  wire [10:0] _T_63097; // @[Modules.scala 50:57:@10273.4]
  wire [10:0] buffer_2_512; // @[Modules.scala 50:57:@10274.4]
  wire [10:0] buffer_2_242; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63099; // @[Modules.scala 50:57:@10276.4]
  wire [10:0] _T_63100; // @[Modules.scala 50:57:@10277.4]
  wire [10:0] buffer_2_513; // @[Modules.scala 50:57:@10278.4]
  wire [10:0] buffer_2_244; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63102; // @[Modules.scala 50:57:@10280.4]
  wire [10:0] _T_63103; // @[Modules.scala 50:57:@10281.4]
  wire [10:0] buffer_2_514; // @[Modules.scala 50:57:@10282.4]
  wire [10:0] buffer_2_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63108; // @[Modules.scala 50:57:@10288.4]
  wire [10:0] _T_63109; // @[Modules.scala 50:57:@10289.4]
  wire [10:0] buffer_2_516; // @[Modules.scala 50:57:@10290.4]
  wire [10:0] buffer_2_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63114; // @[Modules.scala 50:57:@10296.4]
  wire [10:0] _T_63115; // @[Modules.scala 50:57:@10297.4]
  wire [10:0] buffer_2_518; // @[Modules.scala 50:57:@10298.4]
  wire [10:0] buffer_2_258; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63123; // @[Modules.scala 50:57:@10308.4]
  wire [10:0] _T_63124; // @[Modules.scala 50:57:@10309.4]
  wire [10:0] buffer_2_521; // @[Modules.scala 50:57:@10310.4]
  wire [10:0] buffer_2_260; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63126; // @[Modules.scala 50:57:@10312.4]
  wire [10:0] _T_63127; // @[Modules.scala 50:57:@10313.4]
  wire [10:0] buffer_2_522; // @[Modules.scala 50:57:@10314.4]
  wire [10:0] buffer_2_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63129; // @[Modules.scala 50:57:@10316.4]
  wire [10:0] _T_63130; // @[Modules.scala 50:57:@10317.4]
  wire [10:0] buffer_2_523; // @[Modules.scala 50:57:@10318.4]
  wire [10:0] buffer_2_266; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_267; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63135; // @[Modules.scala 50:57:@10324.4]
  wire [10:0] _T_63136; // @[Modules.scala 50:57:@10325.4]
  wire [10:0] buffer_2_525; // @[Modules.scala 50:57:@10326.4]
  wire [10:0] buffer_2_272; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63144; // @[Modules.scala 50:57:@10336.4]
  wire [10:0] _T_63145; // @[Modules.scala 50:57:@10337.4]
  wire [10:0] buffer_2_528; // @[Modules.scala 50:57:@10338.4]
  wire [10:0] buffer_2_274; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63147; // @[Modules.scala 50:57:@10340.4]
  wire [10:0] _T_63148; // @[Modules.scala 50:57:@10341.4]
  wire [10:0] buffer_2_529; // @[Modules.scala 50:57:@10342.4]
  wire [10:0] buffer_2_276; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63150; // @[Modules.scala 50:57:@10344.4]
  wire [10:0] _T_63151; // @[Modules.scala 50:57:@10345.4]
  wire [10:0] buffer_2_530; // @[Modules.scala 50:57:@10346.4]
  wire [11:0] _T_63153; // @[Modules.scala 50:57:@10348.4]
  wire [10:0] _T_63154; // @[Modules.scala 50:57:@10349.4]
  wire [10:0] buffer_2_531; // @[Modules.scala 50:57:@10350.4]
  wire [10:0] buffer_2_280; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63156; // @[Modules.scala 50:57:@10352.4]
  wire [10:0] _T_63157; // @[Modules.scala 50:57:@10353.4]
  wire [10:0] buffer_2_532; // @[Modules.scala 50:57:@10354.4]
  wire [10:0] buffer_2_286; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63165; // @[Modules.scala 50:57:@10364.4]
  wire [10:0] _T_63166; // @[Modules.scala 50:57:@10365.4]
  wire [10:0] buffer_2_535; // @[Modules.scala 50:57:@10366.4]
  wire [11:0] _T_63168; // @[Modules.scala 50:57:@10368.4]
  wire [10:0] _T_63169; // @[Modules.scala 50:57:@10369.4]
  wire [10:0] buffer_2_536; // @[Modules.scala 50:57:@10370.4]
  wire [10:0] buffer_2_290; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63171; // @[Modules.scala 50:57:@10372.4]
  wire [10:0] _T_63172; // @[Modules.scala 50:57:@10373.4]
  wire [10:0] buffer_2_537; // @[Modules.scala 50:57:@10374.4]
  wire [10:0] buffer_2_294; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_295; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63177; // @[Modules.scala 50:57:@10380.4]
  wire [10:0] _T_63178; // @[Modules.scala 50:57:@10381.4]
  wire [10:0] buffer_2_539; // @[Modules.scala 50:57:@10382.4]
  wire [10:0] buffer_2_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63180; // @[Modules.scala 50:57:@10384.4]
  wire [10:0] _T_63181; // @[Modules.scala 50:57:@10385.4]
  wire [10:0] buffer_2_540; // @[Modules.scala 50:57:@10386.4]
  wire [10:0] buffer_2_298; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63183; // @[Modules.scala 50:57:@10388.4]
  wire [10:0] _T_63184; // @[Modules.scala 50:57:@10389.4]
  wire [10:0] buffer_2_541; // @[Modules.scala 50:57:@10390.4]
  wire [10:0] buffer_2_300; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63186; // @[Modules.scala 50:57:@10392.4]
  wire [10:0] _T_63187; // @[Modules.scala 50:57:@10393.4]
  wire [10:0] buffer_2_542; // @[Modules.scala 50:57:@10394.4]
  wire [10:0] buffer_2_302; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_303; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63189; // @[Modules.scala 50:57:@10396.4]
  wire [10:0] _T_63190; // @[Modules.scala 50:57:@10397.4]
  wire [10:0] buffer_2_543; // @[Modules.scala 50:57:@10398.4]
  wire [10:0] buffer_2_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63192; // @[Modules.scala 50:57:@10400.4]
  wire [10:0] _T_63193; // @[Modules.scala 50:57:@10401.4]
  wire [10:0] buffer_2_544; // @[Modules.scala 50:57:@10402.4]
  wire [10:0] buffer_2_308; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63198; // @[Modules.scala 50:57:@10408.4]
  wire [10:0] _T_63199; // @[Modules.scala 50:57:@10409.4]
  wire [10:0] buffer_2_546; // @[Modules.scala 50:57:@10410.4]
  wire [10:0] buffer_2_312; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63204; // @[Modules.scala 50:57:@10416.4]
  wire [10:0] _T_63205; // @[Modules.scala 50:57:@10417.4]
  wire [10:0] buffer_2_548; // @[Modules.scala 50:57:@10418.4]
  wire [10:0] buffer_2_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63210; // @[Modules.scala 50:57:@10424.4]
  wire [10:0] _T_63211; // @[Modules.scala 50:57:@10425.4]
  wire [10:0] buffer_2_550; // @[Modules.scala 50:57:@10426.4]
  wire [10:0] buffer_2_322; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_323; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63219; // @[Modules.scala 50:57:@10436.4]
  wire [10:0] _T_63220; // @[Modules.scala 50:57:@10437.4]
  wire [10:0] buffer_2_553; // @[Modules.scala 50:57:@10438.4]
  wire [10:0] buffer_2_324; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63222; // @[Modules.scala 50:57:@10440.4]
  wire [10:0] _T_63223; // @[Modules.scala 50:57:@10441.4]
  wire [10:0] buffer_2_554; // @[Modules.scala 50:57:@10442.4]
  wire [11:0] _T_63225; // @[Modules.scala 50:57:@10444.4]
  wire [10:0] _T_63226; // @[Modules.scala 50:57:@10445.4]
  wire [10:0] buffer_2_555; // @[Modules.scala 50:57:@10446.4]
  wire [10:0] buffer_2_328; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63228; // @[Modules.scala 50:57:@10448.4]
  wire [10:0] _T_63229; // @[Modules.scala 50:57:@10449.4]
  wire [10:0] buffer_2_556; // @[Modules.scala 50:57:@10450.4]
  wire [10:0] buffer_2_330; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63231; // @[Modules.scala 50:57:@10452.4]
  wire [10:0] _T_63232; // @[Modules.scala 50:57:@10453.4]
  wire [10:0] buffer_2_557; // @[Modules.scala 50:57:@10454.4]
  wire [10:0] buffer_2_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63237; // @[Modules.scala 50:57:@10460.4]
  wire [10:0] _T_63238; // @[Modules.scala 50:57:@10461.4]
  wire [10:0] buffer_2_559; // @[Modules.scala 50:57:@10462.4]
  wire [11:0] _T_63240; // @[Modules.scala 50:57:@10464.4]
  wire [10:0] _T_63241; // @[Modules.scala 50:57:@10465.4]
  wire [10:0] buffer_2_560; // @[Modules.scala 50:57:@10466.4]
  wire [10:0] buffer_2_338; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63243; // @[Modules.scala 50:57:@10468.4]
  wire [10:0] _T_63244; // @[Modules.scala 50:57:@10469.4]
  wire [10:0] buffer_2_561; // @[Modules.scala 50:57:@10470.4]
  wire [10:0] buffer_2_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63246; // @[Modules.scala 50:57:@10472.4]
  wire [10:0] _T_63247; // @[Modules.scala 50:57:@10473.4]
  wire [10:0] buffer_2_562; // @[Modules.scala 50:57:@10474.4]
  wire [10:0] buffer_2_342; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63249; // @[Modules.scala 50:57:@10476.4]
  wire [10:0] _T_63250; // @[Modules.scala 50:57:@10477.4]
  wire [10:0] buffer_2_563; // @[Modules.scala 50:57:@10478.4]
  wire [10:0] buffer_2_344; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63252; // @[Modules.scala 50:57:@10480.4]
  wire [10:0] _T_63253; // @[Modules.scala 50:57:@10481.4]
  wire [10:0] buffer_2_564; // @[Modules.scala 50:57:@10482.4]
  wire [10:0] buffer_2_348; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63258; // @[Modules.scala 50:57:@10488.4]
  wire [10:0] _T_63259; // @[Modules.scala 50:57:@10489.4]
  wire [10:0] buffer_2_566; // @[Modules.scala 50:57:@10490.4]
  wire [10:0] buffer_2_350; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63261; // @[Modules.scala 50:57:@10492.4]
  wire [10:0] _T_63262; // @[Modules.scala 50:57:@10493.4]
  wire [10:0] buffer_2_567; // @[Modules.scala 50:57:@10494.4]
  wire [10:0] buffer_2_352; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_353; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63264; // @[Modules.scala 50:57:@10496.4]
  wire [10:0] _T_63265; // @[Modules.scala 50:57:@10497.4]
  wire [10:0] buffer_2_568; // @[Modules.scala 50:57:@10498.4]
  wire [10:0] buffer_2_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63267; // @[Modules.scala 50:57:@10500.4]
  wire [10:0] _T_63268; // @[Modules.scala 50:57:@10501.4]
  wire [10:0] buffer_2_569; // @[Modules.scala 50:57:@10502.4]
  wire [10:0] buffer_2_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63270; // @[Modules.scala 50:57:@10504.4]
  wire [10:0] _T_63271; // @[Modules.scala 50:57:@10505.4]
  wire [10:0] buffer_2_570; // @[Modules.scala 50:57:@10506.4]
  wire [10:0] buffer_2_358; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63273; // @[Modules.scala 50:57:@10508.4]
  wire [10:0] _T_63274; // @[Modules.scala 50:57:@10509.4]
  wire [10:0] buffer_2_571; // @[Modules.scala 50:57:@10510.4]
  wire [10:0] buffer_2_364; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63282; // @[Modules.scala 50:57:@10520.4]
  wire [10:0] _T_63283; // @[Modules.scala 50:57:@10521.4]
  wire [10:0] buffer_2_574; // @[Modules.scala 50:57:@10522.4]
  wire [10:0] buffer_2_366; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63285; // @[Modules.scala 50:57:@10524.4]
  wire [10:0] _T_63286; // @[Modules.scala 50:57:@10525.4]
  wire [10:0] buffer_2_575; // @[Modules.scala 50:57:@10526.4]
  wire [10:0] buffer_2_374; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63297; // @[Modules.scala 50:57:@10540.4]
  wire [10:0] _T_63298; // @[Modules.scala 50:57:@10541.4]
  wire [10:0] buffer_2_579; // @[Modules.scala 50:57:@10542.4]
  wire [10:0] buffer_2_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63300; // @[Modules.scala 50:57:@10544.4]
  wire [10:0] _T_63301; // @[Modules.scala 50:57:@10545.4]
  wire [10:0] buffer_2_580; // @[Modules.scala 50:57:@10546.4]
  wire [10:0] buffer_2_378; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63303; // @[Modules.scala 50:57:@10548.4]
  wire [10:0] _T_63304; // @[Modules.scala 50:57:@10549.4]
  wire [10:0] buffer_2_581; // @[Modules.scala 50:57:@10550.4]
  wire [10:0] buffer_2_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63321; // @[Modules.scala 50:57:@10572.4]
  wire [10:0] _T_63322; // @[Modules.scala 50:57:@10573.4]
  wire [10:0] buffer_2_587; // @[Modules.scala 50:57:@10574.4]
  wire [11:0] _T_63324; // @[Modules.scala 53:83:@10576.4]
  wire [10:0] _T_63325; // @[Modules.scala 53:83:@10577.4]
  wire [10:0] buffer_2_588; // @[Modules.scala 53:83:@10578.4]
  wire [11:0] _T_63327; // @[Modules.scala 53:83:@10580.4]
  wire [10:0] _T_63328; // @[Modules.scala 53:83:@10581.4]
  wire [10:0] buffer_2_589; // @[Modules.scala 53:83:@10582.4]
  wire [11:0] _T_63330; // @[Modules.scala 53:83:@10584.4]
  wire [10:0] _T_63331; // @[Modules.scala 53:83:@10585.4]
  wire [10:0] buffer_2_590; // @[Modules.scala 53:83:@10586.4]
  wire [11:0] _T_63333; // @[Modules.scala 53:83:@10588.4]
  wire [10:0] _T_63334; // @[Modules.scala 53:83:@10589.4]
  wire [10:0] buffer_2_591; // @[Modules.scala 53:83:@10590.4]
  wire [11:0] _T_63336; // @[Modules.scala 53:83:@10592.4]
  wire [10:0] _T_63337; // @[Modules.scala 53:83:@10593.4]
  wire [10:0] buffer_2_592; // @[Modules.scala 53:83:@10594.4]
  wire [11:0] _T_63339; // @[Modules.scala 53:83:@10596.4]
  wire [10:0] _T_63340; // @[Modules.scala 53:83:@10597.4]
  wire [10:0] buffer_2_593; // @[Modules.scala 53:83:@10598.4]
  wire [11:0] _T_63342; // @[Modules.scala 53:83:@10600.4]
  wire [10:0] _T_63343; // @[Modules.scala 53:83:@10601.4]
  wire [10:0] buffer_2_594; // @[Modules.scala 53:83:@10602.4]
  wire [11:0] _T_63345; // @[Modules.scala 53:83:@10604.4]
  wire [10:0] _T_63346; // @[Modules.scala 53:83:@10605.4]
  wire [10:0] buffer_2_595; // @[Modules.scala 53:83:@10606.4]
  wire [11:0] _T_63348; // @[Modules.scala 53:83:@10608.4]
  wire [10:0] _T_63349; // @[Modules.scala 53:83:@10609.4]
  wire [10:0] buffer_2_596; // @[Modules.scala 53:83:@10610.4]
  wire [11:0] _T_63351; // @[Modules.scala 53:83:@10612.4]
  wire [10:0] _T_63352; // @[Modules.scala 53:83:@10613.4]
  wire [10:0] buffer_2_597; // @[Modules.scala 53:83:@10614.4]
  wire [11:0] _T_63354; // @[Modules.scala 53:83:@10616.4]
  wire [10:0] _T_63355; // @[Modules.scala 53:83:@10617.4]
  wire [10:0] buffer_2_598; // @[Modules.scala 53:83:@10618.4]
  wire [11:0] _T_63357; // @[Modules.scala 53:83:@10620.4]
  wire [10:0] _T_63358; // @[Modules.scala 53:83:@10621.4]
  wire [10:0] buffer_2_599; // @[Modules.scala 53:83:@10622.4]
  wire [11:0] _T_63360; // @[Modules.scala 53:83:@10624.4]
  wire [10:0] _T_63361; // @[Modules.scala 53:83:@10625.4]
  wire [10:0] buffer_2_600; // @[Modules.scala 53:83:@10626.4]
  wire [11:0] _T_63363; // @[Modules.scala 53:83:@10628.4]
  wire [10:0] _T_63364; // @[Modules.scala 53:83:@10629.4]
  wire [10:0] buffer_2_601; // @[Modules.scala 53:83:@10630.4]
  wire [11:0] _T_63366; // @[Modules.scala 53:83:@10632.4]
  wire [10:0] _T_63367; // @[Modules.scala 53:83:@10633.4]
  wire [10:0] buffer_2_602; // @[Modules.scala 53:83:@10634.4]
  wire [11:0] _T_63372; // @[Modules.scala 53:83:@10640.4]
  wire [10:0] _T_63373; // @[Modules.scala 53:83:@10641.4]
  wire [10:0] buffer_2_604; // @[Modules.scala 53:83:@10642.4]
  wire [11:0] _T_63375; // @[Modules.scala 53:83:@10644.4]
  wire [10:0] _T_63376; // @[Modules.scala 53:83:@10645.4]
  wire [10:0] buffer_2_605; // @[Modules.scala 53:83:@10646.4]
  wire [11:0] _T_63378; // @[Modules.scala 53:83:@10648.4]
  wire [10:0] _T_63379; // @[Modules.scala 53:83:@10649.4]
  wire [10:0] buffer_2_606; // @[Modules.scala 53:83:@10650.4]
  wire [11:0] _T_63381; // @[Modules.scala 53:83:@10652.4]
  wire [10:0] _T_63382; // @[Modules.scala 53:83:@10653.4]
  wire [10:0] buffer_2_607; // @[Modules.scala 53:83:@10654.4]
  wire [11:0] _T_63384; // @[Modules.scala 53:83:@10656.4]
  wire [10:0] _T_63385; // @[Modules.scala 53:83:@10657.4]
  wire [10:0] buffer_2_608; // @[Modules.scala 53:83:@10658.4]
  wire [11:0] _T_63387; // @[Modules.scala 53:83:@10660.4]
  wire [10:0] _T_63388; // @[Modules.scala 53:83:@10661.4]
  wire [10:0] buffer_2_609; // @[Modules.scala 53:83:@10662.4]
  wire [11:0] _T_63393; // @[Modules.scala 53:83:@10668.4]
  wire [10:0] _T_63394; // @[Modules.scala 53:83:@10669.4]
  wire [10:0] buffer_2_611; // @[Modules.scala 53:83:@10670.4]
  wire [11:0] _T_63396; // @[Modules.scala 53:83:@10672.4]
  wire [10:0] _T_63397; // @[Modules.scala 53:83:@10673.4]
  wire [10:0] buffer_2_612; // @[Modules.scala 53:83:@10674.4]
  wire [11:0] _T_63399; // @[Modules.scala 53:83:@10676.4]
  wire [10:0] _T_63400; // @[Modules.scala 53:83:@10677.4]
  wire [10:0] buffer_2_613; // @[Modules.scala 53:83:@10678.4]
  wire [11:0] _T_63402; // @[Modules.scala 53:83:@10680.4]
  wire [10:0] _T_63403; // @[Modules.scala 53:83:@10681.4]
  wire [10:0] buffer_2_614; // @[Modules.scala 53:83:@10682.4]
  wire [11:0] _T_63405; // @[Modules.scala 53:83:@10684.4]
  wire [10:0] _T_63406; // @[Modules.scala 53:83:@10685.4]
  wire [10:0] buffer_2_615; // @[Modules.scala 53:83:@10686.4]
  wire [11:0] _T_63411; // @[Modules.scala 53:83:@10692.4]
  wire [10:0] _T_63412; // @[Modules.scala 53:83:@10693.4]
  wire [10:0] buffer_2_617; // @[Modules.scala 53:83:@10694.4]
  wire [11:0] _T_63414; // @[Modules.scala 53:83:@10696.4]
  wire [10:0] _T_63415; // @[Modules.scala 53:83:@10697.4]
  wire [10:0] buffer_2_618; // @[Modules.scala 53:83:@10698.4]
  wire [11:0] _T_63417; // @[Modules.scala 53:83:@10700.4]
  wire [10:0] _T_63418; // @[Modules.scala 53:83:@10701.4]
  wire [10:0] buffer_2_619; // @[Modules.scala 53:83:@10702.4]
  wire [11:0] _T_63420; // @[Modules.scala 53:83:@10704.4]
  wire [10:0] _T_63421; // @[Modules.scala 53:83:@10705.4]
  wire [10:0] buffer_2_620; // @[Modules.scala 53:83:@10706.4]
  wire [11:0] _T_63426; // @[Modules.scala 53:83:@10712.4]
  wire [10:0] _T_63427; // @[Modules.scala 53:83:@10713.4]
  wire [10:0] buffer_2_622; // @[Modules.scala 53:83:@10714.4]
  wire [11:0] _T_63429; // @[Modules.scala 53:83:@10716.4]
  wire [10:0] _T_63430; // @[Modules.scala 53:83:@10717.4]
  wire [10:0] buffer_2_623; // @[Modules.scala 53:83:@10718.4]
  wire [11:0] _T_63432; // @[Modules.scala 53:83:@10720.4]
  wire [10:0] _T_63433; // @[Modules.scala 53:83:@10721.4]
  wire [10:0] buffer_2_624; // @[Modules.scala 53:83:@10722.4]
  wire [11:0] _T_63438; // @[Modules.scala 53:83:@10728.4]
  wire [10:0] _T_63439; // @[Modules.scala 53:83:@10729.4]
  wire [10:0] buffer_2_626; // @[Modules.scala 53:83:@10730.4]
  wire [11:0] _T_63441; // @[Modules.scala 53:83:@10732.4]
  wire [10:0] _T_63442; // @[Modules.scala 53:83:@10733.4]
  wire [10:0] buffer_2_627; // @[Modules.scala 53:83:@10734.4]
  wire [11:0] _T_63444; // @[Modules.scala 53:83:@10736.4]
  wire [10:0] _T_63445; // @[Modules.scala 53:83:@10737.4]
  wire [10:0] buffer_2_628; // @[Modules.scala 53:83:@10738.4]
  wire [11:0] _T_63447; // @[Modules.scala 53:83:@10740.4]
  wire [10:0] _T_63448; // @[Modules.scala 53:83:@10741.4]
  wire [10:0] buffer_2_629; // @[Modules.scala 53:83:@10742.4]
  wire [11:0] _T_63456; // @[Modules.scala 53:83:@10752.4]
  wire [10:0] _T_63457; // @[Modules.scala 53:83:@10753.4]
  wire [10:0] buffer_2_632; // @[Modules.scala 53:83:@10754.4]
  wire [11:0] _T_63459; // @[Modules.scala 53:83:@10756.4]
  wire [10:0] _T_63460; // @[Modules.scala 53:83:@10757.4]
  wire [10:0] buffer_2_633; // @[Modules.scala 53:83:@10758.4]
  wire [11:0] _T_63468; // @[Modules.scala 53:83:@10768.4]
  wire [10:0] _T_63469; // @[Modules.scala 53:83:@10769.4]
  wire [10:0] buffer_2_636; // @[Modules.scala 53:83:@10770.4]
  wire [11:0] _T_63471; // @[Modules.scala 53:83:@10772.4]
  wire [10:0] _T_63472; // @[Modules.scala 53:83:@10773.4]
  wire [10:0] buffer_2_637; // @[Modules.scala 53:83:@10774.4]
  wire [11:0] _T_63477; // @[Modules.scala 53:83:@10780.4]
  wire [10:0] _T_63478; // @[Modules.scala 53:83:@10781.4]
  wire [10:0] buffer_2_639; // @[Modules.scala 53:83:@10782.4]
  wire [11:0] _T_63480; // @[Modules.scala 53:83:@10784.4]
  wire [10:0] _T_63481; // @[Modules.scala 53:83:@10785.4]
  wire [10:0] buffer_2_640; // @[Modules.scala 53:83:@10786.4]
  wire [11:0] _T_63483; // @[Modules.scala 53:83:@10788.4]
  wire [10:0] _T_63484; // @[Modules.scala 53:83:@10789.4]
  wire [10:0] buffer_2_641; // @[Modules.scala 53:83:@10790.4]
  wire [11:0] _T_63486; // @[Modules.scala 53:83:@10792.4]
  wire [10:0] _T_63487; // @[Modules.scala 53:83:@10793.4]
  wire [10:0] buffer_2_642; // @[Modules.scala 53:83:@10794.4]
  wire [11:0] _T_63489; // @[Modules.scala 53:83:@10796.4]
  wire [10:0] _T_63490; // @[Modules.scala 53:83:@10797.4]
  wire [10:0] buffer_2_643; // @[Modules.scala 53:83:@10798.4]
  wire [11:0] _T_63492; // @[Modules.scala 53:83:@10800.4]
  wire [10:0] _T_63493; // @[Modules.scala 53:83:@10801.4]
  wire [10:0] buffer_2_644; // @[Modules.scala 53:83:@10802.4]
  wire [11:0] _T_63495; // @[Modules.scala 53:83:@10804.4]
  wire [10:0] _T_63496; // @[Modules.scala 53:83:@10805.4]
  wire [10:0] buffer_2_645; // @[Modules.scala 53:83:@10806.4]
  wire [11:0] _T_63498; // @[Modules.scala 53:83:@10808.4]
  wire [10:0] _T_63499; // @[Modules.scala 53:83:@10809.4]
  wire [10:0] buffer_2_646; // @[Modules.scala 53:83:@10810.4]
  wire [11:0] _T_63501; // @[Modules.scala 53:83:@10812.4]
  wire [10:0] _T_63502; // @[Modules.scala 53:83:@10813.4]
  wire [10:0] buffer_2_647; // @[Modules.scala 53:83:@10814.4]
  wire [11:0] _T_63504; // @[Modules.scala 53:83:@10816.4]
  wire [10:0] _T_63505; // @[Modules.scala 53:83:@10817.4]
  wire [10:0] buffer_2_648; // @[Modules.scala 53:83:@10818.4]
  wire [11:0] _T_63507; // @[Modules.scala 53:83:@10820.4]
  wire [10:0] _T_63508; // @[Modules.scala 53:83:@10821.4]
  wire [10:0] buffer_2_649; // @[Modules.scala 53:83:@10822.4]
  wire [11:0] _T_63510; // @[Modules.scala 53:83:@10824.4]
  wire [10:0] _T_63511; // @[Modules.scala 53:83:@10825.4]
  wire [10:0] buffer_2_650; // @[Modules.scala 53:83:@10826.4]
  wire [11:0] _T_63513; // @[Modules.scala 53:83:@10828.4]
  wire [10:0] _T_63514; // @[Modules.scala 53:83:@10829.4]
  wire [10:0] buffer_2_651; // @[Modules.scala 53:83:@10830.4]
  wire [11:0] _T_63516; // @[Modules.scala 53:83:@10832.4]
  wire [10:0] _T_63517; // @[Modules.scala 53:83:@10833.4]
  wire [10:0] buffer_2_652; // @[Modules.scala 53:83:@10834.4]
  wire [11:0] _T_63519; // @[Modules.scala 53:83:@10836.4]
  wire [10:0] _T_63520; // @[Modules.scala 53:83:@10837.4]
  wire [10:0] buffer_2_653; // @[Modules.scala 53:83:@10838.4]
  wire [11:0] _T_63522; // @[Modules.scala 53:83:@10840.4]
  wire [10:0] _T_63523; // @[Modules.scala 53:83:@10841.4]
  wire [10:0] buffer_2_654; // @[Modules.scala 53:83:@10842.4]
  wire [11:0] _T_63528; // @[Modules.scala 53:83:@10848.4]
  wire [10:0] _T_63529; // @[Modules.scala 53:83:@10849.4]
  wire [10:0] buffer_2_656; // @[Modules.scala 53:83:@10850.4]
  wire [11:0] _T_63531; // @[Modules.scala 53:83:@10852.4]
  wire [10:0] _T_63532; // @[Modules.scala 53:83:@10853.4]
  wire [10:0] buffer_2_657; // @[Modules.scala 53:83:@10854.4]
  wire [11:0] _T_63534; // @[Modules.scala 53:83:@10856.4]
  wire [10:0] _T_63535; // @[Modules.scala 53:83:@10857.4]
  wire [10:0] buffer_2_658; // @[Modules.scala 53:83:@10858.4]
  wire [11:0] _T_63537; // @[Modules.scala 53:83:@10860.4]
  wire [10:0] _T_63538; // @[Modules.scala 53:83:@10861.4]
  wire [10:0] buffer_2_659; // @[Modules.scala 53:83:@10862.4]
  wire [11:0] _T_63540; // @[Modules.scala 53:83:@10864.4]
  wire [10:0] _T_63541; // @[Modules.scala 53:83:@10865.4]
  wire [10:0] buffer_2_660; // @[Modules.scala 53:83:@10866.4]
  wire [11:0] _T_63543; // @[Modules.scala 53:83:@10868.4]
  wire [10:0] _T_63544; // @[Modules.scala 53:83:@10869.4]
  wire [10:0] buffer_2_661; // @[Modules.scala 53:83:@10870.4]
  wire [11:0] _T_63546; // @[Modules.scala 53:83:@10872.4]
  wire [10:0] _T_63547; // @[Modules.scala 53:83:@10873.4]
  wire [10:0] buffer_2_662; // @[Modules.scala 53:83:@10874.4]
  wire [11:0] _T_63549; // @[Modules.scala 53:83:@10876.4]
  wire [10:0] _T_63550; // @[Modules.scala 53:83:@10877.4]
  wire [10:0] buffer_2_663; // @[Modules.scala 53:83:@10878.4]
  wire [11:0] _T_63552; // @[Modules.scala 53:83:@10880.4]
  wire [10:0] _T_63553; // @[Modules.scala 53:83:@10881.4]
  wire [10:0] buffer_2_664; // @[Modules.scala 53:83:@10882.4]
  wire [11:0] _T_63555; // @[Modules.scala 53:83:@10884.4]
  wire [10:0] _T_63556; // @[Modules.scala 53:83:@10885.4]
  wire [10:0] buffer_2_665; // @[Modules.scala 53:83:@10886.4]
  wire [11:0] _T_63558; // @[Modules.scala 53:83:@10888.4]
  wire [10:0] _T_63559; // @[Modules.scala 53:83:@10889.4]
  wire [10:0] buffer_2_666; // @[Modules.scala 53:83:@10890.4]
  wire [11:0] _T_63561; // @[Modules.scala 53:83:@10892.4]
  wire [10:0] _T_63562; // @[Modules.scala 53:83:@10893.4]
  wire [10:0] buffer_2_667; // @[Modules.scala 53:83:@10894.4]
  wire [11:0] _T_63564; // @[Modules.scala 53:83:@10896.4]
  wire [10:0] _T_63565; // @[Modules.scala 53:83:@10897.4]
  wire [10:0] buffer_2_668; // @[Modules.scala 53:83:@10898.4]
  wire [11:0] _T_63567; // @[Modules.scala 53:83:@10900.4]
  wire [10:0] _T_63568; // @[Modules.scala 53:83:@10901.4]
  wire [10:0] buffer_2_669; // @[Modules.scala 53:83:@10902.4]
  wire [11:0] _T_63570; // @[Modules.scala 53:83:@10904.4]
  wire [10:0] _T_63571; // @[Modules.scala 53:83:@10905.4]
  wire [10:0] buffer_2_670; // @[Modules.scala 53:83:@10906.4]
  wire [11:0] _T_63573; // @[Modules.scala 53:83:@10908.4]
  wire [10:0] _T_63574; // @[Modules.scala 53:83:@10909.4]
  wire [10:0] buffer_2_671; // @[Modules.scala 53:83:@10910.4]
  wire [11:0] _T_63576; // @[Modules.scala 53:83:@10912.4]
  wire [10:0] _T_63577; // @[Modules.scala 53:83:@10913.4]
  wire [10:0] buffer_2_672; // @[Modules.scala 53:83:@10914.4]
  wire [11:0] _T_63579; // @[Modules.scala 53:83:@10916.4]
  wire [10:0] _T_63580; // @[Modules.scala 53:83:@10917.4]
  wire [10:0] buffer_2_673; // @[Modules.scala 53:83:@10918.4]
  wire [11:0] _T_63582; // @[Modules.scala 53:83:@10920.4]
  wire [10:0] _T_63583; // @[Modules.scala 53:83:@10921.4]
  wire [10:0] buffer_2_674; // @[Modules.scala 53:83:@10922.4]
  wire [11:0] _T_63585; // @[Modules.scala 53:83:@10924.4]
  wire [10:0] _T_63586; // @[Modules.scala 53:83:@10925.4]
  wire [10:0] buffer_2_675; // @[Modules.scala 53:83:@10926.4]
  wire [11:0] _T_63588; // @[Modules.scala 53:83:@10928.4]
  wire [10:0] _T_63589; // @[Modules.scala 53:83:@10929.4]
  wire [10:0] buffer_2_676; // @[Modules.scala 53:83:@10930.4]
  wire [11:0] _T_63591; // @[Modules.scala 53:83:@10932.4]
  wire [10:0] _T_63592; // @[Modules.scala 53:83:@10933.4]
  wire [10:0] buffer_2_677; // @[Modules.scala 53:83:@10934.4]
  wire [11:0] _T_63597; // @[Modules.scala 53:83:@10940.4]
  wire [10:0] _T_63598; // @[Modules.scala 53:83:@10941.4]
  wire [10:0] buffer_2_679; // @[Modules.scala 53:83:@10942.4]
  wire [11:0] _T_63603; // @[Modules.scala 53:83:@10948.4]
  wire [10:0] _T_63604; // @[Modules.scala 53:83:@10949.4]
  wire [10:0] buffer_2_681; // @[Modules.scala 53:83:@10950.4]
  wire [11:0] _T_63606; // @[Modules.scala 53:83:@10952.4]
  wire [10:0] _T_63607; // @[Modules.scala 53:83:@10953.4]
  wire [10:0] buffer_2_682; // @[Modules.scala 53:83:@10954.4]
  wire [11:0] _T_63615; // @[Modules.scala 53:83:@10964.4]
  wire [10:0] _T_63616; // @[Modules.scala 53:83:@10965.4]
  wire [10:0] buffer_2_685; // @[Modules.scala 53:83:@10966.4]
  wire [11:0] _T_63618; // @[Modules.scala 56:109:@10968.4]
  wire [10:0] _T_63619; // @[Modules.scala 56:109:@10969.4]
  wire [10:0] buffer_2_686; // @[Modules.scala 56:109:@10970.4]
  wire [11:0] _T_63621; // @[Modules.scala 56:109:@10972.4]
  wire [10:0] _T_63622; // @[Modules.scala 56:109:@10973.4]
  wire [10:0] buffer_2_687; // @[Modules.scala 56:109:@10974.4]
  wire [11:0] _T_63624; // @[Modules.scala 56:109:@10976.4]
  wire [10:0] _T_63625; // @[Modules.scala 56:109:@10977.4]
  wire [10:0] buffer_2_688; // @[Modules.scala 56:109:@10978.4]
  wire [11:0] _T_63627; // @[Modules.scala 56:109:@10980.4]
  wire [10:0] _T_63628; // @[Modules.scala 56:109:@10981.4]
  wire [10:0] buffer_2_689; // @[Modules.scala 56:109:@10982.4]
  wire [11:0] _T_63630; // @[Modules.scala 56:109:@10984.4]
  wire [10:0] _T_63631; // @[Modules.scala 56:109:@10985.4]
  wire [10:0] buffer_2_690; // @[Modules.scala 56:109:@10986.4]
  wire [11:0] _T_63633; // @[Modules.scala 56:109:@10988.4]
  wire [10:0] _T_63634; // @[Modules.scala 56:109:@10989.4]
  wire [10:0] buffer_2_691; // @[Modules.scala 56:109:@10990.4]
  wire [11:0] _T_63636; // @[Modules.scala 56:109:@10992.4]
  wire [10:0] _T_63637; // @[Modules.scala 56:109:@10993.4]
  wire [10:0] buffer_2_692; // @[Modules.scala 56:109:@10994.4]
  wire [11:0] _T_63639; // @[Modules.scala 56:109:@10996.4]
  wire [10:0] _T_63640; // @[Modules.scala 56:109:@10997.4]
  wire [10:0] buffer_2_693; // @[Modules.scala 56:109:@10998.4]
  wire [11:0] _T_63642; // @[Modules.scala 56:109:@11000.4]
  wire [10:0] _T_63643; // @[Modules.scala 56:109:@11001.4]
  wire [10:0] buffer_2_694; // @[Modules.scala 56:109:@11002.4]
  wire [11:0] _T_63645; // @[Modules.scala 56:109:@11004.4]
  wire [10:0] _T_63646; // @[Modules.scala 56:109:@11005.4]
  wire [10:0] buffer_2_695; // @[Modules.scala 56:109:@11006.4]
  wire [11:0] _T_63648; // @[Modules.scala 56:109:@11008.4]
  wire [10:0] _T_63649; // @[Modules.scala 56:109:@11009.4]
  wire [10:0] buffer_2_696; // @[Modules.scala 56:109:@11010.4]
  wire [11:0] _T_63651; // @[Modules.scala 56:109:@11012.4]
  wire [10:0] _T_63652; // @[Modules.scala 56:109:@11013.4]
  wire [10:0] buffer_2_697; // @[Modules.scala 56:109:@11014.4]
  wire [11:0] _T_63654; // @[Modules.scala 56:109:@11016.4]
  wire [10:0] _T_63655; // @[Modules.scala 56:109:@11017.4]
  wire [10:0] buffer_2_698; // @[Modules.scala 56:109:@11018.4]
  wire [11:0] _T_63657; // @[Modules.scala 56:109:@11020.4]
  wire [10:0] _T_63658; // @[Modules.scala 56:109:@11021.4]
  wire [10:0] buffer_2_699; // @[Modules.scala 56:109:@11022.4]
  wire [11:0] _T_63660; // @[Modules.scala 56:109:@11024.4]
  wire [10:0] _T_63661; // @[Modules.scala 56:109:@11025.4]
  wire [10:0] buffer_2_700; // @[Modules.scala 56:109:@11026.4]
  wire [11:0] _T_63663; // @[Modules.scala 56:109:@11028.4]
  wire [10:0] _T_63664; // @[Modules.scala 56:109:@11029.4]
  wire [10:0] buffer_2_701; // @[Modules.scala 56:109:@11030.4]
  wire [11:0] _T_63666; // @[Modules.scala 56:109:@11032.4]
  wire [10:0] _T_63667; // @[Modules.scala 56:109:@11033.4]
  wire [10:0] buffer_2_702; // @[Modules.scala 56:109:@11034.4]
  wire [11:0] _T_63669; // @[Modules.scala 56:109:@11036.4]
  wire [10:0] _T_63670; // @[Modules.scala 56:109:@11037.4]
  wire [10:0] buffer_2_703; // @[Modules.scala 56:109:@11038.4]
  wire [11:0] _T_63672; // @[Modules.scala 56:109:@11040.4]
  wire [10:0] _T_63673; // @[Modules.scala 56:109:@11041.4]
  wire [10:0] buffer_2_704; // @[Modules.scala 56:109:@11042.4]
  wire [11:0] _T_63675; // @[Modules.scala 56:109:@11044.4]
  wire [10:0] _T_63676; // @[Modules.scala 56:109:@11045.4]
  wire [10:0] buffer_2_705; // @[Modules.scala 56:109:@11046.4]
  wire [11:0] _T_63678; // @[Modules.scala 56:109:@11048.4]
  wire [10:0] _T_63679; // @[Modules.scala 56:109:@11049.4]
  wire [10:0] buffer_2_706; // @[Modules.scala 56:109:@11050.4]
  wire [11:0] _T_63684; // @[Modules.scala 56:109:@11056.4]
  wire [10:0] _T_63685; // @[Modules.scala 56:109:@11057.4]
  wire [10:0] buffer_2_708; // @[Modules.scala 56:109:@11058.4]
  wire [11:0] _T_63687; // @[Modules.scala 56:109:@11060.4]
  wire [10:0] _T_63688; // @[Modules.scala 56:109:@11061.4]
  wire [10:0] buffer_2_709; // @[Modules.scala 56:109:@11062.4]
  wire [11:0] _T_63690; // @[Modules.scala 56:109:@11064.4]
  wire [10:0] _T_63691; // @[Modules.scala 56:109:@11065.4]
  wire [10:0] buffer_2_710; // @[Modules.scala 56:109:@11066.4]
  wire [11:0] _T_63693; // @[Modules.scala 56:109:@11068.4]
  wire [10:0] _T_63694; // @[Modules.scala 56:109:@11069.4]
  wire [10:0] buffer_2_711; // @[Modules.scala 56:109:@11070.4]
  wire [11:0] _T_63696; // @[Modules.scala 56:109:@11072.4]
  wire [10:0] _T_63697; // @[Modules.scala 56:109:@11073.4]
  wire [10:0] buffer_2_712; // @[Modules.scala 56:109:@11074.4]
  wire [11:0] _T_63699; // @[Modules.scala 56:109:@11076.4]
  wire [10:0] _T_63700; // @[Modules.scala 56:109:@11077.4]
  wire [10:0] buffer_2_713; // @[Modules.scala 56:109:@11078.4]
  wire [11:0] _T_63702; // @[Modules.scala 56:109:@11080.4]
  wire [10:0] _T_63703; // @[Modules.scala 56:109:@11081.4]
  wire [10:0] buffer_2_714; // @[Modules.scala 56:109:@11082.4]
  wire [11:0] _T_63705; // @[Modules.scala 56:109:@11084.4]
  wire [10:0] _T_63706; // @[Modules.scala 56:109:@11085.4]
  wire [10:0] buffer_2_715; // @[Modules.scala 56:109:@11086.4]
  wire [11:0] _T_63708; // @[Modules.scala 56:109:@11088.4]
  wire [10:0] _T_63709; // @[Modules.scala 56:109:@11089.4]
  wire [10:0] buffer_2_716; // @[Modules.scala 56:109:@11090.4]
  wire [11:0] _T_63711; // @[Modules.scala 56:109:@11092.4]
  wire [10:0] _T_63712; // @[Modules.scala 56:109:@11093.4]
  wire [10:0] buffer_2_717; // @[Modules.scala 56:109:@11094.4]
  wire [11:0] _T_63714; // @[Modules.scala 56:109:@11096.4]
  wire [10:0] _T_63715; // @[Modules.scala 56:109:@11097.4]
  wire [10:0] buffer_2_718; // @[Modules.scala 56:109:@11098.4]
  wire [11:0] _T_63717; // @[Modules.scala 56:109:@11100.4]
  wire [10:0] _T_63718; // @[Modules.scala 56:109:@11101.4]
  wire [10:0] buffer_2_719; // @[Modules.scala 56:109:@11102.4]
  wire [11:0] _T_63720; // @[Modules.scala 56:109:@11104.4]
  wire [10:0] _T_63721; // @[Modules.scala 56:109:@11105.4]
  wire [10:0] buffer_2_720; // @[Modules.scala 56:109:@11106.4]
  wire [11:0] _T_63723; // @[Modules.scala 56:109:@11108.4]
  wire [10:0] _T_63724; // @[Modules.scala 56:109:@11109.4]
  wire [10:0] buffer_2_721; // @[Modules.scala 56:109:@11110.4]
  wire [11:0] _T_63726; // @[Modules.scala 56:109:@11112.4]
  wire [10:0] _T_63727; // @[Modules.scala 56:109:@11113.4]
  wire [10:0] buffer_2_722; // @[Modules.scala 56:109:@11114.4]
  wire [11:0] _T_63729; // @[Modules.scala 56:109:@11116.4]
  wire [10:0] _T_63730; // @[Modules.scala 56:109:@11117.4]
  wire [10:0] buffer_2_723; // @[Modules.scala 56:109:@11118.4]
  wire [11:0] _T_63732; // @[Modules.scala 56:109:@11120.4]
  wire [10:0] _T_63733; // @[Modules.scala 56:109:@11121.4]
  wire [10:0] buffer_2_724; // @[Modules.scala 56:109:@11122.4]
  wire [11:0] _T_63735; // @[Modules.scala 56:109:@11124.4]
  wire [10:0] _T_63736; // @[Modules.scala 56:109:@11125.4]
  wire [10:0] buffer_2_725; // @[Modules.scala 56:109:@11126.4]
  wire [11:0] _T_63738; // @[Modules.scala 56:109:@11128.4]
  wire [10:0] _T_63739; // @[Modules.scala 56:109:@11129.4]
  wire [10:0] buffer_2_726; // @[Modules.scala 56:109:@11130.4]
  wire [11:0] _T_63741; // @[Modules.scala 56:109:@11132.4]
  wire [10:0] _T_63742; // @[Modules.scala 56:109:@11133.4]
  wire [10:0] buffer_2_727; // @[Modules.scala 56:109:@11134.4]
  wire [11:0] _T_63744; // @[Modules.scala 56:109:@11136.4]
  wire [10:0] _T_63745; // @[Modules.scala 56:109:@11137.4]
  wire [10:0] buffer_2_728; // @[Modules.scala 56:109:@11138.4]
  wire [11:0] _T_63747; // @[Modules.scala 56:109:@11140.4]
  wire [10:0] _T_63748; // @[Modules.scala 56:109:@11141.4]
  wire [10:0] buffer_2_729; // @[Modules.scala 56:109:@11142.4]
  wire [11:0] _T_63750; // @[Modules.scala 56:109:@11144.4]
  wire [10:0] _T_63751; // @[Modules.scala 56:109:@11145.4]
  wire [10:0] buffer_2_730; // @[Modules.scala 56:109:@11146.4]
  wire [11:0] _T_63753; // @[Modules.scala 56:109:@11148.4]
  wire [10:0] _T_63754; // @[Modules.scala 56:109:@11149.4]
  wire [10:0] buffer_2_731; // @[Modules.scala 56:109:@11150.4]
  wire [11:0] _T_63756; // @[Modules.scala 56:109:@11152.4]
  wire [10:0] _T_63757; // @[Modules.scala 56:109:@11153.4]
  wire [10:0] buffer_2_732; // @[Modules.scala 56:109:@11154.4]
  wire [11:0] _T_63759; // @[Modules.scala 56:109:@11156.4]
  wire [10:0] _T_63760; // @[Modules.scala 56:109:@11157.4]
  wire [10:0] buffer_2_733; // @[Modules.scala 56:109:@11158.4]
  wire [11:0] _T_63762; // @[Modules.scala 56:109:@11160.4]
  wire [10:0] _T_63763; // @[Modules.scala 56:109:@11161.4]
  wire [10:0] buffer_2_734; // @[Modules.scala 56:109:@11162.4]
  wire [11:0] _T_63765; // @[Modules.scala 63:156:@11165.4]
  wire [10:0] _T_63766; // @[Modules.scala 63:156:@11166.4]
  wire [10:0] buffer_2_736; // @[Modules.scala 63:156:@11167.4]
  wire [11:0] _T_63768; // @[Modules.scala 63:156:@11169.4]
  wire [10:0] _T_63769; // @[Modules.scala 63:156:@11170.4]
  wire [10:0] buffer_2_737; // @[Modules.scala 63:156:@11171.4]
  wire [11:0] _T_63771; // @[Modules.scala 63:156:@11173.4]
  wire [10:0] _T_63772; // @[Modules.scala 63:156:@11174.4]
  wire [10:0] buffer_2_738; // @[Modules.scala 63:156:@11175.4]
  wire [11:0] _T_63774; // @[Modules.scala 63:156:@11177.4]
  wire [10:0] _T_63775; // @[Modules.scala 63:156:@11178.4]
  wire [10:0] buffer_2_739; // @[Modules.scala 63:156:@11179.4]
  wire [11:0] _T_63777; // @[Modules.scala 63:156:@11181.4]
  wire [10:0] _T_63778; // @[Modules.scala 63:156:@11182.4]
  wire [10:0] buffer_2_740; // @[Modules.scala 63:156:@11183.4]
  wire [11:0] _T_63780; // @[Modules.scala 63:156:@11185.4]
  wire [10:0] _T_63781; // @[Modules.scala 63:156:@11186.4]
  wire [10:0] buffer_2_741; // @[Modules.scala 63:156:@11187.4]
  wire [11:0] _T_63783; // @[Modules.scala 63:156:@11189.4]
  wire [10:0] _T_63784; // @[Modules.scala 63:156:@11190.4]
  wire [10:0] buffer_2_742; // @[Modules.scala 63:156:@11191.4]
  wire [11:0] _T_63786; // @[Modules.scala 63:156:@11193.4]
  wire [10:0] _T_63787; // @[Modules.scala 63:156:@11194.4]
  wire [10:0] buffer_2_743; // @[Modules.scala 63:156:@11195.4]
  wire [11:0] _T_63789; // @[Modules.scala 63:156:@11197.4]
  wire [10:0] _T_63790; // @[Modules.scala 63:156:@11198.4]
  wire [10:0] buffer_2_744; // @[Modules.scala 63:156:@11199.4]
  wire [11:0] _T_63792; // @[Modules.scala 63:156:@11201.4]
  wire [10:0] _T_63793; // @[Modules.scala 63:156:@11202.4]
  wire [10:0] buffer_2_745; // @[Modules.scala 63:156:@11203.4]
  wire [11:0] _T_63795; // @[Modules.scala 63:156:@11205.4]
  wire [10:0] _T_63796; // @[Modules.scala 63:156:@11206.4]
  wire [10:0] buffer_2_746; // @[Modules.scala 63:156:@11207.4]
  wire [11:0] _T_63798; // @[Modules.scala 63:156:@11209.4]
  wire [10:0] _T_63799; // @[Modules.scala 63:156:@11210.4]
  wire [10:0] buffer_2_747; // @[Modules.scala 63:156:@11211.4]
  wire [11:0] _T_63801; // @[Modules.scala 63:156:@11213.4]
  wire [10:0] _T_63802; // @[Modules.scala 63:156:@11214.4]
  wire [10:0] buffer_2_748; // @[Modules.scala 63:156:@11215.4]
  wire [11:0] _T_63804; // @[Modules.scala 63:156:@11217.4]
  wire [10:0] _T_63805; // @[Modules.scala 63:156:@11218.4]
  wire [10:0] buffer_2_749; // @[Modules.scala 63:156:@11219.4]
  wire [11:0] _T_63807; // @[Modules.scala 63:156:@11221.4]
  wire [10:0] _T_63808; // @[Modules.scala 63:156:@11222.4]
  wire [10:0] buffer_2_750; // @[Modules.scala 63:156:@11223.4]
  wire [11:0] _T_63810; // @[Modules.scala 63:156:@11225.4]
  wire [10:0] _T_63811; // @[Modules.scala 63:156:@11226.4]
  wire [10:0] buffer_2_751; // @[Modules.scala 63:156:@11227.4]
  wire [11:0] _T_63813; // @[Modules.scala 63:156:@11229.4]
  wire [10:0] _T_63814; // @[Modules.scala 63:156:@11230.4]
  wire [10:0] buffer_2_752; // @[Modules.scala 63:156:@11231.4]
  wire [11:0] _T_63816; // @[Modules.scala 63:156:@11233.4]
  wire [10:0] _T_63817; // @[Modules.scala 63:156:@11234.4]
  wire [10:0] buffer_2_753; // @[Modules.scala 63:156:@11235.4]
  wire [11:0] _T_63819; // @[Modules.scala 63:156:@11237.4]
  wire [10:0] _T_63820; // @[Modules.scala 63:156:@11238.4]
  wire [10:0] buffer_2_754; // @[Modules.scala 63:156:@11239.4]
  wire [11:0] _T_63822; // @[Modules.scala 63:156:@11241.4]
  wire [10:0] _T_63823; // @[Modules.scala 63:156:@11242.4]
  wire [10:0] buffer_2_755; // @[Modules.scala 63:156:@11243.4]
  wire [11:0] _T_63825; // @[Modules.scala 63:156:@11245.4]
  wire [10:0] _T_63826; // @[Modules.scala 63:156:@11246.4]
  wire [10:0] buffer_2_756; // @[Modules.scala 63:156:@11247.4]
  wire [11:0] _T_63828; // @[Modules.scala 63:156:@11249.4]
  wire [10:0] _T_63829; // @[Modules.scala 63:156:@11250.4]
  wire [10:0] buffer_2_757; // @[Modules.scala 63:156:@11251.4]
  wire [11:0] _T_63831; // @[Modules.scala 63:156:@11253.4]
  wire [10:0] _T_63832; // @[Modules.scala 63:156:@11254.4]
  wire [10:0] buffer_2_758; // @[Modules.scala 63:156:@11255.4]
  wire [11:0] _T_63834; // @[Modules.scala 63:156:@11257.4]
  wire [10:0] _T_63835; // @[Modules.scala 63:156:@11258.4]
  wire [10:0] buffer_2_759; // @[Modules.scala 63:156:@11259.4]
  wire [11:0] _T_63837; // @[Modules.scala 63:156:@11261.4]
  wire [10:0] _T_63838; // @[Modules.scala 63:156:@11262.4]
  wire [10:0] buffer_2_760; // @[Modules.scala 63:156:@11263.4]
  wire [11:0] _T_63840; // @[Modules.scala 63:156:@11265.4]
  wire [10:0] _T_63841; // @[Modules.scala 63:156:@11266.4]
  wire [10:0] buffer_2_761; // @[Modules.scala 63:156:@11267.4]
  wire [11:0] _T_63843; // @[Modules.scala 63:156:@11269.4]
  wire [10:0] _T_63844; // @[Modules.scala 63:156:@11270.4]
  wire [10:0] buffer_2_762; // @[Modules.scala 63:156:@11271.4]
  wire [11:0] _T_63846; // @[Modules.scala 63:156:@11273.4]
  wire [10:0] _T_63847; // @[Modules.scala 63:156:@11274.4]
  wire [10:0] buffer_2_763; // @[Modules.scala 63:156:@11275.4]
  wire [11:0] _T_63849; // @[Modules.scala 63:156:@11277.4]
  wire [10:0] _T_63850; // @[Modules.scala 63:156:@11278.4]
  wire [10:0] buffer_2_764; // @[Modules.scala 63:156:@11279.4]
  wire [11:0] _T_63852; // @[Modules.scala 63:156:@11281.4]
  wire [10:0] _T_63853; // @[Modules.scala 63:156:@11282.4]
  wire [10:0] buffer_2_765; // @[Modules.scala 63:156:@11283.4]
  wire [11:0] _T_63855; // @[Modules.scala 63:156:@11285.4]
  wire [10:0] _T_63856; // @[Modules.scala 63:156:@11286.4]
  wire [10:0] buffer_2_766; // @[Modules.scala 63:156:@11287.4]
  wire [11:0] _T_63858; // @[Modules.scala 63:156:@11289.4]
  wire [10:0] _T_63859; // @[Modules.scala 63:156:@11290.4]
  wire [10:0] buffer_2_767; // @[Modules.scala 63:156:@11291.4]
  wire [11:0] _T_63861; // @[Modules.scala 63:156:@11293.4]
  wire [10:0] _T_63862; // @[Modules.scala 63:156:@11294.4]
  wire [10:0] buffer_2_768; // @[Modules.scala 63:156:@11295.4]
  wire [11:0] _T_63864; // @[Modules.scala 63:156:@11297.4]
  wire [10:0] _T_63865; // @[Modules.scala 63:156:@11298.4]
  wire [10:0] buffer_2_769; // @[Modules.scala 63:156:@11299.4]
  wire [11:0] _T_63867; // @[Modules.scala 63:156:@11301.4]
  wire [10:0] _T_63868; // @[Modules.scala 63:156:@11302.4]
  wire [10:0] buffer_2_770; // @[Modules.scala 63:156:@11303.4]
  wire [11:0] _T_63870; // @[Modules.scala 63:156:@11305.4]
  wire [10:0] _T_63871; // @[Modules.scala 63:156:@11306.4]
  wire [10:0] buffer_2_771; // @[Modules.scala 63:156:@11307.4]
  wire [11:0] _T_63873; // @[Modules.scala 63:156:@11309.4]
  wire [10:0] _T_63874; // @[Modules.scala 63:156:@11310.4]
  wire [10:0] buffer_2_772; // @[Modules.scala 63:156:@11311.4]
  wire [11:0] _T_63876; // @[Modules.scala 63:156:@11313.4]
  wire [10:0] _T_63877; // @[Modules.scala 63:156:@11314.4]
  wire [10:0] buffer_2_773; // @[Modules.scala 63:156:@11315.4]
  wire [11:0] _T_63879; // @[Modules.scala 63:156:@11317.4]
  wire [10:0] _T_63880; // @[Modules.scala 63:156:@11318.4]
  wire [10:0] buffer_2_774; // @[Modules.scala 63:156:@11319.4]
  wire [11:0] _T_63882; // @[Modules.scala 63:156:@11321.4]
  wire [10:0] _T_63883; // @[Modules.scala 63:156:@11322.4]
  wire [10:0] buffer_2_775; // @[Modules.scala 63:156:@11323.4]
  wire [11:0] _T_63885; // @[Modules.scala 63:156:@11325.4]
  wire [10:0] _T_63886; // @[Modules.scala 63:156:@11326.4]
  wire [10:0] buffer_2_776; // @[Modules.scala 63:156:@11327.4]
  wire [11:0] _T_63888; // @[Modules.scala 63:156:@11329.4]
  wire [10:0] _T_63889; // @[Modules.scala 63:156:@11330.4]
  wire [10:0] buffer_2_777; // @[Modules.scala 63:156:@11331.4]
  wire [11:0] _T_63891; // @[Modules.scala 63:156:@11333.4]
  wire [10:0] _T_63892; // @[Modules.scala 63:156:@11334.4]
  wire [10:0] buffer_2_778; // @[Modules.scala 63:156:@11335.4]
  wire [11:0] _T_63894; // @[Modules.scala 63:156:@11337.4]
  wire [10:0] _T_63895; // @[Modules.scala 63:156:@11338.4]
  wire [10:0] buffer_2_779; // @[Modules.scala 63:156:@11339.4]
  wire [11:0] _T_63897; // @[Modules.scala 63:156:@11341.4]
  wire [10:0] _T_63898; // @[Modules.scala 63:156:@11342.4]
  wire [10:0] buffer_2_780; // @[Modules.scala 63:156:@11343.4]
  wire [11:0] _T_63900; // @[Modules.scala 63:156:@11345.4]
  wire [10:0] _T_63901; // @[Modules.scala 63:156:@11346.4]
  wire [10:0] buffer_2_781; // @[Modules.scala 63:156:@11347.4]
  wire [11:0] _T_63903; // @[Modules.scala 63:156:@11349.4]
  wire [10:0] _T_63904; // @[Modules.scala 63:156:@11350.4]
  wire [10:0] buffer_2_782; // @[Modules.scala 63:156:@11351.4]
  wire [11:0] _T_63906; // @[Modules.scala 63:156:@11353.4]
  wire [10:0] _T_63907; // @[Modules.scala 63:156:@11354.4]
  wire [10:0] buffer_2_783; // @[Modules.scala 63:156:@11355.4]
  wire [5:0] _T_63909; // @[Modules.scala 40:46:@11358.4]
  wire [4:0] _T_63910; // @[Modules.scala 40:46:@11359.4]
  wire [4:0] _T_63911; // @[Modules.scala 40:46:@11360.4]
  wire [5:0] _T_63912; // @[Modules.scala 40:46:@11362.4]
  wire [4:0] _T_63913; // @[Modules.scala 40:46:@11363.4]
  wire [4:0] _T_63914; // @[Modules.scala 40:46:@11364.4]
  wire [5:0] _T_63925; // @[Modules.scala 46:47:@11377.4]
  wire [4:0] _T_63926; // @[Modules.scala 46:47:@11378.4]
  wire [4:0] _T_63927; // @[Modules.scala 46:47:@11379.4]
  wire [5:0] _T_63928; // @[Modules.scala 40:46:@11381.4]
  wire [4:0] _T_63929; // @[Modules.scala 40:46:@11382.4]
  wire [4:0] _T_63930; // @[Modules.scala 40:46:@11383.4]
  wire [5:0] _T_63957; // @[Modules.scala 40:46:@11415.4]
  wire [4:0] _T_63958; // @[Modules.scala 40:46:@11416.4]
  wire [4:0] _T_63959; // @[Modules.scala 40:46:@11417.4]
  wire [5:0] _T_63960; // @[Modules.scala 37:46:@11419.4]
  wire [4:0] _T_63961; // @[Modules.scala 37:46:@11420.4]
  wire [4:0] _T_63962; // @[Modules.scala 37:46:@11421.4]
  wire [5:0] _T_63963; // @[Modules.scala 37:46:@11423.4]
  wire [4:0] _T_63964; // @[Modules.scala 37:46:@11424.4]
  wire [4:0] _T_63965; // @[Modules.scala 37:46:@11425.4]
  wire [5:0] _T_63970; // @[Modules.scala 46:47:@11430.4]
  wire [4:0] _T_63971; // @[Modules.scala 46:47:@11431.4]
  wire [4:0] _T_63972; // @[Modules.scala 46:47:@11432.4]
  wire [5:0] _T_63973; // @[Modules.scala 40:46:@11434.4]
  wire [4:0] _T_63974; // @[Modules.scala 40:46:@11435.4]
  wire [4:0] _T_63975; // @[Modules.scala 40:46:@11436.4]
  wire [5:0] _T_64031; // @[Modules.scala 43:47:@11495.4]
  wire [4:0] _T_64032; // @[Modules.scala 43:47:@11496.4]
  wire [4:0] _T_64033; // @[Modules.scala 43:47:@11497.4]
  wire [5:0] _T_64038; // @[Modules.scala 46:47:@11502.4]
  wire [4:0] _T_64039; // @[Modules.scala 46:47:@11503.4]
  wire [4:0] _T_64040; // @[Modules.scala 46:47:@11504.4]
  wire [5:0] _T_64045; // @[Modules.scala 46:47:@11509.4]
  wire [4:0] _T_64046; // @[Modules.scala 46:47:@11510.4]
  wire [4:0] _T_64047; // @[Modules.scala 46:47:@11511.4]
  wire [5:0] _T_64048; // @[Modules.scala 40:46:@11513.4]
  wire [4:0] _T_64049; // @[Modules.scala 40:46:@11514.4]
  wire [4:0] _T_64050; // @[Modules.scala 40:46:@11515.4]
  wire [5:0] _T_64055; // @[Modules.scala 43:47:@11520.4]
  wire [4:0] _T_64056; // @[Modules.scala 43:47:@11521.4]
  wire [4:0] _T_64057; // @[Modules.scala 43:47:@11522.4]
  wire [5:0] _T_64069; // @[Modules.scala 46:47:@11534.4]
  wire [4:0] _T_64070; // @[Modules.scala 46:47:@11535.4]
  wire [4:0] _T_64071; // @[Modules.scala 46:47:@11536.4]
  wire [5:0] _T_64104; // @[Modules.scala 46:47:@11569.4]
  wire [4:0] _T_64105; // @[Modules.scala 46:47:@11570.4]
  wire [4:0] _T_64106; // @[Modules.scala 46:47:@11571.4]
  wire [5:0] _T_64108; // @[Modules.scala 46:37:@11573.4]
  wire [4:0] _T_64109; // @[Modules.scala 46:37:@11574.4]
  wire [4:0] _T_64110; // @[Modules.scala 46:37:@11575.4]
  wire [5:0] _T_64111; // @[Modules.scala 46:47:@11576.4]
  wire [4:0] _T_64112; // @[Modules.scala 46:47:@11577.4]
  wire [4:0] _T_64113; // @[Modules.scala 46:47:@11578.4]
  wire [5:0] _T_64115; // @[Modules.scala 46:37:@11580.4]
  wire [4:0] _T_64116; // @[Modules.scala 46:37:@11581.4]
  wire [4:0] _T_64117; // @[Modules.scala 46:37:@11582.4]
  wire [5:0] _T_64118; // @[Modules.scala 46:47:@11583.4]
  wire [4:0] _T_64119; // @[Modules.scala 46:47:@11584.4]
  wire [4:0] _T_64120; // @[Modules.scala 46:47:@11585.4]
  wire [5:0] _T_64130; // @[Modules.scala 40:46:@11599.4]
  wire [4:0] _T_64131; // @[Modules.scala 40:46:@11600.4]
  wire [4:0] _T_64132; // @[Modules.scala 40:46:@11601.4]
  wire [5:0] _T_64134; // @[Modules.scala 46:37:@11603.4]
  wire [4:0] _T_64135; // @[Modules.scala 46:37:@11604.4]
  wire [4:0] _T_64136; // @[Modules.scala 46:37:@11605.4]
  wire [5:0] _T_64137; // @[Modules.scala 46:47:@11606.4]
  wire [4:0] _T_64138; // @[Modules.scala 46:47:@11607.4]
  wire [4:0] _T_64139; // @[Modules.scala 46:47:@11608.4]
  wire [5:0] _T_64141; // @[Modules.scala 46:37:@11610.4]
  wire [4:0] _T_64142; // @[Modules.scala 46:37:@11611.4]
  wire [4:0] _T_64143; // @[Modules.scala 46:37:@11612.4]
  wire [5:0] _T_64144; // @[Modules.scala 46:47:@11613.4]
  wire [4:0] _T_64145; // @[Modules.scala 46:47:@11614.4]
  wire [4:0] _T_64146; // @[Modules.scala 46:47:@11615.4]
  wire [5:0] _T_64151; // @[Modules.scala 46:47:@11620.4]
  wire [4:0] _T_64152; // @[Modules.scala 46:47:@11621.4]
  wire [4:0] _T_64153; // @[Modules.scala 46:47:@11622.4]
  wire [5:0] _T_64160; // @[Modules.scala 40:46:@11632.4]
  wire [4:0] _T_64161; // @[Modules.scala 40:46:@11633.4]
  wire [4:0] _T_64162; // @[Modules.scala 40:46:@11634.4]
  wire [5:0] _T_64167; // @[Modules.scala 46:37:@11640.4]
  wire [4:0] _T_64168; // @[Modules.scala 46:37:@11641.4]
  wire [4:0] _T_64169; // @[Modules.scala 46:37:@11642.4]
  wire [5:0] _T_64170; // @[Modules.scala 46:47:@11643.4]
  wire [4:0] _T_64171; // @[Modules.scala 46:47:@11644.4]
  wire [4:0] _T_64172; // @[Modules.scala 46:47:@11645.4]
  wire [5:0] _T_64174; // @[Modules.scala 46:37:@11647.4]
  wire [4:0] _T_64175; // @[Modules.scala 46:37:@11648.4]
  wire [4:0] _T_64176; // @[Modules.scala 46:37:@11649.4]
  wire [5:0] _T_64177; // @[Modules.scala 46:47:@11650.4]
  wire [4:0] _T_64178; // @[Modules.scala 46:47:@11651.4]
  wire [4:0] _T_64179; // @[Modules.scala 46:47:@11652.4]
  wire [5:0] _T_64181; // @[Modules.scala 46:37:@11654.4]
  wire [4:0] _T_64182; // @[Modules.scala 46:37:@11655.4]
  wire [4:0] _T_64183; // @[Modules.scala 46:37:@11656.4]
  wire [5:0] _T_64184; // @[Modules.scala 46:47:@11657.4]
  wire [4:0] _T_64185; // @[Modules.scala 46:47:@11658.4]
  wire [4:0] _T_64186; // @[Modules.scala 46:47:@11659.4]
  wire [5:0] _T_64191; // @[Modules.scala 43:47:@11664.4]
  wire [4:0] _T_64192; // @[Modules.scala 43:47:@11665.4]
  wire [4:0] _T_64193; // @[Modules.scala 43:47:@11666.4]
  wire [5:0] _T_64194; // @[Modules.scala 40:46:@11668.4]
  wire [4:0] _T_64195; // @[Modules.scala 40:46:@11669.4]
  wire [4:0] _T_64196; // @[Modules.scala 40:46:@11670.4]
  wire [5:0] _T_64197; // @[Modules.scala 40:46:@11672.4]
  wire [4:0] _T_64198; // @[Modules.scala 40:46:@11673.4]
  wire [4:0] _T_64199; // @[Modules.scala 40:46:@11674.4]
  wire [5:0] _T_64200; // @[Modules.scala 37:46:@11676.4]
  wire [4:0] _T_64201; // @[Modules.scala 37:46:@11677.4]
  wire [4:0] _T_64202; // @[Modules.scala 37:46:@11678.4]
  wire [5:0] _T_64213; // @[Modules.scala 37:46:@11691.4]
  wire [4:0] _T_64214; // @[Modules.scala 37:46:@11692.4]
  wire [4:0] _T_64215; // @[Modules.scala 37:46:@11693.4]
  wire [5:0] _T_64216; // @[Modules.scala 37:46:@11695.4]
  wire [4:0] _T_64217; // @[Modules.scala 37:46:@11696.4]
  wire [4:0] _T_64218; // @[Modules.scala 37:46:@11697.4]
  wire [5:0] _T_64219; // @[Modules.scala 37:46:@11699.4]
  wire [4:0] _T_64220; // @[Modules.scala 37:46:@11700.4]
  wire [4:0] _T_64221; // @[Modules.scala 37:46:@11701.4]
  wire [5:0] _T_64222; // @[Modules.scala 37:46:@11703.4]
  wire [4:0] _T_64223; // @[Modules.scala 37:46:@11704.4]
  wire [4:0] _T_64224; // @[Modules.scala 37:46:@11705.4]
  wire [5:0] _T_64235; // @[Modules.scala 46:47:@11718.4]
  wire [4:0] _T_64236; // @[Modules.scala 46:47:@11719.4]
  wire [4:0] _T_64237; // @[Modules.scala 46:47:@11720.4]
  wire [5:0] _T_64238; // @[Modules.scala 40:46:@11722.4]
  wire [4:0] _T_64239; // @[Modules.scala 40:46:@11723.4]
  wire [4:0] _T_64240; // @[Modules.scala 40:46:@11724.4]
  wire [5:0] _T_64244; // @[Modules.scala 40:46:@11730.4]
  wire [4:0] _T_64245; // @[Modules.scala 40:46:@11731.4]
  wire [4:0] _T_64246; // @[Modules.scala 40:46:@11732.4]
  wire [5:0] _T_64261; // @[Modules.scala 43:47:@11748.4]
  wire [4:0] _T_64262; // @[Modules.scala 43:47:@11749.4]
  wire [4:0] _T_64263; // @[Modules.scala 43:47:@11750.4]
  wire [5:0] _T_64270; // @[Modules.scala 37:46:@11760.4]
  wire [4:0] _T_64271; // @[Modules.scala 37:46:@11761.4]
  wire [4:0] _T_64272; // @[Modules.scala 37:46:@11762.4]
  wire [5:0] _T_64277; // @[Modules.scala 43:47:@11767.4]
  wire [4:0] _T_64278; // @[Modules.scala 43:47:@11768.4]
  wire [4:0] _T_64279; // @[Modules.scala 43:47:@11769.4]
  wire [5:0] _T_64280; // @[Modules.scala 37:46:@11771.4]
  wire [4:0] _T_64281; // @[Modules.scala 37:46:@11772.4]
  wire [4:0] _T_64282; // @[Modules.scala 37:46:@11773.4]
  wire [5:0] _T_64286; // @[Modules.scala 37:46:@11779.4]
  wire [4:0] _T_64287; // @[Modules.scala 37:46:@11780.4]
  wire [4:0] _T_64288; // @[Modules.scala 37:46:@11781.4]
  wire [5:0] _T_64311; // @[Modules.scala 37:46:@11810.4]
  wire [4:0] _T_64312; // @[Modules.scala 37:46:@11811.4]
  wire [4:0] _T_64313; // @[Modules.scala 37:46:@11812.4]
  wire [5:0] _T_64320; // @[Modules.scala 37:46:@11822.4]
  wire [4:0] _T_64321; // @[Modules.scala 37:46:@11823.4]
  wire [4:0] _T_64322; // @[Modules.scala 37:46:@11824.4]
  wire [5:0] _T_64323; // @[Modules.scala 37:46:@11826.4]
  wire [4:0] _T_64324; // @[Modules.scala 37:46:@11827.4]
  wire [4:0] _T_64325; // @[Modules.scala 37:46:@11828.4]
  wire [5:0] _T_64333; // @[Modules.scala 40:46:@11837.4]
  wire [4:0] _T_64334; // @[Modules.scala 40:46:@11838.4]
  wire [4:0] _T_64335; // @[Modules.scala 40:46:@11839.4]
  wire [5:0] _T_64336; // @[Modules.scala 40:46:@11841.4]
  wire [4:0] _T_64337; // @[Modules.scala 40:46:@11842.4]
  wire [4:0] _T_64338; // @[Modules.scala 40:46:@11843.4]
  wire [5:0] _T_64352; // @[Modules.scala 43:37:@11861.4]
  wire [4:0] _T_64353; // @[Modules.scala 43:37:@11862.4]
  wire [4:0] _T_64354; // @[Modules.scala 43:37:@11863.4]
  wire [5:0] _T_64355; // @[Modules.scala 43:47:@11864.4]
  wire [4:0] _T_64356; // @[Modules.scala 43:47:@11865.4]
  wire [4:0] _T_64357; // @[Modules.scala 43:47:@11866.4]
  wire [5:0] _T_64358; // @[Modules.scala 37:46:@11868.4]
  wire [4:0] _T_64359; // @[Modules.scala 37:46:@11869.4]
  wire [4:0] _T_64360; // @[Modules.scala 37:46:@11870.4]
  wire [5:0] _T_64361; // @[Modules.scala 37:46:@11872.4]
  wire [4:0] _T_64362; // @[Modules.scala 37:46:@11873.4]
  wire [4:0] _T_64363; // @[Modules.scala 37:46:@11874.4]
  wire [5:0] _T_64374; // @[Modules.scala 37:46:@11887.4]
  wire [4:0] _T_64375; // @[Modules.scala 37:46:@11888.4]
  wire [4:0] _T_64376; // @[Modules.scala 37:46:@11889.4]
  wire [5:0] _T_64377; // @[Modules.scala 37:46:@11891.4]
  wire [4:0] _T_64378; // @[Modules.scala 37:46:@11892.4]
  wire [4:0] _T_64379; // @[Modules.scala 37:46:@11893.4]
  wire [5:0] _T_64380; // @[Modules.scala 40:46:@11895.4]
  wire [4:0] _T_64381; // @[Modules.scala 40:46:@11896.4]
  wire [4:0] _T_64382; // @[Modules.scala 40:46:@11897.4]
  wire [5:0] _T_64383; // @[Modules.scala 37:46:@11899.4]
  wire [4:0] _T_64384; // @[Modules.scala 37:46:@11900.4]
  wire [4:0] _T_64385; // @[Modules.scala 37:46:@11901.4]
  wire [5:0] _T_64396; // @[Modules.scala 40:46:@11914.4]
  wire [4:0] _T_64397; // @[Modules.scala 40:46:@11915.4]
  wire [4:0] _T_64398; // @[Modules.scala 40:46:@11916.4]
  wire [5:0] _T_64408; // @[Modules.scala 37:46:@11930.4]
  wire [4:0] _T_64409; // @[Modules.scala 37:46:@11931.4]
  wire [4:0] _T_64410; // @[Modules.scala 37:46:@11932.4]
  wire [5:0] _T_64411; // @[Modules.scala 37:46:@11934.4]
  wire [4:0] _T_64412; // @[Modules.scala 37:46:@11935.4]
  wire [4:0] _T_64413; // @[Modules.scala 37:46:@11936.4]
  wire [5:0] _T_64418; // @[Modules.scala 43:47:@11941.4]
  wire [4:0] _T_64419; // @[Modules.scala 43:47:@11942.4]
  wire [4:0] _T_64420; // @[Modules.scala 43:47:@11943.4]
  wire [5:0] _T_64421; // @[Modules.scala 40:46:@11945.4]
  wire [4:0] _T_64422; // @[Modules.scala 40:46:@11946.4]
  wire [4:0] _T_64423; // @[Modules.scala 40:46:@11947.4]
  wire [5:0] _T_64424; // @[Modules.scala 37:46:@11949.4]
  wire [4:0] _T_64425; // @[Modules.scala 37:46:@11950.4]
  wire [4:0] _T_64426; // @[Modules.scala 37:46:@11951.4]
  wire [5:0] _T_64427; // @[Modules.scala 37:46:@11953.4]
  wire [4:0] _T_64428; // @[Modules.scala 37:46:@11954.4]
  wire [4:0] _T_64429; // @[Modules.scala 37:46:@11955.4]
  wire [5:0] _T_64430; // @[Modules.scala 37:46:@11957.4]
  wire [4:0] _T_64431; // @[Modules.scala 37:46:@11958.4]
  wire [4:0] _T_64432; // @[Modules.scala 37:46:@11959.4]
  wire [5:0] _T_64436; // @[Modules.scala 37:46:@11965.4]
  wire [4:0] _T_64437; // @[Modules.scala 37:46:@11966.4]
  wire [4:0] _T_64438; // @[Modules.scala 37:46:@11967.4]
  wire [5:0] _T_64439; // @[Modules.scala 40:46:@11969.4]
  wire [4:0] _T_64440; // @[Modules.scala 40:46:@11970.4]
  wire [4:0] _T_64441; // @[Modules.scala 40:46:@11971.4]
  wire [5:0] _T_64442; // @[Modules.scala 37:46:@11973.4]
  wire [4:0] _T_64443; // @[Modules.scala 37:46:@11974.4]
  wire [4:0] _T_64444; // @[Modules.scala 37:46:@11975.4]
  wire [5:0] _T_64451; // @[Modules.scala 37:46:@11985.4]
  wire [4:0] _T_64452; // @[Modules.scala 37:46:@11986.4]
  wire [4:0] _T_64453; // @[Modules.scala 37:46:@11987.4]
  wire [5:0] _T_64454; // @[Modules.scala 37:46:@11989.4]
  wire [4:0] _T_64455; // @[Modules.scala 37:46:@11990.4]
  wire [4:0] _T_64456; // @[Modules.scala 37:46:@11991.4]
  wire [5:0] _T_64457; // @[Modules.scala 37:46:@11993.4]
  wire [4:0] _T_64458; // @[Modules.scala 37:46:@11994.4]
  wire [4:0] _T_64459; // @[Modules.scala 37:46:@11995.4]
  wire [5:0] _T_64481; // @[Modules.scala 37:46:@12018.4]
  wire [4:0] _T_64482; // @[Modules.scala 37:46:@12019.4]
  wire [4:0] _T_64483; // @[Modules.scala 37:46:@12020.4]
  wire [5:0] _T_64487; // @[Modules.scala 37:46:@12026.4]
  wire [4:0] _T_64488; // @[Modules.scala 37:46:@12027.4]
  wire [4:0] _T_64489; // @[Modules.scala 37:46:@12028.4]
  wire [5:0] _T_64490; // @[Modules.scala 37:46:@12030.4]
  wire [4:0] _T_64491; // @[Modules.scala 37:46:@12031.4]
  wire [4:0] _T_64492; // @[Modules.scala 37:46:@12032.4]
  wire [5:0] _T_64493; // @[Modules.scala 37:46:@12034.4]
  wire [4:0] _T_64494; // @[Modules.scala 37:46:@12035.4]
  wire [4:0] _T_64495; // @[Modules.scala 37:46:@12036.4]
  wire [5:0] _T_64496; // @[Modules.scala 37:46:@12038.4]
  wire [4:0] _T_64497; // @[Modules.scala 37:46:@12039.4]
  wire [4:0] _T_64498; // @[Modules.scala 37:46:@12040.4]
  wire [5:0] _T_64505; // @[Modules.scala 37:46:@12050.4]
  wire [4:0] _T_64506; // @[Modules.scala 37:46:@12051.4]
  wire [4:0] _T_64507; // @[Modules.scala 37:46:@12052.4]
  wire [5:0] _T_64508; // @[Modules.scala 37:46:@12054.4]
  wire [4:0] _T_64509; // @[Modules.scala 37:46:@12055.4]
  wire [4:0] _T_64510; // @[Modules.scala 37:46:@12056.4]
  wire [5:0] _T_64511; // @[Modules.scala 40:46:@12058.4]
  wire [4:0] _T_64512; // @[Modules.scala 40:46:@12059.4]
  wire [4:0] _T_64513; // @[Modules.scala 40:46:@12060.4]
  wire [5:0] _T_64525; // @[Modules.scala 46:47:@12072.4]
  wire [4:0] _T_64526; // @[Modules.scala 46:47:@12073.4]
  wire [4:0] _T_64527; // @[Modules.scala 46:47:@12074.4]
  wire [5:0] _T_64546; // @[Modules.scala 43:47:@12093.4]
  wire [4:0] _T_64547; // @[Modules.scala 43:47:@12094.4]
  wire [4:0] _T_64548; // @[Modules.scala 43:47:@12095.4]
  wire [5:0] _T_64549; // @[Modules.scala 37:46:@12097.4]
  wire [4:0] _T_64550; // @[Modules.scala 37:46:@12098.4]
  wire [4:0] _T_64551; // @[Modules.scala 37:46:@12099.4]
  wire [5:0] _T_64552; // @[Modules.scala 40:46:@12101.4]
  wire [4:0] _T_64553; // @[Modules.scala 40:46:@12102.4]
  wire [4:0] _T_64554; // @[Modules.scala 40:46:@12103.4]
  wire [5:0] _T_64555; // @[Modules.scala 40:46:@12105.4]
  wire [4:0] _T_64556; // @[Modules.scala 40:46:@12106.4]
  wire [4:0] _T_64557; // @[Modules.scala 40:46:@12107.4]
  wire [5:0] _T_64575; // @[Modules.scala 43:47:@12127.4]
  wire [4:0] _T_64576; // @[Modules.scala 43:47:@12128.4]
  wire [4:0] _T_64577; // @[Modules.scala 43:47:@12129.4]
  wire [5:0] _T_64578; // @[Modules.scala 37:46:@12131.4]
  wire [4:0] _T_64579; // @[Modules.scala 37:46:@12132.4]
  wire [4:0] _T_64580; // @[Modules.scala 37:46:@12133.4]
  wire [5:0] _T_64592; // @[Modules.scala 46:47:@12145.4]
  wire [4:0] _T_64593; // @[Modules.scala 46:47:@12146.4]
  wire [4:0] _T_64594; // @[Modules.scala 46:47:@12147.4]
  wire [5:0] _T_64603; // @[Modules.scala 46:37:@12156.4]
  wire [4:0] _T_64604; // @[Modules.scala 46:37:@12157.4]
  wire [4:0] _T_64605; // @[Modules.scala 46:37:@12158.4]
  wire [5:0] _T_64606; // @[Modules.scala 46:47:@12159.4]
  wire [4:0] _T_64607; // @[Modules.scala 46:47:@12160.4]
  wire [4:0] _T_64608; // @[Modules.scala 46:47:@12161.4]
  wire [5:0] _T_64658; // @[Modules.scala 40:46:@12212.4]
  wire [4:0] _T_64659; // @[Modules.scala 40:46:@12213.4]
  wire [4:0] _T_64660; // @[Modules.scala 40:46:@12214.4]
  wire [5:0] _T_64662; // @[Modules.scala 43:37:@12216.4]
  wire [4:0] _T_64663; // @[Modules.scala 43:37:@12217.4]
  wire [4:0] _T_64664; // @[Modules.scala 43:37:@12218.4]
  wire [5:0] _T_64665; // @[Modules.scala 43:47:@12219.4]
  wire [4:0] _T_64666; // @[Modules.scala 43:47:@12220.4]
  wire [4:0] _T_64667; // @[Modules.scala 43:47:@12221.4]
  wire [5:0] _T_64668; // @[Modules.scala 40:46:@12223.4]
  wire [4:0] _T_64669; // @[Modules.scala 40:46:@12224.4]
  wire [4:0] _T_64670; // @[Modules.scala 40:46:@12225.4]
  wire [5:0] _T_64675; // @[Modules.scala 46:47:@12230.4]
  wire [4:0] _T_64676; // @[Modules.scala 46:47:@12231.4]
  wire [4:0] _T_64677; // @[Modules.scala 46:47:@12232.4]
  wire [5:0] _T_64679; // @[Modules.scala 46:37:@12234.4]
  wire [4:0] _T_64680; // @[Modules.scala 46:37:@12235.4]
  wire [4:0] _T_64681; // @[Modules.scala 46:37:@12236.4]
  wire [5:0] _T_64682; // @[Modules.scala 46:47:@12237.4]
  wire [4:0] _T_64683; // @[Modules.scala 46:47:@12238.4]
  wire [4:0] _T_64684; // @[Modules.scala 46:47:@12239.4]
  wire [5:0] _T_64686; // @[Modules.scala 46:37:@12241.4]
  wire [4:0] _T_64687; // @[Modules.scala 46:37:@12242.4]
  wire [4:0] _T_64688; // @[Modules.scala 46:37:@12243.4]
  wire [5:0] _T_64689; // @[Modules.scala 46:47:@12244.4]
  wire [4:0] _T_64690; // @[Modules.scala 46:47:@12245.4]
  wire [4:0] _T_64691; // @[Modules.scala 46:47:@12246.4]
  wire [5:0] _T_64693; // @[Modules.scala 46:37:@12248.4]
  wire [4:0] _T_64694; // @[Modules.scala 46:37:@12249.4]
  wire [4:0] _T_64695; // @[Modules.scala 46:37:@12250.4]
  wire [5:0] _T_64696; // @[Modules.scala 46:47:@12251.4]
  wire [4:0] _T_64697; // @[Modules.scala 46:47:@12252.4]
  wire [4:0] _T_64698; // @[Modules.scala 46:47:@12253.4]
  wire [5:0] _T_64700; // @[Modules.scala 46:37:@12255.4]
  wire [4:0] _T_64701; // @[Modules.scala 46:37:@12256.4]
  wire [4:0] _T_64702; // @[Modules.scala 46:37:@12257.4]
  wire [5:0] _T_64703; // @[Modules.scala 46:47:@12258.4]
  wire [4:0] _T_64704; // @[Modules.scala 46:47:@12259.4]
  wire [4:0] _T_64705; // @[Modules.scala 46:47:@12260.4]
  wire [5:0] _T_64755; // @[Modules.scala 43:47:@12311.4]
  wire [4:0] _T_64756; // @[Modules.scala 43:47:@12312.4]
  wire [4:0] _T_64757; // @[Modules.scala 43:47:@12313.4]
  wire [5:0] _T_64758; // @[Modules.scala 40:46:@12315.4]
  wire [4:0] _T_64759; // @[Modules.scala 40:46:@12316.4]
  wire [4:0] _T_64760; // @[Modules.scala 40:46:@12317.4]
  wire [5:0] _T_64765; // @[Modules.scala 46:47:@12322.4]
  wire [4:0] _T_64766; // @[Modules.scala 46:47:@12323.4]
  wire [4:0] _T_64767; // @[Modules.scala 46:47:@12324.4]
  wire [5:0] _T_64769; // @[Modules.scala 46:37:@12326.4]
  wire [4:0] _T_64770; // @[Modules.scala 46:37:@12327.4]
  wire [4:0] _T_64771; // @[Modules.scala 46:37:@12328.4]
  wire [5:0] _T_64772; // @[Modules.scala 46:47:@12329.4]
  wire [4:0] _T_64773; // @[Modules.scala 46:47:@12330.4]
  wire [4:0] _T_64774; // @[Modules.scala 46:47:@12331.4]
  wire [5:0] _T_64776; // @[Modules.scala 46:37:@12333.4]
  wire [4:0] _T_64777; // @[Modules.scala 46:37:@12334.4]
  wire [4:0] _T_64778; // @[Modules.scala 46:37:@12335.4]
  wire [5:0] _T_64779; // @[Modules.scala 46:47:@12336.4]
  wire [4:0] _T_64780; // @[Modules.scala 46:47:@12337.4]
  wire [4:0] _T_64781; // @[Modules.scala 46:47:@12338.4]
  wire [5:0] _T_64783; // @[Modules.scala 43:37:@12340.4]
  wire [4:0] _T_64784; // @[Modules.scala 43:37:@12341.4]
  wire [4:0] _T_64785; // @[Modules.scala 43:37:@12342.4]
  wire [5:0] _T_64786; // @[Modules.scala 43:47:@12343.4]
  wire [4:0] _T_64787; // @[Modules.scala 43:47:@12344.4]
  wire [4:0] _T_64788; // @[Modules.scala 43:47:@12345.4]
  wire [5:0] _T_64790; // @[Modules.scala 46:37:@12347.4]
  wire [4:0] _T_64791; // @[Modules.scala 46:37:@12348.4]
  wire [4:0] _T_64792; // @[Modules.scala 46:37:@12349.4]
  wire [5:0] _T_64793; // @[Modules.scala 46:47:@12350.4]
  wire [4:0] _T_64794; // @[Modules.scala 46:47:@12351.4]
  wire [4:0] _T_64795; // @[Modules.scala 46:47:@12352.4]
  wire [5:0] _T_64807; // @[Modules.scala 43:47:@12364.4]
  wire [4:0] _T_64808; // @[Modules.scala 43:47:@12365.4]
  wire [4:0] _T_64809; // @[Modules.scala 43:47:@12366.4]
  wire [5:0] _T_64821; // @[Modules.scala 46:47:@12378.4]
  wire [4:0] _T_64822; // @[Modules.scala 46:47:@12379.4]
  wire [4:0] _T_64823; // @[Modules.scala 46:47:@12380.4]
  wire [5:0] _T_64838; // @[Modules.scala 37:46:@12396.4]
  wire [4:0] _T_64839; // @[Modules.scala 37:46:@12397.4]
  wire [4:0] _T_64840; // @[Modules.scala 37:46:@12398.4]
  wire [5:0] _T_64844; // @[Modules.scala 40:46:@12404.4]
  wire [4:0] _T_64845; // @[Modules.scala 40:46:@12405.4]
  wire [4:0] _T_64846; // @[Modules.scala 40:46:@12406.4]
  wire [5:0] _T_64851; // @[Modules.scala 46:47:@12411.4]
  wire [4:0] _T_64852; // @[Modules.scala 46:47:@12412.4]
  wire [4:0] _T_64853; // @[Modules.scala 46:47:@12413.4]
  wire [5:0] _T_64855; // @[Modules.scala 46:37:@12415.4]
  wire [4:0] _T_64856; // @[Modules.scala 46:37:@12416.4]
  wire [4:0] _T_64857; // @[Modules.scala 46:37:@12417.4]
  wire [5:0] _T_64858; // @[Modules.scala 46:47:@12418.4]
  wire [4:0] _T_64859; // @[Modules.scala 46:47:@12419.4]
  wire [4:0] _T_64860; // @[Modules.scala 46:47:@12420.4]
  wire [5:0] _T_64862; // @[Modules.scala 43:37:@12422.4]
  wire [4:0] _T_64863; // @[Modules.scala 43:37:@12423.4]
  wire [4:0] _T_64864; // @[Modules.scala 43:37:@12424.4]
  wire [5:0] _T_64865; // @[Modules.scala 43:47:@12425.4]
  wire [4:0] _T_64866; // @[Modules.scala 43:47:@12426.4]
  wire [4:0] _T_64867; // @[Modules.scala 43:47:@12427.4]
  wire [5:0] _T_64868; // @[Modules.scala 40:46:@12429.4]
  wire [4:0] _T_64869; // @[Modules.scala 40:46:@12430.4]
  wire [4:0] _T_64870; // @[Modules.scala 40:46:@12431.4]
  wire [5:0] _T_64872; // @[Modules.scala 46:37:@12433.4]
  wire [4:0] _T_64873; // @[Modules.scala 46:37:@12434.4]
  wire [4:0] _T_64874; // @[Modules.scala 46:37:@12435.4]
  wire [5:0] _T_64875; // @[Modules.scala 46:47:@12436.4]
  wire [4:0] _T_64876; // @[Modules.scala 46:47:@12437.4]
  wire [4:0] _T_64877; // @[Modules.scala 46:47:@12438.4]
  wire [5:0] _T_64886; // @[Modules.scala 46:37:@12447.4]
  wire [4:0] _T_64887; // @[Modules.scala 46:37:@12448.4]
  wire [4:0] _T_64888; // @[Modules.scala 46:37:@12449.4]
  wire [5:0] _T_64889; // @[Modules.scala 46:47:@12450.4]
  wire [4:0] _T_64890; // @[Modules.scala 46:47:@12451.4]
  wire [4:0] _T_64891; // @[Modules.scala 46:47:@12452.4]
  wire [5:0] _T_64892; // @[Modules.scala 40:46:@12454.4]
  wire [4:0] _T_64893; // @[Modules.scala 40:46:@12455.4]
  wire [4:0] _T_64894; // @[Modules.scala 40:46:@12456.4]
  wire [5:0] _T_64896; // @[Modules.scala 46:37:@12458.4]
  wire [4:0] _T_64897; // @[Modules.scala 46:37:@12459.4]
  wire [4:0] _T_64898; // @[Modules.scala 46:37:@12460.4]
  wire [5:0] _T_64899; // @[Modules.scala 46:47:@12461.4]
  wire [4:0] _T_64900; // @[Modules.scala 46:47:@12462.4]
  wire [4:0] _T_64901; // @[Modules.scala 46:47:@12463.4]
  wire [5:0] _T_64903; // @[Modules.scala 46:37:@12465.4]
  wire [4:0] _T_64904; // @[Modules.scala 46:37:@12466.4]
  wire [4:0] _T_64905; // @[Modules.scala 46:37:@12467.4]
  wire [5:0] _T_64906; // @[Modules.scala 46:47:@12468.4]
  wire [4:0] _T_64907; // @[Modules.scala 46:47:@12469.4]
  wire [4:0] _T_64908; // @[Modules.scala 46:47:@12470.4]
  wire [5:0] _T_64913; // @[Modules.scala 43:47:@12475.4]
  wire [4:0] _T_64914; // @[Modules.scala 43:47:@12476.4]
  wire [4:0] _T_64915; // @[Modules.scala 43:47:@12477.4]
  wire [5:0] _T_64916; // @[Modules.scala 37:46:@12479.4]
  wire [4:0] _T_64917; // @[Modules.scala 37:46:@12480.4]
  wire [4:0] _T_64918; // @[Modules.scala 37:46:@12481.4]
  wire [5:0] _T_64919; // @[Modules.scala 40:46:@12483.4]
  wire [4:0] _T_64920; // @[Modules.scala 40:46:@12484.4]
  wire [4:0] _T_64921; // @[Modules.scala 40:46:@12485.4]
  wire [5:0] _T_64925; // @[Modules.scala 37:46:@12491.4]
  wire [4:0] _T_64926; // @[Modules.scala 37:46:@12492.4]
  wire [4:0] _T_64927; // @[Modules.scala 37:46:@12493.4]
  wire [5:0] _T_64932; // @[Modules.scala 43:47:@12498.4]
  wire [4:0] _T_64933; // @[Modules.scala 43:47:@12499.4]
  wire [4:0] _T_64934; // @[Modules.scala 43:47:@12500.4]
  wire [5:0] _T_64977; // @[Modules.scala 43:47:@12544.4]
  wire [4:0] _T_64978; // @[Modules.scala 43:47:@12545.4]
  wire [4:0] _T_64979; // @[Modules.scala 43:47:@12546.4]
  wire [5:0] _T_64984; // @[Modules.scala 46:47:@12551.4]
  wire [4:0] _T_64985; // @[Modules.scala 46:47:@12552.4]
  wire [4:0] _T_64986; // @[Modules.scala 46:47:@12553.4]
  wire [5:0] _T_64987; // @[Modules.scala 37:46:@12555.4]
  wire [4:0] _T_64988; // @[Modules.scala 37:46:@12556.4]
  wire [4:0] _T_64989; // @[Modules.scala 37:46:@12557.4]
  wire [5:0] _T_64990; // @[Modules.scala 37:46:@12559.4]
  wire [4:0] _T_64991; // @[Modules.scala 37:46:@12560.4]
  wire [4:0] _T_64992; // @[Modules.scala 37:46:@12561.4]
  wire [5:0] _T_64993; // @[Modules.scala 40:46:@12563.4]
  wire [4:0] _T_64994; // @[Modules.scala 40:46:@12564.4]
  wire [4:0] _T_64995; // @[Modules.scala 40:46:@12565.4]
  wire [5:0] _T_64999; // @[Modules.scala 37:46:@12571.4]
  wire [4:0] _T_65000; // @[Modules.scala 37:46:@12572.4]
  wire [4:0] _T_65001; // @[Modules.scala 37:46:@12573.4]
  wire [5:0] _T_65009; // @[Modules.scala 46:47:@12582.4]
  wire [4:0] _T_65010; // @[Modules.scala 46:47:@12583.4]
  wire [4:0] _T_65011; // @[Modules.scala 46:47:@12584.4]
  wire [5:0] _T_65049; // @[Modules.scala 37:46:@12626.4]
  wire [4:0] _T_65050; // @[Modules.scala 37:46:@12627.4]
  wire [4:0] _T_65051; // @[Modules.scala 37:46:@12628.4]
  wire [5:0] _T_65052; // @[Modules.scala 37:46:@12630.4]
  wire [4:0] _T_65053; // @[Modules.scala 37:46:@12631.4]
  wire [4:0] _T_65054; // @[Modules.scala 37:46:@12632.4]
  wire [5:0] _T_65065; // @[Modules.scala 37:46:@12645.4]
  wire [4:0] _T_65066; // @[Modules.scala 37:46:@12646.4]
  wire [4:0] _T_65067; // @[Modules.scala 37:46:@12647.4]
  wire [5:0] _T_65068; // @[Modules.scala 40:46:@12649.4]
  wire [4:0] _T_65069; // @[Modules.scala 40:46:@12650.4]
  wire [4:0] _T_65070; // @[Modules.scala 40:46:@12651.4]
  wire [5:0] _T_65103; // @[Modules.scala 43:47:@12684.4]
  wire [4:0] _T_65104; // @[Modules.scala 43:47:@12685.4]
  wire [4:0] _T_65105; // @[Modules.scala 43:47:@12686.4]
  wire [5:0] _T_65115; // @[Modules.scala 37:46:@12700.4]
  wire [4:0] _T_65116; // @[Modules.scala 37:46:@12701.4]
  wire [4:0] _T_65117; // @[Modules.scala 37:46:@12702.4]
  wire [5:0] _T_65118; // @[Modules.scala 37:46:@12704.4]
  wire [4:0] _T_65119; // @[Modules.scala 37:46:@12705.4]
  wire [4:0] _T_65120; // @[Modules.scala 37:46:@12706.4]
  wire [5:0] _T_65121; // @[Modules.scala 40:46:@12708.4]
  wire [4:0] _T_65122; // @[Modules.scala 40:46:@12709.4]
  wire [4:0] _T_65123; // @[Modules.scala 40:46:@12710.4]
  wire [5:0] _T_65127; // @[Modules.scala 37:46:@12716.4]
  wire [4:0] _T_65128; // @[Modules.scala 37:46:@12717.4]
  wire [4:0] _T_65129; // @[Modules.scala 37:46:@12718.4]
  wire [5:0] _T_65141; // @[Modules.scala 46:37:@12731.4]
  wire [4:0] _T_65142; // @[Modules.scala 46:37:@12732.4]
  wire [4:0] _T_65143; // @[Modules.scala 46:37:@12733.4]
  wire [5:0] _T_65144; // @[Modules.scala 46:47:@12734.4]
  wire [4:0] _T_65145; // @[Modules.scala 46:47:@12735.4]
  wire [4:0] _T_65146; // @[Modules.scala 46:47:@12736.4]
  wire [5:0] _T_65180; // @[Modules.scala 37:46:@12775.4]
  wire [4:0] _T_65181; // @[Modules.scala 37:46:@12776.4]
  wire [4:0] _T_65182; // @[Modules.scala 37:46:@12777.4]
  wire [5:0] _T_65195; // @[Modules.scala 40:46:@12795.4]
  wire [4:0] _T_65196; // @[Modules.scala 40:46:@12796.4]
  wire [4:0] _T_65197; // @[Modules.scala 40:46:@12797.4]
  wire [5:0] _T_65202; // @[Modules.scala 46:47:@12802.4]
  wire [4:0] _T_65203; // @[Modules.scala 46:47:@12803.4]
  wire [4:0] _T_65204; // @[Modules.scala 46:47:@12804.4]
  wire [5:0] _T_65212; // @[Modules.scala 40:46:@12813.4]
  wire [4:0] _T_65213; // @[Modules.scala 40:46:@12814.4]
  wire [4:0] _T_65214; // @[Modules.scala 40:46:@12815.4]
  wire [5:0] _T_65226; // @[Modules.scala 46:47:@12827.4]
  wire [4:0] _T_65227; // @[Modules.scala 46:47:@12828.4]
  wire [4:0] _T_65228; // @[Modules.scala 46:47:@12829.4]
  wire [5:0] _T_65232; // @[Modules.scala 37:46:@12835.4]
  wire [4:0] _T_65233; // @[Modules.scala 37:46:@12836.4]
  wire [4:0] _T_65234; // @[Modules.scala 37:46:@12837.4]
  wire [5:0] _T_65235; // @[Modules.scala 37:46:@12839.4]
  wire [4:0] _T_65236; // @[Modules.scala 37:46:@12840.4]
  wire [4:0] _T_65237; // @[Modules.scala 37:46:@12841.4]
  wire [5:0] _T_65238; // @[Modules.scala 40:46:@12843.4]
  wire [4:0] _T_65239; // @[Modules.scala 40:46:@12844.4]
  wire [4:0] _T_65240; // @[Modules.scala 40:46:@12845.4]
  wire [5:0] _T_65250; // @[Modules.scala 37:46:@12859.4]
  wire [4:0] _T_65251; // @[Modules.scala 37:46:@12860.4]
  wire [4:0] _T_65252; // @[Modules.scala 37:46:@12861.4]
  wire [5:0] _T_65259; // @[Modules.scala 40:46:@12871.4]
  wire [4:0] _T_65260; // @[Modules.scala 40:46:@12872.4]
  wire [4:0] _T_65261; // @[Modules.scala 40:46:@12873.4]
  wire [5:0] _T_65278; // @[Modules.scala 37:46:@12894.4]
  wire [4:0] _T_65279; // @[Modules.scala 37:46:@12895.4]
  wire [4:0] _T_65280; // @[Modules.scala 37:46:@12896.4]
  wire [5:0] _T_65284; // @[Modules.scala 37:46:@12902.4]
  wire [4:0] _T_65285; // @[Modules.scala 37:46:@12903.4]
  wire [4:0] _T_65286; // @[Modules.scala 37:46:@12904.4]
  wire [5:0] _T_65300; // @[Modules.scala 37:46:@12921.4]
  wire [4:0] _T_65301; // @[Modules.scala 37:46:@12922.4]
  wire [4:0] _T_65302; // @[Modules.scala 37:46:@12923.4]
  wire [5:0] _T_65321; // @[Modules.scala 46:37:@12943.4]
  wire [4:0] _T_65322; // @[Modules.scala 46:37:@12944.4]
  wire [4:0] _T_65323; // @[Modules.scala 46:37:@12945.4]
  wire [5:0] _T_65324; // @[Modules.scala 46:47:@12946.4]
  wire [4:0] _T_65325; // @[Modules.scala 46:47:@12947.4]
  wire [4:0] _T_65326; // @[Modules.scala 46:47:@12948.4]
  wire [5:0] _T_65341; // @[Modules.scala 43:47:@12964.4]
  wire [4:0] _T_65342; // @[Modules.scala 43:47:@12965.4]
  wire [4:0] _T_65343; // @[Modules.scala 43:47:@12966.4]
  wire [5:0] _T_65344; // @[Modules.scala 37:46:@12968.4]
  wire [4:0] _T_65345; // @[Modules.scala 37:46:@12969.4]
  wire [4:0] _T_65346; // @[Modules.scala 37:46:@12970.4]
  wire [5:0] _T_65350; // @[Modules.scala 40:46:@12976.4]
  wire [4:0] _T_65351; // @[Modules.scala 40:46:@12977.4]
  wire [4:0] _T_65352; // @[Modules.scala 40:46:@12978.4]
  wire [5:0] _T_65363; // @[Modules.scala 37:46:@12991.4]
  wire [4:0] _T_65364; // @[Modules.scala 37:46:@12992.4]
  wire [4:0] _T_65365; // @[Modules.scala 37:46:@12993.4]
  wire [5:0] _T_65380; // @[Modules.scala 43:47:@13009.4]
  wire [4:0] _T_65381; // @[Modules.scala 43:47:@13010.4]
  wire [4:0] _T_65382; // @[Modules.scala 43:47:@13011.4]
  wire [5:0] _T_65386; // @[Modules.scala 40:46:@13017.4]
  wire [4:0] _T_65387; // @[Modules.scala 40:46:@13018.4]
  wire [4:0] _T_65388; // @[Modules.scala 40:46:@13019.4]
  wire [5:0] _T_65389; // @[Modules.scala 40:46:@13021.4]
  wire [4:0] _T_65390; // @[Modules.scala 40:46:@13022.4]
  wire [4:0] _T_65391; // @[Modules.scala 40:46:@13023.4]
  wire [5:0] _T_65396; // @[Modules.scala 43:47:@13028.4]
  wire [4:0] _T_65397; // @[Modules.scala 43:47:@13029.4]
  wire [4:0] _T_65398; // @[Modules.scala 43:47:@13030.4]
  wire [5:0] _T_65402; // @[Modules.scala 37:46:@13036.4]
  wire [4:0] _T_65403; // @[Modules.scala 37:46:@13037.4]
  wire [4:0] _T_65404; // @[Modules.scala 37:46:@13038.4]
  wire [5:0] _T_65408; // @[Modules.scala 40:46:@13044.4]
  wire [4:0] _T_65409; // @[Modules.scala 40:46:@13045.4]
  wire [4:0] _T_65410; // @[Modules.scala 40:46:@13046.4]
  wire [5:0] _T_65424; // @[Modules.scala 43:47:@13063.4]
  wire [4:0] _T_65425; // @[Modules.scala 43:47:@13064.4]
  wire [4:0] _T_65426; // @[Modules.scala 43:47:@13065.4]
  wire [5:0] _T_65431; // @[Modules.scala 43:47:@13070.4]
  wire [4:0] _T_65432; // @[Modules.scala 43:47:@13071.4]
  wire [4:0] _T_65433; // @[Modules.scala 43:47:@13072.4]
  wire [5:0] _T_65458; // @[Modules.scala 46:47:@13099.4]
  wire [4:0] _T_65459; // @[Modules.scala 46:47:@13100.4]
  wire [4:0] _T_65460; // @[Modules.scala 46:47:@13101.4]
  wire [5:0] _T_65468; // @[Modules.scala 40:46:@13110.4]
  wire [4:0] _T_65469; // @[Modules.scala 40:46:@13111.4]
  wire [4:0] _T_65470; // @[Modules.scala 40:46:@13112.4]
  wire [5:0] _T_65474; // @[Modules.scala 40:46:@13118.4]
  wire [4:0] _T_65475; // @[Modules.scala 40:46:@13119.4]
  wire [4:0] _T_65476; // @[Modules.scala 40:46:@13120.4]
  wire [5:0] _T_65477; // @[Modules.scala 40:46:@13122.4]
  wire [4:0] _T_65478; // @[Modules.scala 40:46:@13123.4]
  wire [4:0] _T_65479; // @[Modules.scala 40:46:@13124.4]
  wire [5:0] _T_65481; // @[Modules.scala 43:37:@13126.4]
  wire [4:0] _T_65482; // @[Modules.scala 43:37:@13127.4]
  wire [4:0] _T_65483; // @[Modules.scala 43:37:@13128.4]
  wire [5:0] _T_65484; // @[Modules.scala 43:47:@13129.4]
  wire [4:0] _T_65485; // @[Modules.scala 43:47:@13130.4]
  wire [4:0] _T_65486; // @[Modules.scala 43:47:@13131.4]
  wire [5:0] _T_65503; // @[Modules.scala 43:47:@13152.4]
  wire [4:0] _T_65504; // @[Modules.scala 43:47:@13153.4]
  wire [4:0] _T_65505; // @[Modules.scala 43:47:@13154.4]
  wire [5:0] _T_65506; // @[Modules.scala 37:46:@13156.4]
  wire [4:0] _T_65507; // @[Modules.scala 37:46:@13157.4]
  wire [4:0] _T_65508; // @[Modules.scala 37:46:@13158.4]
  wire [5:0] _T_65513; // @[Modules.scala 46:47:@13163.4]
  wire [4:0] _T_65514; // @[Modules.scala 46:47:@13164.4]
  wire [4:0] _T_65515; // @[Modules.scala 46:47:@13165.4]
  wire [5:0] _T_65517; // @[Modules.scala 46:37:@13167.4]
  wire [4:0] _T_65518; // @[Modules.scala 46:37:@13168.4]
  wire [4:0] _T_65519; // @[Modules.scala 46:37:@13169.4]
  wire [5:0] _T_65520; // @[Modules.scala 46:47:@13170.4]
  wire [4:0] _T_65521; // @[Modules.scala 46:47:@13171.4]
  wire [4:0] _T_65522; // @[Modules.scala 46:47:@13172.4]
  wire [5:0] _T_65534; // @[Modules.scala 46:47:@13184.4]
  wire [4:0] _T_65535; // @[Modules.scala 46:47:@13185.4]
  wire [4:0] _T_65536; // @[Modules.scala 46:47:@13186.4]
  wire [5:0] _T_65544; // @[Modules.scala 37:46:@13195.4]
  wire [4:0] _T_65545; // @[Modules.scala 37:46:@13196.4]
  wire [4:0] _T_65546; // @[Modules.scala 37:46:@13197.4]
  wire [5:0] _T_65555; // @[Modules.scala 43:37:@13206.4]
  wire [4:0] _T_65556; // @[Modules.scala 43:37:@13207.4]
  wire [4:0] _T_65557; // @[Modules.scala 43:37:@13208.4]
  wire [5:0] _T_65558; // @[Modules.scala 43:47:@13209.4]
  wire [4:0] _T_65559; // @[Modules.scala 43:47:@13210.4]
  wire [4:0] _T_65560; // @[Modules.scala 43:47:@13211.4]
  wire [5:0] _T_65570; // @[Modules.scala 37:46:@13225.4]
  wire [4:0] _T_65571; // @[Modules.scala 37:46:@13226.4]
  wire [4:0] _T_65572; // @[Modules.scala 37:46:@13227.4]
  wire [5:0] _T_65597; // @[Modules.scala 46:37:@13255.4]
  wire [4:0] _T_65598; // @[Modules.scala 46:37:@13256.4]
  wire [4:0] _T_65599; // @[Modules.scala 46:37:@13257.4]
  wire [5:0] _T_65600; // @[Modules.scala 46:47:@13258.4]
  wire [4:0] _T_65601; // @[Modules.scala 46:47:@13259.4]
  wire [4:0] _T_65602; // @[Modules.scala 46:47:@13260.4]
  wire [5:0] _T_65612; // @[Modules.scala 40:46:@13274.4]
  wire [4:0] _T_65613; // @[Modules.scala 40:46:@13275.4]
  wire [4:0] _T_65614; // @[Modules.scala 40:46:@13276.4]
  wire [5:0] _T_65621; // @[Modules.scala 37:46:@13286.4]
  wire [4:0] _T_65622; // @[Modules.scala 37:46:@13287.4]
  wire [4:0] _T_65623; // @[Modules.scala 37:46:@13288.4]
  wire [5:0] _T_65624; // @[Modules.scala 37:46:@13290.4]
  wire [4:0] _T_65625; // @[Modules.scala 37:46:@13291.4]
  wire [4:0] _T_65626; // @[Modules.scala 37:46:@13292.4]
  wire [5:0] _T_65627; // @[Modules.scala 37:46:@13294.4]
  wire [4:0] _T_65628; // @[Modules.scala 37:46:@13295.4]
  wire [4:0] _T_65629; // @[Modules.scala 37:46:@13296.4]
  wire [5:0] _T_65634; // @[Modules.scala 43:47:@13301.4]
  wire [4:0] _T_65635; // @[Modules.scala 43:47:@13302.4]
  wire [4:0] _T_65636; // @[Modules.scala 43:47:@13303.4]
  wire [5:0] _T_65637; // @[Modules.scala 37:46:@13305.4]
  wire [4:0] _T_65638; // @[Modules.scala 37:46:@13306.4]
  wire [4:0] _T_65639; // @[Modules.scala 37:46:@13307.4]
  wire [5:0] _T_65640; // @[Modules.scala 37:46:@13309.4]
  wire [4:0] _T_65641; // @[Modules.scala 37:46:@13310.4]
  wire [4:0] _T_65642; // @[Modules.scala 37:46:@13311.4]
  wire [5:0] _T_65644; // @[Modules.scala 46:37:@13313.4]
  wire [4:0] _T_65645; // @[Modules.scala 46:37:@13314.4]
  wire [4:0] _T_65646; // @[Modules.scala 46:37:@13315.4]
  wire [5:0] _T_65647; // @[Modules.scala 46:47:@13316.4]
  wire [4:0] _T_65648; // @[Modules.scala 46:47:@13317.4]
  wire [4:0] _T_65649; // @[Modules.scala 46:47:@13318.4]
  wire [5:0] _T_65653; // @[Modules.scala 40:46:@13324.4]
  wire [4:0] _T_65654; // @[Modules.scala 40:46:@13325.4]
  wire [4:0] _T_65655; // @[Modules.scala 40:46:@13326.4]
  wire [5:0] _T_65657; // @[Modules.scala 43:37:@13328.4]
  wire [4:0] _T_65658; // @[Modules.scala 43:37:@13329.4]
  wire [4:0] _T_65659; // @[Modules.scala 43:37:@13330.4]
  wire [5:0] _T_65660; // @[Modules.scala 43:47:@13331.4]
  wire [4:0] _T_65661; // @[Modules.scala 43:47:@13332.4]
  wire [4:0] _T_65662; // @[Modules.scala 43:47:@13333.4]
  wire [5:0] _T_65663; // @[Modules.scala 37:46:@13335.4]
  wire [4:0] _T_65664; // @[Modules.scala 37:46:@13336.4]
  wire [4:0] _T_65665; // @[Modules.scala 37:46:@13337.4]
  wire [5:0] _T_65679; // @[Modules.scala 37:46:@13354.4]
  wire [4:0] _T_65680; // @[Modules.scala 37:46:@13355.4]
  wire [4:0] _T_65681; // @[Modules.scala 37:46:@13356.4]
  wire [5:0] _T_65685; // @[Modules.scala 37:46:@13362.4]
  wire [4:0] _T_65686; // @[Modules.scala 37:46:@13363.4]
  wire [4:0] _T_65687; // @[Modules.scala 37:46:@13364.4]
  wire [5:0] _T_65688; // @[Modules.scala 37:46:@13366.4]
  wire [4:0] _T_65689; // @[Modules.scala 37:46:@13367.4]
  wire [4:0] _T_65690; // @[Modules.scala 37:46:@13368.4]
  wire [5:0] _T_65691; // @[Modules.scala 37:46:@13370.4]
  wire [4:0] _T_65692; // @[Modules.scala 37:46:@13371.4]
  wire [4:0] _T_65693; // @[Modules.scala 37:46:@13372.4]
  wire [5:0] _T_65694; // @[Modules.scala 37:46:@13374.4]
  wire [4:0] _T_65695; // @[Modules.scala 37:46:@13375.4]
  wire [4:0] _T_65696; // @[Modules.scala 37:46:@13376.4]
  wire [5:0] _T_65708; // @[Modules.scala 43:47:@13388.4]
  wire [4:0] _T_65709; // @[Modules.scala 43:47:@13389.4]
  wire [4:0] _T_65710; // @[Modules.scala 43:47:@13390.4]
  wire [10:0] buffer_3_0; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65717; // @[Modules.scala 50:57:@13400.4]
  wire [10:0] _T_65718; // @[Modules.scala 50:57:@13401.4]
  wire [10:0] buffer_3_392; // @[Modules.scala 50:57:@13402.4]
  wire [10:0] buffer_3_4; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65723; // @[Modules.scala 50:57:@13408.4]
  wire [10:0] _T_65724; // @[Modules.scala 50:57:@13409.4]
  wire [10:0] buffer_3_394; // @[Modules.scala 50:57:@13410.4]
  wire [11:0] _T_65729; // @[Modules.scala 50:57:@13416.4]
  wire [10:0] _T_65730; // @[Modules.scala 50:57:@13417.4]
  wire [10:0] buffer_3_396; // @[Modules.scala 50:57:@13418.4]
  wire [11:0] _T_65732; // @[Modules.scala 50:57:@13420.4]
  wire [10:0] _T_65733; // @[Modules.scala 50:57:@13421.4]
  wire [10:0] buffer_3_397; // @[Modules.scala 50:57:@13422.4]
  wire [10:0] buffer_3_12; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65735; // @[Modules.scala 50:57:@13424.4]
  wire [10:0] _T_65736; // @[Modules.scala 50:57:@13425.4]
  wire [10:0] buffer_3_398; // @[Modules.scala 50:57:@13426.4]
  wire [10:0] buffer_3_14; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65738; // @[Modules.scala 50:57:@13428.4]
  wire [10:0] _T_65739; // @[Modules.scala 50:57:@13429.4]
  wire [10:0] buffer_3_399; // @[Modules.scala 50:57:@13430.4]
  wire [10:0] buffer_3_16; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65741; // @[Modules.scala 50:57:@13432.4]
  wire [10:0] _T_65742; // @[Modules.scala 50:57:@13433.4]
  wire [10:0] buffer_3_400; // @[Modules.scala 50:57:@13434.4]
  wire [11:0] _T_65750; // @[Modules.scala 50:57:@13444.4]
  wire [10:0] _T_65751; // @[Modules.scala 50:57:@13445.4]
  wire [10:0] buffer_3_403; // @[Modules.scala 50:57:@13446.4]
  wire [11:0] _T_65753; // @[Modules.scala 50:57:@13448.4]
  wire [10:0] _T_65754; // @[Modules.scala 50:57:@13449.4]
  wire [10:0] buffer_3_404; // @[Modules.scala 50:57:@13450.4]
  wire [10:0] buffer_3_26; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65756; // @[Modules.scala 50:57:@13452.4]
  wire [10:0] _T_65757; // @[Modules.scala 50:57:@13453.4]
  wire [10:0] buffer_3_405; // @[Modules.scala 50:57:@13454.4]
  wire [10:0] buffer_3_28; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65759; // @[Modules.scala 50:57:@13456.4]
  wire [10:0] _T_65760; // @[Modules.scala 50:57:@13457.4]
  wire [10:0] buffer_3_406; // @[Modules.scala 50:57:@13458.4]
  wire [10:0] buffer_3_30; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65762; // @[Modules.scala 50:57:@13460.4]
  wire [10:0] _T_65763; // @[Modules.scala 50:57:@13461.4]
  wire [10:0] buffer_3_407; // @[Modules.scala 50:57:@13462.4]
  wire [10:0] buffer_3_32; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65765; // @[Modules.scala 50:57:@13464.4]
  wire [10:0] _T_65766; // @[Modules.scala 50:57:@13465.4]
  wire [10:0] buffer_3_408; // @[Modules.scala 50:57:@13466.4]
  wire [10:0] buffer_3_37; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65771; // @[Modules.scala 50:57:@13472.4]
  wire [10:0] _T_65772; // @[Modules.scala 50:57:@13473.4]
  wire [10:0] buffer_3_410; // @[Modules.scala 50:57:@13474.4]
  wire [10:0] buffer_3_38; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_39; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65774; // @[Modules.scala 50:57:@13476.4]
  wire [10:0] _T_65775; // @[Modules.scala 50:57:@13477.4]
  wire [10:0] buffer_3_411; // @[Modules.scala 50:57:@13478.4]
  wire [11:0] _T_65777; // @[Modules.scala 50:57:@13480.4]
  wire [10:0] _T_65778; // @[Modules.scala 50:57:@13481.4]
  wire [10:0] buffer_3_412; // @[Modules.scala 50:57:@13482.4]
  wire [10:0] buffer_3_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65780; // @[Modules.scala 50:57:@13484.4]
  wire [10:0] _T_65781; // @[Modules.scala 50:57:@13485.4]
  wire [10:0] buffer_3_413; // @[Modules.scala 50:57:@13486.4]
  wire [10:0] buffer_3_44; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_45; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65783; // @[Modules.scala 50:57:@13488.4]
  wire [10:0] _T_65784; // @[Modules.scala 50:57:@13489.4]
  wire [10:0] buffer_3_414; // @[Modules.scala 50:57:@13490.4]
  wire [10:0] buffer_3_46; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65786; // @[Modules.scala 50:57:@13492.4]
  wire [10:0] _T_65787; // @[Modules.scala 50:57:@13493.4]
  wire [10:0] buffer_3_415; // @[Modules.scala 50:57:@13494.4]
  wire [10:0] buffer_3_49; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65789; // @[Modules.scala 50:57:@13496.4]
  wire [10:0] _T_65790; // @[Modules.scala 50:57:@13497.4]
  wire [10:0] buffer_3_416; // @[Modules.scala 50:57:@13498.4]
  wire [10:0] buffer_3_51; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65792; // @[Modules.scala 50:57:@13500.4]
  wire [10:0] _T_65793; // @[Modules.scala 50:57:@13501.4]
  wire [10:0] buffer_3_417; // @[Modules.scala 50:57:@13502.4]
  wire [10:0] buffer_3_52; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_53; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65795; // @[Modules.scala 50:57:@13504.4]
  wire [10:0] _T_65796; // @[Modules.scala 50:57:@13505.4]
  wire [10:0] buffer_3_418; // @[Modules.scala 50:57:@13506.4]
  wire [10:0] buffer_3_54; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65798; // @[Modules.scala 50:57:@13508.4]
  wire [10:0] _T_65799; // @[Modules.scala 50:57:@13509.4]
  wire [10:0] buffer_3_419; // @[Modules.scala 50:57:@13510.4]
  wire [10:0] buffer_3_56; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65801; // @[Modules.scala 50:57:@13512.4]
  wire [10:0] _T_65802; // @[Modules.scala 50:57:@13513.4]
  wire [10:0] buffer_3_420; // @[Modules.scala 50:57:@13514.4]
  wire [11:0] _T_65804; // @[Modules.scala 50:57:@13516.4]
  wire [10:0] _T_65805; // @[Modules.scala 50:57:@13517.4]
  wire [10:0] buffer_3_421; // @[Modules.scala 50:57:@13518.4]
  wire [10:0] buffer_3_60; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65807; // @[Modules.scala 50:57:@13520.4]
  wire [10:0] _T_65808; // @[Modules.scala 50:57:@13521.4]
  wire [10:0] buffer_3_422; // @[Modules.scala 50:57:@13522.4]
  wire [10:0] buffer_3_62; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65810; // @[Modules.scala 50:57:@13524.4]
  wire [10:0] _T_65811; // @[Modules.scala 50:57:@13525.4]
  wire [10:0] buffer_3_423; // @[Modules.scala 50:57:@13526.4]
  wire [10:0] buffer_3_66; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_67; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65816; // @[Modules.scala 50:57:@13532.4]
  wire [10:0] _T_65817; // @[Modules.scala 50:57:@13533.4]
  wire [10:0] buffer_3_425; // @[Modules.scala 50:57:@13534.4]
  wire [10:0] buffer_3_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65819; // @[Modules.scala 50:57:@13536.4]
  wire [10:0] _T_65820; // @[Modules.scala 50:57:@13537.4]
  wire [10:0] buffer_3_426; // @[Modules.scala 50:57:@13538.4]
  wire [11:0] _T_65822; // @[Modules.scala 50:57:@13540.4]
  wire [10:0] _T_65823; // @[Modules.scala 50:57:@13541.4]
  wire [10:0] buffer_3_427; // @[Modules.scala 50:57:@13542.4]
  wire [10:0] buffer_3_72; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65825; // @[Modules.scala 50:57:@13544.4]
  wire [10:0] _T_65826; // @[Modules.scala 50:57:@13545.4]
  wire [10:0] buffer_3_428; // @[Modules.scala 50:57:@13546.4]
  wire [10:0] buffer_3_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65828; // @[Modules.scala 50:57:@13548.4]
  wire [10:0] _T_65829; // @[Modules.scala 50:57:@13549.4]
  wire [10:0] buffer_3_429; // @[Modules.scala 50:57:@13550.4]
  wire [10:0] buffer_3_76; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_77; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65831; // @[Modules.scala 50:57:@13552.4]
  wire [10:0] _T_65832; // @[Modules.scala 50:57:@13553.4]
  wire [10:0] buffer_3_430; // @[Modules.scala 50:57:@13554.4]
  wire [10:0] buffer_3_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65834; // @[Modules.scala 50:57:@13556.4]
  wire [10:0] _T_65835; // @[Modules.scala 50:57:@13557.4]
  wire [10:0] buffer_3_431; // @[Modules.scala 50:57:@13558.4]
  wire [10:0] buffer_3_86; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65846; // @[Modules.scala 50:57:@13572.4]
  wire [10:0] _T_65847; // @[Modules.scala 50:57:@13573.4]
  wire [10:0] buffer_3_435; // @[Modules.scala 50:57:@13574.4]
  wire [10:0] buffer_3_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65849; // @[Modules.scala 50:57:@13576.4]
  wire [10:0] _T_65850; // @[Modules.scala 50:57:@13577.4]
  wire [10:0] buffer_3_436; // @[Modules.scala 50:57:@13578.4]
  wire [10:0] buffer_3_90; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65852; // @[Modules.scala 50:57:@13580.4]
  wire [10:0] _T_65853; // @[Modules.scala 50:57:@13581.4]
  wire [10:0] buffer_3_437; // @[Modules.scala 50:57:@13582.4]
  wire [10:0] buffer_3_92; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65855; // @[Modules.scala 50:57:@13584.4]
  wire [10:0] _T_65856; // @[Modules.scala 50:57:@13585.4]
  wire [10:0] buffer_3_438; // @[Modules.scala 50:57:@13586.4]
  wire [11:0] _T_65858; // @[Modules.scala 50:57:@13588.4]
  wire [10:0] _T_65859; // @[Modules.scala 50:57:@13589.4]
  wire [10:0] buffer_3_439; // @[Modules.scala 50:57:@13590.4]
  wire [10:0] buffer_3_98; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65864; // @[Modules.scala 50:57:@13596.4]
  wire [10:0] _T_65865; // @[Modules.scala 50:57:@13597.4]
  wire [10:0] buffer_3_441; // @[Modules.scala 50:57:@13598.4]
  wire [10:0] buffer_3_100; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65867; // @[Modules.scala 50:57:@13600.4]
  wire [10:0] _T_65868; // @[Modules.scala 50:57:@13601.4]
  wire [10:0] buffer_3_442; // @[Modules.scala 50:57:@13602.4]
  wire [10:0] buffer_3_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65870; // @[Modules.scala 50:57:@13604.4]
  wire [10:0] _T_65871; // @[Modules.scala 50:57:@13605.4]
  wire [10:0] buffer_3_443; // @[Modules.scala 50:57:@13606.4]
  wire [10:0] buffer_3_104; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65873; // @[Modules.scala 50:57:@13608.4]
  wire [10:0] _T_65874; // @[Modules.scala 50:57:@13609.4]
  wire [10:0] buffer_3_444; // @[Modules.scala 50:57:@13610.4]
  wire [10:0] buffer_3_106; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65876; // @[Modules.scala 50:57:@13612.4]
  wire [10:0] _T_65877; // @[Modules.scala 50:57:@13613.4]
  wire [10:0] buffer_3_445; // @[Modules.scala 50:57:@13614.4]
  wire [10:0] buffer_3_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65879; // @[Modules.scala 50:57:@13616.4]
  wire [10:0] _T_65880; // @[Modules.scala 50:57:@13617.4]
  wire [10:0] buffer_3_446; // @[Modules.scala 50:57:@13618.4]
  wire [10:0] buffer_3_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65885; // @[Modules.scala 50:57:@13624.4]
  wire [10:0] _T_65886; // @[Modules.scala 50:57:@13625.4]
  wire [10:0] buffer_3_448; // @[Modules.scala 50:57:@13626.4]
  wire [10:0] buffer_3_114; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65888; // @[Modules.scala 50:57:@13628.4]
  wire [10:0] _T_65889; // @[Modules.scala 50:57:@13629.4]
  wire [10:0] buffer_3_449; // @[Modules.scala 50:57:@13630.4]
  wire [10:0] buffer_3_116; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65891; // @[Modules.scala 50:57:@13632.4]
  wire [10:0] _T_65892; // @[Modules.scala 50:57:@13633.4]
  wire [10:0] buffer_3_450; // @[Modules.scala 50:57:@13634.4]
  wire [10:0] buffer_3_118; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65894; // @[Modules.scala 50:57:@13636.4]
  wire [10:0] _T_65895; // @[Modules.scala 50:57:@13637.4]
  wire [10:0] buffer_3_451; // @[Modules.scala 50:57:@13638.4]
  wire [10:0] buffer_3_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65897; // @[Modules.scala 50:57:@13640.4]
  wire [10:0] _T_65898; // @[Modules.scala 50:57:@13641.4]
  wire [10:0] buffer_3_452; // @[Modules.scala 50:57:@13642.4]
  wire [10:0] buffer_3_122; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65900; // @[Modules.scala 50:57:@13644.4]
  wire [10:0] _T_65901; // @[Modules.scala 50:57:@13645.4]
  wire [10:0] buffer_3_453; // @[Modules.scala 50:57:@13646.4]
  wire [10:0] buffer_3_126; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_127; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65906; // @[Modules.scala 50:57:@13652.4]
  wire [10:0] _T_65907; // @[Modules.scala 50:57:@13653.4]
  wire [10:0] buffer_3_455; // @[Modules.scala 50:57:@13654.4]
  wire [10:0] buffer_3_128; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65909; // @[Modules.scala 50:57:@13656.4]
  wire [10:0] _T_65910; // @[Modules.scala 50:57:@13657.4]
  wire [10:0] buffer_3_456; // @[Modules.scala 50:57:@13658.4]
  wire [10:0] buffer_3_132; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65915; // @[Modules.scala 50:57:@13664.4]
  wire [10:0] _T_65916; // @[Modules.scala 50:57:@13665.4]
  wire [10:0] buffer_3_458; // @[Modules.scala 50:57:@13666.4]
  wire [10:0] buffer_3_134; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65918; // @[Modules.scala 50:57:@13668.4]
  wire [10:0] _T_65919; // @[Modules.scala 50:57:@13669.4]
  wire [10:0] buffer_3_459; // @[Modules.scala 50:57:@13670.4]
  wire [10:0] buffer_3_136; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65921; // @[Modules.scala 50:57:@13672.4]
  wire [10:0] _T_65922; // @[Modules.scala 50:57:@13673.4]
  wire [10:0] buffer_3_460; // @[Modules.scala 50:57:@13674.4]
  wire [10:0] buffer_3_140; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65927; // @[Modules.scala 50:57:@13680.4]
  wire [10:0] _T_65928; // @[Modules.scala 50:57:@13681.4]
  wire [10:0] buffer_3_462; // @[Modules.scala 50:57:@13682.4]
  wire [10:0] buffer_3_142; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65930; // @[Modules.scala 50:57:@13684.4]
  wire [10:0] _T_65931; // @[Modules.scala 50:57:@13685.4]
  wire [10:0] buffer_3_463; // @[Modules.scala 50:57:@13686.4]
  wire [10:0] buffer_3_144; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65933; // @[Modules.scala 50:57:@13688.4]
  wire [10:0] _T_65934; // @[Modules.scala 50:57:@13689.4]
  wire [10:0] buffer_3_464; // @[Modules.scala 50:57:@13690.4]
  wire [10:0] buffer_3_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65936; // @[Modules.scala 50:57:@13692.4]
  wire [10:0] _T_65937; // @[Modules.scala 50:57:@13693.4]
  wire [10:0] buffer_3_465; // @[Modules.scala 50:57:@13694.4]
  wire [10:0] buffer_3_148; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_149; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65939; // @[Modules.scala 50:57:@13696.4]
  wire [10:0] _T_65940; // @[Modules.scala 50:57:@13697.4]
  wire [10:0] buffer_3_466; // @[Modules.scala 50:57:@13698.4]
  wire [10:0] buffer_3_150; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65942; // @[Modules.scala 50:57:@13700.4]
  wire [10:0] _T_65943; // @[Modules.scala 50:57:@13701.4]
  wire [10:0] buffer_3_467; // @[Modules.scala 50:57:@13702.4]
  wire [10:0] buffer_3_154; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65948; // @[Modules.scala 50:57:@13708.4]
  wire [10:0] _T_65949; // @[Modules.scala 50:57:@13709.4]
  wire [10:0] buffer_3_469; // @[Modules.scala 50:57:@13710.4]
  wire [10:0] buffer_3_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65951; // @[Modules.scala 50:57:@13712.4]
  wire [10:0] _T_65952; // @[Modules.scala 50:57:@13713.4]
  wire [10:0] buffer_3_470; // @[Modules.scala 50:57:@13714.4]
  wire [10:0] buffer_3_159; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65954; // @[Modules.scala 50:57:@13716.4]
  wire [10:0] _T_65955; // @[Modules.scala 50:57:@13717.4]
  wire [10:0] buffer_3_471; // @[Modules.scala 50:57:@13718.4]
  wire [10:0] buffer_3_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65966; // @[Modules.scala 50:57:@13732.4]
  wire [10:0] _T_65967; // @[Modules.scala 50:57:@13733.4]
  wire [10:0] buffer_3_475; // @[Modules.scala 50:57:@13734.4]
  wire [10:0] buffer_3_168; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65969; // @[Modules.scala 50:57:@13736.4]
  wire [10:0] _T_65970; // @[Modules.scala 50:57:@13737.4]
  wire [10:0] buffer_3_476; // @[Modules.scala 50:57:@13738.4]
  wire [10:0] buffer_3_170; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65972; // @[Modules.scala 50:57:@13740.4]
  wire [10:0] _T_65973; // @[Modules.scala 50:57:@13741.4]
  wire [10:0] buffer_3_477; // @[Modules.scala 50:57:@13742.4]
  wire [10:0] buffer_3_172; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65975; // @[Modules.scala 50:57:@13744.4]
  wire [10:0] _T_65976; // @[Modules.scala 50:57:@13745.4]
  wire [10:0] buffer_3_478; // @[Modules.scala 50:57:@13746.4]
  wire [10:0] buffer_3_174; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65978; // @[Modules.scala 50:57:@13748.4]
  wire [10:0] _T_65979; // @[Modules.scala 50:57:@13749.4]
  wire [10:0] buffer_3_479; // @[Modules.scala 50:57:@13750.4]
  wire [11:0] _T_65987; // @[Modules.scala 50:57:@13760.4]
  wire [10:0] _T_65988; // @[Modules.scala 50:57:@13761.4]
  wire [10:0] buffer_3_482; // @[Modules.scala 50:57:@13762.4]
  wire [10:0] buffer_3_182; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65990; // @[Modules.scala 50:57:@13764.4]
  wire [10:0] _T_65991; // @[Modules.scala 50:57:@13765.4]
  wire [10:0] buffer_3_483; // @[Modules.scala 50:57:@13766.4]
  wire [10:0] buffer_3_184; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65993; // @[Modules.scala 50:57:@13768.4]
  wire [10:0] _T_65994; // @[Modules.scala 50:57:@13769.4]
  wire [10:0] buffer_3_484; // @[Modules.scala 50:57:@13770.4]
  wire [10:0] buffer_3_186; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_187; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65996; // @[Modules.scala 50:57:@13772.4]
  wire [10:0] _T_65997; // @[Modules.scala 50:57:@13773.4]
  wire [10:0] buffer_3_485; // @[Modules.scala 50:57:@13774.4]
  wire [10:0] buffer_3_188; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65999; // @[Modules.scala 50:57:@13776.4]
  wire [10:0] _T_66000; // @[Modules.scala 50:57:@13777.4]
  wire [10:0] buffer_3_486; // @[Modules.scala 50:57:@13778.4]
  wire [10:0] buffer_3_190; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66002; // @[Modules.scala 50:57:@13780.4]
  wire [10:0] _T_66003; // @[Modules.scala 50:57:@13781.4]
  wire [10:0] buffer_3_487; // @[Modules.scala 50:57:@13782.4]
  wire [10:0] buffer_3_192; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66005; // @[Modules.scala 50:57:@13784.4]
  wire [10:0] _T_66006; // @[Modules.scala 50:57:@13785.4]
  wire [10:0] buffer_3_488; // @[Modules.scala 50:57:@13786.4]
  wire [10:0] buffer_3_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66008; // @[Modules.scala 50:57:@13788.4]
  wire [10:0] _T_66009; // @[Modules.scala 50:57:@13789.4]
  wire [10:0] buffer_3_489; // @[Modules.scala 50:57:@13790.4]
  wire [10:0] buffer_3_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66011; // @[Modules.scala 50:57:@13792.4]
  wire [10:0] _T_66012; // @[Modules.scala 50:57:@13793.4]
  wire [10:0] buffer_3_490; // @[Modules.scala 50:57:@13794.4]
  wire [10:0] buffer_3_198; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66014; // @[Modules.scala 50:57:@13796.4]
  wire [10:0] _T_66015; // @[Modules.scala 50:57:@13797.4]
  wire [10:0] buffer_3_491; // @[Modules.scala 50:57:@13798.4]
  wire [10:0] buffer_3_200; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_201; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66017; // @[Modules.scala 50:57:@13800.4]
  wire [10:0] _T_66018; // @[Modules.scala 50:57:@13801.4]
  wire [10:0] buffer_3_492; // @[Modules.scala 50:57:@13802.4]
  wire [10:0] buffer_3_202; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66020; // @[Modules.scala 50:57:@13804.4]
  wire [10:0] _T_66021; // @[Modules.scala 50:57:@13805.4]
  wire [10:0] buffer_3_493; // @[Modules.scala 50:57:@13806.4]
  wire [10:0] buffer_3_204; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66023; // @[Modules.scala 50:57:@13808.4]
  wire [10:0] _T_66024; // @[Modules.scala 50:57:@13809.4]
  wire [10:0] buffer_3_494; // @[Modules.scala 50:57:@13810.4]
  wire [10:0] buffer_3_206; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_207; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66026; // @[Modules.scala 50:57:@13812.4]
  wire [10:0] _T_66027; // @[Modules.scala 50:57:@13813.4]
  wire [10:0] buffer_3_495; // @[Modules.scala 50:57:@13814.4]
  wire [10:0] buffer_3_208; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66029; // @[Modules.scala 50:57:@13816.4]
  wire [10:0] _T_66030; // @[Modules.scala 50:57:@13817.4]
  wire [10:0] buffer_3_496; // @[Modules.scala 50:57:@13818.4]
  wire [10:0] buffer_3_210; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66032; // @[Modules.scala 50:57:@13820.4]
  wire [10:0] _T_66033; // @[Modules.scala 50:57:@13821.4]
  wire [10:0] buffer_3_497; // @[Modules.scala 50:57:@13822.4]
  wire [10:0] buffer_3_212; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66035; // @[Modules.scala 50:57:@13824.4]
  wire [10:0] _T_66036; // @[Modules.scala 50:57:@13825.4]
  wire [10:0] buffer_3_498; // @[Modules.scala 50:57:@13826.4]
  wire [10:0] buffer_3_220; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66047; // @[Modules.scala 50:57:@13840.4]
  wire [10:0] _T_66048; // @[Modules.scala 50:57:@13841.4]
  wire [10:0] buffer_3_502; // @[Modules.scala 50:57:@13842.4]
  wire [10:0] buffer_3_222; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_223; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66050; // @[Modules.scala 50:57:@13844.4]
  wire [10:0] _T_66051; // @[Modules.scala 50:57:@13845.4]
  wire [10:0] buffer_3_503; // @[Modules.scala 50:57:@13846.4]
  wire [10:0] buffer_3_224; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66053; // @[Modules.scala 50:57:@13848.4]
  wire [10:0] _T_66054; // @[Modules.scala 50:57:@13849.4]
  wire [10:0] buffer_3_504; // @[Modules.scala 50:57:@13850.4]
  wire [10:0] buffer_3_226; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66056; // @[Modules.scala 50:57:@13852.4]
  wire [10:0] _T_66057; // @[Modules.scala 50:57:@13853.4]
  wire [10:0] buffer_3_505; // @[Modules.scala 50:57:@13854.4]
  wire [10:0] buffer_3_228; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66059; // @[Modules.scala 50:57:@13856.4]
  wire [10:0] _T_66060; // @[Modules.scala 50:57:@13857.4]
  wire [10:0] buffer_3_506; // @[Modules.scala 50:57:@13858.4]
  wire [11:0] _T_66065; // @[Modules.scala 50:57:@13864.4]
  wire [10:0] _T_66066; // @[Modules.scala 50:57:@13865.4]
  wire [10:0] buffer_3_508; // @[Modules.scala 50:57:@13866.4]
  wire [10:0] buffer_3_236; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_237; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66071; // @[Modules.scala 50:57:@13872.4]
  wire [10:0] _T_66072; // @[Modules.scala 50:57:@13873.4]
  wire [10:0] buffer_3_510; // @[Modules.scala 50:57:@13874.4]
  wire [11:0] _T_66074; // @[Modules.scala 50:57:@13876.4]
  wire [10:0] _T_66075; // @[Modules.scala 50:57:@13877.4]
  wire [10:0] buffer_3_511; // @[Modules.scala 50:57:@13878.4]
  wire [10:0] buffer_3_240; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66077; // @[Modules.scala 50:57:@13880.4]
  wire [10:0] _T_66078; // @[Modules.scala 50:57:@13881.4]
  wire [10:0] buffer_3_512; // @[Modules.scala 50:57:@13882.4]
  wire [10:0] buffer_3_246; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66086; // @[Modules.scala 50:57:@13892.4]
  wire [10:0] _T_66087; // @[Modules.scala 50:57:@13893.4]
  wire [10:0] buffer_3_515; // @[Modules.scala 50:57:@13894.4]
  wire [10:0] buffer_3_250; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_251; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66092; // @[Modules.scala 50:57:@13900.4]
  wire [10:0] _T_66093; // @[Modules.scala 50:57:@13901.4]
  wire [10:0] buffer_3_517; // @[Modules.scala 50:57:@13902.4]
  wire [10:0] buffer_3_252; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66095; // @[Modules.scala 50:57:@13904.4]
  wire [10:0] _T_66096; // @[Modules.scala 50:57:@13905.4]
  wire [10:0] buffer_3_518; // @[Modules.scala 50:57:@13906.4]
  wire [10:0] buffer_3_254; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66098; // @[Modules.scala 50:57:@13908.4]
  wire [10:0] _T_66099; // @[Modules.scala 50:57:@13909.4]
  wire [10:0] buffer_3_519; // @[Modules.scala 50:57:@13910.4]
  wire [10:0] buffer_3_257; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66101; // @[Modules.scala 50:57:@13912.4]
  wire [10:0] _T_66102; // @[Modules.scala 50:57:@13913.4]
  wire [10:0] buffer_3_520; // @[Modules.scala 50:57:@13914.4]
  wire [10:0] buffer_3_265; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66113; // @[Modules.scala 50:57:@13928.4]
  wire [10:0] _T_66114; // @[Modules.scala 50:57:@13929.4]
  wire [10:0] buffer_3_524; // @[Modules.scala 50:57:@13930.4]
  wire [10:0] buffer_3_270; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_271; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66122; // @[Modules.scala 50:57:@13940.4]
  wire [10:0] _T_66123; // @[Modules.scala 50:57:@13941.4]
  wire [10:0] buffer_3_527; // @[Modules.scala 50:57:@13942.4]
  wire [10:0] buffer_3_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66125; // @[Modules.scala 50:57:@13944.4]
  wire [10:0] _T_66126; // @[Modules.scala 50:57:@13945.4]
  wire [10:0] buffer_3_528; // @[Modules.scala 50:57:@13946.4]
  wire [10:0] buffer_3_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66128; // @[Modules.scala 50:57:@13948.4]
  wire [10:0] _T_66129; // @[Modules.scala 50:57:@13949.4]
  wire [10:0] buffer_3_529; // @[Modules.scala 50:57:@13950.4]
  wire [10:0] buffer_3_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66131; // @[Modules.scala 50:57:@13952.4]
  wire [10:0] _T_66132; // @[Modules.scala 50:57:@13953.4]
  wire [10:0] buffer_3_530; // @[Modules.scala 50:57:@13954.4]
  wire [10:0] buffer_3_278; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66134; // @[Modules.scala 50:57:@13956.4]
  wire [10:0] _T_66135; // @[Modules.scala 50:57:@13957.4]
  wire [10:0] buffer_3_531; // @[Modules.scala 50:57:@13958.4]
  wire [11:0] _T_66137; // @[Modules.scala 50:57:@13960.4]
  wire [10:0] _T_66138; // @[Modules.scala 50:57:@13961.4]
  wire [10:0] buffer_3_532; // @[Modules.scala 50:57:@13962.4]
  wire [10:0] buffer_3_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66140; // @[Modules.scala 50:57:@13964.4]
  wire [10:0] _T_66141; // @[Modules.scala 50:57:@13965.4]
  wire [10:0] buffer_3_533; // @[Modules.scala 50:57:@13966.4]
  wire [10:0] buffer_3_286; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66146; // @[Modules.scala 50:57:@13972.4]
  wire [10:0] _T_66147; // @[Modules.scala 50:57:@13973.4]
  wire [10:0] buffer_3_535; // @[Modules.scala 50:57:@13974.4]
  wire [11:0] _T_66149; // @[Modules.scala 50:57:@13976.4]
  wire [10:0] _T_66150; // @[Modules.scala 50:57:@13977.4]
  wire [10:0] buffer_3_536; // @[Modules.scala 50:57:@13978.4]
  wire [10:0] buffer_3_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66152; // @[Modules.scala 50:57:@13980.4]
  wire [10:0] _T_66153; // @[Modules.scala 50:57:@13981.4]
  wire [10:0] buffer_3_537; // @[Modules.scala 50:57:@13982.4]
  wire [10:0] buffer_3_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66155; // @[Modules.scala 50:57:@13984.4]
  wire [10:0] _T_66156; // @[Modules.scala 50:57:@13985.4]
  wire [10:0] buffer_3_538; // @[Modules.scala 50:57:@13986.4]
  wire [10:0] buffer_3_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66161; // @[Modules.scala 50:57:@13992.4]
  wire [10:0] _T_66162; // @[Modules.scala 50:57:@13993.4]
  wire [10:0] buffer_3_540; // @[Modules.scala 50:57:@13994.4]
  wire [11:0] _T_66164; // @[Modules.scala 50:57:@13996.4]
  wire [10:0] _T_66165; // @[Modules.scala 50:57:@13997.4]
  wire [10:0] buffer_3_541; // @[Modules.scala 50:57:@13998.4]
  wire [10:0] buffer_3_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66167; // @[Modules.scala 50:57:@14000.4]
  wire [10:0] _T_66168; // @[Modules.scala 50:57:@14001.4]
  wire [10:0] buffer_3_542; // @[Modules.scala 50:57:@14002.4]
  wire [11:0] _T_66170; // @[Modules.scala 50:57:@14004.4]
  wire [10:0] _T_66171; // @[Modules.scala 50:57:@14005.4]
  wire [10:0] buffer_3_543; // @[Modules.scala 50:57:@14006.4]
  wire [10:0] buffer_3_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66173; // @[Modules.scala 50:57:@14008.4]
  wire [10:0] _T_66174; // @[Modules.scala 50:57:@14009.4]
  wire [10:0] buffer_3_544; // @[Modules.scala 50:57:@14010.4]
  wire [10:0] buffer_3_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66176; // @[Modules.scala 50:57:@14012.4]
  wire [10:0] _T_66177; // @[Modules.scala 50:57:@14013.4]
  wire [10:0] buffer_3_545; // @[Modules.scala 50:57:@14014.4]
  wire [10:0] buffer_3_310; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66182; // @[Modules.scala 50:57:@14020.4]
  wire [10:0] _T_66183; // @[Modules.scala 50:57:@14021.4]
  wire [10:0] buffer_3_547; // @[Modules.scala 50:57:@14022.4]
  wire [10:0] buffer_3_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66185; // @[Modules.scala 50:57:@14024.4]
  wire [10:0] _T_66186; // @[Modules.scala 50:57:@14025.4]
  wire [10:0] buffer_3_548; // @[Modules.scala 50:57:@14026.4]
  wire [10:0] buffer_3_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66188; // @[Modules.scala 50:57:@14028.4]
  wire [10:0] _T_66189; // @[Modules.scala 50:57:@14029.4]
  wire [10:0] buffer_3_549; // @[Modules.scala 50:57:@14030.4]
  wire [10:0] buffer_3_316; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66191; // @[Modules.scala 50:57:@14032.4]
  wire [10:0] _T_66192; // @[Modules.scala 50:57:@14033.4]
  wire [10:0] buffer_3_550; // @[Modules.scala 50:57:@14034.4]
  wire [10:0] buffer_3_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66194; // @[Modules.scala 50:57:@14036.4]
  wire [10:0] _T_66195; // @[Modules.scala 50:57:@14037.4]
  wire [10:0] buffer_3_551; // @[Modules.scala 50:57:@14038.4]
  wire [10:0] buffer_3_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66197; // @[Modules.scala 50:57:@14040.4]
  wire [10:0] _T_66198; // @[Modules.scala 50:57:@14041.4]
  wire [10:0] buffer_3_552; // @[Modules.scala 50:57:@14042.4]
  wire [11:0] _T_66200; // @[Modules.scala 50:57:@14044.4]
  wire [10:0] _T_66201; // @[Modules.scala 50:57:@14045.4]
  wire [10:0] buffer_3_553; // @[Modules.scala 50:57:@14046.4]
  wire [10:0] buffer_3_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66203; // @[Modules.scala 50:57:@14048.4]
  wire [10:0] _T_66204; // @[Modules.scala 50:57:@14049.4]
  wire [10:0] buffer_3_554; // @[Modules.scala 50:57:@14050.4]
  wire [10:0] buffer_3_326; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66206; // @[Modules.scala 50:57:@14052.4]
  wire [10:0] _T_66207; // @[Modules.scala 50:57:@14053.4]
  wire [10:0] buffer_3_555; // @[Modules.scala 50:57:@14054.4]
  wire [11:0] _T_66209; // @[Modules.scala 50:57:@14056.4]
  wire [10:0] _T_66210; // @[Modules.scala 50:57:@14057.4]
  wire [10:0] buffer_3_556; // @[Modules.scala 50:57:@14058.4]
  wire [10:0] buffer_3_331; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66212; // @[Modules.scala 50:57:@14060.4]
  wire [10:0] _T_66213; // @[Modules.scala 50:57:@14061.4]
  wire [10:0] buffer_3_557; // @[Modules.scala 50:57:@14062.4]
  wire [10:0] buffer_3_333; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66215; // @[Modules.scala 50:57:@14064.4]
  wire [10:0] _T_66216; // @[Modules.scala 50:57:@14065.4]
  wire [10:0] buffer_3_558; // @[Modules.scala 50:57:@14066.4]
  wire [10:0] buffer_3_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66218; // @[Modules.scala 50:57:@14068.4]
  wire [10:0] _T_66219; // @[Modules.scala 50:57:@14069.4]
  wire [10:0] buffer_3_559; // @[Modules.scala 50:57:@14070.4]
  wire [10:0] buffer_3_336; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66221; // @[Modules.scala 50:57:@14072.4]
  wire [10:0] _T_66222; // @[Modules.scala 50:57:@14073.4]
  wire [10:0] buffer_3_560; // @[Modules.scala 50:57:@14074.4]
  wire [11:0] _T_66227; // @[Modules.scala 50:57:@14080.4]
  wire [10:0] _T_66228; // @[Modules.scala 50:57:@14081.4]
  wire [10:0] buffer_3_562; // @[Modules.scala 50:57:@14082.4]
  wire [10:0] buffer_3_342; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66230; // @[Modules.scala 50:57:@14084.4]
  wire [10:0] _T_66231; // @[Modules.scala 50:57:@14085.4]
  wire [10:0] buffer_3_563; // @[Modules.scala 50:57:@14086.4]
  wire [10:0] buffer_3_344; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66233; // @[Modules.scala 50:57:@14088.4]
  wire [10:0] _T_66234; // @[Modules.scala 50:57:@14089.4]
  wire [10:0] buffer_3_564; // @[Modules.scala 50:57:@14090.4]
  wire [10:0] buffer_3_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66236; // @[Modules.scala 50:57:@14092.4]
  wire [10:0] _T_66237; // @[Modules.scala 50:57:@14093.4]
  wire [10:0] buffer_3_565; // @[Modules.scala 50:57:@14094.4]
  wire [10:0] buffer_3_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66239; // @[Modules.scala 50:57:@14096.4]
  wire [10:0] _T_66240; // @[Modules.scala 50:57:@14097.4]
  wire [10:0] buffer_3_566; // @[Modules.scala 50:57:@14098.4]
  wire [10:0] buffer_3_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66242; // @[Modules.scala 50:57:@14100.4]
  wire [10:0] _T_66243; // @[Modules.scala 50:57:@14101.4]
  wire [10:0] buffer_3_567; // @[Modules.scala 50:57:@14102.4]
  wire [10:0] buffer_3_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66248; // @[Modules.scala 50:57:@14108.4]
  wire [10:0] _T_66249; // @[Modules.scala 50:57:@14109.4]
  wire [10:0] buffer_3_569; // @[Modules.scala 50:57:@14110.4]
  wire [10:0] buffer_3_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66257; // @[Modules.scala 50:57:@14120.4]
  wire [10:0] _T_66258; // @[Modules.scala 50:57:@14121.4]
  wire [10:0] buffer_3_572; // @[Modules.scala 50:57:@14122.4]
  wire [11:0] _T_66260; // @[Modules.scala 50:57:@14124.4]
  wire [10:0] _T_66261; // @[Modules.scala 50:57:@14125.4]
  wire [10:0] buffer_3_573; // @[Modules.scala 50:57:@14126.4]
  wire [10:0] buffer_3_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66263; // @[Modules.scala 50:57:@14128.4]
  wire [10:0] _T_66264; // @[Modules.scala 50:57:@14129.4]
  wire [10:0] buffer_3_574; // @[Modules.scala 50:57:@14130.4]
  wire [10:0] buffer_3_368; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_369; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66269; // @[Modules.scala 50:57:@14136.4]
  wire [10:0] _T_66270; // @[Modules.scala 50:57:@14137.4]
  wire [10:0] buffer_3_576; // @[Modules.scala 50:57:@14138.4]
  wire [10:0] buffer_3_370; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66272; // @[Modules.scala 50:57:@14140.4]
  wire [10:0] _T_66273; // @[Modules.scala 50:57:@14141.4]
  wire [10:0] buffer_3_577; // @[Modules.scala 50:57:@14142.4]
  wire [10:0] buffer_3_372; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_373; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66275; // @[Modules.scala 50:57:@14144.4]
  wire [10:0] _T_66276; // @[Modules.scala 50:57:@14145.4]
  wire [10:0] buffer_3_578; // @[Modules.scala 50:57:@14146.4]
  wire [10:0] buffer_3_374; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66278; // @[Modules.scala 50:57:@14148.4]
  wire [10:0] _T_66279; // @[Modules.scala 50:57:@14149.4]
  wire [10:0] buffer_3_579; // @[Modules.scala 50:57:@14150.4]
  wire [10:0] buffer_3_376; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66281; // @[Modules.scala 50:57:@14152.4]
  wire [10:0] _T_66282; // @[Modules.scala 50:57:@14153.4]
  wire [10:0] buffer_3_580; // @[Modules.scala 50:57:@14154.4]
  wire [10:0] buffer_3_378; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66284; // @[Modules.scala 50:57:@14156.4]
  wire [10:0] _T_66285; // @[Modules.scala 50:57:@14157.4]
  wire [10:0] buffer_3_581; // @[Modules.scala 50:57:@14158.4]
  wire [10:0] buffer_3_382; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66290; // @[Modules.scala 50:57:@14164.4]
  wire [10:0] _T_66291; // @[Modules.scala 50:57:@14165.4]
  wire [10:0] buffer_3_583; // @[Modules.scala 50:57:@14166.4]
  wire [10:0] buffer_3_384; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_385; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66293; // @[Modules.scala 50:57:@14168.4]
  wire [10:0] _T_66294; // @[Modules.scala 50:57:@14169.4]
  wire [10:0] buffer_3_584; // @[Modules.scala 50:57:@14170.4]
  wire [10:0] buffer_3_386; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_387; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66296; // @[Modules.scala 50:57:@14172.4]
  wire [10:0] _T_66297; // @[Modules.scala 50:57:@14173.4]
  wire [10:0] buffer_3_585; // @[Modules.scala 50:57:@14174.4]
  wire [10:0] buffer_3_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66299; // @[Modules.scala 50:57:@14176.4]
  wire [10:0] _T_66300; // @[Modules.scala 50:57:@14177.4]
  wire [10:0] buffer_3_586; // @[Modules.scala 50:57:@14178.4]
  wire [11:0] _T_66302; // @[Modules.scala 50:57:@14180.4]
  wire [10:0] _T_66303; // @[Modules.scala 50:57:@14181.4]
  wire [10:0] buffer_3_587; // @[Modules.scala 50:57:@14182.4]
  wire [11:0] _T_66305; // @[Modules.scala 53:83:@14184.4]
  wire [10:0] _T_66306; // @[Modules.scala 53:83:@14185.4]
  wire [10:0] buffer_3_588; // @[Modules.scala 53:83:@14186.4]
  wire [11:0] _T_66308; // @[Modules.scala 53:83:@14188.4]
  wire [10:0] _T_66309; // @[Modules.scala 53:83:@14189.4]
  wire [10:0] buffer_3_589; // @[Modules.scala 53:83:@14190.4]
  wire [11:0] _T_66311; // @[Modules.scala 53:83:@14192.4]
  wire [10:0] _T_66312; // @[Modules.scala 53:83:@14193.4]
  wire [10:0] buffer_3_590; // @[Modules.scala 53:83:@14194.4]
  wire [11:0] _T_66314; // @[Modules.scala 53:83:@14196.4]
  wire [10:0] _T_66315; // @[Modules.scala 53:83:@14197.4]
  wire [10:0] buffer_3_591; // @[Modules.scala 53:83:@14198.4]
  wire [11:0] _T_66317; // @[Modules.scala 53:83:@14200.4]
  wire [10:0] _T_66318; // @[Modules.scala 53:83:@14201.4]
  wire [10:0] buffer_3_592; // @[Modules.scala 53:83:@14202.4]
  wire [11:0] _T_66320; // @[Modules.scala 53:83:@14204.4]
  wire [10:0] _T_66321; // @[Modules.scala 53:83:@14205.4]
  wire [10:0] buffer_3_593; // @[Modules.scala 53:83:@14206.4]
  wire [11:0] _T_66323; // @[Modules.scala 53:83:@14208.4]
  wire [10:0] _T_66324; // @[Modules.scala 53:83:@14209.4]
  wire [10:0] buffer_3_594; // @[Modules.scala 53:83:@14210.4]
  wire [11:0] _T_66326; // @[Modules.scala 53:83:@14212.4]
  wire [10:0] _T_66327; // @[Modules.scala 53:83:@14213.4]
  wire [10:0] buffer_3_595; // @[Modules.scala 53:83:@14214.4]
  wire [11:0] _T_66329; // @[Modules.scala 53:83:@14216.4]
  wire [10:0] _T_66330; // @[Modules.scala 53:83:@14217.4]
  wire [10:0] buffer_3_596; // @[Modules.scala 53:83:@14218.4]
  wire [11:0] _T_66332; // @[Modules.scala 53:83:@14220.4]
  wire [10:0] _T_66333; // @[Modules.scala 53:83:@14221.4]
  wire [10:0] buffer_3_597; // @[Modules.scala 53:83:@14222.4]
  wire [11:0] _T_66335; // @[Modules.scala 53:83:@14224.4]
  wire [10:0] _T_66336; // @[Modules.scala 53:83:@14225.4]
  wire [10:0] buffer_3_598; // @[Modules.scala 53:83:@14226.4]
  wire [11:0] _T_66338; // @[Modules.scala 53:83:@14228.4]
  wire [10:0] _T_66339; // @[Modules.scala 53:83:@14229.4]
  wire [10:0] buffer_3_599; // @[Modules.scala 53:83:@14230.4]
  wire [11:0] _T_66341; // @[Modules.scala 53:83:@14232.4]
  wire [10:0] _T_66342; // @[Modules.scala 53:83:@14233.4]
  wire [10:0] buffer_3_600; // @[Modules.scala 53:83:@14234.4]
  wire [11:0] _T_66344; // @[Modules.scala 53:83:@14236.4]
  wire [10:0] _T_66345; // @[Modules.scala 53:83:@14237.4]
  wire [10:0] buffer_3_601; // @[Modules.scala 53:83:@14238.4]
  wire [11:0] _T_66347; // @[Modules.scala 53:83:@14240.4]
  wire [10:0] _T_66348; // @[Modules.scala 53:83:@14241.4]
  wire [10:0] buffer_3_602; // @[Modules.scala 53:83:@14242.4]
  wire [11:0] _T_66350; // @[Modules.scala 53:83:@14244.4]
  wire [10:0] _T_66351; // @[Modules.scala 53:83:@14245.4]
  wire [10:0] buffer_3_603; // @[Modules.scala 53:83:@14246.4]
  wire [11:0] _T_66353; // @[Modules.scala 53:83:@14248.4]
  wire [10:0] _T_66354; // @[Modules.scala 53:83:@14249.4]
  wire [10:0] buffer_3_604; // @[Modules.scala 53:83:@14250.4]
  wire [11:0] _T_66356; // @[Modules.scala 53:83:@14252.4]
  wire [10:0] _T_66357; // @[Modules.scala 53:83:@14253.4]
  wire [10:0] buffer_3_605; // @[Modules.scala 53:83:@14254.4]
  wire [11:0] _T_66359; // @[Modules.scala 53:83:@14256.4]
  wire [10:0] _T_66360; // @[Modules.scala 53:83:@14257.4]
  wire [10:0] buffer_3_606; // @[Modules.scala 53:83:@14258.4]
  wire [11:0] _T_66362; // @[Modules.scala 53:83:@14260.4]
  wire [10:0] _T_66363; // @[Modules.scala 53:83:@14261.4]
  wire [10:0] buffer_3_607; // @[Modules.scala 53:83:@14262.4]
  wire [11:0] _T_66368; // @[Modules.scala 53:83:@14268.4]
  wire [10:0] _T_66369; // @[Modules.scala 53:83:@14269.4]
  wire [10:0] buffer_3_609; // @[Modules.scala 53:83:@14270.4]
  wire [11:0] _T_66371; // @[Modules.scala 53:83:@14272.4]
  wire [10:0] _T_66372; // @[Modules.scala 53:83:@14273.4]
  wire [10:0] buffer_3_610; // @[Modules.scala 53:83:@14274.4]
  wire [11:0] _T_66374; // @[Modules.scala 53:83:@14276.4]
  wire [10:0] _T_66375; // @[Modules.scala 53:83:@14277.4]
  wire [10:0] buffer_3_611; // @[Modules.scala 53:83:@14278.4]
  wire [11:0] _T_66377; // @[Modules.scala 53:83:@14280.4]
  wire [10:0] _T_66378; // @[Modules.scala 53:83:@14281.4]
  wire [10:0] buffer_3_612; // @[Modules.scala 53:83:@14282.4]
  wire [11:0] _T_66380; // @[Modules.scala 53:83:@14284.4]
  wire [10:0] _T_66381; // @[Modules.scala 53:83:@14285.4]
  wire [10:0] buffer_3_613; // @[Modules.scala 53:83:@14286.4]
  wire [11:0] _T_66383; // @[Modules.scala 53:83:@14288.4]
  wire [10:0] _T_66384; // @[Modules.scala 53:83:@14289.4]
  wire [10:0] buffer_3_614; // @[Modules.scala 53:83:@14290.4]
  wire [11:0] _T_66386; // @[Modules.scala 53:83:@14292.4]
  wire [10:0] _T_66387; // @[Modules.scala 53:83:@14293.4]
  wire [10:0] buffer_3_615; // @[Modules.scala 53:83:@14294.4]
  wire [11:0] _T_66389; // @[Modules.scala 53:83:@14296.4]
  wire [10:0] _T_66390; // @[Modules.scala 53:83:@14297.4]
  wire [10:0] buffer_3_616; // @[Modules.scala 53:83:@14298.4]
  wire [11:0] _T_66392; // @[Modules.scala 53:83:@14300.4]
  wire [10:0] _T_66393; // @[Modules.scala 53:83:@14301.4]
  wire [10:0] buffer_3_617; // @[Modules.scala 53:83:@14302.4]
  wire [11:0] _T_66395; // @[Modules.scala 53:83:@14304.4]
  wire [10:0] _T_66396; // @[Modules.scala 53:83:@14305.4]
  wire [10:0] buffer_3_618; // @[Modules.scala 53:83:@14306.4]
  wire [11:0] _T_66398; // @[Modules.scala 53:83:@14308.4]
  wire [10:0] _T_66399; // @[Modules.scala 53:83:@14309.4]
  wire [10:0] buffer_3_619; // @[Modules.scala 53:83:@14310.4]
  wire [11:0] _T_66401; // @[Modules.scala 53:83:@14312.4]
  wire [10:0] _T_66402; // @[Modules.scala 53:83:@14313.4]
  wire [10:0] buffer_3_620; // @[Modules.scala 53:83:@14314.4]
  wire [11:0] _T_66404; // @[Modules.scala 53:83:@14316.4]
  wire [10:0] _T_66405; // @[Modules.scala 53:83:@14317.4]
  wire [10:0] buffer_3_621; // @[Modules.scala 53:83:@14318.4]
  wire [11:0] _T_66407; // @[Modules.scala 53:83:@14320.4]
  wire [10:0] _T_66408; // @[Modules.scala 53:83:@14321.4]
  wire [10:0] buffer_3_622; // @[Modules.scala 53:83:@14322.4]
  wire [11:0] _T_66410; // @[Modules.scala 53:83:@14324.4]
  wire [10:0] _T_66411; // @[Modules.scala 53:83:@14325.4]
  wire [10:0] buffer_3_623; // @[Modules.scala 53:83:@14326.4]
  wire [11:0] _T_66413; // @[Modules.scala 53:83:@14328.4]
  wire [10:0] _T_66414; // @[Modules.scala 53:83:@14329.4]
  wire [10:0] buffer_3_624; // @[Modules.scala 53:83:@14330.4]
  wire [11:0] _T_66416; // @[Modules.scala 53:83:@14332.4]
  wire [10:0] _T_66417; // @[Modules.scala 53:83:@14333.4]
  wire [10:0] buffer_3_625; // @[Modules.scala 53:83:@14334.4]
  wire [11:0] _T_66419; // @[Modules.scala 53:83:@14336.4]
  wire [10:0] _T_66420; // @[Modules.scala 53:83:@14337.4]
  wire [10:0] buffer_3_626; // @[Modules.scala 53:83:@14338.4]
  wire [11:0] _T_66422; // @[Modules.scala 53:83:@14340.4]
  wire [10:0] _T_66423; // @[Modules.scala 53:83:@14341.4]
  wire [10:0] buffer_3_627; // @[Modules.scala 53:83:@14342.4]
  wire [11:0] _T_66425; // @[Modules.scala 53:83:@14344.4]
  wire [10:0] _T_66426; // @[Modules.scala 53:83:@14345.4]
  wire [10:0] buffer_3_628; // @[Modules.scala 53:83:@14346.4]
  wire [11:0] _T_66428; // @[Modules.scala 53:83:@14348.4]
  wire [10:0] _T_66429; // @[Modules.scala 53:83:@14349.4]
  wire [10:0] buffer_3_629; // @[Modules.scala 53:83:@14350.4]
  wire [11:0] _T_66431; // @[Modules.scala 53:83:@14352.4]
  wire [10:0] _T_66432; // @[Modules.scala 53:83:@14353.4]
  wire [10:0] buffer_3_630; // @[Modules.scala 53:83:@14354.4]
  wire [11:0] _T_66434; // @[Modules.scala 53:83:@14356.4]
  wire [10:0] _T_66435; // @[Modules.scala 53:83:@14357.4]
  wire [10:0] buffer_3_631; // @[Modules.scala 53:83:@14358.4]
  wire [11:0] _T_66440; // @[Modules.scala 53:83:@14364.4]
  wire [10:0] _T_66441; // @[Modules.scala 53:83:@14365.4]
  wire [10:0] buffer_3_633; // @[Modules.scala 53:83:@14366.4]
  wire [11:0] _T_66443; // @[Modules.scala 53:83:@14368.4]
  wire [10:0] _T_66444; // @[Modules.scala 53:83:@14369.4]
  wire [10:0] buffer_3_634; // @[Modules.scala 53:83:@14370.4]
  wire [11:0] _T_66446; // @[Modules.scala 53:83:@14372.4]
  wire [10:0] _T_66447; // @[Modules.scala 53:83:@14373.4]
  wire [10:0] buffer_3_635; // @[Modules.scala 53:83:@14374.4]
  wire [11:0] _T_66449; // @[Modules.scala 53:83:@14376.4]
  wire [10:0] _T_66450; // @[Modules.scala 53:83:@14377.4]
  wire [10:0] buffer_3_636; // @[Modules.scala 53:83:@14378.4]
  wire [11:0] _T_66452; // @[Modules.scala 53:83:@14380.4]
  wire [10:0] _T_66453; // @[Modules.scala 53:83:@14381.4]
  wire [10:0] buffer_3_637; // @[Modules.scala 53:83:@14382.4]
  wire [11:0] _T_66455; // @[Modules.scala 53:83:@14384.4]
  wire [10:0] _T_66456; // @[Modules.scala 53:83:@14385.4]
  wire [10:0] buffer_3_638; // @[Modules.scala 53:83:@14386.4]
  wire [11:0] _T_66458; // @[Modules.scala 53:83:@14388.4]
  wire [10:0] _T_66459; // @[Modules.scala 53:83:@14389.4]
  wire [10:0] buffer_3_639; // @[Modules.scala 53:83:@14390.4]
  wire [11:0] _T_66461; // @[Modules.scala 53:83:@14392.4]
  wire [10:0] _T_66462; // @[Modules.scala 53:83:@14393.4]
  wire [10:0] buffer_3_640; // @[Modules.scala 53:83:@14394.4]
  wire [11:0] _T_66464; // @[Modules.scala 53:83:@14396.4]
  wire [10:0] _T_66465; // @[Modules.scala 53:83:@14397.4]
  wire [10:0] buffer_3_641; // @[Modules.scala 53:83:@14398.4]
  wire [11:0] _T_66467; // @[Modules.scala 53:83:@14400.4]
  wire [10:0] _T_66468; // @[Modules.scala 53:83:@14401.4]
  wire [10:0] buffer_3_642; // @[Modules.scala 53:83:@14402.4]
  wire [11:0] _T_66470; // @[Modules.scala 53:83:@14404.4]
  wire [10:0] _T_66471; // @[Modules.scala 53:83:@14405.4]
  wire [10:0] buffer_3_643; // @[Modules.scala 53:83:@14406.4]
  wire [11:0] _T_66473; // @[Modules.scala 53:83:@14408.4]
  wire [10:0] _T_66474; // @[Modules.scala 53:83:@14409.4]
  wire [10:0] buffer_3_644; // @[Modules.scala 53:83:@14410.4]
  wire [11:0] _T_66476; // @[Modules.scala 53:83:@14412.4]
  wire [10:0] _T_66477; // @[Modules.scala 53:83:@14413.4]
  wire [10:0] buffer_3_645; // @[Modules.scala 53:83:@14414.4]
  wire [11:0] _T_66479; // @[Modules.scala 53:83:@14416.4]
  wire [10:0] _T_66480; // @[Modules.scala 53:83:@14417.4]
  wire [10:0] buffer_3_646; // @[Modules.scala 53:83:@14418.4]
  wire [11:0] _T_66482; // @[Modules.scala 53:83:@14420.4]
  wire [10:0] _T_66483; // @[Modules.scala 53:83:@14421.4]
  wire [10:0] buffer_3_647; // @[Modules.scala 53:83:@14422.4]
  wire [11:0] _T_66485; // @[Modules.scala 53:83:@14424.4]
  wire [10:0] _T_66486; // @[Modules.scala 53:83:@14425.4]
  wire [10:0] buffer_3_648; // @[Modules.scala 53:83:@14426.4]
  wire [11:0] _T_66488; // @[Modules.scala 53:83:@14428.4]
  wire [10:0] _T_66489; // @[Modules.scala 53:83:@14429.4]
  wire [10:0] buffer_3_649; // @[Modules.scala 53:83:@14430.4]
  wire [11:0] _T_66491; // @[Modules.scala 53:83:@14432.4]
  wire [10:0] _T_66492; // @[Modules.scala 53:83:@14433.4]
  wire [10:0] buffer_3_650; // @[Modules.scala 53:83:@14434.4]
  wire [11:0] _T_66494; // @[Modules.scala 53:83:@14436.4]
  wire [10:0] _T_66495; // @[Modules.scala 53:83:@14437.4]
  wire [10:0] buffer_3_651; // @[Modules.scala 53:83:@14438.4]
  wire [11:0] _T_66497; // @[Modules.scala 53:83:@14440.4]
  wire [10:0] _T_66498; // @[Modules.scala 53:83:@14441.4]
  wire [10:0] buffer_3_652; // @[Modules.scala 53:83:@14442.4]
  wire [11:0] _T_66500; // @[Modules.scala 53:83:@14444.4]
  wire [10:0] _T_66501; // @[Modules.scala 53:83:@14445.4]
  wire [10:0] buffer_3_653; // @[Modules.scala 53:83:@14446.4]
  wire [11:0] _T_66503; // @[Modules.scala 53:83:@14448.4]
  wire [10:0] _T_66504; // @[Modules.scala 53:83:@14449.4]
  wire [10:0] buffer_3_654; // @[Modules.scala 53:83:@14450.4]
  wire [11:0] _T_66506; // @[Modules.scala 53:83:@14452.4]
  wire [10:0] _T_66507; // @[Modules.scala 53:83:@14453.4]
  wire [10:0] buffer_3_655; // @[Modules.scala 53:83:@14454.4]
  wire [11:0] _T_66509; // @[Modules.scala 53:83:@14456.4]
  wire [10:0] _T_66510; // @[Modules.scala 53:83:@14457.4]
  wire [10:0] buffer_3_656; // @[Modules.scala 53:83:@14458.4]
  wire [11:0] _T_66512; // @[Modules.scala 53:83:@14460.4]
  wire [10:0] _T_66513; // @[Modules.scala 53:83:@14461.4]
  wire [10:0] buffer_3_657; // @[Modules.scala 53:83:@14462.4]
  wire [11:0] _T_66515; // @[Modules.scala 53:83:@14464.4]
  wire [10:0] _T_66516; // @[Modules.scala 53:83:@14465.4]
  wire [10:0] buffer_3_658; // @[Modules.scala 53:83:@14466.4]
  wire [11:0] _T_66518; // @[Modules.scala 53:83:@14468.4]
  wire [10:0] _T_66519; // @[Modules.scala 53:83:@14469.4]
  wire [10:0] buffer_3_659; // @[Modules.scala 53:83:@14470.4]
  wire [11:0] _T_66521; // @[Modules.scala 53:83:@14472.4]
  wire [10:0] _T_66522; // @[Modules.scala 53:83:@14473.4]
  wire [10:0] buffer_3_660; // @[Modules.scala 53:83:@14474.4]
  wire [11:0] _T_66524; // @[Modules.scala 53:83:@14476.4]
  wire [10:0] _T_66525; // @[Modules.scala 53:83:@14477.4]
  wire [10:0] buffer_3_661; // @[Modules.scala 53:83:@14478.4]
  wire [11:0] _T_66527; // @[Modules.scala 53:83:@14480.4]
  wire [10:0] _T_66528; // @[Modules.scala 53:83:@14481.4]
  wire [10:0] buffer_3_662; // @[Modules.scala 53:83:@14482.4]
  wire [11:0] _T_66530; // @[Modules.scala 53:83:@14484.4]
  wire [10:0] _T_66531; // @[Modules.scala 53:83:@14485.4]
  wire [10:0] buffer_3_663; // @[Modules.scala 53:83:@14486.4]
  wire [11:0] _T_66533; // @[Modules.scala 53:83:@14488.4]
  wire [10:0] _T_66534; // @[Modules.scala 53:83:@14489.4]
  wire [10:0] buffer_3_664; // @[Modules.scala 53:83:@14490.4]
  wire [11:0] _T_66536; // @[Modules.scala 53:83:@14492.4]
  wire [10:0] _T_66537; // @[Modules.scala 53:83:@14493.4]
  wire [10:0] buffer_3_665; // @[Modules.scala 53:83:@14494.4]
  wire [11:0] _T_66539; // @[Modules.scala 53:83:@14496.4]
  wire [10:0] _T_66540; // @[Modules.scala 53:83:@14497.4]
  wire [10:0] buffer_3_666; // @[Modules.scala 53:83:@14498.4]
  wire [11:0] _T_66542; // @[Modules.scala 53:83:@14500.4]
  wire [10:0] _T_66543; // @[Modules.scala 53:83:@14501.4]
  wire [10:0] buffer_3_667; // @[Modules.scala 53:83:@14502.4]
  wire [11:0] _T_66545; // @[Modules.scala 53:83:@14504.4]
  wire [10:0] _T_66546; // @[Modules.scala 53:83:@14505.4]
  wire [10:0] buffer_3_668; // @[Modules.scala 53:83:@14506.4]
  wire [11:0] _T_66548; // @[Modules.scala 53:83:@14508.4]
  wire [10:0] _T_66549; // @[Modules.scala 53:83:@14509.4]
  wire [10:0] buffer_3_669; // @[Modules.scala 53:83:@14510.4]
  wire [11:0] _T_66551; // @[Modules.scala 53:83:@14512.4]
  wire [10:0] _T_66552; // @[Modules.scala 53:83:@14513.4]
  wire [10:0] buffer_3_670; // @[Modules.scala 53:83:@14514.4]
  wire [11:0] _T_66554; // @[Modules.scala 53:83:@14516.4]
  wire [10:0] _T_66555; // @[Modules.scala 53:83:@14517.4]
  wire [10:0] buffer_3_671; // @[Modules.scala 53:83:@14518.4]
  wire [11:0] _T_66557; // @[Modules.scala 53:83:@14520.4]
  wire [10:0] _T_66558; // @[Modules.scala 53:83:@14521.4]
  wire [10:0] buffer_3_672; // @[Modules.scala 53:83:@14522.4]
  wire [11:0] _T_66560; // @[Modules.scala 53:83:@14524.4]
  wire [10:0] _T_66561; // @[Modules.scala 53:83:@14525.4]
  wire [10:0] buffer_3_673; // @[Modules.scala 53:83:@14526.4]
  wire [11:0] _T_66563; // @[Modules.scala 53:83:@14528.4]
  wire [10:0] _T_66564; // @[Modules.scala 53:83:@14529.4]
  wire [10:0] buffer_3_674; // @[Modules.scala 53:83:@14530.4]
  wire [11:0] _T_66566; // @[Modules.scala 53:83:@14532.4]
  wire [10:0] _T_66567; // @[Modules.scala 53:83:@14533.4]
  wire [10:0] buffer_3_675; // @[Modules.scala 53:83:@14534.4]
  wire [11:0] _T_66569; // @[Modules.scala 53:83:@14536.4]
  wire [10:0] _T_66570; // @[Modules.scala 53:83:@14537.4]
  wire [10:0] buffer_3_676; // @[Modules.scala 53:83:@14538.4]
  wire [11:0] _T_66572; // @[Modules.scala 53:83:@14540.4]
  wire [10:0] _T_66573; // @[Modules.scala 53:83:@14541.4]
  wire [10:0] buffer_3_677; // @[Modules.scala 53:83:@14542.4]
  wire [11:0] _T_66575; // @[Modules.scala 53:83:@14544.4]
  wire [10:0] _T_66576; // @[Modules.scala 53:83:@14545.4]
  wire [10:0] buffer_3_678; // @[Modules.scala 53:83:@14546.4]
  wire [11:0] _T_66578; // @[Modules.scala 53:83:@14548.4]
  wire [10:0] _T_66579; // @[Modules.scala 53:83:@14549.4]
  wire [10:0] buffer_3_679; // @[Modules.scala 53:83:@14550.4]
  wire [11:0] _T_66581; // @[Modules.scala 53:83:@14552.4]
  wire [10:0] _T_66582; // @[Modules.scala 53:83:@14553.4]
  wire [10:0] buffer_3_680; // @[Modules.scala 53:83:@14554.4]
  wire [11:0] _T_66584; // @[Modules.scala 53:83:@14556.4]
  wire [10:0] _T_66585; // @[Modules.scala 53:83:@14557.4]
  wire [10:0] buffer_3_681; // @[Modules.scala 53:83:@14558.4]
  wire [11:0] _T_66587; // @[Modules.scala 53:83:@14560.4]
  wire [10:0] _T_66588; // @[Modules.scala 53:83:@14561.4]
  wire [10:0] buffer_3_682; // @[Modules.scala 53:83:@14562.4]
  wire [11:0] _T_66590; // @[Modules.scala 53:83:@14564.4]
  wire [10:0] _T_66591; // @[Modules.scala 53:83:@14565.4]
  wire [10:0] buffer_3_683; // @[Modules.scala 53:83:@14566.4]
  wire [11:0] _T_66593; // @[Modules.scala 53:83:@14568.4]
  wire [10:0] _T_66594; // @[Modules.scala 53:83:@14569.4]
  wire [10:0] buffer_3_684; // @[Modules.scala 53:83:@14570.4]
  wire [11:0] _T_66596; // @[Modules.scala 53:83:@14572.4]
  wire [10:0] _T_66597; // @[Modules.scala 53:83:@14573.4]
  wire [10:0] buffer_3_685; // @[Modules.scala 53:83:@14574.4]
  wire [11:0] _T_66599; // @[Modules.scala 56:109:@14576.4]
  wire [10:0] _T_66600; // @[Modules.scala 56:109:@14577.4]
  wire [10:0] buffer_3_686; // @[Modules.scala 56:109:@14578.4]
  wire [11:0] _T_66602; // @[Modules.scala 56:109:@14580.4]
  wire [10:0] _T_66603; // @[Modules.scala 56:109:@14581.4]
  wire [10:0] buffer_3_687; // @[Modules.scala 56:109:@14582.4]
  wire [11:0] _T_66605; // @[Modules.scala 56:109:@14584.4]
  wire [10:0] _T_66606; // @[Modules.scala 56:109:@14585.4]
  wire [10:0] buffer_3_688; // @[Modules.scala 56:109:@14586.4]
  wire [11:0] _T_66608; // @[Modules.scala 56:109:@14588.4]
  wire [10:0] _T_66609; // @[Modules.scala 56:109:@14589.4]
  wire [10:0] buffer_3_689; // @[Modules.scala 56:109:@14590.4]
  wire [11:0] _T_66611; // @[Modules.scala 56:109:@14592.4]
  wire [10:0] _T_66612; // @[Modules.scala 56:109:@14593.4]
  wire [10:0] buffer_3_690; // @[Modules.scala 56:109:@14594.4]
  wire [11:0] _T_66614; // @[Modules.scala 56:109:@14596.4]
  wire [10:0] _T_66615; // @[Modules.scala 56:109:@14597.4]
  wire [10:0] buffer_3_691; // @[Modules.scala 56:109:@14598.4]
  wire [11:0] _T_66617; // @[Modules.scala 56:109:@14600.4]
  wire [10:0] _T_66618; // @[Modules.scala 56:109:@14601.4]
  wire [10:0] buffer_3_692; // @[Modules.scala 56:109:@14602.4]
  wire [11:0] _T_66620; // @[Modules.scala 56:109:@14604.4]
  wire [10:0] _T_66621; // @[Modules.scala 56:109:@14605.4]
  wire [10:0] buffer_3_693; // @[Modules.scala 56:109:@14606.4]
  wire [11:0] _T_66623; // @[Modules.scala 56:109:@14608.4]
  wire [10:0] _T_66624; // @[Modules.scala 56:109:@14609.4]
  wire [10:0] buffer_3_694; // @[Modules.scala 56:109:@14610.4]
  wire [11:0] _T_66626; // @[Modules.scala 56:109:@14612.4]
  wire [10:0] _T_66627; // @[Modules.scala 56:109:@14613.4]
  wire [10:0] buffer_3_695; // @[Modules.scala 56:109:@14614.4]
  wire [11:0] _T_66629; // @[Modules.scala 56:109:@14616.4]
  wire [10:0] _T_66630; // @[Modules.scala 56:109:@14617.4]
  wire [10:0] buffer_3_696; // @[Modules.scala 56:109:@14618.4]
  wire [11:0] _T_66632; // @[Modules.scala 56:109:@14620.4]
  wire [10:0] _T_66633; // @[Modules.scala 56:109:@14621.4]
  wire [10:0] buffer_3_697; // @[Modules.scala 56:109:@14622.4]
  wire [11:0] _T_66635; // @[Modules.scala 56:109:@14624.4]
  wire [10:0] _T_66636; // @[Modules.scala 56:109:@14625.4]
  wire [10:0] buffer_3_698; // @[Modules.scala 56:109:@14626.4]
  wire [11:0] _T_66638; // @[Modules.scala 56:109:@14628.4]
  wire [10:0] _T_66639; // @[Modules.scala 56:109:@14629.4]
  wire [10:0] buffer_3_699; // @[Modules.scala 56:109:@14630.4]
  wire [11:0] _T_66641; // @[Modules.scala 56:109:@14632.4]
  wire [10:0] _T_66642; // @[Modules.scala 56:109:@14633.4]
  wire [10:0] buffer_3_700; // @[Modules.scala 56:109:@14634.4]
  wire [11:0] _T_66644; // @[Modules.scala 56:109:@14636.4]
  wire [10:0] _T_66645; // @[Modules.scala 56:109:@14637.4]
  wire [10:0] buffer_3_701; // @[Modules.scala 56:109:@14638.4]
  wire [11:0] _T_66647; // @[Modules.scala 56:109:@14640.4]
  wire [10:0] _T_66648; // @[Modules.scala 56:109:@14641.4]
  wire [10:0] buffer_3_702; // @[Modules.scala 56:109:@14642.4]
  wire [11:0] _T_66650; // @[Modules.scala 56:109:@14644.4]
  wire [10:0] _T_66651; // @[Modules.scala 56:109:@14645.4]
  wire [10:0] buffer_3_703; // @[Modules.scala 56:109:@14646.4]
  wire [11:0] _T_66653; // @[Modules.scala 56:109:@14648.4]
  wire [10:0] _T_66654; // @[Modules.scala 56:109:@14649.4]
  wire [10:0] buffer_3_704; // @[Modules.scala 56:109:@14650.4]
  wire [11:0] _T_66656; // @[Modules.scala 56:109:@14652.4]
  wire [10:0] _T_66657; // @[Modules.scala 56:109:@14653.4]
  wire [10:0] buffer_3_705; // @[Modules.scala 56:109:@14654.4]
  wire [11:0] _T_66659; // @[Modules.scala 56:109:@14656.4]
  wire [10:0] _T_66660; // @[Modules.scala 56:109:@14657.4]
  wire [10:0] buffer_3_706; // @[Modules.scala 56:109:@14658.4]
  wire [11:0] _T_66662; // @[Modules.scala 56:109:@14660.4]
  wire [10:0] _T_66663; // @[Modules.scala 56:109:@14661.4]
  wire [10:0] buffer_3_707; // @[Modules.scala 56:109:@14662.4]
  wire [11:0] _T_66665; // @[Modules.scala 56:109:@14664.4]
  wire [10:0] _T_66666; // @[Modules.scala 56:109:@14665.4]
  wire [10:0] buffer_3_708; // @[Modules.scala 56:109:@14666.4]
  wire [11:0] _T_66668; // @[Modules.scala 56:109:@14668.4]
  wire [10:0] _T_66669; // @[Modules.scala 56:109:@14669.4]
  wire [10:0] buffer_3_709; // @[Modules.scala 56:109:@14670.4]
  wire [11:0] _T_66671; // @[Modules.scala 56:109:@14672.4]
  wire [10:0] _T_66672; // @[Modules.scala 56:109:@14673.4]
  wire [10:0] buffer_3_710; // @[Modules.scala 56:109:@14674.4]
  wire [11:0] _T_66674; // @[Modules.scala 56:109:@14676.4]
  wire [10:0] _T_66675; // @[Modules.scala 56:109:@14677.4]
  wire [10:0] buffer_3_711; // @[Modules.scala 56:109:@14678.4]
  wire [11:0] _T_66677; // @[Modules.scala 56:109:@14680.4]
  wire [10:0] _T_66678; // @[Modules.scala 56:109:@14681.4]
  wire [10:0] buffer_3_712; // @[Modules.scala 56:109:@14682.4]
  wire [11:0] _T_66680; // @[Modules.scala 56:109:@14684.4]
  wire [10:0] _T_66681; // @[Modules.scala 56:109:@14685.4]
  wire [10:0] buffer_3_713; // @[Modules.scala 56:109:@14686.4]
  wire [11:0] _T_66683; // @[Modules.scala 56:109:@14688.4]
  wire [10:0] _T_66684; // @[Modules.scala 56:109:@14689.4]
  wire [10:0] buffer_3_714; // @[Modules.scala 56:109:@14690.4]
  wire [11:0] _T_66686; // @[Modules.scala 56:109:@14692.4]
  wire [10:0] _T_66687; // @[Modules.scala 56:109:@14693.4]
  wire [10:0] buffer_3_715; // @[Modules.scala 56:109:@14694.4]
  wire [11:0] _T_66689; // @[Modules.scala 56:109:@14696.4]
  wire [10:0] _T_66690; // @[Modules.scala 56:109:@14697.4]
  wire [10:0] buffer_3_716; // @[Modules.scala 56:109:@14698.4]
  wire [11:0] _T_66692; // @[Modules.scala 56:109:@14700.4]
  wire [10:0] _T_66693; // @[Modules.scala 56:109:@14701.4]
  wire [10:0] buffer_3_717; // @[Modules.scala 56:109:@14702.4]
  wire [11:0] _T_66695; // @[Modules.scala 56:109:@14704.4]
  wire [10:0] _T_66696; // @[Modules.scala 56:109:@14705.4]
  wire [10:0] buffer_3_718; // @[Modules.scala 56:109:@14706.4]
  wire [11:0] _T_66698; // @[Modules.scala 56:109:@14708.4]
  wire [10:0] _T_66699; // @[Modules.scala 56:109:@14709.4]
  wire [10:0] buffer_3_719; // @[Modules.scala 56:109:@14710.4]
  wire [11:0] _T_66701; // @[Modules.scala 56:109:@14712.4]
  wire [10:0] _T_66702; // @[Modules.scala 56:109:@14713.4]
  wire [10:0] buffer_3_720; // @[Modules.scala 56:109:@14714.4]
  wire [11:0] _T_66704; // @[Modules.scala 56:109:@14716.4]
  wire [10:0] _T_66705; // @[Modules.scala 56:109:@14717.4]
  wire [10:0] buffer_3_721; // @[Modules.scala 56:109:@14718.4]
  wire [11:0] _T_66707; // @[Modules.scala 56:109:@14720.4]
  wire [10:0] _T_66708; // @[Modules.scala 56:109:@14721.4]
  wire [10:0] buffer_3_722; // @[Modules.scala 56:109:@14722.4]
  wire [11:0] _T_66710; // @[Modules.scala 56:109:@14724.4]
  wire [10:0] _T_66711; // @[Modules.scala 56:109:@14725.4]
  wire [10:0] buffer_3_723; // @[Modules.scala 56:109:@14726.4]
  wire [11:0] _T_66713; // @[Modules.scala 56:109:@14728.4]
  wire [10:0] _T_66714; // @[Modules.scala 56:109:@14729.4]
  wire [10:0] buffer_3_724; // @[Modules.scala 56:109:@14730.4]
  wire [11:0] _T_66716; // @[Modules.scala 56:109:@14732.4]
  wire [10:0] _T_66717; // @[Modules.scala 56:109:@14733.4]
  wire [10:0] buffer_3_725; // @[Modules.scala 56:109:@14734.4]
  wire [11:0] _T_66719; // @[Modules.scala 56:109:@14736.4]
  wire [10:0] _T_66720; // @[Modules.scala 56:109:@14737.4]
  wire [10:0] buffer_3_726; // @[Modules.scala 56:109:@14738.4]
  wire [11:0] _T_66722; // @[Modules.scala 56:109:@14740.4]
  wire [10:0] _T_66723; // @[Modules.scala 56:109:@14741.4]
  wire [10:0] buffer_3_727; // @[Modules.scala 56:109:@14742.4]
  wire [11:0] _T_66725; // @[Modules.scala 56:109:@14744.4]
  wire [10:0] _T_66726; // @[Modules.scala 56:109:@14745.4]
  wire [10:0] buffer_3_728; // @[Modules.scala 56:109:@14746.4]
  wire [11:0] _T_66728; // @[Modules.scala 56:109:@14748.4]
  wire [10:0] _T_66729; // @[Modules.scala 56:109:@14749.4]
  wire [10:0] buffer_3_729; // @[Modules.scala 56:109:@14750.4]
  wire [11:0] _T_66731; // @[Modules.scala 56:109:@14752.4]
  wire [10:0] _T_66732; // @[Modules.scala 56:109:@14753.4]
  wire [10:0] buffer_3_730; // @[Modules.scala 56:109:@14754.4]
  wire [11:0] _T_66734; // @[Modules.scala 56:109:@14756.4]
  wire [10:0] _T_66735; // @[Modules.scala 56:109:@14757.4]
  wire [10:0] buffer_3_731; // @[Modules.scala 56:109:@14758.4]
  wire [11:0] _T_66737; // @[Modules.scala 56:109:@14760.4]
  wire [10:0] _T_66738; // @[Modules.scala 56:109:@14761.4]
  wire [10:0] buffer_3_732; // @[Modules.scala 56:109:@14762.4]
  wire [11:0] _T_66740; // @[Modules.scala 56:109:@14764.4]
  wire [10:0] _T_66741; // @[Modules.scala 56:109:@14765.4]
  wire [10:0] buffer_3_733; // @[Modules.scala 56:109:@14766.4]
  wire [11:0] _T_66743; // @[Modules.scala 56:109:@14768.4]
  wire [10:0] _T_66744; // @[Modules.scala 56:109:@14769.4]
  wire [10:0] buffer_3_734; // @[Modules.scala 56:109:@14770.4]
  wire [11:0] _T_66746; // @[Modules.scala 63:156:@14773.4]
  wire [10:0] _T_66747; // @[Modules.scala 63:156:@14774.4]
  wire [10:0] buffer_3_736; // @[Modules.scala 63:156:@14775.4]
  wire [11:0] _T_66749; // @[Modules.scala 63:156:@14777.4]
  wire [10:0] _T_66750; // @[Modules.scala 63:156:@14778.4]
  wire [10:0] buffer_3_737; // @[Modules.scala 63:156:@14779.4]
  wire [11:0] _T_66752; // @[Modules.scala 63:156:@14781.4]
  wire [10:0] _T_66753; // @[Modules.scala 63:156:@14782.4]
  wire [10:0] buffer_3_738; // @[Modules.scala 63:156:@14783.4]
  wire [11:0] _T_66755; // @[Modules.scala 63:156:@14785.4]
  wire [10:0] _T_66756; // @[Modules.scala 63:156:@14786.4]
  wire [10:0] buffer_3_739; // @[Modules.scala 63:156:@14787.4]
  wire [11:0] _T_66758; // @[Modules.scala 63:156:@14789.4]
  wire [10:0] _T_66759; // @[Modules.scala 63:156:@14790.4]
  wire [10:0] buffer_3_740; // @[Modules.scala 63:156:@14791.4]
  wire [11:0] _T_66761; // @[Modules.scala 63:156:@14793.4]
  wire [10:0] _T_66762; // @[Modules.scala 63:156:@14794.4]
  wire [10:0] buffer_3_741; // @[Modules.scala 63:156:@14795.4]
  wire [11:0] _T_66764; // @[Modules.scala 63:156:@14797.4]
  wire [10:0] _T_66765; // @[Modules.scala 63:156:@14798.4]
  wire [10:0] buffer_3_742; // @[Modules.scala 63:156:@14799.4]
  wire [11:0] _T_66767; // @[Modules.scala 63:156:@14801.4]
  wire [10:0] _T_66768; // @[Modules.scala 63:156:@14802.4]
  wire [10:0] buffer_3_743; // @[Modules.scala 63:156:@14803.4]
  wire [11:0] _T_66770; // @[Modules.scala 63:156:@14805.4]
  wire [10:0] _T_66771; // @[Modules.scala 63:156:@14806.4]
  wire [10:0] buffer_3_744; // @[Modules.scala 63:156:@14807.4]
  wire [11:0] _T_66773; // @[Modules.scala 63:156:@14809.4]
  wire [10:0] _T_66774; // @[Modules.scala 63:156:@14810.4]
  wire [10:0] buffer_3_745; // @[Modules.scala 63:156:@14811.4]
  wire [11:0] _T_66776; // @[Modules.scala 63:156:@14813.4]
  wire [10:0] _T_66777; // @[Modules.scala 63:156:@14814.4]
  wire [10:0] buffer_3_746; // @[Modules.scala 63:156:@14815.4]
  wire [11:0] _T_66779; // @[Modules.scala 63:156:@14817.4]
  wire [10:0] _T_66780; // @[Modules.scala 63:156:@14818.4]
  wire [10:0] buffer_3_747; // @[Modules.scala 63:156:@14819.4]
  wire [11:0] _T_66782; // @[Modules.scala 63:156:@14821.4]
  wire [10:0] _T_66783; // @[Modules.scala 63:156:@14822.4]
  wire [10:0] buffer_3_748; // @[Modules.scala 63:156:@14823.4]
  wire [11:0] _T_66785; // @[Modules.scala 63:156:@14825.4]
  wire [10:0] _T_66786; // @[Modules.scala 63:156:@14826.4]
  wire [10:0] buffer_3_749; // @[Modules.scala 63:156:@14827.4]
  wire [11:0] _T_66788; // @[Modules.scala 63:156:@14829.4]
  wire [10:0] _T_66789; // @[Modules.scala 63:156:@14830.4]
  wire [10:0] buffer_3_750; // @[Modules.scala 63:156:@14831.4]
  wire [11:0] _T_66791; // @[Modules.scala 63:156:@14833.4]
  wire [10:0] _T_66792; // @[Modules.scala 63:156:@14834.4]
  wire [10:0] buffer_3_751; // @[Modules.scala 63:156:@14835.4]
  wire [11:0] _T_66794; // @[Modules.scala 63:156:@14837.4]
  wire [10:0] _T_66795; // @[Modules.scala 63:156:@14838.4]
  wire [10:0] buffer_3_752; // @[Modules.scala 63:156:@14839.4]
  wire [11:0] _T_66797; // @[Modules.scala 63:156:@14841.4]
  wire [10:0] _T_66798; // @[Modules.scala 63:156:@14842.4]
  wire [10:0] buffer_3_753; // @[Modules.scala 63:156:@14843.4]
  wire [11:0] _T_66800; // @[Modules.scala 63:156:@14845.4]
  wire [10:0] _T_66801; // @[Modules.scala 63:156:@14846.4]
  wire [10:0] buffer_3_754; // @[Modules.scala 63:156:@14847.4]
  wire [11:0] _T_66803; // @[Modules.scala 63:156:@14849.4]
  wire [10:0] _T_66804; // @[Modules.scala 63:156:@14850.4]
  wire [10:0] buffer_3_755; // @[Modules.scala 63:156:@14851.4]
  wire [11:0] _T_66806; // @[Modules.scala 63:156:@14853.4]
  wire [10:0] _T_66807; // @[Modules.scala 63:156:@14854.4]
  wire [10:0] buffer_3_756; // @[Modules.scala 63:156:@14855.4]
  wire [11:0] _T_66809; // @[Modules.scala 63:156:@14857.4]
  wire [10:0] _T_66810; // @[Modules.scala 63:156:@14858.4]
  wire [10:0] buffer_3_757; // @[Modules.scala 63:156:@14859.4]
  wire [11:0] _T_66812; // @[Modules.scala 63:156:@14861.4]
  wire [10:0] _T_66813; // @[Modules.scala 63:156:@14862.4]
  wire [10:0] buffer_3_758; // @[Modules.scala 63:156:@14863.4]
  wire [11:0] _T_66815; // @[Modules.scala 63:156:@14865.4]
  wire [10:0] _T_66816; // @[Modules.scala 63:156:@14866.4]
  wire [10:0] buffer_3_759; // @[Modules.scala 63:156:@14867.4]
  wire [11:0] _T_66818; // @[Modules.scala 63:156:@14869.4]
  wire [10:0] _T_66819; // @[Modules.scala 63:156:@14870.4]
  wire [10:0] buffer_3_760; // @[Modules.scala 63:156:@14871.4]
  wire [11:0] _T_66821; // @[Modules.scala 63:156:@14873.4]
  wire [10:0] _T_66822; // @[Modules.scala 63:156:@14874.4]
  wire [10:0] buffer_3_761; // @[Modules.scala 63:156:@14875.4]
  wire [11:0] _T_66824; // @[Modules.scala 63:156:@14877.4]
  wire [10:0] _T_66825; // @[Modules.scala 63:156:@14878.4]
  wire [10:0] buffer_3_762; // @[Modules.scala 63:156:@14879.4]
  wire [11:0] _T_66827; // @[Modules.scala 63:156:@14881.4]
  wire [10:0] _T_66828; // @[Modules.scala 63:156:@14882.4]
  wire [10:0] buffer_3_763; // @[Modules.scala 63:156:@14883.4]
  wire [11:0] _T_66830; // @[Modules.scala 63:156:@14885.4]
  wire [10:0] _T_66831; // @[Modules.scala 63:156:@14886.4]
  wire [10:0] buffer_3_764; // @[Modules.scala 63:156:@14887.4]
  wire [11:0] _T_66833; // @[Modules.scala 63:156:@14889.4]
  wire [10:0] _T_66834; // @[Modules.scala 63:156:@14890.4]
  wire [10:0] buffer_3_765; // @[Modules.scala 63:156:@14891.4]
  wire [11:0] _T_66836; // @[Modules.scala 63:156:@14893.4]
  wire [10:0] _T_66837; // @[Modules.scala 63:156:@14894.4]
  wire [10:0] buffer_3_766; // @[Modules.scala 63:156:@14895.4]
  wire [11:0] _T_66839; // @[Modules.scala 63:156:@14897.4]
  wire [10:0] _T_66840; // @[Modules.scala 63:156:@14898.4]
  wire [10:0] buffer_3_767; // @[Modules.scala 63:156:@14899.4]
  wire [11:0] _T_66842; // @[Modules.scala 63:156:@14901.4]
  wire [10:0] _T_66843; // @[Modules.scala 63:156:@14902.4]
  wire [10:0] buffer_3_768; // @[Modules.scala 63:156:@14903.4]
  wire [11:0] _T_66845; // @[Modules.scala 63:156:@14905.4]
  wire [10:0] _T_66846; // @[Modules.scala 63:156:@14906.4]
  wire [10:0] buffer_3_769; // @[Modules.scala 63:156:@14907.4]
  wire [11:0] _T_66848; // @[Modules.scala 63:156:@14909.4]
  wire [10:0] _T_66849; // @[Modules.scala 63:156:@14910.4]
  wire [10:0] buffer_3_770; // @[Modules.scala 63:156:@14911.4]
  wire [11:0] _T_66851; // @[Modules.scala 63:156:@14913.4]
  wire [10:0] _T_66852; // @[Modules.scala 63:156:@14914.4]
  wire [10:0] buffer_3_771; // @[Modules.scala 63:156:@14915.4]
  wire [11:0] _T_66854; // @[Modules.scala 63:156:@14917.4]
  wire [10:0] _T_66855; // @[Modules.scala 63:156:@14918.4]
  wire [10:0] buffer_3_772; // @[Modules.scala 63:156:@14919.4]
  wire [11:0] _T_66857; // @[Modules.scala 63:156:@14921.4]
  wire [10:0] _T_66858; // @[Modules.scala 63:156:@14922.4]
  wire [10:0] buffer_3_773; // @[Modules.scala 63:156:@14923.4]
  wire [11:0] _T_66860; // @[Modules.scala 63:156:@14925.4]
  wire [10:0] _T_66861; // @[Modules.scala 63:156:@14926.4]
  wire [10:0] buffer_3_774; // @[Modules.scala 63:156:@14927.4]
  wire [11:0] _T_66863; // @[Modules.scala 63:156:@14929.4]
  wire [10:0] _T_66864; // @[Modules.scala 63:156:@14930.4]
  wire [10:0] buffer_3_775; // @[Modules.scala 63:156:@14931.4]
  wire [11:0] _T_66866; // @[Modules.scala 63:156:@14933.4]
  wire [10:0] _T_66867; // @[Modules.scala 63:156:@14934.4]
  wire [10:0] buffer_3_776; // @[Modules.scala 63:156:@14935.4]
  wire [11:0] _T_66869; // @[Modules.scala 63:156:@14937.4]
  wire [10:0] _T_66870; // @[Modules.scala 63:156:@14938.4]
  wire [10:0] buffer_3_777; // @[Modules.scala 63:156:@14939.4]
  wire [11:0] _T_66872; // @[Modules.scala 63:156:@14941.4]
  wire [10:0] _T_66873; // @[Modules.scala 63:156:@14942.4]
  wire [10:0] buffer_3_778; // @[Modules.scala 63:156:@14943.4]
  wire [11:0] _T_66875; // @[Modules.scala 63:156:@14945.4]
  wire [10:0] _T_66876; // @[Modules.scala 63:156:@14946.4]
  wire [10:0] buffer_3_779; // @[Modules.scala 63:156:@14947.4]
  wire [11:0] _T_66878; // @[Modules.scala 63:156:@14949.4]
  wire [10:0] _T_66879; // @[Modules.scala 63:156:@14950.4]
  wire [10:0] buffer_3_780; // @[Modules.scala 63:156:@14951.4]
  wire [11:0] _T_66881; // @[Modules.scala 63:156:@14953.4]
  wire [10:0] _T_66882; // @[Modules.scala 63:156:@14954.4]
  wire [10:0] buffer_3_781; // @[Modules.scala 63:156:@14955.4]
  wire [11:0] _T_66884; // @[Modules.scala 63:156:@14957.4]
  wire [10:0] _T_66885; // @[Modules.scala 63:156:@14958.4]
  wire [10:0] buffer_3_782; // @[Modules.scala 63:156:@14959.4]
  wire [11:0] _T_66887; // @[Modules.scala 63:156:@14961.4]
  wire [10:0] _T_66888; // @[Modules.scala 63:156:@14962.4]
  wire [10:0] buffer_3_783; // @[Modules.scala 63:156:@14963.4]
  wire [5:0] _T_66897; // @[Modules.scala 43:47:@14973.4]
  wire [4:0] _T_66898; // @[Modules.scala 43:47:@14974.4]
  wire [4:0] _T_66899; // @[Modules.scala 43:47:@14975.4]
  wire [5:0] _T_66921; // @[Modules.scala 43:47:@14998.4]
  wire [4:0] _T_66922; // @[Modules.scala 43:47:@14999.4]
  wire [4:0] _T_66923; // @[Modules.scala 43:47:@15000.4]
  wire [5:0] _T_66935; // @[Modules.scala 46:37:@15013.4]
  wire [4:0] _T_66936; // @[Modules.scala 46:37:@15014.4]
  wire [4:0] _T_66937; // @[Modules.scala 46:37:@15015.4]
  wire [5:0] _T_66938; // @[Modules.scala 46:47:@15016.4]
  wire [4:0] _T_66939; // @[Modules.scala 46:47:@15017.4]
  wire [4:0] _T_66940; // @[Modules.scala 46:47:@15018.4]
  wire [5:0] _T_66951; // @[Modules.scala 46:47:@15031.4]
  wire [4:0] _T_66952; // @[Modules.scala 46:47:@15032.4]
  wire [4:0] _T_66953; // @[Modules.scala 46:47:@15033.4]
  wire [5:0] _T_66961; // @[Modules.scala 43:47:@15042.4]
  wire [4:0] _T_66962; // @[Modules.scala 43:47:@15043.4]
  wire [4:0] _T_66963; // @[Modules.scala 43:47:@15044.4]
  wire [5:0] _T_66968; // @[Modules.scala 43:47:@15049.4]
  wire [4:0] _T_66969; // @[Modules.scala 43:47:@15050.4]
  wire [4:0] _T_66970; // @[Modules.scala 43:47:@15051.4]
  wire [5:0] _T_67000; // @[Modules.scala 37:46:@15087.4]
  wire [4:0] _T_67001; // @[Modules.scala 37:46:@15088.4]
  wire [4:0] _T_67002; // @[Modules.scala 37:46:@15089.4]
  wire [5:0] _T_67102; // @[Modules.scala 43:47:@15202.4]
  wire [4:0] _T_67103; // @[Modules.scala 43:47:@15203.4]
  wire [4:0] _T_67104; // @[Modules.scala 43:47:@15204.4]
  wire [5:0] _T_67156; // @[Modules.scala 43:47:@15267.4]
  wire [4:0] _T_67157; // @[Modules.scala 43:47:@15268.4]
  wire [4:0] _T_67158; // @[Modules.scala 43:47:@15269.4]
  wire [5:0] _T_67163; // @[Modules.scala 43:47:@15274.4]
  wire [4:0] _T_67164; // @[Modules.scala 43:47:@15275.4]
  wire [4:0] _T_67165; // @[Modules.scala 43:47:@15276.4]
  wire [5:0] _T_67169; // @[Modules.scala 40:46:@15282.4]
  wire [4:0] _T_67170; // @[Modules.scala 40:46:@15283.4]
  wire [4:0] _T_67171; // @[Modules.scala 40:46:@15284.4]
  wire [5:0] _T_67182; // @[Modules.scala 40:46:@15297.4]
  wire [4:0] _T_67183; // @[Modules.scala 40:46:@15298.4]
  wire [4:0] _T_67184; // @[Modules.scala 40:46:@15299.4]
  wire [5:0] _T_67200; // @[Modules.scala 46:37:@15315.4]
  wire [4:0] _T_67201; // @[Modules.scala 46:37:@15316.4]
  wire [4:0] _T_67202; // @[Modules.scala 46:37:@15317.4]
  wire [5:0] _T_67203; // @[Modules.scala 46:47:@15318.4]
  wire [4:0] _T_67204; // @[Modules.scala 46:47:@15319.4]
  wire [4:0] _T_67205; // @[Modules.scala 46:47:@15320.4]
  wire [5:0] _T_67209; // @[Modules.scala 37:46:@15326.4]
  wire [4:0] _T_67210; // @[Modules.scala 37:46:@15327.4]
  wire [4:0] _T_67211; // @[Modules.scala 37:46:@15328.4]
  wire [5:0] _T_67226; // @[Modules.scala 37:46:@15344.4]
  wire [4:0] _T_67227; // @[Modules.scala 37:46:@15345.4]
  wire [4:0] _T_67228; // @[Modules.scala 37:46:@15346.4]
  wire [5:0] _T_67238; // @[Modules.scala 37:46:@15360.4]
  wire [4:0] _T_67239; // @[Modules.scala 37:46:@15361.4]
  wire [4:0] _T_67240; // @[Modules.scala 37:46:@15362.4]
  wire [5:0] _T_67244; // @[Modules.scala 37:46:@15368.4]
  wire [4:0] _T_67245; // @[Modules.scala 37:46:@15369.4]
  wire [4:0] _T_67246; // @[Modules.scala 37:46:@15370.4]
  wire [5:0] _T_67250; // @[Modules.scala 40:46:@15376.4]
  wire [4:0] _T_67251; // @[Modules.scala 40:46:@15377.4]
  wire [4:0] _T_67252; // @[Modules.scala 40:46:@15378.4]
  wire [5:0] _T_67266; // @[Modules.scala 37:46:@15395.4]
  wire [4:0] _T_67267; // @[Modules.scala 37:46:@15396.4]
  wire [4:0] _T_67268; // @[Modules.scala 37:46:@15397.4]
  wire [5:0] _T_67306; // @[Modules.scala 43:47:@15439.4]
  wire [4:0] _T_67307; // @[Modules.scala 43:47:@15440.4]
  wire [4:0] _T_67308; // @[Modules.scala 43:47:@15441.4]
  wire [5:0] _T_67312; // @[Modules.scala 37:46:@15447.4]
  wire [4:0] _T_67313; // @[Modules.scala 37:46:@15448.4]
  wire [4:0] _T_67314; // @[Modules.scala 37:46:@15449.4]
  wire [5:0] _T_67345; // @[Modules.scala 43:47:@15484.4]
  wire [4:0] _T_67346; // @[Modules.scala 43:47:@15485.4]
  wire [4:0] _T_67347; // @[Modules.scala 43:47:@15486.4]
  wire [5:0] _T_67348; // @[Modules.scala 40:46:@15488.4]
  wire [4:0] _T_67349; // @[Modules.scala 40:46:@15489.4]
  wire [4:0] _T_67350; // @[Modules.scala 40:46:@15490.4]
  wire [5:0] _T_67362; // @[Modules.scala 46:37:@15503.4]
  wire [4:0] _T_67363; // @[Modules.scala 46:37:@15504.4]
  wire [4:0] _T_67364; // @[Modules.scala 46:37:@15505.4]
  wire [5:0] _T_67365; // @[Modules.scala 46:47:@15506.4]
  wire [4:0] _T_67366; // @[Modules.scala 46:47:@15507.4]
  wire [4:0] _T_67367; // @[Modules.scala 46:47:@15508.4]
  wire [5:0] _T_67372; // @[Modules.scala 46:47:@15513.4]
  wire [4:0] _T_67373; // @[Modules.scala 46:47:@15514.4]
  wire [4:0] _T_67374; // @[Modules.scala 46:47:@15515.4]
  wire [5:0] _T_67412; // @[Modules.scala 43:47:@15557.4]
  wire [4:0] _T_67413; // @[Modules.scala 43:47:@15558.4]
  wire [4:0] _T_67414; // @[Modules.scala 43:47:@15559.4]
  wire [5:0] _T_67422; // @[Modules.scala 37:46:@15568.4]
  wire [4:0] _T_67423; // @[Modules.scala 37:46:@15569.4]
  wire [4:0] _T_67424; // @[Modules.scala 37:46:@15570.4]
  wire [5:0] _T_67453; // @[Modules.scala 43:47:@15600.4]
  wire [4:0] _T_67454; // @[Modules.scala 43:47:@15601.4]
  wire [4:0] _T_67455; // @[Modules.scala 43:47:@15602.4]
  wire [5:0] _T_67456; // @[Modules.scala 37:46:@15604.4]
  wire [4:0] _T_67457; // @[Modules.scala 37:46:@15605.4]
  wire [4:0] _T_67458; // @[Modules.scala 37:46:@15606.4]
  wire [5:0] _T_67486; // @[Modules.scala 43:47:@15637.4]
  wire [4:0] _T_67487; // @[Modules.scala 43:47:@15638.4]
  wire [4:0] _T_67488; // @[Modules.scala 43:47:@15639.4]
  wire [5:0] _T_67489; // @[Modules.scala 37:46:@15641.4]
  wire [4:0] _T_67490; // @[Modules.scala 37:46:@15642.4]
  wire [4:0] _T_67491; // @[Modules.scala 37:46:@15643.4]
  wire [5:0] _T_67492; // @[Modules.scala 37:46:@15645.4]
  wire [4:0] _T_67493; // @[Modules.scala 37:46:@15646.4]
  wire [4:0] _T_67494; // @[Modules.scala 37:46:@15647.4]
  wire [5:0] _T_67594; // @[Modules.scala 43:47:@15753.4]
  wire [4:0] _T_67595; // @[Modules.scala 43:47:@15754.4]
  wire [4:0] _T_67596; // @[Modules.scala 43:47:@15755.4]
  wire [5:0] _T_67597; // @[Modules.scala 37:46:@15757.4]
  wire [4:0] _T_67598; // @[Modules.scala 37:46:@15758.4]
  wire [4:0] _T_67599; // @[Modules.scala 37:46:@15759.4]
  wire [5:0] _T_67607; // @[Modules.scala 37:46:@15768.4]
  wire [4:0] _T_67608; // @[Modules.scala 37:46:@15769.4]
  wire [4:0] _T_67609; // @[Modules.scala 37:46:@15770.4]
  wire [5:0] _T_67616; // @[Modules.scala 40:46:@15780.4]
  wire [4:0] _T_67617; // @[Modules.scala 40:46:@15781.4]
  wire [4:0] _T_67618; // @[Modules.scala 40:46:@15782.4]
  wire [5:0] _T_67623; // @[Modules.scala 43:47:@15787.4]
  wire [4:0] _T_67624; // @[Modules.scala 43:47:@15788.4]
  wire [4:0] _T_67625; // @[Modules.scala 43:47:@15789.4]
  wire [5:0] _T_67718; // @[Modules.scala 40:46:@15888.4]
  wire [4:0] _T_67719; // @[Modules.scala 40:46:@15889.4]
  wire [4:0] _T_67720; // @[Modules.scala 40:46:@15890.4]
  wire [5:0] _T_67734; // @[Modules.scala 40:46:@15907.4]
  wire [4:0] _T_67735; // @[Modules.scala 40:46:@15908.4]
  wire [4:0] _T_67736; // @[Modules.scala 40:46:@15909.4]
  wire [5:0] _T_67764; // @[Modules.scala 40:46:@15940.4]
  wire [4:0] _T_67765; // @[Modules.scala 40:46:@15941.4]
  wire [4:0] _T_67766; // @[Modules.scala 40:46:@15942.4]
  wire [5:0] _T_67781; // @[Modules.scala 40:46:@15958.4]
  wire [4:0] _T_67782; // @[Modules.scala 40:46:@15959.4]
  wire [4:0] _T_67783; // @[Modules.scala 40:46:@15960.4]
  wire [5:0] _T_67800; // @[Modules.scala 40:46:@15981.4]
  wire [4:0] _T_67801; // @[Modules.scala 40:46:@15982.4]
  wire [4:0] _T_67802; // @[Modules.scala 40:46:@15983.4]
  wire [5:0] _T_67820; // @[Modules.scala 37:46:@16003.4]
  wire [4:0] _T_67821; // @[Modules.scala 37:46:@16004.4]
  wire [4:0] _T_67822; // @[Modules.scala 37:46:@16005.4]
  wire [5:0] _T_67823; // @[Modules.scala 40:46:@16007.4]
  wire [4:0] _T_67824; // @[Modules.scala 40:46:@16008.4]
  wire [4:0] _T_67825; // @[Modules.scala 40:46:@16009.4]
  wire [5:0] _T_67826; // @[Modules.scala 40:46:@16011.4]
  wire [4:0] _T_67827; // @[Modules.scala 40:46:@16012.4]
  wire [4:0] _T_67828; // @[Modules.scala 40:46:@16013.4]
  wire [5:0] _T_67847; // @[Modules.scala 43:47:@16032.4]
  wire [4:0] _T_67848; // @[Modules.scala 43:47:@16033.4]
  wire [4:0] _T_67849; // @[Modules.scala 43:47:@16034.4]
  wire [5:0] _T_67867; // @[Modules.scala 43:47:@16054.4]
  wire [4:0] _T_67868; // @[Modules.scala 43:47:@16055.4]
  wire [4:0] _T_67869; // @[Modules.scala 43:47:@16056.4]
  wire [5:0] _T_67876; // @[Modules.scala 40:46:@16066.4]
  wire [4:0] _T_67877; // @[Modules.scala 40:46:@16067.4]
  wire [4:0] _T_67878; // @[Modules.scala 40:46:@16068.4]
  wire [5:0] _T_67882; // @[Modules.scala 37:46:@16074.4]
  wire [4:0] _T_67883; // @[Modules.scala 37:46:@16075.4]
  wire [4:0] _T_67884; // @[Modules.scala 37:46:@16076.4]
  wire [5:0] _T_67885; // @[Modules.scala 40:46:@16078.4]
  wire [4:0] _T_67886; // @[Modules.scala 40:46:@16079.4]
  wire [4:0] _T_67887; // @[Modules.scala 40:46:@16080.4]
  wire [5:0] _T_67888; // @[Modules.scala 37:46:@16082.4]
  wire [4:0] _T_67889; // @[Modules.scala 37:46:@16083.4]
  wire [4:0] _T_67890; // @[Modules.scala 37:46:@16084.4]
  wire [5:0] _T_67910; // @[Modules.scala 40:46:@16109.4]
  wire [4:0] _T_67911; // @[Modules.scala 40:46:@16110.4]
  wire [4:0] _T_67912; // @[Modules.scala 40:46:@16111.4]
  wire [5:0] _T_67916; // @[Modules.scala 40:46:@16117.4]
  wire [4:0] _T_67917; // @[Modules.scala 40:46:@16118.4]
  wire [4:0] _T_67918; // @[Modules.scala 40:46:@16119.4]
  wire [5:0] _T_67959; // @[Modules.scala 40:46:@16165.4]
  wire [4:0] _T_67960; // @[Modules.scala 40:46:@16166.4]
  wire [4:0] _T_67961; // @[Modules.scala 40:46:@16167.4]
  wire [5:0] _T_67979; // @[Modules.scala 43:47:@16187.4]
  wire [4:0] _T_67980; // @[Modules.scala 43:47:@16188.4]
  wire [4:0] _T_67981; // @[Modules.scala 43:47:@16189.4]
  wire [5:0] _T_68027; // @[Modules.scala 43:47:@16244.4]
  wire [4:0] _T_68028; // @[Modules.scala 43:47:@16245.4]
  wire [4:0] _T_68029; // @[Modules.scala 43:47:@16246.4]
  wire [5:0] _T_68044; // @[Modules.scala 37:46:@16262.4]
  wire [4:0] _T_68045; // @[Modules.scala 37:46:@16263.4]
  wire [4:0] _T_68046; // @[Modules.scala 37:46:@16264.4]
  wire [5:0] _T_68048; // @[Modules.scala 43:37:@16266.4]
  wire [4:0] _T_68049; // @[Modules.scala 43:37:@16267.4]
  wire [4:0] _T_68050; // @[Modules.scala 43:37:@16268.4]
  wire [5:0] _T_68051; // @[Modules.scala 43:47:@16269.4]
  wire [4:0] _T_68052; // @[Modules.scala 43:47:@16270.4]
  wire [4:0] _T_68053; // @[Modules.scala 43:47:@16271.4]
  wire [5:0] _T_68082; // @[Modules.scala 40:46:@16308.4]
  wire [4:0] _T_68083; // @[Modules.scala 40:46:@16309.4]
  wire [4:0] _T_68084; // @[Modules.scala 40:46:@16310.4]
  wire [5:0] _T_68085; // @[Modules.scala 40:46:@16312.4]
  wire [4:0] _T_68086; // @[Modules.scala 40:46:@16313.4]
  wire [4:0] _T_68087; // @[Modules.scala 40:46:@16314.4]
  wire [5:0] _T_68095; // @[Modules.scala 43:47:@16323.4]
  wire [4:0] _T_68096; // @[Modules.scala 43:47:@16324.4]
  wire [4:0] _T_68097; // @[Modules.scala 43:47:@16325.4]
  wire [5:0] _T_68098; // @[Modules.scala 40:46:@16327.4]
  wire [4:0] _T_68099; // @[Modules.scala 40:46:@16328.4]
  wire [4:0] _T_68100; // @[Modules.scala 40:46:@16329.4]
  wire [5:0] _T_68146; // @[Modules.scala 40:46:@16384.4]
  wire [4:0] _T_68147; // @[Modules.scala 40:46:@16385.4]
  wire [4:0] _T_68148; // @[Modules.scala 40:46:@16386.4]
  wire [5:0] _T_68149; // @[Modules.scala 37:46:@16388.4]
  wire [4:0] _T_68150; // @[Modules.scala 37:46:@16389.4]
  wire [4:0] _T_68151; // @[Modules.scala 37:46:@16390.4]
  wire [5:0] _T_68212; // @[Modules.scala 37:46:@16465.4]
  wire [4:0] _T_68213; // @[Modules.scala 37:46:@16466.4]
  wire [4:0] _T_68214; // @[Modules.scala 37:46:@16467.4]
  wire [5:0] _T_68218; // @[Modules.scala 40:46:@16473.4]
  wire [4:0] _T_68219; // @[Modules.scala 40:46:@16474.4]
  wire [4:0] _T_68220; // @[Modules.scala 40:46:@16475.4]
  wire [5:0] _T_68225; // @[Modules.scala 46:47:@16480.4]
  wire [4:0] _T_68226; // @[Modules.scala 46:47:@16481.4]
  wire [4:0] _T_68227; // @[Modules.scala 46:47:@16482.4]
  wire [5:0] _T_68268; // @[Modules.scala 40:46:@16535.4]
  wire [4:0] _T_68269; // @[Modules.scala 40:46:@16536.4]
  wire [4:0] _T_68270; // @[Modules.scala 40:46:@16537.4]
  wire [5:0] _T_68271; // @[Modules.scala 37:46:@16539.4]
  wire [4:0] _T_68272; // @[Modules.scala 37:46:@16540.4]
  wire [4:0] _T_68273; // @[Modules.scala 37:46:@16541.4]
  wire [5:0] _T_68287; // @[Modules.scala 37:46:@16558.4]
  wire [4:0] _T_68288; // @[Modules.scala 37:46:@16559.4]
  wire [4:0] _T_68289; // @[Modules.scala 37:46:@16560.4]
  wire [5:0] _T_68310; // @[Modules.scala 43:47:@16584.4]
  wire [4:0] _T_68311; // @[Modules.scala 43:47:@16585.4]
  wire [4:0] _T_68312; // @[Modules.scala 43:47:@16586.4]
  wire [5:0] _T_68346; // @[Modules.scala 40:46:@16625.4]
  wire [4:0] _T_68347; // @[Modules.scala 40:46:@16626.4]
  wire [4:0] _T_68348; // @[Modules.scala 40:46:@16627.4]
  wire [5:0] _T_68368; // @[Modules.scala 40:46:@16652.4]
  wire [4:0] _T_68369; // @[Modules.scala 40:46:@16653.4]
  wire [4:0] _T_68370; // @[Modules.scala 40:46:@16654.4]
  wire [5:0] _T_68388; // @[Modules.scala 43:47:@16674.4]
  wire [4:0] _T_68389; // @[Modules.scala 43:47:@16675.4]
  wire [4:0] _T_68390; // @[Modules.scala 43:47:@16676.4]
  wire [5:0] _T_68395; // @[Modules.scala 43:47:@16681.4]
  wire [4:0] _T_68396; // @[Modules.scala 43:47:@16682.4]
  wire [4:0] _T_68397; // @[Modules.scala 43:47:@16683.4]
  wire [5:0] _T_68398; // @[Modules.scala 37:46:@16685.4]
  wire [4:0] _T_68399; // @[Modules.scala 37:46:@16686.4]
  wire [4:0] _T_68400; // @[Modules.scala 37:46:@16687.4]
  wire [5:0] _T_68404; // @[Modules.scala 40:46:@16693.4]
  wire [4:0] _T_68405; // @[Modules.scala 40:46:@16694.4]
  wire [4:0] _T_68406; // @[Modules.scala 40:46:@16695.4]
  wire [5:0] _T_68411; // @[Modules.scala 43:47:@16700.4]
  wire [4:0] _T_68412; // @[Modules.scala 43:47:@16701.4]
  wire [4:0] _T_68413; // @[Modules.scala 43:47:@16702.4]
  wire [5:0] _T_68454; // @[Modules.scala 43:47:@16748.4]
  wire [4:0] _T_68455; // @[Modules.scala 43:47:@16749.4]
  wire [4:0] _T_68456; // @[Modules.scala 43:47:@16750.4]
  wire [5:0] _T_68457; // @[Modules.scala 40:46:@16752.4]
  wire [4:0] _T_68458; // @[Modules.scala 40:46:@16753.4]
  wire [4:0] _T_68459; // @[Modules.scala 40:46:@16754.4]
  wire [5:0] _T_68466; // @[Modules.scala 40:46:@16764.4]
  wire [4:0] _T_68467; // @[Modules.scala 40:46:@16765.4]
  wire [4:0] _T_68468; // @[Modules.scala 40:46:@16766.4]
  wire [5:0] _T_68533; // @[Modules.scala 46:37:@16831.4]
  wire [4:0] _T_68534; // @[Modules.scala 46:37:@16832.4]
  wire [4:0] _T_68535; // @[Modules.scala 46:37:@16833.4]
  wire [5:0] _T_68536; // @[Modules.scala 46:47:@16834.4]
  wire [4:0] _T_68537; // @[Modules.scala 46:47:@16835.4]
  wire [4:0] _T_68538; // @[Modules.scala 46:47:@16836.4]
  wire [5:0] _T_68539; // @[Modules.scala 37:46:@16838.4]
  wire [4:0] _T_68540; // @[Modules.scala 37:46:@16839.4]
  wire [4:0] _T_68541; // @[Modules.scala 37:46:@16840.4]
  wire [5:0] _T_68611; // @[Modules.scala 46:47:@16913.4]
  wire [4:0] _T_68612; // @[Modules.scala 46:47:@16914.4]
  wire [4:0] _T_68613; // @[Modules.scala 46:47:@16915.4]
  wire [5:0] _T_68615; // @[Modules.scala 43:37:@16917.4]
  wire [4:0] _T_68616; // @[Modules.scala 43:37:@16918.4]
  wire [4:0] _T_68617; // @[Modules.scala 43:37:@16919.4]
  wire [5:0] _T_68618; // @[Modules.scala 43:47:@16920.4]
  wire [4:0] _T_68619; // @[Modules.scala 43:47:@16921.4]
  wire [4:0] _T_68620; // @[Modules.scala 43:47:@16922.4]
  wire [5:0] _T_68659; // @[Modules.scala 43:47:@16963.4]
  wire [4:0] _T_68660; // @[Modules.scala 43:47:@16964.4]
  wire [4:0] _T_68661; // @[Modules.scala 43:47:@16965.4]
  wire [5:0] _T_68672; // @[Modules.scala 40:46:@16978.4]
  wire [4:0] _T_68673; // @[Modules.scala 40:46:@16979.4]
  wire [4:0] _T_68674; // @[Modules.scala 40:46:@16980.4]
  wire [5:0] _T_68700; // @[Modules.scala 46:47:@17006.4]
  wire [4:0] _T_68701; // @[Modules.scala 46:47:@17007.4]
  wire [4:0] _T_68702; // @[Modules.scala 46:47:@17008.4]
  wire [10:0] buffer_4_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68710; // @[Modules.scala 50:57:@17017.4]
  wire [10:0] _T_68711; // @[Modules.scala 50:57:@17018.4]
  wire [10:0] buffer_4_392; // @[Modules.scala 50:57:@17019.4]
  wire [11:0] _T_68713; // @[Modules.scala 50:57:@17021.4]
  wire [10:0] _T_68714; // @[Modules.scala 50:57:@17022.4]
  wire [10:0] buffer_4_393; // @[Modules.scala 50:57:@17023.4]
  wire [10:0] buffer_4_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68716; // @[Modules.scala 50:57:@17025.4]
  wire [10:0] _T_68717; // @[Modules.scala 50:57:@17026.4]
  wire [10:0] buffer_4_394; // @[Modules.scala 50:57:@17027.4]
  wire [11:0] _T_68719; // @[Modules.scala 50:57:@17029.4]
  wire [10:0] _T_68720; // @[Modules.scala 50:57:@17030.4]
  wire [10:0] buffer_4_395; // @[Modules.scala 50:57:@17031.4]
  wire [10:0] buffer_4_8; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68722; // @[Modules.scala 50:57:@17033.4]
  wire [10:0] _T_68723; // @[Modules.scala 50:57:@17034.4]
  wire [10:0] buffer_4_396; // @[Modules.scala 50:57:@17035.4]
  wire [10:0] buffer_4_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68725; // @[Modules.scala 50:57:@17037.4]
  wire [10:0] _T_68726; // @[Modules.scala 50:57:@17038.4]
  wire [10:0] buffer_4_397; // @[Modules.scala 50:57:@17039.4]
  wire [10:0] buffer_4_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68728; // @[Modules.scala 50:57:@17041.4]
  wire [10:0] _T_68729; // @[Modules.scala 50:57:@17042.4]
  wire [10:0] buffer_4_398; // @[Modules.scala 50:57:@17043.4]
  wire [10:0] buffer_4_14; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68731; // @[Modules.scala 50:57:@17045.4]
  wire [10:0] _T_68732; // @[Modules.scala 50:57:@17046.4]
  wire [10:0] buffer_4_399; // @[Modules.scala 50:57:@17047.4]
  wire [11:0] _T_68740; // @[Modules.scala 50:57:@17057.4]
  wire [10:0] _T_68741; // @[Modules.scala 50:57:@17058.4]
  wire [10:0] buffer_4_402; // @[Modules.scala 50:57:@17059.4]
  wire [10:0] buffer_4_22; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68743; // @[Modules.scala 50:57:@17061.4]
  wire [10:0] _T_68744; // @[Modules.scala 50:57:@17062.4]
  wire [10:0] buffer_4_403; // @[Modules.scala 50:57:@17063.4]
  wire [11:0] _T_68749; // @[Modules.scala 50:57:@17069.4]
  wire [10:0] _T_68750; // @[Modules.scala 50:57:@17070.4]
  wire [10:0] buffer_4_405; // @[Modules.scala 50:57:@17071.4]
  wire [11:0] _T_68773; // @[Modules.scala 50:57:@17101.4]
  wire [10:0] _T_68774; // @[Modules.scala 50:57:@17102.4]
  wire [10:0] buffer_4_413; // @[Modules.scala 50:57:@17103.4]
  wire [10:0] buffer_4_44; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68776; // @[Modules.scala 50:57:@17105.4]
  wire [10:0] _T_68777; // @[Modules.scala 50:57:@17106.4]
  wire [10:0] buffer_4_414; // @[Modules.scala 50:57:@17107.4]
  wire [11:0] _T_68794; // @[Modules.scala 50:57:@17129.4]
  wire [10:0] _T_68795; // @[Modules.scala 50:57:@17130.4]
  wire [10:0] buffer_4_420; // @[Modules.scala 50:57:@17131.4]
  wire [10:0] buffer_4_58; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_59; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68797; // @[Modules.scala 50:57:@17133.4]
  wire [10:0] _T_68798; // @[Modules.scala 50:57:@17134.4]
  wire [10:0] buffer_4_421; // @[Modules.scala 50:57:@17135.4]
  wire [10:0] buffer_4_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68800; // @[Modules.scala 50:57:@17137.4]
  wire [10:0] _T_68801; // @[Modules.scala 50:57:@17138.4]
  wire [10:0] buffer_4_422; // @[Modules.scala 50:57:@17139.4]
  wire [11:0] _T_68803; // @[Modules.scala 50:57:@17141.4]
  wire [10:0] _T_68804; // @[Modules.scala 50:57:@17142.4]
  wire [10:0] buffer_4_423; // @[Modules.scala 50:57:@17143.4]
  wire [10:0] buffer_4_64; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68806; // @[Modules.scala 50:57:@17145.4]
  wire [10:0] _T_68807; // @[Modules.scala 50:57:@17146.4]
  wire [10:0] buffer_4_424; // @[Modules.scala 50:57:@17147.4]
  wire [10:0] buffer_4_67; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68809; // @[Modules.scala 50:57:@17149.4]
  wire [10:0] _T_68810; // @[Modules.scala 50:57:@17150.4]
  wire [10:0] buffer_4_425; // @[Modules.scala 50:57:@17151.4]
  wire [10:0] buffer_4_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68812; // @[Modules.scala 50:57:@17153.4]
  wire [10:0] _T_68813; // @[Modules.scala 50:57:@17154.4]
  wire [10:0] buffer_4_426; // @[Modules.scala 50:57:@17155.4]
  wire [11:0] _T_68815; // @[Modules.scala 50:57:@17157.4]
  wire [10:0] _T_68816; // @[Modules.scala 50:57:@17158.4]
  wire [10:0] buffer_4_427; // @[Modules.scala 50:57:@17159.4]
  wire [10:0] buffer_4_72; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68818; // @[Modules.scala 50:57:@17161.4]
  wire [10:0] _T_68819; // @[Modules.scala 50:57:@17162.4]
  wire [10:0] buffer_4_428; // @[Modules.scala 50:57:@17163.4]
  wire [10:0] buffer_4_76; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68824; // @[Modules.scala 50:57:@17169.4]
  wire [10:0] _T_68825; // @[Modules.scala 50:57:@17170.4]
  wire [10:0] buffer_4_430; // @[Modules.scala 50:57:@17171.4]
  wire [10:0] buffer_4_78; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68827; // @[Modules.scala 50:57:@17173.4]
  wire [10:0] _T_68828; // @[Modules.scala 50:57:@17174.4]
  wire [10:0] buffer_4_431; // @[Modules.scala 50:57:@17175.4]
  wire [10:0] buffer_4_80; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68830; // @[Modules.scala 50:57:@17177.4]
  wire [10:0] _T_68831; // @[Modules.scala 50:57:@17178.4]
  wire [10:0] buffer_4_432; // @[Modules.scala 50:57:@17179.4]
  wire [10:0] buffer_4_84; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68836; // @[Modules.scala 50:57:@17185.4]
  wire [10:0] _T_68837; // @[Modules.scala 50:57:@17186.4]
  wire [10:0] buffer_4_434; // @[Modules.scala 50:57:@17187.4]
  wire [10:0] buffer_4_92; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68848; // @[Modules.scala 50:57:@17201.4]
  wire [10:0] _T_68849; // @[Modules.scala 50:57:@17202.4]
  wire [10:0] buffer_4_438; // @[Modules.scala 50:57:@17203.4]
  wire [10:0] buffer_4_94; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68851; // @[Modules.scala 50:57:@17205.4]
  wire [10:0] _T_68852; // @[Modules.scala 50:57:@17206.4]
  wire [10:0] buffer_4_439; // @[Modules.scala 50:57:@17207.4]
  wire [11:0] _T_68857; // @[Modules.scala 50:57:@17213.4]
  wire [10:0] _T_68858; // @[Modules.scala 50:57:@17214.4]
  wire [10:0] buffer_4_441; // @[Modules.scala 50:57:@17215.4]
  wire [10:0] buffer_4_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68860; // @[Modules.scala 50:57:@17217.4]
  wire [10:0] _T_68861; // @[Modules.scala 50:57:@17218.4]
  wire [10:0] buffer_4_442; // @[Modules.scala 50:57:@17219.4]
  wire [10:0] buffer_4_102; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68863; // @[Modules.scala 50:57:@17221.4]
  wire [10:0] _T_68864; // @[Modules.scala 50:57:@17222.4]
  wire [10:0] buffer_4_443; // @[Modules.scala 50:57:@17223.4]
  wire [10:0] buffer_4_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68866; // @[Modules.scala 50:57:@17225.4]
  wire [10:0] _T_68867; // @[Modules.scala 50:57:@17226.4]
  wire [10:0] buffer_4_444; // @[Modules.scala 50:57:@17227.4]
  wire [10:0] buffer_4_106; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68869; // @[Modules.scala 50:57:@17229.4]
  wire [10:0] _T_68870; // @[Modules.scala 50:57:@17230.4]
  wire [10:0] buffer_4_445; // @[Modules.scala 50:57:@17231.4]
  wire [10:0] buffer_4_114; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68881; // @[Modules.scala 50:57:@17245.4]
  wire [10:0] _T_68882; // @[Modules.scala 50:57:@17246.4]
  wire [10:0] buffer_4_449; // @[Modules.scala 50:57:@17247.4]
  wire [10:0] buffer_4_116; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68884; // @[Modules.scala 50:57:@17249.4]
  wire [10:0] _T_68885; // @[Modules.scala 50:57:@17250.4]
  wire [10:0] buffer_4_450; // @[Modules.scala 50:57:@17251.4]
  wire [10:0] buffer_4_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68890; // @[Modules.scala 50:57:@17257.4]
  wire [10:0] _T_68891; // @[Modules.scala 50:57:@17258.4]
  wire [10:0] buffer_4_452; // @[Modules.scala 50:57:@17259.4]
  wire [10:0] buffer_4_122; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68893; // @[Modules.scala 50:57:@17261.4]
  wire [10:0] _T_68894; // @[Modules.scala 50:57:@17262.4]
  wire [10:0] buffer_4_453; // @[Modules.scala 50:57:@17263.4]
  wire [10:0] buffer_4_128; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68902; // @[Modules.scala 50:57:@17273.4]
  wire [10:0] _T_68903; // @[Modules.scala 50:57:@17274.4]
  wire [10:0] buffer_4_456; // @[Modules.scala 50:57:@17275.4]
  wire [10:0] buffer_4_130; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68905; // @[Modules.scala 50:57:@17277.4]
  wire [10:0] _T_68906; // @[Modules.scala 50:57:@17278.4]
  wire [10:0] buffer_4_457; // @[Modules.scala 50:57:@17279.4]
  wire [11:0] _T_68920; // @[Modules.scala 50:57:@17297.4]
  wire [10:0] _T_68921; // @[Modules.scala 50:57:@17298.4]
  wire [10:0] buffer_4_462; // @[Modules.scala 50:57:@17299.4]
  wire [11:0] _T_68923; // @[Modules.scala 50:57:@17301.4]
  wire [10:0] _T_68924; // @[Modules.scala 50:57:@17302.4]
  wire [10:0] buffer_4_463; // @[Modules.scala 50:57:@17303.4]
  wire [10:0] buffer_4_148; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_149; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68932; // @[Modules.scala 50:57:@17313.4]
  wire [10:0] _T_68933; // @[Modules.scala 50:57:@17314.4]
  wire [10:0] buffer_4_466; // @[Modules.scala 50:57:@17315.4]
  wire [10:0] buffer_4_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68935; // @[Modules.scala 50:57:@17317.4]
  wire [10:0] _T_68936; // @[Modules.scala 50:57:@17318.4]
  wire [10:0] buffer_4_467; // @[Modules.scala 50:57:@17319.4]
  wire [10:0] buffer_4_154; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68941; // @[Modules.scala 50:57:@17325.4]
  wire [10:0] _T_68942; // @[Modules.scala 50:57:@17326.4]
  wire [10:0] buffer_4_469; // @[Modules.scala 50:57:@17327.4]
  wire [11:0] _T_68950; // @[Modules.scala 50:57:@17337.4]
  wire [10:0] _T_68951; // @[Modules.scala 50:57:@17338.4]
  wire [10:0] buffer_4_472; // @[Modules.scala 50:57:@17339.4]
  wire [11:0] _T_68959; // @[Modules.scala 50:57:@17349.4]
  wire [10:0] _T_68960; // @[Modules.scala 50:57:@17350.4]
  wire [10:0] buffer_4_475; // @[Modules.scala 50:57:@17351.4]
  wire [10:0] buffer_4_172; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68968; // @[Modules.scala 50:57:@17361.4]
  wire [10:0] _T_68969; // @[Modules.scala 50:57:@17362.4]
  wire [10:0] buffer_4_478; // @[Modules.scala 50:57:@17363.4]
  wire [10:0] buffer_4_176; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68974; // @[Modules.scala 50:57:@17369.4]
  wire [10:0] _T_68975; // @[Modules.scala 50:57:@17370.4]
  wire [10:0] buffer_4_480; // @[Modules.scala 50:57:@17371.4]
  wire [11:0] _T_68980; // @[Modules.scala 50:57:@17377.4]
  wire [10:0] _T_68981; // @[Modules.scala 50:57:@17378.4]
  wire [10:0] buffer_4_482; // @[Modules.scala 50:57:@17379.4]
  wire [10:0] buffer_4_182; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68983; // @[Modules.scala 50:57:@17381.4]
  wire [10:0] _T_68984; // @[Modules.scala 50:57:@17382.4]
  wire [10:0] buffer_4_483; // @[Modules.scala 50:57:@17383.4]
  wire [10:0] buffer_4_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68986; // @[Modules.scala 50:57:@17385.4]
  wire [10:0] _T_68987; // @[Modules.scala 50:57:@17386.4]
  wire [10:0] buffer_4_484; // @[Modules.scala 50:57:@17387.4]
  wire [10:0] buffer_4_190; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68995; // @[Modules.scala 50:57:@17397.4]
  wire [10:0] _T_68996; // @[Modules.scala 50:57:@17398.4]
  wire [10:0] buffer_4_487; // @[Modules.scala 50:57:@17399.4]
  wire [11:0] _T_68998; // @[Modules.scala 50:57:@17401.4]
  wire [10:0] _T_68999; // @[Modules.scala 50:57:@17402.4]
  wire [10:0] buffer_4_488; // @[Modules.scala 50:57:@17403.4]
  wire [10:0] buffer_4_194; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69001; // @[Modules.scala 50:57:@17405.4]
  wire [10:0] _T_69002; // @[Modules.scala 50:57:@17406.4]
  wire [10:0] buffer_4_489; // @[Modules.scala 50:57:@17407.4]
  wire [10:0] buffer_4_196; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69004; // @[Modules.scala 50:57:@17409.4]
  wire [10:0] _T_69005; // @[Modules.scala 50:57:@17410.4]
  wire [10:0] buffer_4_490; // @[Modules.scala 50:57:@17411.4]
  wire [10:0] buffer_4_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69007; // @[Modules.scala 50:57:@17413.4]
  wire [10:0] _T_69008; // @[Modules.scala 50:57:@17414.4]
  wire [10:0] buffer_4_491; // @[Modules.scala 50:57:@17415.4]
  wire [11:0] _T_69010; // @[Modules.scala 50:57:@17417.4]
  wire [10:0] _T_69011; // @[Modules.scala 50:57:@17418.4]
  wire [10:0] buffer_4_492; // @[Modules.scala 50:57:@17419.4]
  wire [10:0] buffer_4_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69013; // @[Modules.scala 50:57:@17421.4]
  wire [10:0] _T_69014; // @[Modules.scala 50:57:@17422.4]
  wire [10:0] buffer_4_493; // @[Modules.scala 50:57:@17423.4]
  wire [11:0] _T_69016; // @[Modules.scala 50:57:@17425.4]
  wire [10:0] _T_69017; // @[Modules.scala 50:57:@17426.4]
  wire [10:0] buffer_4_494; // @[Modules.scala 50:57:@17427.4]
  wire [10:0] buffer_4_206; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69019; // @[Modules.scala 50:57:@17429.4]
  wire [10:0] _T_69020; // @[Modules.scala 50:57:@17430.4]
  wire [10:0] buffer_4_495; // @[Modules.scala 50:57:@17431.4]
  wire [10:0] buffer_4_208; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69022; // @[Modules.scala 50:57:@17433.4]
  wire [10:0] _T_69023; // @[Modules.scala 50:57:@17434.4]
  wire [10:0] buffer_4_496; // @[Modules.scala 50:57:@17435.4]
  wire [10:0] buffer_4_210; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69025; // @[Modules.scala 50:57:@17437.4]
  wire [10:0] _T_69026; // @[Modules.scala 50:57:@17438.4]
  wire [10:0] buffer_4_497; // @[Modules.scala 50:57:@17439.4]
  wire [10:0] buffer_4_216; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69034; // @[Modules.scala 50:57:@17449.4]
  wire [10:0] _T_69035; // @[Modules.scala 50:57:@17450.4]
  wire [10:0] buffer_4_500; // @[Modules.scala 50:57:@17451.4]
  wire [10:0] buffer_4_218; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69037; // @[Modules.scala 50:57:@17453.4]
  wire [10:0] _T_69038; // @[Modules.scala 50:57:@17454.4]
  wire [10:0] buffer_4_501; // @[Modules.scala 50:57:@17455.4]
  wire [11:0] _T_69040; // @[Modules.scala 50:57:@17457.4]
  wire [10:0] _T_69041; // @[Modules.scala 50:57:@17458.4]
  wire [10:0] buffer_4_502; // @[Modules.scala 50:57:@17459.4]
  wire [10:0] buffer_4_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69049; // @[Modules.scala 50:57:@17469.4]
  wire [10:0] _T_69050; // @[Modules.scala 50:57:@17470.4]
  wire [10:0] buffer_4_505; // @[Modules.scala 50:57:@17471.4]
  wire [10:0] buffer_4_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69055; // @[Modules.scala 50:57:@17477.4]
  wire [10:0] _T_69056; // @[Modules.scala 50:57:@17478.4]
  wire [10:0] buffer_4_507; // @[Modules.scala 50:57:@17479.4]
  wire [11:0] _T_69058; // @[Modules.scala 50:57:@17481.4]
  wire [10:0] _T_69059; // @[Modules.scala 50:57:@17482.4]
  wire [10:0] buffer_4_508; // @[Modules.scala 50:57:@17483.4]
  wire [11:0] _T_69067; // @[Modules.scala 50:57:@17493.4]
  wire [10:0] _T_69068; // @[Modules.scala 50:57:@17494.4]
  wire [10:0] buffer_4_511; // @[Modules.scala 50:57:@17495.4]
  wire [11:0] _T_69070; // @[Modules.scala 50:57:@17497.4]
  wire [10:0] _T_69071; // @[Modules.scala 50:57:@17498.4]
  wire [10:0] buffer_4_512; // @[Modules.scala 50:57:@17499.4]
  wire [10:0] buffer_4_243; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69073; // @[Modules.scala 50:57:@17501.4]
  wire [10:0] _T_69074; // @[Modules.scala 50:57:@17502.4]
  wire [10:0] buffer_4_513; // @[Modules.scala 50:57:@17503.4]
  wire [10:0] buffer_4_246; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69079; // @[Modules.scala 50:57:@17509.4]
  wire [10:0] _T_69080; // @[Modules.scala 50:57:@17510.4]
  wire [10:0] buffer_4_515; // @[Modules.scala 50:57:@17511.4]
  wire [11:0] _T_69088; // @[Modules.scala 50:57:@17521.4]
  wire [10:0] _T_69089; // @[Modules.scala 50:57:@17522.4]
  wire [10:0] buffer_4_518; // @[Modules.scala 50:57:@17523.4]
  wire [10:0] buffer_4_256; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_257; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69094; // @[Modules.scala 50:57:@17529.4]
  wire [10:0] _T_69095; // @[Modules.scala 50:57:@17530.4]
  wire [10:0] buffer_4_520; // @[Modules.scala 50:57:@17531.4]
  wire [10:0] buffer_4_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69097; // @[Modules.scala 50:57:@17533.4]
  wire [10:0] _T_69098; // @[Modules.scala 50:57:@17534.4]
  wire [10:0] buffer_4_521; // @[Modules.scala 50:57:@17535.4]
  wire [10:0] buffer_4_260; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69100; // @[Modules.scala 50:57:@17537.4]
  wire [10:0] _T_69101; // @[Modules.scala 50:57:@17538.4]
  wire [10:0] buffer_4_522; // @[Modules.scala 50:57:@17539.4]
  wire [11:0] _T_69103; // @[Modules.scala 50:57:@17541.4]
  wire [10:0] _T_69104; // @[Modules.scala 50:57:@17542.4]
  wire [10:0] buffer_4_523; // @[Modules.scala 50:57:@17543.4]
  wire [11:0] _T_69109; // @[Modules.scala 50:57:@17549.4]
  wire [10:0] _T_69110; // @[Modules.scala 50:57:@17550.4]
  wire [10:0] buffer_4_525; // @[Modules.scala 50:57:@17551.4]
  wire [10:0] buffer_4_272; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69118; // @[Modules.scala 50:57:@17561.4]
  wire [10:0] _T_69119; // @[Modules.scala 50:57:@17562.4]
  wire [10:0] buffer_4_528; // @[Modules.scala 50:57:@17563.4]
  wire [11:0] _T_69127; // @[Modules.scala 50:57:@17573.4]
  wire [10:0] _T_69128; // @[Modules.scala 50:57:@17574.4]
  wire [10:0] buffer_4_531; // @[Modules.scala 50:57:@17575.4]
  wire [11:0] _T_69139; // @[Modules.scala 50:57:@17589.4]
  wire [10:0] _T_69140; // @[Modules.scala 50:57:@17590.4]
  wire [10:0] buffer_4_535; // @[Modules.scala 50:57:@17591.4]
  wire [10:0] buffer_4_290; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69145; // @[Modules.scala 50:57:@17597.4]
  wire [10:0] _T_69146; // @[Modules.scala 50:57:@17598.4]
  wire [10:0] buffer_4_537; // @[Modules.scala 50:57:@17599.4]
  wire [10:0] buffer_4_292; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69148; // @[Modules.scala 50:57:@17601.4]
  wire [10:0] _T_69149; // @[Modules.scala 50:57:@17602.4]
  wire [10:0] buffer_4_538; // @[Modules.scala 50:57:@17603.4]
  wire [11:0] _T_69151; // @[Modules.scala 50:57:@17605.4]
  wire [10:0] _T_69152; // @[Modules.scala 50:57:@17606.4]
  wire [10:0] buffer_4_539; // @[Modules.scala 50:57:@17607.4]
  wire [11:0] _T_69157; // @[Modules.scala 50:57:@17613.4]
  wire [10:0] _T_69158; // @[Modules.scala 50:57:@17614.4]
  wire [10:0] buffer_4_541; // @[Modules.scala 50:57:@17615.4]
  wire [11:0] _T_69166; // @[Modules.scala 50:57:@17625.4]
  wire [10:0] _T_69167; // @[Modules.scala 50:57:@17626.4]
  wire [10:0] buffer_4_544; // @[Modules.scala 50:57:@17627.4]
  wire [10:0] buffer_4_306; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69169; // @[Modules.scala 50:57:@17629.4]
  wire [10:0] _T_69170; // @[Modules.scala 50:57:@17630.4]
  wire [10:0] buffer_4_545; // @[Modules.scala 50:57:@17631.4]
  wire [10:0] buffer_4_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69175; // @[Modules.scala 50:57:@17637.4]
  wire [10:0] _T_69176; // @[Modules.scala 50:57:@17638.4]
  wire [10:0] buffer_4_547; // @[Modules.scala 50:57:@17639.4]
  wire [11:0] _T_69178; // @[Modules.scala 50:57:@17641.4]
  wire [10:0] _T_69179; // @[Modules.scala 50:57:@17642.4]
  wire [10:0] buffer_4_548; // @[Modules.scala 50:57:@17643.4]
  wire [10:0] buffer_4_316; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69184; // @[Modules.scala 50:57:@17649.4]
  wire [10:0] _T_69185; // @[Modules.scala 50:57:@17650.4]
  wire [10:0] buffer_4_550; // @[Modules.scala 50:57:@17651.4]
  wire [11:0] _T_69190; // @[Modules.scala 50:57:@17657.4]
  wire [10:0] _T_69191; // @[Modules.scala 50:57:@17658.4]
  wire [10:0] buffer_4_552; // @[Modules.scala 50:57:@17659.4]
  wire [10:0] buffer_4_324; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69196; // @[Modules.scala 50:57:@17665.4]
  wire [10:0] _T_69197; // @[Modules.scala 50:57:@17666.4]
  wire [10:0] buffer_4_554; // @[Modules.scala 50:57:@17667.4]
  wire [10:0] buffer_4_330; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69205; // @[Modules.scala 50:57:@17677.4]
  wire [10:0] _T_69206; // @[Modules.scala 50:57:@17678.4]
  wire [10:0] buffer_4_557; // @[Modules.scala 50:57:@17679.4]
  wire [11:0] _T_69208; // @[Modules.scala 50:57:@17681.4]
  wire [10:0] _T_69209; // @[Modules.scala 50:57:@17682.4]
  wire [10:0] buffer_4_558; // @[Modules.scala 50:57:@17683.4]
  wire [10:0] buffer_4_334; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69211; // @[Modules.scala 50:57:@17685.4]
  wire [10:0] _T_69212; // @[Modules.scala 50:57:@17686.4]
  wire [10:0] buffer_4_559; // @[Modules.scala 50:57:@17687.4]
  wire [10:0] buffer_4_336; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69214; // @[Modules.scala 50:57:@17689.4]
  wire [10:0] _T_69215; // @[Modules.scala 50:57:@17690.4]
  wire [10:0] buffer_4_560; // @[Modules.scala 50:57:@17691.4]
  wire [10:0] buffer_4_338; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69217; // @[Modules.scala 50:57:@17693.4]
  wire [10:0] _T_69218; // @[Modules.scala 50:57:@17694.4]
  wire [10:0] buffer_4_561; // @[Modules.scala 50:57:@17695.4]
  wire [11:0] _T_69223; // @[Modules.scala 50:57:@17701.4]
  wire [10:0] _T_69224; // @[Modules.scala 50:57:@17702.4]
  wire [10:0] buffer_4_563; // @[Modules.scala 50:57:@17703.4]
  wire [11:0] _T_69226; // @[Modules.scala 50:57:@17705.4]
  wire [10:0] _T_69227; // @[Modules.scala 50:57:@17706.4]
  wire [10:0] buffer_4_564; // @[Modules.scala 50:57:@17707.4]
  wire [10:0] buffer_4_348; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69232; // @[Modules.scala 50:57:@17713.4]
  wire [10:0] _T_69233; // @[Modules.scala 50:57:@17714.4]
  wire [10:0] buffer_4_566; // @[Modules.scala 50:57:@17715.4]
  wire [10:0] buffer_4_352; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69238; // @[Modules.scala 50:57:@17721.4]
  wire [10:0] _T_69239; // @[Modules.scala 50:57:@17722.4]
  wire [10:0] buffer_4_568; // @[Modules.scala 50:57:@17723.4]
  wire [10:0] buffer_4_362; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69253; // @[Modules.scala 50:57:@17741.4]
  wire [10:0] _T_69254; // @[Modules.scala 50:57:@17742.4]
  wire [10:0] buffer_4_573; // @[Modules.scala 50:57:@17743.4]
  wire [10:0] buffer_4_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69271; // @[Modules.scala 50:57:@17765.4]
  wire [10:0] _T_69272; // @[Modules.scala 50:57:@17766.4]
  wire [10:0] buffer_4_579; // @[Modules.scala 50:57:@17767.4]
  wire [10:0] buffer_4_376; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69274; // @[Modules.scala 50:57:@17769.4]
  wire [10:0] _T_69275; // @[Modules.scala 50:57:@17770.4]
  wire [10:0] buffer_4_580; // @[Modules.scala 50:57:@17771.4]
  wire [11:0] _T_69277; // @[Modules.scala 50:57:@17773.4]
  wire [10:0] _T_69278; // @[Modules.scala 50:57:@17774.4]
  wire [10:0] buffer_4_581; // @[Modules.scala 50:57:@17775.4]
  wire [11:0] _T_69280; // @[Modules.scala 50:57:@17777.4]
  wire [10:0] _T_69281; // @[Modules.scala 50:57:@17778.4]
  wire [10:0] buffer_4_582; // @[Modules.scala 50:57:@17779.4]
  wire [10:0] buffer_4_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69283; // @[Modules.scala 50:57:@17781.4]
  wire [10:0] _T_69284; // @[Modules.scala 50:57:@17782.4]
  wire [10:0] buffer_4_583; // @[Modules.scala 50:57:@17783.4]
  wire [11:0] _T_69286; // @[Modules.scala 50:57:@17785.4]
  wire [10:0] _T_69287; // @[Modules.scala 50:57:@17786.4]
  wire [10:0] buffer_4_584; // @[Modules.scala 50:57:@17787.4]
  wire [10:0] buffer_4_386; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69289; // @[Modules.scala 50:57:@17789.4]
  wire [10:0] _T_69290; // @[Modules.scala 50:57:@17790.4]
  wire [10:0] buffer_4_585; // @[Modules.scala 50:57:@17791.4]
  wire [10:0] buffer_4_390; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69295; // @[Modules.scala 50:57:@17797.4]
  wire [10:0] _T_69296; // @[Modules.scala 50:57:@17798.4]
  wire [10:0] buffer_4_587; // @[Modules.scala 50:57:@17799.4]
  wire [11:0] _T_69298; // @[Modules.scala 53:83:@17801.4]
  wire [10:0] _T_69299; // @[Modules.scala 53:83:@17802.4]
  wire [10:0] buffer_4_588; // @[Modules.scala 53:83:@17803.4]
  wire [11:0] _T_69301; // @[Modules.scala 53:83:@17805.4]
  wire [10:0] _T_69302; // @[Modules.scala 53:83:@17806.4]
  wire [10:0] buffer_4_589; // @[Modules.scala 53:83:@17807.4]
  wire [11:0] _T_69304; // @[Modules.scala 53:83:@17809.4]
  wire [10:0] _T_69305; // @[Modules.scala 53:83:@17810.4]
  wire [10:0] buffer_4_590; // @[Modules.scala 53:83:@17811.4]
  wire [11:0] _T_69307; // @[Modules.scala 53:83:@17813.4]
  wire [10:0] _T_69308; // @[Modules.scala 53:83:@17814.4]
  wire [10:0] buffer_4_591; // @[Modules.scala 53:83:@17815.4]
  wire [11:0] _T_69310; // @[Modules.scala 53:83:@17817.4]
  wire [10:0] _T_69311; // @[Modules.scala 53:83:@17818.4]
  wire [10:0] buffer_4_592; // @[Modules.scala 53:83:@17819.4]
  wire [11:0] _T_69313; // @[Modules.scala 53:83:@17821.4]
  wire [10:0] _T_69314; // @[Modules.scala 53:83:@17822.4]
  wire [10:0] buffer_4_593; // @[Modules.scala 53:83:@17823.4]
  wire [11:0] _T_69316; // @[Modules.scala 53:83:@17825.4]
  wire [10:0] _T_69317; // @[Modules.scala 53:83:@17826.4]
  wire [10:0] buffer_4_594; // @[Modules.scala 53:83:@17827.4]
  wire [11:0] _T_69319; // @[Modules.scala 53:83:@17829.4]
  wire [10:0] _T_69320; // @[Modules.scala 53:83:@17830.4]
  wire [10:0] buffer_4_595; // @[Modules.scala 53:83:@17831.4]
  wire [11:0] _T_69328; // @[Modules.scala 53:83:@17841.4]
  wire [10:0] _T_69329; // @[Modules.scala 53:83:@17842.4]
  wire [10:0] buffer_4_598; // @[Modules.scala 53:83:@17843.4]
  wire [11:0] _T_69331; // @[Modules.scala 53:83:@17845.4]
  wire [10:0] _T_69332; // @[Modules.scala 53:83:@17846.4]
  wire [10:0] buffer_4_599; // @[Modules.scala 53:83:@17847.4]
  wire [11:0] _T_69340; // @[Modules.scala 53:83:@17857.4]
  wire [10:0] _T_69341; // @[Modules.scala 53:83:@17858.4]
  wire [10:0] buffer_4_602; // @[Modules.scala 53:83:@17859.4]
  wire [11:0] _T_69343; // @[Modules.scala 53:83:@17861.4]
  wire [10:0] _T_69344; // @[Modules.scala 53:83:@17862.4]
  wire [10:0] buffer_4_603; // @[Modules.scala 53:83:@17863.4]
  wire [11:0] _T_69346; // @[Modules.scala 53:83:@17865.4]
  wire [10:0] _T_69347; // @[Modules.scala 53:83:@17866.4]
  wire [10:0] buffer_4_604; // @[Modules.scala 53:83:@17867.4]
  wire [11:0] _T_69349; // @[Modules.scala 53:83:@17869.4]
  wire [10:0] _T_69350; // @[Modules.scala 53:83:@17870.4]
  wire [10:0] buffer_4_605; // @[Modules.scala 53:83:@17871.4]
  wire [11:0] _T_69352; // @[Modules.scala 53:83:@17873.4]
  wire [10:0] _T_69353; // @[Modules.scala 53:83:@17874.4]
  wire [10:0] buffer_4_606; // @[Modules.scala 53:83:@17875.4]
  wire [11:0] _T_69355; // @[Modules.scala 53:83:@17877.4]
  wire [10:0] _T_69356; // @[Modules.scala 53:83:@17878.4]
  wire [10:0] buffer_4_607; // @[Modules.scala 53:83:@17879.4]
  wire [11:0] _T_69358; // @[Modules.scala 53:83:@17881.4]
  wire [10:0] _T_69359; // @[Modules.scala 53:83:@17882.4]
  wire [10:0] buffer_4_608; // @[Modules.scala 53:83:@17883.4]
  wire [11:0] _T_69361; // @[Modules.scala 53:83:@17885.4]
  wire [10:0] _T_69362; // @[Modules.scala 53:83:@17886.4]
  wire [10:0] buffer_4_609; // @[Modules.scala 53:83:@17887.4]
  wire [11:0] _T_69364; // @[Modules.scala 53:83:@17889.4]
  wire [10:0] _T_69365; // @[Modules.scala 53:83:@17890.4]
  wire [10:0] buffer_4_610; // @[Modules.scala 53:83:@17891.4]
  wire [11:0] _T_69367; // @[Modules.scala 53:83:@17893.4]
  wire [10:0] _T_69368; // @[Modules.scala 53:83:@17894.4]
  wire [10:0] buffer_4_611; // @[Modules.scala 53:83:@17895.4]
  wire [11:0] _T_69370; // @[Modules.scala 53:83:@17897.4]
  wire [10:0] _T_69371; // @[Modules.scala 53:83:@17898.4]
  wire [10:0] buffer_4_612; // @[Modules.scala 53:83:@17899.4]
  wire [11:0] _T_69373; // @[Modules.scala 53:83:@17901.4]
  wire [10:0] _T_69374; // @[Modules.scala 53:83:@17902.4]
  wire [10:0] buffer_4_613; // @[Modules.scala 53:83:@17903.4]
  wire [11:0] _T_69376; // @[Modules.scala 53:83:@17905.4]
  wire [10:0] _T_69377; // @[Modules.scala 53:83:@17906.4]
  wire [10:0] buffer_4_614; // @[Modules.scala 53:83:@17907.4]
  wire [11:0] _T_69382; // @[Modules.scala 53:83:@17913.4]
  wire [10:0] _T_69383; // @[Modules.scala 53:83:@17914.4]
  wire [10:0] buffer_4_616; // @[Modules.scala 53:83:@17915.4]
  wire [11:0] _T_69385; // @[Modules.scala 53:83:@17917.4]
  wire [10:0] _T_69386; // @[Modules.scala 53:83:@17918.4]
  wire [10:0] buffer_4_617; // @[Modules.scala 53:83:@17919.4]
  wire [11:0] _T_69388; // @[Modules.scala 53:83:@17921.4]
  wire [10:0] _T_69389; // @[Modules.scala 53:83:@17922.4]
  wire [10:0] buffer_4_618; // @[Modules.scala 53:83:@17923.4]
  wire [11:0] _T_69394; // @[Modules.scala 53:83:@17929.4]
  wire [10:0] _T_69395; // @[Modules.scala 53:83:@17930.4]
  wire [10:0] buffer_4_620; // @[Modules.scala 53:83:@17931.4]
  wire [11:0] _T_69403; // @[Modules.scala 53:83:@17941.4]
  wire [10:0] _T_69404; // @[Modules.scala 53:83:@17942.4]
  wire [10:0] buffer_4_623; // @[Modules.scala 53:83:@17943.4]
  wire [11:0] _T_69409; // @[Modules.scala 53:83:@17949.4]
  wire [10:0] _T_69410; // @[Modules.scala 53:83:@17950.4]
  wire [10:0] buffer_4_625; // @[Modules.scala 53:83:@17951.4]
  wire [11:0] _T_69412; // @[Modules.scala 53:83:@17953.4]
  wire [10:0] _T_69413; // @[Modules.scala 53:83:@17954.4]
  wire [10:0] buffer_4_626; // @[Modules.scala 53:83:@17955.4]
  wire [11:0] _T_69415; // @[Modules.scala 53:83:@17957.4]
  wire [10:0] _T_69416; // @[Modules.scala 53:83:@17958.4]
  wire [10:0] buffer_4_627; // @[Modules.scala 53:83:@17959.4]
  wire [11:0] _T_69418; // @[Modules.scala 53:83:@17961.4]
  wire [10:0] _T_69419; // @[Modules.scala 53:83:@17962.4]
  wire [10:0] buffer_4_628; // @[Modules.scala 53:83:@17963.4]
  wire [11:0] _T_69421; // @[Modules.scala 53:83:@17965.4]
  wire [10:0] _T_69422; // @[Modules.scala 53:83:@17966.4]
  wire [10:0] buffer_4_629; // @[Modules.scala 53:83:@17967.4]
  wire [11:0] _T_69424; // @[Modules.scala 53:83:@17969.4]
  wire [10:0] _T_69425; // @[Modules.scala 53:83:@17970.4]
  wire [10:0] buffer_4_630; // @[Modules.scala 53:83:@17971.4]
  wire [11:0] _T_69427; // @[Modules.scala 53:83:@17973.4]
  wire [10:0] _T_69428; // @[Modules.scala 53:83:@17974.4]
  wire [10:0] buffer_4_631; // @[Modules.scala 53:83:@17975.4]
  wire [11:0] _T_69430; // @[Modules.scala 53:83:@17977.4]
  wire [10:0] _T_69431; // @[Modules.scala 53:83:@17978.4]
  wire [10:0] buffer_4_632; // @[Modules.scala 53:83:@17979.4]
  wire [11:0] _T_69433; // @[Modules.scala 53:83:@17981.4]
  wire [10:0] _T_69434; // @[Modules.scala 53:83:@17982.4]
  wire [10:0] buffer_4_633; // @[Modules.scala 53:83:@17983.4]
  wire [11:0] _T_69436; // @[Modules.scala 53:83:@17985.4]
  wire [10:0] _T_69437; // @[Modules.scala 53:83:@17986.4]
  wire [10:0] buffer_4_634; // @[Modules.scala 53:83:@17987.4]
  wire [11:0] _T_69439; // @[Modules.scala 53:83:@17989.4]
  wire [10:0] _T_69440; // @[Modules.scala 53:83:@17990.4]
  wire [10:0] buffer_4_635; // @[Modules.scala 53:83:@17991.4]
  wire [11:0] _T_69442; // @[Modules.scala 53:83:@17993.4]
  wire [10:0] _T_69443; // @[Modules.scala 53:83:@17994.4]
  wire [10:0] buffer_4_636; // @[Modules.scala 53:83:@17995.4]
  wire [11:0] _T_69445; // @[Modules.scala 53:83:@17997.4]
  wire [10:0] _T_69446; // @[Modules.scala 53:83:@17998.4]
  wire [10:0] buffer_4_637; // @[Modules.scala 53:83:@17999.4]
  wire [11:0] _T_69448; // @[Modules.scala 53:83:@18001.4]
  wire [10:0] _T_69449; // @[Modules.scala 53:83:@18002.4]
  wire [10:0] buffer_4_638; // @[Modules.scala 53:83:@18003.4]
  wire [11:0] _T_69451; // @[Modules.scala 53:83:@18005.4]
  wire [10:0] _T_69452; // @[Modules.scala 53:83:@18006.4]
  wire [10:0] buffer_4_639; // @[Modules.scala 53:83:@18007.4]
  wire [11:0] _T_69454; // @[Modules.scala 53:83:@18009.4]
  wire [10:0] _T_69455; // @[Modules.scala 53:83:@18010.4]
  wire [10:0] buffer_4_640; // @[Modules.scala 53:83:@18011.4]
  wire [11:0] _T_69457; // @[Modules.scala 53:83:@18013.4]
  wire [10:0] _T_69458; // @[Modules.scala 53:83:@18014.4]
  wire [10:0] buffer_4_641; // @[Modules.scala 53:83:@18015.4]
  wire [11:0] _T_69460; // @[Modules.scala 53:83:@18017.4]
  wire [10:0] _T_69461; // @[Modules.scala 53:83:@18018.4]
  wire [10:0] buffer_4_642; // @[Modules.scala 53:83:@18019.4]
  wire [11:0] _T_69463; // @[Modules.scala 53:83:@18021.4]
  wire [10:0] _T_69464; // @[Modules.scala 53:83:@18022.4]
  wire [10:0] buffer_4_643; // @[Modules.scala 53:83:@18023.4]
  wire [11:0] _T_69466; // @[Modules.scala 53:83:@18025.4]
  wire [10:0] _T_69467; // @[Modules.scala 53:83:@18026.4]
  wire [10:0] buffer_4_644; // @[Modules.scala 53:83:@18027.4]
  wire [11:0] _T_69469; // @[Modules.scala 53:83:@18029.4]
  wire [10:0] _T_69470; // @[Modules.scala 53:83:@18030.4]
  wire [10:0] buffer_4_645; // @[Modules.scala 53:83:@18031.4]
  wire [11:0] _T_69472; // @[Modules.scala 53:83:@18033.4]
  wire [10:0] _T_69473; // @[Modules.scala 53:83:@18034.4]
  wire [10:0] buffer_4_646; // @[Modules.scala 53:83:@18035.4]
  wire [11:0] _T_69475; // @[Modules.scala 53:83:@18037.4]
  wire [10:0] _T_69476; // @[Modules.scala 53:83:@18038.4]
  wire [10:0] buffer_4_647; // @[Modules.scala 53:83:@18039.4]
  wire [11:0] _T_69478; // @[Modules.scala 53:83:@18041.4]
  wire [10:0] _T_69479; // @[Modules.scala 53:83:@18042.4]
  wire [10:0] buffer_4_648; // @[Modules.scala 53:83:@18043.4]
  wire [11:0] _T_69481; // @[Modules.scala 53:83:@18045.4]
  wire [10:0] _T_69482; // @[Modules.scala 53:83:@18046.4]
  wire [10:0] buffer_4_649; // @[Modules.scala 53:83:@18047.4]
  wire [11:0] _T_69487; // @[Modules.scala 53:83:@18053.4]
  wire [10:0] _T_69488; // @[Modules.scala 53:83:@18054.4]
  wire [10:0] buffer_4_651; // @[Modules.scala 53:83:@18055.4]
  wire [11:0] _T_69490; // @[Modules.scala 53:83:@18057.4]
  wire [10:0] _T_69491; // @[Modules.scala 53:83:@18058.4]
  wire [10:0] buffer_4_652; // @[Modules.scala 53:83:@18059.4]
  wire [11:0] _T_69493; // @[Modules.scala 53:83:@18061.4]
  wire [10:0] _T_69494; // @[Modules.scala 53:83:@18062.4]
  wire [10:0] buffer_4_653; // @[Modules.scala 53:83:@18063.4]
  wire [11:0] _T_69496; // @[Modules.scala 53:83:@18065.4]
  wire [10:0] _T_69497; // @[Modules.scala 53:83:@18066.4]
  wire [10:0] buffer_4_654; // @[Modules.scala 53:83:@18067.4]
  wire [11:0] _T_69502; // @[Modules.scala 53:83:@18073.4]
  wire [10:0] _T_69503; // @[Modules.scala 53:83:@18074.4]
  wire [10:0] buffer_4_656; // @[Modules.scala 53:83:@18075.4]
  wire [11:0] _T_69505; // @[Modules.scala 53:83:@18077.4]
  wire [10:0] _T_69506; // @[Modules.scala 53:83:@18078.4]
  wire [10:0] buffer_4_657; // @[Modules.scala 53:83:@18079.4]
  wire [11:0] _T_69508; // @[Modules.scala 53:83:@18081.4]
  wire [10:0] _T_69509; // @[Modules.scala 53:83:@18082.4]
  wire [10:0] buffer_4_658; // @[Modules.scala 53:83:@18083.4]
  wire [11:0] _T_69511; // @[Modules.scala 53:83:@18085.4]
  wire [10:0] _T_69512; // @[Modules.scala 53:83:@18086.4]
  wire [10:0] buffer_4_659; // @[Modules.scala 53:83:@18087.4]
  wire [11:0] _T_69514; // @[Modules.scala 53:83:@18089.4]
  wire [10:0] _T_69515; // @[Modules.scala 53:83:@18090.4]
  wire [10:0] buffer_4_660; // @[Modules.scala 53:83:@18091.4]
  wire [11:0] _T_69517; // @[Modules.scala 53:83:@18093.4]
  wire [10:0] _T_69518; // @[Modules.scala 53:83:@18094.4]
  wire [10:0] buffer_4_661; // @[Modules.scala 53:83:@18095.4]
  wire [11:0] _T_69520; // @[Modules.scala 53:83:@18097.4]
  wire [10:0] _T_69521; // @[Modules.scala 53:83:@18098.4]
  wire [10:0] buffer_4_662; // @[Modules.scala 53:83:@18099.4]
  wire [11:0] _T_69526; // @[Modules.scala 53:83:@18105.4]
  wire [10:0] _T_69527; // @[Modules.scala 53:83:@18106.4]
  wire [10:0] buffer_4_664; // @[Modules.scala 53:83:@18107.4]
  wire [11:0] _T_69529; // @[Modules.scala 53:83:@18109.4]
  wire [10:0] _T_69530; // @[Modules.scala 53:83:@18110.4]
  wire [10:0] buffer_4_665; // @[Modules.scala 53:83:@18111.4]
  wire [11:0] _T_69532; // @[Modules.scala 53:83:@18113.4]
  wire [10:0] _T_69533; // @[Modules.scala 53:83:@18114.4]
  wire [10:0] buffer_4_666; // @[Modules.scala 53:83:@18115.4]
  wire [11:0] _T_69535; // @[Modules.scala 53:83:@18117.4]
  wire [10:0] _T_69536; // @[Modules.scala 53:83:@18118.4]
  wire [10:0] buffer_4_667; // @[Modules.scala 53:83:@18119.4]
  wire [11:0] _T_69538; // @[Modules.scala 53:83:@18121.4]
  wire [10:0] _T_69539; // @[Modules.scala 53:83:@18122.4]
  wire [10:0] buffer_4_668; // @[Modules.scala 53:83:@18123.4]
  wire [11:0] _T_69541; // @[Modules.scala 53:83:@18125.4]
  wire [10:0] _T_69542; // @[Modules.scala 53:83:@18126.4]
  wire [10:0] buffer_4_669; // @[Modules.scala 53:83:@18127.4]
  wire [11:0] _T_69544; // @[Modules.scala 53:83:@18129.4]
  wire [10:0] _T_69545; // @[Modules.scala 53:83:@18130.4]
  wire [10:0] buffer_4_670; // @[Modules.scala 53:83:@18131.4]
  wire [11:0] _T_69547; // @[Modules.scala 53:83:@18133.4]
  wire [10:0] _T_69548; // @[Modules.scala 53:83:@18134.4]
  wire [10:0] buffer_4_671; // @[Modules.scala 53:83:@18135.4]
  wire [11:0] _T_69550; // @[Modules.scala 53:83:@18137.4]
  wire [10:0] _T_69551; // @[Modules.scala 53:83:@18138.4]
  wire [10:0] buffer_4_672; // @[Modules.scala 53:83:@18139.4]
  wire [11:0] _T_69553; // @[Modules.scala 53:83:@18141.4]
  wire [10:0] _T_69554; // @[Modules.scala 53:83:@18142.4]
  wire [10:0] buffer_4_673; // @[Modules.scala 53:83:@18143.4]
  wire [11:0] _T_69556; // @[Modules.scala 53:83:@18145.4]
  wire [10:0] _T_69557; // @[Modules.scala 53:83:@18146.4]
  wire [10:0] buffer_4_674; // @[Modules.scala 53:83:@18147.4]
  wire [11:0] _T_69559; // @[Modules.scala 53:83:@18149.4]
  wire [10:0] _T_69560; // @[Modules.scala 53:83:@18150.4]
  wire [10:0] buffer_4_675; // @[Modules.scala 53:83:@18151.4]
  wire [11:0] _T_69562; // @[Modules.scala 53:83:@18153.4]
  wire [10:0] _T_69563; // @[Modules.scala 53:83:@18154.4]
  wire [10:0] buffer_4_676; // @[Modules.scala 53:83:@18155.4]
  wire [11:0] _T_69568; // @[Modules.scala 53:83:@18161.4]
  wire [10:0] _T_69569; // @[Modules.scala 53:83:@18162.4]
  wire [10:0] buffer_4_678; // @[Modules.scala 53:83:@18163.4]
  wire [11:0] _T_69571; // @[Modules.scala 53:83:@18165.4]
  wire [10:0] _T_69572; // @[Modules.scala 53:83:@18166.4]
  wire [10:0] buffer_4_679; // @[Modules.scala 53:83:@18167.4]
  wire [11:0] _T_69577; // @[Modules.scala 53:83:@18173.4]
  wire [10:0] _T_69578; // @[Modules.scala 53:83:@18174.4]
  wire [10:0] buffer_4_681; // @[Modules.scala 53:83:@18175.4]
  wire [11:0] _T_69580; // @[Modules.scala 53:83:@18177.4]
  wire [10:0] _T_69581; // @[Modules.scala 53:83:@18178.4]
  wire [10:0] buffer_4_682; // @[Modules.scala 53:83:@18179.4]
  wire [11:0] _T_69583; // @[Modules.scala 53:83:@18181.4]
  wire [10:0] _T_69584; // @[Modules.scala 53:83:@18182.4]
  wire [10:0] buffer_4_683; // @[Modules.scala 53:83:@18183.4]
  wire [11:0] _T_69586; // @[Modules.scala 53:83:@18185.4]
  wire [10:0] _T_69587; // @[Modules.scala 53:83:@18186.4]
  wire [10:0] buffer_4_684; // @[Modules.scala 53:83:@18187.4]
  wire [11:0] _T_69589; // @[Modules.scala 53:83:@18189.4]
  wire [10:0] _T_69590; // @[Modules.scala 53:83:@18190.4]
  wire [10:0] buffer_4_685; // @[Modules.scala 53:83:@18191.4]
  wire [11:0] _T_69592; // @[Modules.scala 56:109:@18193.4]
  wire [10:0] _T_69593; // @[Modules.scala 56:109:@18194.4]
  wire [10:0] buffer_4_686; // @[Modules.scala 56:109:@18195.4]
  wire [11:0] _T_69595; // @[Modules.scala 56:109:@18197.4]
  wire [10:0] _T_69596; // @[Modules.scala 56:109:@18198.4]
  wire [10:0] buffer_4_687; // @[Modules.scala 56:109:@18199.4]
  wire [11:0] _T_69598; // @[Modules.scala 56:109:@18201.4]
  wire [10:0] _T_69599; // @[Modules.scala 56:109:@18202.4]
  wire [10:0] buffer_4_688; // @[Modules.scala 56:109:@18203.4]
  wire [11:0] _T_69601; // @[Modules.scala 56:109:@18205.4]
  wire [10:0] _T_69602; // @[Modules.scala 56:109:@18206.4]
  wire [10:0] buffer_4_689; // @[Modules.scala 56:109:@18207.4]
  wire [11:0] _T_69607; // @[Modules.scala 56:109:@18213.4]
  wire [10:0] _T_69608; // @[Modules.scala 56:109:@18214.4]
  wire [10:0] buffer_4_691; // @[Modules.scala 56:109:@18215.4]
  wire [11:0] _T_69613; // @[Modules.scala 56:109:@18221.4]
  wire [10:0] _T_69614; // @[Modules.scala 56:109:@18222.4]
  wire [10:0] buffer_4_693; // @[Modules.scala 56:109:@18223.4]
  wire [11:0] _T_69616; // @[Modules.scala 56:109:@18225.4]
  wire [10:0] _T_69617; // @[Modules.scala 56:109:@18226.4]
  wire [10:0] buffer_4_694; // @[Modules.scala 56:109:@18227.4]
  wire [11:0] _T_69619; // @[Modules.scala 56:109:@18229.4]
  wire [10:0] _T_69620; // @[Modules.scala 56:109:@18230.4]
  wire [10:0] buffer_4_695; // @[Modules.scala 56:109:@18231.4]
  wire [11:0] _T_69622; // @[Modules.scala 56:109:@18233.4]
  wire [10:0] _T_69623; // @[Modules.scala 56:109:@18234.4]
  wire [10:0] buffer_4_696; // @[Modules.scala 56:109:@18235.4]
  wire [11:0] _T_69625; // @[Modules.scala 56:109:@18237.4]
  wire [10:0] _T_69626; // @[Modules.scala 56:109:@18238.4]
  wire [10:0] buffer_4_697; // @[Modules.scala 56:109:@18239.4]
  wire [11:0] _T_69628; // @[Modules.scala 56:109:@18241.4]
  wire [10:0] _T_69629; // @[Modules.scala 56:109:@18242.4]
  wire [10:0] buffer_4_698; // @[Modules.scala 56:109:@18243.4]
  wire [11:0] _T_69631; // @[Modules.scala 56:109:@18245.4]
  wire [10:0] _T_69632; // @[Modules.scala 56:109:@18246.4]
  wire [10:0] buffer_4_699; // @[Modules.scala 56:109:@18247.4]
  wire [11:0] _T_69634; // @[Modules.scala 56:109:@18249.4]
  wire [10:0] _T_69635; // @[Modules.scala 56:109:@18250.4]
  wire [10:0] buffer_4_700; // @[Modules.scala 56:109:@18251.4]
  wire [11:0] _T_69637; // @[Modules.scala 56:109:@18253.4]
  wire [10:0] _T_69638; // @[Modules.scala 56:109:@18254.4]
  wire [10:0] buffer_4_701; // @[Modules.scala 56:109:@18255.4]
  wire [11:0] _T_69640; // @[Modules.scala 56:109:@18257.4]
  wire [10:0] _T_69641; // @[Modules.scala 56:109:@18258.4]
  wire [10:0] buffer_4_702; // @[Modules.scala 56:109:@18259.4]
  wire [11:0] _T_69643; // @[Modules.scala 56:109:@18261.4]
  wire [10:0] _T_69644; // @[Modules.scala 56:109:@18262.4]
  wire [10:0] buffer_4_703; // @[Modules.scala 56:109:@18263.4]
  wire [11:0] _T_69646; // @[Modules.scala 56:109:@18265.4]
  wire [10:0] _T_69647; // @[Modules.scala 56:109:@18266.4]
  wire [10:0] buffer_4_704; // @[Modules.scala 56:109:@18267.4]
  wire [11:0] _T_69649; // @[Modules.scala 56:109:@18269.4]
  wire [10:0] _T_69650; // @[Modules.scala 56:109:@18270.4]
  wire [10:0] buffer_4_705; // @[Modules.scala 56:109:@18271.4]
  wire [11:0] _T_69652; // @[Modules.scala 56:109:@18273.4]
  wire [10:0] _T_69653; // @[Modules.scala 56:109:@18274.4]
  wire [10:0] buffer_4_706; // @[Modules.scala 56:109:@18275.4]
  wire [11:0] _T_69655; // @[Modules.scala 56:109:@18277.4]
  wire [10:0] _T_69656; // @[Modules.scala 56:109:@18278.4]
  wire [10:0] buffer_4_707; // @[Modules.scala 56:109:@18279.4]
  wire [11:0] _T_69658; // @[Modules.scala 56:109:@18281.4]
  wire [10:0] _T_69659; // @[Modules.scala 56:109:@18282.4]
  wire [10:0] buffer_4_708; // @[Modules.scala 56:109:@18283.4]
  wire [11:0] _T_69661; // @[Modules.scala 56:109:@18285.4]
  wire [10:0] _T_69662; // @[Modules.scala 56:109:@18286.4]
  wire [10:0] buffer_4_709; // @[Modules.scala 56:109:@18287.4]
  wire [11:0] _T_69664; // @[Modules.scala 56:109:@18289.4]
  wire [10:0] _T_69665; // @[Modules.scala 56:109:@18290.4]
  wire [10:0] buffer_4_710; // @[Modules.scala 56:109:@18291.4]
  wire [11:0] _T_69667; // @[Modules.scala 56:109:@18293.4]
  wire [10:0] _T_69668; // @[Modules.scala 56:109:@18294.4]
  wire [10:0] buffer_4_711; // @[Modules.scala 56:109:@18295.4]
  wire [11:0] _T_69670; // @[Modules.scala 56:109:@18297.4]
  wire [10:0] _T_69671; // @[Modules.scala 56:109:@18298.4]
  wire [10:0] buffer_4_712; // @[Modules.scala 56:109:@18299.4]
  wire [11:0] _T_69673; // @[Modules.scala 56:109:@18301.4]
  wire [10:0] _T_69674; // @[Modules.scala 56:109:@18302.4]
  wire [10:0] buffer_4_713; // @[Modules.scala 56:109:@18303.4]
  wire [11:0] _T_69676; // @[Modules.scala 56:109:@18305.4]
  wire [10:0] _T_69677; // @[Modules.scala 56:109:@18306.4]
  wire [10:0] buffer_4_714; // @[Modules.scala 56:109:@18307.4]
  wire [11:0] _T_69679; // @[Modules.scala 56:109:@18309.4]
  wire [10:0] _T_69680; // @[Modules.scala 56:109:@18310.4]
  wire [10:0] buffer_4_715; // @[Modules.scala 56:109:@18311.4]
  wire [11:0] _T_69682; // @[Modules.scala 56:109:@18313.4]
  wire [10:0] _T_69683; // @[Modules.scala 56:109:@18314.4]
  wire [10:0] buffer_4_716; // @[Modules.scala 56:109:@18315.4]
  wire [11:0] _T_69685; // @[Modules.scala 56:109:@18317.4]
  wire [10:0] _T_69686; // @[Modules.scala 56:109:@18318.4]
  wire [10:0] buffer_4_717; // @[Modules.scala 56:109:@18319.4]
  wire [11:0] _T_69688; // @[Modules.scala 56:109:@18321.4]
  wire [10:0] _T_69689; // @[Modules.scala 56:109:@18322.4]
  wire [10:0] buffer_4_718; // @[Modules.scala 56:109:@18323.4]
  wire [11:0] _T_69691; // @[Modules.scala 56:109:@18325.4]
  wire [10:0] _T_69692; // @[Modules.scala 56:109:@18326.4]
  wire [10:0] buffer_4_719; // @[Modules.scala 56:109:@18327.4]
  wire [11:0] _T_69694; // @[Modules.scala 56:109:@18329.4]
  wire [10:0] _T_69695; // @[Modules.scala 56:109:@18330.4]
  wire [10:0] buffer_4_720; // @[Modules.scala 56:109:@18331.4]
  wire [11:0] _T_69697; // @[Modules.scala 56:109:@18333.4]
  wire [10:0] _T_69698; // @[Modules.scala 56:109:@18334.4]
  wire [10:0] buffer_4_721; // @[Modules.scala 56:109:@18335.4]
  wire [11:0] _T_69700; // @[Modules.scala 56:109:@18337.4]
  wire [10:0] _T_69701; // @[Modules.scala 56:109:@18338.4]
  wire [10:0] buffer_4_722; // @[Modules.scala 56:109:@18339.4]
  wire [11:0] _T_69703; // @[Modules.scala 56:109:@18341.4]
  wire [10:0] _T_69704; // @[Modules.scala 56:109:@18342.4]
  wire [10:0] buffer_4_723; // @[Modules.scala 56:109:@18343.4]
  wire [11:0] _T_69706; // @[Modules.scala 56:109:@18345.4]
  wire [10:0] _T_69707; // @[Modules.scala 56:109:@18346.4]
  wire [10:0] buffer_4_724; // @[Modules.scala 56:109:@18347.4]
  wire [11:0] _T_69709; // @[Modules.scala 56:109:@18349.4]
  wire [10:0] _T_69710; // @[Modules.scala 56:109:@18350.4]
  wire [10:0] buffer_4_725; // @[Modules.scala 56:109:@18351.4]
  wire [11:0] _T_69712; // @[Modules.scala 56:109:@18353.4]
  wire [10:0] _T_69713; // @[Modules.scala 56:109:@18354.4]
  wire [10:0] buffer_4_726; // @[Modules.scala 56:109:@18355.4]
  wire [11:0] _T_69715; // @[Modules.scala 56:109:@18357.4]
  wire [10:0] _T_69716; // @[Modules.scala 56:109:@18358.4]
  wire [10:0] buffer_4_727; // @[Modules.scala 56:109:@18359.4]
  wire [11:0] _T_69718; // @[Modules.scala 56:109:@18361.4]
  wire [10:0] _T_69719; // @[Modules.scala 56:109:@18362.4]
  wire [10:0] buffer_4_728; // @[Modules.scala 56:109:@18363.4]
  wire [11:0] _T_69721; // @[Modules.scala 56:109:@18365.4]
  wire [10:0] _T_69722; // @[Modules.scala 56:109:@18366.4]
  wire [10:0] buffer_4_729; // @[Modules.scala 56:109:@18367.4]
  wire [11:0] _T_69724; // @[Modules.scala 56:109:@18369.4]
  wire [10:0] _T_69725; // @[Modules.scala 56:109:@18370.4]
  wire [10:0] buffer_4_730; // @[Modules.scala 56:109:@18371.4]
  wire [11:0] _T_69727; // @[Modules.scala 56:109:@18373.4]
  wire [10:0] _T_69728; // @[Modules.scala 56:109:@18374.4]
  wire [10:0] buffer_4_731; // @[Modules.scala 56:109:@18375.4]
  wire [11:0] _T_69730; // @[Modules.scala 56:109:@18377.4]
  wire [10:0] _T_69731; // @[Modules.scala 56:109:@18378.4]
  wire [10:0] buffer_4_732; // @[Modules.scala 56:109:@18379.4]
  wire [11:0] _T_69733; // @[Modules.scala 56:109:@18381.4]
  wire [10:0] _T_69734; // @[Modules.scala 56:109:@18382.4]
  wire [10:0] buffer_4_733; // @[Modules.scala 56:109:@18383.4]
  wire [11:0] _T_69736; // @[Modules.scala 56:109:@18385.4]
  wire [10:0] _T_69737; // @[Modules.scala 56:109:@18386.4]
  wire [10:0] buffer_4_734; // @[Modules.scala 56:109:@18387.4]
  wire [11:0] _T_69739; // @[Modules.scala 63:156:@18390.4]
  wire [10:0] _T_69740; // @[Modules.scala 63:156:@18391.4]
  wire [10:0] buffer_4_736; // @[Modules.scala 63:156:@18392.4]
  wire [11:0] _T_69742; // @[Modules.scala 63:156:@18394.4]
  wire [10:0] _T_69743; // @[Modules.scala 63:156:@18395.4]
  wire [10:0] buffer_4_737; // @[Modules.scala 63:156:@18396.4]
  wire [11:0] _T_69745; // @[Modules.scala 63:156:@18398.4]
  wire [10:0] _T_69746; // @[Modules.scala 63:156:@18399.4]
  wire [10:0] buffer_4_738; // @[Modules.scala 63:156:@18400.4]
  wire [11:0] _T_69748; // @[Modules.scala 63:156:@18402.4]
  wire [10:0] _T_69749; // @[Modules.scala 63:156:@18403.4]
  wire [10:0] buffer_4_739; // @[Modules.scala 63:156:@18404.4]
  wire [11:0] _T_69751; // @[Modules.scala 63:156:@18406.4]
  wire [10:0] _T_69752; // @[Modules.scala 63:156:@18407.4]
  wire [10:0] buffer_4_740; // @[Modules.scala 63:156:@18408.4]
  wire [11:0] _T_69754; // @[Modules.scala 63:156:@18410.4]
  wire [10:0] _T_69755; // @[Modules.scala 63:156:@18411.4]
  wire [10:0] buffer_4_741; // @[Modules.scala 63:156:@18412.4]
  wire [11:0] _T_69757; // @[Modules.scala 63:156:@18414.4]
  wire [10:0] _T_69758; // @[Modules.scala 63:156:@18415.4]
  wire [10:0] buffer_4_742; // @[Modules.scala 63:156:@18416.4]
  wire [11:0] _T_69760; // @[Modules.scala 63:156:@18418.4]
  wire [10:0] _T_69761; // @[Modules.scala 63:156:@18419.4]
  wire [10:0] buffer_4_743; // @[Modules.scala 63:156:@18420.4]
  wire [11:0] _T_69763; // @[Modules.scala 63:156:@18422.4]
  wire [10:0] _T_69764; // @[Modules.scala 63:156:@18423.4]
  wire [10:0] buffer_4_744; // @[Modules.scala 63:156:@18424.4]
  wire [11:0] _T_69766; // @[Modules.scala 63:156:@18426.4]
  wire [10:0] _T_69767; // @[Modules.scala 63:156:@18427.4]
  wire [10:0] buffer_4_745; // @[Modules.scala 63:156:@18428.4]
  wire [11:0] _T_69769; // @[Modules.scala 63:156:@18430.4]
  wire [10:0] _T_69770; // @[Modules.scala 63:156:@18431.4]
  wire [10:0] buffer_4_746; // @[Modules.scala 63:156:@18432.4]
  wire [11:0] _T_69772; // @[Modules.scala 63:156:@18434.4]
  wire [10:0] _T_69773; // @[Modules.scala 63:156:@18435.4]
  wire [10:0] buffer_4_747; // @[Modules.scala 63:156:@18436.4]
  wire [11:0] _T_69775; // @[Modules.scala 63:156:@18438.4]
  wire [10:0] _T_69776; // @[Modules.scala 63:156:@18439.4]
  wire [10:0] buffer_4_748; // @[Modules.scala 63:156:@18440.4]
  wire [11:0] _T_69778; // @[Modules.scala 63:156:@18442.4]
  wire [10:0] _T_69779; // @[Modules.scala 63:156:@18443.4]
  wire [10:0] buffer_4_749; // @[Modules.scala 63:156:@18444.4]
  wire [11:0] _T_69781; // @[Modules.scala 63:156:@18446.4]
  wire [10:0] _T_69782; // @[Modules.scala 63:156:@18447.4]
  wire [10:0] buffer_4_750; // @[Modules.scala 63:156:@18448.4]
  wire [11:0] _T_69784; // @[Modules.scala 63:156:@18450.4]
  wire [10:0] _T_69785; // @[Modules.scala 63:156:@18451.4]
  wire [10:0] buffer_4_751; // @[Modules.scala 63:156:@18452.4]
  wire [11:0] _T_69787; // @[Modules.scala 63:156:@18454.4]
  wire [10:0] _T_69788; // @[Modules.scala 63:156:@18455.4]
  wire [10:0] buffer_4_752; // @[Modules.scala 63:156:@18456.4]
  wire [11:0] _T_69790; // @[Modules.scala 63:156:@18458.4]
  wire [10:0] _T_69791; // @[Modules.scala 63:156:@18459.4]
  wire [10:0] buffer_4_753; // @[Modules.scala 63:156:@18460.4]
  wire [11:0] _T_69793; // @[Modules.scala 63:156:@18462.4]
  wire [10:0] _T_69794; // @[Modules.scala 63:156:@18463.4]
  wire [10:0] buffer_4_754; // @[Modules.scala 63:156:@18464.4]
  wire [11:0] _T_69796; // @[Modules.scala 63:156:@18466.4]
  wire [10:0] _T_69797; // @[Modules.scala 63:156:@18467.4]
  wire [10:0] buffer_4_755; // @[Modules.scala 63:156:@18468.4]
  wire [11:0] _T_69799; // @[Modules.scala 63:156:@18470.4]
  wire [10:0] _T_69800; // @[Modules.scala 63:156:@18471.4]
  wire [10:0] buffer_4_756; // @[Modules.scala 63:156:@18472.4]
  wire [11:0] _T_69802; // @[Modules.scala 63:156:@18474.4]
  wire [10:0] _T_69803; // @[Modules.scala 63:156:@18475.4]
  wire [10:0] buffer_4_757; // @[Modules.scala 63:156:@18476.4]
  wire [11:0] _T_69805; // @[Modules.scala 63:156:@18478.4]
  wire [10:0] _T_69806; // @[Modules.scala 63:156:@18479.4]
  wire [10:0] buffer_4_758; // @[Modules.scala 63:156:@18480.4]
  wire [11:0] _T_69808; // @[Modules.scala 63:156:@18482.4]
  wire [10:0] _T_69809; // @[Modules.scala 63:156:@18483.4]
  wire [10:0] buffer_4_759; // @[Modules.scala 63:156:@18484.4]
  wire [11:0] _T_69811; // @[Modules.scala 63:156:@18486.4]
  wire [10:0] _T_69812; // @[Modules.scala 63:156:@18487.4]
  wire [10:0] buffer_4_760; // @[Modules.scala 63:156:@18488.4]
  wire [11:0] _T_69814; // @[Modules.scala 63:156:@18490.4]
  wire [10:0] _T_69815; // @[Modules.scala 63:156:@18491.4]
  wire [10:0] buffer_4_761; // @[Modules.scala 63:156:@18492.4]
  wire [11:0] _T_69817; // @[Modules.scala 63:156:@18494.4]
  wire [10:0] _T_69818; // @[Modules.scala 63:156:@18495.4]
  wire [10:0] buffer_4_762; // @[Modules.scala 63:156:@18496.4]
  wire [11:0] _T_69820; // @[Modules.scala 63:156:@18498.4]
  wire [10:0] _T_69821; // @[Modules.scala 63:156:@18499.4]
  wire [10:0] buffer_4_763; // @[Modules.scala 63:156:@18500.4]
  wire [11:0] _T_69823; // @[Modules.scala 63:156:@18502.4]
  wire [10:0] _T_69824; // @[Modules.scala 63:156:@18503.4]
  wire [10:0] buffer_4_764; // @[Modules.scala 63:156:@18504.4]
  wire [11:0] _T_69826; // @[Modules.scala 63:156:@18506.4]
  wire [10:0] _T_69827; // @[Modules.scala 63:156:@18507.4]
  wire [10:0] buffer_4_765; // @[Modules.scala 63:156:@18508.4]
  wire [11:0] _T_69829; // @[Modules.scala 63:156:@18510.4]
  wire [10:0] _T_69830; // @[Modules.scala 63:156:@18511.4]
  wire [10:0] buffer_4_766; // @[Modules.scala 63:156:@18512.4]
  wire [11:0] _T_69832; // @[Modules.scala 63:156:@18514.4]
  wire [10:0] _T_69833; // @[Modules.scala 63:156:@18515.4]
  wire [10:0] buffer_4_767; // @[Modules.scala 63:156:@18516.4]
  wire [11:0] _T_69835; // @[Modules.scala 63:156:@18518.4]
  wire [10:0] _T_69836; // @[Modules.scala 63:156:@18519.4]
  wire [10:0] buffer_4_768; // @[Modules.scala 63:156:@18520.4]
  wire [11:0] _T_69838; // @[Modules.scala 63:156:@18522.4]
  wire [10:0] _T_69839; // @[Modules.scala 63:156:@18523.4]
  wire [10:0] buffer_4_769; // @[Modules.scala 63:156:@18524.4]
  wire [11:0] _T_69841; // @[Modules.scala 63:156:@18526.4]
  wire [10:0] _T_69842; // @[Modules.scala 63:156:@18527.4]
  wire [10:0] buffer_4_770; // @[Modules.scala 63:156:@18528.4]
  wire [11:0] _T_69844; // @[Modules.scala 63:156:@18530.4]
  wire [10:0] _T_69845; // @[Modules.scala 63:156:@18531.4]
  wire [10:0] buffer_4_771; // @[Modules.scala 63:156:@18532.4]
  wire [11:0] _T_69847; // @[Modules.scala 63:156:@18534.4]
  wire [10:0] _T_69848; // @[Modules.scala 63:156:@18535.4]
  wire [10:0] buffer_4_772; // @[Modules.scala 63:156:@18536.4]
  wire [11:0] _T_69850; // @[Modules.scala 63:156:@18538.4]
  wire [10:0] _T_69851; // @[Modules.scala 63:156:@18539.4]
  wire [10:0] buffer_4_773; // @[Modules.scala 63:156:@18540.4]
  wire [11:0] _T_69853; // @[Modules.scala 63:156:@18542.4]
  wire [10:0] _T_69854; // @[Modules.scala 63:156:@18543.4]
  wire [10:0] buffer_4_774; // @[Modules.scala 63:156:@18544.4]
  wire [11:0] _T_69856; // @[Modules.scala 63:156:@18546.4]
  wire [10:0] _T_69857; // @[Modules.scala 63:156:@18547.4]
  wire [10:0] buffer_4_775; // @[Modules.scala 63:156:@18548.4]
  wire [11:0] _T_69859; // @[Modules.scala 63:156:@18550.4]
  wire [10:0] _T_69860; // @[Modules.scala 63:156:@18551.4]
  wire [10:0] buffer_4_776; // @[Modules.scala 63:156:@18552.4]
  wire [11:0] _T_69862; // @[Modules.scala 63:156:@18554.4]
  wire [10:0] _T_69863; // @[Modules.scala 63:156:@18555.4]
  wire [10:0] buffer_4_777; // @[Modules.scala 63:156:@18556.4]
  wire [11:0] _T_69865; // @[Modules.scala 63:156:@18558.4]
  wire [10:0] _T_69866; // @[Modules.scala 63:156:@18559.4]
  wire [10:0] buffer_4_778; // @[Modules.scala 63:156:@18560.4]
  wire [11:0] _T_69868; // @[Modules.scala 63:156:@18562.4]
  wire [10:0] _T_69869; // @[Modules.scala 63:156:@18563.4]
  wire [10:0] buffer_4_779; // @[Modules.scala 63:156:@18564.4]
  wire [11:0] _T_69871; // @[Modules.scala 63:156:@18566.4]
  wire [10:0] _T_69872; // @[Modules.scala 63:156:@18567.4]
  wire [10:0] buffer_4_780; // @[Modules.scala 63:156:@18568.4]
  wire [11:0] _T_69874; // @[Modules.scala 63:156:@18570.4]
  wire [10:0] _T_69875; // @[Modules.scala 63:156:@18571.4]
  wire [10:0] buffer_4_781; // @[Modules.scala 63:156:@18572.4]
  wire [11:0] _T_69877; // @[Modules.scala 63:156:@18574.4]
  wire [10:0] _T_69878; // @[Modules.scala 63:156:@18575.4]
  wire [10:0] buffer_4_782; // @[Modules.scala 63:156:@18576.4]
  wire [11:0] _T_69880; // @[Modules.scala 63:156:@18578.4]
  wire [10:0] _T_69881; // @[Modules.scala 63:156:@18579.4]
  wire [10:0] buffer_4_783; // @[Modules.scala 63:156:@18580.4]
  wire [5:0] _T_69930; // @[Modules.scala 43:37:@18635.4]
  wire [4:0] _T_69931; // @[Modules.scala 43:37:@18636.4]
  wire [4:0] _T_69932; // @[Modules.scala 43:37:@18637.4]
  wire [5:0] _T_69933; // @[Modules.scala 43:47:@18638.4]
  wire [4:0] _T_69934; // @[Modules.scala 43:47:@18639.4]
  wire [4:0] _T_69935; // @[Modules.scala 43:47:@18640.4]
  wire [5:0] _T_69967; // @[Modules.scala 43:47:@18674.4]
  wire [4:0] _T_69968; // @[Modules.scala 43:47:@18675.4]
  wire [4:0] _T_69969; // @[Modules.scala 43:47:@18676.4]
  wire [5:0] _T_70002; // @[Modules.scala 43:47:@18709.4]
  wire [4:0] _T_70003; // @[Modules.scala 43:47:@18710.4]
  wire [4:0] _T_70004; // @[Modules.scala 43:47:@18711.4]
  wire [5:0] _T_70095; // @[Modules.scala 43:47:@18805.4]
  wire [4:0] _T_70096; // @[Modules.scala 43:47:@18806.4]
  wire [4:0] _T_70097; // @[Modules.scala 43:47:@18807.4]
  wire [5:0] _T_70125; // @[Modules.scala 37:46:@18838.4]
  wire [4:0] _T_70126; // @[Modules.scala 37:46:@18839.4]
  wire [4:0] _T_70127; // @[Modules.scala 37:46:@18840.4]
  wire [5:0] _T_70202; // @[Modules.scala 40:46:@18922.4]
  wire [4:0] _T_70203; // @[Modules.scala 40:46:@18923.4]
  wire [4:0] _T_70204; // @[Modules.scala 40:46:@18924.4]
  wire [5:0] _T_70205; // @[Modules.scala 37:46:@18926.4]
  wire [4:0] _T_70206; // @[Modules.scala 37:46:@18927.4]
  wire [4:0] _T_70207; // @[Modules.scala 37:46:@18928.4]
  wire [5:0] _T_70233; // @[Modules.scala 40:46:@18961.4]
  wire [4:0] _T_70234; // @[Modules.scala 40:46:@18962.4]
  wire [4:0] _T_70235; // @[Modules.scala 40:46:@18963.4]
  wire [5:0] _T_70244; // @[Modules.scala 43:37:@18972.4]
  wire [4:0] _T_70245; // @[Modules.scala 43:37:@18973.4]
  wire [4:0] _T_70246; // @[Modules.scala 43:37:@18974.4]
  wire [5:0] _T_70247; // @[Modules.scala 43:47:@18975.4]
  wire [4:0] _T_70248; // @[Modules.scala 43:47:@18976.4]
  wire [4:0] _T_70249; // @[Modules.scala 43:47:@18977.4]
  wire [5:0] _T_70260; // @[Modules.scala 37:46:@18990.4]
  wire [4:0] _T_70261; // @[Modules.scala 37:46:@18991.4]
  wire [4:0] _T_70262; // @[Modules.scala 37:46:@18992.4]
  wire [5:0] _T_70270; // @[Modules.scala 43:47:@19001.4]
  wire [4:0] _T_70271; // @[Modules.scala 43:47:@19002.4]
  wire [4:0] _T_70272; // @[Modules.scala 43:47:@19003.4]
  wire [5:0] _T_70299; // @[Modules.scala 43:47:@19035.4]
  wire [4:0] _T_70300; // @[Modules.scala 43:47:@19036.4]
  wire [4:0] _T_70301; // @[Modules.scala 43:47:@19037.4]
  wire [5:0] _T_70306; // @[Modules.scala 46:47:@19042.4]
  wire [4:0] _T_70307; // @[Modules.scala 46:47:@19043.4]
  wire [4:0] _T_70308; // @[Modules.scala 46:47:@19044.4]
  wire [5:0] _T_70313; // @[Modules.scala 43:47:@19049.4]
  wire [4:0] _T_70314; // @[Modules.scala 43:47:@19050.4]
  wire [4:0] _T_70315; // @[Modules.scala 43:47:@19051.4]
  wire [5:0] _T_70316; // @[Modules.scala 40:46:@19053.4]
  wire [4:0] _T_70317; // @[Modules.scala 40:46:@19054.4]
  wire [4:0] _T_70318; // @[Modules.scala 40:46:@19055.4]
  wire [5:0] _T_70332; // @[Modules.scala 40:46:@19072.4]
  wire [4:0] _T_70333; // @[Modules.scala 40:46:@19073.4]
  wire [4:0] _T_70334; // @[Modules.scala 40:46:@19074.4]
  wire [5:0] _T_70344; // @[Modules.scala 37:46:@19088.4]
  wire [4:0] _T_70345; // @[Modules.scala 37:46:@19089.4]
  wire [4:0] _T_70346; // @[Modules.scala 37:46:@19090.4]
  wire [5:0] _T_70347; // @[Modules.scala 37:46:@19092.4]
  wire [4:0] _T_70348; // @[Modules.scala 37:46:@19093.4]
  wire [4:0] _T_70349; // @[Modules.scala 37:46:@19094.4]
  wire [5:0] _T_70360; // @[Modules.scala 46:47:@19107.4]
  wire [4:0] _T_70361; // @[Modules.scala 46:47:@19108.4]
  wire [4:0] _T_70362; // @[Modules.scala 46:47:@19109.4]
  wire [5:0] _T_70390; // @[Modules.scala 40:46:@19140.4]
  wire [4:0] _T_70391; // @[Modules.scala 40:46:@19141.4]
  wire [4:0] _T_70392; // @[Modules.scala 40:46:@19142.4]
  wire [5:0] _T_70419; // @[Modules.scala 40:46:@19174.4]
  wire [4:0] _T_70420; // @[Modules.scala 40:46:@19175.4]
  wire [4:0] _T_70421; // @[Modules.scala 40:46:@19176.4]
  wire [5:0] _T_70436; // @[Modules.scala 40:46:@19192.4]
  wire [4:0] _T_70437; // @[Modules.scala 40:46:@19193.4]
  wire [4:0] _T_70438; // @[Modules.scala 40:46:@19194.4]
  wire [5:0] _T_70450; // @[Modules.scala 43:47:@19206.4]
  wire [4:0] _T_70451; // @[Modules.scala 43:47:@19207.4]
  wire [4:0] _T_70452; // @[Modules.scala 43:47:@19208.4]
  wire [5:0] _T_70456; // @[Modules.scala 37:46:@19214.4]
  wire [4:0] _T_70457; // @[Modules.scala 37:46:@19215.4]
  wire [4:0] _T_70458; // @[Modules.scala 37:46:@19216.4]
  wire [5:0] _T_70497; // @[Modules.scala 40:46:@19264.4]
  wire [4:0] _T_70498; // @[Modules.scala 40:46:@19265.4]
  wire [4:0] _T_70499; // @[Modules.scala 40:46:@19266.4]
  wire [5:0] _T_70535; // @[Modules.scala 43:47:@19303.4]
  wire [4:0] _T_70536; // @[Modules.scala 43:47:@19304.4]
  wire [4:0] _T_70537; // @[Modules.scala 43:47:@19305.4]
  wire [5:0] _T_70544; // @[Modules.scala 40:46:@19315.4]
  wire [4:0] _T_70545; // @[Modules.scala 40:46:@19316.4]
  wire [4:0] _T_70546; // @[Modules.scala 40:46:@19317.4]
  wire [5:0] _T_70547; // @[Modules.scala 40:46:@19319.4]
  wire [4:0] _T_70548; // @[Modules.scala 40:46:@19320.4]
  wire [4:0] _T_70549; // @[Modules.scala 40:46:@19321.4]
  wire [5:0] _T_70550; // @[Modules.scala 40:46:@19323.4]
  wire [4:0] _T_70551; // @[Modules.scala 40:46:@19324.4]
  wire [4:0] _T_70552; // @[Modules.scala 40:46:@19325.4]
  wire [5:0] _T_70560; // @[Modules.scala 40:46:@19334.4]
  wire [4:0] _T_70561; // @[Modules.scala 40:46:@19335.4]
  wire [4:0] _T_70562; // @[Modules.scala 40:46:@19336.4]
  wire [5:0] _T_70563; // @[Modules.scala 40:46:@19338.4]
  wire [4:0] _T_70564; // @[Modules.scala 40:46:@19339.4]
  wire [4:0] _T_70565; // @[Modules.scala 40:46:@19340.4]
  wire [5:0] _T_70580; // @[Modules.scala 40:46:@19356.4]
  wire [4:0] _T_70581; // @[Modules.scala 40:46:@19357.4]
  wire [4:0] _T_70582; // @[Modules.scala 40:46:@19358.4]
  wire [5:0] _T_70604; // @[Modules.scala 37:46:@19381.4]
  wire [4:0] _T_70605; // @[Modules.scala 37:46:@19382.4]
  wire [4:0] _T_70606; // @[Modules.scala 37:46:@19383.4]
  wire [5:0] _T_70607; // @[Modules.scala 40:46:@19385.4]
  wire [4:0] _T_70608; // @[Modules.scala 40:46:@19386.4]
  wire [4:0] _T_70609; // @[Modules.scala 40:46:@19387.4]
  wire [5:0] _T_70613; // @[Modules.scala 37:46:@19393.4]
  wire [4:0] _T_70614; // @[Modules.scala 37:46:@19394.4]
  wire [4:0] _T_70615; // @[Modules.scala 37:46:@19395.4]
  wire [5:0] _T_70616; // @[Modules.scala 40:46:@19397.4]
  wire [4:0] _T_70617; // @[Modules.scala 40:46:@19398.4]
  wire [4:0] _T_70618; // @[Modules.scala 40:46:@19399.4]
  wire [5:0] _T_70630; // @[Modules.scala 43:47:@19411.4]
  wire [4:0] _T_70631; // @[Modules.scala 43:47:@19412.4]
  wire [4:0] _T_70632; // @[Modules.scala 43:47:@19413.4]
  wire [5:0] _T_70678; // @[Modules.scala 37:46:@19461.4]
  wire [4:0] _T_70679; // @[Modules.scala 37:46:@19462.4]
  wire [4:0] _T_70680; // @[Modules.scala 37:46:@19463.4]
  wire [5:0] _T_70681; // @[Modules.scala 40:46:@19465.4]
  wire [4:0] _T_70682; // @[Modules.scala 40:46:@19466.4]
  wire [4:0] _T_70683; // @[Modules.scala 40:46:@19467.4]
  wire [5:0] _T_70684; // @[Modules.scala 37:46:@19469.4]
  wire [4:0] _T_70685; // @[Modules.scala 37:46:@19470.4]
  wire [4:0] _T_70686; // @[Modules.scala 37:46:@19471.4]
  wire [5:0] _T_70690; // @[Modules.scala 37:46:@19477.4]
  wire [4:0] _T_70691; // @[Modules.scala 37:46:@19478.4]
  wire [4:0] _T_70692; // @[Modules.scala 37:46:@19479.4]
  wire [5:0] _T_70703; // @[Modules.scala 37:46:@19492.4]
  wire [4:0] _T_70704; // @[Modules.scala 37:46:@19493.4]
  wire [4:0] _T_70705; // @[Modules.scala 37:46:@19494.4]
  wire [5:0] _T_70710; // @[Modules.scala 43:47:@19499.4]
  wire [4:0] _T_70711; // @[Modules.scala 43:47:@19500.4]
  wire [4:0] _T_70712; // @[Modules.scala 43:47:@19501.4]
  wire [5:0] _T_70713; // @[Modules.scala 40:46:@19503.4]
  wire [4:0] _T_70714; // @[Modules.scala 40:46:@19504.4]
  wire [4:0] _T_70715; // @[Modules.scala 40:46:@19505.4]
  wire [5:0] _T_70754; // @[Modules.scala 43:47:@19546.4]
  wire [4:0] _T_70755; // @[Modules.scala 43:47:@19547.4]
  wire [4:0] _T_70756; // @[Modules.scala 43:47:@19548.4]
  wire [5:0] _T_70757; // @[Modules.scala 40:46:@19550.4]
  wire [4:0] _T_70758; // @[Modules.scala 40:46:@19551.4]
  wire [4:0] _T_70759; // @[Modules.scala 40:46:@19552.4]
  wire [5:0] _T_70788; // @[Modules.scala 43:47:@19582.4]
  wire [4:0] _T_70789; // @[Modules.scala 43:47:@19583.4]
  wire [4:0] _T_70790; // @[Modules.scala 43:47:@19584.4]
  wire [5:0] _T_70805; // @[Modules.scala 40:46:@19600.4]
  wire [4:0] _T_70806; // @[Modules.scala 40:46:@19601.4]
  wire [4:0] _T_70807; // @[Modules.scala 40:46:@19602.4]
  wire [5:0] _T_70812; // @[Modules.scala 46:47:@19607.4]
  wire [4:0] _T_70813; // @[Modules.scala 46:47:@19608.4]
  wire [4:0] _T_70814; // @[Modules.scala 46:47:@19609.4]
  wire [5:0] _T_70819; // @[Modules.scala 43:47:@19614.4]
  wire [4:0] _T_70820; // @[Modules.scala 43:47:@19615.4]
  wire [4:0] _T_70821; // @[Modules.scala 43:47:@19616.4]
  wire [5:0] _T_70849; // @[Modules.scala 43:47:@19647.4]
  wire [4:0] _T_70850; // @[Modules.scala 43:47:@19648.4]
  wire [4:0] _T_70851; // @[Modules.scala 43:47:@19649.4]
  wire [5:0] _T_70866; // @[Modules.scala 43:47:@19665.4]
  wire [4:0] _T_70867; // @[Modules.scala 43:47:@19666.4]
  wire [4:0] _T_70868; // @[Modules.scala 43:47:@19667.4]
  wire [5:0] _T_70887; // @[Modules.scala 46:47:@19686.4]
  wire [4:0] _T_70888; // @[Modules.scala 46:47:@19687.4]
  wire [4:0] _T_70889; // @[Modules.scala 46:47:@19688.4]
  wire [5:0] _T_70891; // @[Modules.scala 46:37:@19690.4]
  wire [4:0] _T_70892; // @[Modules.scala 46:37:@19691.4]
  wire [4:0] _T_70893; // @[Modules.scala 46:37:@19692.4]
  wire [5:0] _T_70894; // @[Modules.scala 46:47:@19693.4]
  wire [4:0] _T_70895; // @[Modules.scala 46:47:@19694.4]
  wire [4:0] _T_70896; // @[Modules.scala 46:47:@19695.4]
  wire [5:0] _T_70937; // @[Modules.scala 46:47:@19741.4]
  wire [4:0] _T_70938; // @[Modules.scala 46:47:@19742.4]
  wire [4:0] _T_70939; // @[Modules.scala 46:47:@19743.4]
  wire [5:0] _T_70944; // @[Modules.scala 43:47:@19748.4]
  wire [4:0] _T_70945; // @[Modules.scala 43:47:@19749.4]
  wire [4:0] _T_70946; // @[Modules.scala 43:47:@19750.4]
  wire [5:0] _T_70947; // @[Modules.scala 40:46:@19752.4]
  wire [4:0] _T_70948; // @[Modules.scala 40:46:@19753.4]
  wire [4:0] _T_70949; // @[Modules.scala 40:46:@19754.4]
  wire [5:0] _T_70958; // @[Modules.scala 46:37:@19763.4]
  wire [4:0] _T_70959; // @[Modules.scala 46:37:@19764.4]
  wire [4:0] _T_70960; // @[Modules.scala 46:37:@19765.4]
  wire [5:0] _T_70961; // @[Modules.scala 46:47:@19766.4]
  wire [4:0] _T_70962; // @[Modules.scala 46:47:@19767.4]
  wire [4:0] _T_70963; // @[Modules.scala 46:47:@19768.4]
  wire [5:0] _T_70981; // @[Modules.scala 43:47:@19788.4]
  wire [4:0] _T_70982; // @[Modules.scala 43:47:@19789.4]
  wire [4:0] _T_70983; // @[Modules.scala 43:47:@19790.4]
  wire [5:0] _T_71009; // @[Modules.scala 43:47:@19816.4]
  wire [4:0] _T_71010; // @[Modules.scala 43:47:@19817.4]
  wire [4:0] _T_71011; // @[Modules.scala 43:47:@19818.4]
  wire [5:0] _T_71044; // @[Modules.scala 40:46:@19858.4]
  wire [4:0] _T_71045; // @[Modules.scala 40:46:@19859.4]
  wire [4:0] _T_71046; // @[Modules.scala 40:46:@19860.4]
  wire [5:0] _T_71047; // @[Modules.scala 40:46:@19862.4]
  wire [4:0] _T_71048; // @[Modules.scala 40:46:@19863.4]
  wire [4:0] _T_71049; // @[Modules.scala 40:46:@19864.4]
  wire [5:0] _T_71054; // @[Modules.scala 46:47:@19869.4]
  wire [4:0] _T_71055; // @[Modules.scala 46:47:@19870.4]
  wire [4:0] _T_71056; // @[Modules.scala 46:47:@19871.4]
  wire [5:0] _T_71075; // @[Modules.scala 43:47:@19890.4]
  wire [4:0] _T_71076; // @[Modules.scala 43:47:@19891.4]
  wire [4:0] _T_71077; // @[Modules.scala 43:47:@19892.4]
  wire [5:0] _T_71101; // @[Modules.scala 40:46:@19920.4]
  wire [4:0] _T_71102; // @[Modules.scala 40:46:@19921.4]
  wire [4:0] _T_71103; // @[Modules.scala 40:46:@19922.4]
  wire [5:0] _T_71160; // @[Modules.scala 40:46:@19987.4]
  wire [4:0] _T_71161; // @[Modules.scala 40:46:@19988.4]
  wire [4:0] _T_71162; // @[Modules.scala 40:46:@19989.4]
  wire [5:0] _T_71167; // @[Modules.scala 43:47:@19994.4]
  wire [4:0] _T_71168; // @[Modules.scala 43:47:@19995.4]
  wire [4:0] _T_71169; // @[Modules.scala 43:47:@19996.4]
  wire [5:0] _T_71215; // @[Modules.scala 40:46:@20051.4]
  wire [4:0] _T_71216; // @[Modules.scala 40:46:@20052.4]
  wire [4:0] _T_71217; // @[Modules.scala 40:46:@20053.4]
  wire [5:0] _T_71222; // @[Modules.scala 43:47:@20058.4]
  wire [4:0] _T_71223; // @[Modules.scala 43:47:@20059.4]
  wire [4:0] _T_71224; // @[Modules.scala 43:47:@20060.4]
  wire [5:0] _T_71229; // @[Modules.scala 43:47:@20065.4]
  wire [4:0] _T_71230; // @[Modules.scala 43:47:@20066.4]
  wire [4:0] _T_71231; // @[Modules.scala 43:47:@20067.4]
  wire [5:0] _T_71270; // @[Modules.scala 43:47:@20108.4]
  wire [4:0] _T_71271; // @[Modules.scala 43:47:@20109.4]
  wire [4:0] _T_71272; // @[Modules.scala 43:47:@20110.4]
  wire [5:0] _T_71276; // @[Modules.scala 37:46:@20116.4]
  wire [4:0] _T_71277; // @[Modules.scala 37:46:@20117.4]
  wire [4:0] _T_71278; // @[Modules.scala 37:46:@20118.4]
  wire [5:0] _T_71290; // @[Modules.scala 43:47:@20130.4]
  wire [4:0] _T_71291; // @[Modules.scala 43:47:@20131.4]
  wire [4:0] _T_71292; // @[Modules.scala 43:47:@20132.4]
  wire [5:0] _T_71293; // @[Modules.scala 40:46:@20134.4]
  wire [4:0] _T_71294; // @[Modules.scala 40:46:@20135.4]
  wire [4:0] _T_71295; // @[Modules.scala 40:46:@20136.4]
  wire [5:0] _T_71310; // @[Modules.scala 46:47:@20152.4]
  wire [4:0] _T_71311; // @[Modules.scala 46:47:@20153.4]
  wire [4:0] _T_71312; // @[Modules.scala 46:47:@20154.4]
  wire [5:0] _T_71324; // @[Modules.scala 46:47:@20166.4]
  wire [4:0] _T_71325; // @[Modules.scala 46:47:@20167.4]
  wire [4:0] _T_71326; // @[Modules.scala 46:47:@20168.4]
  wire [5:0] _T_71328; // @[Modules.scala 46:37:@20170.4]
  wire [4:0] _T_71329; // @[Modules.scala 46:37:@20171.4]
  wire [4:0] _T_71330; // @[Modules.scala 46:37:@20172.4]
  wire [5:0] _T_71331; // @[Modules.scala 46:47:@20173.4]
  wire [4:0] _T_71332; // @[Modules.scala 46:47:@20174.4]
  wire [4:0] _T_71333; // @[Modules.scala 46:47:@20175.4]
  wire [5:0] _T_71335; // @[Modules.scala 43:37:@20177.4]
  wire [4:0] _T_71336; // @[Modules.scala 43:37:@20178.4]
  wire [4:0] _T_71337; // @[Modules.scala 43:37:@20179.4]
  wire [5:0] _T_71338; // @[Modules.scala 43:47:@20180.4]
  wire [4:0] _T_71339; // @[Modules.scala 43:47:@20181.4]
  wire [4:0] _T_71340; // @[Modules.scala 43:47:@20182.4]
  wire [5:0] _T_71345; // @[Modules.scala 43:47:@20187.4]
  wire [4:0] _T_71346; // @[Modules.scala 43:47:@20188.4]
  wire [4:0] _T_71347; // @[Modules.scala 43:47:@20189.4]
  wire [5:0] _T_71352; // @[Modules.scala 43:47:@20194.4]
  wire [4:0] _T_71353; // @[Modules.scala 43:47:@20195.4]
  wire [4:0] _T_71354; // @[Modules.scala 43:47:@20196.4]
  wire [5:0] _T_71391; // @[Modules.scala 46:47:@20239.4]
  wire [4:0] _T_71392; // @[Modules.scala 46:47:@20240.4]
  wire [4:0] _T_71393; // @[Modules.scala 46:47:@20241.4]
  wire [5:0] _T_71401; // @[Modules.scala 40:46:@20250.4]
  wire [4:0] _T_71402; // @[Modules.scala 40:46:@20251.4]
  wire [4:0] _T_71403; // @[Modules.scala 40:46:@20252.4]
  wire [5:0] _T_71446; // @[Modules.scala 40:46:@20303.4]
  wire [4:0] _T_71447; // @[Modules.scala 40:46:@20304.4]
  wire [4:0] _T_71448; // @[Modules.scala 40:46:@20305.4]
  wire [5:0] _T_71449; // @[Modules.scala 40:46:@20307.4]
  wire [4:0] _T_71450; // @[Modules.scala 40:46:@20308.4]
  wire [4:0] _T_71451; // @[Modules.scala 40:46:@20309.4]
  wire [5:0] _T_71479; // @[Modules.scala 40:46:@20340.4]
  wire [4:0] _T_71480; // @[Modules.scala 40:46:@20341.4]
  wire [4:0] _T_71481; // @[Modules.scala 40:46:@20342.4]
  wire [5:0] _T_71505; // @[Modules.scala 40:46:@20370.4]
  wire [4:0] _T_71506; // @[Modules.scala 40:46:@20371.4]
  wire [4:0] _T_71507; // @[Modules.scala 40:46:@20372.4]
  wire [5:0] _T_71519; // @[Modules.scala 43:47:@20384.4]
  wire [4:0] _T_71520; // @[Modules.scala 43:47:@20385.4]
  wire [4:0] _T_71521; // @[Modules.scala 43:47:@20386.4]
  wire [5:0] _T_71522; // @[Modules.scala 40:46:@20388.4]
  wire [4:0] _T_71523; // @[Modules.scala 40:46:@20389.4]
  wire [4:0] _T_71524; // @[Modules.scala 40:46:@20390.4]
  wire [5:0] _T_71539; // @[Modules.scala 43:47:@20406.4]
  wire [4:0] _T_71540; // @[Modules.scala 43:47:@20407.4]
  wire [4:0] _T_71541; // @[Modules.scala 43:47:@20408.4]
  wire [5:0] _T_71568; // @[Modules.scala 40:46:@20440.4]
  wire [4:0] _T_71569; // @[Modules.scala 40:46:@20441.4]
  wire [4:0] _T_71570; // @[Modules.scala 40:46:@20442.4]
  wire [5:0] _T_71571; // @[Modules.scala 40:46:@20444.4]
  wire [4:0] _T_71572; // @[Modules.scala 40:46:@20445.4]
  wire [4:0] _T_71573; // @[Modules.scala 40:46:@20446.4]
  wire [5:0] _T_71578; // @[Modules.scala 43:47:@20451.4]
  wire [4:0] _T_71579; // @[Modules.scala 43:47:@20452.4]
  wire [4:0] _T_71580; // @[Modules.scala 43:47:@20453.4]
  wire [5:0] _T_71592; // @[Modules.scala 43:47:@20465.4]
  wire [4:0] _T_71593; // @[Modules.scala 43:47:@20466.4]
  wire [4:0] _T_71594; // @[Modules.scala 43:47:@20467.4]
  wire [5:0] _T_71613; // @[Modules.scala 40:46:@20493.4]
  wire [4:0] _T_71614; // @[Modules.scala 40:46:@20494.4]
  wire [4:0] _T_71615; // @[Modules.scala 40:46:@20495.4]
  wire [5:0] _T_71620; // @[Modules.scala 46:47:@20500.4]
  wire [4:0] _T_71621; // @[Modules.scala 46:47:@20501.4]
  wire [4:0] _T_71622; // @[Modules.scala 46:47:@20502.4]
  wire [5:0] _T_71627; // @[Modules.scala 43:47:@20507.4]
  wire [4:0] _T_71628; // @[Modules.scala 43:47:@20508.4]
  wire [4:0] _T_71629; // @[Modules.scala 43:47:@20509.4]
  wire [5:0] _T_71654; // @[Modules.scala 40:46:@20543.4]
  wire [4:0] _T_71655; // @[Modules.scala 40:46:@20544.4]
  wire [4:0] _T_71656; // @[Modules.scala 40:46:@20545.4]
  wire [5:0] _T_71676; // @[Modules.scala 40:46:@20570.4]
  wire [4:0] _T_71677; // @[Modules.scala 40:46:@20571.4]
  wire [4:0] _T_71678; // @[Modules.scala 40:46:@20572.4]
  wire [5:0] _T_71688; // @[Modules.scala 37:46:@20586.4]
  wire [4:0] _T_71689; // @[Modules.scala 37:46:@20587.4]
  wire [4:0] _T_71690; // @[Modules.scala 37:46:@20588.4]
  wire [5:0] _T_71700; // @[Modules.scala 37:46:@20602.4]
  wire [4:0] _T_71701; // @[Modules.scala 37:46:@20603.4]
  wire [4:0] _T_71702; // @[Modules.scala 37:46:@20604.4]
  wire [5:0] _T_71720; // @[Modules.scala 46:37:@20625.4]
  wire [4:0] _T_71721; // @[Modules.scala 46:37:@20626.4]
  wire [4:0] _T_71722; // @[Modules.scala 46:37:@20627.4]
  wire [5:0] _T_71723; // @[Modules.scala 46:47:@20628.4]
  wire [4:0] _T_71724; // @[Modules.scala 46:47:@20629.4]
  wire [4:0] _T_71725; // @[Modules.scala 46:47:@20630.4]
  wire [5:0] _T_71740; // @[Modules.scala 40:46:@20646.4]
  wire [4:0] _T_71741; // @[Modules.scala 40:46:@20647.4]
  wire [4:0] _T_71742; // @[Modules.scala 40:46:@20648.4]
  wire [5:0] _T_71758; // @[Modules.scala 37:46:@20670.4]
  wire [4:0] _T_71759; // @[Modules.scala 37:46:@20671.4]
  wire [4:0] _T_71760; // @[Modules.scala 37:46:@20672.4]
  wire [11:0] _T_71767; // @[Modules.scala 50:57:@20682.4]
  wire [10:0] _T_71768; // @[Modules.scala 50:57:@20683.4]
  wire [10:0] buffer_5_392; // @[Modules.scala 50:57:@20684.4]
  wire [11:0] _T_71770; // @[Modules.scala 50:57:@20686.4]
  wire [10:0] _T_71771; // @[Modules.scala 50:57:@20687.4]
  wire [10:0] buffer_5_393; // @[Modules.scala 50:57:@20688.4]
  wire [11:0] _T_71773; // @[Modules.scala 50:57:@20690.4]
  wire [10:0] _T_71774; // @[Modules.scala 50:57:@20691.4]
  wire [10:0] buffer_5_394; // @[Modules.scala 50:57:@20692.4]
  wire [10:0] buffer_5_10; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71782; // @[Modules.scala 50:57:@20702.4]
  wire [10:0] _T_71783; // @[Modules.scala 50:57:@20703.4]
  wire [10:0] buffer_5_397; // @[Modules.scala 50:57:@20704.4]
  wire [11:0] _T_71788; // @[Modules.scala 50:57:@20710.4]
  wire [10:0] _T_71789; // @[Modules.scala 50:57:@20711.4]
  wire [10:0] buffer_5_399; // @[Modules.scala 50:57:@20712.4]
  wire [10:0] buffer_5_16; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71791; // @[Modules.scala 50:57:@20714.4]
  wire [10:0] _T_71792; // @[Modules.scala 50:57:@20715.4]
  wire [10:0] buffer_5_400; // @[Modules.scala 50:57:@20716.4]
  wire [10:0] buffer_5_21; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71797; // @[Modules.scala 50:57:@20722.4]
  wire [10:0] _T_71798; // @[Modules.scala 50:57:@20723.4]
  wire [10:0] buffer_5_402; // @[Modules.scala 50:57:@20724.4]
  wire [11:0] _T_71809; // @[Modules.scala 50:57:@20738.4]
  wire [10:0] _T_71810; // @[Modules.scala 50:57:@20739.4]
  wire [10:0] buffer_5_406; // @[Modules.scala 50:57:@20740.4]
  wire [11:0] _T_71818; // @[Modules.scala 50:57:@20750.4]
  wire [10:0] _T_71819; // @[Modules.scala 50:57:@20751.4]
  wire [10:0] buffer_5_409; // @[Modules.scala 50:57:@20752.4]
  wire [10:0] buffer_5_36; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71821; // @[Modules.scala 50:57:@20754.4]
  wire [10:0] _T_71822; // @[Modules.scala 50:57:@20755.4]
  wire [10:0] buffer_5_410; // @[Modules.scala 50:57:@20756.4]
  wire [11:0] _T_71827; // @[Modules.scala 50:57:@20762.4]
  wire [10:0] _T_71828; // @[Modules.scala 50:57:@20763.4]
  wire [10:0] buffer_5_412; // @[Modules.scala 50:57:@20764.4]
  wire [10:0] buffer_5_42; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71830; // @[Modules.scala 50:57:@20766.4]
  wire [10:0] _T_71831; // @[Modules.scala 50:57:@20767.4]
  wire [10:0] buffer_5_413; // @[Modules.scala 50:57:@20768.4]
  wire [11:0] _T_71842; // @[Modules.scala 50:57:@20782.4]
  wire [10:0] _T_71843; // @[Modules.scala 50:57:@20783.4]
  wire [10:0] buffer_5_417; // @[Modules.scala 50:57:@20784.4]
  wire [11:0] _T_71848; // @[Modules.scala 50:57:@20790.4]
  wire [10:0] _T_71849; // @[Modules.scala 50:57:@20791.4]
  wire [10:0] buffer_5_419; // @[Modules.scala 50:57:@20792.4]
  wire [10:0] buffer_5_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71851; // @[Modules.scala 50:57:@20794.4]
  wire [10:0] _T_71852; // @[Modules.scala 50:57:@20795.4]
  wire [10:0] buffer_5_420; // @[Modules.scala 50:57:@20796.4]
  wire [10:0] buffer_5_58; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71854; // @[Modules.scala 50:57:@20798.4]
  wire [10:0] _T_71855; // @[Modules.scala 50:57:@20799.4]
  wire [10:0] buffer_5_421; // @[Modules.scala 50:57:@20800.4]
  wire [11:0] _T_71863; // @[Modules.scala 50:57:@20810.4]
  wire [10:0] _T_71864; // @[Modules.scala 50:57:@20811.4]
  wire [10:0] buffer_5_424; // @[Modules.scala 50:57:@20812.4]
  wire [10:0] buffer_5_66; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71866; // @[Modules.scala 50:57:@20814.4]
  wire [10:0] _T_71867; // @[Modules.scala 50:57:@20815.4]
  wire [10:0] buffer_5_425; // @[Modules.scala 50:57:@20816.4]
  wire [10:0] buffer_5_68; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71869; // @[Modules.scala 50:57:@20818.4]
  wire [10:0] _T_71870; // @[Modules.scala 50:57:@20819.4]
  wire [10:0] buffer_5_426; // @[Modules.scala 50:57:@20820.4]
  wire [10:0] buffer_5_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71872; // @[Modules.scala 50:57:@20822.4]
  wire [10:0] _T_71873; // @[Modules.scala 50:57:@20823.4]
  wire [10:0] buffer_5_427; // @[Modules.scala 50:57:@20824.4]
  wire [10:0] buffer_5_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71875; // @[Modules.scala 50:57:@20826.4]
  wire [10:0] _T_71876; // @[Modules.scala 50:57:@20827.4]
  wire [10:0] buffer_5_428; // @[Modules.scala 50:57:@20828.4]
  wire [10:0] buffer_5_80; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_81; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71887; // @[Modules.scala 50:57:@20842.4]
  wire [10:0] _T_71888; // @[Modules.scala 50:57:@20843.4]
  wire [10:0] buffer_5_432; // @[Modules.scala 50:57:@20844.4]
  wire [10:0] buffer_5_82; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71890; // @[Modules.scala 50:57:@20846.4]
  wire [10:0] _T_71891; // @[Modules.scala 50:57:@20847.4]
  wire [10:0] buffer_5_433; // @[Modules.scala 50:57:@20848.4]
  wire [11:0] _T_71893; // @[Modules.scala 50:57:@20850.4]
  wire [10:0] _T_71894; // @[Modules.scala 50:57:@20851.4]
  wire [10:0] buffer_5_434; // @[Modules.scala 50:57:@20852.4]
  wire [10:0] buffer_5_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71896; // @[Modules.scala 50:57:@20854.4]
  wire [10:0] _T_71897; // @[Modules.scala 50:57:@20855.4]
  wire [10:0] buffer_5_435; // @[Modules.scala 50:57:@20856.4]
  wire [10:0] buffer_5_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71902; // @[Modules.scala 50:57:@20862.4]
  wire [10:0] _T_71903; // @[Modules.scala 50:57:@20863.4]
  wire [10:0] buffer_5_437; // @[Modules.scala 50:57:@20864.4]
  wire [10:0] buffer_5_92; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71905; // @[Modules.scala 50:57:@20866.4]
  wire [10:0] _T_71906; // @[Modules.scala 50:57:@20867.4]
  wire [10:0] buffer_5_438; // @[Modules.scala 50:57:@20868.4]
  wire [10:0] buffer_5_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71908; // @[Modules.scala 50:57:@20870.4]
  wire [10:0] _T_71909; // @[Modules.scala 50:57:@20871.4]
  wire [10:0] buffer_5_439; // @[Modules.scala 50:57:@20872.4]
  wire [11:0] _T_71911; // @[Modules.scala 50:57:@20874.4]
  wire [10:0] _T_71912; // @[Modules.scala 50:57:@20875.4]
  wire [10:0] buffer_5_440; // @[Modules.scala 50:57:@20876.4]
  wire [10:0] buffer_5_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71917; // @[Modules.scala 50:57:@20882.4]
  wire [10:0] _T_71918; // @[Modules.scala 50:57:@20883.4]
  wire [10:0] buffer_5_442; // @[Modules.scala 50:57:@20884.4]
  wire [11:0] _T_71920; // @[Modules.scala 50:57:@20886.4]
  wire [10:0] _T_71921; // @[Modules.scala 50:57:@20887.4]
  wire [10:0] buffer_5_443; // @[Modules.scala 50:57:@20888.4]
  wire [11:0] _T_71923; // @[Modules.scala 50:57:@20890.4]
  wire [10:0] _T_71924; // @[Modules.scala 50:57:@20891.4]
  wire [10:0] buffer_5_444; // @[Modules.scala 50:57:@20892.4]
  wire [11:0] _T_71926; // @[Modules.scala 50:57:@20894.4]
  wire [10:0] _T_71927; // @[Modules.scala 50:57:@20895.4]
  wire [10:0] buffer_5_445; // @[Modules.scala 50:57:@20896.4]
  wire [10:0] buffer_5_108; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71929; // @[Modules.scala 50:57:@20898.4]
  wire [10:0] _T_71930; // @[Modules.scala 50:57:@20899.4]
  wire [10:0] buffer_5_446; // @[Modules.scala 50:57:@20900.4]
  wire [10:0] buffer_5_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71932; // @[Modules.scala 50:57:@20902.4]
  wire [10:0] _T_71933; // @[Modules.scala 50:57:@20903.4]
  wire [10:0] buffer_5_447; // @[Modules.scala 50:57:@20904.4]
  wire [10:0] buffer_5_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71935; // @[Modules.scala 50:57:@20906.4]
  wire [10:0] _T_71936; // @[Modules.scala 50:57:@20907.4]
  wire [10:0] buffer_5_448; // @[Modules.scala 50:57:@20908.4]
  wire [10:0] buffer_5_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71938; // @[Modules.scala 50:57:@20910.4]
  wire [10:0] _T_71939; // @[Modules.scala 50:57:@20911.4]
  wire [10:0] buffer_5_449; // @[Modules.scala 50:57:@20912.4]
  wire [11:0] _T_71950; // @[Modules.scala 50:57:@20926.4]
  wire [10:0] _T_71951; // @[Modules.scala 50:57:@20927.4]
  wire [10:0] buffer_5_453; // @[Modules.scala 50:57:@20928.4]
  wire [11:0] _T_71953; // @[Modules.scala 50:57:@20930.4]
  wire [10:0] _T_71954; // @[Modules.scala 50:57:@20931.4]
  wire [10:0] buffer_5_454; // @[Modules.scala 50:57:@20932.4]
  wire [10:0] buffer_5_126; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71956; // @[Modules.scala 50:57:@20934.4]
  wire [10:0] _T_71957; // @[Modules.scala 50:57:@20935.4]
  wire [10:0] buffer_5_455; // @[Modules.scala 50:57:@20936.4]
  wire [11:0] _T_71962; // @[Modules.scala 50:57:@20942.4]
  wire [10:0] _T_71963; // @[Modules.scala 50:57:@20943.4]
  wire [10:0] buffer_5_457; // @[Modules.scala 50:57:@20944.4]
  wire [10:0] buffer_5_132; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71965; // @[Modules.scala 50:57:@20946.4]
  wire [10:0] _T_71966; // @[Modules.scala 50:57:@20947.4]
  wire [10:0] buffer_5_458; // @[Modules.scala 50:57:@20948.4]
  wire [10:0] buffer_5_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71968; // @[Modules.scala 50:57:@20950.4]
  wire [10:0] _T_71969; // @[Modules.scala 50:57:@20951.4]
  wire [10:0] buffer_5_459; // @[Modules.scala 50:57:@20952.4]
  wire [10:0] buffer_5_136; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71971; // @[Modules.scala 50:57:@20954.4]
  wire [10:0] _T_71972; // @[Modules.scala 50:57:@20955.4]
  wire [10:0] buffer_5_460; // @[Modules.scala 50:57:@20956.4]
  wire [10:0] buffer_5_139; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71974; // @[Modules.scala 50:57:@20958.4]
  wire [10:0] _T_71975; // @[Modules.scala 50:57:@20959.4]
  wire [10:0] buffer_5_461; // @[Modules.scala 50:57:@20960.4]
  wire [10:0] buffer_5_140; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71977; // @[Modules.scala 50:57:@20962.4]
  wire [10:0] _T_71978; // @[Modules.scala 50:57:@20963.4]
  wire [10:0] buffer_5_462; // @[Modules.scala 50:57:@20964.4]
  wire [10:0] buffer_5_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71980; // @[Modules.scala 50:57:@20966.4]
  wire [10:0] _T_71981; // @[Modules.scala 50:57:@20967.4]
  wire [10:0] buffer_5_463; // @[Modules.scala 50:57:@20968.4]
  wire [10:0] buffer_5_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71986; // @[Modules.scala 50:57:@20974.4]
  wire [10:0] _T_71987; // @[Modules.scala 50:57:@20975.4]
  wire [10:0] buffer_5_465; // @[Modules.scala 50:57:@20976.4]
  wire [10:0] buffer_5_148; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71989; // @[Modules.scala 50:57:@20978.4]
  wire [10:0] _T_71990; // @[Modules.scala 50:57:@20979.4]
  wire [10:0] buffer_5_466; // @[Modules.scala 50:57:@20980.4]
  wire [10:0] buffer_5_150; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71992; // @[Modules.scala 50:57:@20982.4]
  wire [10:0] _T_71993; // @[Modules.scala 50:57:@20983.4]
  wire [10:0] buffer_5_467; // @[Modules.scala 50:57:@20984.4]
  wire [10:0] buffer_5_153; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_71995; // @[Modules.scala 50:57:@20986.4]
  wire [10:0] _T_71996; // @[Modules.scala 50:57:@20987.4]
  wire [10:0] buffer_5_468; // @[Modules.scala 50:57:@20988.4]
  wire [11:0] _T_71998; // @[Modules.scala 50:57:@20990.4]
  wire [10:0] _T_71999; // @[Modules.scala 50:57:@20991.4]
  wire [10:0] buffer_5_469; // @[Modules.scala 50:57:@20992.4]
  wire [10:0] buffer_5_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72007; // @[Modules.scala 50:57:@21002.4]
  wire [10:0] _T_72008; // @[Modules.scala 50:57:@21003.4]
  wire [10:0] buffer_5_472; // @[Modules.scala 50:57:@21004.4]
  wire [10:0] buffer_5_162; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_163; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72010; // @[Modules.scala 50:57:@21006.4]
  wire [10:0] _T_72011; // @[Modules.scala 50:57:@21007.4]
  wire [10:0] buffer_5_473; // @[Modules.scala 50:57:@21008.4]
  wire [10:0] buffer_5_165; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72013; // @[Modules.scala 50:57:@21010.4]
  wire [10:0] _T_72014; // @[Modules.scala 50:57:@21011.4]
  wire [10:0] buffer_5_474; // @[Modules.scala 50:57:@21012.4]
  wire [10:0] buffer_5_168; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72019; // @[Modules.scala 50:57:@21018.4]
  wire [10:0] _T_72020; // @[Modules.scala 50:57:@21019.4]
  wire [10:0] buffer_5_476; // @[Modules.scala 50:57:@21020.4]
  wire [10:0] buffer_5_170; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72022; // @[Modules.scala 50:57:@21022.4]
  wire [10:0] _T_72023; // @[Modules.scala 50:57:@21023.4]
  wire [10:0] buffer_5_477; // @[Modules.scala 50:57:@21024.4]
  wire [11:0] _T_72028; // @[Modules.scala 50:57:@21030.4]
  wire [10:0] _T_72029; // @[Modules.scala 50:57:@21031.4]
  wire [10:0] buffer_5_479; // @[Modules.scala 50:57:@21032.4]
  wire [10:0] buffer_5_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72031; // @[Modules.scala 50:57:@21034.4]
  wire [10:0] _T_72032; // @[Modules.scala 50:57:@21035.4]
  wire [10:0] buffer_5_480; // @[Modules.scala 50:57:@21036.4]
  wire [10:0] buffer_5_178; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72034; // @[Modules.scala 50:57:@21038.4]
  wire [10:0] _T_72035; // @[Modules.scala 50:57:@21039.4]
  wire [10:0] buffer_5_481; // @[Modules.scala 50:57:@21040.4]
  wire [10:0] buffer_5_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72040; // @[Modules.scala 50:57:@21046.4]
  wire [10:0] _T_72041; // @[Modules.scala 50:57:@21047.4]
  wire [10:0] buffer_5_483; // @[Modules.scala 50:57:@21048.4]
  wire [10:0] buffer_5_186; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_187; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72046; // @[Modules.scala 50:57:@21054.4]
  wire [10:0] _T_72047; // @[Modules.scala 50:57:@21055.4]
  wire [10:0] buffer_5_485; // @[Modules.scala 50:57:@21056.4]
  wire [10:0] buffer_5_188; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72049; // @[Modules.scala 50:57:@21058.4]
  wire [10:0] _T_72050; // @[Modules.scala 50:57:@21059.4]
  wire [10:0] buffer_5_486; // @[Modules.scala 50:57:@21060.4]
  wire [10:0] buffer_5_194; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72058; // @[Modules.scala 50:57:@21070.4]
  wire [10:0] _T_72059; // @[Modules.scala 50:57:@21071.4]
  wire [10:0] buffer_5_489; // @[Modules.scala 50:57:@21072.4]
  wire [10:0] buffer_5_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72061; // @[Modules.scala 50:57:@21074.4]
  wire [10:0] _T_72062; // @[Modules.scala 50:57:@21075.4]
  wire [10:0] buffer_5_490; // @[Modules.scala 50:57:@21076.4]
  wire [10:0] buffer_5_200; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_201; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72067; // @[Modules.scala 50:57:@21082.4]
  wire [10:0] _T_72068; // @[Modules.scala 50:57:@21083.4]
  wire [10:0] buffer_5_492; // @[Modules.scala 50:57:@21084.4]
  wire [11:0] _T_72079; // @[Modules.scala 50:57:@21098.4]
  wire [10:0] _T_72080; // @[Modules.scala 50:57:@21099.4]
  wire [10:0] buffer_5_496; // @[Modules.scala 50:57:@21100.4]
  wire [10:0] buffer_5_210; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72082; // @[Modules.scala 50:57:@21102.4]
  wire [10:0] _T_72083; // @[Modules.scala 50:57:@21103.4]
  wire [10:0] buffer_5_497; // @[Modules.scala 50:57:@21104.4]
  wire [10:0] buffer_5_212; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72085; // @[Modules.scala 50:57:@21106.4]
  wire [10:0] _T_72086; // @[Modules.scala 50:57:@21107.4]
  wire [10:0] buffer_5_498; // @[Modules.scala 50:57:@21108.4]
  wire [10:0] buffer_5_214; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72088; // @[Modules.scala 50:57:@21110.4]
  wire [10:0] _T_72089; // @[Modules.scala 50:57:@21111.4]
  wire [10:0] buffer_5_499; // @[Modules.scala 50:57:@21112.4]
  wire [10:0] buffer_5_218; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72094; // @[Modules.scala 50:57:@21118.4]
  wire [10:0] _T_72095; // @[Modules.scala 50:57:@21119.4]
  wire [10:0] buffer_5_501; // @[Modules.scala 50:57:@21120.4]
  wire [11:0] _T_72097; // @[Modules.scala 50:57:@21122.4]
  wire [10:0] _T_72098; // @[Modules.scala 50:57:@21123.4]
  wire [10:0] buffer_5_502; // @[Modules.scala 50:57:@21124.4]
  wire [10:0] buffer_5_222; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72100; // @[Modules.scala 50:57:@21126.4]
  wire [10:0] _T_72101; // @[Modules.scala 50:57:@21127.4]
  wire [10:0] buffer_5_503; // @[Modules.scala 50:57:@21128.4]
  wire [11:0] _T_72106; // @[Modules.scala 50:57:@21134.4]
  wire [10:0] _T_72107; // @[Modules.scala 50:57:@21135.4]
  wire [10:0] buffer_5_505; // @[Modules.scala 50:57:@21136.4]
  wire [10:0] buffer_5_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72112; // @[Modules.scala 50:57:@21142.4]
  wire [10:0] _T_72113; // @[Modules.scala 50:57:@21143.4]
  wire [10:0] buffer_5_507; // @[Modules.scala 50:57:@21144.4]
  wire [10:0] buffer_5_232; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72115; // @[Modules.scala 50:57:@21146.4]
  wire [10:0] _T_72116; // @[Modules.scala 50:57:@21147.4]
  wire [10:0] buffer_5_508; // @[Modules.scala 50:57:@21148.4]
  wire [11:0] _T_72118; // @[Modules.scala 50:57:@21150.4]
  wire [10:0] _T_72119; // @[Modules.scala 50:57:@21151.4]
  wire [10:0] buffer_5_509; // @[Modules.scala 50:57:@21152.4]
  wire [10:0] buffer_5_236; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72121; // @[Modules.scala 50:57:@21154.4]
  wire [10:0] _T_72122; // @[Modules.scala 50:57:@21155.4]
  wire [10:0] buffer_5_510; // @[Modules.scala 50:57:@21156.4]
  wire [11:0] _T_72127; // @[Modules.scala 50:57:@21162.4]
  wire [10:0] _T_72128; // @[Modules.scala 50:57:@21163.4]
  wire [10:0] buffer_5_512; // @[Modules.scala 50:57:@21164.4]
  wire [10:0] buffer_5_242; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72130; // @[Modules.scala 50:57:@21166.4]
  wire [10:0] _T_72131; // @[Modules.scala 50:57:@21167.4]
  wire [10:0] buffer_5_513; // @[Modules.scala 50:57:@21168.4]
  wire [11:0] _T_72136; // @[Modules.scala 50:57:@21174.4]
  wire [10:0] _T_72137; // @[Modules.scala 50:57:@21175.4]
  wire [10:0] buffer_5_515; // @[Modules.scala 50:57:@21176.4]
  wire [11:0] _T_72139; // @[Modules.scala 50:57:@21178.4]
  wire [10:0] _T_72140; // @[Modules.scala 50:57:@21179.4]
  wire [10:0] buffer_5_516; // @[Modules.scala 50:57:@21180.4]
  wire [10:0] buffer_5_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72148; // @[Modules.scala 50:57:@21190.4]
  wire [10:0] _T_72149; // @[Modules.scala 50:57:@21191.4]
  wire [10:0] buffer_5_519; // @[Modules.scala 50:57:@21192.4]
  wire [10:0] buffer_5_256; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72151; // @[Modules.scala 50:57:@21194.4]
  wire [10:0] _T_72152; // @[Modules.scala 50:57:@21195.4]
  wire [10:0] buffer_5_520; // @[Modules.scala 50:57:@21196.4]
  wire [11:0] _T_72154; // @[Modules.scala 50:57:@21198.4]
  wire [10:0] _T_72155; // @[Modules.scala 50:57:@21199.4]
  wire [10:0] buffer_5_521; // @[Modules.scala 50:57:@21200.4]
  wire [11:0] _T_72157; // @[Modules.scala 50:57:@21202.4]
  wire [10:0] _T_72158; // @[Modules.scala 50:57:@21203.4]
  wire [10:0] buffer_5_522; // @[Modules.scala 50:57:@21204.4]
  wire [10:0] buffer_5_268; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72169; // @[Modules.scala 50:57:@21218.4]
  wire [10:0] _T_72170; // @[Modules.scala 50:57:@21219.4]
  wire [10:0] buffer_5_526; // @[Modules.scala 50:57:@21220.4]
  wire [10:0] buffer_5_270; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72172; // @[Modules.scala 50:57:@21222.4]
  wire [10:0] _T_72173; // @[Modules.scala 50:57:@21223.4]
  wire [10:0] buffer_5_527; // @[Modules.scala 50:57:@21224.4]
  wire [11:0] _T_72175; // @[Modules.scala 50:57:@21226.4]
  wire [10:0] _T_72176; // @[Modules.scala 50:57:@21227.4]
  wire [10:0] buffer_5_528; // @[Modules.scala 50:57:@21228.4]
  wire [11:0] _T_72178; // @[Modules.scala 50:57:@21230.4]
  wire [10:0] _T_72179; // @[Modules.scala 50:57:@21231.4]
  wire [10:0] buffer_5_529; // @[Modules.scala 50:57:@21232.4]
  wire [10:0] buffer_5_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72181; // @[Modules.scala 50:57:@21234.4]
  wire [10:0] _T_72182; // @[Modules.scala 50:57:@21235.4]
  wire [10:0] buffer_5_530; // @[Modules.scala 50:57:@21236.4]
  wire [10:0] buffer_5_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72184; // @[Modules.scala 50:57:@21238.4]
  wire [10:0] _T_72185; // @[Modules.scala 50:57:@21239.4]
  wire [10:0] buffer_5_531; // @[Modules.scala 50:57:@21240.4]
  wire [10:0] buffer_5_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72187; // @[Modules.scala 50:57:@21242.4]
  wire [10:0] _T_72188; // @[Modules.scala 50:57:@21243.4]
  wire [10:0] buffer_5_532; // @[Modules.scala 50:57:@21244.4]
  wire [10:0] buffer_5_282; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72190; // @[Modules.scala 50:57:@21246.4]
  wire [10:0] _T_72191; // @[Modules.scala 50:57:@21247.4]
  wire [10:0] buffer_5_533; // @[Modules.scala 50:57:@21248.4]
  wire [10:0] buffer_5_285; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72193; // @[Modules.scala 50:57:@21250.4]
  wire [10:0] _T_72194; // @[Modules.scala 50:57:@21251.4]
  wire [10:0] buffer_5_534; // @[Modules.scala 50:57:@21252.4]
  wire [10:0] buffer_5_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72196; // @[Modules.scala 50:57:@21254.4]
  wire [10:0] _T_72197; // @[Modules.scala 50:57:@21255.4]
  wire [10:0] buffer_5_535; // @[Modules.scala 50:57:@21256.4]
  wire [10:0] buffer_5_288; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72199; // @[Modules.scala 50:57:@21258.4]
  wire [10:0] _T_72200; // @[Modules.scala 50:57:@21259.4]
  wire [10:0] buffer_5_536; // @[Modules.scala 50:57:@21260.4]
  wire [10:0] buffer_5_290; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72202; // @[Modules.scala 50:57:@21262.4]
  wire [10:0] _T_72203; // @[Modules.scala 50:57:@21263.4]
  wire [10:0] buffer_5_537; // @[Modules.scala 50:57:@21264.4]
  wire [11:0] _T_72214; // @[Modules.scala 50:57:@21278.4]
  wire [10:0] _T_72215; // @[Modules.scala 50:57:@21279.4]
  wire [10:0] buffer_5_541; // @[Modules.scala 50:57:@21280.4]
  wire [10:0] buffer_5_300; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72217; // @[Modules.scala 50:57:@21282.4]
  wire [10:0] _T_72218; // @[Modules.scala 50:57:@21283.4]
  wire [10:0] buffer_5_542; // @[Modules.scala 50:57:@21284.4]
  wire [10:0] buffer_5_302; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72220; // @[Modules.scala 50:57:@21286.4]
  wire [10:0] _T_72221; // @[Modules.scala 50:57:@21287.4]
  wire [10:0] buffer_5_543; // @[Modules.scala 50:57:@21288.4]
  wire [10:0] buffer_5_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72235; // @[Modules.scala 50:57:@21306.4]
  wire [10:0] _T_72236; // @[Modules.scala 50:57:@21307.4]
  wire [10:0] buffer_5_548; // @[Modules.scala 50:57:@21308.4]
  wire [10:0] buffer_5_314; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72238; // @[Modules.scala 50:57:@21310.4]
  wire [10:0] _T_72239; // @[Modules.scala 50:57:@21311.4]
  wire [10:0] buffer_5_549; // @[Modules.scala 50:57:@21312.4]
  wire [11:0] _T_72241; // @[Modules.scala 50:57:@21314.4]
  wire [10:0] _T_72242; // @[Modules.scala 50:57:@21315.4]
  wire [10:0] buffer_5_550; // @[Modules.scala 50:57:@21316.4]
  wire [10:0] buffer_5_320; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72247; // @[Modules.scala 50:57:@21322.4]
  wire [10:0] _T_72248; // @[Modules.scala 50:57:@21323.4]
  wire [10:0] buffer_5_552; // @[Modules.scala 50:57:@21324.4]
  wire [11:0] _T_72253; // @[Modules.scala 50:57:@21330.4]
  wire [10:0] _T_72254; // @[Modules.scala 50:57:@21331.4]
  wire [10:0] buffer_5_554; // @[Modules.scala 50:57:@21332.4]
  wire [10:0] buffer_5_326; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72256; // @[Modules.scala 50:57:@21334.4]
  wire [10:0] _T_72257; // @[Modules.scala 50:57:@21335.4]
  wire [10:0] buffer_5_555; // @[Modules.scala 50:57:@21336.4]
  wire [10:0] buffer_5_328; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72259; // @[Modules.scala 50:57:@21338.4]
  wire [10:0] _T_72260; // @[Modules.scala 50:57:@21339.4]
  wire [10:0] buffer_5_556; // @[Modules.scala 50:57:@21340.4]
  wire [11:0] _T_72262; // @[Modules.scala 50:57:@21342.4]
  wire [10:0] _T_72263; // @[Modules.scala 50:57:@21343.4]
  wire [10:0] buffer_5_557; // @[Modules.scala 50:57:@21344.4]
  wire [10:0] buffer_5_332; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72265; // @[Modules.scala 50:57:@21346.4]
  wire [10:0] _T_72266; // @[Modules.scala 50:57:@21347.4]
  wire [10:0] buffer_5_558; // @[Modules.scala 50:57:@21348.4]
  wire [11:0] _T_72271; // @[Modules.scala 50:57:@21354.4]
  wire [10:0] _T_72272; // @[Modules.scala 50:57:@21355.4]
  wire [10:0] buffer_5_560; // @[Modules.scala 50:57:@21356.4]
  wire [10:0] buffer_5_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72274; // @[Modules.scala 50:57:@21358.4]
  wire [10:0] _T_72275; // @[Modules.scala 50:57:@21359.4]
  wire [10:0] buffer_5_561; // @[Modules.scala 50:57:@21360.4]
  wire [10:0] buffer_5_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72277; // @[Modules.scala 50:57:@21362.4]
  wire [10:0] _T_72278; // @[Modules.scala 50:57:@21363.4]
  wire [10:0] buffer_5_562; // @[Modules.scala 50:57:@21364.4]
  wire [10:0] buffer_5_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72280; // @[Modules.scala 50:57:@21366.4]
  wire [10:0] _T_72281; // @[Modules.scala 50:57:@21367.4]
  wire [10:0] buffer_5_563; // @[Modules.scala 50:57:@21368.4]
  wire [11:0] _T_72289; // @[Modules.scala 50:57:@21378.4]
  wire [10:0] _T_72290; // @[Modules.scala 50:57:@21379.4]
  wire [10:0] buffer_5_566; // @[Modules.scala 50:57:@21380.4]
  wire [10:0] buffer_5_350; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72292; // @[Modules.scala 50:57:@21382.4]
  wire [10:0] _T_72293; // @[Modules.scala 50:57:@21383.4]
  wire [10:0] buffer_5_567; // @[Modules.scala 50:57:@21384.4]
  wire [10:0] buffer_5_352; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72295; // @[Modules.scala 50:57:@21386.4]
  wire [10:0] _T_72296; // @[Modules.scala 50:57:@21387.4]
  wire [10:0] buffer_5_568; // @[Modules.scala 50:57:@21388.4]
  wire [10:0] buffer_5_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72307; // @[Modules.scala 50:57:@21402.4]
  wire [10:0] _T_72308; // @[Modules.scala 50:57:@21403.4]
  wire [10:0] buffer_5_572; // @[Modules.scala 50:57:@21404.4]
  wire [10:0] buffer_5_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72316; // @[Modules.scala 50:57:@21414.4]
  wire [10:0] _T_72317; // @[Modules.scala 50:57:@21415.4]
  wire [10:0] buffer_5_575; // @[Modules.scala 50:57:@21416.4]
  wire [10:0] buffer_5_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72322; // @[Modules.scala 50:57:@21422.4]
  wire [10:0] _T_72323; // @[Modules.scala 50:57:@21423.4]
  wire [10:0] buffer_5_577; // @[Modules.scala 50:57:@21424.4]
  wire [10:0] buffer_5_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72328; // @[Modules.scala 50:57:@21430.4]
  wire [10:0] _T_72329; // @[Modules.scala 50:57:@21431.4]
  wire [10:0] buffer_5_579; // @[Modules.scala 50:57:@21432.4]
  wire [10:0] buffer_5_380; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72337; // @[Modules.scala 50:57:@21442.4]
  wire [10:0] _T_72338; // @[Modules.scala 50:57:@21443.4]
  wire [10:0] buffer_5_582; // @[Modules.scala 50:57:@21444.4]
  wire [10:0] buffer_5_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72340; // @[Modules.scala 50:57:@21446.4]
  wire [10:0] _T_72341; // @[Modules.scala 50:57:@21447.4]
  wire [10:0] buffer_5_583; // @[Modules.scala 50:57:@21448.4]
  wire [10:0] buffer_5_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72349; // @[Modules.scala 50:57:@21458.4]
  wire [10:0] _T_72350; // @[Modules.scala 50:57:@21459.4]
  wire [10:0] buffer_5_586; // @[Modules.scala 50:57:@21460.4]
  wire [11:0] _T_72355; // @[Modules.scala 53:83:@21466.4]
  wire [10:0] _T_72356; // @[Modules.scala 53:83:@21467.4]
  wire [10:0] buffer_5_588; // @[Modules.scala 53:83:@21468.4]
  wire [11:0] _T_72358; // @[Modules.scala 53:83:@21470.4]
  wire [10:0] _T_72359; // @[Modules.scala 53:83:@21471.4]
  wire [10:0] buffer_5_589; // @[Modules.scala 53:83:@21472.4]
  wire [11:0] _T_72361; // @[Modules.scala 53:83:@21474.4]
  wire [10:0] _T_72362; // @[Modules.scala 53:83:@21475.4]
  wire [10:0] buffer_5_590; // @[Modules.scala 53:83:@21476.4]
  wire [11:0] _T_72364; // @[Modules.scala 53:83:@21478.4]
  wire [10:0] _T_72365; // @[Modules.scala 53:83:@21479.4]
  wire [10:0] buffer_5_591; // @[Modules.scala 53:83:@21480.4]
  wire [11:0] _T_72367; // @[Modules.scala 53:83:@21482.4]
  wire [10:0] _T_72368; // @[Modules.scala 53:83:@21483.4]
  wire [10:0] buffer_5_592; // @[Modules.scala 53:83:@21484.4]
  wire [11:0] _T_72370; // @[Modules.scala 53:83:@21486.4]
  wire [10:0] _T_72371; // @[Modules.scala 53:83:@21487.4]
  wire [10:0] buffer_5_593; // @[Modules.scala 53:83:@21488.4]
  wire [11:0] _T_72373; // @[Modules.scala 53:83:@21490.4]
  wire [10:0] _T_72374; // @[Modules.scala 53:83:@21491.4]
  wire [10:0] buffer_5_594; // @[Modules.scala 53:83:@21492.4]
  wire [11:0] _T_72376; // @[Modules.scala 53:83:@21494.4]
  wire [10:0] _T_72377; // @[Modules.scala 53:83:@21495.4]
  wire [10:0] buffer_5_595; // @[Modules.scala 53:83:@21496.4]
  wire [11:0] _T_72379; // @[Modules.scala 53:83:@21498.4]
  wire [10:0] _T_72380; // @[Modules.scala 53:83:@21499.4]
  wire [10:0] buffer_5_596; // @[Modules.scala 53:83:@21500.4]
  wire [11:0] _T_72382; // @[Modules.scala 53:83:@21502.4]
  wire [10:0] _T_72383; // @[Modules.scala 53:83:@21503.4]
  wire [10:0] buffer_5_597; // @[Modules.scala 53:83:@21504.4]
  wire [11:0] _T_72385; // @[Modules.scala 53:83:@21506.4]
  wire [10:0] _T_72386; // @[Modules.scala 53:83:@21507.4]
  wire [10:0] buffer_5_598; // @[Modules.scala 53:83:@21508.4]
  wire [11:0] _T_72391; // @[Modules.scala 53:83:@21514.4]
  wire [10:0] _T_72392; // @[Modules.scala 53:83:@21515.4]
  wire [10:0] buffer_5_600; // @[Modules.scala 53:83:@21516.4]
  wire [11:0] _T_72394; // @[Modules.scala 53:83:@21518.4]
  wire [10:0] _T_72395; // @[Modules.scala 53:83:@21519.4]
  wire [10:0] buffer_5_601; // @[Modules.scala 53:83:@21520.4]
  wire [11:0] _T_72397; // @[Modules.scala 53:83:@21522.4]
  wire [10:0] _T_72398; // @[Modules.scala 53:83:@21523.4]
  wire [10:0] buffer_5_602; // @[Modules.scala 53:83:@21524.4]
  wire [11:0] _T_72403; // @[Modules.scala 53:83:@21530.4]
  wire [10:0] _T_72404; // @[Modules.scala 53:83:@21531.4]
  wire [10:0] buffer_5_604; // @[Modules.scala 53:83:@21532.4]
  wire [11:0] _T_72406; // @[Modules.scala 53:83:@21534.4]
  wire [10:0] _T_72407; // @[Modules.scala 53:83:@21535.4]
  wire [10:0] buffer_5_605; // @[Modules.scala 53:83:@21536.4]
  wire [11:0] _T_72409; // @[Modules.scala 53:83:@21538.4]
  wire [10:0] _T_72410; // @[Modules.scala 53:83:@21539.4]
  wire [10:0] buffer_5_606; // @[Modules.scala 53:83:@21540.4]
  wire [11:0] _T_72412; // @[Modules.scala 53:83:@21542.4]
  wire [10:0] _T_72413; // @[Modules.scala 53:83:@21543.4]
  wire [10:0] buffer_5_607; // @[Modules.scala 53:83:@21544.4]
  wire [11:0] _T_72415; // @[Modules.scala 53:83:@21546.4]
  wire [10:0] _T_72416; // @[Modules.scala 53:83:@21547.4]
  wire [10:0] buffer_5_608; // @[Modules.scala 53:83:@21548.4]
  wire [11:0] _T_72418; // @[Modules.scala 53:83:@21550.4]
  wire [10:0] _T_72419; // @[Modules.scala 53:83:@21551.4]
  wire [10:0] buffer_5_609; // @[Modules.scala 53:83:@21552.4]
  wire [11:0] _T_72421; // @[Modules.scala 53:83:@21554.4]
  wire [10:0] _T_72422; // @[Modules.scala 53:83:@21555.4]
  wire [10:0] buffer_5_610; // @[Modules.scala 53:83:@21556.4]
  wire [11:0] _T_72424; // @[Modules.scala 53:83:@21558.4]
  wire [10:0] _T_72425; // @[Modules.scala 53:83:@21559.4]
  wire [10:0] buffer_5_611; // @[Modules.scala 53:83:@21560.4]
  wire [11:0] _T_72427; // @[Modules.scala 53:83:@21562.4]
  wire [10:0] _T_72428; // @[Modules.scala 53:83:@21563.4]
  wire [10:0] buffer_5_612; // @[Modules.scala 53:83:@21564.4]
  wire [11:0] _T_72430; // @[Modules.scala 53:83:@21566.4]
  wire [10:0] _T_72431; // @[Modules.scala 53:83:@21567.4]
  wire [10:0] buffer_5_613; // @[Modules.scala 53:83:@21568.4]
  wire [11:0] _T_72433; // @[Modules.scala 53:83:@21570.4]
  wire [10:0] _T_72434; // @[Modules.scala 53:83:@21571.4]
  wire [10:0] buffer_5_614; // @[Modules.scala 53:83:@21572.4]
  wire [11:0] _T_72436; // @[Modules.scala 53:83:@21574.4]
  wire [10:0] _T_72437; // @[Modules.scala 53:83:@21575.4]
  wire [10:0] buffer_5_615; // @[Modules.scala 53:83:@21576.4]
  wire [11:0] _T_72439; // @[Modules.scala 53:83:@21578.4]
  wire [10:0] _T_72440; // @[Modules.scala 53:83:@21579.4]
  wire [10:0] buffer_5_616; // @[Modules.scala 53:83:@21580.4]
  wire [11:0] _T_72442; // @[Modules.scala 53:83:@21582.4]
  wire [10:0] _T_72443; // @[Modules.scala 53:83:@21583.4]
  wire [10:0] buffer_5_617; // @[Modules.scala 53:83:@21584.4]
  wire [11:0] _T_72445; // @[Modules.scala 53:83:@21586.4]
  wire [10:0] _T_72446; // @[Modules.scala 53:83:@21587.4]
  wire [10:0] buffer_5_618; // @[Modules.scala 53:83:@21588.4]
  wire [11:0] _T_72448; // @[Modules.scala 53:83:@21590.4]
  wire [10:0] _T_72449; // @[Modules.scala 53:83:@21591.4]
  wire [10:0] buffer_5_619; // @[Modules.scala 53:83:@21592.4]
  wire [11:0] _T_72451; // @[Modules.scala 53:83:@21594.4]
  wire [10:0] _T_72452; // @[Modules.scala 53:83:@21595.4]
  wire [10:0] buffer_5_620; // @[Modules.scala 53:83:@21596.4]
  wire [11:0] _T_72454; // @[Modules.scala 53:83:@21598.4]
  wire [10:0] _T_72455; // @[Modules.scala 53:83:@21599.4]
  wire [10:0] buffer_5_621; // @[Modules.scala 53:83:@21600.4]
  wire [11:0] _T_72457; // @[Modules.scala 53:83:@21602.4]
  wire [10:0] _T_72458; // @[Modules.scala 53:83:@21603.4]
  wire [10:0] buffer_5_622; // @[Modules.scala 53:83:@21604.4]
  wire [11:0] _T_72460; // @[Modules.scala 53:83:@21606.4]
  wire [10:0] _T_72461; // @[Modules.scala 53:83:@21607.4]
  wire [10:0] buffer_5_623; // @[Modules.scala 53:83:@21608.4]
  wire [11:0] _T_72463; // @[Modules.scala 53:83:@21610.4]
  wire [10:0] _T_72464; // @[Modules.scala 53:83:@21611.4]
  wire [10:0] buffer_5_624; // @[Modules.scala 53:83:@21612.4]
  wire [11:0] _T_72466; // @[Modules.scala 53:83:@21614.4]
  wire [10:0] _T_72467; // @[Modules.scala 53:83:@21615.4]
  wire [10:0] buffer_5_625; // @[Modules.scala 53:83:@21616.4]
  wire [11:0] _T_72469; // @[Modules.scala 53:83:@21618.4]
  wire [10:0] _T_72470; // @[Modules.scala 53:83:@21619.4]
  wire [10:0] buffer_5_626; // @[Modules.scala 53:83:@21620.4]
  wire [11:0] _T_72475; // @[Modules.scala 53:83:@21626.4]
  wire [10:0] _T_72476; // @[Modules.scala 53:83:@21627.4]
  wire [10:0] buffer_5_628; // @[Modules.scala 53:83:@21628.4]
  wire [11:0] _T_72478; // @[Modules.scala 53:83:@21630.4]
  wire [10:0] _T_72479; // @[Modules.scala 53:83:@21631.4]
  wire [10:0] buffer_5_629; // @[Modules.scala 53:83:@21632.4]
  wire [11:0] _T_72481; // @[Modules.scala 53:83:@21634.4]
  wire [10:0] _T_72482; // @[Modules.scala 53:83:@21635.4]
  wire [10:0] buffer_5_630; // @[Modules.scala 53:83:@21636.4]
  wire [11:0] _T_72484; // @[Modules.scala 53:83:@21638.4]
  wire [10:0] _T_72485; // @[Modules.scala 53:83:@21639.4]
  wire [10:0] buffer_5_631; // @[Modules.scala 53:83:@21640.4]
  wire [11:0] _T_72487; // @[Modules.scala 53:83:@21642.4]
  wire [10:0] _T_72488; // @[Modules.scala 53:83:@21643.4]
  wire [10:0] buffer_5_632; // @[Modules.scala 53:83:@21644.4]
  wire [11:0] _T_72490; // @[Modules.scala 53:83:@21646.4]
  wire [10:0] _T_72491; // @[Modules.scala 53:83:@21647.4]
  wire [10:0] buffer_5_633; // @[Modules.scala 53:83:@21648.4]
  wire [11:0] _T_72493; // @[Modules.scala 53:83:@21650.4]
  wire [10:0] _T_72494; // @[Modules.scala 53:83:@21651.4]
  wire [10:0] buffer_5_634; // @[Modules.scala 53:83:@21652.4]
  wire [11:0] _T_72496; // @[Modules.scala 53:83:@21654.4]
  wire [10:0] _T_72497; // @[Modules.scala 53:83:@21655.4]
  wire [10:0] buffer_5_635; // @[Modules.scala 53:83:@21656.4]
  wire [11:0] _T_72499; // @[Modules.scala 53:83:@21658.4]
  wire [10:0] _T_72500; // @[Modules.scala 53:83:@21659.4]
  wire [10:0] buffer_5_636; // @[Modules.scala 53:83:@21660.4]
  wire [11:0] _T_72502; // @[Modules.scala 53:83:@21662.4]
  wire [10:0] _T_72503; // @[Modules.scala 53:83:@21663.4]
  wire [10:0] buffer_5_637; // @[Modules.scala 53:83:@21664.4]
  wire [11:0] _T_72505; // @[Modules.scala 53:83:@21666.4]
  wire [10:0] _T_72506; // @[Modules.scala 53:83:@21667.4]
  wire [10:0] buffer_5_638; // @[Modules.scala 53:83:@21668.4]
  wire [11:0] _T_72508; // @[Modules.scala 53:83:@21670.4]
  wire [10:0] _T_72509; // @[Modules.scala 53:83:@21671.4]
  wire [10:0] buffer_5_639; // @[Modules.scala 53:83:@21672.4]
  wire [11:0] _T_72511; // @[Modules.scala 53:83:@21674.4]
  wire [10:0] _T_72512; // @[Modules.scala 53:83:@21675.4]
  wire [10:0] buffer_5_640; // @[Modules.scala 53:83:@21676.4]
  wire [11:0] _T_72514; // @[Modules.scala 53:83:@21678.4]
  wire [10:0] _T_72515; // @[Modules.scala 53:83:@21679.4]
  wire [10:0] buffer_5_641; // @[Modules.scala 53:83:@21680.4]
  wire [11:0] _T_72517; // @[Modules.scala 53:83:@21682.4]
  wire [10:0] _T_72518; // @[Modules.scala 53:83:@21683.4]
  wire [10:0] buffer_5_642; // @[Modules.scala 53:83:@21684.4]
  wire [11:0] _T_72520; // @[Modules.scala 53:83:@21686.4]
  wire [10:0] _T_72521; // @[Modules.scala 53:83:@21687.4]
  wire [10:0] buffer_5_643; // @[Modules.scala 53:83:@21688.4]
  wire [11:0] _T_72523; // @[Modules.scala 53:83:@21690.4]
  wire [10:0] _T_72524; // @[Modules.scala 53:83:@21691.4]
  wire [10:0] buffer_5_644; // @[Modules.scala 53:83:@21692.4]
  wire [11:0] _T_72526; // @[Modules.scala 53:83:@21694.4]
  wire [10:0] _T_72527; // @[Modules.scala 53:83:@21695.4]
  wire [10:0] buffer_5_645; // @[Modules.scala 53:83:@21696.4]
  wire [11:0] _T_72529; // @[Modules.scala 53:83:@21698.4]
  wire [10:0] _T_72530; // @[Modules.scala 53:83:@21699.4]
  wire [10:0] buffer_5_646; // @[Modules.scala 53:83:@21700.4]
  wire [11:0] _T_72532; // @[Modules.scala 53:83:@21702.4]
  wire [10:0] _T_72533; // @[Modules.scala 53:83:@21703.4]
  wire [10:0] buffer_5_647; // @[Modules.scala 53:83:@21704.4]
  wire [11:0] _T_72535; // @[Modules.scala 53:83:@21706.4]
  wire [10:0] _T_72536; // @[Modules.scala 53:83:@21707.4]
  wire [10:0] buffer_5_648; // @[Modules.scala 53:83:@21708.4]
  wire [11:0] _T_72538; // @[Modules.scala 53:83:@21710.4]
  wire [10:0] _T_72539; // @[Modules.scala 53:83:@21711.4]
  wire [10:0] buffer_5_649; // @[Modules.scala 53:83:@21712.4]
  wire [11:0] _T_72541; // @[Modules.scala 53:83:@21714.4]
  wire [10:0] _T_72542; // @[Modules.scala 53:83:@21715.4]
  wire [10:0] buffer_5_650; // @[Modules.scala 53:83:@21716.4]
  wire [11:0] _T_72544; // @[Modules.scala 53:83:@21718.4]
  wire [10:0] _T_72545; // @[Modules.scala 53:83:@21719.4]
  wire [10:0] buffer_5_651; // @[Modules.scala 53:83:@21720.4]
  wire [11:0] _T_72547; // @[Modules.scala 53:83:@21722.4]
  wire [10:0] _T_72548; // @[Modules.scala 53:83:@21723.4]
  wire [10:0] buffer_5_652; // @[Modules.scala 53:83:@21724.4]
  wire [11:0] _T_72550; // @[Modules.scala 53:83:@21726.4]
  wire [10:0] _T_72551; // @[Modules.scala 53:83:@21727.4]
  wire [10:0] buffer_5_653; // @[Modules.scala 53:83:@21728.4]
  wire [11:0] _T_72553; // @[Modules.scala 53:83:@21730.4]
  wire [10:0] _T_72554; // @[Modules.scala 53:83:@21731.4]
  wire [10:0] buffer_5_654; // @[Modules.scala 53:83:@21732.4]
  wire [11:0] _T_72556; // @[Modules.scala 53:83:@21734.4]
  wire [10:0] _T_72557; // @[Modules.scala 53:83:@21735.4]
  wire [10:0] buffer_5_655; // @[Modules.scala 53:83:@21736.4]
  wire [11:0] _T_72559; // @[Modules.scala 53:83:@21738.4]
  wire [10:0] _T_72560; // @[Modules.scala 53:83:@21739.4]
  wire [10:0] buffer_5_656; // @[Modules.scala 53:83:@21740.4]
  wire [11:0] _T_72562; // @[Modules.scala 53:83:@21742.4]
  wire [10:0] _T_72563; // @[Modules.scala 53:83:@21743.4]
  wire [10:0] buffer_5_657; // @[Modules.scala 53:83:@21744.4]
  wire [11:0] _T_72565; // @[Modules.scala 53:83:@21746.4]
  wire [10:0] _T_72566; // @[Modules.scala 53:83:@21747.4]
  wire [10:0] buffer_5_658; // @[Modules.scala 53:83:@21748.4]
  wire [11:0] _T_72568; // @[Modules.scala 53:83:@21750.4]
  wire [10:0] _T_72569; // @[Modules.scala 53:83:@21751.4]
  wire [10:0] buffer_5_659; // @[Modules.scala 53:83:@21752.4]
  wire [11:0] _T_72571; // @[Modules.scala 53:83:@21754.4]
  wire [10:0] _T_72572; // @[Modules.scala 53:83:@21755.4]
  wire [10:0] buffer_5_660; // @[Modules.scala 53:83:@21756.4]
  wire [11:0] _T_72574; // @[Modules.scala 53:83:@21758.4]
  wire [10:0] _T_72575; // @[Modules.scala 53:83:@21759.4]
  wire [10:0] buffer_5_661; // @[Modules.scala 53:83:@21760.4]
  wire [11:0] _T_72577; // @[Modules.scala 53:83:@21762.4]
  wire [10:0] _T_72578; // @[Modules.scala 53:83:@21763.4]
  wire [10:0] buffer_5_662; // @[Modules.scala 53:83:@21764.4]
  wire [11:0] _T_72580; // @[Modules.scala 53:83:@21766.4]
  wire [10:0] _T_72581; // @[Modules.scala 53:83:@21767.4]
  wire [10:0] buffer_5_663; // @[Modules.scala 53:83:@21768.4]
  wire [11:0] _T_72583; // @[Modules.scala 53:83:@21770.4]
  wire [10:0] _T_72584; // @[Modules.scala 53:83:@21771.4]
  wire [10:0] buffer_5_664; // @[Modules.scala 53:83:@21772.4]
  wire [11:0] _T_72586; // @[Modules.scala 53:83:@21774.4]
  wire [10:0] _T_72587; // @[Modules.scala 53:83:@21775.4]
  wire [10:0] buffer_5_665; // @[Modules.scala 53:83:@21776.4]
  wire [11:0] _T_72589; // @[Modules.scala 53:83:@21778.4]
  wire [10:0] _T_72590; // @[Modules.scala 53:83:@21779.4]
  wire [10:0] buffer_5_666; // @[Modules.scala 53:83:@21780.4]
  wire [11:0] _T_72592; // @[Modules.scala 53:83:@21782.4]
  wire [10:0] _T_72593; // @[Modules.scala 53:83:@21783.4]
  wire [10:0] buffer_5_667; // @[Modules.scala 53:83:@21784.4]
  wire [11:0] _T_72595; // @[Modules.scala 53:83:@21786.4]
  wire [10:0] _T_72596; // @[Modules.scala 53:83:@21787.4]
  wire [10:0] buffer_5_668; // @[Modules.scala 53:83:@21788.4]
  wire [11:0] _T_72598; // @[Modules.scala 53:83:@21790.4]
  wire [10:0] _T_72599; // @[Modules.scala 53:83:@21791.4]
  wire [10:0] buffer_5_669; // @[Modules.scala 53:83:@21792.4]
  wire [11:0] _T_72601; // @[Modules.scala 53:83:@21794.4]
  wire [10:0] _T_72602; // @[Modules.scala 53:83:@21795.4]
  wire [10:0] buffer_5_670; // @[Modules.scala 53:83:@21796.4]
  wire [11:0] _T_72604; // @[Modules.scala 53:83:@21798.4]
  wire [10:0] _T_72605; // @[Modules.scala 53:83:@21799.4]
  wire [10:0] buffer_5_671; // @[Modules.scala 53:83:@21800.4]
  wire [11:0] _T_72607; // @[Modules.scala 53:83:@21802.4]
  wire [10:0] _T_72608; // @[Modules.scala 53:83:@21803.4]
  wire [10:0] buffer_5_672; // @[Modules.scala 53:83:@21804.4]
  wire [11:0] _T_72610; // @[Modules.scala 53:83:@21806.4]
  wire [10:0] _T_72611; // @[Modules.scala 53:83:@21807.4]
  wire [10:0] buffer_5_673; // @[Modules.scala 53:83:@21808.4]
  wire [11:0] _T_72616; // @[Modules.scala 53:83:@21814.4]
  wire [10:0] _T_72617; // @[Modules.scala 53:83:@21815.4]
  wire [10:0] buffer_5_675; // @[Modules.scala 53:83:@21816.4]
  wire [11:0] _T_72619; // @[Modules.scala 53:83:@21818.4]
  wire [10:0] _T_72620; // @[Modules.scala 53:83:@21819.4]
  wire [10:0] buffer_5_676; // @[Modules.scala 53:83:@21820.4]
  wire [11:0] _T_72625; // @[Modules.scala 53:83:@21826.4]
  wire [10:0] _T_72626; // @[Modules.scala 53:83:@21827.4]
  wire [10:0] buffer_5_678; // @[Modules.scala 53:83:@21828.4]
  wire [11:0] _T_72628; // @[Modules.scala 53:83:@21830.4]
  wire [10:0] _T_72629; // @[Modules.scala 53:83:@21831.4]
  wire [10:0] buffer_5_679; // @[Modules.scala 53:83:@21832.4]
  wire [11:0] _T_72631; // @[Modules.scala 53:83:@21834.4]
  wire [10:0] _T_72632; // @[Modules.scala 53:83:@21835.4]
  wire [10:0] buffer_5_680; // @[Modules.scala 53:83:@21836.4]
  wire [11:0] _T_72634; // @[Modules.scala 53:83:@21838.4]
  wire [10:0] _T_72635; // @[Modules.scala 53:83:@21839.4]
  wire [10:0] buffer_5_681; // @[Modules.scala 53:83:@21840.4]
  wire [11:0] _T_72637; // @[Modules.scala 53:83:@21842.4]
  wire [10:0] _T_72638; // @[Modules.scala 53:83:@21843.4]
  wire [10:0] buffer_5_682; // @[Modules.scala 53:83:@21844.4]
  wire [11:0] _T_72640; // @[Modules.scala 53:83:@21846.4]
  wire [10:0] _T_72641; // @[Modules.scala 53:83:@21847.4]
  wire [10:0] buffer_5_683; // @[Modules.scala 53:83:@21848.4]
  wire [11:0] _T_72646; // @[Modules.scala 53:83:@21854.4]
  wire [10:0] _T_72647; // @[Modules.scala 53:83:@21855.4]
  wire [10:0] buffer_5_685; // @[Modules.scala 53:83:@21856.4]
  wire [11:0] _T_72649; // @[Modules.scala 56:109:@21858.4]
  wire [10:0] _T_72650; // @[Modules.scala 56:109:@21859.4]
  wire [10:0] buffer_5_686; // @[Modules.scala 56:109:@21860.4]
  wire [11:0] _T_72652; // @[Modules.scala 56:109:@21862.4]
  wire [10:0] _T_72653; // @[Modules.scala 56:109:@21863.4]
  wire [10:0] buffer_5_687; // @[Modules.scala 56:109:@21864.4]
  wire [11:0] _T_72655; // @[Modules.scala 56:109:@21866.4]
  wire [10:0] _T_72656; // @[Modules.scala 56:109:@21867.4]
  wire [10:0] buffer_5_688; // @[Modules.scala 56:109:@21868.4]
  wire [11:0] _T_72658; // @[Modules.scala 56:109:@21870.4]
  wire [10:0] _T_72659; // @[Modules.scala 56:109:@21871.4]
  wire [10:0] buffer_5_689; // @[Modules.scala 56:109:@21872.4]
  wire [11:0] _T_72661; // @[Modules.scala 56:109:@21874.4]
  wire [10:0] _T_72662; // @[Modules.scala 56:109:@21875.4]
  wire [10:0] buffer_5_690; // @[Modules.scala 56:109:@21876.4]
  wire [11:0] _T_72664; // @[Modules.scala 56:109:@21878.4]
  wire [10:0] _T_72665; // @[Modules.scala 56:109:@21879.4]
  wire [10:0] buffer_5_691; // @[Modules.scala 56:109:@21880.4]
  wire [11:0] _T_72667; // @[Modules.scala 56:109:@21882.4]
  wire [10:0] _T_72668; // @[Modules.scala 56:109:@21883.4]
  wire [10:0] buffer_5_692; // @[Modules.scala 56:109:@21884.4]
  wire [11:0] _T_72670; // @[Modules.scala 56:109:@21886.4]
  wire [10:0] _T_72671; // @[Modules.scala 56:109:@21887.4]
  wire [10:0] buffer_5_693; // @[Modules.scala 56:109:@21888.4]
  wire [11:0] _T_72673; // @[Modules.scala 56:109:@21890.4]
  wire [10:0] _T_72674; // @[Modules.scala 56:109:@21891.4]
  wire [10:0] buffer_5_694; // @[Modules.scala 56:109:@21892.4]
  wire [11:0] _T_72676; // @[Modules.scala 56:109:@21894.4]
  wire [10:0] _T_72677; // @[Modules.scala 56:109:@21895.4]
  wire [10:0] buffer_5_695; // @[Modules.scala 56:109:@21896.4]
  wire [11:0] _T_72679; // @[Modules.scala 56:109:@21898.4]
  wire [10:0] _T_72680; // @[Modules.scala 56:109:@21899.4]
  wire [10:0] buffer_5_696; // @[Modules.scala 56:109:@21900.4]
  wire [11:0] _T_72682; // @[Modules.scala 56:109:@21902.4]
  wire [10:0] _T_72683; // @[Modules.scala 56:109:@21903.4]
  wire [10:0] buffer_5_697; // @[Modules.scala 56:109:@21904.4]
  wire [11:0] _T_72685; // @[Modules.scala 56:109:@21906.4]
  wire [10:0] _T_72686; // @[Modules.scala 56:109:@21907.4]
  wire [10:0] buffer_5_698; // @[Modules.scala 56:109:@21908.4]
  wire [11:0] _T_72688; // @[Modules.scala 56:109:@21910.4]
  wire [10:0] _T_72689; // @[Modules.scala 56:109:@21911.4]
  wire [10:0] buffer_5_699; // @[Modules.scala 56:109:@21912.4]
  wire [11:0] _T_72691; // @[Modules.scala 56:109:@21914.4]
  wire [10:0] _T_72692; // @[Modules.scala 56:109:@21915.4]
  wire [10:0] buffer_5_700; // @[Modules.scala 56:109:@21916.4]
  wire [11:0] _T_72694; // @[Modules.scala 56:109:@21918.4]
  wire [10:0] _T_72695; // @[Modules.scala 56:109:@21919.4]
  wire [10:0] buffer_5_701; // @[Modules.scala 56:109:@21920.4]
  wire [11:0] _T_72697; // @[Modules.scala 56:109:@21922.4]
  wire [10:0] _T_72698; // @[Modules.scala 56:109:@21923.4]
  wire [10:0] buffer_5_702; // @[Modules.scala 56:109:@21924.4]
  wire [11:0] _T_72700; // @[Modules.scala 56:109:@21926.4]
  wire [10:0] _T_72701; // @[Modules.scala 56:109:@21927.4]
  wire [10:0] buffer_5_703; // @[Modules.scala 56:109:@21928.4]
  wire [11:0] _T_72703; // @[Modules.scala 56:109:@21930.4]
  wire [10:0] _T_72704; // @[Modules.scala 56:109:@21931.4]
  wire [10:0] buffer_5_704; // @[Modules.scala 56:109:@21932.4]
  wire [11:0] _T_72706; // @[Modules.scala 56:109:@21934.4]
  wire [10:0] _T_72707; // @[Modules.scala 56:109:@21935.4]
  wire [10:0] buffer_5_705; // @[Modules.scala 56:109:@21936.4]
  wire [11:0] _T_72709; // @[Modules.scala 56:109:@21938.4]
  wire [10:0] _T_72710; // @[Modules.scala 56:109:@21939.4]
  wire [10:0] buffer_5_706; // @[Modules.scala 56:109:@21940.4]
  wire [11:0] _T_72712; // @[Modules.scala 56:109:@21942.4]
  wire [10:0] _T_72713; // @[Modules.scala 56:109:@21943.4]
  wire [10:0] buffer_5_707; // @[Modules.scala 56:109:@21944.4]
  wire [11:0] _T_72715; // @[Modules.scala 56:109:@21946.4]
  wire [10:0] _T_72716; // @[Modules.scala 56:109:@21947.4]
  wire [10:0] buffer_5_708; // @[Modules.scala 56:109:@21948.4]
  wire [11:0] _T_72718; // @[Modules.scala 56:109:@21950.4]
  wire [10:0] _T_72719; // @[Modules.scala 56:109:@21951.4]
  wire [10:0] buffer_5_709; // @[Modules.scala 56:109:@21952.4]
  wire [11:0] _T_72721; // @[Modules.scala 56:109:@21954.4]
  wire [10:0] _T_72722; // @[Modules.scala 56:109:@21955.4]
  wire [10:0] buffer_5_710; // @[Modules.scala 56:109:@21956.4]
  wire [11:0] _T_72724; // @[Modules.scala 56:109:@21958.4]
  wire [10:0] _T_72725; // @[Modules.scala 56:109:@21959.4]
  wire [10:0] buffer_5_711; // @[Modules.scala 56:109:@21960.4]
  wire [11:0] _T_72727; // @[Modules.scala 56:109:@21962.4]
  wire [10:0] _T_72728; // @[Modules.scala 56:109:@21963.4]
  wire [10:0] buffer_5_712; // @[Modules.scala 56:109:@21964.4]
  wire [11:0] _T_72730; // @[Modules.scala 56:109:@21966.4]
  wire [10:0] _T_72731; // @[Modules.scala 56:109:@21967.4]
  wire [10:0] buffer_5_713; // @[Modules.scala 56:109:@21968.4]
  wire [11:0] _T_72733; // @[Modules.scala 56:109:@21970.4]
  wire [10:0] _T_72734; // @[Modules.scala 56:109:@21971.4]
  wire [10:0] buffer_5_714; // @[Modules.scala 56:109:@21972.4]
  wire [11:0] _T_72736; // @[Modules.scala 56:109:@21974.4]
  wire [10:0] _T_72737; // @[Modules.scala 56:109:@21975.4]
  wire [10:0] buffer_5_715; // @[Modules.scala 56:109:@21976.4]
  wire [11:0] _T_72739; // @[Modules.scala 56:109:@21978.4]
  wire [10:0] _T_72740; // @[Modules.scala 56:109:@21979.4]
  wire [10:0] buffer_5_716; // @[Modules.scala 56:109:@21980.4]
  wire [11:0] _T_72742; // @[Modules.scala 56:109:@21982.4]
  wire [10:0] _T_72743; // @[Modules.scala 56:109:@21983.4]
  wire [10:0] buffer_5_717; // @[Modules.scala 56:109:@21984.4]
  wire [11:0] _T_72745; // @[Modules.scala 56:109:@21986.4]
  wire [10:0] _T_72746; // @[Modules.scala 56:109:@21987.4]
  wire [10:0] buffer_5_718; // @[Modules.scala 56:109:@21988.4]
  wire [11:0] _T_72748; // @[Modules.scala 56:109:@21990.4]
  wire [10:0] _T_72749; // @[Modules.scala 56:109:@21991.4]
  wire [10:0] buffer_5_719; // @[Modules.scala 56:109:@21992.4]
  wire [11:0] _T_72751; // @[Modules.scala 56:109:@21994.4]
  wire [10:0] _T_72752; // @[Modules.scala 56:109:@21995.4]
  wire [10:0] buffer_5_720; // @[Modules.scala 56:109:@21996.4]
  wire [11:0] _T_72754; // @[Modules.scala 56:109:@21998.4]
  wire [10:0] _T_72755; // @[Modules.scala 56:109:@21999.4]
  wire [10:0] buffer_5_721; // @[Modules.scala 56:109:@22000.4]
  wire [11:0] _T_72757; // @[Modules.scala 56:109:@22002.4]
  wire [10:0] _T_72758; // @[Modules.scala 56:109:@22003.4]
  wire [10:0] buffer_5_722; // @[Modules.scala 56:109:@22004.4]
  wire [11:0] _T_72760; // @[Modules.scala 56:109:@22006.4]
  wire [10:0] _T_72761; // @[Modules.scala 56:109:@22007.4]
  wire [10:0] buffer_5_723; // @[Modules.scala 56:109:@22008.4]
  wire [11:0] _T_72763; // @[Modules.scala 56:109:@22010.4]
  wire [10:0] _T_72764; // @[Modules.scala 56:109:@22011.4]
  wire [10:0] buffer_5_724; // @[Modules.scala 56:109:@22012.4]
  wire [11:0] _T_72766; // @[Modules.scala 56:109:@22014.4]
  wire [10:0] _T_72767; // @[Modules.scala 56:109:@22015.4]
  wire [10:0] buffer_5_725; // @[Modules.scala 56:109:@22016.4]
  wire [11:0] _T_72769; // @[Modules.scala 56:109:@22018.4]
  wire [10:0] _T_72770; // @[Modules.scala 56:109:@22019.4]
  wire [10:0] buffer_5_726; // @[Modules.scala 56:109:@22020.4]
  wire [11:0] _T_72772; // @[Modules.scala 56:109:@22022.4]
  wire [10:0] _T_72773; // @[Modules.scala 56:109:@22023.4]
  wire [10:0] buffer_5_727; // @[Modules.scala 56:109:@22024.4]
  wire [11:0] _T_72775; // @[Modules.scala 56:109:@22026.4]
  wire [10:0] _T_72776; // @[Modules.scala 56:109:@22027.4]
  wire [10:0] buffer_5_728; // @[Modules.scala 56:109:@22028.4]
  wire [11:0] _T_72778; // @[Modules.scala 56:109:@22030.4]
  wire [10:0] _T_72779; // @[Modules.scala 56:109:@22031.4]
  wire [10:0] buffer_5_729; // @[Modules.scala 56:109:@22032.4]
  wire [11:0] _T_72781; // @[Modules.scala 56:109:@22034.4]
  wire [10:0] _T_72782; // @[Modules.scala 56:109:@22035.4]
  wire [10:0] buffer_5_730; // @[Modules.scala 56:109:@22036.4]
  wire [11:0] _T_72784; // @[Modules.scala 56:109:@22038.4]
  wire [10:0] _T_72785; // @[Modules.scala 56:109:@22039.4]
  wire [10:0] buffer_5_731; // @[Modules.scala 56:109:@22040.4]
  wire [11:0] _T_72787; // @[Modules.scala 56:109:@22042.4]
  wire [10:0] _T_72788; // @[Modules.scala 56:109:@22043.4]
  wire [10:0] buffer_5_732; // @[Modules.scala 56:109:@22044.4]
  wire [11:0] _T_72790; // @[Modules.scala 56:109:@22046.4]
  wire [10:0] _T_72791; // @[Modules.scala 56:109:@22047.4]
  wire [10:0] buffer_5_733; // @[Modules.scala 56:109:@22048.4]
  wire [11:0] _T_72793; // @[Modules.scala 56:109:@22050.4]
  wire [10:0] _T_72794; // @[Modules.scala 56:109:@22051.4]
  wire [10:0] buffer_5_734; // @[Modules.scala 56:109:@22052.4]
  wire [11:0] _T_72796; // @[Modules.scala 63:156:@22055.4]
  wire [10:0] _T_72797; // @[Modules.scala 63:156:@22056.4]
  wire [10:0] buffer_5_736; // @[Modules.scala 63:156:@22057.4]
  wire [11:0] _T_72799; // @[Modules.scala 63:156:@22059.4]
  wire [10:0] _T_72800; // @[Modules.scala 63:156:@22060.4]
  wire [10:0] buffer_5_737; // @[Modules.scala 63:156:@22061.4]
  wire [11:0] _T_72802; // @[Modules.scala 63:156:@22063.4]
  wire [10:0] _T_72803; // @[Modules.scala 63:156:@22064.4]
  wire [10:0] buffer_5_738; // @[Modules.scala 63:156:@22065.4]
  wire [11:0] _T_72805; // @[Modules.scala 63:156:@22067.4]
  wire [10:0] _T_72806; // @[Modules.scala 63:156:@22068.4]
  wire [10:0] buffer_5_739; // @[Modules.scala 63:156:@22069.4]
  wire [11:0] _T_72808; // @[Modules.scala 63:156:@22071.4]
  wire [10:0] _T_72809; // @[Modules.scala 63:156:@22072.4]
  wire [10:0] buffer_5_740; // @[Modules.scala 63:156:@22073.4]
  wire [11:0] _T_72811; // @[Modules.scala 63:156:@22075.4]
  wire [10:0] _T_72812; // @[Modules.scala 63:156:@22076.4]
  wire [10:0] buffer_5_741; // @[Modules.scala 63:156:@22077.4]
  wire [11:0] _T_72814; // @[Modules.scala 63:156:@22079.4]
  wire [10:0] _T_72815; // @[Modules.scala 63:156:@22080.4]
  wire [10:0] buffer_5_742; // @[Modules.scala 63:156:@22081.4]
  wire [11:0] _T_72817; // @[Modules.scala 63:156:@22083.4]
  wire [10:0] _T_72818; // @[Modules.scala 63:156:@22084.4]
  wire [10:0] buffer_5_743; // @[Modules.scala 63:156:@22085.4]
  wire [11:0] _T_72820; // @[Modules.scala 63:156:@22087.4]
  wire [10:0] _T_72821; // @[Modules.scala 63:156:@22088.4]
  wire [10:0] buffer_5_744; // @[Modules.scala 63:156:@22089.4]
  wire [11:0] _T_72823; // @[Modules.scala 63:156:@22091.4]
  wire [10:0] _T_72824; // @[Modules.scala 63:156:@22092.4]
  wire [10:0] buffer_5_745; // @[Modules.scala 63:156:@22093.4]
  wire [11:0] _T_72826; // @[Modules.scala 63:156:@22095.4]
  wire [10:0] _T_72827; // @[Modules.scala 63:156:@22096.4]
  wire [10:0] buffer_5_746; // @[Modules.scala 63:156:@22097.4]
  wire [11:0] _T_72829; // @[Modules.scala 63:156:@22099.4]
  wire [10:0] _T_72830; // @[Modules.scala 63:156:@22100.4]
  wire [10:0] buffer_5_747; // @[Modules.scala 63:156:@22101.4]
  wire [11:0] _T_72832; // @[Modules.scala 63:156:@22103.4]
  wire [10:0] _T_72833; // @[Modules.scala 63:156:@22104.4]
  wire [10:0] buffer_5_748; // @[Modules.scala 63:156:@22105.4]
  wire [11:0] _T_72835; // @[Modules.scala 63:156:@22107.4]
  wire [10:0] _T_72836; // @[Modules.scala 63:156:@22108.4]
  wire [10:0] buffer_5_749; // @[Modules.scala 63:156:@22109.4]
  wire [11:0] _T_72838; // @[Modules.scala 63:156:@22111.4]
  wire [10:0] _T_72839; // @[Modules.scala 63:156:@22112.4]
  wire [10:0] buffer_5_750; // @[Modules.scala 63:156:@22113.4]
  wire [11:0] _T_72841; // @[Modules.scala 63:156:@22115.4]
  wire [10:0] _T_72842; // @[Modules.scala 63:156:@22116.4]
  wire [10:0] buffer_5_751; // @[Modules.scala 63:156:@22117.4]
  wire [11:0] _T_72844; // @[Modules.scala 63:156:@22119.4]
  wire [10:0] _T_72845; // @[Modules.scala 63:156:@22120.4]
  wire [10:0] buffer_5_752; // @[Modules.scala 63:156:@22121.4]
  wire [11:0] _T_72847; // @[Modules.scala 63:156:@22123.4]
  wire [10:0] _T_72848; // @[Modules.scala 63:156:@22124.4]
  wire [10:0] buffer_5_753; // @[Modules.scala 63:156:@22125.4]
  wire [11:0] _T_72850; // @[Modules.scala 63:156:@22127.4]
  wire [10:0] _T_72851; // @[Modules.scala 63:156:@22128.4]
  wire [10:0] buffer_5_754; // @[Modules.scala 63:156:@22129.4]
  wire [11:0] _T_72853; // @[Modules.scala 63:156:@22131.4]
  wire [10:0] _T_72854; // @[Modules.scala 63:156:@22132.4]
  wire [10:0] buffer_5_755; // @[Modules.scala 63:156:@22133.4]
  wire [11:0] _T_72856; // @[Modules.scala 63:156:@22135.4]
  wire [10:0] _T_72857; // @[Modules.scala 63:156:@22136.4]
  wire [10:0] buffer_5_756; // @[Modules.scala 63:156:@22137.4]
  wire [11:0] _T_72859; // @[Modules.scala 63:156:@22139.4]
  wire [10:0] _T_72860; // @[Modules.scala 63:156:@22140.4]
  wire [10:0] buffer_5_757; // @[Modules.scala 63:156:@22141.4]
  wire [11:0] _T_72862; // @[Modules.scala 63:156:@22143.4]
  wire [10:0] _T_72863; // @[Modules.scala 63:156:@22144.4]
  wire [10:0] buffer_5_758; // @[Modules.scala 63:156:@22145.4]
  wire [11:0] _T_72865; // @[Modules.scala 63:156:@22147.4]
  wire [10:0] _T_72866; // @[Modules.scala 63:156:@22148.4]
  wire [10:0] buffer_5_759; // @[Modules.scala 63:156:@22149.4]
  wire [11:0] _T_72868; // @[Modules.scala 63:156:@22151.4]
  wire [10:0] _T_72869; // @[Modules.scala 63:156:@22152.4]
  wire [10:0] buffer_5_760; // @[Modules.scala 63:156:@22153.4]
  wire [11:0] _T_72871; // @[Modules.scala 63:156:@22155.4]
  wire [10:0] _T_72872; // @[Modules.scala 63:156:@22156.4]
  wire [10:0] buffer_5_761; // @[Modules.scala 63:156:@22157.4]
  wire [11:0] _T_72874; // @[Modules.scala 63:156:@22159.4]
  wire [10:0] _T_72875; // @[Modules.scala 63:156:@22160.4]
  wire [10:0] buffer_5_762; // @[Modules.scala 63:156:@22161.4]
  wire [11:0] _T_72877; // @[Modules.scala 63:156:@22163.4]
  wire [10:0] _T_72878; // @[Modules.scala 63:156:@22164.4]
  wire [10:0] buffer_5_763; // @[Modules.scala 63:156:@22165.4]
  wire [11:0] _T_72880; // @[Modules.scala 63:156:@22167.4]
  wire [10:0] _T_72881; // @[Modules.scala 63:156:@22168.4]
  wire [10:0] buffer_5_764; // @[Modules.scala 63:156:@22169.4]
  wire [11:0] _T_72883; // @[Modules.scala 63:156:@22171.4]
  wire [10:0] _T_72884; // @[Modules.scala 63:156:@22172.4]
  wire [10:0] buffer_5_765; // @[Modules.scala 63:156:@22173.4]
  wire [11:0] _T_72886; // @[Modules.scala 63:156:@22175.4]
  wire [10:0] _T_72887; // @[Modules.scala 63:156:@22176.4]
  wire [10:0] buffer_5_766; // @[Modules.scala 63:156:@22177.4]
  wire [11:0] _T_72889; // @[Modules.scala 63:156:@22179.4]
  wire [10:0] _T_72890; // @[Modules.scala 63:156:@22180.4]
  wire [10:0] buffer_5_767; // @[Modules.scala 63:156:@22181.4]
  wire [11:0] _T_72892; // @[Modules.scala 63:156:@22183.4]
  wire [10:0] _T_72893; // @[Modules.scala 63:156:@22184.4]
  wire [10:0] buffer_5_768; // @[Modules.scala 63:156:@22185.4]
  wire [11:0] _T_72895; // @[Modules.scala 63:156:@22187.4]
  wire [10:0] _T_72896; // @[Modules.scala 63:156:@22188.4]
  wire [10:0] buffer_5_769; // @[Modules.scala 63:156:@22189.4]
  wire [11:0] _T_72898; // @[Modules.scala 63:156:@22191.4]
  wire [10:0] _T_72899; // @[Modules.scala 63:156:@22192.4]
  wire [10:0] buffer_5_770; // @[Modules.scala 63:156:@22193.4]
  wire [11:0] _T_72901; // @[Modules.scala 63:156:@22195.4]
  wire [10:0] _T_72902; // @[Modules.scala 63:156:@22196.4]
  wire [10:0] buffer_5_771; // @[Modules.scala 63:156:@22197.4]
  wire [11:0] _T_72904; // @[Modules.scala 63:156:@22199.4]
  wire [10:0] _T_72905; // @[Modules.scala 63:156:@22200.4]
  wire [10:0] buffer_5_772; // @[Modules.scala 63:156:@22201.4]
  wire [11:0] _T_72907; // @[Modules.scala 63:156:@22203.4]
  wire [10:0] _T_72908; // @[Modules.scala 63:156:@22204.4]
  wire [10:0] buffer_5_773; // @[Modules.scala 63:156:@22205.4]
  wire [11:0] _T_72910; // @[Modules.scala 63:156:@22207.4]
  wire [10:0] _T_72911; // @[Modules.scala 63:156:@22208.4]
  wire [10:0] buffer_5_774; // @[Modules.scala 63:156:@22209.4]
  wire [11:0] _T_72913; // @[Modules.scala 63:156:@22211.4]
  wire [10:0] _T_72914; // @[Modules.scala 63:156:@22212.4]
  wire [10:0] buffer_5_775; // @[Modules.scala 63:156:@22213.4]
  wire [11:0] _T_72916; // @[Modules.scala 63:156:@22215.4]
  wire [10:0] _T_72917; // @[Modules.scala 63:156:@22216.4]
  wire [10:0] buffer_5_776; // @[Modules.scala 63:156:@22217.4]
  wire [11:0] _T_72919; // @[Modules.scala 63:156:@22219.4]
  wire [10:0] _T_72920; // @[Modules.scala 63:156:@22220.4]
  wire [10:0] buffer_5_777; // @[Modules.scala 63:156:@22221.4]
  wire [11:0] _T_72922; // @[Modules.scala 63:156:@22223.4]
  wire [10:0] _T_72923; // @[Modules.scala 63:156:@22224.4]
  wire [10:0] buffer_5_778; // @[Modules.scala 63:156:@22225.4]
  wire [11:0] _T_72925; // @[Modules.scala 63:156:@22227.4]
  wire [10:0] _T_72926; // @[Modules.scala 63:156:@22228.4]
  wire [10:0] buffer_5_779; // @[Modules.scala 63:156:@22229.4]
  wire [11:0] _T_72928; // @[Modules.scala 63:156:@22231.4]
  wire [10:0] _T_72929; // @[Modules.scala 63:156:@22232.4]
  wire [10:0] buffer_5_780; // @[Modules.scala 63:156:@22233.4]
  wire [11:0] _T_72931; // @[Modules.scala 63:156:@22235.4]
  wire [10:0] _T_72932; // @[Modules.scala 63:156:@22236.4]
  wire [10:0] buffer_5_781; // @[Modules.scala 63:156:@22237.4]
  wire [11:0] _T_72934; // @[Modules.scala 63:156:@22239.4]
  wire [10:0] _T_72935; // @[Modules.scala 63:156:@22240.4]
  wire [10:0] buffer_5_782; // @[Modules.scala 63:156:@22241.4]
  wire [11:0] _T_72937; // @[Modules.scala 63:156:@22243.4]
  wire [10:0] _T_72938; // @[Modules.scala 63:156:@22244.4]
  wire [10:0] buffer_5_783; // @[Modules.scala 63:156:@22245.4]
  wire [5:0] _T_73239; // @[Modules.scala 46:37:@22559.4]
  wire [4:0] _T_73240; // @[Modules.scala 46:37:@22560.4]
  wire [4:0] _T_73241; // @[Modules.scala 46:37:@22561.4]
  wire [5:0] _T_73242; // @[Modules.scala 46:47:@22562.4]
  wire [4:0] _T_73243; // @[Modules.scala 46:47:@22563.4]
  wire [4:0] _T_73244; // @[Modules.scala 46:47:@22564.4]
  wire [5:0] _T_73259; // @[Modules.scala 40:46:@22580.4]
  wire [4:0] _T_73260; // @[Modules.scala 40:46:@22581.4]
  wire [4:0] _T_73261; // @[Modules.scala 40:46:@22582.4]
  wire [5:0] _T_73328; // @[Modules.scala 46:47:@22651.4]
  wire [4:0] _T_73329; // @[Modules.scala 46:47:@22652.4]
  wire [4:0] _T_73330; // @[Modules.scala 46:47:@22653.4]
  wire [5:0] _T_73375; // @[Modules.scala 40:46:@22702.4]
  wire [4:0] _T_73376; // @[Modules.scala 40:46:@22703.4]
  wire [4:0] _T_73377; // @[Modules.scala 40:46:@22704.4]
  wire [5:0] _T_73382; // @[Modules.scala 43:47:@22709.4]
  wire [4:0] _T_73383; // @[Modules.scala 43:47:@22710.4]
  wire [4:0] _T_73384; // @[Modules.scala 43:47:@22711.4]
  wire [5:0] _T_73437; // @[Modules.scala 46:47:@22766.4]
  wire [4:0] _T_73438; // @[Modules.scala 46:47:@22767.4]
  wire [4:0] _T_73439; // @[Modules.scala 46:47:@22768.4]
  wire [5:0] _T_73454; // @[Modules.scala 43:47:@22784.4]
  wire [4:0] _T_73455; // @[Modules.scala 43:47:@22785.4]
  wire [4:0] _T_73456; // @[Modules.scala 43:47:@22786.4]
  wire [5:0] _T_73490; // @[Modules.scala 43:47:@22825.4]
  wire [4:0] _T_73491; // @[Modules.scala 43:47:@22826.4]
  wire [4:0] _T_73492; // @[Modules.scala 43:47:@22827.4]
  wire [5:0] _T_73507; // @[Modules.scala 40:46:@22843.4]
  wire [4:0] _T_73508; // @[Modules.scala 40:46:@22844.4]
  wire [4:0] _T_73509; // @[Modules.scala 40:46:@22845.4]
  wire [5:0] _T_73514; // @[Modules.scala 46:47:@22850.4]
  wire [4:0] _T_73515; // @[Modules.scala 46:47:@22851.4]
  wire [4:0] _T_73516; // @[Modules.scala 46:47:@22852.4]
  wire [5:0] _T_73530; // @[Modules.scala 37:46:@22869.4]
  wire [4:0] _T_73531; // @[Modules.scala 37:46:@22870.4]
  wire [4:0] _T_73532; // @[Modules.scala 37:46:@22871.4]
  wire [5:0] _T_73549; // @[Modules.scala 40:46:@22892.4]
  wire [4:0] _T_73550; // @[Modules.scala 40:46:@22893.4]
  wire [4:0] _T_73551; // @[Modules.scala 40:46:@22894.4]
  wire [5:0] _T_73608; // @[Modules.scala 43:47:@22959.4]
  wire [4:0] _T_73609; // @[Modules.scala 43:47:@22960.4]
  wire [4:0] _T_73610; // @[Modules.scala 43:47:@22961.4]
  wire [5:0] _T_73611; // @[Modules.scala 40:46:@22963.4]
  wire [4:0] _T_73612; // @[Modules.scala 40:46:@22964.4]
  wire [4:0] _T_73613; // @[Modules.scala 40:46:@22965.4]
  wire [5:0] _T_73617; // @[Modules.scala 40:46:@22971.4]
  wire [4:0] _T_73618; // @[Modules.scala 40:46:@22972.4]
  wire [4:0] _T_73619; // @[Modules.scala 40:46:@22973.4]
  wire [5:0] _T_73651; // @[Modules.scala 40:46:@23007.4]
  wire [4:0] _T_73652; // @[Modules.scala 40:46:@23008.4]
  wire [4:0] _T_73653; // @[Modules.scala 40:46:@23009.4]
  wire [5:0] _T_73657; // @[Modules.scala 37:46:@23015.4]
  wire [4:0] _T_73658; // @[Modules.scala 37:46:@23016.4]
  wire [4:0] _T_73659; // @[Modules.scala 37:46:@23017.4]
  wire [5:0] _T_73727; // @[Modules.scala 40:46:@23092.4]
  wire [4:0] _T_73728; // @[Modules.scala 40:46:@23093.4]
  wire [4:0] _T_73729; // @[Modules.scala 40:46:@23094.4]
  wire [5:0] _T_73750; // @[Modules.scala 43:47:@23118.4]
  wire [4:0] _T_73751; // @[Modules.scala 43:47:@23119.4]
  wire [4:0] _T_73752; // @[Modules.scala 43:47:@23120.4]
  wire [5:0] _T_73792; // @[Modules.scala 43:47:@23160.4]
  wire [4:0] _T_73793; // @[Modules.scala 43:47:@23161.4]
  wire [4:0] _T_73794; // @[Modules.scala 43:47:@23162.4]
  wire [5:0] _T_73806; // @[Modules.scala 43:47:@23174.4]
  wire [4:0] _T_73807; // @[Modules.scala 43:47:@23175.4]
  wire [4:0] _T_73808; // @[Modules.scala 43:47:@23176.4]
  wire [5:0] _T_73819; // @[Modules.scala 43:47:@23189.4]
  wire [4:0] _T_73820; // @[Modules.scala 43:47:@23190.4]
  wire [4:0] _T_73821; // @[Modules.scala 43:47:@23191.4]
  wire [5:0] _T_73822; // @[Modules.scala 37:46:@23193.4]
  wire [4:0] _T_73823; // @[Modules.scala 37:46:@23194.4]
  wire [4:0] _T_73824; // @[Modules.scala 37:46:@23195.4]
  wire [5:0] _T_73849; // @[Modules.scala 46:47:@23222.4]
  wire [4:0] _T_73850; // @[Modules.scala 46:47:@23223.4]
  wire [4:0] _T_73851; // @[Modules.scala 46:47:@23224.4]
  wire [5:0] _T_73859; // @[Modules.scala 37:46:@23233.4]
  wire [4:0] _T_73860; // @[Modules.scala 37:46:@23234.4]
  wire [4:0] _T_73861; // @[Modules.scala 37:46:@23235.4]
  wire [5:0] _T_73862; // @[Modules.scala 37:46:@23237.4]
  wire [4:0] _T_73863; // @[Modules.scala 37:46:@23238.4]
  wire [4:0] _T_73864; // @[Modules.scala 37:46:@23239.4]
  wire [5:0] _T_73869; // @[Modules.scala 43:47:@23244.4]
  wire [4:0] _T_73870; // @[Modules.scala 43:47:@23245.4]
  wire [4:0] _T_73871; // @[Modules.scala 43:47:@23246.4]
  wire [5:0] _T_73879; // @[Modules.scala 43:47:@23255.4]
  wire [4:0] _T_73880; // @[Modules.scala 43:47:@23256.4]
  wire [4:0] _T_73881; // @[Modules.scala 43:47:@23257.4]
  wire [5:0] _T_73893; // @[Modules.scala 43:47:@23269.4]
  wire [4:0] _T_73894; // @[Modules.scala 43:47:@23270.4]
  wire [4:0] _T_73895; // @[Modules.scala 43:47:@23271.4]
  wire [5:0] _T_73906; // @[Modules.scala 43:47:@23284.4]
  wire [4:0] _T_73907; // @[Modules.scala 43:47:@23285.4]
  wire [4:0] _T_73908; // @[Modules.scala 43:47:@23286.4]
  wire [5:0] _T_73909; // @[Modules.scala 40:46:@23288.4]
  wire [4:0] _T_73910; // @[Modules.scala 40:46:@23289.4]
  wire [4:0] _T_73911; // @[Modules.scala 40:46:@23290.4]
  wire [5:0] _T_73959; // @[Modules.scala 43:47:@23343.4]
  wire [4:0] _T_73960; // @[Modules.scala 43:47:@23344.4]
  wire [4:0] _T_73961; // @[Modules.scala 43:47:@23345.4]
  wire [5:0] _T_73992; // @[Modules.scala 43:47:@23380.4]
  wire [4:0] _T_73993; // @[Modules.scala 43:47:@23381.4]
  wire [4:0] _T_73994; // @[Modules.scala 43:47:@23382.4]
  wire [5:0] _T_74045; // @[Modules.scala 40:46:@23439.4]
  wire [4:0] _T_74046; // @[Modules.scala 40:46:@23440.4]
  wire [4:0] _T_74047; // @[Modules.scala 40:46:@23441.4]
  wire [5:0] _T_74079; // @[Modules.scala 40:46:@23475.4]
  wire [4:0] _T_74080; // @[Modules.scala 40:46:@23476.4]
  wire [4:0] _T_74081; // @[Modules.scala 40:46:@23477.4]
  wire [5:0] _T_74082; // @[Modules.scala 40:46:@23479.4]
  wire [4:0] _T_74083; // @[Modules.scala 40:46:@23480.4]
  wire [4:0] _T_74084; // @[Modules.scala 40:46:@23481.4]
  wire [5:0] _T_74089; // @[Modules.scala 43:47:@23486.4]
  wire [4:0] _T_74090; // @[Modules.scala 43:47:@23487.4]
  wire [4:0] _T_74091; // @[Modules.scala 43:47:@23488.4]
  wire [5:0] _T_74099; // @[Modules.scala 43:47:@23497.4]
  wire [4:0] _T_74100; // @[Modules.scala 43:47:@23498.4]
  wire [4:0] _T_74101; // @[Modules.scala 43:47:@23499.4]
  wire [5:0] _T_74105; // @[Modules.scala 37:46:@23505.4]
  wire [4:0] _T_74106; // @[Modules.scala 37:46:@23506.4]
  wire [4:0] _T_74107; // @[Modules.scala 37:46:@23507.4]
  wire [5:0] _T_74111; // @[Modules.scala 40:46:@23513.4]
  wire [4:0] _T_74112; // @[Modules.scala 40:46:@23514.4]
  wire [4:0] _T_74113; // @[Modules.scala 40:46:@23515.4]
  wire [5:0] _T_74151; // @[Modules.scala 43:47:@23557.4]
  wire [4:0] _T_74152; // @[Modules.scala 43:47:@23558.4]
  wire [4:0] _T_74153; // @[Modules.scala 43:47:@23559.4]
  wire [5:0] _T_74167; // @[Modules.scala 40:46:@23576.4]
  wire [4:0] _T_74168; // @[Modules.scala 40:46:@23577.4]
  wire [4:0] _T_74169; // @[Modules.scala 40:46:@23578.4]
  wire [5:0] _T_74173; // @[Modules.scala 40:46:@23584.4]
  wire [4:0] _T_74174; // @[Modules.scala 40:46:@23585.4]
  wire [4:0] _T_74175; // @[Modules.scala 40:46:@23586.4]
  wire [5:0] _T_74211; // @[Modules.scala 43:47:@23623.4]
  wire [4:0] _T_74212; // @[Modules.scala 43:47:@23624.4]
  wire [4:0] _T_74213; // @[Modules.scala 43:47:@23625.4]
  wire [5:0] _T_74260; // @[Modules.scala 37:46:@23679.4]
  wire [4:0] _T_74261; // @[Modules.scala 37:46:@23680.4]
  wire [4:0] _T_74262; // @[Modules.scala 37:46:@23681.4]
  wire [5:0] _T_74263; // @[Modules.scala 40:46:@23683.4]
  wire [4:0] _T_74264; // @[Modules.scala 40:46:@23684.4]
  wire [4:0] _T_74265; // @[Modules.scala 40:46:@23685.4]
  wire [5:0] _T_74315; // @[Modules.scala 46:47:@23736.4]
  wire [4:0] _T_74316; // @[Modules.scala 46:47:@23737.4]
  wire [4:0] _T_74317; // @[Modules.scala 46:47:@23738.4]
  wire [5:0] _T_74417; // @[Modules.scala 46:37:@23838.4]
  wire [4:0] _T_74418; // @[Modules.scala 46:37:@23839.4]
  wire [4:0] _T_74419; // @[Modules.scala 46:37:@23840.4]
  wire [5:0] _T_74420; // @[Modules.scala 46:47:@23841.4]
  wire [4:0] _T_74421; // @[Modules.scala 46:47:@23842.4]
  wire [4:0] _T_74422; // @[Modules.scala 46:47:@23843.4]
  wire [5:0] _T_74511; // @[Modules.scala 46:47:@23932.4]
  wire [4:0] _T_74512; // @[Modules.scala 46:47:@23933.4]
  wire [4:0] _T_74513; // @[Modules.scala 46:47:@23934.4]
  wire [5:0] _T_74542; // @[Modules.scala 37:46:@23964.4]
  wire [4:0] _T_74543; // @[Modules.scala 37:46:@23965.4]
  wire [4:0] _T_74544; // @[Modules.scala 37:46:@23966.4]
  wire [5:0] _T_74598; // @[Modules.scala 46:47:@24020.4]
  wire [4:0] _T_74599; // @[Modules.scala 46:47:@24021.4]
  wire [4:0] _T_74600; // @[Modules.scala 46:47:@24022.4]
  wire [5:0] _T_74626; // @[Modules.scala 43:47:@24048.4]
  wire [4:0] _T_74627; // @[Modules.scala 43:47:@24049.4]
  wire [4:0] _T_74628; // @[Modules.scala 43:47:@24050.4]
  wire [5:0] _T_74664; // @[Modules.scala 43:47:@24087.4]
  wire [4:0] _T_74665; // @[Modules.scala 43:47:@24088.4]
  wire [4:0] _T_74666; // @[Modules.scala 43:47:@24089.4]
  wire [5:0] _T_74681; // @[Modules.scala 43:47:@24105.4]
  wire [4:0] _T_74682; // @[Modules.scala 43:47:@24106.4]
  wire [4:0] _T_74683; // @[Modules.scala 43:47:@24107.4]
  wire [5:0] _T_74709; // @[Modules.scala 46:47:@24133.4]
  wire [4:0] _T_74710; // @[Modules.scala 46:47:@24134.4]
  wire [4:0] _T_74711; // @[Modules.scala 46:47:@24135.4]
  wire [5:0] _T_74730; // @[Modules.scala 46:37:@24155.4]
  wire [4:0] _T_74731; // @[Modules.scala 46:37:@24156.4]
  wire [4:0] _T_74732; // @[Modules.scala 46:37:@24157.4]
  wire [5:0] _T_74733; // @[Modules.scala 46:47:@24158.4]
  wire [4:0] _T_74734; // @[Modules.scala 46:47:@24159.4]
  wire [4:0] _T_74735; // @[Modules.scala 46:47:@24160.4]
  wire [5:0] _T_74749; // @[Modules.scala 40:46:@24177.4]
  wire [4:0] _T_74750; // @[Modules.scala 40:46:@24178.4]
  wire [4:0] _T_74751; // @[Modules.scala 40:46:@24179.4]
  wire [5:0] _T_74815; // @[Modules.scala 46:47:@24244.4]
  wire [4:0] _T_74816; // @[Modules.scala 46:47:@24245.4]
  wire [4:0] _T_74817; // @[Modules.scala 46:47:@24246.4]
  wire [5:0] _T_74927; // @[Modules.scala 40:46:@24363.4]
  wire [4:0] _T_74928; // @[Modules.scala 40:46:@24364.4]
  wire [4:0] _T_74929; // @[Modules.scala 40:46:@24365.4]
  wire [5:0] _T_74941; // @[Modules.scala 43:47:@24377.4]
  wire [4:0] _T_74942; // @[Modules.scala 43:47:@24378.4]
  wire [4:0] _T_74943; // @[Modules.scala 43:47:@24379.4]
  wire [5:0] _T_75056; // @[Modules.scala 43:47:@24507.4]
  wire [4:0] _T_75057; // @[Modules.scala 43:47:@24508.4]
  wire [4:0] _T_75058; // @[Modules.scala 43:47:@24509.4]
  wire [5:0] _T_75080; // @[Modules.scala 43:47:@24532.4]
  wire [4:0] _T_75081; // @[Modules.scala 43:47:@24533.4]
  wire [4:0] _T_75082; // @[Modules.scala 43:47:@24534.4]
  wire [11:0] _T_75103; // @[Modules.scala 50:57:@24558.4]
  wire [10:0] _T_75104; // @[Modules.scala 50:57:@24559.4]
  wire [10:0] buffer_6_393; // @[Modules.scala 50:57:@24560.4]
  wire [11:0] _T_75106; // @[Modules.scala 50:57:@24562.4]
  wire [10:0] _T_75107; // @[Modules.scala 50:57:@24563.4]
  wire [10:0] buffer_6_394; // @[Modules.scala 50:57:@24564.4]
  wire [11:0] _T_75139; // @[Modules.scala 50:57:@24606.4]
  wire [10:0] _T_75140; // @[Modules.scala 50:57:@24607.4]
  wire [10:0] buffer_6_405; // @[Modules.scala 50:57:@24608.4]
  wire [11:0] _T_75142; // @[Modules.scala 50:57:@24610.4]
  wire [10:0] _T_75143; // @[Modules.scala 50:57:@24611.4]
  wire [10:0] buffer_6_406; // @[Modules.scala 50:57:@24612.4]
  wire [11:0] _T_75163; // @[Modules.scala 50:57:@24638.4]
  wire [10:0] _T_75164; // @[Modules.scala 50:57:@24639.4]
  wire [10:0] buffer_6_413; // @[Modules.scala 50:57:@24640.4]
  wire [11:0] _T_75169; // @[Modules.scala 50:57:@24646.4]
  wire [10:0] _T_75170; // @[Modules.scala 50:57:@24647.4]
  wire [10:0] buffer_6_415; // @[Modules.scala 50:57:@24648.4]
  wire [10:0] buffer_6_50; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75175; // @[Modules.scala 50:57:@24654.4]
  wire [10:0] _T_75176; // @[Modules.scala 50:57:@24655.4]
  wire [10:0] buffer_6_417; // @[Modules.scala 50:57:@24656.4]
  wire [10:0] buffer_6_53; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75178; // @[Modules.scala 50:57:@24658.4]
  wire [10:0] _T_75179; // @[Modules.scala 50:57:@24659.4]
  wire [10:0] buffer_6_418; // @[Modules.scala 50:57:@24660.4]
  wire [11:0] _T_75181; // @[Modules.scala 50:57:@24662.4]
  wire [10:0] _T_75182; // @[Modules.scala 50:57:@24663.4]
  wire [10:0] buffer_6_419; // @[Modules.scala 50:57:@24664.4]
  wire [10:0] buffer_6_64; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75196; // @[Modules.scala 50:57:@24682.4]
  wire [10:0] _T_75197; // @[Modules.scala 50:57:@24683.4]
  wire [10:0] buffer_6_424; // @[Modules.scala 50:57:@24684.4]
  wire [10:0] buffer_6_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75208; // @[Modules.scala 50:57:@24698.4]
  wire [10:0] _T_75209; // @[Modules.scala 50:57:@24699.4]
  wire [10:0] buffer_6_428; // @[Modules.scala 50:57:@24700.4]
  wire [10:0] buffer_6_74; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75211; // @[Modules.scala 50:57:@24702.4]
  wire [10:0] _T_75212; // @[Modules.scala 50:57:@24703.4]
  wire [10:0] buffer_6_429; // @[Modules.scala 50:57:@24704.4]
  wire [10:0] buffer_6_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75223; // @[Modules.scala 50:57:@24718.4]
  wire [10:0] _T_75224; // @[Modules.scala 50:57:@24719.4]
  wire [10:0] buffer_6_433; // @[Modules.scala 50:57:@24720.4]
  wire [10:0] buffer_6_86; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75229; // @[Modules.scala 50:57:@24726.4]
  wire [10:0] _T_75230; // @[Modules.scala 50:57:@24727.4]
  wire [10:0] buffer_6_435; // @[Modules.scala 50:57:@24728.4]
  wire [11:0] _T_75232; // @[Modules.scala 50:57:@24730.4]
  wire [10:0] _T_75233; // @[Modules.scala 50:57:@24731.4]
  wire [10:0] buffer_6_436; // @[Modules.scala 50:57:@24732.4]
  wire [10:0] buffer_6_94; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75241; // @[Modules.scala 50:57:@24742.4]
  wire [10:0] _T_75242; // @[Modules.scala 50:57:@24743.4]
  wire [10:0] buffer_6_439; // @[Modules.scala 50:57:@24744.4]
  wire [10:0] buffer_6_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75244; // @[Modules.scala 50:57:@24746.4]
  wire [10:0] _T_75245; // @[Modules.scala 50:57:@24747.4]
  wire [10:0] buffer_6_440; // @[Modules.scala 50:57:@24748.4]
  wire [10:0] buffer_6_98; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75247; // @[Modules.scala 50:57:@24750.4]
  wire [10:0] _T_75248; // @[Modules.scala 50:57:@24751.4]
  wire [10:0] buffer_6_441; // @[Modules.scala 50:57:@24752.4]
  wire [11:0] _T_75250; // @[Modules.scala 50:57:@24754.4]
  wire [10:0] _T_75251; // @[Modules.scala 50:57:@24755.4]
  wire [10:0] buffer_6_442; // @[Modules.scala 50:57:@24756.4]
  wire [10:0] buffer_6_102; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75253; // @[Modules.scala 50:57:@24758.4]
  wire [10:0] _T_75254; // @[Modules.scala 50:57:@24759.4]
  wire [10:0] buffer_6_443; // @[Modules.scala 50:57:@24760.4]
  wire [11:0] _T_75256; // @[Modules.scala 50:57:@24762.4]
  wire [10:0] _T_75257; // @[Modules.scala 50:57:@24763.4]
  wire [10:0] buffer_6_444; // @[Modules.scala 50:57:@24764.4]
  wire [10:0] buffer_6_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75259; // @[Modules.scala 50:57:@24766.4]
  wire [10:0] _T_75260; // @[Modules.scala 50:57:@24767.4]
  wire [10:0] buffer_6_445; // @[Modules.scala 50:57:@24768.4]
  wire [11:0] _T_75262; // @[Modules.scala 50:57:@24770.4]
  wire [10:0] _T_75263; // @[Modules.scala 50:57:@24771.4]
  wire [10:0] buffer_6_446; // @[Modules.scala 50:57:@24772.4]
  wire [11:0] _T_75268; // @[Modules.scala 50:57:@24778.4]
  wire [10:0] _T_75269; // @[Modules.scala 50:57:@24779.4]
  wire [10:0] buffer_6_448; // @[Modules.scala 50:57:@24780.4]
  wire [11:0] _T_75274; // @[Modules.scala 50:57:@24786.4]
  wire [10:0] _T_75275; // @[Modules.scala 50:57:@24787.4]
  wire [10:0] buffer_6_450; // @[Modules.scala 50:57:@24788.4]
  wire [10:0] buffer_6_120; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75280; // @[Modules.scala 50:57:@24794.4]
  wire [10:0] _T_75281; // @[Modules.scala 50:57:@24795.4]
  wire [10:0] buffer_6_452; // @[Modules.scala 50:57:@24796.4]
  wire [10:0] buffer_6_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75283; // @[Modules.scala 50:57:@24798.4]
  wire [10:0] _T_75284; // @[Modules.scala 50:57:@24799.4]
  wire [10:0] buffer_6_453; // @[Modules.scala 50:57:@24800.4]
  wire [11:0] _T_75289; // @[Modules.scala 50:57:@24806.4]
  wire [10:0] _T_75290; // @[Modules.scala 50:57:@24807.4]
  wire [10:0] buffer_6_455; // @[Modules.scala 50:57:@24808.4]
  wire [10:0] buffer_6_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75292; // @[Modules.scala 50:57:@24810.4]
  wire [10:0] _T_75293; // @[Modules.scala 50:57:@24811.4]
  wire [10:0] buffer_6_456; // @[Modules.scala 50:57:@24812.4]
  wire [10:0] buffer_6_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75295; // @[Modules.scala 50:57:@24814.4]
  wire [10:0] _T_75296; // @[Modules.scala 50:57:@24815.4]
  wire [10:0] buffer_6_457; // @[Modules.scala 50:57:@24816.4]
  wire [11:0] _T_75304; // @[Modules.scala 50:57:@24826.4]
  wire [10:0] _T_75305; // @[Modules.scala 50:57:@24827.4]
  wire [10:0] buffer_6_460; // @[Modules.scala 50:57:@24828.4]
  wire [11:0] _T_75310; // @[Modules.scala 50:57:@24834.4]
  wire [10:0] _T_75311; // @[Modules.scala 50:57:@24835.4]
  wire [10:0] buffer_6_462; // @[Modules.scala 50:57:@24836.4]
  wire [10:0] buffer_6_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75316; // @[Modules.scala 50:57:@24842.4]
  wire [10:0] _T_75317; // @[Modules.scala 50:57:@24843.4]
  wire [10:0] buffer_6_464; // @[Modules.scala 50:57:@24844.4]
  wire [11:0] _T_75319; // @[Modules.scala 50:57:@24846.4]
  wire [10:0] _T_75320; // @[Modules.scala 50:57:@24847.4]
  wire [10:0] buffer_6_465; // @[Modules.scala 50:57:@24848.4]
  wire [11:0] _T_75322; // @[Modules.scala 50:57:@24850.4]
  wire [10:0] _T_75323; // @[Modules.scala 50:57:@24851.4]
  wire [10:0] buffer_6_466; // @[Modules.scala 50:57:@24852.4]
  wire [10:0] buffer_6_150; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75325; // @[Modules.scala 50:57:@24854.4]
  wire [10:0] _T_75326; // @[Modules.scala 50:57:@24855.4]
  wire [10:0] buffer_6_467; // @[Modules.scala 50:57:@24856.4]
  wire [11:0] _T_75331; // @[Modules.scala 50:57:@24862.4]
  wire [10:0] _T_75332; // @[Modules.scala 50:57:@24863.4]
  wire [10:0] buffer_6_469; // @[Modules.scala 50:57:@24864.4]
  wire [10:0] buffer_6_156; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75334; // @[Modules.scala 50:57:@24866.4]
  wire [10:0] _T_75335; // @[Modules.scala 50:57:@24867.4]
  wire [10:0] buffer_6_470; // @[Modules.scala 50:57:@24868.4]
  wire [10:0] buffer_6_158; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75337; // @[Modules.scala 50:57:@24870.4]
  wire [10:0] _T_75338; // @[Modules.scala 50:57:@24871.4]
  wire [10:0] buffer_6_471; // @[Modules.scala 50:57:@24872.4]
  wire [10:0] buffer_6_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75340; // @[Modules.scala 50:57:@24874.4]
  wire [10:0] _T_75341; // @[Modules.scala 50:57:@24875.4]
  wire [10:0] buffer_6_472; // @[Modules.scala 50:57:@24876.4]
  wire [10:0] buffer_6_162; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75343; // @[Modules.scala 50:57:@24878.4]
  wire [10:0] _T_75344; // @[Modules.scala 50:57:@24879.4]
  wire [10:0] buffer_6_473; // @[Modules.scala 50:57:@24880.4]
  wire [10:0] buffer_6_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75349; // @[Modules.scala 50:57:@24886.4]
  wire [10:0] _T_75350; // @[Modules.scala 50:57:@24887.4]
  wire [10:0] buffer_6_475; // @[Modules.scala 50:57:@24888.4]
  wire [10:0] buffer_6_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75352; // @[Modules.scala 50:57:@24890.4]
  wire [10:0] _T_75353; // @[Modules.scala 50:57:@24891.4]
  wire [10:0] buffer_6_476; // @[Modules.scala 50:57:@24892.4]
  wire [10:0] buffer_6_170; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75355; // @[Modules.scala 50:57:@24894.4]
  wire [10:0] _T_75356; // @[Modules.scala 50:57:@24895.4]
  wire [10:0] buffer_6_477; // @[Modules.scala 50:57:@24896.4]
  wire [10:0] buffer_6_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75358; // @[Modules.scala 50:57:@24898.4]
  wire [10:0] _T_75359; // @[Modules.scala 50:57:@24899.4]
  wire [10:0] buffer_6_478; // @[Modules.scala 50:57:@24900.4]
  wire [10:0] buffer_6_175; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75361; // @[Modules.scala 50:57:@24902.4]
  wire [10:0] _T_75362; // @[Modules.scala 50:57:@24903.4]
  wire [10:0] buffer_6_479; // @[Modules.scala 50:57:@24904.4]
  wire [10:0] buffer_6_178; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75367; // @[Modules.scala 50:57:@24910.4]
  wire [10:0] _T_75368; // @[Modules.scala 50:57:@24911.4]
  wire [10:0] buffer_6_481; // @[Modules.scala 50:57:@24912.4]
  wire [11:0] _T_75373; // @[Modules.scala 50:57:@24918.4]
  wire [10:0] _T_75374; // @[Modules.scala 50:57:@24919.4]
  wire [10:0] buffer_6_483; // @[Modules.scala 50:57:@24920.4]
  wire [11:0] _T_75379; // @[Modules.scala 50:57:@24926.4]
  wire [10:0] _T_75380; // @[Modules.scala 50:57:@24927.4]
  wire [10:0] buffer_6_485; // @[Modules.scala 50:57:@24928.4]
  wire [10:0] buffer_6_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75382; // @[Modules.scala 50:57:@24930.4]
  wire [10:0] _T_75383; // @[Modules.scala 50:57:@24931.4]
  wire [10:0] buffer_6_486; // @[Modules.scala 50:57:@24932.4]
  wire [10:0] buffer_6_196; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75394; // @[Modules.scala 50:57:@24946.4]
  wire [10:0] _T_75395; // @[Modules.scala 50:57:@24947.4]
  wire [10:0] buffer_6_490; // @[Modules.scala 50:57:@24948.4]
  wire [11:0] _T_75400; // @[Modules.scala 50:57:@24954.4]
  wire [10:0] _T_75401; // @[Modules.scala 50:57:@24955.4]
  wire [10:0] buffer_6_492; // @[Modules.scala 50:57:@24956.4]
  wire [11:0] _T_75403; // @[Modules.scala 50:57:@24958.4]
  wire [10:0] _T_75404; // @[Modules.scala 50:57:@24959.4]
  wire [10:0] buffer_6_493; // @[Modules.scala 50:57:@24960.4]
  wire [10:0] buffer_6_207; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75409; // @[Modules.scala 50:57:@24966.4]
  wire [10:0] _T_75410; // @[Modules.scala 50:57:@24967.4]
  wire [10:0] buffer_6_495; // @[Modules.scala 50:57:@24968.4]
  wire [11:0] _T_75412; // @[Modules.scala 50:57:@24970.4]
  wire [10:0] _T_75413; // @[Modules.scala 50:57:@24971.4]
  wire [10:0] buffer_6_496; // @[Modules.scala 50:57:@24972.4]
  wire [11:0] _T_75415; // @[Modules.scala 50:57:@24974.4]
  wire [10:0] _T_75416; // @[Modules.scala 50:57:@24975.4]
  wire [10:0] buffer_6_497; // @[Modules.scala 50:57:@24976.4]
  wire [10:0] buffer_6_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75418; // @[Modules.scala 50:57:@24978.4]
  wire [10:0] _T_75419; // @[Modules.scala 50:57:@24979.4]
  wire [10:0] buffer_6_498; // @[Modules.scala 50:57:@24980.4]
  wire [10:0] buffer_6_214; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75421; // @[Modules.scala 50:57:@24982.4]
  wire [10:0] _T_75422; // @[Modules.scala 50:57:@24983.4]
  wire [10:0] buffer_6_499; // @[Modules.scala 50:57:@24984.4]
  wire [10:0] buffer_6_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75424; // @[Modules.scala 50:57:@24986.4]
  wire [10:0] _T_75425; // @[Modules.scala 50:57:@24987.4]
  wire [10:0] buffer_6_500; // @[Modules.scala 50:57:@24988.4]
  wire [10:0] buffer_6_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75427; // @[Modules.scala 50:57:@24990.4]
  wire [10:0] _T_75428; // @[Modules.scala 50:57:@24991.4]
  wire [10:0] buffer_6_501; // @[Modules.scala 50:57:@24992.4]
  wire [10:0] buffer_6_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75430; // @[Modules.scala 50:57:@24994.4]
  wire [10:0] _T_75431; // @[Modules.scala 50:57:@24995.4]
  wire [10:0] buffer_6_502; // @[Modules.scala 50:57:@24996.4]
  wire [11:0] _T_75436; // @[Modules.scala 50:57:@25002.4]
  wire [10:0] _T_75437; // @[Modules.scala 50:57:@25003.4]
  wire [10:0] buffer_6_504; // @[Modules.scala 50:57:@25004.4]
  wire [10:0] buffer_6_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75442; // @[Modules.scala 50:57:@25010.4]
  wire [10:0] _T_75443; // @[Modules.scala 50:57:@25011.4]
  wire [10:0] buffer_6_506; // @[Modules.scala 50:57:@25012.4]
  wire [11:0] _T_75445; // @[Modules.scala 50:57:@25014.4]
  wire [10:0] _T_75446; // @[Modules.scala 50:57:@25015.4]
  wire [10:0] buffer_6_507; // @[Modules.scala 50:57:@25016.4]
  wire [10:0] buffer_6_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75448; // @[Modules.scala 50:57:@25018.4]
  wire [10:0] _T_75449; // @[Modules.scala 50:57:@25019.4]
  wire [10:0] buffer_6_508; // @[Modules.scala 50:57:@25020.4]
  wire [10:0] buffer_6_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75451; // @[Modules.scala 50:57:@25022.4]
  wire [10:0] _T_75452; // @[Modules.scala 50:57:@25023.4]
  wire [10:0] buffer_6_509; // @[Modules.scala 50:57:@25024.4]
  wire [11:0] _T_75457; // @[Modules.scala 50:57:@25030.4]
  wire [10:0] _T_75458; // @[Modules.scala 50:57:@25031.4]
  wire [10:0] buffer_6_511; // @[Modules.scala 50:57:@25032.4]
  wire [10:0] buffer_6_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75460; // @[Modules.scala 50:57:@25034.4]
  wire [10:0] _T_75461; // @[Modules.scala 50:57:@25035.4]
  wire [10:0] buffer_6_512; // @[Modules.scala 50:57:@25036.4]
  wire [11:0] _T_75463; // @[Modules.scala 50:57:@25038.4]
  wire [10:0] _T_75464; // @[Modules.scala 50:57:@25039.4]
  wire [10:0] buffer_6_513; // @[Modules.scala 50:57:@25040.4]
  wire [11:0] _T_75469; // @[Modules.scala 50:57:@25046.4]
  wire [10:0] _T_75470; // @[Modules.scala 50:57:@25047.4]
  wire [10:0] buffer_6_515; // @[Modules.scala 50:57:@25048.4]
  wire [10:0] buffer_6_252; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75478; // @[Modules.scala 50:57:@25058.4]
  wire [10:0] _T_75479; // @[Modules.scala 50:57:@25059.4]
  wire [10:0] buffer_6_518; // @[Modules.scala 50:57:@25060.4]
  wire [11:0] _T_75487; // @[Modules.scala 50:57:@25070.4]
  wire [10:0] _T_75488; // @[Modules.scala 50:57:@25071.4]
  wire [10:0] buffer_6_521; // @[Modules.scala 50:57:@25072.4]
  wire [10:0] buffer_6_261; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75490; // @[Modules.scala 50:57:@25074.4]
  wire [10:0] _T_75491; // @[Modules.scala 50:57:@25075.4]
  wire [10:0] buffer_6_522; // @[Modules.scala 50:57:@25076.4]
  wire [11:0] _T_75505; // @[Modules.scala 50:57:@25094.4]
  wire [10:0] _T_75506; // @[Modules.scala 50:57:@25095.4]
  wire [10:0] buffer_6_527; // @[Modules.scala 50:57:@25096.4]
  wire [10:0] buffer_6_276; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75514; // @[Modules.scala 50:57:@25106.4]
  wire [10:0] _T_75515; // @[Modules.scala 50:57:@25107.4]
  wire [10:0] buffer_6_530; // @[Modules.scala 50:57:@25108.4]
  wire [10:0] buffer_6_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75532; // @[Modules.scala 50:57:@25130.4]
  wire [10:0] _T_75533; // @[Modules.scala 50:57:@25131.4]
  wire [10:0] buffer_6_536; // @[Modules.scala 50:57:@25132.4]
  wire [11:0] _T_75538; // @[Modules.scala 50:57:@25138.4]
  wire [10:0] _T_75539; // @[Modules.scala 50:57:@25139.4]
  wire [10:0] buffer_6_538; // @[Modules.scala 50:57:@25140.4]
  wire [10:0] buffer_6_294; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75541; // @[Modules.scala 50:57:@25142.4]
  wire [10:0] _T_75542; // @[Modules.scala 50:57:@25143.4]
  wire [10:0] buffer_6_539; // @[Modules.scala 50:57:@25144.4]
  wire [10:0] buffer_6_302; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75553; // @[Modules.scala 50:57:@25158.4]
  wire [10:0] _T_75554; // @[Modules.scala 50:57:@25159.4]
  wire [10:0] buffer_6_543; // @[Modules.scala 50:57:@25160.4]
  wire [10:0] buffer_6_306; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75559; // @[Modules.scala 50:57:@25166.4]
  wire [10:0] _T_75560; // @[Modules.scala 50:57:@25167.4]
  wire [10:0] buffer_6_545; // @[Modules.scala 50:57:@25168.4]
  wire [10:0] buffer_6_312; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75568; // @[Modules.scala 50:57:@25178.4]
  wire [10:0] _T_75569; // @[Modules.scala 50:57:@25179.4]
  wire [10:0] buffer_6_548; // @[Modules.scala 50:57:@25180.4]
  wire [10:0] buffer_6_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75571; // @[Modules.scala 50:57:@25182.4]
  wire [10:0] _T_75572; // @[Modules.scala 50:57:@25183.4]
  wire [10:0] buffer_6_549; // @[Modules.scala 50:57:@25184.4]
  wire [10:0] buffer_6_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75577; // @[Modules.scala 50:57:@25190.4]
  wire [10:0] _T_75578; // @[Modules.scala 50:57:@25191.4]
  wire [10:0] buffer_6_551; // @[Modules.scala 50:57:@25192.4]
  wire [10:0] buffer_6_323; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75583; // @[Modules.scala 50:57:@25198.4]
  wire [10:0] _T_75584; // @[Modules.scala 50:57:@25199.4]
  wire [10:0] buffer_6_553; // @[Modules.scala 50:57:@25200.4]
  wire [11:0] _T_75586; // @[Modules.scala 50:57:@25202.4]
  wire [10:0] _T_75587; // @[Modules.scala 50:57:@25203.4]
  wire [10:0] buffer_6_554; // @[Modules.scala 50:57:@25204.4]
  wire [10:0] buffer_6_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75589; // @[Modules.scala 50:57:@25206.4]
  wire [10:0] _T_75590; // @[Modules.scala 50:57:@25207.4]
  wire [10:0] buffer_6_555; // @[Modules.scala 50:57:@25208.4]
  wire [11:0] _T_75601; // @[Modules.scala 50:57:@25222.4]
  wire [10:0] _T_75602; // @[Modules.scala 50:57:@25223.4]
  wire [10:0] buffer_6_559; // @[Modules.scala 50:57:@25224.4]
  wire [10:0] buffer_6_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75604; // @[Modules.scala 50:57:@25226.4]
  wire [10:0] _T_75605; // @[Modules.scala 50:57:@25227.4]
  wire [10:0] buffer_6_560; // @[Modules.scala 50:57:@25228.4]
  wire [11:0] _T_75616; // @[Modules.scala 50:57:@25242.4]
  wire [10:0] _T_75617; // @[Modules.scala 50:57:@25243.4]
  wire [10:0] buffer_6_564; // @[Modules.scala 50:57:@25244.4]
  wire [11:0] _T_75619; // @[Modules.scala 50:57:@25246.4]
  wire [10:0] _T_75620; // @[Modules.scala 50:57:@25247.4]
  wire [10:0] buffer_6_565; // @[Modules.scala 50:57:@25248.4]
  wire [11:0] _T_75631; // @[Modules.scala 50:57:@25262.4]
  wire [10:0] _T_75632; // @[Modules.scala 50:57:@25263.4]
  wire [10:0] buffer_6_569; // @[Modules.scala 50:57:@25264.4]
  wire [10:0] buffer_6_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75634; // @[Modules.scala 50:57:@25266.4]
  wire [10:0] _T_75635; // @[Modules.scala 50:57:@25267.4]
  wire [10:0] buffer_6_570; // @[Modules.scala 50:57:@25268.4]
  wire [10:0] buffer_6_359; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75637; // @[Modules.scala 50:57:@25270.4]
  wire [10:0] _T_75638; // @[Modules.scala 50:57:@25271.4]
  wire [10:0] buffer_6_571; // @[Modules.scala 50:57:@25272.4]
  wire [11:0] _T_75643; // @[Modules.scala 50:57:@25278.4]
  wire [10:0] _T_75644; // @[Modules.scala 50:57:@25279.4]
  wire [10:0] buffer_6_573; // @[Modules.scala 50:57:@25280.4]
  wire [11:0] _T_75646; // @[Modules.scala 50:57:@25282.4]
  wire [10:0] _T_75647; // @[Modules.scala 50:57:@25283.4]
  wire [10:0] buffer_6_574; // @[Modules.scala 50:57:@25284.4]
  wire [11:0] _T_75661; // @[Modules.scala 50:57:@25302.4]
  wire [10:0] _T_75662; // @[Modules.scala 50:57:@25303.4]
  wire [10:0] buffer_6_579; // @[Modules.scala 50:57:@25304.4]
  wire [10:0] buffer_6_384; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75676; // @[Modules.scala 50:57:@25322.4]
  wire [10:0] _T_75677; // @[Modules.scala 50:57:@25323.4]
  wire [10:0] buffer_6_584; // @[Modules.scala 50:57:@25324.4]
  wire [10:0] buffer_6_388; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75682; // @[Modules.scala 50:57:@25330.4]
  wire [10:0] _T_75683; // @[Modules.scala 50:57:@25331.4]
  wire [10:0] buffer_6_586; // @[Modules.scala 50:57:@25332.4]
  wire [11:0] _T_75688; // @[Modules.scala 53:83:@25338.4]
  wire [10:0] _T_75689; // @[Modules.scala 53:83:@25339.4]
  wire [10:0] buffer_6_588; // @[Modules.scala 53:83:@25340.4]
  wire [11:0] _T_75691; // @[Modules.scala 53:83:@25342.4]
  wire [10:0] _T_75692; // @[Modules.scala 53:83:@25343.4]
  wire [10:0] buffer_6_589; // @[Modules.scala 53:83:@25344.4]
  wire [11:0] _T_75694; // @[Modules.scala 53:83:@25346.4]
  wire [10:0] _T_75695; // @[Modules.scala 53:83:@25347.4]
  wire [10:0] buffer_6_590; // @[Modules.scala 53:83:@25348.4]
  wire [11:0] _T_75697; // @[Modules.scala 53:83:@25350.4]
  wire [10:0] _T_75698; // @[Modules.scala 53:83:@25351.4]
  wire [10:0] buffer_6_591; // @[Modules.scala 53:83:@25352.4]
  wire [11:0] _T_75700; // @[Modules.scala 53:83:@25354.4]
  wire [10:0] _T_75701; // @[Modules.scala 53:83:@25355.4]
  wire [10:0] buffer_6_592; // @[Modules.scala 53:83:@25356.4]
  wire [11:0] _T_75706; // @[Modules.scala 53:83:@25362.4]
  wire [10:0] _T_75707; // @[Modules.scala 53:83:@25363.4]
  wire [10:0] buffer_6_594; // @[Modules.scala 53:83:@25364.4]
  wire [11:0] _T_75709; // @[Modules.scala 53:83:@25366.4]
  wire [10:0] _T_75710; // @[Modules.scala 53:83:@25367.4]
  wire [10:0] buffer_6_595; // @[Modules.scala 53:83:@25368.4]
  wire [11:0] _T_75718; // @[Modules.scala 53:83:@25378.4]
  wire [10:0] _T_75719; // @[Modules.scala 53:83:@25379.4]
  wire [10:0] buffer_6_598; // @[Modules.scala 53:83:@25380.4]
  wire [11:0] _T_75721; // @[Modules.scala 53:83:@25382.4]
  wire [10:0] _T_75722; // @[Modules.scala 53:83:@25383.4]
  wire [10:0] buffer_6_599; // @[Modules.scala 53:83:@25384.4]
  wire [11:0] _T_75724; // @[Modules.scala 53:83:@25386.4]
  wire [10:0] _T_75725; // @[Modules.scala 53:83:@25387.4]
  wire [10:0] buffer_6_600; // @[Modules.scala 53:83:@25388.4]
  wire [11:0] _T_75727; // @[Modules.scala 53:83:@25390.4]
  wire [10:0] _T_75728; // @[Modules.scala 53:83:@25391.4]
  wire [10:0] buffer_6_601; // @[Modules.scala 53:83:@25392.4]
  wire [11:0] _T_75730; // @[Modules.scala 53:83:@25394.4]
  wire [10:0] _T_75731; // @[Modules.scala 53:83:@25395.4]
  wire [10:0] buffer_6_602; // @[Modules.scala 53:83:@25396.4]
  wire [11:0] _T_75736; // @[Modules.scala 53:83:@25402.4]
  wire [10:0] _T_75737; // @[Modules.scala 53:83:@25403.4]
  wire [10:0] buffer_6_604; // @[Modules.scala 53:83:@25404.4]
  wire [11:0] _T_75739; // @[Modules.scala 53:83:@25406.4]
  wire [10:0] _T_75740; // @[Modules.scala 53:83:@25407.4]
  wire [10:0] buffer_6_605; // @[Modules.scala 53:83:@25408.4]
  wire [11:0] _T_75742; // @[Modules.scala 53:83:@25410.4]
  wire [10:0] _T_75743; // @[Modules.scala 53:83:@25411.4]
  wire [10:0] buffer_6_606; // @[Modules.scala 53:83:@25412.4]
  wire [11:0] _T_75748; // @[Modules.scala 53:83:@25418.4]
  wire [10:0] _T_75749; // @[Modules.scala 53:83:@25419.4]
  wire [10:0] buffer_6_608; // @[Modules.scala 53:83:@25420.4]
  wire [11:0] _T_75751; // @[Modules.scala 53:83:@25422.4]
  wire [10:0] _T_75752; // @[Modules.scala 53:83:@25423.4]
  wire [10:0] buffer_6_609; // @[Modules.scala 53:83:@25424.4]
  wire [11:0] _T_75754; // @[Modules.scala 53:83:@25426.4]
  wire [10:0] _T_75755; // @[Modules.scala 53:83:@25427.4]
  wire [10:0] buffer_6_610; // @[Modules.scala 53:83:@25428.4]
  wire [11:0] _T_75757; // @[Modules.scala 53:83:@25430.4]
  wire [10:0] _T_75758; // @[Modules.scala 53:83:@25431.4]
  wire [10:0] buffer_6_611; // @[Modules.scala 53:83:@25432.4]
  wire [11:0] _T_75760; // @[Modules.scala 53:83:@25434.4]
  wire [10:0] _T_75761; // @[Modules.scala 53:83:@25435.4]
  wire [10:0] buffer_6_612; // @[Modules.scala 53:83:@25436.4]
  wire [11:0] _T_75763; // @[Modules.scala 53:83:@25438.4]
  wire [10:0] _T_75764; // @[Modules.scala 53:83:@25439.4]
  wire [10:0] buffer_6_613; // @[Modules.scala 53:83:@25440.4]
  wire [11:0] _T_75766; // @[Modules.scala 53:83:@25442.4]
  wire [10:0] _T_75767; // @[Modules.scala 53:83:@25443.4]
  wire [10:0] buffer_6_614; // @[Modules.scala 53:83:@25444.4]
  wire [11:0] _T_75769; // @[Modules.scala 53:83:@25446.4]
  wire [10:0] _T_75770; // @[Modules.scala 53:83:@25447.4]
  wire [10:0] buffer_6_615; // @[Modules.scala 53:83:@25448.4]
  wire [11:0] _T_75772; // @[Modules.scala 53:83:@25450.4]
  wire [10:0] _T_75773; // @[Modules.scala 53:83:@25451.4]
  wire [10:0] buffer_6_616; // @[Modules.scala 53:83:@25452.4]
  wire [11:0] _T_75775; // @[Modules.scala 53:83:@25454.4]
  wire [10:0] _T_75776; // @[Modules.scala 53:83:@25455.4]
  wire [10:0] buffer_6_617; // @[Modules.scala 53:83:@25456.4]
  wire [11:0] _T_75778; // @[Modules.scala 53:83:@25458.4]
  wire [10:0] _T_75779; // @[Modules.scala 53:83:@25459.4]
  wire [10:0] buffer_6_618; // @[Modules.scala 53:83:@25460.4]
  wire [11:0] _T_75781; // @[Modules.scala 53:83:@25462.4]
  wire [10:0] _T_75782; // @[Modules.scala 53:83:@25463.4]
  wire [10:0] buffer_6_619; // @[Modules.scala 53:83:@25464.4]
  wire [11:0] _T_75784; // @[Modules.scala 53:83:@25466.4]
  wire [10:0] _T_75785; // @[Modules.scala 53:83:@25467.4]
  wire [10:0] buffer_6_620; // @[Modules.scala 53:83:@25468.4]
  wire [11:0] _T_75790; // @[Modules.scala 53:83:@25474.4]
  wire [10:0] _T_75791; // @[Modules.scala 53:83:@25475.4]
  wire [10:0] buffer_6_622; // @[Modules.scala 53:83:@25476.4]
  wire [11:0] _T_75793; // @[Modules.scala 53:83:@25478.4]
  wire [10:0] _T_75794; // @[Modules.scala 53:83:@25479.4]
  wire [10:0] buffer_6_623; // @[Modules.scala 53:83:@25480.4]
  wire [11:0] _T_75796; // @[Modules.scala 53:83:@25482.4]
  wire [10:0] _T_75797; // @[Modules.scala 53:83:@25483.4]
  wire [10:0] buffer_6_624; // @[Modules.scala 53:83:@25484.4]
  wire [11:0] _T_75799; // @[Modules.scala 53:83:@25486.4]
  wire [10:0] _T_75800; // @[Modules.scala 53:83:@25487.4]
  wire [10:0] buffer_6_625; // @[Modules.scala 53:83:@25488.4]
  wire [11:0] _T_75802; // @[Modules.scala 53:83:@25490.4]
  wire [10:0] _T_75803; // @[Modules.scala 53:83:@25491.4]
  wire [10:0] buffer_6_626; // @[Modules.scala 53:83:@25492.4]
  wire [11:0] _T_75805; // @[Modules.scala 53:83:@25494.4]
  wire [10:0] _T_75806; // @[Modules.scala 53:83:@25495.4]
  wire [10:0] buffer_6_627; // @[Modules.scala 53:83:@25496.4]
  wire [11:0] _T_75808; // @[Modules.scala 53:83:@25498.4]
  wire [10:0] _T_75809; // @[Modules.scala 53:83:@25499.4]
  wire [10:0] buffer_6_628; // @[Modules.scala 53:83:@25500.4]
  wire [11:0] _T_75811; // @[Modules.scala 53:83:@25502.4]
  wire [10:0] _T_75812; // @[Modules.scala 53:83:@25503.4]
  wire [10:0] buffer_6_629; // @[Modules.scala 53:83:@25504.4]
  wire [11:0] _T_75814; // @[Modules.scala 53:83:@25506.4]
  wire [10:0] _T_75815; // @[Modules.scala 53:83:@25507.4]
  wire [10:0] buffer_6_630; // @[Modules.scala 53:83:@25508.4]
  wire [11:0] _T_75817; // @[Modules.scala 53:83:@25510.4]
  wire [10:0] _T_75818; // @[Modules.scala 53:83:@25511.4]
  wire [10:0] buffer_6_631; // @[Modules.scala 53:83:@25512.4]
  wire [11:0] _T_75820; // @[Modules.scala 53:83:@25514.4]
  wire [10:0] _T_75821; // @[Modules.scala 53:83:@25515.4]
  wire [10:0] buffer_6_632; // @[Modules.scala 53:83:@25516.4]
  wire [11:0] _T_75823; // @[Modules.scala 53:83:@25518.4]
  wire [10:0] _T_75824; // @[Modules.scala 53:83:@25519.4]
  wire [10:0] buffer_6_633; // @[Modules.scala 53:83:@25520.4]
  wire [11:0] _T_75826; // @[Modules.scala 53:83:@25522.4]
  wire [10:0] _T_75827; // @[Modules.scala 53:83:@25523.4]
  wire [10:0] buffer_6_634; // @[Modules.scala 53:83:@25524.4]
  wire [11:0] _T_75829; // @[Modules.scala 53:83:@25526.4]
  wire [10:0] _T_75830; // @[Modules.scala 53:83:@25527.4]
  wire [10:0] buffer_6_635; // @[Modules.scala 53:83:@25528.4]
  wire [11:0] _T_75832; // @[Modules.scala 53:83:@25530.4]
  wire [10:0] _T_75833; // @[Modules.scala 53:83:@25531.4]
  wire [10:0] buffer_6_636; // @[Modules.scala 53:83:@25532.4]
  wire [11:0] _T_75835; // @[Modules.scala 53:83:@25534.4]
  wire [10:0] _T_75836; // @[Modules.scala 53:83:@25535.4]
  wire [10:0] buffer_6_637; // @[Modules.scala 53:83:@25536.4]
  wire [11:0] _T_75838; // @[Modules.scala 53:83:@25538.4]
  wire [10:0] _T_75839; // @[Modules.scala 53:83:@25539.4]
  wire [10:0] buffer_6_638; // @[Modules.scala 53:83:@25540.4]
  wire [11:0] _T_75841; // @[Modules.scala 53:83:@25542.4]
  wire [10:0] _T_75842; // @[Modules.scala 53:83:@25543.4]
  wire [10:0] buffer_6_639; // @[Modules.scala 53:83:@25544.4]
  wire [11:0] _T_75844; // @[Modules.scala 53:83:@25546.4]
  wire [10:0] _T_75845; // @[Modules.scala 53:83:@25547.4]
  wire [10:0] buffer_6_640; // @[Modules.scala 53:83:@25548.4]
  wire [11:0] _T_75847; // @[Modules.scala 53:83:@25550.4]
  wire [10:0] _T_75848; // @[Modules.scala 53:83:@25551.4]
  wire [10:0] buffer_6_641; // @[Modules.scala 53:83:@25552.4]
  wire [11:0] _T_75850; // @[Modules.scala 53:83:@25554.4]
  wire [10:0] _T_75851; // @[Modules.scala 53:83:@25555.4]
  wire [10:0] buffer_6_642; // @[Modules.scala 53:83:@25556.4]
  wire [11:0] _T_75853; // @[Modules.scala 53:83:@25558.4]
  wire [10:0] _T_75854; // @[Modules.scala 53:83:@25559.4]
  wire [10:0] buffer_6_643; // @[Modules.scala 53:83:@25560.4]
  wire [11:0] _T_75856; // @[Modules.scala 53:83:@25562.4]
  wire [10:0] _T_75857; // @[Modules.scala 53:83:@25563.4]
  wire [10:0] buffer_6_644; // @[Modules.scala 53:83:@25564.4]
  wire [11:0] _T_75859; // @[Modules.scala 53:83:@25566.4]
  wire [10:0] _T_75860; // @[Modules.scala 53:83:@25567.4]
  wire [10:0] buffer_6_645; // @[Modules.scala 53:83:@25568.4]
  wire [11:0] _T_75862; // @[Modules.scala 53:83:@25570.4]
  wire [10:0] _T_75863; // @[Modules.scala 53:83:@25571.4]
  wire [10:0] buffer_6_646; // @[Modules.scala 53:83:@25572.4]
  wire [11:0] _T_75865; // @[Modules.scala 53:83:@25574.4]
  wire [10:0] _T_75866; // @[Modules.scala 53:83:@25575.4]
  wire [10:0] buffer_6_647; // @[Modules.scala 53:83:@25576.4]
  wire [11:0] _T_75868; // @[Modules.scala 53:83:@25578.4]
  wire [10:0] _T_75869; // @[Modules.scala 53:83:@25579.4]
  wire [10:0] buffer_6_648; // @[Modules.scala 53:83:@25580.4]
  wire [11:0] _T_75871; // @[Modules.scala 53:83:@25582.4]
  wire [10:0] _T_75872; // @[Modules.scala 53:83:@25583.4]
  wire [10:0] buffer_6_649; // @[Modules.scala 53:83:@25584.4]
  wire [11:0] _T_75874; // @[Modules.scala 53:83:@25586.4]
  wire [10:0] _T_75875; // @[Modules.scala 53:83:@25587.4]
  wire [10:0] buffer_6_650; // @[Modules.scala 53:83:@25588.4]
  wire [11:0] _T_75877; // @[Modules.scala 53:83:@25590.4]
  wire [10:0] _T_75878; // @[Modules.scala 53:83:@25591.4]
  wire [10:0] buffer_6_651; // @[Modules.scala 53:83:@25592.4]
  wire [11:0] _T_75880; // @[Modules.scala 53:83:@25594.4]
  wire [10:0] _T_75881; // @[Modules.scala 53:83:@25595.4]
  wire [10:0] buffer_6_652; // @[Modules.scala 53:83:@25596.4]
  wire [11:0] _T_75883; // @[Modules.scala 53:83:@25598.4]
  wire [10:0] _T_75884; // @[Modules.scala 53:83:@25599.4]
  wire [10:0] buffer_6_653; // @[Modules.scala 53:83:@25600.4]
  wire [11:0] _T_75889; // @[Modules.scala 53:83:@25606.4]
  wire [10:0] _T_75890; // @[Modules.scala 53:83:@25607.4]
  wire [10:0] buffer_6_655; // @[Modules.scala 53:83:@25608.4]
  wire [11:0] _T_75892; // @[Modules.scala 53:83:@25610.4]
  wire [10:0] _T_75893; // @[Modules.scala 53:83:@25611.4]
  wire [10:0] buffer_6_656; // @[Modules.scala 53:83:@25612.4]
  wire [11:0] _T_75895; // @[Modules.scala 53:83:@25614.4]
  wire [10:0] _T_75896; // @[Modules.scala 53:83:@25615.4]
  wire [10:0] buffer_6_657; // @[Modules.scala 53:83:@25616.4]
  wire [11:0] _T_75904; // @[Modules.scala 53:83:@25626.4]
  wire [10:0] _T_75905; // @[Modules.scala 53:83:@25627.4]
  wire [10:0] buffer_6_660; // @[Modules.scala 53:83:@25628.4]
  wire [11:0] _T_75907; // @[Modules.scala 53:83:@25630.4]
  wire [10:0] _T_75908; // @[Modules.scala 53:83:@25631.4]
  wire [10:0] buffer_6_661; // @[Modules.scala 53:83:@25632.4]
  wire [11:0] _T_75913; // @[Modules.scala 53:83:@25638.4]
  wire [10:0] _T_75914; // @[Modules.scala 53:83:@25639.4]
  wire [10:0] buffer_6_663; // @[Modules.scala 53:83:@25640.4]
  wire [11:0] _T_75916; // @[Modules.scala 53:83:@25642.4]
  wire [10:0] _T_75917; // @[Modules.scala 53:83:@25643.4]
  wire [10:0] buffer_6_664; // @[Modules.scala 53:83:@25644.4]
  wire [11:0] _T_75922; // @[Modules.scala 53:83:@25650.4]
  wire [10:0] _T_75923; // @[Modules.scala 53:83:@25651.4]
  wire [10:0] buffer_6_666; // @[Modules.scala 53:83:@25652.4]
  wire [11:0] _T_75925; // @[Modules.scala 53:83:@25654.4]
  wire [10:0] _T_75926; // @[Modules.scala 53:83:@25655.4]
  wire [10:0] buffer_6_667; // @[Modules.scala 53:83:@25656.4]
  wire [11:0] _T_75928; // @[Modules.scala 53:83:@25658.4]
  wire [10:0] _T_75929; // @[Modules.scala 53:83:@25659.4]
  wire [10:0] buffer_6_668; // @[Modules.scala 53:83:@25660.4]
  wire [11:0] _T_75931; // @[Modules.scala 53:83:@25662.4]
  wire [10:0] _T_75932; // @[Modules.scala 53:83:@25663.4]
  wire [10:0] buffer_6_669; // @[Modules.scala 53:83:@25664.4]
  wire [11:0] _T_75934; // @[Modules.scala 53:83:@25666.4]
  wire [10:0] _T_75935; // @[Modules.scala 53:83:@25667.4]
  wire [10:0] buffer_6_670; // @[Modules.scala 53:83:@25668.4]
  wire [11:0] _T_75937; // @[Modules.scala 53:83:@25670.4]
  wire [10:0] _T_75938; // @[Modules.scala 53:83:@25671.4]
  wire [10:0] buffer_6_671; // @[Modules.scala 53:83:@25672.4]
  wire [11:0] _T_75940; // @[Modules.scala 53:83:@25674.4]
  wire [10:0] _T_75941; // @[Modules.scala 53:83:@25675.4]
  wire [10:0] buffer_6_672; // @[Modules.scala 53:83:@25676.4]
  wire [11:0] _T_75943; // @[Modules.scala 53:83:@25678.4]
  wire [10:0] _T_75944; // @[Modules.scala 53:83:@25679.4]
  wire [10:0] buffer_6_673; // @[Modules.scala 53:83:@25680.4]
  wire [11:0] _T_75946; // @[Modules.scala 53:83:@25682.4]
  wire [10:0] _T_75947; // @[Modules.scala 53:83:@25683.4]
  wire [10:0] buffer_6_674; // @[Modules.scala 53:83:@25684.4]
  wire [11:0] _T_75949; // @[Modules.scala 53:83:@25686.4]
  wire [10:0] _T_75950; // @[Modules.scala 53:83:@25687.4]
  wire [10:0] buffer_6_675; // @[Modules.scala 53:83:@25688.4]
  wire [11:0] _T_75952; // @[Modules.scala 53:83:@25690.4]
  wire [10:0] _T_75953; // @[Modules.scala 53:83:@25691.4]
  wire [10:0] buffer_6_676; // @[Modules.scala 53:83:@25692.4]
  wire [11:0] _T_75955; // @[Modules.scala 53:83:@25694.4]
  wire [10:0] _T_75956; // @[Modules.scala 53:83:@25695.4]
  wire [10:0] buffer_6_677; // @[Modules.scala 53:83:@25696.4]
  wire [11:0] _T_75958; // @[Modules.scala 53:83:@25698.4]
  wire [10:0] _T_75959; // @[Modules.scala 53:83:@25699.4]
  wire [10:0] buffer_6_678; // @[Modules.scala 53:83:@25700.4]
  wire [11:0] _T_75961; // @[Modules.scala 53:83:@25702.4]
  wire [10:0] _T_75962; // @[Modules.scala 53:83:@25703.4]
  wire [10:0] buffer_6_679; // @[Modules.scala 53:83:@25704.4]
  wire [11:0] _T_75967; // @[Modules.scala 53:83:@25710.4]
  wire [10:0] _T_75968; // @[Modules.scala 53:83:@25711.4]
  wire [10:0] buffer_6_681; // @[Modules.scala 53:83:@25712.4]
  wire [11:0] _T_75970; // @[Modules.scala 53:83:@25714.4]
  wire [10:0] _T_75971; // @[Modules.scala 53:83:@25715.4]
  wire [10:0] buffer_6_682; // @[Modules.scala 53:83:@25716.4]
  wire [11:0] _T_75973; // @[Modules.scala 53:83:@25718.4]
  wire [10:0] _T_75974; // @[Modules.scala 53:83:@25719.4]
  wire [10:0] buffer_6_683; // @[Modules.scala 53:83:@25720.4]
  wire [11:0] _T_75976; // @[Modules.scala 53:83:@25722.4]
  wire [10:0] _T_75977; // @[Modules.scala 53:83:@25723.4]
  wire [10:0] buffer_6_684; // @[Modules.scala 53:83:@25724.4]
  wire [11:0] _T_75979; // @[Modules.scala 53:83:@25726.4]
  wire [10:0] _T_75980; // @[Modules.scala 53:83:@25727.4]
  wire [10:0] buffer_6_685; // @[Modules.scala 53:83:@25728.4]
  wire [11:0] _T_75982; // @[Modules.scala 56:109:@25730.4]
  wire [10:0] _T_75983; // @[Modules.scala 56:109:@25731.4]
  wire [10:0] buffer_6_686; // @[Modules.scala 56:109:@25732.4]
  wire [11:0] _T_75985; // @[Modules.scala 56:109:@25734.4]
  wire [10:0] _T_75986; // @[Modules.scala 56:109:@25735.4]
  wire [10:0] buffer_6_687; // @[Modules.scala 56:109:@25736.4]
  wire [11:0] _T_75988; // @[Modules.scala 56:109:@25738.4]
  wire [10:0] _T_75989; // @[Modules.scala 56:109:@25739.4]
  wire [10:0] buffer_6_688; // @[Modules.scala 56:109:@25740.4]
  wire [11:0] _T_75991; // @[Modules.scala 56:109:@25742.4]
  wire [10:0] _T_75992; // @[Modules.scala 56:109:@25743.4]
  wire [10:0] buffer_6_689; // @[Modules.scala 56:109:@25744.4]
  wire [11:0] _T_75997; // @[Modules.scala 56:109:@25750.4]
  wire [10:0] _T_75998; // @[Modules.scala 56:109:@25751.4]
  wire [10:0] buffer_6_691; // @[Modules.scala 56:109:@25752.4]
  wire [11:0] _T_76000; // @[Modules.scala 56:109:@25754.4]
  wire [10:0] _T_76001; // @[Modules.scala 56:109:@25755.4]
  wire [10:0] buffer_6_692; // @[Modules.scala 56:109:@25756.4]
  wire [11:0] _T_76003; // @[Modules.scala 56:109:@25758.4]
  wire [10:0] _T_76004; // @[Modules.scala 56:109:@25759.4]
  wire [10:0] buffer_6_693; // @[Modules.scala 56:109:@25760.4]
  wire [11:0] _T_76006; // @[Modules.scala 56:109:@25762.4]
  wire [10:0] _T_76007; // @[Modules.scala 56:109:@25763.4]
  wire [10:0] buffer_6_694; // @[Modules.scala 56:109:@25764.4]
  wire [11:0] _T_76009; // @[Modules.scala 56:109:@25766.4]
  wire [10:0] _T_76010; // @[Modules.scala 56:109:@25767.4]
  wire [10:0] buffer_6_695; // @[Modules.scala 56:109:@25768.4]
  wire [11:0] _T_76012; // @[Modules.scala 56:109:@25770.4]
  wire [10:0] _T_76013; // @[Modules.scala 56:109:@25771.4]
  wire [10:0] buffer_6_696; // @[Modules.scala 56:109:@25772.4]
  wire [11:0] _T_76015; // @[Modules.scala 56:109:@25774.4]
  wire [10:0] _T_76016; // @[Modules.scala 56:109:@25775.4]
  wire [10:0] buffer_6_697; // @[Modules.scala 56:109:@25776.4]
  wire [11:0] _T_76018; // @[Modules.scala 56:109:@25778.4]
  wire [10:0] _T_76019; // @[Modules.scala 56:109:@25779.4]
  wire [10:0] buffer_6_698; // @[Modules.scala 56:109:@25780.4]
  wire [11:0] _T_76021; // @[Modules.scala 56:109:@25782.4]
  wire [10:0] _T_76022; // @[Modules.scala 56:109:@25783.4]
  wire [10:0] buffer_6_699; // @[Modules.scala 56:109:@25784.4]
  wire [11:0] _T_76024; // @[Modules.scala 56:109:@25786.4]
  wire [10:0] _T_76025; // @[Modules.scala 56:109:@25787.4]
  wire [10:0] buffer_6_700; // @[Modules.scala 56:109:@25788.4]
  wire [11:0] _T_76027; // @[Modules.scala 56:109:@25790.4]
  wire [10:0] _T_76028; // @[Modules.scala 56:109:@25791.4]
  wire [10:0] buffer_6_701; // @[Modules.scala 56:109:@25792.4]
  wire [11:0] _T_76030; // @[Modules.scala 56:109:@25794.4]
  wire [10:0] _T_76031; // @[Modules.scala 56:109:@25795.4]
  wire [10:0] buffer_6_702; // @[Modules.scala 56:109:@25796.4]
  wire [11:0] _T_76033; // @[Modules.scala 56:109:@25798.4]
  wire [10:0] _T_76034; // @[Modules.scala 56:109:@25799.4]
  wire [10:0] buffer_6_703; // @[Modules.scala 56:109:@25800.4]
  wire [11:0] _T_76036; // @[Modules.scala 56:109:@25802.4]
  wire [10:0] _T_76037; // @[Modules.scala 56:109:@25803.4]
  wire [10:0] buffer_6_704; // @[Modules.scala 56:109:@25804.4]
  wire [11:0] _T_76039; // @[Modules.scala 56:109:@25806.4]
  wire [10:0] _T_76040; // @[Modules.scala 56:109:@25807.4]
  wire [10:0] buffer_6_705; // @[Modules.scala 56:109:@25808.4]
  wire [11:0] _T_76042; // @[Modules.scala 56:109:@25810.4]
  wire [10:0] _T_76043; // @[Modules.scala 56:109:@25811.4]
  wire [10:0] buffer_6_706; // @[Modules.scala 56:109:@25812.4]
  wire [11:0] _T_76045; // @[Modules.scala 56:109:@25814.4]
  wire [10:0] _T_76046; // @[Modules.scala 56:109:@25815.4]
  wire [10:0] buffer_6_707; // @[Modules.scala 56:109:@25816.4]
  wire [11:0] _T_76048; // @[Modules.scala 56:109:@25818.4]
  wire [10:0] _T_76049; // @[Modules.scala 56:109:@25819.4]
  wire [10:0] buffer_6_708; // @[Modules.scala 56:109:@25820.4]
  wire [11:0] _T_76051; // @[Modules.scala 56:109:@25822.4]
  wire [10:0] _T_76052; // @[Modules.scala 56:109:@25823.4]
  wire [10:0] buffer_6_709; // @[Modules.scala 56:109:@25824.4]
  wire [11:0] _T_76054; // @[Modules.scala 56:109:@25826.4]
  wire [10:0] _T_76055; // @[Modules.scala 56:109:@25827.4]
  wire [10:0] buffer_6_710; // @[Modules.scala 56:109:@25828.4]
  wire [11:0] _T_76057; // @[Modules.scala 56:109:@25830.4]
  wire [10:0] _T_76058; // @[Modules.scala 56:109:@25831.4]
  wire [10:0] buffer_6_711; // @[Modules.scala 56:109:@25832.4]
  wire [11:0] _T_76060; // @[Modules.scala 56:109:@25834.4]
  wire [10:0] _T_76061; // @[Modules.scala 56:109:@25835.4]
  wire [10:0] buffer_6_712; // @[Modules.scala 56:109:@25836.4]
  wire [11:0] _T_76063; // @[Modules.scala 56:109:@25838.4]
  wire [10:0] _T_76064; // @[Modules.scala 56:109:@25839.4]
  wire [10:0] buffer_6_713; // @[Modules.scala 56:109:@25840.4]
  wire [11:0] _T_76066; // @[Modules.scala 56:109:@25842.4]
  wire [10:0] _T_76067; // @[Modules.scala 56:109:@25843.4]
  wire [10:0] buffer_6_714; // @[Modules.scala 56:109:@25844.4]
  wire [11:0] _T_76069; // @[Modules.scala 56:109:@25846.4]
  wire [10:0] _T_76070; // @[Modules.scala 56:109:@25847.4]
  wire [10:0] buffer_6_715; // @[Modules.scala 56:109:@25848.4]
  wire [11:0] _T_76072; // @[Modules.scala 56:109:@25850.4]
  wire [10:0] _T_76073; // @[Modules.scala 56:109:@25851.4]
  wire [10:0] buffer_6_716; // @[Modules.scala 56:109:@25852.4]
  wire [11:0] _T_76075; // @[Modules.scala 56:109:@25854.4]
  wire [10:0] _T_76076; // @[Modules.scala 56:109:@25855.4]
  wire [10:0] buffer_6_717; // @[Modules.scala 56:109:@25856.4]
  wire [11:0] _T_76078; // @[Modules.scala 56:109:@25858.4]
  wire [10:0] _T_76079; // @[Modules.scala 56:109:@25859.4]
  wire [10:0] buffer_6_718; // @[Modules.scala 56:109:@25860.4]
  wire [11:0] _T_76081; // @[Modules.scala 56:109:@25862.4]
  wire [10:0] _T_76082; // @[Modules.scala 56:109:@25863.4]
  wire [10:0] buffer_6_719; // @[Modules.scala 56:109:@25864.4]
  wire [11:0] _T_76084; // @[Modules.scala 56:109:@25866.4]
  wire [10:0] _T_76085; // @[Modules.scala 56:109:@25867.4]
  wire [10:0] buffer_6_720; // @[Modules.scala 56:109:@25868.4]
  wire [11:0] _T_76087; // @[Modules.scala 56:109:@25870.4]
  wire [10:0] _T_76088; // @[Modules.scala 56:109:@25871.4]
  wire [10:0] buffer_6_721; // @[Modules.scala 56:109:@25872.4]
  wire [11:0] _T_76090; // @[Modules.scala 56:109:@25874.4]
  wire [10:0] _T_76091; // @[Modules.scala 56:109:@25875.4]
  wire [10:0] buffer_6_722; // @[Modules.scala 56:109:@25876.4]
  wire [11:0] _T_76093; // @[Modules.scala 56:109:@25878.4]
  wire [10:0] _T_76094; // @[Modules.scala 56:109:@25879.4]
  wire [10:0] buffer_6_723; // @[Modules.scala 56:109:@25880.4]
  wire [11:0] _T_76096; // @[Modules.scala 56:109:@25882.4]
  wire [10:0] _T_76097; // @[Modules.scala 56:109:@25883.4]
  wire [10:0] buffer_6_724; // @[Modules.scala 56:109:@25884.4]
  wire [11:0] _T_76099; // @[Modules.scala 56:109:@25886.4]
  wire [10:0] _T_76100; // @[Modules.scala 56:109:@25887.4]
  wire [10:0] buffer_6_725; // @[Modules.scala 56:109:@25888.4]
  wire [11:0] _T_76102; // @[Modules.scala 56:109:@25890.4]
  wire [10:0] _T_76103; // @[Modules.scala 56:109:@25891.4]
  wire [10:0] buffer_6_726; // @[Modules.scala 56:109:@25892.4]
  wire [11:0] _T_76105; // @[Modules.scala 56:109:@25894.4]
  wire [10:0] _T_76106; // @[Modules.scala 56:109:@25895.4]
  wire [10:0] buffer_6_727; // @[Modules.scala 56:109:@25896.4]
  wire [11:0] _T_76108; // @[Modules.scala 56:109:@25898.4]
  wire [10:0] _T_76109; // @[Modules.scala 56:109:@25899.4]
  wire [10:0] buffer_6_728; // @[Modules.scala 56:109:@25900.4]
  wire [11:0] _T_76111; // @[Modules.scala 56:109:@25902.4]
  wire [10:0] _T_76112; // @[Modules.scala 56:109:@25903.4]
  wire [10:0] buffer_6_729; // @[Modules.scala 56:109:@25904.4]
  wire [11:0] _T_76114; // @[Modules.scala 56:109:@25906.4]
  wire [10:0] _T_76115; // @[Modules.scala 56:109:@25907.4]
  wire [10:0] buffer_6_730; // @[Modules.scala 56:109:@25908.4]
  wire [11:0] _T_76117; // @[Modules.scala 56:109:@25910.4]
  wire [10:0] _T_76118; // @[Modules.scala 56:109:@25911.4]
  wire [10:0] buffer_6_731; // @[Modules.scala 56:109:@25912.4]
  wire [11:0] _T_76120; // @[Modules.scala 56:109:@25914.4]
  wire [10:0] _T_76121; // @[Modules.scala 56:109:@25915.4]
  wire [10:0] buffer_6_732; // @[Modules.scala 56:109:@25916.4]
  wire [11:0] _T_76123; // @[Modules.scala 56:109:@25918.4]
  wire [10:0] _T_76124; // @[Modules.scala 56:109:@25919.4]
  wire [10:0] buffer_6_733; // @[Modules.scala 56:109:@25920.4]
  wire [11:0] _T_76126; // @[Modules.scala 56:109:@25922.4]
  wire [10:0] _T_76127; // @[Modules.scala 56:109:@25923.4]
  wire [10:0] buffer_6_734; // @[Modules.scala 56:109:@25924.4]
  wire [11:0] _T_76129; // @[Modules.scala 63:156:@25927.4]
  wire [10:0] _T_76130; // @[Modules.scala 63:156:@25928.4]
  wire [10:0] buffer_6_736; // @[Modules.scala 63:156:@25929.4]
  wire [11:0] _T_76132; // @[Modules.scala 63:156:@25931.4]
  wire [10:0] _T_76133; // @[Modules.scala 63:156:@25932.4]
  wire [10:0] buffer_6_737; // @[Modules.scala 63:156:@25933.4]
  wire [11:0] _T_76135; // @[Modules.scala 63:156:@25935.4]
  wire [10:0] _T_76136; // @[Modules.scala 63:156:@25936.4]
  wire [10:0] buffer_6_738; // @[Modules.scala 63:156:@25937.4]
  wire [11:0] _T_76138; // @[Modules.scala 63:156:@25939.4]
  wire [10:0] _T_76139; // @[Modules.scala 63:156:@25940.4]
  wire [10:0] buffer_6_739; // @[Modules.scala 63:156:@25941.4]
  wire [11:0] _T_76141; // @[Modules.scala 63:156:@25943.4]
  wire [10:0] _T_76142; // @[Modules.scala 63:156:@25944.4]
  wire [10:0] buffer_6_740; // @[Modules.scala 63:156:@25945.4]
  wire [11:0] _T_76144; // @[Modules.scala 63:156:@25947.4]
  wire [10:0] _T_76145; // @[Modules.scala 63:156:@25948.4]
  wire [10:0] buffer_6_741; // @[Modules.scala 63:156:@25949.4]
  wire [11:0] _T_76147; // @[Modules.scala 63:156:@25951.4]
  wire [10:0] _T_76148; // @[Modules.scala 63:156:@25952.4]
  wire [10:0] buffer_6_742; // @[Modules.scala 63:156:@25953.4]
  wire [11:0] _T_76150; // @[Modules.scala 63:156:@25955.4]
  wire [10:0] _T_76151; // @[Modules.scala 63:156:@25956.4]
  wire [10:0] buffer_6_743; // @[Modules.scala 63:156:@25957.4]
  wire [11:0] _T_76153; // @[Modules.scala 63:156:@25959.4]
  wire [10:0] _T_76154; // @[Modules.scala 63:156:@25960.4]
  wire [10:0] buffer_6_744; // @[Modules.scala 63:156:@25961.4]
  wire [11:0] _T_76156; // @[Modules.scala 63:156:@25963.4]
  wire [10:0] _T_76157; // @[Modules.scala 63:156:@25964.4]
  wire [10:0] buffer_6_745; // @[Modules.scala 63:156:@25965.4]
  wire [11:0] _T_76159; // @[Modules.scala 63:156:@25967.4]
  wire [10:0] _T_76160; // @[Modules.scala 63:156:@25968.4]
  wire [10:0] buffer_6_746; // @[Modules.scala 63:156:@25969.4]
  wire [11:0] _T_76162; // @[Modules.scala 63:156:@25971.4]
  wire [10:0] _T_76163; // @[Modules.scala 63:156:@25972.4]
  wire [10:0] buffer_6_747; // @[Modules.scala 63:156:@25973.4]
  wire [11:0] _T_76165; // @[Modules.scala 63:156:@25975.4]
  wire [10:0] _T_76166; // @[Modules.scala 63:156:@25976.4]
  wire [10:0] buffer_6_748; // @[Modules.scala 63:156:@25977.4]
  wire [11:0] _T_76168; // @[Modules.scala 63:156:@25979.4]
  wire [10:0] _T_76169; // @[Modules.scala 63:156:@25980.4]
  wire [10:0] buffer_6_749; // @[Modules.scala 63:156:@25981.4]
  wire [11:0] _T_76171; // @[Modules.scala 63:156:@25983.4]
  wire [10:0] _T_76172; // @[Modules.scala 63:156:@25984.4]
  wire [10:0] buffer_6_750; // @[Modules.scala 63:156:@25985.4]
  wire [11:0] _T_76174; // @[Modules.scala 63:156:@25987.4]
  wire [10:0] _T_76175; // @[Modules.scala 63:156:@25988.4]
  wire [10:0] buffer_6_751; // @[Modules.scala 63:156:@25989.4]
  wire [11:0] _T_76177; // @[Modules.scala 63:156:@25991.4]
  wire [10:0] _T_76178; // @[Modules.scala 63:156:@25992.4]
  wire [10:0] buffer_6_752; // @[Modules.scala 63:156:@25993.4]
  wire [11:0] _T_76180; // @[Modules.scala 63:156:@25995.4]
  wire [10:0] _T_76181; // @[Modules.scala 63:156:@25996.4]
  wire [10:0] buffer_6_753; // @[Modules.scala 63:156:@25997.4]
  wire [11:0] _T_76183; // @[Modules.scala 63:156:@25999.4]
  wire [10:0] _T_76184; // @[Modules.scala 63:156:@26000.4]
  wire [10:0] buffer_6_754; // @[Modules.scala 63:156:@26001.4]
  wire [11:0] _T_76186; // @[Modules.scala 63:156:@26003.4]
  wire [10:0] _T_76187; // @[Modules.scala 63:156:@26004.4]
  wire [10:0] buffer_6_755; // @[Modules.scala 63:156:@26005.4]
  wire [11:0] _T_76189; // @[Modules.scala 63:156:@26007.4]
  wire [10:0] _T_76190; // @[Modules.scala 63:156:@26008.4]
  wire [10:0] buffer_6_756; // @[Modules.scala 63:156:@26009.4]
  wire [11:0] _T_76192; // @[Modules.scala 63:156:@26011.4]
  wire [10:0] _T_76193; // @[Modules.scala 63:156:@26012.4]
  wire [10:0] buffer_6_757; // @[Modules.scala 63:156:@26013.4]
  wire [11:0] _T_76195; // @[Modules.scala 63:156:@26015.4]
  wire [10:0] _T_76196; // @[Modules.scala 63:156:@26016.4]
  wire [10:0] buffer_6_758; // @[Modules.scala 63:156:@26017.4]
  wire [11:0] _T_76198; // @[Modules.scala 63:156:@26019.4]
  wire [10:0] _T_76199; // @[Modules.scala 63:156:@26020.4]
  wire [10:0] buffer_6_759; // @[Modules.scala 63:156:@26021.4]
  wire [11:0] _T_76201; // @[Modules.scala 63:156:@26023.4]
  wire [10:0] _T_76202; // @[Modules.scala 63:156:@26024.4]
  wire [10:0] buffer_6_760; // @[Modules.scala 63:156:@26025.4]
  wire [11:0] _T_76204; // @[Modules.scala 63:156:@26027.4]
  wire [10:0] _T_76205; // @[Modules.scala 63:156:@26028.4]
  wire [10:0] buffer_6_761; // @[Modules.scala 63:156:@26029.4]
  wire [11:0] _T_76207; // @[Modules.scala 63:156:@26031.4]
  wire [10:0] _T_76208; // @[Modules.scala 63:156:@26032.4]
  wire [10:0] buffer_6_762; // @[Modules.scala 63:156:@26033.4]
  wire [11:0] _T_76210; // @[Modules.scala 63:156:@26035.4]
  wire [10:0] _T_76211; // @[Modules.scala 63:156:@26036.4]
  wire [10:0] buffer_6_763; // @[Modules.scala 63:156:@26037.4]
  wire [11:0] _T_76213; // @[Modules.scala 63:156:@26039.4]
  wire [10:0] _T_76214; // @[Modules.scala 63:156:@26040.4]
  wire [10:0] buffer_6_764; // @[Modules.scala 63:156:@26041.4]
  wire [11:0] _T_76216; // @[Modules.scala 63:156:@26043.4]
  wire [10:0] _T_76217; // @[Modules.scala 63:156:@26044.4]
  wire [10:0] buffer_6_765; // @[Modules.scala 63:156:@26045.4]
  wire [11:0] _T_76219; // @[Modules.scala 63:156:@26047.4]
  wire [10:0] _T_76220; // @[Modules.scala 63:156:@26048.4]
  wire [10:0] buffer_6_766; // @[Modules.scala 63:156:@26049.4]
  wire [11:0] _T_76222; // @[Modules.scala 63:156:@26051.4]
  wire [10:0] _T_76223; // @[Modules.scala 63:156:@26052.4]
  wire [10:0] buffer_6_767; // @[Modules.scala 63:156:@26053.4]
  wire [11:0] _T_76225; // @[Modules.scala 63:156:@26055.4]
  wire [10:0] _T_76226; // @[Modules.scala 63:156:@26056.4]
  wire [10:0] buffer_6_768; // @[Modules.scala 63:156:@26057.4]
  wire [11:0] _T_76228; // @[Modules.scala 63:156:@26059.4]
  wire [10:0] _T_76229; // @[Modules.scala 63:156:@26060.4]
  wire [10:0] buffer_6_769; // @[Modules.scala 63:156:@26061.4]
  wire [11:0] _T_76231; // @[Modules.scala 63:156:@26063.4]
  wire [10:0] _T_76232; // @[Modules.scala 63:156:@26064.4]
  wire [10:0] buffer_6_770; // @[Modules.scala 63:156:@26065.4]
  wire [11:0] _T_76234; // @[Modules.scala 63:156:@26067.4]
  wire [10:0] _T_76235; // @[Modules.scala 63:156:@26068.4]
  wire [10:0] buffer_6_771; // @[Modules.scala 63:156:@26069.4]
  wire [11:0] _T_76237; // @[Modules.scala 63:156:@26071.4]
  wire [10:0] _T_76238; // @[Modules.scala 63:156:@26072.4]
  wire [10:0] buffer_6_772; // @[Modules.scala 63:156:@26073.4]
  wire [11:0] _T_76240; // @[Modules.scala 63:156:@26075.4]
  wire [10:0] _T_76241; // @[Modules.scala 63:156:@26076.4]
  wire [10:0] buffer_6_773; // @[Modules.scala 63:156:@26077.4]
  wire [11:0] _T_76243; // @[Modules.scala 63:156:@26079.4]
  wire [10:0] _T_76244; // @[Modules.scala 63:156:@26080.4]
  wire [10:0] buffer_6_774; // @[Modules.scala 63:156:@26081.4]
  wire [11:0] _T_76246; // @[Modules.scala 63:156:@26083.4]
  wire [10:0] _T_76247; // @[Modules.scala 63:156:@26084.4]
  wire [10:0] buffer_6_775; // @[Modules.scala 63:156:@26085.4]
  wire [11:0] _T_76249; // @[Modules.scala 63:156:@26087.4]
  wire [10:0] _T_76250; // @[Modules.scala 63:156:@26088.4]
  wire [10:0] buffer_6_776; // @[Modules.scala 63:156:@26089.4]
  wire [11:0] _T_76252; // @[Modules.scala 63:156:@26091.4]
  wire [10:0] _T_76253; // @[Modules.scala 63:156:@26092.4]
  wire [10:0] buffer_6_777; // @[Modules.scala 63:156:@26093.4]
  wire [11:0] _T_76255; // @[Modules.scala 63:156:@26095.4]
  wire [10:0] _T_76256; // @[Modules.scala 63:156:@26096.4]
  wire [10:0] buffer_6_778; // @[Modules.scala 63:156:@26097.4]
  wire [11:0] _T_76258; // @[Modules.scala 63:156:@26099.4]
  wire [10:0] _T_76259; // @[Modules.scala 63:156:@26100.4]
  wire [10:0] buffer_6_779; // @[Modules.scala 63:156:@26101.4]
  wire [11:0] _T_76261; // @[Modules.scala 63:156:@26103.4]
  wire [10:0] _T_76262; // @[Modules.scala 63:156:@26104.4]
  wire [10:0] buffer_6_780; // @[Modules.scala 63:156:@26105.4]
  wire [11:0] _T_76264; // @[Modules.scala 63:156:@26107.4]
  wire [10:0] _T_76265; // @[Modules.scala 63:156:@26108.4]
  wire [10:0] buffer_6_781; // @[Modules.scala 63:156:@26109.4]
  wire [11:0] _T_76267; // @[Modules.scala 63:156:@26111.4]
  wire [10:0] _T_76268; // @[Modules.scala 63:156:@26112.4]
  wire [10:0] buffer_6_782; // @[Modules.scala 63:156:@26113.4]
  wire [11:0] _T_76270; // @[Modules.scala 63:156:@26115.4]
  wire [10:0] _T_76271; // @[Modules.scala 63:156:@26116.4]
  wire [10:0] buffer_6_783; // @[Modules.scala 63:156:@26117.4]
  wire [5:0] _T_76273; // @[Modules.scala 37:46:@26120.4]
  wire [4:0] _T_76274; // @[Modules.scala 37:46:@26121.4]
  wire [4:0] _T_76275; // @[Modules.scala 37:46:@26122.4]
  wire [5:0] _T_76317; // @[Modules.scala 43:47:@26167.4]
  wire [4:0] _T_76318; // @[Modules.scala 43:47:@26168.4]
  wire [4:0] _T_76319; // @[Modules.scala 43:47:@26169.4]
  wire [5:0] _T_76331; // @[Modules.scala 46:47:@26181.4]
  wire [4:0] _T_76332; // @[Modules.scala 46:47:@26182.4]
  wire [4:0] _T_76333; // @[Modules.scala 46:47:@26183.4]
  wire [5:0] _T_76372; // @[Modules.scala 43:47:@26224.4]
  wire [4:0] _T_76373; // @[Modules.scala 43:47:@26225.4]
  wire [4:0] _T_76374; // @[Modules.scala 43:47:@26226.4]
  wire [5:0] _T_76410; // @[Modules.scala 37:46:@26270.4]
  wire [4:0] _T_76411; // @[Modules.scala 37:46:@26271.4]
  wire [4:0] _T_76412; // @[Modules.scala 37:46:@26272.4]
  wire [5:0] _T_76562; // @[Modules.scala 40:46:@26447.4]
  wire [4:0] _T_76563; // @[Modules.scala 40:46:@26448.4]
  wire [4:0] _T_76564; // @[Modules.scala 40:46:@26449.4]
  wire [5:0] _T_76625; // @[Modules.scala 40:46:@26517.4]
  wire [4:0] _T_76626; // @[Modules.scala 40:46:@26518.4]
  wire [4:0] _T_76627; // @[Modules.scala 40:46:@26519.4]
  wire [5:0] _T_76666; // @[Modules.scala 43:47:@26567.4]
  wire [4:0] _T_76667; // @[Modules.scala 43:47:@26568.4]
  wire [4:0] _T_76668; // @[Modules.scala 43:47:@26569.4]
  wire [5:0] _T_76680; // @[Modules.scala 43:47:@26581.4]
  wire [4:0] _T_76681; // @[Modules.scala 43:47:@26582.4]
  wire [4:0] _T_76682; // @[Modules.scala 43:47:@26583.4]
  wire [5:0] _T_76781; // @[Modules.scala 37:46:@26690.4]
  wire [4:0] _T_76782; // @[Modules.scala 37:46:@26691.4]
  wire [4:0] _T_76783; // @[Modules.scala 37:46:@26692.4]
  wire [5:0] _T_76825; // @[Modules.scala 43:47:@26737.4]
  wire [4:0] _T_76826; // @[Modules.scala 43:47:@26738.4]
  wire [4:0] _T_76827; // @[Modules.scala 43:47:@26739.4]
  wire [5:0] _T_76828; // @[Modules.scala 40:46:@26741.4]
  wire [4:0] _T_76829; // @[Modules.scala 40:46:@26742.4]
  wire [4:0] _T_76830; // @[Modules.scala 40:46:@26743.4]
  wire [5:0] _T_76945; // @[Modules.scala 43:47:@26862.4]
  wire [4:0] _T_76946; // @[Modules.scala 43:47:@26863.4]
  wire [4:0] _T_76947; // @[Modules.scala 43:47:@26864.4]
  wire [5:0] _T_76971; // @[Modules.scala 37:46:@26892.4]
  wire [4:0] _T_76972; // @[Modules.scala 37:46:@26893.4]
  wire [4:0] _T_76973; // @[Modules.scala 37:46:@26894.4]
  wire [5:0] _T_76974; // @[Modules.scala 37:46:@26896.4]
  wire [4:0] _T_76975; // @[Modules.scala 37:46:@26897.4]
  wire [4:0] _T_76976; // @[Modules.scala 37:46:@26898.4]
  wire [5:0] _T_76977; // @[Modules.scala 40:46:@26900.4]
  wire [4:0] _T_76978; // @[Modules.scala 40:46:@26901.4]
  wire [4:0] _T_76979; // @[Modules.scala 40:46:@26902.4]
  wire [5:0] _T_76983; // @[Modules.scala 40:46:@26908.4]
  wire [4:0] _T_76984; // @[Modules.scala 40:46:@26909.4]
  wire [4:0] _T_76985; // @[Modules.scala 40:46:@26910.4]
  wire [5:0] _T_77041; // @[Modules.scala 37:46:@26969.4]
  wire [4:0] _T_77042; // @[Modules.scala 37:46:@26970.4]
  wire [4:0] _T_77043; // @[Modules.scala 37:46:@26971.4]
  wire [5:0] _T_77117; // @[Modules.scala 46:47:@27047.4]
  wire [4:0] _T_77118; // @[Modules.scala 46:47:@27048.4]
  wire [4:0] _T_77119; // @[Modules.scala 46:47:@27049.4]
  wire [5:0] _T_77191; // @[Modules.scala 37:46:@27127.4]
  wire [4:0] _T_77192; // @[Modules.scala 37:46:@27128.4]
  wire [4:0] _T_77193; // @[Modules.scala 37:46:@27129.4]
  wire [5:0] _T_77234; // @[Modules.scala 43:47:@27175.4]
  wire [4:0] _T_77235; // @[Modules.scala 43:47:@27176.4]
  wire [4:0] _T_77236; // @[Modules.scala 43:47:@27177.4]
  wire [5:0] _T_77271; // @[Modules.scala 40:46:@27215.4]
  wire [4:0] _T_77272; // @[Modules.scala 40:46:@27216.4]
  wire [4:0] _T_77273; // @[Modules.scala 40:46:@27217.4]
  wire [5:0] _T_77274; // @[Modules.scala 40:46:@27219.4]
  wire [4:0] _T_77275; // @[Modules.scala 40:46:@27220.4]
  wire [4:0] _T_77276; // @[Modules.scala 40:46:@27221.4]
  wire [5:0] _T_77389; // @[Modules.scala 46:47:@27349.4]
  wire [4:0] _T_77390; // @[Modules.scala 46:47:@27350.4]
  wire [4:0] _T_77391; // @[Modules.scala 46:47:@27351.4]
  wire [5:0] _T_77396; // @[Modules.scala 43:47:@27356.4]
  wire [4:0] _T_77397; // @[Modules.scala 43:47:@27357.4]
  wire [4:0] _T_77398; // @[Modules.scala 43:47:@27358.4]
  wire [5:0] _T_77443; // @[Modules.scala 43:47:@27407.4]
  wire [4:0] _T_77444; // @[Modules.scala 43:47:@27408.4]
  wire [4:0] _T_77445; // @[Modules.scala 43:47:@27409.4]
  wire [5:0] _T_77467; // @[Modules.scala 46:37:@27433.4]
  wire [4:0] _T_77468; // @[Modules.scala 46:37:@27434.4]
  wire [4:0] _T_77469; // @[Modules.scala 46:37:@27435.4]
  wire [5:0] _T_77470; // @[Modules.scala 46:47:@27436.4]
  wire [4:0] _T_77471; // @[Modules.scala 46:47:@27437.4]
  wire [4:0] _T_77472; // @[Modules.scala 46:47:@27438.4]
  wire [5:0] _T_77473; // @[Modules.scala 40:46:@27440.4]
  wire [4:0] _T_77474; // @[Modules.scala 40:46:@27441.4]
  wire [4:0] _T_77475; // @[Modules.scala 40:46:@27442.4]
  wire [5:0] _T_77502; // @[Modules.scala 46:47:@27474.4]
  wire [4:0] _T_77503; // @[Modules.scala 46:47:@27475.4]
  wire [4:0] _T_77504; // @[Modules.scala 46:47:@27476.4]
  wire [5:0] _T_77522; // @[Modules.scala 40:46:@27496.4]
  wire [4:0] _T_77523; // @[Modules.scala 40:46:@27497.4]
  wire [4:0] _T_77524; // @[Modules.scala 40:46:@27498.4]
  wire [5:0] _T_77567; // @[Modules.scala 40:46:@27549.4]
  wire [4:0] _T_77568; // @[Modules.scala 40:46:@27550.4]
  wire [4:0] _T_77569; // @[Modules.scala 40:46:@27551.4]
  wire [5:0] _T_77574; // @[Modules.scala 43:47:@27556.4]
  wire [4:0] _T_77575; // @[Modules.scala 43:47:@27557.4]
  wire [4:0] _T_77576; // @[Modules.scala 43:47:@27558.4]
  wire [5:0] _T_77604; // @[Modules.scala 40:46:@27589.4]
  wire [4:0] _T_77605; // @[Modules.scala 40:46:@27590.4]
  wire [4:0] _T_77606; // @[Modules.scala 40:46:@27591.4]
  wire [5:0] _T_77629; // @[Modules.scala 43:47:@27620.4]
  wire [4:0] _T_77630; // @[Modules.scala 43:47:@27621.4]
  wire [4:0] _T_77631; // @[Modules.scala 43:47:@27622.4]
  wire [5:0] _T_77692; // @[Modules.scala 40:46:@27697.4]
  wire [4:0] _T_77693; // @[Modules.scala 40:46:@27698.4]
  wire [4:0] _T_77694; // @[Modules.scala 40:46:@27699.4]
  wire [5:0] _T_77730; // @[Modules.scala 43:47:@27736.4]
  wire [4:0] _T_77731; // @[Modules.scala 43:47:@27737.4]
  wire [4:0] _T_77732; // @[Modules.scala 43:47:@27738.4]
  wire [5:0] _T_77744; // @[Modules.scala 43:47:@27750.4]
  wire [4:0] _T_77745; // @[Modules.scala 43:47:@27751.4]
  wire [4:0] _T_77746; // @[Modules.scala 43:47:@27752.4]
  wire [5:0] _T_77774; // @[Modules.scala 46:47:@27783.4]
  wire [4:0] _T_77775; // @[Modules.scala 46:47:@27784.4]
  wire [4:0] _T_77776; // @[Modules.scala 46:47:@27785.4]
  wire [5:0] _T_77794; // @[Modules.scala 40:46:@27805.4]
  wire [4:0] _T_77795; // @[Modules.scala 40:46:@27806.4]
  wire [4:0] _T_77796; // @[Modules.scala 40:46:@27807.4]
  wire [5:0] _T_77960; // @[Modules.scala 43:47:@27989.4]
  wire [4:0] _T_77961; // @[Modules.scala 43:47:@27990.4]
  wire [4:0] _T_77962; // @[Modules.scala 43:47:@27991.4]
  wire [5:0] _T_78189; // @[Modules.scala 43:47:@28222.4]
  wire [4:0] _T_78190; // @[Modules.scala 43:47:@28223.4]
  wire [4:0] _T_78191; // @[Modules.scala 43:47:@28224.4]
  wire [5:0] _T_78255; // @[Modules.scala 37:46:@28289.4]
  wire [4:0] _T_78256; // @[Modules.scala 37:46:@28290.4]
  wire [4:0] _T_78257; // @[Modules.scala 37:46:@28291.4]
  wire [10:0] buffer_7_0; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78265; // @[Modules.scala 50:57:@28300.4]
  wire [10:0] _T_78266; // @[Modules.scala 50:57:@28301.4]
  wire [10:0] buffer_7_392; // @[Modules.scala 50:57:@28302.4]
  wire [11:0] _T_78268; // @[Modules.scala 50:57:@28304.4]
  wire [10:0] _T_78269; // @[Modules.scala 50:57:@28305.4]
  wire [10:0] buffer_7_393; // @[Modules.scala 50:57:@28306.4]
  wire [10:0] buffer_7_8; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78277; // @[Modules.scala 50:57:@28316.4]
  wire [10:0] _T_78278; // @[Modules.scala 50:57:@28317.4]
  wire [10:0] buffer_7_396; // @[Modules.scala 50:57:@28318.4]
  wire [10:0] buffer_7_10; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78280; // @[Modules.scala 50:57:@28320.4]
  wire [10:0] _T_78281; // @[Modules.scala 50:57:@28321.4]
  wire [10:0] buffer_7_397; // @[Modules.scala 50:57:@28322.4]
  wire [11:0] _T_78286; // @[Modules.scala 50:57:@28328.4]
  wire [10:0] _T_78287; // @[Modules.scala 50:57:@28329.4]
  wire [10:0] buffer_7_399; // @[Modules.scala 50:57:@28330.4]
  wire [10:0] buffer_7_17; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78289; // @[Modules.scala 50:57:@28332.4]
  wire [10:0] _T_78290; // @[Modules.scala 50:57:@28333.4]
  wire [10:0] buffer_7_400; // @[Modules.scala 50:57:@28334.4]
  wire [10:0] buffer_7_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78304; // @[Modules.scala 50:57:@28352.4]
  wire [10:0] _T_78305; // @[Modules.scala 50:57:@28353.4]
  wire [10:0] buffer_7_405; // @[Modules.scala 50:57:@28354.4]
  wire [11:0] _T_78310; // @[Modules.scala 50:57:@28360.4]
  wire [10:0] _T_78311; // @[Modules.scala 50:57:@28361.4]
  wire [10:0] buffer_7_407; // @[Modules.scala 50:57:@28362.4]
  wire [11:0] _T_78337; // @[Modules.scala 50:57:@28396.4]
  wire [10:0] _T_78338; // @[Modules.scala 50:57:@28397.4]
  wire [10:0] buffer_7_416; // @[Modules.scala 50:57:@28398.4]
  wire [11:0] _T_78352; // @[Modules.scala 50:57:@28416.4]
  wire [10:0] _T_78353; // @[Modules.scala 50:57:@28417.4]
  wire [10:0] buffer_7_421; // @[Modules.scala 50:57:@28418.4]
  wire [11:0] _T_78355; // @[Modules.scala 50:57:@28420.4]
  wire [10:0] _T_78356; // @[Modules.scala 50:57:@28421.4]
  wire [10:0] buffer_7_422; // @[Modules.scala 50:57:@28422.4]
  wire [10:0] buffer_7_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78358; // @[Modules.scala 50:57:@28424.4]
  wire [10:0] _T_78359; // @[Modules.scala 50:57:@28425.4]
  wire [10:0] buffer_7_423; // @[Modules.scala 50:57:@28426.4]
  wire [11:0] _T_78364; // @[Modules.scala 50:57:@28432.4]
  wire [10:0] _T_78365; // @[Modules.scala 50:57:@28433.4]
  wire [10:0] buffer_7_425; // @[Modules.scala 50:57:@28434.4]
  wire [11:0] _T_78373; // @[Modules.scala 50:57:@28444.4]
  wire [10:0] _T_78374; // @[Modules.scala 50:57:@28445.4]
  wire [10:0] buffer_7_428; // @[Modules.scala 50:57:@28446.4]
  wire [11:0] _T_78376; // @[Modules.scala 50:57:@28448.4]
  wire [10:0] _T_78377; // @[Modules.scala 50:57:@28449.4]
  wire [10:0] buffer_7_429; // @[Modules.scala 50:57:@28450.4]
  wire [10:0] buffer_7_76; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78379; // @[Modules.scala 50:57:@28452.4]
  wire [10:0] _T_78380; // @[Modules.scala 50:57:@28453.4]
  wire [10:0] buffer_7_430; // @[Modules.scala 50:57:@28454.4]
  wire [10:0] buffer_7_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78394; // @[Modules.scala 50:57:@28472.4]
  wire [10:0] _T_78395; // @[Modules.scala 50:57:@28473.4]
  wire [10:0] buffer_7_435; // @[Modules.scala 50:57:@28474.4]
  wire [10:0] buffer_7_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78397; // @[Modules.scala 50:57:@28476.4]
  wire [10:0] _T_78398; // @[Modules.scala 50:57:@28477.4]
  wire [10:0] buffer_7_436; // @[Modules.scala 50:57:@28478.4]
  wire [11:0] _T_78406; // @[Modules.scala 50:57:@28488.4]
  wire [10:0] _T_78407; // @[Modules.scala 50:57:@28489.4]
  wire [10:0] buffer_7_439; // @[Modules.scala 50:57:@28490.4]
  wire [10:0] buffer_7_108; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78427; // @[Modules.scala 50:57:@28516.4]
  wire [10:0] _T_78428; // @[Modules.scala 50:57:@28517.4]
  wire [10:0] buffer_7_446; // @[Modules.scala 50:57:@28518.4]
  wire [11:0] _T_78436; // @[Modules.scala 50:57:@28528.4]
  wire [10:0] _T_78437; // @[Modules.scala 50:57:@28529.4]
  wire [10:0] buffer_7_449; // @[Modules.scala 50:57:@28530.4]
  wire [10:0] buffer_7_116; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78439; // @[Modules.scala 50:57:@28532.4]
  wire [10:0] _T_78440; // @[Modules.scala 50:57:@28533.4]
  wire [10:0] buffer_7_450; // @[Modules.scala 50:57:@28534.4]
  wire [11:0] _T_78448; // @[Modules.scala 50:57:@28544.4]
  wire [10:0] _T_78449; // @[Modules.scala 50:57:@28545.4]
  wire [10:0] buffer_7_453; // @[Modules.scala 50:57:@28546.4]
  wire [11:0] _T_78466; // @[Modules.scala 50:57:@28568.4]
  wire [10:0] _T_78467; // @[Modules.scala 50:57:@28569.4]
  wire [10:0] buffer_7_459; // @[Modules.scala 50:57:@28570.4]
  wire [10:0] buffer_7_136; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78469; // @[Modules.scala 50:57:@28572.4]
  wire [10:0] _T_78470; // @[Modules.scala 50:57:@28573.4]
  wire [10:0] buffer_7_460; // @[Modules.scala 50:57:@28574.4]
  wire [10:0] buffer_7_142; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78478; // @[Modules.scala 50:57:@28584.4]
  wire [10:0] _T_78479; // @[Modules.scala 50:57:@28585.4]
  wire [10:0] buffer_7_463; // @[Modules.scala 50:57:@28586.4]
  wire [10:0] buffer_7_144; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78481; // @[Modules.scala 50:57:@28588.4]
  wire [10:0] _T_78482; // @[Modules.scala 50:57:@28589.4]
  wire [10:0] buffer_7_464; // @[Modules.scala 50:57:@28590.4]
  wire [10:0] buffer_7_146; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78484; // @[Modules.scala 50:57:@28592.4]
  wire [10:0] _T_78485; // @[Modules.scala 50:57:@28593.4]
  wire [10:0] buffer_7_465; // @[Modules.scala 50:57:@28594.4]
  wire [10:0] buffer_7_156; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78499; // @[Modules.scala 50:57:@28612.4]
  wire [10:0] _T_78500; // @[Modules.scala 50:57:@28613.4]
  wire [10:0] buffer_7_470; // @[Modules.scala 50:57:@28614.4]
  wire [11:0] _T_78502; // @[Modules.scala 50:57:@28616.4]
  wire [10:0] _T_78503; // @[Modules.scala 50:57:@28617.4]
  wire [10:0] buffer_7_471; // @[Modules.scala 50:57:@28618.4]
  wire [10:0] buffer_7_168; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78517; // @[Modules.scala 50:57:@28636.4]
  wire [10:0] _T_78518; // @[Modules.scala 50:57:@28637.4]
  wire [10:0] buffer_7_476; // @[Modules.scala 50:57:@28638.4]
  wire [11:0] _T_78532; // @[Modules.scala 50:57:@28656.4]
  wire [10:0] _T_78533; // @[Modules.scala 50:57:@28657.4]
  wire [10:0] buffer_7_481; // @[Modules.scala 50:57:@28658.4]
  wire [10:0] buffer_7_182; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78538; // @[Modules.scala 50:57:@28664.4]
  wire [10:0] _T_78539; // @[Modules.scala 50:57:@28665.4]
  wire [10:0] buffer_7_483; // @[Modules.scala 50:57:@28666.4]
  wire [10:0] buffer_7_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78550; // @[Modules.scala 50:57:@28680.4]
  wire [10:0] _T_78551; // @[Modules.scala 50:57:@28681.4]
  wire [10:0] buffer_7_487; // @[Modules.scala 50:57:@28682.4]
  wire [11:0] _T_78559; // @[Modules.scala 50:57:@28692.4]
  wire [10:0] _T_78560; // @[Modules.scala 50:57:@28693.4]
  wire [10:0] buffer_7_490; // @[Modules.scala 50:57:@28694.4]
  wire [10:0] buffer_7_198; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78562; // @[Modules.scala 50:57:@28696.4]
  wire [10:0] _T_78563; // @[Modules.scala 50:57:@28697.4]
  wire [10:0] buffer_7_491; // @[Modules.scala 50:57:@28698.4]
  wire [11:0] _T_78565; // @[Modules.scala 50:57:@28700.4]
  wire [10:0] _T_78566; // @[Modules.scala 50:57:@28701.4]
  wire [10:0] buffer_7_492; // @[Modules.scala 50:57:@28702.4]
  wire [11:0] _T_78571; // @[Modules.scala 50:57:@28708.4]
  wire [10:0] _T_78572; // @[Modules.scala 50:57:@28709.4]
  wire [10:0] buffer_7_494; // @[Modules.scala 50:57:@28710.4]
  wire [11:0] _T_78580; // @[Modules.scala 50:57:@28720.4]
  wire [10:0] _T_78581; // @[Modules.scala 50:57:@28721.4]
  wire [10:0] buffer_7_497; // @[Modules.scala 50:57:@28722.4]
  wire [11:0] _T_78583; // @[Modules.scala 50:57:@28724.4]
  wire [10:0] _T_78584; // @[Modules.scala 50:57:@28725.4]
  wire [10:0] buffer_7_498; // @[Modules.scala 50:57:@28726.4]
  wire [11:0] _T_78586; // @[Modules.scala 50:57:@28728.4]
  wire [10:0] _T_78587; // @[Modules.scala 50:57:@28729.4]
  wire [10:0] buffer_7_499; // @[Modules.scala 50:57:@28730.4]
  wire [11:0] _T_78592; // @[Modules.scala 50:57:@28736.4]
  wire [10:0] _T_78593; // @[Modules.scala 50:57:@28737.4]
  wire [10:0] buffer_7_501; // @[Modules.scala 50:57:@28738.4]
  wire [10:0] buffer_7_224; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78601; // @[Modules.scala 50:57:@28748.4]
  wire [10:0] _T_78602; // @[Modules.scala 50:57:@28749.4]
  wire [10:0] buffer_7_504; // @[Modules.scala 50:57:@28750.4]
  wire [11:0] _T_78607; // @[Modules.scala 50:57:@28756.4]
  wire [10:0] _T_78608; // @[Modules.scala 50:57:@28757.4]
  wire [10:0] buffer_7_506; // @[Modules.scala 50:57:@28758.4]
  wire [10:0] buffer_7_234; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78616; // @[Modules.scala 50:57:@28768.4]
  wire [10:0] _T_78617; // @[Modules.scala 50:57:@28769.4]
  wire [10:0] buffer_7_509; // @[Modules.scala 50:57:@28770.4]
  wire [10:0] buffer_7_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78622; // @[Modules.scala 50:57:@28776.4]
  wire [10:0] _T_78623; // @[Modules.scala 50:57:@28777.4]
  wire [10:0] buffer_7_511; // @[Modules.scala 50:57:@28778.4]
  wire [10:0] buffer_7_240; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78625; // @[Modules.scala 50:57:@28780.4]
  wire [10:0] _T_78626; // @[Modules.scala 50:57:@28781.4]
  wire [10:0] buffer_7_512; // @[Modules.scala 50:57:@28782.4]
  wire [10:0] buffer_7_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78634; // @[Modules.scala 50:57:@28792.4]
  wire [10:0] _T_78635; // @[Modules.scala 50:57:@28793.4]
  wire [10:0] buffer_7_515; // @[Modules.scala 50:57:@28794.4]
  wire [10:0] buffer_7_251; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78640; // @[Modules.scala 50:57:@28800.4]
  wire [10:0] _T_78641; // @[Modules.scala 50:57:@28801.4]
  wire [10:0] buffer_7_517; // @[Modules.scala 50:57:@28802.4]
  wire [11:0] _T_78655; // @[Modules.scala 50:57:@28820.4]
  wire [10:0] _T_78656; // @[Modules.scala 50:57:@28821.4]
  wire [10:0] buffer_7_522; // @[Modules.scala 50:57:@28822.4]
  wire [10:0] buffer_7_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78658; // @[Modules.scala 50:57:@28824.4]
  wire [10:0] _T_78659; // @[Modules.scala 50:57:@28825.4]
  wire [10:0] buffer_7_523; // @[Modules.scala 50:57:@28826.4]
  wire [10:0] buffer_7_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78667; // @[Modules.scala 50:57:@28836.4]
  wire [10:0] _T_78668; // @[Modules.scala 50:57:@28837.4]
  wire [10:0] buffer_7_526; // @[Modules.scala 50:57:@28838.4]
  wire [11:0] _T_78673; // @[Modules.scala 50:57:@28844.4]
  wire [10:0] _T_78674; // @[Modules.scala 50:57:@28845.4]
  wire [10:0] buffer_7_528; // @[Modules.scala 50:57:@28846.4]
  wire [11:0] _T_78676; // @[Modules.scala 50:57:@28848.4]
  wire [10:0] _T_78677; // @[Modules.scala 50:57:@28849.4]
  wire [10:0] buffer_7_529; // @[Modules.scala 50:57:@28850.4]
  wire [10:0] buffer_7_276; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78679; // @[Modules.scala 50:57:@28852.4]
  wire [10:0] _T_78680; // @[Modules.scala 50:57:@28853.4]
  wire [10:0] buffer_7_530; // @[Modules.scala 50:57:@28854.4]
  wire [11:0] _T_78688; // @[Modules.scala 50:57:@28864.4]
  wire [10:0] _T_78689; // @[Modules.scala 50:57:@28865.4]
  wire [10:0] buffer_7_533; // @[Modules.scala 50:57:@28866.4]
  wire [10:0] buffer_7_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78703; // @[Modules.scala 50:57:@28884.4]
  wire [10:0] _T_78704; // @[Modules.scala 50:57:@28885.4]
  wire [10:0] buffer_7_538; // @[Modules.scala 50:57:@28886.4]
  wire [11:0] _T_78706; // @[Modules.scala 50:57:@28888.4]
  wire [10:0] _T_78707; // @[Modules.scala 50:57:@28889.4]
  wire [10:0] buffer_7_539; // @[Modules.scala 50:57:@28890.4]
  wire [10:0] buffer_7_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78712; // @[Modules.scala 50:57:@28896.4]
  wire [10:0] _T_78713; // @[Modules.scala 50:57:@28897.4]
  wire [10:0] buffer_7_541; // @[Modules.scala 50:57:@28898.4]
  wire [10:0] buffer_7_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78715; // @[Modules.scala 50:57:@28900.4]
  wire [10:0] _T_78716; // @[Modules.scala 50:57:@28901.4]
  wire [10:0] buffer_7_542; // @[Modules.scala 50:57:@28902.4]
  wire [10:0] buffer_7_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78724; // @[Modules.scala 50:57:@28912.4]
  wire [10:0] _T_78725; // @[Modules.scala 50:57:@28913.4]
  wire [10:0] buffer_7_545; // @[Modules.scala 50:57:@28914.4]
  wire [11:0] _T_78727; // @[Modules.scala 50:57:@28916.4]
  wire [10:0] _T_78728; // @[Modules.scala 50:57:@28917.4]
  wire [10:0] buffer_7_546; // @[Modules.scala 50:57:@28918.4]
  wire [10:0] buffer_7_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78730; // @[Modules.scala 50:57:@28920.4]
  wire [10:0] _T_78731; // @[Modules.scala 50:57:@28921.4]
  wire [10:0] buffer_7_547; // @[Modules.scala 50:57:@28922.4]
  wire [11:0] _T_78733; // @[Modules.scala 50:57:@28924.4]
  wire [10:0] _T_78734; // @[Modules.scala 50:57:@28925.4]
  wire [10:0] buffer_7_548; // @[Modules.scala 50:57:@28926.4]
  wire [11:0] _T_78739; // @[Modules.scala 50:57:@28932.4]
  wire [10:0] _T_78740; // @[Modules.scala 50:57:@28933.4]
  wire [10:0] buffer_7_550; // @[Modules.scala 50:57:@28934.4]
  wire [11:0] _T_78748; // @[Modules.scala 50:57:@28944.4]
  wire [10:0] _T_78749; // @[Modules.scala 50:57:@28945.4]
  wire [10:0] buffer_7_553; // @[Modules.scala 50:57:@28946.4]
  wire [11:0] _T_78757; // @[Modules.scala 50:57:@28956.4]
  wire [10:0] _T_78758; // @[Modules.scala 50:57:@28957.4]
  wire [10:0] buffer_7_556; // @[Modules.scala 50:57:@28958.4]
  wire [11:0] _T_78763; // @[Modules.scala 50:57:@28964.4]
  wire [10:0] _T_78764; // @[Modules.scala 50:57:@28965.4]
  wire [10:0] buffer_7_558; // @[Modules.scala 50:57:@28966.4]
  wire [11:0] _T_78766; // @[Modules.scala 50:57:@28968.4]
  wire [10:0] _T_78767; // @[Modules.scala 50:57:@28969.4]
  wire [10:0] buffer_7_559; // @[Modules.scala 50:57:@28970.4]
  wire [11:0] _T_78769; // @[Modules.scala 50:57:@28972.4]
  wire [10:0] _T_78770; // @[Modules.scala 50:57:@28973.4]
  wire [10:0] buffer_7_560; // @[Modules.scala 50:57:@28974.4]
  wire [11:0] _T_78778; // @[Modules.scala 50:57:@28984.4]
  wire [10:0] _T_78779; // @[Modules.scala 50:57:@28985.4]
  wire [10:0] buffer_7_563; // @[Modules.scala 50:57:@28986.4]
  wire [10:0] buffer_7_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78781; // @[Modules.scala 50:57:@28988.4]
  wire [10:0] _T_78782; // @[Modules.scala 50:57:@28989.4]
  wire [10:0] buffer_7_564; // @[Modules.scala 50:57:@28990.4]
  wire [11:0] _T_78787; // @[Modules.scala 50:57:@28996.4]
  wire [10:0] _T_78788; // @[Modules.scala 50:57:@28997.4]
  wire [10:0] buffer_7_566; // @[Modules.scala 50:57:@28998.4]
  wire [11:0] _T_78790; // @[Modules.scala 50:57:@29000.4]
  wire [10:0] _T_78791; // @[Modules.scala 50:57:@29001.4]
  wire [10:0] buffer_7_567; // @[Modules.scala 50:57:@29002.4]
  wire [11:0] _T_78808; // @[Modules.scala 50:57:@29024.4]
  wire [10:0] _T_78809; // @[Modules.scala 50:57:@29025.4]
  wire [10:0] buffer_7_573; // @[Modules.scala 50:57:@29026.4]
  wire [11:0] _T_78829; // @[Modules.scala 50:57:@29052.4]
  wire [10:0] _T_78830; // @[Modules.scala 50:57:@29053.4]
  wire [10:0] buffer_7_580; // @[Modules.scala 50:57:@29054.4]
  wire [10:0] buffer_7_380; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78835; // @[Modules.scala 50:57:@29060.4]
  wire [10:0] _T_78836; // @[Modules.scala 50:57:@29061.4]
  wire [10:0] buffer_7_582; // @[Modules.scala 50:57:@29062.4]
  wire [10:0] buffer_7_390; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_78850; // @[Modules.scala 50:57:@29080.4]
  wire [10:0] _T_78851; // @[Modules.scala 50:57:@29081.4]
  wire [10:0] buffer_7_587; // @[Modules.scala 50:57:@29082.4]
  wire [11:0] _T_78853; // @[Modules.scala 53:83:@29084.4]
  wire [10:0] _T_78854; // @[Modules.scala 53:83:@29085.4]
  wire [10:0] buffer_7_588; // @[Modules.scala 53:83:@29086.4]
  wire [11:0] _T_78859; // @[Modules.scala 53:83:@29092.4]
  wire [10:0] _T_78860; // @[Modules.scala 53:83:@29093.4]
  wire [10:0] buffer_7_590; // @[Modules.scala 53:83:@29094.4]
  wire [11:0] _T_78862; // @[Modules.scala 53:83:@29096.4]
  wire [10:0] _T_78863; // @[Modules.scala 53:83:@29097.4]
  wire [10:0] buffer_7_591; // @[Modules.scala 53:83:@29098.4]
  wire [11:0] _T_78865; // @[Modules.scala 53:83:@29100.4]
  wire [10:0] _T_78866; // @[Modules.scala 53:83:@29101.4]
  wire [10:0] buffer_7_592; // @[Modules.scala 53:83:@29102.4]
  wire [11:0] _T_78868; // @[Modules.scala 53:83:@29104.4]
  wire [10:0] _T_78869; // @[Modules.scala 53:83:@29105.4]
  wire [10:0] buffer_7_593; // @[Modules.scala 53:83:@29106.4]
  wire [11:0] _T_78871; // @[Modules.scala 53:83:@29108.4]
  wire [10:0] _T_78872; // @[Modules.scala 53:83:@29109.4]
  wire [10:0] buffer_7_594; // @[Modules.scala 53:83:@29110.4]
  wire [11:0] _T_78874; // @[Modules.scala 53:83:@29112.4]
  wire [10:0] _T_78875; // @[Modules.scala 53:83:@29113.4]
  wire [10:0] buffer_7_595; // @[Modules.scala 53:83:@29114.4]
  wire [11:0] _T_78883; // @[Modules.scala 53:83:@29124.4]
  wire [10:0] _T_78884; // @[Modules.scala 53:83:@29125.4]
  wire [10:0] buffer_7_598; // @[Modules.scala 53:83:@29126.4]
  wire [11:0] _T_78886; // @[Modules.scala 53:83:@29128.4]
  wire [10:0] _T_78887; // @[Modules.scala 53:83:@29129.4]
  wire [10:0] buffer_7_599; // @[Modules.scala 53:83:@29130.4]
  wire [11:0] _T_78889; // @[Modules.scala 53:83:@29132.4]
  wire [10:0] _T_78890; // @[Modules.scala 53:83:@29133.4]
  wire [10:0] buffer_7_600; // @[Modules.scala 53:83:@29134.4]
  wire [11:0] _T_78892; // @[Modules.scala 53:83:@29136.4]
  wire [10:0] _T_78893; // @[Modules.scala 53:83:@29137.4]
  wire [10:0] buffer_7_601; // @[Modules.scala 53:83:@29138.4]
  wire [11:0] _T_78895; // @[Modules.scala 53:83:@29140.4]
  wire [10:0] _T_78896; // @[Modules.scala 53:83:@29141.4]
  wire [10:0] buffer_7_602; // @[Modules.scala 53:83:@29142.4]
  wire [11:0] _T_78898; // @[Modules.scala 53:83:@29144.4]
  wire [10:0] _T_78899; // @[Modules.scala 53:83:@29145.4]
  wire [10:0] buffer_7_603; // @[Modules.scala 53:83:@29146.4]
  wire [11:0] _T_78901; // @[Modules.scala 53:83:@29148.4]
  wire [10:0] _T_78902; // @[Modules.scala 53:83:@29149.4]
  wire [10:0] buffer_7_604; // @[Modules.scala 53:83:@29150.4]
  wire [11:0] _T_78904; // @[Modules.scala 53:83:@29152.4]
  wire [10:0] _T_78905; // @[Modules.scala 53:83:@29153.4]
  wire [10:0] buffer_7_605; // @[Modules.scala 53:83:@29154.4]
  wire [11:0] _T_78907; // @[Modules.scala 53:83:@29156.4]
  wire [10:0] _T_78908; // @[Modules.scala 53:83:@29157.4]
  wire [10:0] buffer_7_606; // @[Modules.scala 53:83:@29158.4]
  wire [11:0] _T_78910; // @[Modules.scala 53:83:@29160.4]
  wire [10:0] _T_78911; // @[Modules.scala 53:83:@29161.4]
  wire [10:0] buffer_7_607; // @[Modules.scala 53:83:@29162.4]
  wire [11:0] _T_78916; // @[Modules.scala 53:83:@29168.4]
  wire [10:0] _T_78917; // @[Modules.scala 53:83:@29169.4]
  wire [10:0] buffer_7_609; // @[Modules.scala 53:83:@29170.4]
  wire [11:0] _T_78919; // @[Modules.scala 53:83:@29172.4]
  wire [10:0] _T_78920; // @[Modules.scala 53:83:@29173.4]
  wire [10:0] buffer_7_610; // @[Modules.scala 53:83:@29174.4]
  wire [11:0] _T_78922; // @[Modules.scala 53:83:@29176.4]
  wire [10:0] _T_78923; // @[Modules.scala 53:83:@29177.4]
  wire [10:0] buffer_7_611; // @[Modules.scala 53:83:@29178.4]
  wire [11:0] _T_78925; // @[Modules.scala 53:83:@29180.4]
  wire [10:0] _T_78926; // @[Modules.scala 53:83:@29181.4]
  wire [10:0] buffer_7_612; // @[Modules.scala 53:83:@29182.4]
  wire [11:0] _T_78928; // @[Modules.scala 53:83:@29184.4]
  wire [10:0] _T_78929; // @[Modules.scala 53:83:@29185.4]
  wire [10:0] buffer_7_613; // @[Modules.scala 53:83:@29186.4]
  wire [11:0] _T_78934; // @[Modules.scala 53:83:@29192.4]
  wire [10:0] _T_78935; // @[Modules.scala 53:83:@29193.4]
  wire [10:0] buffer_7_615; // @[Modules.scala 53:83:@29194.4]
  wire [11:0] _T_78937; // @[Modules.scala 53:83:@29196.4]
  wire [10:0] _T_78938; // @[Modules.scala 53:83:@29197.4]
  wire [10:0] buffer_7_616; // @[Modules.scala 53:83:@29198.4]
  wire [11:0] _T_78940; // @[Modules.scala 53:83:@29200.4]
  wire [10:0] _T_78941; // @[Modules.scala 53:83:@29201.4]
  wire [10:0] buffer_7_617; // @[Modules.scala 53:83:@29202.4]
  wire [11:0] _T_78943; // @[Modules.scala 53:83:@29204.4]
  wire [10:0] _T_78944; // @[Modules.scala 53:83:@29205.4]
  wire [10:0] buffer_7_618; // @[Modules.scala 53:83:@29206.4]
  wire [11:0] _T_78952; // @[Modules.scala 53:83:@29216.4]
  wire [10:0] _T_78953; // @[Modules.scala 53:83:@29217.4]
  wire [10:0] buffer_7_621; // @[Modules.scala 53:83:@29218.4]
  wire [11:0] _T_78955; // @[Modules.scala 53:83:@29220.4]
  wire [10:0] _T_78956; // @[Modules.scala 53:83:@29221.4]
  wire [10:0] buffer_7_622; // @[Modules.scala 53:83:@29222.4]
  wire [11:0] _T_78958; // @[Modules.scala 53:83:@29224.4]
  wire [10:0] _T_78959; // @[Modules.scala 53:83:@29225.4]
  wire [10:0] buffer_7_623; // @[Modules.scala 53:83:@29226.4]
  wire [11:0] _T_78961; // @[Modules.scala 53:83:@29228.4]
  wire [10:0] _T_78962; // @[Modules.scala 53:83:@29229.4]
  wire [10:0] buffer_7_624; // @[Modules.scala 53:83:@29230.4]
  wire [11:0] _T_78970; // @[Modules.scala 53:83:@29240.4]
  wire [10:0] _T_78971; // @[Modules.scala 53:83:@29241.4]
  wire [10:0] buffer_7_627; // @[Modules.scala 53:83:@29242.4]
  wire [11:0] _T_78979; // @[Modules.scala 53:83:@29252.4]
  wire [10:0] _T_78980; // @[Modules.scala 53:83:@29253.4]
  wire [10:0] buffer_7_630; // @[Modules.scala 53:83:@29254.4]
  wire [11:0] _T_78985; // @[Modules.scala 53:83:@29260.4]
  wire [10:0] _T_78986; // @[Modules.scala 53:83:@29261.4]
  wire [10:0] buffer_7_632; // @[Modules.scala 53:83:@29262.4]
  wire [11:0] _T_78988; // @[Modules.scala 53:83:@29264.4]
  wire [10:0] _T_78989; // @[Modules.scala 53:83:@29265.4]
  wire [10:0] buffer_7_633; // @[Modules.scala 53:83:@29266.4]
  wire [11:0] _T_78994; // @[Modules.scala 53:83:@29272.4]
  wire [10:0] _T_78995; // @[Modules.scala 53:83:@29273.4]
  wire [10:0] buffer_7_635; // @[Modules.scala 53:83:@29274.4]
  wire [11:0] _T_79000; // @[Modules.scala 53:83:@29280.4]
  wire [10:0] _T_79001; // @[Modules.scala 53:83:@29281.4]
  wire [10:0] buffer_7_637; // @[Modules.scala 53:83:@29282.4]
  wire [11:0] _T_79003; // @[Modules.scala 53:83:@29284.4]
  wire [10:0] _T_79004; // @[Modules.scala 53:83:@29285.4]
  wire [10:0] buffer_7_638; // @[Modules.scala 53:83:@29286.4]
  wire [11:0] _T_79006; // @[Modules.scala 53:83:@29288.4]
  wire [10:0] _T_79007; // @[Modules.scala 53:83:@29289.4]
  wire [10:0] buffer_7_639; // @[Modules.scala 53:83:@29290.4]
  wire [11:0] _T_79009; // @[Modules.scala 53:83:@29292.4]
  wire [10:0] _T_79010; // @[Modules.scala 53:83:@29293.4]
  wire [10:0] buffer_7_640; // @[Modules.scala 53:83:@29294.4]
  wire [11:0] _T_79012; // @[Modules.scala 53:83:@29296.4]
  wire [10:0] _T_79013; // @[Modules.scala 53:83:@29297.4]
  wire [10:0] buffer_7_641; // @[Modules.scala 53:83:@29298.4]
  wire [11:0] _T_79015; // @[Modules.scala 53:83:@29300.4]
  wire [10:0] _T_79016; // @[Modules.scala 53:83:@29301.4]
  wire [10:0] buffer_7_642; // @[Modules.scala 53:83:@29302.4]
  wire [11:0] _T_79018; // @[Modules.scala 53:83:@29304.4]
  wire [10:0] _T_79019; // @[Modules.scala 53:83:@29305.4]
  wire [10:0] buffer_7_643; // @[Modules.scala 53:83:@29306.4]
  wire [11:0] _T_79021; // @[Modules.scala 53:83:@29308.4]
  wire [10:0] _T_79022; // @[Modules.scala 53:83:@29309.4]
  wire [10:0] buffer_7_644; // @[Modules.scala 53:83:@29310.4]
  wire [11:0] _T_79024; // @[Modules.scala 53:83:@29312.4]
  wire [10:0] _T_79025; // @[Modules.scala 53:83:@29313.4]
  wire [10:0] buffer_7_645; // @[Modules.scala 53:83:@29314.4]
  wire [11:0] _T_79027; // @[Modules.scala 53:83:@29316.4]
  wire [10:0] _T_79028; // @[Modules.scala 53:83:@29317.4]
  wire [10:0] buffer_7_646; // @[Modules.scala 53:83:@29318.4]
  wire [11:0] _T_79030; // @[Modules.scala 53:83:@29320.4]
  wire [10:0] _T_79031; // @[Modules.scala 53:83:@29321.4]
  wire [10:0] buffer_7_647; // @[Modules.scala 53:83:@29322.4]
  wire [11:0] _T_79033; // @[Modules.scala 53:83:@29324.4]
  wire [10:0] _T_79034; // @[Modules.scala 53:83:@29325.4]
  wire [10:0] buffer_7_648; // @[Modules.scala 53:83:@29326.4]
  wire [11:0] _T_79036; // @[Modules.scala 53:83:@29328.4]
  wire [10:0] _T_79037; // @[Modules.scala 53:83:@29329.4]
  wire [10:0] buffer_7_649; // @[Modules.scala 53:83:@29330.4]
  wire [11:0] _T_79039; // @[Modules.scala 53:83:@29332.4]
  wire [10:0] _T_79040; // @[Modules.scala 53:83:@29333.4]
  wire [10:0] buffer_7_650; // @[Modules.scala 53:83:@29334.4]
  wire [11:0] _T_79042; // @[Modules.scala 53:83:@29336.4]
  wire [10:0] _T_79043; // @[Modules.scala 53:83:@29337.4]
  wire [10:0] buffer_7_651; // @[Modules.scala 53:83:@29338.4]
  wire [11:0] _T_79045; // @[Modules.scala 53:83:@29340.4]
  wire [10:0] _T_79046; // @[Modules.scala 53:83:@29341.4]
  wire [10:0] buffer_7_652; // @[Modules.scala 53:83:@29342.4]
  wire [11:0] _T_79048; // @[Modules.scala 53:83:@29344.4]
  wire [10:0] _T_79049; // @[Modules.scala 53:83:@29345.4]
  wire [10:0] buffer_7_653; // @[Modules.scala 53:83:@29346.4]
  wire [11:0] _T_79051; // @[Modules.scala 53:83:@29348.4]
  wire [10:0] _T_79052; // @[Modules.scala 53:83:@29349.4]
  wire [10:0] buffer_7_654; // @[Modules.scala 53:83:@29350.4]
  wire [11:0] _T_79054; // @[Modules.scala 53:83:@29352.4]
  wire [10:0] _T_79055; // @[Modules.scala 53:83:@29353.4]
  wire [10:0] buffer_7_655; // @[Modules.scala 53:83:@29354.4]
  wire [11:0] _T_79057; // @[Modules.scala 53:83:@29356.4]
  wire [10:0] _T_79058; // @[Modules.scala 53:83:@29357.4]
  wire [10:0] buffer_7_656; // @[Modules.scala 53:83:@29358.4]
  wire [11:0] _T_79060; // @[Modules.scala 53:83:@29360.4]
  wire [10:0] _T_79061; // @[Modules.scala 53:83:@29361.4]
  wire [10:0] buffer_7_657; // @[Modules.scala 53:83:@29362.4]
  wire [11:0] _T_79063; // @[Modules.scala 53:83:@29364.4]
  wire [10:0] _T_79064; // @[Modules.scala 53:83:@29365.4]
  wire [10:0] buffer_7_658; // @[Modules.scala 53:83:@29366.4]
  wire [11:0] _T_79069; // @[Modules.scala 53:83:@29372.4]
  wire [10:0] _T_79070; // @[Modules.scala 53:83:@29373.4]
  wire [10:0] buffer_7_660; // @[Modules.scala 53:83:@29374.4]
  wire [11:0] _T_79072; // @[Modules.scala 53:83:@29376.4]
  wire [10:0] _T_79073; // @[Modules.scala 53:83:@29377.4]
  wire [10:0] buffer_7_661; // @[Modules.scala 53:83:@29378.4]
  wire [11:0] _T_79075; // @[Modules.scala 53:83:@29380.4]
  wire [10:0] _T_79076; // @[Modules.scala 53:83:@29381.4]
  wire [10:0] buffer_7_662; // @[Modules.scala 53:83:@29382.4]
  wire [11:0] _T_79078; // @[Modules.scala 53:83:@29384.4]
  wire [10:0] _T_79079; // @[Modules.scala 53:83:@29385.4]
  wire [10:0] buffer_7_663; // @[Modules.scala 53:83:@29386.4]
  wire [11:0] _T_79081; // @[Modules.scala 53:83:@29388.4]
  wire [10:0] _T_79082; // @[Modules.scala 53:83:@29389.4]
  wire [10:0] buffer_7_664; // @[Modules.scala 53:83:@29390.4]
  wire [11:0] _T_79084; // @[Modules.scala 53:83:@29392.4]
  wire [10:0] _T_79085; // @[Modules.scala 53:83:@29393.4]
  wire [10:0] buffer_7_665; // @[Modules.scala 53:83:@29394.4]
  wire [11:0] _T_79087; // @[Modules.scala 53:83:@29396.4]
  wire [10:0] _T_79088; // @[Modules.scala 53:83:@29397.4]
  wire [10:0] buffer_7_666; // @[Modules.scala 53:83:@29398.4]
  wire [11:0] _T_79090; // @[Modules.scala 53:83:@29400.4]
  wire [10:0] _T_79091; // @[Modules.scala 53:83:@29401.4]
  wire [10:0] buffer_7_667; // @[Modules.scala 53:83:@29402.4]
  wire [11:0] _T_79093; // @[Modules.scala 53:83:@29404.4]
  wire [10:0] _T_79094; // @[Modules.scala 53:83:@29405.4]
  wire [10:0] buffer_7_668; // @[Modules.scala 53:83:@29406.4]
  wire [11:0] _T_79096; // @[Modules.scala 53:83:@29408.4]
  wire [10:0] _T_79097; // @[Modules.scala 53:83:@29409.4]
  wire [10:0] buffer_7_669; // @[Modules.scala 53:83:@29410.4]
  wire [11:0] _T_79099; // @[Modules.scala 53:83:@29412.4]
  wire [10:0] _T_79100; // @[Modules.scala 53:83:@29413.4]
  wire [10:0] buffer_7_670; // @[Modules.scala 53:83:@29414.4]
  wire [11:0] _T_79102; // @[Modules.scala 53:83:@29416.4]
  wire [10:0] _T_79103; // @[Modules.scala 53:83:@29417.4]
  wire [10:0] buffer_7_671; // @[Modules.scala 53:83:@29418.4]
  wire [11:0] _T_79105; // @[Modules.scala 53:83:@29420.4]
  wire [10:0] _T_79106; // @[Modules.scala 53:83:@29421.4]
  wire [10:0] buffer_7_672; // @[Modules.scala 53:83:@29422.4]
  wire [11:0] _T_79108; // @[Modules.scala 53:83:@29424.4]
  wire [10:0] _T_79109; // @[Modules.scala 53:83:@29425.4]
  wire [10:0] buffer_7_673; // @[Modules.scala 53:83:@29426.4]
  wire [11:0] _T_79111; // @[Modules.scala 53:83:@29428.4]
  wire [10:0] _T_79112; // @[Modules.scala 53:83:@29429.4]
  wire [10:0] buffer_7_674; // @[Modules.scala 53:83:@29430.4]
  wire [11:0] _T_79114; // @[Modules.scala 53:83:@29432.4]
  wire [10:0] _T_79115; // @[Modules.scala 53:83:@29433.4]
  wire [10:0] buffer_7_675; // @[Modules.scala 53:83:@29434.4]
  wire [11:0] _T_79123; // @[Modules.scala 53:83:@29444.4]
  wire [10:0] _T_79124; // @[Modules.scala 53:83:@29445.4]
  wire [10:0] buffer_7_678; // @[Modules.scala 53:83:@29446.4]
  wire [11:0] _T_79135; // @[Modules.scala 53:83:@29460.4]
  wire [10:0] _T_79136; // @[Modules.scala 53:83:@29461.4]
  wire [10:0] buffer_7_682; // @[Modules.scala 53:83:@29462.4]
  wire [11:0] _T_79138; // @[Modules.scala 53:83:@29464.4]
  wire [10:0] _T_79139; // @[Modules.scala 53:83:@29465.4]
  wire [10:0] buffer_7_683; // @[Modules.scala 53:83:@29466.4]
  wire [11:0] _T_79144; // @[Modules.scala 53:83:@29472.4]
  wire [10:0] _T_79145; // @[Modules.scala 53:83:@29473.4]
  wire [10:0] buffer_7_685; // @[Modules.scala 53:83:@29474.4]
  wire [11:0] _T_79147; // @[Modules.scala 56:109:@29476.4]
  wire [10:0] _T_79148; // @[Modules.scala 56:109:@29477.4]
  wire [10:0] buffer_7_686; // @[Modules.scala 56:109:@29478.4]
  wire [11:0] _T_79150; // @[Modules.scala 56:109:@29480.4]
  wire [10:0] _T_79151; // @[Modules.scala 56:109:@29481.4]
  wire [10:0] buffer_7_687; // @[Modules.scala 56:109:@29482.4]
  wire [11:0] _T_79153; // @[Modules.scala 56:109:@29484.4]
  wire [10:0] _T_79154; // @[Modules.scala 56:109:@29485.4]
  wire [10:0] buffer_7_688; // @[Modules.scala 56:109:@29486.4]
  wire [11:0] _T_79156; // @[Modules.scala 56:109:@29488.4]
  wire [10:0] _T_79157; // @[Modules.scala 56:109:@29489.4]
  wire [10:0] buffer_7_689; // @[Modules.scala 56:109:@29490.4]
  wire [11:0] _T_79162; // @[Modules.scala 56:109:@29496.4]
  wire [10:0] _T_79163; // @[Modules.scala 56:109:@29497.4]
  wire [10:0] buffer_7_691; // @[Modules.scala 56:109:@29498.4]
  wire [11:0] _T_79165; // @[Modules.scala 56:109:@29500.4]
  wire [10:0] _T_79166; // @[Modules.scala 56:109:@29501.4]
  wire [10:0] buffer_7_692; // @[Modules.scala 56:109:@29502.4]
  wire [11:0] _T_79168; // @[Modules.scala 56:109:@29504.4]
  wire [10:0] _T_79169; // @[Modules.scala 56:109:@29505.4]
  wire [10:0] buffer_7_693; // @[Modules.scala 56:109:@29506.4]
  wire [11:0] _T_79171; // @[Modules.scala 56:109:@29508.4]
  wire [10:0] _T_79172; // @[Modules.scala 56:109:@29509.4]
  wire [10:0] buffer_7_694; // @[Modules.scala 56:109:@29510.4]
  wire [11:0] _T_79174; // @[Modules.scala 56:109:@29512.4]
  wire [10:0] _T_79175; // @[Modules.scala 56:109:@29513.4]
  wire [10:0] buffer_7_695; // @[Modules.scala 56:109:@29514.4]
  wire [11:0] _T_79177; // @[Modules.scala 56:109:@29516.4]
  wire [10:0] _T_79178; // @[Modules.scala 56:109:@29517.4]
  wire [10:0] buffer_7_696; // @[Modules.scala 56:109:@29518.4]
  wire [11:0] _T_79180; // @[Modules.scala 56:109:@29520.4]
  wire [10:0] _T_79181; // @[Modules.scala 56:109:@29521.4]
  wire [10:0] buffer_7_697; // @[Modules.scala 56:109:@29522.4]
  wire [11:0] _T_79183; // @[Modules.scala 56:109:@29524.4]
  wire [10:0] _T_79184; // @[Modules.scala 56:109:@29525.4]
  wire [10:0] buffer_7_698; // @[Modules.scala 56:109:@29526.4]
  wire [11:0] _T_79186; // @[Modules.scala 56:109:@29528.4]
  wire [10:0] _T_79187; // @[Modules.scala 56:109:@29529.4]
  wire [10:0] buffer_7_699; // @[Modules.scala 56:109:@29530.4]
  wire [11:0] _T_79189; // @[Modules.scala 56:109:@29532.4]
  wire [10:0] _T_79190; // @[Modules.scala 56:109:@29533.4]
  wire [10:0] buffer_7_700; // @[Modules.scala 56:109:@29534.4]
  wire [11:0] _T_79192; // @[Modules.scala 56:109:@29536.4]
  wire [10:0] _T_79193; // @[Modules.scala 56:109:@29537.4]
  wire [10:0] buffer_7_701; // @[Modules.scala 56:109:@29538.4]
  wire [11:0] _T_79195; // @[Modules.scala 56:109:@29540.4]
  wire [10:0] _T_79196; // @[Modules.scala 56:109:@29541.4]
  wire [10:0] buffer_7_702; // @[Modules.scala 56:109:@29542.4]
  wire [11:0] _T_79198; // @[Modules.scala 56:109:@29544.4]
  wire [10:0] _T_79199; // @[Modules.scala 56:109:@29545.4]
  wire [10:0] buffer_7_703; // @[Modules.scala 56:109:@29546.4]
  wire [11:0] _T_79201; // @[Modules.scala 56:109:@29548.4]
  wire [10:0] _T_79202; // @[Modules.scala 56:109:@29549.4]
  wire [10:0] buffer_7_704; // @[Modules.scala 56:109:@29550.4]
  wire [11:0] _T_79204; // @[Modules.scala 56:109:@29552.4]
  wire [10:0] _T_79205; // @[Modules.scala 56:109:@29553.4]
  wire [10:0] buffer_7_705; // @[Modules.scala 56:109:@29554.4]
  wire [11:0] _T_79207; // @[Modules.scala 56:109:@29556.4]
  wire [10:0] _T_79208; // @[Modules.scala 56:109:@29557.4]
  wire [10:0] buffer_7_706; // @[Modules.scala 56:109:@29558.4]
  wire [11:0] _T_79210; // @[Modules.scala 56:109:@29560.4]
  wire [10:0] _T_79211; // @[Modules.scala 56:109:@29561.4]
  wire [10:0] buffer_7_707; // @[Modules.scala 56:109:@29562.4]
  wire [11:0] _T_79213; // @[Modules.scala 56:109:@29564.4]
  wire [10:0] _T_79214; // @[Modules.scala 56:109:@29565.4]
  wire [10:0] buffer_7_708; // @[Modules.scala 56:109:@29566.4]
  wire [11:0] _T_79216; // @[Modules.scala 56:109:@29568.4]
  wire [10:0] _T_79217; // @[Modules.scala 56:109:@29569.4]
  wire [10:0] buffer_7_709; // @[Modules.scala 56:109:@29570.4]
  wire [11:0] _T_79219; // @[Modules.scala 56:109:@29572.4]
  wire [10:0] _T_79220; // @[Modules.scala 56:109:@29573.4]
  wire [10:0] buffer_7_710; // @[Modules.scala 56:109:@29574.4]
  wire [11:0] _T_79222; // @[Modules.scala 56:109:@29576.4]
  wire [10:0] _T_79223; // @[Modules.scala 56:109:@29577.4]
  wire [10:0] buffer_7_711; // @[Modules.scala 56:109:@29578.4]
  wire [11:0] _T_79225; // @[Modules.scala 56:109:@29580.4]
  wire [10:0] _T_79226; // @[Modules.scala 56:109:@29581.4]
  wire [10:0] buffer_7_712; // @[Modules.scala 56:109:@29582.4]
  wire [11:0] _T_79228; // @[Modules.scala 56:109:@29584.4]
  wire [10:0] _T_79229; // @[Modules.scala 56:109:@29585.4]
  wire [10:0] buffer_7_713; // @[Modules.scala 56:109:@29586.4]
  wire [11:0] _T_79231; // @[Modules.scala 56:109:@29588.4]
  wire [10:0] _T_79232; // @[Modules.scala 56:109:@29589.4]
  wire [10:0] buffer_7_714; // @[Modules.scala 56:109:@29590.4]
  wire [11:0] _T_79234; // @[Modules.scala 56:109:@29592.4]
  wire [10:0] _T_79235; // @[Modules.scala 56:109:@29593.4]
  wire [10:0] buffer_7_715; // @[Modules.scala 56:109:@29594.4]
  wire [11:0] _T_79237; // @[Modules.scala 56:109:@29596.4]
  wire [10:0] _T_79238; // @[Modules.scala 56:109:@29597.4]
  wire [10:0] buffer_7_716; // @[Modules.scala 56:109:@29598.4]
  wire [11:0] _T_79240; // @[Modules.scala 56:109:@29600.4]
  wire [10:0] _T_79241; // @[Modules.scala 56:109:@29601.4]
  wire [10:0] buffer_7_717; // @[Modules.scala 56:109:@29602.4]
  wire [11:0] _T_79243; // @[Modules.scala 56:109:@29604.4]
  wire [10:0] _T_79244; // @[Modules.scala 56:109:@29605.4]
  wire [10:0] buffer_7_718; // @[Modules.scala 56:109:@29606.4]
  wire [11:0] _T_79246; // @[Modules.scala 56:109:@29608.4]
  wire [10:0] _T_79247; // @[Modules.scala 56:109:@29609.4]
  wire [10:0] buffer_7_719; // @[Modules.scala 56:109:@29610.4]
  wire [11:0] _T_79249; // @[Modules.scala 56:109:@29612.4]
  wire [10:0] _T_79250; // @[Modules.scala 56:109:@29613.4]
  wire [10:0] buffer_7_720; // @[Modules.scala 56:109:@29614.4]
  wire [11:0] _T_79252; // @[Modules.scala 56:109:@29616.4]
  wire [10:0] _T_79253; // @[Modules.scala 56:109:@29617.4]
  wire [10:0] buffer_7_721; // @[Modules.scala 56:109:@29618.4]
  wire [11:0] _T_79255; // @[Modules.scala 56:109:@29620.4]
  wire [10:0] _T_79256; // @[Modules.scala 56:109:@29621.4]
  wire [10:0] buffer_7_722; // @[Modules.scala 56:109:@29622.4]
  wire [11:0] _T_79258; // @[Modules.scala 56:109:@29624.4]
  wire [10:0] _T_79259; // @[Modules.scala 56:109:@29625.4]
  wire [10:0] buffer_7_723; // @[Modules.scala 56:109:@29626.4]
  wire [11:0] _T_79261; // @[Modules.scala 56:109:@29628.4]
  wire [10:0] _T_79262; // @[Modules.scala 56:109:@29629.4]
  wire [10:0] buffer_7_724; // @[Modules.scala 56:109:@29630.4]
  wire [11:0] _T_79264; // @[Modules.scala 56:109:@29632.4]
  wire [10:0] _T_79265; // @[Modules.scala 56:109:@29633.4]
  wire [10:0] buffer_7_725; // @[Modules.scala 56:109:@29634.4]
  wire [11:0] _T_79267; // @[Modules.scala 56:109:@29636.4]
  wire [10:0] _T_79268; // @[Modules.scala 56:109:@29637.4]
  wire [10:0] buffer_7_726; // @[Modules.scala 56:109:@29638.4]
  wire [11:0] _T_79270; // @[Modules.scala 56:109:@29640.4]
  wire [10:0] _T_79271; // @[Modules.scala 56:109:@29641.4]
  wire [10:0] buffer_7_727; // @[Modules.scala 56:109:@29642.4]
  wire [11:0] _T_79273; // @[Modules.scala 56:109:@29644.4]
  wire [10:0] _T_79274; // @[Modules.scala 56:109:@29645.4]
  wire [10:0] buffer_7_728; // @[Modules.scala 56:109:@29646.4]
  wire [11:0] _T_79276; // @[Modules.scala 56:109:@29648.4]
  wire [10:0] _T_79277; // @[Modules.scala 56:109:@29649.4]
  wire [10:0] buffer_7_729; // @[Modules.scala 56:109:@29650.4]
  wire [11:0] _T_79282; // @[Modules.scala 56:109:@29656.4]
  wire [10:0] _T_79283; // @[Modules.scala 56:109:@29657.4]
  wire [10:0] buffer_7_731; // @[Modules.scala 56:109:@29658.4]
  wire [11:0] _T_79288; // @[Modules.scala 56:109:@29664.4]
  wire [10:0] _T_79289; // @[Modules.scala 56:109:@29665.4]
  wire [10:0] buffer_7_733; // @[Modules.scala 56:109:@29666.4]
  wire [11:0] _T_79291; // @[Modules.scala 56:109:@29668.4]
  wire [10:0] _T_79292; // @[Modules.scala 56:109:@29669.4]
  wire [10:0] buffer_7_734; // @[Modules.scala 56:109:@29670.4]
  wire [11:0] _T_79294; // @[Modules.scala 63:156:@29673.4]
  wire [10:0] _T_79295; // @[Modules.scala 63:156:@29674.4]
  wire [10:0] buffer_7_736; // @[Modules.scala 63:156:@29675.4]
  wire [11:0] _T_79297; // @[Modules.scala 63:156:@29677.4]
  wire [10:0] _T_79298; // @[Modules.scala 63:156:@29678.4]
  wire [10:0] buffer_7_737; // @[Modules.scala 63:156:@29679.4]
  wire [11:0] _T_79300; // @[Modules.scala 63:156:@29681.4]
  wire [10:0] _T_79301; // @[Modules.scala 63:156:@29682.4]
  wire [10:0] buffer_7_738; // @[Modules.scala 63:156:@29683.4]
  wire [11:0] _T_79303; // @[Modules.scala 63:156:@29685.4]
  wire [10:0] _T_79304; // @[Modules.scala 63:156:@29686.4]
  wire [10:0] buffer_7_739; // @[Modules.scala 63:156:@29687.4]
  wire [11:0] _T_79306; // @[Modules.scala 63:156:@29689.4]
  wire [10:0] _T_79307; // @[Modules.scala 63:156:@29690.4]
  wire [10:0] buffer_7_740; // @[Modules.scala 63:156:@29691.4]
  wire [11:0] _T_79309; // @[Modules.scala 63:156:@29693.4]
  wire [10:0] _T_79310; // @[Modules.scala 63:156:@29694.4]
  wire [10:0] buffer_7_741; // @[Modules.scala 63:156:@29695.4]
  wire [11:0] _T_79312; // @[Modules.scala 63:156:@29697.4]
  wire [10:0] _T_79313; // @[Modules.scala 63:156:@29698.4]
  wire [10:0] buffer_7_742; // @[Modules.scala 63:156:@29699.4]
  wire [11:0] _T_79315; // @[Modules.scala 63:156:@29701.4]
  wire [10:0] _T_79316; // @[Modules.scala 63:156:@29702.4]
  wire [10:0] buffer_7_743; // @[Modules.scala 63:156:@29703.4]
  wire [11:0] _T_79318; // @[Modules.scala 63:156:@29705.4]
  wire [10:0] _T_79319; // @[Modules.scala 63:156:@29706.4]
  wire [10:0] buffer_7_744; // @[Modules.scala 63:156:@29707.4]
  wire [11:0] _T_79321; // @[Modules.scala 63:156:@29709.4]
  wire [10:0] _T_79322; // @[Modules.scala 63:156:@29710.4]
  wire [10:0] buffer_7_745; // @[Modules.scala 63:156:@29711.4]
  wire [11:0] _T_79324; // @[Modules.scala 63:156:@29713.4]
  wire [10:0] _T_79325; // @[Modules.scala 63:156:@29714.4]
  wire [10:0] buffer_7_746; // @[Modules.scala 63:156:@29715.4]
  wire [11:0] _T_79327; // @[Modules.scala 63:156:@29717.4]
  wire [10:0] _T_79328; // @[Modules.scala 63:156:@29718.4]
  wire [10:0] buffer_7_747; // @[Modules.scala 63:156:@29719.4]
  wire [11:0] _T_79330; // @[Modules.scala 63:156:@29721.4]
  wire [10:0] _T_79331; // @[Modules.scala 63:156:@29722.4]
  wire [10:0] buffer_7_748; // @[Modules.scala 63:156:@29723.4]
  wire [11:0] _T_79333; // @[Modules.scala 63:156:@29725.4]
  wire [10:0] _T_79334; // @[Modules.scala 63:156:@29726.4]
  wire [10:0] buffer_7_749; // @[Modules.scala 63:156:@29727.4]
  wire [11:0] _T_79336; // @[Modules.scala 63:156:@29729.4]
  wire [10:0] _T_79337; // @[Modules.scala 63:156:@29730.4]
  wire [10:0] buffer_7_750; // @[Modules.scala 63:156:@29731.4]
  wire [11:0] _T_79339; // @[Modules.scala 63:156:@29733.4]
  wire [10:0] _T_79340; // @[Modules.scala 63:156:@29734.4]
  wire [10:0] buffer_7_751; // @[Modules.scala 63:156:@29735.4]
  wire [11:0] _T_79342; // @[Modules.scala 63:156:@29737.4]
  wire [10:0] _T_79343; // @[Modules.scala 63:156:@29738.4]
  wire [10:0] buffer_7_752; // @[Modules.scala 63:156:@29739.4]
  wire [11:0] _T_79345; // @[Modules.scala 63:156:@29741.4]
  wire [10:0] _T_79346; // @[Modules.scala 63:156:@29742.4]
  wire [10:0] buffer_7_753; // @[Modules.scala 63:156:@29743.4]
  wire [11:0] _T_79348; // @[Modules.scala 63:156:@29745.4]
  wire [10:0] _T_79349; // @[Modules.scala 63:156:@29746.4]
  wire [10:0] buffer_7_754; // @[Modules.scala 63:156:@29747.4]
  wire [11:0] _T_79351; // @[Modules.scala 63:156:@29749.4]
  wire [10:0] _T_79352; // @[Modules.scala 63:156:@29750.4]
  wire [10:0] buffer_7_755; // @[Modules.scala 63:156:@29751.4]
  wire [11:0] _T_79354; // @[Modules.scala 63:156:@29753.4]
  wire [10:0] _T_79355; // @[Modules.scala 63:156:@29754.4]
  wire [10:0] buffer_7_756; // @[Modules.scala 63:156:@29755.4]
  wire [11:0] _T_79357; // @[Modules.scala 63:156:@29757.4]
  wire [10:0] _T_79358; // @[Modules.scala 63:156:@29758.4]
  wire [10:0] buffer_7_757; // @[Modules.scala 63:156:@29759.4]
  wire [11:0] _T_79360; // @[Modules.scala 63:156:@29761.4]
  wire [10:0] _T_79361; // @[Modules.scala 63:156:@29762.4]
  wire [10:0] buffer_7_758; // @[Modules.scala 63:156:@29763.4]
  wire [11:0] _T_79363; // @[Modules.scala 63:156:@29765.4]
  wire [10:0] _T_79364; // @[Modules.scala 63:156:@29766.4]
  wire [10:0] buffer_7_759; // @[Modules.scala 63:156:@29767.4]
  wire [11:0] _T_79366; // @[Modules.scala 63:156:@29769.4]
  wire [10:0] _T_79367; // @[Modules.scala 63:156:@29770.4]
  wire [10:0] buffer_7_760; // @[Modules.scala 63:156:@29771.4]
  wire [11:0] _T_79369; // @[Modules.scala 63:156:@29773.4]
  wire [10:0] _T_79370; // @[Modules.scala 63:156:@29774.4]
  wire [10:0] buffer_7_761; // @[Modules.scala 63:156:@29775.4]
  wire [11:0] _T_79372; // @[Modules.scala 63:156:@29777.4]
  wire [10:0] _T_79373; // @[Modules.scala 63:156:@29778.4]
  wire [10:0] buffer_7_762; // @[Modules.scala 63:156:@29779.4]
  wire [11:0] _T_79375; // @[Modules.scala 63:156:@29781.4]
  wire [10:0] _T_79376; // @[Modules.scala 63:156:@29782.4]
  wire [10:0] buffer_7_763; // @[Modules.scala 63:156:@29783.4]
  wire [11:0] _T_79378; // @[Modules.scala 63:156:@29785.4]
  wire [10:0] _T_79379; // @[Modules.scala 63:156:@29786.4]
  wire [10:0] buffer_7_764; // @[Modules.scala 63:156:@29787.4]
  wire [11:0] _T_79381; // @[Modules.scala 63:156:@29789.4]
  wire [10:0] _T_79382; // @[Modules.scala 63:156:@29790.4]
  wire [10:0] buffer_7_765; // @[Modules.scala 63:156:@29791.4]
  wire [11:0] _T_79384; // @[Modules.scala 63:156:@29793.4]
  wire [10:0] _T_79385; // @[Modules.scala 63:156:@29794.4]
  wire [10:0] buffer_7_766; // @[Modules.scala 63:156:@29795.4]
  wire [11:0] _T_79387; // @[Modules.scala 63:156:@29797.4]
  wire [10:0] _T_79388; // @[Modules.scala 63:156:@29798.4]
  wire [10:0] buffer_7_767; // @[Modules.scala 63:156:@29799.4]
  wire [11:0] _T_79390; // @[Modules.scala 63:156:@29801.4]
  wire [10:0] _T_79391; // @[Modules.scala 63:156:@29802.4]
  wire [10:0] buffer_7_768; // @[Modules.scala 63:156:@29803.4]
  wire [11:0] _T_79393; // @[Modules.scala 63:156:@29805.4]
  wire [10:0] _T_79394; // @[Modules.scala 63:156:@29806.4]
  wire [10:0] buffer_7_769; // @[Modules.scala 63:156:@29807.4]
  wire [11:0] _T_79396; // @[Modules.scala 63:156:@29809.4]
  wire [10:0] _T_79397; // @[Modules.scala 63:156:@29810.4]
  wire [10:0] buffer_7_770; // @[Modules.scala 63:156:@29811.4]
  wire [11:0] _T_79399; // @[Modules.scala 63:156:@29813.4]
  wire [10:0] _T_79400; // @[Modules.scala 63:156:@29814.4]
  wire [10:0] buffer_7_771; // @[Modules.scala 63:156:@29815.4]
  wire [11:0] _T_79402; // @[Modules.scala 63:156:@29817.4]
  wire [10:0] _T_79403; // @[Modules.scala 63:156:@29818.4]
  wire [10:0] buffer_7_772; // @[Modules.scala 63:156:@29819.4]
  wire [11:0] _T_79405; // @[Modules.scala 63:156:@29821.4]
  wire [10:0] _T_79406; // @[Modules.scala 63:156:@29822.4]
  wire [10:0] buffer_7_773; // @[Modules.scala 63:156:@29823.4]
  wire [11:0] _T_79408; // @[Modules.scala 63:156:@29825.4]
  wire [10:0] _T_79409; // @[Modules.scala 63:156:@29826.4]
  wire [10:0] buffer_7_774; // @[Modules.scala 63:156:@29827.4]
  wire [11:0] _T_79411; // @[Modules.scala 63:156:@29829.4]
  wire [10:0] _T_79412; // @[Modules.scala 63:156:@29830.4]
  wire [10:0] buffer_7_775; // @[Modules.scala 63:156:@29831.4]
  wire [11:0] _T_79414; // @[Modules.scala 63:156:@29833.4]
  wire [10:0] _T_79415; // @[Modules.scala 63:156:@29834.4]
  wire [10:0] buffer_7_776; // @[Modules.scala 63:156:@29835.4]
  wire [11:0] _T_79417; // @[Modules.scala 63:156:@29837.4]
  wire [10:0] _T_79418; // @[Modules.scala 63:156:@29838.4]
  wire [10:0] buffer_7_777; // @[Modules.scala 63:156:@29839.4]
  wire [11:0] _T_79420; // @[Modules.scala 63:156:@29841.4]
  wire [10:0] _T_79421; // @[Modules.scala 63:156:@29842.4]
  wire [10:0] buffer_7_778; // @[Modules.scala 63:156:@29843.4]
  wire [11:0] _T_79423; // @[Modules.scala 63:156:@29845.4]
  wire [10:0] _T_79424; // @[Modules.scala 63:156:@29846.4]
  wire [10:0] buffer_7_779; // @[Modules.scala 63:156:@29847.4]
  wire [11:0] _T_79426; // @[Modules.scala 63:156:@29849.4]
  wire [10:0] _T_79427; // @[Modules.scala 63:156:@29850.4]
  wire [10:0] buffer_7_780; // @[Modules.scala 63:156:@29851.4]
  wire [11:0] _T_79429; // @[Modules.scala 63:156:@29853.4]
  wire [10:0] _T_79430; // @[Modules.scala 63:156:@29854.4]
  wire [10:0] buffer_7_781; // @[Modules.scala 63:156:@29855.4]
  wire [11:0] _T_79432; // @[Modules.scala 63:156:@29857.4]
  wire [10:0] _T_79433; // @[Modules.scala 63:156:@29858.4]
  wire [10:0] buffer_7_782; // @[Modules.scala 63:156:@29859.4]
  wire [11:0] _T_79435; // @[Modules.scala 63:156:@29861.4]
  wire [10:0] _T_79436; // @[Modules.scala 63:156:@29862.4]
  wire [10:0] buffer_7_783; // @[Modules.scala 63:156:@29863.4]
  wire [5:0] _T_79763; // @[Modules.scala 43:47:@30206.4]
  wire [4:0] _T_79764; // @[Modules.scala 43:47:@30207.4]
  wire [4:0] _T_79765; // @[Modules.scala 43:47:@30208.4]
  wire [5:0] _T_79786; // @[Modules.scala 43:47:@30232.4]
  wire [4:0] _T_79787; // @[Modules.scala 43:47:@30233.4]
  wire [4:0] _T_79788; // @[Modules.scala 43:47:@30234.4]
  wire [5:0] _T_79793; // @[Modules.scala 43:47:@30239.4]
  wire [4:0] _T_79794; // @[Modules.scala 43:47:@30240.4]
  wire [4:0] _T_79795; // @[Modules.scala 43:47:@30241.4]
  wire [5:0] _T_79800; // @[Modules.scala 43:47:@30246.4]
  wire [4:0] _T_79801; // @[Modules.scala 43:47:@30247.4]
  wire [4:0] _T_79802; // @[Modules.scala 43:47:@30248.4]
  wire [5:0] _T_79838; // @[Modules.scala 46:47:@30285.4]
  wire [4:0] _T_79839; // @[Modules.scala 46:47:@30286.4]
  wire [4:0] _T_79840; // @[Modules.scala 46:47:@30287.4]
  wire [5:0] _T_79958; // @[Modules.scala 40:46:@30424.4]
  wire [4:0] _T_79959; // @[Modules.scala 40:46:@30425.4]
  wire [4:0] _T_79960; // @[Modules.scala 40:46:@30426.4]
  wire [5:0] _T_80042; // @[Modules.scala 43:47:@30515.4]
  wire [4:0] _T_80043; // @[Modules.scala 43:47:@30516.4]
  wire [4:0] _T_80044; // @[Modules.scala 43:47:@30517.4]
  wire [5:0] _T_80051; // @[Modules.scala 40:46:@30527.4]
  wire [4:0] _T_80052; // @[Modules.scala 40:46:@30528.4]
  wire [4:0] _T_80053; // @[Modules.scala 40:46:@30529.4]
  wire [5:0] _T_80068; // @[Modules.scala 40:46:@30545.4]
  wire [4:0] _T_80069; // @[Modules.scala 40:46:@30546.4]
  wire [4:0] _T_80070; // @[Modules.scala 40:46:@30547.4]
  wire [5:0] _T_80111; // @[Modules.scala 40:46:@30593.4]
  wire [4:0] _T_80112; // @[Modules.scala 40:46:@30594.4]
  wire [4:0] _T_80113; // @[Modules.scala 40:46:@30595.4]
  wire [5:0] _T_80114; // @[Modules.scala 40:46:@30597.4]
  wire [4:0] _T_80115; // @[Modules.scala 40:46:@30598.4]
  wire [4:0] _T_80116; // @[Modules.scala 40:46:@30599.4]
  wire [5:0] _T_80181; // @[Modules.scala 40:46:@30670.4]
  wire [4:0] _T_80182; // @[Modules.scala 40:46:@30671.4]
  wire [4:0] _T_80183; // @[Modules.scala 40:46:@30672.4]
  wire [5:0] _T_80417; // @[Modules.scala 37:46:@30917.4]
  wire [4:0] _T_80418; // @[Modules.scala 37:46:@30918.4]
  wire [4:0] _T_80419; // @[Modules.scala 37:46:@30919.4]
  wire [5:0] _T_80453; // @[Modules.scala 40:46:@30958.4]
  wire [4:0] _T_80454; // @[Modules.scala 40:46:@30959.4]
  wire [4:0] _T_80455; // @[Modules.scala 40:46:@30960.4]
  wire [5:0] _T_80470; // @[Modules.scala 40:46:@30976.4]
  wire [4:0] _T_80471; // @[Modules.scala 40:46:@30977.4]
  wire [4:0] _T_80472; // @[Modules.scala 40:46:@30978.4]
  wire [5:0] _T_80497; // @[Modules.scala 37:46:@31005.4]
  wire [4:0] _T_80498; // @[Modules.scala 37:46:@31006.4]
  wire [4:0] _T_80499; // @[Modules.scala 37:46:@31007.4]
  wire [5:0] _T_80522; // @[Modules.scala 43:47:@31036.4]
  wire [4:0] _T_80523; // @[Modules.scala 43:47:@31037.4]
  wire [4:0] _T_80524; // @[Modules.scala 43:47:@31038.4]
  wire [5:0] _T_80671; // @[Modules.scala 43:47:@31209.4]
  wire [4:0] _T_80672; // @[Modules.scala 43:47:@31210.4]
  wire [4:0] _T_80673; // @[Modules.scala 43:47:@31211.4]
  wire [5:0] _T_80710; // @[Modules.scala 43:47:@31254.4]
  wire [4:0] _T_80711; // @[Modules.scala 43:47:@31255.4]
  wire [4:0] _T_80712; // @[Modules.scala 43:47:@31256.4]
  wire [5:0] _T_80740; // @[Modules.scala 43:47:@31287.4]
  wire [4:0] _T_80741; // @[Modules.scala 43:47:@31288.4]
  wire [4:0] _T_80742; // @[Modules.scala 43:47:@31289.4]
  wire [5:0] _T_80890; // @[Modules.scala 43:47:@31452.4]
  wire [4:0] _T_80891; // @[Modules.scala 43:47:@31453.4]
  wire [4:0] _T_80892; // @[Modules.scala 43:47:@31454.4]
  wire [5:0] _T_80952; // @[Modules.scala 43:47:@31523.4]
  wire [4:0] _T_80953; // @[Modules.scala 43:47:@31524.4]
  wire [4:0] _T_80954; // @[Modules.scala 43:47:@31525.4]
  wire [5:0] _T_80987; // @[Modules.scala 43:47:@31558.4]
  wire [4:0] _T_80988; // @[Modules.scala 43:47:@31559.4]
  wire [4:0] _T_80989; // @[Modules.scala 43:47:@31560.4]
  wire [5:0] _T_81023; // @[Modules.scala 43:47:@31599.4]
  wire [4:0] _T_81024; // @[Modules.scala 43:47:@31600.4]
  wire [4:0] _T_81025; // @[Modules.scala 43:47:@31601.4]
  wire [5:0] _T_81095; // @[Modules.scala 43:47:@31681.4]
  wire [4:0] _T_81096; // @[Modules.scala 43:47:@31682.4]
  wire [4:0] _T_81097; // @[Modules.scala 43:47:@31683.4]
  wire [5:0] _T_81410; // @[Modules.scala 46:47:@32003.4]
  wire [4:0] _T_81411; // @[Modules.scala 46:47:@32004.4]
  wire [4:0] _T_81412; // @[Modules.scala 46:47:@32005.4]
  wire [5:0] _T_81427; // @[Modules.scala 43:47:@32021.4]
  wire [4:0] _T_81428; // @[Modules.scala 43:47:@32022.4]
  wire [4:0] _T_81429; // @[Modules.scala 43:47:@32023.4]
  wire [5:0] _T_81440; // @[Modules.scala 40:46:@32036.4]
  wire [4:0] _T_81441; // @[Modules.scala 40:46:@32037.4]
  wire [4:0] _T_81442; // @[Modules.scala 40:46:@32038.4]
  wire [11:0] _T_81504; // @[Modules.scala 50:57:@32105.4]
  wire [10:0] _T_81505; // @[Modules.scala 50:57:@32106.4]
  wire [10:0] buffer_8_394; // @[Modules.scala 50:57:@32107.4]
  wire [11:0] _T_81513; // @[Modules.scala 50:57:@32117.4]
  wire [10:0] _T_81514; // @[Modules.scala 50:57:@32118.4]
  wire [10:0] buffer_8_397; // @[Modules.scala 50:57:@32119.4]
  wire [11:0] _T_81519; // @[Modules.scala 50:57:@32125.4]
  wire [10:0] _T_81520; // @[Modules.scala 50:57:@32126.4]
  wire [10:0] buffer_8_399; // @[Modules.scala 50:57:@32127.4]
  wire [11:0] _T_81522; // @[Modules.scala 50:57:@32129.4]
  wire [10:0] _T_81523; // @[Modules.scala 50:57:@32130.4]
  wire [10:0] buffer_8_400; // @[Modules.scala 50:57:@32131.4]
  wire [11:0] _T_81564; // @[Modules.scala 50:57:@32185.4]
  wire [10:0] _T_81565; // @[Modules.scala 50:57:@32186.4]
  wire [10:0] buffer_8_414; // @[Modules.scala 50:57:@32187.4]
  wire [10:0] buffer_8_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81579; // @[Modules.scala 50:57:@32205.4]
  wire [10:0] _T_81580; // @[Modules.scala 50:57:@32206.4]
  wire [10:0] buffer_8_419; // @[Modules.scala 50:57:@32207.4]
  wire [11:0] _T_81582; // @[Modules.scala 50:57:@32209.4]
  wire [10:0] _T_81583; // @[Modules.scala 50:57:@32210.4]
  wire [10:0] buffer_8_420; // @[Modules.scala 50:57:@32211.4]
  wire [10:0] buffer_8_60; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_8_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81588; // @[Modules.scala 50:57:@32217.4]
  wire [10:0] _T_81589; // @[Modules.scala 50:57:@32218.4]
  wire [10:0] buffer_8_422; // @[Modules.scala 50:57:@32219.4]
  wire [10:0] buffer_8_62; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81591; // @[Modules.scala 50:57:@32221.4]
  wire [10:0] _T_81592; // @[Modules.scala 50:57:@32222.4]
  wire [10:0] buffer_8_423; // @[Modules.scala 50:57:@32223.4]
  wire [10:0] buffer_8_68; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81600; // @[Modules.scala 50:57:@32233.4]
  wire [10:0] _T_81601; // @[Modules.scala 50:57:@32234.4]
  wire [10:0] buffer_8_426; // @[Modules.scala 50:57:@32235.4]
  wire [11:0] _T_81603; // @[Modules.scala 50:57:@32237.4]
  wire [10:0] _T_81604; // @[Modules.scala 50:57:@32238.4]
  wire [10:0] buffer_8_427; // @[Modules.scala 50:57:@32239.4]
  wire [11:0] _T_81621; // @[Modules.scala 50:57:@32261.4]
  wire [10:0] _T_81622; // @[Modules.scala 50:57:@32262.4]
  wire [10:0] buffer_8_433; // @[Modules.scala 50:57:@32263.4]
  wire [10:0] buffer_8_96; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81642; // @[Modules.scala 50:57:@32289.4]
  wire [10:0] _T_81643; // @[Modules.scala 50:57:@32290.4]
  wire [10:0] buffer_8_440; // @[Modules.scala 50:57:@32291.4]
  wire [11:0] _T_81651; // @[Modules.scala 50:57:@32301.4]
  wire [10:0] _T_81652; // @[Modules.scala 50:57:@32302.4]
  wire [10:0] buffer_8_443; // @[Modules.scala 50:57:@32303.4]
  wire [11:0] _T_81657; // @[Modules.scala 50:57:@32309.4]
  wire [10:0] _T_81658; // @[Modules.scala 50:57:@32310.4]
  wire [10:0] buffer_8_445; // @[Modules.scala 50:57:@32311.4]
  wire [10:0] buffer_8_112; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81666; // @[Modules.scala 50:57:@32321.4]
  wire [10:0] _T_81667; // @[Modules.scala 50:57:@32322.4]
  wire [10:0] buffer_8_448; // @[Modules.scala 50:57:@32323.4]
  wire [10:0] buffer_8_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81669; // @[Modules.scala 50:57:@32325.4]
  wire [10:0] _T_81670; // @[Modules.scala 50:57:@32326.4]
  wire [10:0] buffer_8_449; // @[Modules.scala 50:57:@32327.4]
  wire [10:0] buffer_8_118; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81675; // @[Modules.scala 50:57:@32333.4]
  wire [10:0] _T_81676; // @[Modules.scala 50:57:@32334.4]
  wire [10:0] buffer_8_451; // @[Modules.scala 50:57:@32335.4]
  wire [11:0] _T_81678; // @[Modules.scala 50:57:@32337.4]
  wire [10:0] _T_81679; // @[Modules.scala 50:57:@32338.4]
  wire [10:0] buffer_8_452; // @[Modules.scala 50:57:@32339.4]
  wire [11:0] _T_81681; // @[Modules.scala 50:57:@32341.4]
  wire [10:0] _T_81682; // @[Modules.scala 50:57:@32342.4]
  wire [10:0] buffer_8_453; // @[Modules.scala 50:57:@32343.4]
  wire [10:0] buffer_8_127; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81687; // @[Modules.scala 50:57:@32349.4]
  wire [10:0] _T_81688; // @[Modules.scala 50:57:@32350.4]
  wire [10:0] buffer_8_455; // @[Modules.scala 50:57:@32351.4]
  wire [10:0] buffer_8_128; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81690; // @[Modules.scala 50:57:@32353.4]
  wire [10:0] _T_81691; // @[Modules.scala 50:57:@32354.4]
  wire [10:0] buffer_8_456; // @[Modules.scala 50:57:@32355.4]
  wire [11:0] _T_81693; // @[Modules.scala 50:57:@32357.4]
  wire [10:0] _T_81694; // @[Modules.scala 50:57:@32358.4]
  wire [10:0] buffer_8_457; // @[Modules.scala 50:57:@32359.4]
  wire [11:0] _T_81702; // @[Modules.scala 50:57:@32369.4]
  wire [10:0] _T_81703; // @[Modules.scala 50:57:@32370.4]
  wire [10:0] buffer_8_460; // @[Modules.scala 50:57:@32371.4]
  wire [10:0] buffer_8_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81708; // @[Modules.scala 50:57:@32377.4]
  wire [10:0] _T_81709; // @[Modules.scala 50:57:@32378.4]
  wire [10:0] buffer_8_462; // @[Modules.scala 50:57:@32379.4]
  wire [11:0] _T_81729; // @[Modules.scala 50:57:@32405.4]
  wire [10:0] _T_81730; // @[Modules.scala 50:57:@32406.4]
  wire [10:0] buffer_8_469; // @[Modules.scala 50:57:@32407.4]
  wire [11:0] _T_81741; // @[Modules.scala 50:57:@32421.4]
  wire [10:0] _T_81742; // @[Modules.scala 50:57:@32422.4]
  wire [10:0] buffer_8_473; // @[Modules.scala 50:57:@32423.4]
  wire [11:0] _T_81750; // @[Modules.scala 50:57:@32433.4]
  wire [10:0] _T_81751; // @[Modules.scala 50:57:@32434.4]
  wire [10:0] buffer_8_476; // @[Modules.scala 50:57:@32435.4]
  wire [11:0] _T_81762; // @[Modules.scala 50:57:@32449.4]
  wire [10:0] _T_81763; // @[Modules.scala 50:57:@32450.4]
  wire [10:0] buffer_8_480; // @[Modules.scala 50:57:@32451.4]
  wire [10:0] buffer_8_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81768; // @[Modules.scala 50:57:@32457.4]
  wire [10:0] _T_81769; // @[Modules.scala 50:57:@32458.4]
  wire [10:0] buffer_8_482; // @[Modules.scala 50:57:@32459.4]
  wire [10:0] buffer_8_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81780; // @[Modules.scala 50:57:@32473.4]
  wire [10:0] _T_81781; // @[Modules.scala 50:57:@32474.4]
  wire [10:0] buffer_8_486; // @[Modules.scala 50:57:@32475.4]
  wire [10:0] buffer_8_192; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81786; // @[Modules.scala 50:57:@32481.4]
  wire [10:0] _T_81787; // @[Modules.scala 50:57:@32482.4]
  wire [10:0] buffer_8_488; // @[Modules.scala 50:57:@32483.4]
  wire [10:0] buffer_8_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81792; // @[Modules.scala 50:57:@32489.4]
  wire [10:0] _T_81793; // @[Modules.scala 50:57:@32490.4]
  wire [10:0] buffer_8_490; // @[Modules.scala 50:57:@32491.4]
  wire [11:0] _T_81798; // @[Modules.scala 50:57:@32497.4]
  wire [10:0] _T_81799; // @[Modules.scala 50:57:@32498.4]
  wire [10:0] buffer_8_492; // @[Modules.scala 50:57:@32499.4]
  wire [10:0] buffer_8_204; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81804; // @[Modules.scala 50:57:@32505.4]
  wire [10:0] _T_81805; // @[Modules.scala 50:57:@32506.4]
  wire [10:0] buffer_8_494; // @[Modules.scala 50:57:@32507.4]
  wire [11:0] _T_81807; // @[Modules.scala 50:57:@32509.4]
  wire [10:0] _T_81808; // @[Modules.scala 50:57:@32510.4]
  wire [10:0] buffer_8_495; // @[Modules.scala 50:57:@32511.4]
  wire [11:0] _T_81828; // @[Modules.scala 50:57:@32537.4]
  wire [10:0] _T_81829; // @[Modules.scala 50:57:@32538.4]
  wire [10:0] buffer_8_502; // @[Modules.scala 50:57:@32539.4]
  wire [11:0] _T_81831; // @[Modules.scala 50:57:@32541.4]
  wire [10:0] _T_81832; // @[Modules.scala 50:57:@32542.4]
  wire [10:0] buffer_8_503; // @[Modules.scala 50:57:@32543.4]
  wire [11:0] _T_81834; // @[Modules.scala 50:57:@32545.4]
  wire [10:0] _T_81835; // @[Modules.scala 50:57:@32546.4]
  wire [10:0] buffer_8_504; // @[Modules.scala 50:57:@32547.4]
  wire [10:0] buffer_8_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81855; // @[Modules.scala 50:57:@32573.4]
  wire [10:0] _T_81856; // @[Modules.scala 50:57:@32574.4]
  wire [10:0] buffer_8_511; // @[Modules.scala 50:57:@32575.4]
  wire [11:0] _T_81867; // @[Modules.scala 50:57:@32589.4]
  wire [10:0] _T_81868; // @[Modules.scala 50:57:@32590.4]
  wire [10:0] buffer_8_515; // @[Modules.scala 50:57:@32591.4]
  wire [10:0] buffer_8_248; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81870; // @[Modules.scala 50:57:@32593.4]
  wire [10:0] _T_81871; // @[Modules.scala 50:57:@32594.4]
  wire [10:0] buffer_8_516; // @[Modules.scala 50:57:@32595.4]
  wire [11:0] _T_81876; // @[Modules.scala 50:57:@32601.4]
  wire [10:0] _T_81877; // @[Modules.scala 50:57:@32602.4]
  wire [10:0] buffer_8_518; // @[Modules.scala 50:57:@32603.4]
  wire [10:0] buffer_8_254; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81879; // @[Modules.scala 50:57:@32605.4]
  wire [10:0] _T_81880; // @[Modules.scala 50:57:@32606.4]
  wire [10:0] buffer_8_519; // @[Modules.scala 50:57:@32607.4]
  wire [11:0] _T_81897; // @[Modules.scala 50:57:@32629.4]
  wire [10:0] _T_81898; // @[Modules.scala 50:57:@32630.4]
  wire [10:0] buffer_8_525; // @[Modules.scala 50:57:@32631.4]
  wire [11:0] _T_81900; // @[Modules.scala 50:57:@32633.4]
  wire [10:0] _T_81901; // @[Modules.scala 50:57:@32634.4]
  wire [10:0] buffer_8_526; // @[Modules.scala 50:57:@32635.4]
  wire [11:0] _T_81906; // @[Modules.scala 50:57:@32641.4]
  wire [10:0] _T_81907; // @[Modules.scala 50:57:@32642.4]
  wire [10:0] buffer_8_528; // @[Modules.scala 50:57:@32643.4]
  wire [11:0] _T_81912; // @[Modules.scala 50:57:@32649.4]
  wire [10:0] _T_81913; // @[Modules.scala 50:57:@32650.4]
  wire [10:0] buffer_8_530; // @[Modules.scala 50:57:@32651.4]
  wire [11:0] _T_81918; // @[Modules.scala 50:57:@32657.4]
  wire [10:0] _T_81919; // @[Modules.scala 50:57:@32658.4]
  wire [10:0] buffer_8_532; // @[Modules.scala 50:57:@32659.4]
  wire [11:0] _T_81921; // @[Modules.scala 50:57:@32661.4]
  wire [10:0] _T_81922; // @[Modules.scala 50:57:@32662.4]
  wire [10:0] buffer_8_533; // @[Modules.scala 50:57:@32663.4]
  wire [10:0] buffer_8_284; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81924; // @[Modules.scala 50:57:@32665.4]
  wire [10:0] _T_81925; // @[Modules.scala 50:57:@32666.4]
  wire [10:0] buffer_8_534; // @[Modules.scala 50:57:@32667.4]
  wire [11:0] _T_81936; // @[Modules.scala 50:57:@32681.4]
  wire [10:0] _T_81937; // @[Modules.scala 50:57:@32682.4]
  wire [10:0] buffer_8_538; // @[Modules.scala 50:57:@32683.4]
  wire [10:0] buffer_8_298; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81945; // @[Modules.scala 50:57:@32693.4]
  wire [10:0] _T_81946; // @[Modules.scala 50:57:@32694.4]
  wire [10:0] buffer_8_541; // @[Modules.scala 50:57:@32695.4]
  wire [11:0] _T_81948; // @[Modules.scala 50:57:@32697.4]
  wire [10:0] _T_81949; // @[Modules.scala 50:57:@32698.4]
  wire [10:0] buffer_8_542; // @[Modules.scala 50:57:@32699.4]
  wire [10:0] buffer_8_303; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81951; // @[Modules.scala 50:57:@32701.4]
  wire [10:0] _T_81952; // @[Modules.scala 50:57:@32702.4]
  wire [10:0] buffer_8_543; // @[Modules.scala 50:57:@32703.4]
  wire [10:0] buffer_8_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81963; // @[Modules.scala 50:57:@32717.4]
  wire [10:0] _T_81964; // @[Modules.scala 50:57:@32718.4]
  wire [10:0] buffer_8_547; // @[Modules.scala 50:57:@32719.4]
  wire [11:0] _T_81966; // @[Modules.scala 50:57:@32721.4]
  wire [10:0] _T_81967; // @[Modules.scala 50:57:@32722.4]
  wire [10:0] buffer_8_548; // @[Modules.scala 50:57:@32723.4]
  wire [11:0] _T_81969; // @[Modules.scala 50:57:@32725.4]
  wire [10:0] _T_81970; // @[Modules.scala 50:57:@32726.4]
  wire [10:0] buffer_8_549; // @[Modules.scala 50:57:@32727.4]
  wire [11:0] _T_81984; // @[Modules.scala 50:57:@32745.4]
  wire [10:0] _T_81985; // @[Modules.scala 50:57:@32746.4]
  wire [10:0] buffer_8_554; // @[Modules.scala 50:57:@32747.4]
  wire [10:0] buffer_8_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81987; // @[Modules.scala 50:57:@32749.4]
  wire [10:0] _T_81988; // @[Modules.scala 50:57:@32750.4]
  wire [10:0] buffer_8_555; // @[Modules.scala 50:57:@32751.4]
  wire [11:0] _T_81993; // @[Modules.scala 50:57:@32757.4]
  wire [10:0] _T_81994; // @[Modules.scala 50:57:@32758.4]
  wire [10:0] buffer_8_557; // @[Modules.scala 50:57:@32759.4]
  wire [11:0] _T_81999; // @[Modules.scala 50:57:@32765.4]
  wire [10:0] _T_82000; // @[Modules.scala 50:57:@32766.4]
  wire [10:0] buffer_8_559; // @[Modules.scala 50:57:@32767.4]
  wire [11:0] _T_82005; // @[Modules.scala 50:57:@32773.4]
  wire [10:0] _T_82006; // @[Modules.scala 50:57:@32774.4]
  wire [10:0] buffer_8_561; // @[Modules.scala 50:57:@32775.4]
  wire [11:0] _T_82023; // @[Modules.scala 50:57:@32797.4]
  wire [10:0] _T_82024; // @[Modules.scala 50:57:@32798.4]
  wire [10:0] buffer_8_567; // @[Modules.scala 50:57:@32799.4]
  wire [10:0] buffer_8_376; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_82062; // @[Modules.scala 50:57:@32849.4]
  wire [10:0] _T_82063; // @[Modules.scala 50:57:@32850.4]
  wire [10:0] buffer_8_580; // @[Modules.scala 50:57:@32851.4]
  wire [10:0] buffer_8_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_82065; // @[Modules.scala 50:57:@32853.4]
  wire [10:0] _T_82066; // @[Modules.scala 50:57:@32854.4]
  wire [10:0] buffer_8_581; // @[Modules.scala 50:57:@32855.4]
  wire [10:0] buffer_8_382; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_82071; // @[Modules.scala 50:57:@32861.4]
  wire [10:0] _T_82072; // @[Modules.scala 50:57:@32862.4]
  wire [10:0] buffer_8_583; // @[Modules.scala 50:57:@32863.4]
  wire [11:0] _T_82080; // @[Modules.scala 50:57:@32873.4]
  wire [10:0] _T_82081; // @[Modules.scala 50:57:@32874.4]
  wire [10:0] buffer_8_586; // @[Modules.scala 50:57:@32875.4]
  wire [11:0] _T_82089; // @[Modules.scala 53:83:@32885.4]
  wire [10:0] _T_82090; // @[Modules.scala 53:83:@32886.4]
  wire [10:0] buffer_8_589; // @[Modules.scala 53:83:@32887.4]
  wire [11:0] _T_82092; // @[Modules.scala 53:83:@32889.4]
  wire [10:0] _T_82093; // @[Modules.scala 53:83:@32890.4]
  wire [10:0] buffer_8_590; // @[Modules.scala 53:83:@32891.4]
  wire [11:0] _T_82095; // @[Modules.scala 53:83:@32893.4]
  wire [10:0] _T_82096; // @[Modules.scala 53:83:@32894.4]
  wire [10:0] buffer_8_591; // @[Modules.scala 53:83:@32895.4]
  wire [11:0] _T_82098; // @[Modules.scala 53:83:@32897.4]
  wire [10:0] _T_82099; // @[Modules.scala 53:83:@32898.4]
  wire [10:0] buffer_8_592; // @[Modules.scala 53:83:@32899.4]
  wire [11:0] _T_82104; // @[Modules.scala 53:83:@32905.4]
  wire [10:0] _T_82105; // @[Modules.scala 53:83:@32906.4]
  wire [10:0] buffer_8_594; // @[Modules.scala 53:83:@32907.4]
  wire [11:0] _T_82116; // @[Modules.scala 53:83:@32921.4]
  wire [10:0] _T_82117; // @[Modules.scala 53:83:@32922.4]
  wire [10:0] buffer_8_598; // @[Modules.scala 53:83:@32923.4]
  wire [11:0] _T_82119; // @[Modules.scala 53:83:@32925.4]
  wire [10:0] _T_82120; // @[Modules.scala 53:83:@32926.4]
  wire [10:0] buffer_8_599; // @[Modules.scala 53:83:@32927.4]
  wire [11:0] _T_82125; // @[Modules.scala 53:83:@32933.4]
  wire [10:0] _T_82126; // @[Modules.scala 53:83:@32934.4]
  wire [10:0] buffer_8_601; // @[Modules.scala 53:83:@32935.4]
  wire [11:0] _T_82128; // @[Modules.scala 53:83:@32937.4]
  wire [10:0] _T_82129; // @[Modules.scala 53:83:@32938.4]
  wire [10:0] buffer_8_602; // @[Modules.scala 53:83:@32939.4]
  wire [11:0] _T_82131; // @[Modules.scala 53:83:@32941.4]
  wire [10:0] _T_82132; // @[Modules.scala 53:83:@32942.4]
  wire [10:0] buffer_8_603; // @[Modules.scala 53:83:@32943.4]
  wire [11:0] _T_82134; // @[Modules.scala 53:83:@32945.4]
  wire [10:0] _T_82135; // @[Modules.scala 53:83:@32946.4]
  wire [10:0] buffer_8_604; // @[Modules.scala 53:83:@32947.4]
  wire [11:0] _T_82137; // @[Modules.scala 53:83:@32949.4]
  wire [10:0] _T_82138; // @[Modules.scala 53:83:@32950.4]
  wire [10:0] buffer_8_605; // @[Modules.scala 53:83:@32951.4]
  wire [11:0] _T_82146; // @[Modules.scala 53:83:@32961.4]
  wire [10:0] _T_82147; // @[Modules.scala 53:83:@32962.4]
  wire [10:0] buffer_8_608; // @[Modules.scala 53:83:@32963.4]
  wire [11:0] _T_82152; // @[Modules.scala 53:83:@32969.4]
  wire [10:0] _T_82153; // @[Modules.scala 53:83:@32970.4]
  wire [10:0] buffer_8_610; // @[Modules.scala 53:83:@32971.4]
  wire [11:0] _T_82155; // @[Modules.scala 53:83:@32973.4]
  wire [10:0] _T_82156; // @[Modules.scala 53:83:@32974.4]
  wire [10:0] buffer_8_611; // @[Modules.scala 53:83:@32975.4]
  wire [11:0] _T_82158; // @[Modules.scala 53:83:@32977.4]
  wire [10:0] _T_82159; // @[Modules.scala 53:83:@32978.4]
  wire [10:0] buffer_8_612; // @[Modules.scala 53:83:@32979.4]
  wire [11:0] _T_82161; // @[Modules.scala 53:83:@32981.4]
  wire [10:0] _T_82162; // @[Modules.scala 53:83:@32982.4]
  wire [10:0] buffer_8_613; // @[Modules.scala 53:83:@32983.4]
  wire [11:0] _T_82164; // @[Modules.scala 53:83:@32985.4]
  wire [10:0] _T_82165; // @[Modules.scala 53:83:@32986.4]
  wire [10:0] buffer_8_614; // @[Modules.scala 53:83:@32987.4]
  wire [11:0] _T_82167; // @[Modules.scala 53:83:@32989.4]
  wire [10:0] _T_82168; // @[Modules.scala 53:83:@32990.4]
  wire [10:0] buffer_8_615; // @[Modules.scala 53:83:@32991.4]
  wire [11:0] _T_82170; // @[Modules.scala 53:83:@32993.4]
  wire [10:0] _T_82171; // @[Modules.scala 53:83:@32994.4]
  wire [10:0] buffer_8_616; // @[Modules.scala 53:83:@32995.4]
  wire [11:0] _T_82173; // @[Modules.scala 53:83:@32997.4]
  wire [10:0] _T_82174; // @[Modules.scala 53:83:@32998.4]
  wire [10:0] buffer_8_617; // @[Modules.scala 53:83:@32999.4]
  wire [11:0] _T_82176; // @[Modules.scala 53:83:@33001.4]
  wire [10:0] _T_82177; // @[Modules.scala 53:83:@33002.4]
  wire [10:0] buffer_8_618; // @[Modules.scala 53:83:@33003.4]
  wire [11:0] _T_82179; // @[Modules.scala 53:83:@33005.4]
  wire [10:0] _T_82180; // @[Modules.scala 53:83:@33006.4]
  wire [10:0] buffer_8_619; // @[Modules.scala 53:83:@33007.4]
  wire [11:0] _T_82182; // @[Modules.scala 53:83:@33009.4]
  wire [10:0] _T_82183; // @[Modules.scala 53:83:@33010.4]
  wire [10:0] buffer_8_620; // @[Modules.scala 53:83:@33011.4]
  wire [11:0] _T_82185; // @[Modules.scala 53:83:@33013.4]
  wire [10:0] _T_82186; // @[Modules.scala 53:83:@33014.4]
  wire [10:0] buffer_8_621; // @[Modules.scala 53:83:@33015.4]
  wire [11:0] _T_82188; // @[Modules.scala 53:83:@33017.4]
  wire [10:0] _T_82189; // @[Modules.scala 53:83:@33018.4]
  wire [10:0] buffer_8_622; // @[Modules.scala 53:83:@33019.4]
  wire [11:0] _T_82191; // @[Modules.scala 53:83:@33021.4]
  wire [10:0] _T_82192; // @[Modules.scala 53:83:@33022.4]
  wire [10:0] buffer_8_623; // @[Modules.scala 53:83:@33023.4]
  wire [11:0] _T_82197; // @[Modules.scala 53:83:@33029.4]
  wire [10:0] _T_82198; // @[Modules.scala 53:83:@33030.4]
  wire [10:0] buffer_8_625; // @[Modules.scala 53:83:@33031.4]
  wire [11:0] _T_82200; // @[Modules.scala 53:83:@33033.4]
  wire [10:0] _T_82201; // @[Modules.scala 53:83:@33034.4]
  wire [10:0] buffer_8_626; // @[Modules.scala 53:83:@33035.4]
  wire [11:0] _T_82206; // @[Modules.scala 53:83:@33041.4]
  wire [10:0] _T_82207; // @[Modules.scala 53:83:@33042.4]
  wire [10:0] buffer_8_628; // @[Modules.scala 53:83:@33043.4]
  wire [11:0] _T_82209; // @[Modules.scala 53:83:@33045.4]
  wire [10:0] _T_82210; // @[Modules.scala 53:83:@33046.4]
  wire [10:0] buffer_8_629; // @[Modules.scala 53:83:@33047.4]
  wire [11:0] _T_82212; // @[Modules.scala 53:83:@33049.4]
  wire [10:0] _T_82213; // @[Modules.scala 53:83:@33050.4]
  wire [10:0] buffer_8_630; // @[Modules.scala 53:83:@33051.4]
  wire [11:0] _T_82218; // @[Modules.scala 53:83:@33057.4]
  wire [10:0] _T_82219; // @[Modules.scala 53:83:@33058.4]
  wire [10:0] buffer_8_632; // @[Modules.scala 53:83:@33059.4]
  wire [11:0] _T_82221; // @[Modules.scala 53:83:@33061.4]
  wire [10:0] _T_82222; // @[Modules.scala 53:83:@33062.4]
  wire [10:0] buffer_8_633; // @[Modules.scala 53:83:@33063.4]
  wire [11:0] _T_82224; // @[Modules.scala 53:83:@33065.4]
  wire [10:0] _T_82225; // @[Modules.scala 53:83:@33066.4]
  wire [10:0] buffer_8_634; // @[Modules.scala 53:83:@33067.4]
  wire [11:0] _T_82227; // @[Modules.scala 53:83:@33069.4]
  wire [10:0] _T_82228; // @[Modules.scala 53:83:@33070.4]
  wire [10:0] buffer_8_635; // @[Modules.scala 53:83:@33071.4]
  wire [11:0] _T_82230; // @[Modules.scala 53:83:@33073.4]
  wire [10:0] _T_82231; // @[Modules.scala 53:83:@33074.4]
  wire [10:0] buffer_8_636; // @[Modules.scala 53:83:@33075.4]
  wire [11:0] _T_82233; // @[Modules.scala 53:83:@33077.4]
  wire [10:0] _T_82234; // @[Modules.scala 53:83:@33078.4]
  wire [10:0] buffer_8_637; // @[Modules.scala 53:83:@33079.4]
  wire [11:0] _T_82236; // @[Modules.scala 53:83:@33081.4]
  wire [10:0] _T_82237; // @[Modules.scala 53:83:@33082.4]
  wire [10:0] buffer_8_638; // @[Modules.scala 53:83:@33083.4]
  wire [11:0] _T_82239; // @[Modules.scala 53:83:@33085.4]
  wire [10:0] _T_82240; // @[Modules.scala 53:83:@33086.4]
  wire [10:0] buffer_8_639; // @[Modules.scala 53:83:@33087.4]
  wire [11:0] _T_82245; // @[Modules.scala 53:83:@33093.4]
  wire [10:0] _T_82246; // @[Modules.scala 53:83:@33094.4]
  wire [10:0] buffer_8_641; // @[Modules.scala 53:83:@33095.4]
  wire [11:0] _T_82248; // @[Modules.scala 53:83:@33097.4]
  wire [10:0] _T_82249; // @[Modules.scala 53:83:@33098.4]
  wire [10:0] buffer_8_642; // @[Modules.scala 53:83:@33099.4]
  wire [11:0] _T_82251; // @[Modules.scala 53:83:@33101.4]
  wire [10:0] _T_82252; // @[Modules.scala 53:83:@33102.4]
  wire [10:0] buffer_8_643; // @[Modules.scala 53:83:@33103.4]
  wire [11:0] _T_82254; // @[Modules.scala 53:83:@33105.4]
  wire [10:0] _T_82255; // @[Modules.scala 53:83:@33106.4]
  wire [10:0] buffer_8_644; // @[Modules.scala 53:83:@33107.4]
  wire [11:0] _T_82260; // @[Modules.scala 53:83:@33113.4]
  wire [10:0] _T_82261; // @[Modules.scala 53:83:@33114.4]
  wire [10:0] buffer_8_646; // @[Modules.scala 53:83:@33115.4]
  wire [11:0] _T_82263; // @[Modules.scala 53:83:@33117.4]
  wire [10:0] _T_82264; // @[Modules.scala 53:83:@33118.4]
  wire [10:0] buffer_8_647; // @[Modules.scala 53:83:@33119.4]
  wire [11:0] _T_82266; // @[Modules.scala 53:83:@33121.4]
  wire [10:0] _T_82267; // @[Modules.scala 53:83:@33122.4]
  wire [10:0] buffer_8_648; // @[Modules.scala 53:83:@33123.4]
  wire [11:0] _T_82269; // @[Modules.scala 53:83:@33125.4]
  wire [10:0] _T_82270; // @[Modules.scala 53:83:@33126.4]
  wire [10:0] buffer_8_649; // @[Modules.scala 53:83:@33127.4]
  wire [11:0] _T_82272; // @[Modules.scala 53:83:@33129.4]
  wire [10:0] _T_82273; // @[Modules.scala 53:83:@33130.4]
  wire [10:0] buffer_8_650; // @[Modules.scala 53:83:@33131.4]
  wire [11:0] _T_82275; // @[Modules.scala 53:83:@33133.4]
  wire [10:0] _T_82276; // @[Modules.scala 53:83:@33134.4]
  wire [10:0] buffer_8_651; // @[Modules.scala 53:83:@33135.4]
  wire [11:0] _T_82278; // @[Modules.scala 53:83:@33137.4]
  wire [10:0] _T_82279; // @[Modules.scala 53:83:@33138.4]
  wire [10:0] buffer_8_652; // @[Modules.scala 53:83:@33139.4]
  wire [11:0] _T_82281; // @[Modules.scala 53:83:@33141.4]
  wire [10:0] _T_82282; // @[Modules.scala 53:83:@33142.4]
  wire [10:0] buffer_8_653; // @[Modules.scala 53:83:@33143.4]
  wire [11:0] _T_82284; // @[Modules.scala 53:83:@33145.4]
  wire [10:0] _T_82285; // @[Modules.scala 53:83:@33146.4]
  wire [10:0] buffer_8_654; // @[Modules.scala 53:83:@33147.4]
  wire [11:0] _T_82287; // @[Modules.scala 53:83:@33149.4]
  wire [10:0] _T_82288; // @[Modules.scala 53:83:@33150.4]
  wire [10:0] buffer_8_655; // @[Modules.scala 53:83:@33151.4]
  wire [11:0] _T_82290; // @[Modules.scala 53:83:@33153.4]
  wire [10:0] _T_82291; // @[Modules.scala 53:83:@33154.4]
  wire [10:0] buffer_8_656; // @[Modules.scala 53:83:@33155.4]
  wire [11:0] _T_82293; // @[Modules.scala 53:83:@33157.4]
  wire [10:0] _T_82294; // @[Modules.scala 53:83:@33158.4]
  wire [10:0] buffer_8_657; // @[Modules.scala 53:83:@33159.4]
  wire [11:0] _T_82296; // @[Modules.scala 53:83:@33161.4]
  wire [10:0] _T_82297; // @[Modules.scala 53:83:@33162.4]
  wire [10:0] buffer_8_658; // @[Modules.scala 53:83:@33163.4]
  wire [11:0] _T_82299; // @[Modules.scala 53:83:@33165.4]
  wire [10:0] _T_82300; // @[Modules.scala 53:83:@33166.4]
  wire [10:0] buffer_8_659; // @[Modules.scala 53:83:@33167.4]
  wire [11:0] _T_82302; // @[Modules.scala 53:83:@33169.4]
  wire [10:0] _T_82303; // @[Modules.scala 53:83:@33170.4]
  wire [10:0] buffer_8_660; // @[Modules.scala 53:83:@33171.4]
  wire [11:0] _T_82305; // @[Modules.scala 53:83:@33173.4]
  wire [10:0] _T_82306; // @[Modules.scala 53:83:@33174.4]
  wire [10:0] buffer_8_661; // @[Modules.scala 53:83:@33175.4]
  wire [11:0] _T_82308; // @[Modules.scala 53:83:@33177.4]
  wire [10:0] _T_82309; // @[Modules.scala 53:83:@33178.4]
  wire [10:0] buffer_8_662; // @[Modules.scala 53:83:@33179.4]
  wire [11:0] _T_82311; // @[Modules.scala 53:83:@33181.4]
  wire [10:0] _T_82312; // @[Modules.scala 53:83:@33182.4]
  wire [10:0] buffer_8_663; // @[Modules.scala 53:83:@33183.4]
  wire [11:0] _T_82317; // @[Modules.scala 53:83:@33189.4]
  wire [10:0] _T_82318; // @[Modules.scala 53:83:@33190.4]
  wire [10:0] buffer_8_665; // @[Modules.scala 53:83:@33191.4]
  wire [11:0] _T_82320; // @[Modules.scala 53:83:@33193.4]
  wire [10:0] _T_82321; // @[Modules.scala 53:83:@33194.4]
  wire [10:0] buffer_8_666; // @[Modules.scala 53:83:@33195.4]
  wire [11:0] _T_82329; // @[Modules.scala 53:83:@33205.4]
  wire [10:0] _T_82330; // @[Modules.scala 53:83:@33206.4]
  wire [10:0] buffer_8_669; // @[Modules.scala 53:83:@33207.4]
  wire [11:0] _T_82332; // @[Modules.scala 53:83:@33209.4]
  wire [10:0] _T_82333; // @[Modules.scala 53:83:@33210.4]
  wire [10:0] buffer_8_670; // @[Modules.scala 53:83:@33211.4]
  wire [11:0] _T_82335; // @[Modules.scala 53:83:@33213.4]
  wire [10:0] _T_82336; // @[Modules.scala 53:83:@33214.4]
  wire [10:0] buffer_8_671; // @[Modules.scala 53:83:@33215.4]
  wire [11:0] _T_82338; // @[Modules.scala 53:83:@33217.4]
  wire [10:0] _T_82339; // @[Modules.scala 53:83:@33218.4]
  wire [10:0] buffer_8_672; // @[Modules.scala 53:83:@33219.4]
  wire [11:0] _T_82347; // @[Modules.scala 53:83:@33229.4]
  wire [10:0] _T_82348; // @[Modules.scala 53:83:@33230.4]
  wire [10:0] buffer_8_675; // @[Modules.scala 53:83:@33231.4]
  wire [11:0] _T_82368; // @[Modules.scala 53:83:@33257.4]
  wire [10:0] _T_82369; // @[Modules.scala 53:83:@33258.4]
  wire [10:0] buffer_8_682; // @[Modules.scala 53:83:@33259.4]
  wire [11:0] _T_82371; // @[Modules.scala 53:83:@33261.4]
  wire [10:0] _T_82372; // @[Modules.scala 53:83:@33262.4]
  wire [10:0] buffer_8_683; // @[Modules.scala 53:83:@33263.4]
  wire [11:0] _T_82377; // @[Modules.scala 53:83:@33269.4]
  wire [10:0] _T_82378; // @[Modules.scala 53:83:@33270.4]
  wire [10:0] buffer_8_685; // @[Modules.scala 53:83:@33271.4]
  wire [11:0] _T_82380; // @[Modules.scala 56:109:@33273.4]
  wire [10:0] _T_82381; // @[Modules.scala 56:109:@33274.4]
  wire [10:0] buffer_8_686; // @[Modules.scala 56:109:@33275.4]
  wire [11:0] _T_82383; // @[Modules.scala 56:109:@33277.4]
  wire [10:0] _T_82384; // @[Modules.scala 56:109:@33278.4]
  wire [10:0] buffer_8_687; // @[Modules.scala 56:109:@33279.4]
  wire [11:0] _T_82386; // @[Modules.scala 56:109:@33281.4]
  wire [10:0] _T_82387; // @[Modules.scala 56:109:@33282.4]
  wire [10:0] buffer_8_688; // @[Modules.scala 56:109:@33283.4]
  wire [11:0] _T_82389; // @[Modules.scala 56:109:@33285.4]
  wire [10:0] _T_82390; // @[Modules.scala 56:109:@33286.4]
  wire [10:0] buffer_8_689; // @[Modules.scala 56:109:@33287.4]
  wire [11:0] _T_82395; // @[Modules.scala 56:109:@33293.4]
  wire [10:0] _T_82396; // @[Modules.scala 56:109:@33294.4]
  wire [10:0] buffer_8_691; // @[Modules.scala 56:109:@33295.4]
  wire [11:0] _T_82398; // @[Modules.scala 56:109:@33297.4]
  wire [10:0] _T_82399; // @[Modules.scala 56:109:@33298.4]
  wire [10:0] buffer_8_692; // @[Modules.scala 56:109:@33299.4]
  wire [11:0] _T_82401; // @[Modules.scala 56:109:@33301.4]
  wire [10:0] _T_82402; // @[Modules.scala 56:109:@33302.4]
  wire [10:0] buffer_8_693; // @[Modules.scala 56:109:@33303.4]
  wire [11:0] _T_82404; // @[Modules.scala 56:109:@33305.4]
  wire [10:0] _T_82405; // @[Modules.scala 56:109:@33306.4]
  wire [10:0] buffer_8_694; // @[Modules.scala 56:109:@33307.4]
  wire [11:0] _T_82410; // @[Modules.scala 56:109:@33313.4]
  wire [10:0] _T_82411; // @[Modules.scala 56:109:@33314.4]
  wire [10:0] buffer_8_696; // @[Modules.scala 56:109:@33315.4]
  wire [11:0] _T_82413; // @[Modules.scala 56:109:@33317.4]
  wire [10:0] _T_82414; // @[Modules.scala 56:109:@33318.4]
  wire [10:0] buffer_8_697; // @[Modules.scala 56:109:@33319.4]
  wire [11:0] _T_82416; // @[Modules.scala 56:109:@33321.4]
  wire [10:0] _T_82417; // @[Modules.scala 56:109:@33322.4]
  wire [10:0] buffer_8_698; // @[Modules.scala 56:109:@33323.4]
  wire [11:0] _T_82419; // @[Modules.scala 56:109:@33325.4]
  wire [10:0] _T_82420; // @[Modules.scala 56:109:@33326.4]
  wire [10:0] buffer_8_699; // @[Modules.scala 56:109:@33327.4]
  wire [11:0] _T_82422; // @[Modules.scala 56:109:@33329.4]
  wire [10:0] _T_82423; // @[Modules.scala 56:109:@33330.4]
  wire [10:0] buffer_8_700; // @[Modules.scala 56:109:@33331.4]
  wire [11:0] _T_82425; // @[Modules.scala 56:109:@33333.4]
  wire [10:0] _T_82426; // @[Modules.scala 56:109:@33334.4]
  wire [10:0] buffer_8_701; // @[Modules.scala 56:109:@33335.4]
  wire [11:0] _T_82428; // @[Modules.scala 56:109:@33337.4]
  wire [10:0] _T_82429; // @[Modules.scala 56:109:@33338.4]
  wire [10:0] buffer_8_702; // @[Modules.scala 56:109:@33339.4]
  wire [11:0] _T_82431; // @[Modules.scala 56:109:@33341.4]
  wire [10:0] _T_82432; // @[Modules.scala 56:109:@33342.4]
  wire [10:0] buffer_8_703; // @[Modules.scala 56:109:@33343.4]
  wire [11:0] _T_82434; // @[Modules.scala 56:109:@33345.4]
  wire [10:0] _T_82435; // @[Modules.scala 56:109:@33346.4]
  wire [10:0] buffer_8_704; // @[Modules.scala 56:109:@33347.4]
  wire [11:0] _T_82437; // @[Modules.scala 56:109:@33349.4]
  wire [10:0] _T_82438; // @[Modules.scala 56:109:@33350.4]
  wire [10:0] buffer_8_705; // @[Modules.scala 56:109:@33351.4]
  wire [11:0] _T_82440; // @[Modules.scala 56:109:@33353.4]
  wire [10:0] _T_82441; // @[Modules.scala 56:109:@33354.4]
  wire [10:0] buffer_8_706; // @[Modules.scala 56:109:@33355.4]
  wire [11:0] _T_82443; // @[Modules.scala 56:109:@33357.4]
  wire [10:0] _T_82444; // @[Modules.scala 56:109:@33358.4]
  wire [10:0] buffer_8_707; // @[Modules.scala 56:109:@33359.4]
  wire [11:0] _T_82446; // @[Modules.scala 56:109:@33361.4]
  wire [10:0] _T_82447; // @[Modules.scala 56:109:@33362.4]
  wire [10:0] buffer_8_708; // @[Modules.scala 56:109:@33363.4]
  wire [11:0] _T_82449; // @[Modules.scala 56:109:@33365.4]
  wire [10:0] _T_82450; // @[Modules.scala 56:109:@33366.4]
  wire [10:0] buffer_8_709; // @[Modules.scala 56:109:@33367.4]
  wire [11:0] _T_82452; // @[Modules.scala 56:109:@33369.4]
  wire [10:0] _T_82453; // @[Modules.scala 56:109:@33370.4]
  wire [10:0] buffer_8_710; // @[Modules.scala 56:109:@33371.4]
  wire [11:0] _T_82455; // @[Modules.scala 56:109:@33373.4]
  wire [10:0] _T_82456; // @[Modules.scala 56:109:@33374.4]
  wire [10:0] buffer_8_711; // @[Modules.scala 56:109:@33375.4]
  wire [11:0] _T_82458; // @[Modules.scala 56:109:@33377.4]
  wire [10:0] _T_82459; // @[Modules.scala 56:109:@33378.4]
  wire [10:0] buffer_8_712; // @[Modules.scala 56:109:@33379.4]
  wire [11:0] _T_82461; // @[Modules.scala 56:109:@33381.4]
  wire [10:0] _T_82462; // @[Modules.scala 56:109:@33382.4]
  wire [10:0] buffer_8_713; // @[Modules.scala 56:109:@33383.4]
  wire [11:0] _T_82464; // @[Modules.scala 56:109:@33385.4]
  wire [10:0] _T_82465; // @[Modules.scala 56:109:@33386.4]
  wire [10:0] buffer_8_714; // @[Modules.scala 56:109:@33387.4]
  wire [11:0] _T_82467; // @[Modules.scala 56:109:@33389.4]
  wire [10:0] _T_82468; // @[Modules.scala 56:109:@33390.4]
  wire [10:0] buffer_8_715; // @[Modules.scala 56:109:@33391.4]
  wire [11:0] _T_82470; // @[Modules.scala 56:109:@33393.4]
  wire [10:0] _T_82471; // @[Modules.scala 56:109:@33394.4]
  wire [10:0] buffer_8_716; // @[Modules.scala 56:109:@33395.4]
  wire [11:0] _T_82473; // @[Modules.scala 56:109:@33397.4]
  wire [10:0] _T_82474; // @[Modules.scala 56:109:@33398.4]
  wire [10:0] buffer_8_717; // @[Modules.scala 56:109:@33399.4]
  wire [11:0] _T_82476; // @[Modules.scala 56:109:@33401.4]
  wire [10:0] _T_82477; // @[Modules.scala 56:109:@33402.4]
  wire [10:0] buffer_8_718; // @[Modules.scala 56:109:@33403.4]
  wire [11:0] _T_82479; // @[Modules.scala 56:109:@33405.4]
  wire [10:0] _T_82480; // @[Modules.scala 56:109:@33406.4]
  wire [10:0] buffer_8_719; // @[Modules.scala 56:109:@33407.4]
  wire [11:0] _T_82482; // @[Modules.scala 56:109:@33409.4]
  wire [10:0] _T_82483; // @[Modules.scala 56:109:@33410.4]
  wire [10:0] buffer_8_720; // @[Modules.scala 56:109:@33411.4]
  wire [11:0] _T_82485; // @[Modules.scala 56:109:@33413.4]
  wire [10:0] _T_82486; // @[Modules.scala 56:109:@33414.4]
  wire [10:0] buffer_8_721; // @[Modules.scala 56:109:@33415.4]
  wire [11:0] _T_82488; // @[Modules.scala 56:109:@33417.4]
  wire [10:0] _T_82489; // @[Modules.scala 56:109:@33418.4]
  wire [10:0] buffer_8_722; // @[Modules.scala 56:109:@33419.4]
  wire [11:0] _T_82491; // @[Modules.scala 56:109:@33421.4]
  wire [10:0] _T_82492; // @[Modules.scala 56:109:@33422.4]
  wire [10:0] buffer_8_723; // @[Modules.scala 56:109:@33423.4]
  wire [11:0] _T_82494; // @[Modules.scala 56:109:@33425.4]
  wire [10:0] _T_82495; // @[Modules.scala 56:109:@33426.4]
  wire [10:0] buffer_8_724; // @[Modules.scala 56:109:@33427.4]
  wire [11:0] _T_82497; // @[Modules.scala 56:109:@33429.4]
  wire [10:0] _T_82498; // @[Modules.scala 56:109:@33430.4]
  wire [10:0] buffer_8_725; // @[Modules.scala 56:109:@33431.4]
  wire [11:0] _T_82500; // @[Modules.scala 56:109:@33433.4]
  wire [10:0] _T_82501; // @[Modules.scala 56:109:@33434.4]
  wire [10:0] buffer_8_726; // @[Modules.scala 56:109:@33435.4]
  wire [11:0] _T_82503; // @[Modules.scala 56:109:@33437.4]
  wire [10:0] _T_82504; // @[Modules.scala 56:109:@33438.4]
  wire [10:0] buffer_8_727; // @[Modules.scala 56:109:@33439.4]
  wire [11:0] _T_82506; // @[Modules.scala 56:109:@33441.4]
  wire [10:0] _T_82507; // @[Modules.scala 56:109:@33442.4]
  wire [10:0] buffer_8_728; // @[Modules.scala 56:109:@33443.4]
  wire [11:0] _T_82509; // @[Modules.scala 56:109:@33445.4]
  wire [10:0] _T_82510; // @[Modules.scala 56:109:@33446.4]
  wire [10:0] buffer_8_729; // @[Modules.scala 56:109:@33447.4]
  wire [11:0] _T_82515; // @[Modules.scala 56:109:@33453.4]
  wire [10:0] _T_82516; // @[Modules.scala 56:109:@33454.4]
  wire [10:0] buffer_8_731; // @[Modules.scala 56:109:@33455.4]
  wire [11:0] _T_82521; // @[Modules.scala 56:109:@33461.4]
  wire [10:0] _T_82522; // @[Modules.scala 56:109:@33462.4]
  wire [10:0] buffer_8_733; // @[Modules.scala 56:109:@33463.4]
  wire [11:0] _T_82524; // @[Modules.scala 56:109:@33465.4]
  wire [10:0] _T_82525; // @[Modules.scala 56:109:@33466.4]
  wire [10:0] buffer_8_734; // @[Modules.scala 56:109:@33467.4]
  wire [11:0] _T_82527; // @[Modules.scala 63:156:@33470.4]
  wire [10:0] _T_82528; // @[Modules.scala 63:156:@33471.4]
  wire [10:0] buffer_8_736; // @[Modules.scala 63:156:@33472.4]
  wire [11:0] _T_82530; // @[Modules.scala 63:156:@33474.4]
  wire [10:0] _T_82531; // @[Modules.scala 63:156:@33475.4]
  wire [10:0] buffer_8_737; // @[Modules.scala 63:156:@33476.4]
  wire [11:0] _T_82533; // @[Modules.scala 63:156:@33478.4]
  wire [10:0] _T_82534; // @[Modules.scala 63:156:@33479.4]
  wire [10:0] buffer_8_738; // @[Modules.scala 63:156:@33480.4]
  wire [11:0] _T_82536; // @[Modules.scala 63:156:@33482.4]
  wire [10:0] _T_82537; // @[Modules.scala 63:156:@33483.4]
  wire [10:0] buffer_8_739; // @[Modules.scala 63:156:@33484.4]
  wire [11:0] _T_82539; // @[Modules.scala 63:156:@33486.4]
  wire [10:0] _T_82540; // @[Modules.scala 63:156:@33487.4]
  wire [10:0] buffer_8_740; // @[Modules.scala 63:156:@33488.4]
  wire [11:0] _T_82542; // @[Modules.scala 63:156:@33490.4]
  wire [10:0] _T_82543; // @[Modules.scala 63:156:@33491.4]
  wire [10:0] buffer_8_741; // @[Modules.scala 63:156:@33492.4]
  wire [11:0] _T_82545; // @[Modules.scala 63:156:@33494.4]
  wire [10:0] _T_82546; // @[Modules.scala 63:156:@33495.4]
  wire [10:0] buffer_8_742; // @[Modules.scala 63:156:@33496.4]
  wire [11:0] _T_82548; // @[Modules.scala 63:156:@33498.4]
  wire [10:0] _T_82549; // @[Modules.scala 63:156:@33499.4]
  wire [10:0] buffer_8_743; // @[Modules.scala 63:156:@33500.4]
  wire [11:0] _T_82551; // @[Modules.scala 63:156:@33502.4]
  wire [10:0] _T_82552; // @[Modules.scala 63:156:@33503.4]
  wire [10:0] buffer_8_744; // @[Modules.scala 63:156:@33504.4]
  wire [11:0] _T_82554; // @[Modules.scala 63:156:@33506.4]
  wire [10:0] _T_82555; // @[Modules.scala 63:156:@33507.4]
  wire [10:0] buffer_8_745; // @[Modules.scala 63:156:@33508.4]
  wire [11:0] _T_82557; // @[Modules.scala 63:156:@33510.4]
  wire [10:0] _T_82558; // @[Modules.scala 63:156:@33511.4]
  wire [10:0] buffer_8_746; // @[Modules.scala 63:156:@33512.4]
  wire [11:0] _T_82560; // @[Modules.scala 63:156:@33514.4]
  wire [10:0] _T_82561; // @[Modules.scala 63:156:@33515.4]
  wire [10:0] buffer_8_747; // @[Modules.scala 63:156:@33516.4]
  wire [11:0] _T_82563; // @[Modules.scala 63:156:@33518.4]
  wire [10:0] _T_82564; // @[Modules.scala 63:156:@33519.4]
  wire [10:0] buffer_8_748; // @[Modules.scala 63:156:@33520.4]
  wire [11:0] _T_82566; // @[Modules.scala 63:156:@33522.4]
  wire [10:0] _T_82567; // @[Modules.scala 63:156:@33523.4]
  wire [10:0] buffer_8_749; // @[Modules.scala 63:156:@33524.4]
  wire [11:0] _T_82569; // @[Modules.scala 63:156:@33526.4]
  wire [10:0] _T_82570; // @[Modules.scala 63:156:@33527.4]
  wire [10:0] buffer_8_750; // @[Modules.scala 63:156:@33528.4]
  wire [11:0] _T_82572; // @[Modules.scala 63:156:@33530.4]
  wire [10:0] _T_82573; // @[Modules.scala 63:156:@33531.4]
  wire [10:0] buffer_8_751; // @[Modules.scala 63:156:@33532.4]
  wire [11:0] _T_82575; // @[Modules.scala 63:156:@33534.4]
  wire [10:0] _T_82576; // @[Modules.scala 63:156:@33535.4]
  wire [10:0] buffer_8_752; // @[Modules.scala 63:156:@33536.4]
  wire [11:0] _T_82578; // @[Modules.scala 63:156:@33538.4]
  wire [10:0] _T_82579; // @[Modules.scala 63:156:@33539.4]
  wire [10:0] buffer_8_753; // @[Modules.scala 63:156:@33540.4]
  wire [11:0] _T_82581; // @[Modules.scala 63:156:@33542.4]
  wire [10:0] _T_82582; // @[Modules.scala 63:156:@33543.4]
  wire [10:0] buffer_8_754; // @[Modules.scala 63:156:@33544.4]
  wire [11:0] _T_82584; // @[Modules.scala 63:156:@33546.4]
  wire [10:0] _T_82585; // @[Modules.scala 63:156:@33547.4]
  wire [10:0] buffer_8_755; // @[Modules.scala 63:156:@33548.4]
  wire [11:0] _T_82587; // @[Modules.scala 63:156:@33550.4]
  wire [10:0] _T_82588; // @[Modules.scala 63:156:@33551.4]
  wire [10:0] buffer_8_756; // @[Modules.scala 63:156:@33552.4]
  wire [11:0] _T_82590; // @[Modules.scala 63:156:@33554.4]
  wire [10:0] _T_82591; // @[Modules.scala 63:156:@33555.4]
  wire [10:0] buffer_8_757; // @[Modules.scala 63:156:@33556.4]
  wire [11:0] _T_82593; // @[Modules.scala 63:156:@33558.4]
  wire [10:0] _T_82594; // @[Modules.scala 63:156:@33559.4]
  wire [10:0] buffer_8_758; // @[Modules.scala 63:156:@33560.4]
  wire [11:0] _T_82596; // @[Modules.scala 63:156:@33562.4]
  wire [10:0] _T_82597; // @[Modules.scala 63:156:@33563.4]
  wire [10:0] buffer_8_759; // @[Modules.scala 63:156:@33564.4]
  wire [11:0] _T_82599; // @[Modules.scala 63:156:@33566.4]
  wire [10:0] _T_82600; // @[Modules.scala 63:156:@33567.4]
  wire [10:0] buffer_8_760; // @[Modules.scala 63:156:@33568.4]
  wire [11:0] _T_82602; // @[Modules.scala 63:156:@33570.4]
  wire [10:0] _T_82603; // @[Modules.scala 63:156:@33571.4]
  wire [10:0] buffer_8_761; // @[Modules.scala 63:156:@33572.4]
  wire [11:0] _T_82605; // @[Modules.scala 63:156:@33574.4]
  wire [10:0] _T_82606; // @[Modules.scala 63:156:@33575.4]
  wire [10:0] buffer_8_762; // @[Modules.scala 63:156:@33576.4]
  wire [11:0] _T_82608; // @[Modules.scala 63:156:@33578.4]
  wire [10:0] _T_82609; // @[Modules.scala 63:156:@33579.4]
  wire [10:0] buffer_8_763; // @[Modules.scala 63:156:@33580.4]
  wire [11:0] _T_82611; // @[Modules.scala 63:156:@33582.4]
  wire [10:0] _T_82612; // @[Modules.scala 63:156:@33583.4]
  wire [10:0] buffer_8_764; // @[Modules.scala 63:156:@33584.4]
  wire [11:0] _T_82614; // @[Modules.scala 63:156:@33586.4]
  wire [10:0] _T_82615; // @[Modules.scala 63:156:@33587.4]
  wire [10:0] buffer_8_765; // @[Modules.scala 63:156:@33588.4]
  wire [11:0] _T_82617; // @[Modules.scala 63:156:@33590.4]
  wire [10:0] _T_82618; // @[Modules.scala 63:156:@33591.4]
  wire [10:0] buffer_8_766; // @[Modules.scala 63:156:@33592.4]
  wire [11:0] _T_82620; // @[Modules.scala 63:156:@33594.4]
  wire [10:0] _T_82621; // @[Modules.scala 63:156:@33595.4]
  wire [10:0] buffer_8_767; // @[Modules.scala 63:156:@33596.4]
  wire [11:0] _T_82623; // @[Modules.scala 63:156:@33598.4]
  wire [10:0] _T_82624; // @[Modules.scala 63:156:@33599.4]
  wire [10:0] buffer_8_768; // @[Modules.scala 63:156:@33600.4]
  wire [11:0] _T_82626; // @[Modules.scala 63:156:@33602.4]
  wire [10:0] _T_82627; // @[Modules.scala 63:156:@33603.4]
  wire [10:0] buffer_8_769; // @[Modules.scala 63:156:@33604.4]
  wire [11:0] _T_82629; // @[Modules.scala 63:156:@33606.4]
  wire [10:0] _T_82630; // @[Modules.scala 63:156:@33607.4]
  wire [10:0] buffer_8_770; // @[Modules.scala 63:156:@33608.4]
  wire [11:0] _T_82632; // @[Modules.scala 63:156:@33610.4]
  wire [10:0] _T_82633; // @[Modules.scala 63:156:@33611.4]
  wire [10:0] buffer_8_771; // @[Modules.scala 63:156:@33612.4]
  wire [11:0] _T_82635; // @[Modules.scala 63:156:@33614.4]
  wire [10:0] _T_82636; // @[Modules.scala 63:156:@33615.4]
  wire [10:0] buffer_8_772; // @[Modules.scala 63:156:@33616.4]
  wire [11:0] _T_82638; // @[Modules.scala 63:156:@33618.4]
  wire [10:0] _T_82639; // @[Modules.scala 63:156:@33619.4]
  wire [10:0] buffer_8_773; // @[Modules.scala 63:156:@33620.4]
  wire [11:0] _T_82641; // @[Modules.scala 63:156:@33622.4]
  wire [10:0] _T_82642; // @[Modules.scala 63:156:@33623.4]
  wire [10:0] buffer_8_774; // @[Modules.scala 63:156:@33624.4]
  wire [11:0] _T_82644; // @[Modules.scala 63:156:@33626.4]
  wire [10:0] _T_82645; // @[Modules.scala 63:156:@33627.4]
  wire [10:0] buffer_8_775; // @[Modules.scala 63:156:@33628.4]
  wire [11:0] _T_82647; // @[Modules.scala 63:156:@33630.4]
  wire [10:0] _T_82648; // @[Modules.scala 63:156:@33631.4]
  wire [10:0] buffer_8_776; // @[Modules.scala 63:156:@33632.4]
  wire [11:0] _T_82650; // @[Modules.scala 63:156:@33634.4]
  wire [10:0] _T_82651; // @[Modules.scala 63:156:@33635.4]
  wire [10:0] buffer_8_777; // @[Modules.scala 63:156:@33636.4]
  wire [11:0] _T_82653; // @[Modules.scala 63:156:@33638.4]
  wire [10:0] _T_82654; // @[Modules.scala 63:156:@33639.4]
  wire [10:0] buffer_8_778; // @[Modules.scala 63:156:@33640.4]
  wire [11:0] _T_82656; // @[Modules.scala 63:156:@33642.4]
  wire [10:0] _T_82657; // @[Modules.scala 63:156:@33643.4]
  wire [10:0] buffer_8_779; // @[Modules.scala 63:156:@33644.4]
  wire [11:0] _T_82659; // @[Modules.scala 63:156:@33646.4]
  wire [10:0] _T_82660; // @[Modules.scala 63:156:@33647.4]
  wire [10:0] buffer_8_780; // @[Modules.scala 63:156:@33648.4]
  wire [11:0] _T_82662; // @[Modules.scala 63:156:@33650.4]
  wire [10:0] _T_82663; // @[Modules.scala 63:156:@33651.4]
  wire [10:0] buffer_8_781; // @[Modules.scala 63:156:@33652.4]
  wire [11:0] _T_82665; // @[Modules.scala 63:156:@33654.4]
  wire [10:0] _T_82666; // @[Modules.scala 63:156:@33655.4]
  wire [10:0] buffer_8_782; // @[Modules.scala 63:156:@33656.4]
  wire [11:0] _T_82668; // @[Modules.scala 63:156:@33658.4]
  wire [10:0] _T_82669; // @[Modules.scala 63:156:@33659.4]
  wire [10:0] buffer_8_783; // @[Modules.scala 63:156:@33660.4]
  wire [5:0] _T_82678; // @[Modules.scala 37:46:@33670.4]
  wire [4:0] _T_82679; // @[Modules.scala 37:46:@33671.4]
  wire [4:0] _T_82680; // @[Modules.scala 37:46:@33672.4]
  wire [5:0] _T_82685; // @[Modules.scala 46:47:@33677.4]
  wire [4:0] _T_82686; // @[Modules.scala 46:47:@33678.4]
  wire [4:0] _T_82687; // @[Modules.scala 46:47:@33679.4]
  wire [5:0] _T_82730; // @[Modules.scala 37:46:@33723.4]
  wire [4:0] _T_82731; // @[Modules.scala 37:46:@33724.4]
  wire [4:0] _T_82732; // @[Modules.scala 37:46:@33725.4]
  wire [5:0] _T_82858; // @[Modules.scala 43:47:@33875.4]
  wire [4:0] _T_82859; // @[Modules.scala 43:47:@33876.4]
  wire [4:0] _T_82860; // @[Modules.scala 43:47:@33877.4]
  wire [5:0] _T_82996; // @[Modules.scala 43:47:@34038.4]
  wire [4:0] _T_82997; // @[Modules.scala 43:47:@34039.4]
  wire [4:0] _T_82998; // @[Modules.scala 43:47:@34040.4]
  wire [5:0] _T_83013; // @[Modules.scala 43:47:@34056.4]
  wire [4:0] _T_83014; // @[Modules.scala 43:47:@34057.4]
  wire [4:0] _T_83015; // @[Modules.scala 43:47:@34058.4]
  wire [5:0] _T_83054; // @[Modules.scala 43:47:@34099.4]
  wire [4:0] _T_83055; // @[Modules.scala 43:47:@34100.4]
  wire [4:0] _T_83056; // @[Modules.scala 43:47:@34101.4]
  wire [5:0] _T_83084; // @[Modules.scala 43:47:@34132.4]
  wire [4:0] _T_83085; // @[Modules.scala 43:47:@34133.4]
  wire [4:0] _T_83086; // @[Modules.scala 43:47:@34134.4]
  wire [5:0] _T_83197; // @[Modules.scala 40:46:@34257.4]
  wire [4:0] _T_83198; // @[Modules.scala 40:46:@34258.4]
  wire [4:0] _T_83199; // @[Modules.scala 40:46:@34259.4]
  wire [5:0] _T_83241; // @[Modules.scala 43:47:@34304.4]
  wire [4:0] _T_83242; // @[Modules.scala 43:47:@34305.4]
  wire [4:0] _T_83243; // @[Modules.scala 43:47:@34306.4]
  wire [5:0] _T_83294; // @[Modules.scala 40:46:@34363.4]
  wire [4:0] _T_83295; // @[Modules.scala 40:46:@34364.4]
  wire [4:0] _T_83296; // @[Modules.scala 40:46:@34365.4]
  wire [5:0] _T_83399; // @[Modules.scala 40:46:@34475.4]
  wire [4:0] _T_83400; // @[Modules.scala 40:46:@34476.4]
  wire [4:0] _T_83401; // @[Modules.scala 40:46:@34477.4]
  wire [5:0] _T_83415; // @[Modules.scala 40:46:@34494.4]
  wire [4:0] _T_83416; // @[Modules.scala 40:46:@34495.4]
  wire [4:0] _T_83417; // @[Modules.scala 40:46:@34496.4]
  wire [5:0] _T_83443; // @[Modules.scala 43:47:@34522.4]
  wire [4:0] _T_83444; // @[Modules.scala 43:47:@34523.4]
  wire [4:0] _T_83445; // @[Modules.scala 43:47:@34524.4]
  wire [5:0] _T_83509; // @[Modules.scala 43:47:@34596.4]
  wire [4:0] _T_83510; // @[Modules.scala 43:47:@34597.4]
  wire [4:0] _T_83511; // @[Modules.scala 43:47:@34598.4]
  wire [5:0] _T_83588; // @[Modules.scala 40:46:@34685.4]
  wire [4:0] _T_83589; // @[Modules.scala 40:46:@34686.4]
  wire [4:0] _T_83590; // @[Modules.scala 40:46:@34687.4]
  wire [5:0] _T_83635; // @[Modules.scala 40:46:@34736.4]
  wire [4:0] _T_83636; // @[Modules.scala 40:46:@34737.4]
  wire [4:0] _T_83637; // @[Modules.scala 40:46:@34738.4]
  wire [5:0] _T_83765; // @[Modules.scala 40:46:@34879.4]
  wire [4:0] _T_83766; // @[Modules.scala 40:46:@34880.4]
  wire [4:0] _T_83767; // @[Modules.scala 40:46:@34881.4]
  wire [5:0] _T_83858; // @[Modules.scala 40:46:@34982.4]
  wire [4:0] _T_83859; // @[Modules.scala 40:46:@34983.4]
  wire [4:0] _T_83860; // @[Modules.scala 40:46:@34984.4]
  wire [5:0] _T_84008; // @[Modules.scala 43:47:@35161.4]
  wire [4:0] _T_84009; // @[Modules.scala 43:47:@35162.4]
  wire [4:0] _T_84010; // @[Modules.scala 43:47:@35163.4]
  wire [5:0] _T_84067; // @[Modules.scala 40:46:@35235.4]
  wire [4:0] _T_84068; // @[Modules.scala 40:46:@35236.4]
  wire [4:0] _T_84069; // @[Modules.scala 40:46:@35237.4]
  wire [5:0] _T_84079; // @[Modules.scala 40:46:@35251.4]
  wire [4:0] _T_84080; // @[Modules.scala 40:46:@35252.4]
  wire [4:0] _T_84081; // @[Modules.scala 40:46:@35253.4]
  wire [5:0] _T_84086; // @[Modules.scala 43:47:@35258.4]
  wire [4:0] _T_84087; // @[Modules.scala 43:47:@35259.4]
  wire [4:0] _T_84088; // @[Modules.scala 43:47:@35260.4]
  wire [5:0] _T_84151; // @[Modules.scala 43:47:@35333.4]
  wire [4:0] _T_84152; // @[Modules.scala 43:47:@35334.4]
  wire [4:0] _T_84153; // @[Modules.scala 43:47:@35335.4]
  wire [5:0] _T_84261; // @[Modules.scala 43:47:@35461.4]
  wire [4:0] _T_84262; // @[Modules.scala 43:47:@35462.4]
  wire [4:0] _T_84263; // @[Modules.scala 43:47:@35463.4]
  wire [5:0] _T_84264; // @[Modules.scala 40:46:@35465.4]
  wire [4:0] _T_84265; // @[Modules.scala 40:46:@35466.4]
  wire [4:0] _T_84266; // @[Modules.scala 40:46:@35467.4]
  wire [5:0] _T_84293; // @[Modules.scala 40:46:@35499.4]
  wire [4:0] _T_84294; // @[Modules.scala 40:46:@35500.4]
  wire [4:0] _T_84295; // @[Modules.scala 40:46:@35501.4]
  wire [5:0] _T_84303; // @[Modules.scala 40:46:@35510.4]
  wire [4:0] _T_84304; // @[Modules.scala 40:46:@35511.4]
  wire [4:0] _T_84305; // @[Modules.scala 40:46:@35512.4]
  wire [5:0] _T_84317; // @[Modules.scala 43:47:@35524.4]
  wire [4:0] _T_84318; // @[Modules.scala 43:47:@35525.4]
  wire [4:0] _T_84319; // @[Modules.scala 43:47:@35526.4]
  wire [5:0] _T_84345; // @[Modules.scala 43:47:@35552.4]
  wire [4:0] _T_84346; // @[Modules.scala 43:47:@35553.4]
  wire [4:0] _T_84347; // @[Modules.scala 43:47:@35554.4]
  wire [5:0] _T_84355; // @[Modules.scala 43:47:@35563.4]
  wire [4:0] _T_84356; // @[Modules.scala 43:47:@35564.4]
  wire [4:0] _T_84357; // @[Modules.scala 43:47:@35565.4]
  wire [5:0] _T_84430; // @[Modules.scala 46:47:@35642.4]
  wire [4:0] _T_84431; // @[Modules.scala 46:47:@35643.4]
  wire [4:0] _T_84432; // @[Modules.scala 46:47:@35644.4]
  wire [5:0] _T_84436; // @[Modules.scala 40:46:@35650.4]
  wire [4:0] _T_84437; // @[Modules.scala 40:46:@35651.4]
  wire [4:0] _T_84438; // @[Modules.scala 40:46:@35652.4]
  wire [5:0] _T_84450; // @[Modules.scala 43:47:@35664.4]
  wire [4:0] _T_84451; // @[Modules.scala 43:47:@35665.4]
  wire [4:0] _T_84452; // @[Modules.scala 43:47:@35666.4]
  wire [5:0] _T_84472; // @[Modules.scala 40:46:@35691.4]
  wire [4:0] _T_84473; // @[Modules.scala 40:46:@35692.4]
  wire [4:0] _T_84474; // @[Modules.scala 40:46:@35693.4]
  wire [10:0] buffer_9_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84487; // @[Modules.scala 50:57:@35711.4]
  wire [10:0] _T_84488; // @[Modules.scala 50:57:@35712.4]
  wire [10:0] buffer_9_392; // @[Modules.scala 50:57:@35713.4]
  wire [10:0] buffer_9_2; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84490; // @[Modules.scala 50:57:@35715.4]
  wire [10:0] _T_84491; // @[Modules.scala 50:57:@35716.4]
  wire [10:0] buffer_9_393; // @[Modules.scala 50:57:@35717.4]
  wire [11:0] _T_84493; // @[Modules.scala 50:57:@35719.4]
  wire [10:0] _T_84494; // @[Modules.scala 50:57:@35720.4]
  wire [10:0] buffer_9_394; // @[Modules.scala 50:57:@35721.4]
  wire [10:0] buffer_9_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84499; // @[Modules.scala 50:57:@35727.4]
  wire [10:0] _T_84500; // @[Modules.scala 50:57:@35728.4]
  wire [10:0] buffer_9_396; // @[Modules.scala 50:57:@35729.4]
  wire [11:0] _T_84505; // @[Modules.scala 50:57:@35735.4]
  wire [10:0] _T_84506; // @[Modules.scala 50:57:@35736.4]
  wire [10:0] buffer_9_398; // @[Modules.scala 50:57:@35737.4]
  wire [11:0] _T_84520; // @[Modules.scala 50:57:@35755.4]
  wire [10:0] _T_84521; // @[Modules.scala 50:57:@35756.4]
  wire [10:0] buffer_9_403; // @[Modules.scala 50:57:@35757.4]
  wire [10:0] buffer_9_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84547; // @[Modules.scala 50:57:@35791.4]
  wire [10:0] _T_84548; // @[Modules.scala 50:57:@35792.4]
  wire [10:0] buffer_9_412; // @[Modules.scala 50:57:@35793.4]
  wire [11:0] _T_84571; // @[Modules.scala 50:57:@35823.4]
  wire [10:0] _T_84572; // @[Modules.scala 50:57:@35824.4]
  wire [10:0] buffer_9_420; // @[Modules.scala 50:57:@35825.4]
  wire [11:0] _T_84589; // @[Modules.scala 50:57:@35847.4]
  wire [10:0] _T_84590; // @[Modules.scala 50:57:@35848.4]
  wire [10:0] buffer_9_426; // @[Modules.scala 50:57:@35849.4]
  wire [10:0] buffer_9_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84598; // @[Modules.scala 50:57:@35859.4]
  wire [10:0] _T_84599; // @[Modules.scala 50:57:@35860.4]
  wire [10:0] buffer_9_429; // @[Modules.scala 50:57:@35861.4]
  wire [11:0] _T_84601; // @[Modules.scala 50:57:@35863.4]
  wire [10:0] _T_84602; // @[Modules.scala 50:57:@35864.4]
  wire [10:0] buffer_9_430; // @[Modules.scala 50:57:@35865.4]
  wire [10:0] buffer_9_78; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84604; // @[Modules.scala 50:57:@35867.4]
  wire [10:0] _T_84605; // @[Modules.scala 50:57:@35868.4]
  wire [10:0] buffer_9_431; // @[Modules.scala 50:57:@35869.4]
  wire [11:0] _T_84607; // @[Modules.scala 50:57:@35871.4]
  wire [10:0] _T_84608; // @[Modules.scala 50:57:@35872.4]
  wire [10:0] buffer_9_432; // @[Modules.scala 50:57:@35873.4]
  wire [10:0] buffer_9_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84613; // @[Modules.scala 50:57:@35879.4]
  wire [10:0] _T_84614; // @[Modules.scala 50:57:@35880.4]
  wire [10:0] buffer_9_434; // @[Modules.scala 50:57:@35881.4]
  wire [10:0] buffer_9_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84622; // @[Modules.scala 50:57:@35891.4]
  wire [10:0] _T_84623; // @[Modules.scala 50:57:@35892.4]
  wire [10:0] buffer_9_437; // @[Modules.scala 50:57:@35893.4]
  wire [11:0] _T_84628; // @[Modules.scala 50:57:@35899.4]
  wire [10:0] _T_84629; // @[Modules.scala 50:57:@35900.4]
  wire [10:0] buffer_9_439; // @[Modules.scala 50:57:@35901.4]
  wire [11:0] _T_84631; // @[Modules.scala 50:57:@35903.4]
  wire [10:0] _T_84632; // @[Modules.scala 50:57:@35904.4]
  wire [10:0] buffer_9_440; // @[Modules.scala 50:57:@35905.4]
  wire [11:0] _T_84640; // @[Modules.scala 50:57:@35915.4]
  wire [10:0] _T_84641; // @[Modules.scala 50:57:@35916.4]
  wire [10:0] buffer_9_443; // @[Modules.scala 50:57:@35917.4]
  wire [11:0] _T_84646; // @[Modules.scala 50:57:@35923.4]
  wire [10:0] _T_84647; // @[Modules.scala 50:57:@35924.4]
  wire [10:0] buffer_9_445; // @[Modules.scala 50:57:@35925.4]
  wire [11:0] _T_84649; // @[Modules.scala 50:57:@35927.4]
  wire [10:0] _T_84650; // @[Modules.scala 50:57:@35928.4]
  wire [10:0] buffer_9_446; // @[Modules.scala 50:57:@35929.4]
  wire [11:0] _T_84652; // @[Modules.scala 50:57:@35931.4]
  wire [10:0] _T_84653; // @[Modules.scala 50:57:@35932.4]
  wire [10:0] buffer_9_447; // @[Modules.scala 50:57:@35933.4]
  wire [11:0] _T_84655; // @[Modules.scala 50:57:@35935.4]
  wire [10:0] _T_84656; // @[Modules.scala 50:57:@35936.4]
  wire [10:0] buffer_9_448; // @[Modules.scala 50:57:@35937.4]
  wire [10:0] buffer_9_114; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84658; // @[Modules.scala 50:57:@35939.4]
  wire [10:0] _T_84659; // @[Modules.scala 50:57:@35940.4]
  wire [10:0] buffer_9_449; // @[Modules.scala 50:57:@35941.4]
  wire [11:0] _T_84664; // @[Modules.scala 50:57:@35947.4]
  wire [10:0] _T_84665; // @[Modules.scala 50:57:@35948.4]
  wire [10:0] buffer_9_451; // @[Modules.scala 50:57:@35949.4]
  wire [10:0] buffer_9_122; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84670; // @[Modules.scala 50:57:@35955.4]
  wire [10:0] _T_84671; // @[Modules.scala 50:57:@35956.4]
  wire [10:0] buffer_9_453; // @[Modules.scala 50:57:@35957.4]
  wire [11:0] _T_84679; // @[Modules.scala 50:57:@35967.4]
  wire [10:0] _T_84680; // @[Modules.scala 50:57:@35968.4]
  wire [10:0] buffer_9_456; // @[Modules.scala 50:57:@35969.4]
  wire [10:0] buffer_9_133; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84685; // @[Modules.scala 50:57:@35975.4]
  wire [10:0] _T_84686; // @[Modules.scala 50:57:@35976.4]
  wire [10:0] buffer_9_458; // @[Modules.scala 50:57:@35977.4]
  wire [11:0] _T_84694; // @[Modules.scala 50:57:@35987.4]
  wire [10:0] _T_84695; // @[Modules.scala 50:57:@35988.4]
  wire [10:0] buffer_9_461; // @[Modules.scala 50:57:@35989.4]
  wire [11:0] _T_84697; // @[Modules.scala 50:57:@35991.4]
  wire [10:0] _T_84698; // @[Modules.scala 50:57:@35992.4]
  wire [10:0] buffer_9_462; // @[Modules.scala 50:57:@35993.4]
  wire [11:0] _T_84700; // @[Modules.scala 50:57:@35995.4]
  wire [10:0] _T_84701; // @[Modules.scala 50:57:@35996.4]
  wire [10:0] buffer_9_463; // @[Modules.scala 50:57:@35997.4]
  wire [11:0] _T_84712; // @[Modules.scala 50:57:@36011.4]
  wire [10:0] _T_84713; // @[Modules.scala 50:57:@36012.4]
  wire [10:0] buffer_9_467; // @[Modules.scala 50:57:@36013.4]
  wire [10:0] buffer_9_152; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84715; // @[Modules.scala 50:57:@36015.4]
  wire [10:0] _T_84716; // @[Modules.scala 50:57:@36016.4]
  wire [10:0] buffer_9_468; // @[Modules.scala 50:57:@36017.4]
  wire [10:0] buffer_9_156; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84721; // @[Modules.scala 50:57:@36023.4]
  wire [10:0] _T_84722; // @[Modules.scala 50:57:@36024.4]
  wire [10:0] buffer_9_470; // @[Modules.scala 50:57:@36025.4]
  wire [10:0] buffer_9_160; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84727; // @[Modules.scala 50:57:@36031.4]
  wire [10:0] _T_84728; // @[Modules.scala 50:57:@36032.4]
  wire [10:0] buffer_9_472; // @[Modules.scala 50:57:@36033.4]
  wire [10:0] buffer_9_174; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84748; // @[Modules.scala 50:57:@36059.4]
  wire [10:0] _T_84749; // @[Modules.scala 50:57:@36060.4]
  wire [10:0] buffer_9_479; // @[Modules.scala 50:57:@36061.4]
  wire [11:0] _T_84751; // @[Modules.scala 50:57:@36063.4]
  wire [10:0] _T_84752; // @[Modules.scala 50:57:@36064.4]
  wire [10:0] buffer_9_480; // @[Modules.scala 50:57:@36065.4]
  wire [11:0] _T_84754; // @[Modules.scala 50:57:@36067.4]
  wire [10:0] _T_84755; // @[Modules.scala 50:57:@36068.4]
  wire [10:0] buffer_9_481; // @[Modules.scala 50:57:@36069.4]
  wire [11:0] _T_84766; // @[Modules.scala 50:57:@36083.4]
  wire [10:0] _T_84767; // @[Modules.scala 50:57:@36084.4]
  wire [10:0] buffer_9_485; // @[Modules.scala 50:57:@36085.4]
  wire [10:0] buffer_9_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84772; // @[Modules.scala 50:57:@36091.4]
  wire [10:0] _T_84773; // @[Modules.scala 50:57:@36092.4]
  wire [10:0] buffer_9_487; // @[Modules.scala 50:57:@36093.4]
  wire [11:0] _T_84778; // @[Modules.scala 50:57:@36099.4]
  wire [10:0] _T_84779; // @[Modules.scala 50:57:@36100.4]
  wire [10:0] buffer_9_489; // @[Modules.scala 50:57:@36101.4]
  wire [11:0] _T_84781; // @[Modules.scala 50:57:@36103.4]
  wire [10:0] _T_84782; // @[Modules.scala 50:57:@36104.4]
  wire [10:0] buffer_9_490; // @[Modules.scala 50:57:@36105.4]
  wire [10:0] buffer_9_200; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84787; // @[Modules.scala 50:57:@36111.4]
  wire [10:0] _T_84788; // @[Modules.scala 50:57:@36112.4]
  wire [10:0] buffer_9_492; // @[Modules.scala 50:57:@36113.4]
  wire [11:0] _T_84805; // @[Modules.scala 50:57:@36135.4]
  wire [10:0] _T_84806; // @[Modules.scala 50:57:@36136.4]
  wire [10:0] buffer_9_498; // @[Modules.scala 50:57:@36137.4]
  wire [11:0] _T_84808; // @[Modules.scala 50:57:@36139.4]
  wire [10:0] _T_84809; // @[Modules.scala 50:57:@36140.4]
  wire [10:0] buffer_9_499; // @[Modules.scala 50:57:@36141.4]
  wire [11:0] _T_84823; // @[Modules.scala 50:57:@36159.4]
  wire [10:0] _T_84824; // @[Modules.scala 50:57:@36160.4]
  wire [10:0] buffer_9_504; // @[Modules.scala 50:57:@36161.4]
  wire [10:0] buffer_9_226; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84826; // @[Modules.scala 50:57:@36163.4]
  wire [10:0] _T_84827; // @[Modules.scala 50:57:@36164.4]
  wire [10:0] buffer_9_505; // @[Modules.scala 50:57:@36165.4]
  wire [11:0] _T_84829; // @[Modules.scala 50:57:@36167.4]
  wire [10:0] _T_84830; // @[Modules.scala 50:57:@36168.4]
  wire [10:0] buffer_9_506; // @[Modules.scala 50:57:@36169.4]
  wire [11:0] _T_84835; // @[Modules.scala 50:57:@36175.4]
  wire [10:0] _T_84836; // @[Modules.scala 50:57:@36176.4]
  wire [10:0] buffer_9_508; // @[Modules.scala 50:57:@36177.4]
  wire [11:0] _T_84847; // @[Modules.scala 50:57:@36191.4]
  wire [10:0] _T_84848; // @[Modules.scala 50:57:@36192.4]
  wire [10:0] buffer_9_512; // @[Modules.scala 50:57:@36193.4]
  wire [10:0] buffer_9_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84853; // @[Modules.scala 50:57:@36199.4]
  wire [10:0] _T_84854; // @[Modules.scala 50:57:@36200.4]
  wire [10:0] buffer_9_514; // @[Modules.scala 50:57:@36201.4]
  wire [11:0] _T_84868; // @[Modules.scala 50:57:@36219.4]
  wire [10:0] _T_84869; // @[Modules.scala 50:57:@36220.4]
  wire [10:0] buffer_9_519; // @[Modules.scala 50:57:@36221.4]
  wire [11:0] _T_84889; // @[Modules.scala 50:57:@36247.4]
  wire [10:0] _T_84890; // @[Modules.scala 50:57:@36248.4]
  wire [10:0] buffer_9_526; // @[Modules.scala 50:57:@36249.4]
  wire [10:0] buffer_9_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84910; // @[Modules.scala 50:57:@36275.4]
  wire [10:0] _T_84911; // @[Modules.scala 50:57:@36276.4]
  wire [10:0] buffer_9_533; // @[Modules.scala 50:57:@36277.4]
  wire [11:0] _T_84913; // @[Modules.scala 50:57:@36279.4]
  wire [10:0] _T_84914; // @[Modules.scala 50:57:@36280.4]
  wire [10:0] buffer_9_534; // @[Modules.scala 50:57:@36281.4]
  wire [11:0] _T_84916; // @[Modules.scala 50:57:@36283.4]
  wire [10:0] _T_84917; // @[Modules.scala 50:57:@36284.4]
  wire [10:0] buffer_9_535; // @[Modules.scala 50:57:@36285.4]
  wire [11:0] _T_84934; // @[Modules.scala 50:57:@36307.4]
  wire [10:0] _T_84935; // @[Modules.scala 50:57:@36308.4]
  wire [10:0] buffer_9_541; // @[Modules.scala 50:57:@36309.4]
  wire [10:0] buffer_9_300; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84937; // @[Modules.scala 50:57:@36311.4]
  wire [10:0] _T_84938; // @[Modules.scala 50:57:@36312.4]
  wire [10:0] buffer_9_542; // @[Modules.scala 50:57:@36313.4]
  wire [10:0] buffer_9_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_9_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84943; // @[Modules.scala 50:57:@36319.4]
  wire [10:0] _T_84944; // @[Modules.scala 50:57:@36320.4]
  wire [10:0] buffer_9_544; // @[Modules.scala 50:57:@36321.4]
  wire [11:0] _T_84955; // @[Modules.scala 50:57:@36335.4]
  wire [10:0] _T_84956; // @[Modules.scala 50:57:@36336.4]
  wire [10:0] buffer_9_548; // @[Modules.scala 50:57:@36337.4]
  wire [11:0] _T_84961; // @[Modules.scala 50:57:@36343.4]
  wire [10:0] _T_84962; // @[Modules.scala 50:57:@36344.4]
  wire [10:0] buffer_9_550; // @[Modules.scala 50:57:@36345.4]
  wire [11:0] _T_84964; // @[Modules.scala 50:57:@36347.4]
  wire [10:0] _T_84965; // @[Modules.scala 50:57:@36348.4]
  wire [10:0] buffer_9_551; // @[Modules.scala 50:57:@36349.4]
  wire [10:0] buffer_9_320; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_84967; // @[Modules.scala 50:57:@36351.4]
  wire [10:0] _T_84968; // @[Modules.scala 50:57:@36352.4]
  wire [10:0] buffer_9_552; // @[Modules.scala 50:57:@36353.4]
  wire [11:0] _T_84976; // @[Modules.scala 50:57:@36363.4]
  wire [10:0] _T_84977; // @[Modules.scala 50:57:@36364.4]
  wire [10:0] buffer_9_555; // @[Modules.scala 50:57:@36365.4]
  wire [11:0] _T_84985; // @[Modules.scala 50:57:@36375.4]
  wire [10:0] _T_84986; // @[Modules.scala 50:57:@36376.4]
  wire [10:0] buffer_9_558; // @[Modules.scala 50:57:@36377.4]
  wire [10:0] buffer_9_346; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_9_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85006; // @[Modules.scala 50:57:@36403.4]
  wire [10:0] _T_85007; // @[Modules.scala 50:57:@36404.4]
  wire [10:0] buffer_9_565; // @[Modules.scala 50:57:@36405.4]
  wire [11:0] _T_85009; // @[Modules.scala 50:57:@36407.4]
  wire [10:0] _T_85010; // @[Modules.scala 50:57:@36408.4]
  wire [10:0] buffer_9_566; // @[Modules.scala 50:57:@36409.4]
  wire [11:0] _T_85012; // @[Modules.scala 50:57:@36411.4]
  wire [10:0] _T_85013; // @[Modules.scala 50:57:@36412.4]
  wire [10:0] buffer_9_567; // @[Modules.scala 50:57:@36413.4]
  wire [10:0] buffer_9_354; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85018; // @[Modules.scala 50:57:@36419.4]
  wire [10:0] _T_85019; // @[Modules.scala 50:57:@36420.4]
  wire [10:0] buffer_9_569; // @[Modules.scala 50:57:@36421.4]
  wire [10:0] buffer_9_356; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85021; // @[Modules.scala 50:57:@36423.4]
  wire [10:0] _T_85022; // @[Modules.scala 50:57:@36424.4]
  wire [10:0] buffer_9_570; // @[Modules.scala 50:57:@36425.4]
  wire [10:0] buffer_9_358; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85024; // @[Modules.scala 50:57:@36427.4]
  wire [10:0] _T_85025; // @[Modules.scala 50:57:@36428.4]
  wire [10:0] buffer_9_571; // @[Modules.scala 50:57:@36429.4]
  wire [10:0] buffer_9_362; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85030; // @[Modules.scala 50:57:@36435.4]
  wire [10:0] _T_85031; // @[Modules.scala 50:57:@36436.4]
  wire [10:0] buffer_9_573; // @[Modules.scala 50:57:@36437.4]
  wire [10:0] buffer_9_364; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85033; // @[Modules.scala 50:57:@36439.4]
  wire [10:0] _T_85034; // @[Modules.scala 50:57:@36440.4]
  wire [10:0] buffer_9_574; // @[Modules.scala 50:57:@36441.4]
  wire [11:0] _T_85045; // @[Modules.scala 50:57:@36455.4]
  wire [10:0] _T_85046; // @[Modules.scala 50:57:@36456.4]
  wire [10:0] buffer_9_578; // @[Modules.scala 50:57:@36457.4]
  wire [11:0] _T_85048; // @[Modules.scala 50:57:@36459.4]
  wire [10:0] _T_85049; // @[Modules.scala 50:57:@36460.4]
  wire [10:0] buffer_9_579; // @[Modules.scala 50:57:@36461.4]
  wire [10:0] buffer_9_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85051; // @[Modules.scala 50:57:@36463.4]
  wire [10:0] _T_85052; // @[Modules.scala 50:57:@36464.4]
  wire [10:0] buffer_9_580; // @[Modules.scala 50:57:@36465.4]
  wire [10:0] buffer_9_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85054; // @[Modules.scala 50:57:@36467.4]
  wire [10:0] _T_85055; // @[Modules.scala 50:57:@36468.4]
  wire [10:0] buffer_9_581; // @[Modules.scala 50:57:@36469.4]
  wire [10:0] buffer_9_381; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85057; // @[Modules.scala 50:57:@36471.4]
  wire [10:0] _T_85058; // @[Modules.scala 50:57:@36472.4]
  wire [10:0] buffer_9_582; // @[Modules.scala 50:57:@36473.4]
  wire [11:0] _T_85060; // @[Modules.scala 50:57:@36475.4]
  wire [10:0] _T_85061; // @[Modules.scala 50:57:@36476.4]
  wire [10:0] buffer_9_583; // @[Modules.scala 50:57:@36477.4]
  wire [10:0] buffer_9_387; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_85066; // @[Modules.scala 50:57:@36483.4]
  wire [10:0] _T_85067; // @[Modules.scala 50:57:@36484.4]
  wire [10:0] buffer_9_585; // @[Modules.scala 50:57:@36485.4]
  wire [11:0] _T_85075; // @[Modules.scala 53:83:@36495.4]
  wire [10:0] _T_85076; // @[Modules.scala 53:83:@36496.4]
  wire [10:0] buffer_9_588; // @[Modules.scala 53:83:@36497.4]
  wire [11:0] _T_85078; // @[Modules.scala 53:83:@36499.4]
  wire [10:0] _T_85079; // @[Modules.scala 53:83:@36500.4]
  wire [10:0] buffer_9_589; // @[Modules.scala 53:83:@36501.4]
  wire [11:0] _T_85081; // @[Modules.scala 53:83:@36503.4]
  wire [10:0] _T_85082; // @[Modules.scala 53:83:@36504.4]
  wire [10:0] buffer_9_590; // @[Modules.scala 53:83:@36505.4]
  wire [11:0] _T_85084; // @[Modules.scala 53:83:@36507.4]
  wire [10:0] _T_85085; // @[Modules.scala 53:83:@36508.4]
  wire [10:0] buffer_9_591; // @[Modules.scala 53:83:@36509.4]
  wire [11:0] _T_85090; // @[Modules.scala 53:83:@36515.4]
  wire [10:0] _T_85091; // @[Modules.scala 53:83:@36516.4]
  wire [10:0] buffer_9_593; // @[Modules.scala 53:83:@36517.4]
  wire [11:0] _T_85093; // @[Modules.scala 53:83:@36519.4]
  wire [10:0] _T_85094; // @[Modules.scala 53:83:@36520.4]
  wire [10:0] buffer_9_594; // @[Modules.scala 53:83:@36521.4]
  wire [11:0] _T_85096; // @[Modules.scala 53:83:@36523.4]
  wire [10:0] _T_85097; // @[Modules.scala 53:83:@36524.4]
  wire [10:0] buffer_9_595; // @[Modules.scala 53:83:@36525.4]
  wire [11:0] _T_85105; // @[Modules.scala 53:83:@36535.4]
  wire [10:0] _T_85106; // @[Modules.scala 53:83:@36536.4]
  wire [10:0] buffer_9_598; // @[Modules.scala 53:83:@36537.4]
  wire [11:0] _T_85117; // @[Modules.scala 53:83:@36551.4]
  wire [10:0] _T_85118; // @[Modules.scala 53:83:@36552.4]
  wire [10:0] buffer_9_602; // @[Modules.scala 53:83:@36553.4]
  wire [11:0] _T_85123; // @[Modules.scala 53:83:@36559.4]
  wire [10:0] _T_85124; // @[Modules.scala 53:83:@36560.4]
  wire [10:0] buffer_9_604; // @[Modules.scala 53:83:@36561.4]
  wire [11:0] _T_85126; // @[Modules.scala 53:83:@36563.4]
  wire [10:0] _T_85127; // @[Modules.scala 53:83:@36564.4]
  wire [10:0] buffer_9_605; // @[Modules.scala 53:83:@36565.4]
  wire [11:0] _T_85129; // @[Modules.scala 53:83:@36567.4]
  wire [10:0] _T_85130; // @[Modules.scala 53:83:@36568.4]
  wire [10:0] buffer_9_606; // @[Modules.scala 53:83:@36569.4]
  wire [11:0] _T_85132; // @[Modules.scala 53:83:@36571.4]
  wire [10:0] _T_85133; // @[Modules.scala 53:83:@36572.4]
  wire [10:0] buffer_9_607; // @[Modules.scala 53:83:@36573.4]
  wire [11:0] _T_85135; // @[Modules.scala 53:83:@36575.4]
  wire [10:0] _T_85136; // @[Modules.scala 53:83:@36576.4]
  wire [10:0] buffer_9_608; // @[Modules.scala 53:83:@36577.4]
  wire [11:0] _T_85138; // @[Modules.scala 53:83:@36579.4]
  wire [10:0] _T_85139; // @[Modules.scala 53:83:@36580.4]
  wire [10:0] buffer_9_609; // @[Modules.scala 53:83:@36581.4]
  wire [11:0] _T_85141; // @[Modules.scala 53:83:@36583.4]
  wire [10:0] _T_85142; // @[Modules.scala 53:83:@36584.4]
  wire [10:0] buffer_9_610; // @[Modules.scala 53:83:@36585.4]
  wire [11:0] _T_85144; // @[Modules.scala 53:83:@36587.4]
  wire [10:0] _T_85145; // @[Modules.scala 53:83:@36588.4]
  wire [10:0] buffer_9_611; // @[Modules.scala 53:83:@36589.4]
  wire [11:0] _T_85147; // @[Modules.scala 53:83:@36591.4]
  wire [10:0] _T_85148; // @[Modules.scala 53:83:@36592.4]
  wire [10:0] buffer_9_612; // @[Modules.scala 53:83:@36593.4]
  wire [11:0] _T_85150; // @[Modules.scala 53:83:@36595.4]
  wire [10:0] _T_85151; // @[Modules.scala 53:83:@36596.4]
  wire [10:0] buffer_9_613; // @[Modules.scala 53:83:@36597.4]
  wire [11:0] _T_85153; // @[Modules.scala 53:83:@36599.4]
  wire [10:0] _T_85154; // @[Modules.scala 53:83:@36600.4]
  wire [10:0] buffer_9_614; // @[Modules.scala 53:83:@36601.4]
  wire [11:0] _T_85156; // @[Modules.scala 53:83:@36603.4]
  wire [10:0] _T_85157; // @[Modules.scala 53:83:@36604.4]
  wire [10:0] buffer_9_615; // @[Modules.scala 53:83:@36605.4]
  wire [11:0] _T_85159; // @[Modules.scala 53:83:@36607.4]
  wire [10:0] _T_85160; // @[Modules.scala 53:83:@36608.4]
  wire [10:0] buffer_9_616; // @[Modules.scala 53:83:@36609.4]
  wire [11:0] _T_85162; // @[Modules.scala 53:83:@36611.4]
  wire [10:0] _T_85163; // @[Modules.scala 53:83:@36612.4]
  wire [10:0] buffer_9_617; // @[Modules.scala 53:83:@36613.4]
  wire [11:0] _T_85165; // @[Modules.scala 53:83:@36615.4]
  wire [10:0] _T_85166; // @[Modules.scala 53:83:@36616.4]
  wire [10:0] buffer_9_618; // @[Modules.scala 53:83:@36617.4]
  wire [11:0] _T_85171; // @[Modules.scala 53:83:@36623.4]
  wire [10:0] _T_85172; // @[Modules.scala 53:83:@36624.4]
  wire [10:0] buffer_9_620; // @[Modules.scala 53:83:@36625.4]
  wire [11:0] _T_85174; // @[Modules.scala 53:83:@36627.4]
  wire [10:0] _T_85175; // @[Modules.scala 53:83:@36628.4]
  wire [10:0] buffer_9_621; // @[Modules.scala 53:83:@36629.4]
  wire [11:0] _T_85177; // @[Modules.scala 53:83:@36631.4]
  wire [10:0] _T_85178; // @[Modules.scala 53:83:@36632.4]
  wire [10:0] buffer_9_622; // @[Modules.scala 53:83:@36633.4]
  wire [11:0] _T_85180; // @[Modules.scala 53:83:@36635.4]
  wire [10:0] _T_85181; // @[Modules.scala 53:83:@36636.4]
  wire [10:0] buffer_9_623; // @[Modules.scala 53:83:@36637.4]
  wire [11:0] _T_85186; // @[Modules.scala 53:83:@36643.4]
  wire [10:0] _T_85187; // @[Modules.scala 53:83:@36644.4]
  wire [10:0] buffer_9_625; // @[Modules.scala 53:83:@36645.4]
  wire [11:0] _T_85189; // @[Modules.scala 53:83:@36647.4]
  wire [10:0] _T_85190; // @[Modules.scala 53:83:@36648.4]
  wire [10:0] buffer_9_626; // @[Modules.scala 53:83:@36649.4]
  wire [11:0] _T_85192; // @[Modules.scala 53:83:@36651.4]
  wire [10:0] _T_85193; // @[Modules.scala 53:83:@36652.4]
  wire [10:0] buffer_9_627; // @[Modules.scala 53:83:@36653.4]
  wire [11:0] _T_85195; // @[Modules.scala 53:83:@36655.4]
  wire [10:0] _T_85196; // @[Modules.scala 53:83:@36656.4]
  wire [10:0] buffer_9_628; // @[Modules.scala 53:83:@36657.4]
  wire [11:0] _T_85198; // @[Modules.scala 53:83:@36659.4]
  wire [10:0] _T_85199; // @[Modules.scala 53:83:@36660.4]
  wire [10:0] buffer_9_629; // @[Modules.scala 53:83:@36661.4]
  wire [11:0] _T_85204; // @[Modules.scala 53:83:@36667.4]
  wire [10:0] _T_85205; // @[Modules.scala 53:83:@36668.4]
  wire [10:0] buffer_9_631; // @[Modules.scala 53:83:@36669.4]
  wire [11:0] _T_85207; // @[Modules.scala 53:83:@36671.4]
  wire [10:0] _T_85208; // @[Modules.scala 53:83:@36672.4]
  wire [10:0] buffer_9_632; // @[Modules.scala 53:83:@36673.4]
  wire [11:0] _T_85213; // @[Modules.scala 53:83:@36679.4]
  wire [10:0] _T_85214; // @[Modules.scala 53:83:@36680.4]
  wire [10:0] buffer_9_634; // @[Modules.scala 53:83:@36681.4]
  wire [11:0] _T_85216; // @[Modules.scala 53:83:@36683.4]
  wire [10:0] _T_85217; // @[Modules.scala 53:83:@36684.4]
  wire [10:0] buffer_9_635; // @[Modules.scala 53:83:@36685.4]
  wire [11:0] _T_85219; // @[Modules.scala 53:83:@36687.4]
  wire [10:0] _T_85220; // @[Modules.scala 53:83:@36688.4]
  wire [10:0] buffer_9_636; // @[Modules.scala 53:83:@36689.4]
  wire [11:0] _T_85222; // @[Modules.scala 53:83:@36691.4]
  wire [10:0] _T_85223; // @[Modules.scala 53:83:@36692.4]
  wire [10:0] buffer_9_637; // @[Modules.scala 53:83:@36693.4]
  wire [11:0] _T_85225; // @[Modules.scala 53:83:@36695.4]
  wire [10:0] _T_85226; // @[Modules.scala 53:83:@36696.4]
  wire [10:0] buffer_9_638; // @[Modules.scala 53:83:@36697.4]
  wire [11:0] _T_85231; // @[Modules.scala 53:83:@36703.4]
  wire [10:0] _T_85232; // @[Modules.scala 53:83:@36704.4]
  wire [10:0] buffer_9_640; // @[Modules.scala 53:83:@36705.4]
  wire [11:0] _T_85234; // @[Modules.scala 53:83:@36707.4]
  wire [10:0] _T_85235; // @[Modules.scala 53:83:@36708.4]
  wire [10:0] buffer_9_641; // @[Modules.scala 53:83:@36709.4]
  wire [11:0] _T_85243; // @[Modules.scala 53:83:@36719.4]
  wire [10:0] _T_85244; // @[Modules.scala 53:83:@36720.4]
  wire [10:0] buffer_9_644; // @[Modules.scala 53:83:@36721.4]
  wire [11:0] _T_85246; // @[Modules.scala 53:83:@36723.4]
  wire [10:0] _T_85247; // @[Modules.scala 53:83:@36724.4]
  wire [10:0] buffer_9_645; // @[Modules.scala 53:83:@36725.4]
  wire [11:0] _T_85249; // @[Modules.scala 53:83:@36727.4]
  wire [10:0] _T_85250; // @[Modules.scala 53:83:@36728.4]
  wire [10:0] buffer_9_646; // @[Modules.scala 53:83:@36729.4]
  wire [11:0] _T_85255; // @[Modules.scala 53:83:@36735.4]
  wire [10:0] _T_85256; // @[Modules.scala 53:83:@36736.4]
  wire [10:0] buffer_9_648; // @[Modules.scala 53:83:@36737.4]
  wire [11:0] _T_85258; // @[Modules.scala 53:83:@36739.4]
  wire [10:0] _T_85259; // @[Modules.scala 53:83:@36740.4]
  wire [10:0] buffer_9_649; // @[Modules.scala 53:83:@36741.4]
  wire [11:0] _T_85264; // @[Modules.scala 53:83:@36747.4]
  wire [10:0] _T_85265; // @[Modules.scala 53:83:@36748.4]
  wire [10:0] buffer_9_651; // @[Modules.scala 53:83:@36749.4]
  wire [11:0] _T_85276; // @[Modules.scala 53:83:@36763.4]
  wire [10:0] _T_85277; // @[Modules.scala 53:83:@36764.4]
  wire [10:0] buffer_9_655; // @[Modules.scala 53:83:@36765.4]
  wire [11:0] _T_85285; // @[Modules.scala 53:83:@36775.4]
  wire [10:0] _T_85286; // @[Modules.scala 53:83:@36776.4]
  wire [10:0] buffer_9_658; // @[Modules.scala 53:83:@36777.4]
  wire [11:0] _T_85288; // @[Modules.scala 53:83:@36779.4]
  wire [10:0] _T_85289; // @[Modules.scala 53:83:@36780.4]
  wire [10:0] buffer_9_659; // @[Modules.scala 53:83:@36781.4]
  wire [11:0] _T_85294; // @[Modules.scala 53:83:@36787.4]
  wire [10:0] _T_85295; // @[Modules.scala 53:83:@36788.4]
  wire [10:0] buffer_9_661; // @[Modules.scala 53:83:@36789.4]
  wire [11:0] _T_85297; // @[Modules.scala 53:83:@36791.4]
  wire [10:0] _T_85298; // @[Modules.scala 53:83:@36792.4]
  wire [10:0] buffer_9_662; // @[Modules.scala 53:83:@36793.4]
  wire [11:0] _T_85300; // @[Modules.scala 53:83:@36795.4]
  wire [10:0] _T_85301; // @[Modules.scala 53:83:@36796.4]
  wire [10:0] buffer_9_663; // @[Modules.scala 53:83:@36797.4]
  wire [11:0] _T_85303; // @[Modules.scala 53:83:@36799.4]
  wire [10:0] _T_85304; // @[Modules.scala 53:83:@36800.4]
  wire [10:0] buffer_9_664; // @[Modules.scala 53:83:@36801.4]
  wire [11:0] _T_85309; // @[Modules.scala 53:83:@36807.4]
  wire [10:0] _T_85310; // @[Modules.scala 53:83:@36808.4]
  wire [10:0] buffer_9_666; // @[Modules.scala 53:83:@36809.4]
  wire [11:0] _T_85312; // @[Modules.scala 53:83:@36811.4]
  wire [10:0] _T_85313; // @[Modules.scala 53:83:@36812.4]
  wire [10:0] buffer_9_667; // @[Modules.scala 53:83:@36813.4]
  wire [11:0] _T_85315; // @[Modules.scala 53:83:@36815.4]
  wire [10:0] _T_85316; // @[Modules.scala 53:83:@36816.4]
  wire [10:0] buffer_9_668; // @[Modules.scala 53:83:@36817.4]
  wire [11:0] _T_85318; // @[Modules.scala 53:83:@36819.4]
  wire [10:0] _T_85319; // @[Modules.scala 53:83:@36820.4]
  wire [10:0] buffer_9_669; // @[Modules.scala 53:83:@36821.4]
  wire [11:0] _T_85324; // @[Modules.scala 53:83:@36827.4]
  wire [10:0] _T_85325; // @[Modules.scala 53:83:@36828.4]
  wire [10:0] buffer_9_671; // @[Modules.scala 53:83:@36829.4]
  wire [11:0] _T_85327; // @[Modules.scala 53:83:@36831.4]
  wire [10:0] _T_85328; // @[Modules.scala 53:83:@36832.4]
  wire [10:0] buffer_9_672; // @[Modules.scala 53:83:@36833.4]
  wire [11:0] _T_85333; // @[Modules.scala 53:83:@36839.4]
  wire [10:0] _T_85334; // @[Modules.scala 53:83:@36840.4]
  wire [10:0] buffer_9_674; // @[Modules.scala 53:83:@36841.4]
  wire [11:0] _T_85336; // @[Modules.scala 53:83:@36843.4]
  wire [10:0] _T_85337; // @[Modules.scala 53:83:@36844.4]
  wire [10:0] buffer_9_675; // @[Modules.scala 53:83:@36845.4]
  wire [11:0] _T_85339; // @[Modules.scala 53:83:@36847.4]
  wire [10:0] _T_85340; // @[Modules.scala 53:83:@36848.4]
  wire [10:0] buffer_9_676; // @[Modules.scala 53:83:@36849.4]
  wire [11:0] _T_85342; // @[Modules.scala 53:83:@36851.4]
  wire [10:0] _T_85343; // @[Modules.scala 53:83:@36852.4]
  wire [10:0] buffer_9_677; // @[Modules.scala 53:83:@36853.4]
  wire [11:0] _T_85345; // @[Modules.scala 53:83:@36855.4]
  wire [10:0] _T_85346; // @[Modules.scala 53:83:@36856.4]
  wire [10:0] buffer_9_678; // @[Modules.scala 53:83:@36857.4]
  wire [11:0] _T_85348; // @[Modules.scala 53:83:@36859.4]
  wire [10:0] _T_85349; // @[Modules.scala 53:83:@36860.4]
  wire [10:0] buffer_9_679; // @[Modules.scala 53:83:@36861.4]
  wire [11:0] _T_85354; // @[Modules.scala 53:83:@36867.4]
  wire [10:0] _T_85355; // @[Modules.scala 53:83:@36868.4]
  wire [10:0] buffer_9_681; // @[Modules.scala 53:83:@36869.4]
  wire [11:0] _T_85357; // @[Modules.scala 53:83:@36871.4]
  wire [10:0] _T_85358; // @[Modules.scala 53:83:@36872.4]
  wire [10:0] buffer_9_682; // @[Modules.scala 53:83:@36873.4]
  wire [11:0] _T_85360; // @[Modules.scala 53:83:@36875.4]
  wire [10:0] _T_85361; // @[Modules.scala 53:83:@36876.4]
  wire [10:0] buffer_9_683; // @[Modules.scala 53:83:@36877.4]
  wire [11:0] _T_85363; // @[Modules.scala 53:83:@36879.4]
  wire [10:0] _T_85364; // @[Modules.scala 53:83:@36880.4]
  wire [10:0] buffer_9_684; // @[Modules.scala 53:83:@36881.4]
  wire [11:0] _T_85369; // @[Modules.scala 56:109:@36887.4]
  wire [10:0] _T_85370; // @[Modules.scala 56:109:@36888.4]
  wire [10:0] buffer_9_686; // @[Modules.scala 56:109:@36889.4]
  wire [11:0] _T_85372; // @[Modules.scala 56:109:@36891.4]
  wire [10:0] _T_85373; // @[Modules.scala 56:109:@36892.4]
  wire [10:0] buffer_9_687; // @[Modules.scala 56:109:@36893.4]
  wire [11:0] _T_85375; // @[Modules.scala 56:109:@36895.4]
  wire [10:0] _T_85376; // @[Modules.scala 56:109:@36896.4]
  wire [10:0] buffer_9_688; // @[Modules.scala 56:109:@36897.4]
  wire [11:0] _T_85378; // @[Modules.scala 56:109:@36899.4]
  wire [10:0] _T_85379; // @[Modules.scala 56:109:@36900.4]
  wire [10:0] buffer_9_689; // @[Modules.scala 56:109:@36901.4]
  wire [11:0] _T_85384; // @[Modules.scala 56:109:@36907.4]
  wire [10:0] _T_85385; // @[Modules.scala 56:109:@36908.4]
  wire [10:0] buffer_9_691; // @[Modules.scala 56:109:@36909.4]
  wire [11:0] _T_85390; // @[Modules.scala 56:109:@36915.4]
  wire [10:0] _T_85391; // @[Modules.scala 56:109:@36916.4]
  wire [10:0] buffer_9_693; // @[Modules.scala 56:109:@36917.4]
  wire [11:0] _T_85393; // @[Modules.scala 56:109:@36919.4]
  wire [10:0] _T_85394; // @[Modules.scala 56:109:@36920.4]
  wire [10:0] buffer_9_694; // @[Modules.scala 56:109:@36921.4]
  wire [11:0] _T_85396; // @[Modules.scala 56:109:@36923.4]
  wire [10:0] _T_85397; // @[Modules.scala 56:109:@36924.4]
  wire [10:0] buffer_9_695; // @[Modules.scala 56:109:@36925.4]
  wire [11:0] _T_85399; // @[Modules.scala 56:109:@36927.4]
  wire [10:0] _T_85400; // @[Modules.scala 56:109:@36928.4]
  wire [10:0] buffer_9_696; // @[Modules.scala 56:109:@36929.4]
  wire [11:0] _T_85402; // @[Modules.scala 56:109:@36931.4]
  wire [10:0] _T_85403; // @[Modules.scala 56:109:@36932.4]
  wire [10:0] buffer_9_697; // @[Modules.scala 56:109:@36933.4]
  wire [11:0] _T_85405; // @[Modules.scala 56:109:@36935.4]
  wire [10:0] _T_85406; // @[Modules.scala 56:109:@36936.4]
  wire [10:0] buffer_9_698; // @[Modules.scala 56:109:@36937.4]
  wire [11:0] _T_85408; // @[Modules.scala 56:109:@36939.4]
  wire [10:0] _T_85409; // @[Modules.scala 56:109:@36940.4]
  wire [10:0] buffer_9_699; // @[Modules.scala 56:109:@36941.4]
  wire [11:0] _T_85411; // @[Modules.scala 56:109:@36943.4]
  wire [10:0] _T_85412; // @[Modules.scala 56:109:@36944.4]
  wire [10:0] buffer_9_700; // @[Modules.scala 56:109:@36945.4]
  wire [11:0] _T_85414; // @[Modules.scala 56:109:@36947.4]
  wire [10:0] _T_85415; // @[Modules.scala 56:109:@36948.4]
  wire [10:0] buffer_9_701; // @[Modules.scala 56:109:@36949.4]
  wire [11:0] _T_85417; // @[Modules.scala 56:109:@36951.4]
  wire [10:0] _T_85418; // @[Modules.scala 56:109:@36952.4]
  wire [10:0] buffer_9_702; // @[Modules.scala 56:109:@36953.4]
  wire [11:0] _T_85420; // @[Modules.scala 56:109:@36955.4]
  wire [10:0] _T_85421; // @[Modules.scala 56:109:@36956.4]
  wire [10:0] buffer_9_703; // @[Modules.scala 56:109:@36957.4]
  wire [11:0] _T_85423; // @[Modules.scala 56:109:@36959.4]
  wire [10:0] _T_85424; // @[Modules.scala 56:109:@36960.4]
  wire [10:0] buffer_9_704; // @[Modules.scala 56:109:@36961.4]
  wire [11:0] _T_85426; // @[Modules.scala 56:109:@36963.4]
  wire [10:0] _T_85427; // @[Modules.scala 56:109:@36964.4]
  wire [10:0] buffer_9_705; // @[Modules.scala 56:109:@36965.4]
  wire [11:0] _T_85429; // @[Modules.scala 56:109:@36967.4]
  wire [10:0] _T_85430; // @[Modules.scala 56:109:@36968.4]
  wire [10:0] buffer_9_706; // @[Modules.scala 56:109:@36969.4]
  wire [11:0] _T_85432; // @[Modules.scala 56:109:@36971.4]
  wire [10:0] _T_85433; // @[Modules.scala 56:109:@36972.4]
  wire [10:0] buffer_9_707; // @[Modules.scala 56:109:@36973.4]
  wire [11:0] _T_85435; // @[Modules.scala 56:109:@36975.4]
  wire [10:0] _T_85436; // @[Modules.scala 56:109:@36976.4]
  wire [10:0] buffer_9_708; // @[Modules.scala 56:109:@36977.4]
  wire [11:0] _T_85438; // @[Modules.scala 56:109:@36979.4]
  wire [10:0] _T_85439; // @[Modules.scala 56:109:@36980.4]
  wire [10:0] buffer_9_709; // @[Modules.scala 56:109:@36981.4]
  wire [11:0] _T_85441; // @[Modules.scala 56:109:@36983.4]
  wire [10:0] _T_85442; // @[Modules.scala 56:109:@36984.4]
  wire [10:0] buffer_9_710; // @[Modules.scala 56:109:@36985.4]
  wire [11:0] _T_85444; // @[Modules.scala 56:109:@36987.4]
  wire [10:0] _T_85445; // @[Modules.scala 56:109:@36988.4]
  wire [10:0] buffer_9_711; // @[Modules.scala 56:109:@36989.4]
  wire [11:0] _T_85447; // @[Modules.scala 56:109:@36991.4]
  wire [10:0] _T_85448; // @[Modules.scala 56:109:@36992.4]
  wire [10:0] buffer_9_712; // @[Modules.scala 56:109:@36993.4]
  wire [11:0] _T_85450; // @[Modules.scala 56:109:@36995.4]
  wire [10:0] _T_85451; // @[Modules.scala 56:109:@36996.4]
  wire [10:0] buffer_9_713; // @[Modules.scala 56:109:@36997.4]
  wire [11:0] _T_85453; // @[Modules.scala 56:109:@36999.4]
  wire [10:0] _T_85454; // @[Modules.scala 56:109:@37000.4]
  wire [10:0] buffer_9_714; // @[Modules.scala 56:109:@37001.4]
  wire [11:0] _T_85456; // @[Modules.scala 56:109:@37003.4]
  wire [10:0] _T_85457; // @[Modules.scala 56:109:@37004.4]
  wire [10:0] buffer_9_715; // @[Modules.scala 56:109:@37005.4]
  wire [11:0] _T_85459; // @[Modules.scala 56:109:@37007.4]
  wire [10:0] _T_85460; // @[Modules.scala 56:109:@37008.4]
  wire [10:0] buffer_9_716; // @[Modules.scala 56:109:@37009.4]
  wire [11:0] _T_85462; // @[Modules.scala 56:109:@37011.4]
  wire [10:0] _T_85463; // @[Modules.scala 56:109:@37012.4]
  wire [10:0] buffer_9_717; // @[Modules.scala 56:109:@37013.4]
  wire [11:0] _T_85465; // @[Modules.scala 56:109:@37015.4]
  wire [10:0] _T_85466; // @[Modules.scala 56:109:@37016.4]
  wire [10:0] buffer_9_718; // @[Modules.scala 56:109:@37017.4]
  wire [11:0] _T_85468; // @[Modules.scala 56:109:@37019.4]
  wire [10:0] _T_85469; // @[Modules.scala 56:109:@37020.4]
  wire [10:0] buffer_9_719; // @[Modules.scala 56:109:@37021.4]
  wire [11:0] _T_85471; // @[Modules.scala 56:109:@37023.4]
  wire [10:0] _T_85472; // @[Modules.scala 56:109:@37024.4]
  wire [10:0] buffer_9_720; // @[Modules.scala 56:109:@37025.4]
  wire [11:0] _T_85474; // @[Modules.scala 56:109:@37027.4]
  wire [10:0] _T_85475; // @[Modules.scala 56:109:@37028.4]
  wire [10:0] buffer_9_721; // @[Modules.scala 56:109:@37029.4]
  wire [11:0] _T_85477; // @[Modules.scala 56:109:@37031.4]
  wire [10:0] _T_85478; // @[Modules.scala 56:109:@37032.4]
  wire [10:0] buffer_9_722; // @[Modules.scala 56:109:@37033.4]
  wire [11:0] _T_85480; // @[Modules.scala 56:109:@37035.4]
  wire [10:0] _T_85481; // @[Modules.scala 56:109:@37036.4]
  wire [10:0] buffer_9_723; // @[Modules.scala 56:109:@37037.4]
  wire [11:0] _T_85483; // @[Modules.scala 56:109:@37039.4]
  wire [10:0] _T_85484; // @[Modules.scala 56:109:@37040.4]
  wire [10:0] buffer_9_724; // @[Modules.scala 56:109:@37041.4]
  wire [11:0] _T_85486; // @[Modules.scala 56:109:@37043.4]
  wire [10:0] _T_85487; // @[Modules.scala 56:109:@37044.4]
  wire [10:0] buffer_9_725; // @[Modules.scala 56:109:@37045.4]
  wire [11:0] _T_85489; // @[Modules.scala 56:109:@37047.4]
  wire [10:0] _T_85490; // @[Modules.scala 56:109:@37048.4]
  wire [10:0] buffer_9_726; // @[Modules.scala 56:109:@37049.4]
  wire [11:0] _T_85492; // @[Modules.scala 56:109:@37051.4]
  wire [10:0] _T_85493; // @[Modules.scala 56:109:@37052.4]
  wire [10:0] buffer_9_727; // @[Modules.scala 56:109:@37053.4]
  wire [11:0] _T_85495; // @[Modules.scala 56:109:@37055.4]
  wire [10:0] _T_85496; // @[Modules.scala 56:109:@37056.4]
  wire [10:0] buffer_9_728; // @[Modules.scala 56:109:@37057.4]
  wire [11:0] _T_85498; // @[Modules.scala 56:109:@37059.4]
  wire [10:0] _T_85499; // @[Modules.scala 56:109:@37060.4]
  wire [10:0] buffer_9_729; // @[Modules.scala 56:109:@37061.4]
  wire [11:0] _T_85501; // @[Modules.scala 56:109:@37063.4]
  wire [10:0] _T_85502; // @[Modules.scala 56:109:@37064.4]
  wire [10:0] buffer_9_730; // @[Modules.scala 56:109:@37065.4]
  wire [11:0] _T_85504; // @[Modules.scala 56:109:@37067.4]
  wire [10:0] _T_85505; // @[Modules.scala 56:109:@37068.4]
  wire [10:0] buffer_9_731; // @[Modules.scala 56:109:@37069.4]
  wire [11:0] _T_85507; // @[Modules.scala 56:109:@37071.4]
  wire [10:0] _T_85508; // @[Modules.scala 56:109:@37072.4]
  wire [10:0] buffer_9_732; // @[Modules.scala 56:109:@37073.4]
  wire [11:0] _T_85510; // @[Modules.scala 56:109:@37075.4]
  wire [10:0] _T_85511; // @[Modules.scala 56:109:@37076.4]
  wire [10:0] buffer_9_733; // @[Modules.scala 56:109:@37077.4]
  wire [11:0] _T_85513; // @[Modules.scala 56:109:@37079.4]
  wire [10:0] _T_85514; // @[Modules.scala 56:109:@37080.4]
  wire [10:0] buffer_9_734; // @[Modules.scala 56:109:@37081.4]
  wire [11:0] _T_85516; // @[Modules.scala 63:156:@37084.4]
  wire [10:0] _T_85517; // @[Modules.scala 63:156:@37085.4]
  wire [10:0] buffer_9_736; // @[Modules.scala 63:156:@37086.4]
  wire [11:0] _T_85519; // @[Modules.scala 63:156:@37088.4]
  wire [10:0] _T_85520; // @[Modules.scala 63:156:@37089.4]
  wire [10:0] buffer_9_737; // @[Modules.scala 63:156:@37090.4]
  wire [11:0] _T_85522; // @[Modules.scala 63:156:@37092.4]
  wire [10:0] _T_85523; // @[Modules.scala 63:156:@37093.4]
  wire [10:0] buffer_9_738; // @[Modules.scala 63:156:@37094.4]
  wire [11:0] _T_85525; // @[Modules.scala 63:156:@37096.4]
  wire [10:0] _T_85526; // @[Modules.scala 63:156:@37097.4]
  wire [10:0] buffer_9_739; // @[Modules.scala 63:156:@37098.4]
  wire [11:0] _T_85528; // @[Modules.scala 63:156:@37100.4]
  wire [10:0] _T_85529; // @[Modules.scala 63:156:@37101.4]
  wire [10:0] buffer_9_740; // @[Modules.scala 63:156:@37102.4]
  wire [11:0] _T_85531; // @[Modules.scala 63:156:@37104.4]
  wire [10:0] _T_85532; // @[Modules.scala 63:156:@37105.4]
  wire [10:0] buffer_9_741; // @[Modules.scala 63:156:@37106.4]
  wire [11:0] _T_85534; // @[Modules.scala 63:156:@37108.4]
  wire [10:0] _T_85535; // @[Modules.scala 63:156:@37109.4]
  wire [10:0] buffer_9_742; // @[Modules.scala 63:156:@37110.4]
  wire [11:0] _T_85537; // @[Modules.scala 63:156:@37112.4]
  wire [10:0] _T_85538; // @[Modules.scala 63:156:@37113.4]
  wire [10:0] buffer_9_743; // @[Modules.scala 63:156:@37114.4]
  wire [11:0] _T_85540; // @[Modules.scala 63:156:@37116.4]
  wire [10:0] _T_85541; // @[Modules.scala 63:156:@37117.4]
  wire [10:0] buffer_9_744; // @[Modules.scala 63:156:@37118.4]
  wire [11:0] _T_85543; // @[Modules.scala 63:156:@37120.4]
  wire [10:0] _T_85544; // @[Modules.scala 63:156:@37121.4]
  wire [10:0] buffer_9_745; // @[Modules.scala 63:156:@37122.4]
  wire [11:0] _T_85546; // @[Modules.scala 63:156:@37124.4]
  wire [10:0] _T_85547; // @[Modules.scala 63:156:@37125.4]
  wire [10:0] buffer_9_746; // @[Modules.scala 63:156:@37126.4]
  wire [11:0] _T_85549; // @[Modules.scala 63:156:@37128.4]
  wire [10:0] _T_85550; // @[Modules.scala 63:156:@37129.4]
  wire [10:0] buffer_9_747; // @[Modules.scala 63:156:@37130.4]
  wire [11:0] _T_85552; // @[Modules.scala 63:156:@37132.4]
  wire [10:0] _T_85553; // @[Modules.scala 63:156:@37133.4]
  wire [10:0] buffer_9_748; // @[Modules.scala 63:156:@37134.4]
  wire [11:0] _T_85555; // @[Modules.scala 63:156:@37136.4]
  wire [10:0] _T_85556; // @[Modules.scala 63:156:@37137.4]
  wire [10:0] buffer_9_749; // @[Modules.scala 63:156:@37138.4]
  wire [11:0] _T_85558; // @[Modules.scala 63:156:@37140.4]
  wire [10:0] _T_85559; // @[Modules.scala 63:156:@37141.4]
  wire [10:0] buffer_9_750; // @[Modules.scala 63:156:@37142.4]
  wire [11:0] _T_85561; // @[Modules.scala 63:156:@37144.4]
  wire [10:0] _T_85562; // @[Modules.scala 63:156:@37145.4]
  wire [10:0] buffer_9_751; // @[Modules.scala 63:156:@37146.4]
  wire [11:0] _T_85564; // @[Modules.scala 63:156:@37148.4]
  wire [10:0] _T_85565; // @[Modules.scala 63:156:@37149.4]
  wire [10:0] buffer_9_752; // @[Modules.scala 63:156:@37150.4]
  wire [11:0] _T_85567; // @[Modules.scala 63:156:@37152.4]
  wire [10:0] _T_85568; // @[Modules.scala 63:156:@37153.4]
  wire [10:0] buffer_9_753; // @[Modules.scala 63:156:@37154.4]
  wire [11:0] _T_85570; // @[Modules.scala 63:156:@37156.4]
  wire [10:0] _T_85571; // @[Modules.scala 63:156:@37157.4]
  wire [10:0] buffer_9_754; // @[Modules.scala 63:156:@37158.4]
  wire [11:0] _T_85573; // @[Modules.scala 63:156:@37160.4]
  wire [10:0] _T_85574; // @[Modules.scala 63:156:@37161.4]
  wire [10:0] buffer_9_755; // @[Modules.scala 63:156:@37162.4]
  wire [11:0] _T_85576; // @[Modules.scala 63:156:@37164.4]
  wire [10:0] _T_85577; // @[Modules.scala 63:156:@37165.4]
  wire [10:0] buffer_9_756; // @[Modules.scala 63:156:@37166.4]
  wire [11:0] _T_85579; // @[Modules.scala 63:156:@37168.4]
  wire [10:0] _T_85580; // @[Modules.scala 63:156:@37169.4]
  wire [10:0] buffer_9_757; // @[Modules.scala 63:156:@37170.4]
  wire [11:0] _T_85582; // @[Modules.scala 63:156:@37172.4]
  wire [10:0] _T_85583; // @[Modules.scala 63:156:@37173.4]
  wire [10:0] buffer_9_758; // @[Modules.scala 63:156:@37174.4]
  wire [11:0] _T_85585; // @[Modules.scala 63:156:@37176.4]
  wire [10:0] _T_85586; // @[Modules.scala 63:156:@37177.4]
  wire [10:0] buffer_9_759; // @[Modules.scala 63:156:@37178.4]
  wire [11:0] _T_85588; // @[Modules.scala 63:156:@37180.4]
  wire [10:0] _T_85589; // @[Modules.scala 63:156:@37181.4]
  wire [10:0] buffer_9_760; // @[Modules.scala 63:156:@37182.4]
  wire [11:0] _T_85591; // @[Modules.scala 63:156:@37184.4]
  wire [10:0] _T_85592; // @[Modules.scala 63:156:@37185.4]
  wire [10:0] buffer_9_761; // @[Modules.scala 63:156:@37186.4]
  wire [11:0] _T_85594; // @[Modules.scala 63:156:@37188.4]
  wire [10:0] _T_85595; // @[Modules.scala 63:156:@37189.4]
  wire [10:0] buffer_9_762; // @[Modules.scala 63:156:@37190.4]
  wire [11:0] _T_85597; // @[Modules.scala 63:156:@37192.4]
  wire [10:0] _T_85598; // @[Modules.scala 63:156:@37193.4]
  wire [10:0] buffer_9_763; // @[Modules.scala 63:156:@37194.4]
  wire [11:0] _T_85600; // @[Modules.scala 63:156:@37196.4]
  wire [10:0] _T_85601; // @[Modules.scala 63:156:@37197.4]
  wire [10:0] buffer_9_764; // @[Modules.scala 63:156:@37198.4]
  wire [11:0] _T_85603; // @[Modules.scala 63:156:@37200.4]
  wire [10:0] _T_85604; // @[Modules.scala 63:156:@37201.4]
  wire [10:0] buffer_9_765; // @[Modules.scala 63:156:@37202.4]
  wire [11:0] _T_85606; // @[Modules.scala 63:156:@37204.4]
  wire [10:0] _T_85607; // @[Modules.scala 63:156:@37205.4]
  wire [10:0] buffer_9_766; // @[Modules.scala 63:156:@37206.4]
  wire [11:0] _T_85609; // @[Modules.scala 63:156:@37208.4]
  wire [10:0] _T_85610; // @[Modules.scala 63:156:@37209.4]
  wire [10:0] buffer_9_767; // @[Modules.scala 63:156:@37210.4]
  wire [11:0] _T_85612; // @[Modules.scala 63:156:@37212.4]
  wire [10:0] _T_85613; // @[Modules.scala 63:156:@37213.4]
  wire [10:0] buffer_9_768; // @[Modules.scala 63:156:@37214.4]
  wire [11:0] _T_85615; // @[Modules.scala 63:156:@37216.4]
  wire [10:0] _T_85616; // @[Modules.scala 63:156:@37217.4]
  wire [10:0] buffer_9_769; // @[Modules.scala 63:156:@37218.4]
  wire [11:0] _T_85618; // @[Modules.scala 63:156:@37220.4]
  wire [10:0] _T_85619; // @[Modules.scala 63:156:@37221.4]
  wire [10:0] buffer_9_770; // @[Modules.scala 63:156:@37222.4]
  wire [11:0] _T_85621; // @[Modules.scala 63:156:@37224.4]
  wire [10:0] _T_85622; // @[Modules.scala 63:156:@37225.4]
  wire [10:0] buffer_9_771; // @[Modules.scala 63:156:@37226.4]
  wire [11:0] _T_85624; // @[Modules.scala 63:156:@37228.4]
  wire [10:0] _T_85625; // @[Modules.scala 63:156:@37229.4]
  wire [10:0] buffer_9_772; // @[Modules.scala 63:156:@37230.4]
  wire [11:0] _T_85627; // @[Modules.scala 63:156:@37232.4]
  wire [10:0] _T_85628; // @[Modules.scala 63:156:@37233.4]
  wire [10:0] buffer_9_773; // @[Modules.scala 63:156:@37234.4]
  wire [11:0] _T_85630; // @[Modules.scala 63:156:@37236.4]
  wire [10:0] _T_85631; // @[Modules.scala 63:156:@37237.4]
  wire [10:0] buffer_9_774; // @[Modules.scala 63:156:@37238.4]
  wire [11:0] _T_85633; // @[Modules.scala 63:156:@37240.4]
  wire [10:0] _T_85634; // @[Modules.scala 63:156:@37241.4]
  wire [10:0] buffer_9_775; // @[Modules.scala 63:156:@37242.4]
  wire [11:0] _T_85636; // @[Modules.scala 63:156:@37244.4]
  wire [10:0] _T_85637; // @[Modules.scala 63:156:@37245.4]
  wire [10:0] buffer_9_776; // @[Modules.scala 63:156:@37246.4]
  wire [11:0] _T_85639; // @[Modules.scala 63:156:@37248.4]
  wire [10:0] _T_85640; // @[Modules.scala 63:156:@37249.4]
  wire [10:0] buffer_9_777; // @[Modules.scala 63:156:@37250.4]
  wire [11:0] _T_85642; // @[Modules.scala 63:156:@37252.4]
  wire [10:0] _T_85643; // @[Modules.scala 63:156:@37253.4]
  wire [10:0] buffer_9_778; // @[Modules.scala 63:156:@37254.4]
  wire [11:0] _T_85645; // @[Modules.scala 63:156:@37256.4]
  wire [10:0] _T_85646; // @[Modules.scala 63:156:@37257.4]
  wire [10:0] buffer_9_779; // @[Modules.scala 63:156:@37258.4]
  wire [11:0] _T_85648; // @[Modules.scala 63:156:@37260.4]
  wire [10:0] _T_85649; // @[Modules.scala 63:156:@37261.4]
  wire [10:0] buffer_9_780; // @[Modules.scala 63:156:@37262.4]
  wire [11:0] _T_85651; // @[Modules.scala 63:156:@37264.4]
  wire [10:0] _T_85652; // @[Modules.scala 63:156:@37265.4]
  wire [10:0] buffer_9_781; // @[Modules.scala 63:156:@37266.4]
  wire [11:0] _T_85654; // @[Modules.scala 63:156:@37268.4]
  wire [10:0] _T_85655; // @[Modules.scala 63:156:@37269.4]
  wire [10:0] buffer_9_782; // @[Modules.scala 63:156:@37270.4]
  wire [11:0] _T_85657; // @[Modules.scala 63:156:@37272.4]
  wire [10:0] _T_85658; // @[Modules.scala 63:156:@37273.4]
  wire [10:0] buffer_9_783; // @[Modules.scala 63:156:@37274.4]
  wire [5:0] _T_85880; // @[Modules.scala 37:46:@37540.4]
  wire [4:0] _T_85881; // @[Modules.scala 37:46:@37541.4]
  wire [4:0] _T_85882; // @[Modules.scala 37:46:@37542.4]
  wire [5:0] _T_85959; // @[Modules.scala 43:47:@37636.4]
  wire [4:0] _T_85960; // @[Modules.scala 43:47:@37637.4]
  wire [4:0] _T_85961; // @[Modules.scala 43:47:@37638.4]
  wire [5:0] _T_86000; // @[Modules.scala 40:46:@37686.4]
  wire [4:0] _T_86001; // @[Modules.scala 40:46:@37687.4]
  wire [4:0] _T_86002; // @[Modules.scala 40:46:@37688.4]
  wire [5:0] _T_86068; // @[Modules.scala 40:46:@37758.4]
  wire [4:0] _T_86069; // @[Modules.scala 40:46:@37759.4]
  wire [4:0] _T_86070; // @[Modules.scala 40:46:@37760.4]
  wire [5:0] _T_86165; // @[Modules.scala 40:46:@37864.4]
  wire [4:0] _T_86166; // @[Modules.scala 40:46:@37865.4]
  wire [4:0] _T_86167; // @[Modules.scala 40:46:@37866.4]
  wire [5:0] _T_86386; // @[Modules.scala 37:46:@38091.4]
  wire [4:0] _T_86387; // @[Modules.scala 37:46:@38092.4]
  wire [4:0] _T_86388; // @[Modules.scala 37:46:@38093.4]
  wire [5:0] _T_86607; // @[Modules.scala 43:47:@38325.4]
  wire [4:0] _T_86608; // @[Modules.scala 43:47:@38326.4]
  wire [4:0] _T_86609; // @[Modules.scala 43:47:@38327.4]
  wire [5:0] _T_86657; // @[Modules.scala 40:46:@38380.4]
  wire [4:0] _T_86658; // @[Modules.scala 40:46:@38381.4]
  wire [4:0] _T_86659; // @[Modules.scala 40:46:@38382.4]
  wire [5:0] _T_86774; // @[Modules.scala 43:47:@38515.4]
  wire [4:0] _T_86775; // @[Modules.scala 43:47:@38516.4]
  wire [4:0] _T_86776; // @[Modules.scala 43:47:@38517.4]
  wire [5:0] _T_86873; // @[Modules.scala 43:47:@38633.4]
  wire [4:0] _T_86874; // @[Modules.scala 43:47:@38634.4]
  wire [4:0] _T_86875; // @[Modules.scala 43:47:@38635.4]
  wire [5:0] _T_87126; // @[Modules.scala 40:46:@38933.4]
  wire [4:0] _T_87127; // @[Modules.scala 40:46:@38934.4]
  wire [4:0] _T_87128; // @[Modules.scala 40:46:@38935.4]
  wire [5:0] _T_87146; // @[Modules.scala 37:46:@38955.4]
  wire [4:0] _T_87147; // @[Modules.scala 37:46:@38956.4]
  wire [4:0] _T_87148; // @[Modules.scala 37:46:@38957.4]
  wire [5:0] _T_87291; // @[Modules.scala 40:46:@39118.4]
  wire [4:0] _T_87292; // @[Modules.scala 40:46:@39119.4]
  wire [4:0] _T_87293; // @[Modules.scala 40:46:@39120.4]
  wire [5:0] _T_87380; // @[Modules.scala 43:47:@39211.4]
  wire [4:0] _T_87381; // @[Modules.scala 43:47:@39212.4]
  wire [4:0] _T_87382; // @[Modules.scala 43:47:@39213.4]
  wire [11:0] _T_87495; // @[Modules.scala 50:57:@39341.4]
  wire [10:0] _T_87496; // @[Modules.scala 50:57:@39342.4]
  wire [10:0] buffer_10_393; // @[Modules.scala 50:57:@39343.4]
  wire [11:0] _T_87498; // @[Modules.scala 50:57:@39345.4]
  wire [10:0] _T_87499; // @[Modules.scala 50:57:@39346.4]
  wire [10:0] buffer_10_394; // @[Modules.scala 50:57:@39347.4]
  wire [11:0] _T_87510; // @[Modules.scala 50:57:@39361.4]
  wire [10:0] _T_87511; // @[Modules.scala 50:57:@39362.4]
  wire [10:0] buffer_10_398; // @[Modules.scala 50:57:@39363.4]
  wire [11:0] _T_87531; // @[Modules.scala 50:57:@39389.4]
  wire [10:0] _T_87532; // @[Modules.scala 50:57:@39390.4]
  wire [10:0] buffer_10_405; // @[Modules.scala 50:57:@39391.4]
  wire [11:0] _T_87537; // @[Modules.scala 50:57:@39397.4]
  wire [10:0] _T_87538; // @[Modules.scala 50:57:@39398.4]
  wire [10:0] buffer_10_407; // @[Modules.scala 50:57:@39399.4]
  wire [11:0] _T_87555; // @[Modules.scala 50:57:@39421.4]
  wire [10:0] _T_87556; // @[Modules.scala 50:57:@39422.4]
  wire [10:0] buffer_10_413; // @[Modules.scala 50:57:@39423.4]
  wire [11:0] _T_87573; // @[Modules.scala 50:57:@39445.4]
  wire [10:0] _T_87574; // @[Modules.scala 50:57:@39446.4]
  wire [10:0] buffer_10_419; // @[Modules.scala 50:57:@39447.4]
  wire [10:0] buffer_10_56; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87576; // @[Modules.scala 50:57:@39449.4]
  wire [10:0] _T_87577; // @[Modules.scala 50:57:@39450.4]
  wire [10:0] buffer_10_420; // @[Modules.scala 50:57:@39451.4]
  wire [11:0] _T_87588; // @[Modules.scala 50:57:@39465.4]
  wire [10:0] _T_87589; // @[Modules.scala 50:57:@39466.4]
  wire [10:0] buffer_10_424; // @[Modules.scala 50:57:@39467.4]
  wire [11:0] _T_87594; // @[Modules.scala 50:57:@39473.4]
  wire [10:0] _T_87595; // @[Modules.scala 50:57:@39474.4]
  wire [10:0] buffer_10_426; // @[Modules.scala 50:57:@39475.4]
  wire [11:0] _T_87597; // @[Modules.scala 50:57:@39477.4]
  wire [10:0] _T_87598; // @[Modules.scala 50:57:@39478.4]
  wire [10:0] buffer_10_427; // @[Modules.scala 50:57:@39479.4]
  wire [11:0] _T_87603; // @[Modules.scala 50:57:@39485.4]
  wire [10:0] _T_87604; // @[Modules.scala 50:57:@39486.4]
  wire [10:0] buffer_10_429; // @[Modules.scala 50:57:@39487.4]
  wire [10:0] buffer_10_77; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87606; // @[Modules.scala 50:57:@39489.4]
  wire [10:0] _T_87607; // @[Modules.scala 50:57:@39490.4]
  wire [10:0] buffer_10_430; // @[Modules.scala 50:57:@39491.4]
  wire [11:0] _T_87609; // @[Modules.scala 50:57:@39493.4]
  wire [10:0] _T_87610; // @[Modules.scala 50:57:@39494.4]
  wire [10:0] buffer_10_431; // @[Modules.scala 50:57:@39495.4]
  wire [11:0] _T_87612; // @[Modules.scala 50:57:@39497.4]
  wire [10:0] _T_87613; // @[Modules.scala 50:57:@39498.4]
  wire [10:0] buffer_10_432; // @[Modules.scala 50:57:@39499.4]
  wire [11:0] _T_87615; // @[Modules.scala 50:57:@39501.4]
  wire [10:0] _T_87616; // @[Modules.scala 50:57:@39502.4]
  wire [10:0] buffer_10_433; // @[Modules.scala 50:57:@39503.4]
  wire [11:0] _T_87618; // @[Modules.scala 50:57:@39505.4]
  wire [10:0] _T_87619; // @[Modules.scala 50:57:@39506.4]
  wire [10:0] buffer_10_434; // @[Modules.scala 50:57:@39507.4]
  wire [11:0] _T_87621; // @[Modules.scala 50:57:@39509.4]
  wire [10:0] _T_87622; // @[Modules.scala 50:57:@39510.4]
  wire [10:0] buffer_10_435; // @[Modules.scala 50:57:@39511.4]
  wire [10:0] buffer_10_88; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87624; // @[Modules.scala 50:57:@39513.4]
  wire [10:0] _T_87625; // @[Modules.scala 50:57:@39514.4]
  wire [10:0] buffer_10_436; // @[Modules.scala 50:57:@39515.4]
  wire [11:0] _T_87636; // @[Modules.scala 50:57:@39529.4]
  wire [10:0] _T_87637; // @[Modules.scala 50:57:@39530.4]
  wire [10:0] buffer_10_440; // @[Modules.scala 50:57:@39531.4]
  wire [10:0] buffer_10_100; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87642; // @[Modules.scala 50:57:@39537.4]
  wire [10:0] _T_87643; // @[Modules.scala 50:57:@39538.4]
  wire [10:0] buffer_10_442; // @[Modules.scala 50:57:@39539.4]
  wire [11:0] _T_87645; // @[Modules.scala 50:57:@39541.4]
  wire [10:0] _T_87646; // @[Modules.scala 50:57:@39542.4]
  wire [10:0] buffer_10_443; // @[Modules.scala 50:57:@39543.4]
  wire [11:0] _T_87648; // @[Modules.scala 50:57:@39545.4]
  wire [10:0] _T_87649; // @[Modules.scala 50:57:@39546.4]
  wire [10:0] buffer_10_444; // @[Modules.scala 50:57:@39547.4]
  wire [11:0] _T_87663; // @[Modules.scala 50:57:@39565.4]
  wire [10:0] _T_87664; // @[Modules.scala 50:57:@39566.4]
  wire [10:0] buffer_10_449; // @[Modules.scala 50:57:@39567.4]
  wire [10:0] buffer_10_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87669; // @[Modules.scala 50:57:@39573.4]
  wire [10:0] _T_87670; // @[Modules.scala 50:57:@39574.4]
  wire [10:0] buffer_10_451; // @[Modules.scala 50:57:@39575.4]
  wire [10:0] buffer_10_154; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87723; // @[Modules.scala 50:57:@39645.4]
  wire [10:0] _T_87724; // @[Modules.scala 50:57:@39646.4]
  wire [10:0] buffer_10_469; // @[Modules.scala 50:57:@39647.4]
  wire [11:0] _T_87735; // @[Modules.scala 50:57:@39661.4]
  wire [10:0] _T_87736; // @[Modules.scala 50:57:@39662.4]
  wire [10:0] buffer_10_473; // @[Modules.scala 50:57:@39663.4]
  wire [11:0] _T_87741; // @[Modules.scala 50:57:@39669.4]
  wire [10:0] _T_87742; // @[Modules.scala 50:57:@39670.4]
  wire [10:0] buffer_10_475; // @[Modules.scala 50:57:@39671.4]
  wire [11:0] _T_87756; // @[Modules.scala 50:57:@39689.4]
  wire [10:0] _T_87757; // @[Modules.scala 50:57:@39690.4]
  wire [10:0] buffer_10_480; // @[Modules.scala 50:57:@39691.4]
  wire [11:0] _T_87777; // @[Modules.scala 50:57:@39717.4]
  wire [10:0] _T_87778; // @[Modules.scala 50:57:@39718.4]
  wire [10:0] buffer_10_487; // @[Modules.scala 50:57:@39719.4]
  wire [10:0] buffer_10_193; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87780; // @[Modules.scala 50:57:@39721.4]
  wire [10:0] _T_87781; // @[Modules.scala 50:57:@39722.4]
  wire [10:0] buffer_10_488; // @[Modules.scala 50:57:@39723.4]
  wire [10:0] buffer_10_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87795; // @[Modules.scala 50:57:@39741.4]
  wire [10:0] _T_87796; // @[Modules.scala 50:57:@39742.4]
  wire [10:0] buffer_10_493; // @[Modules.scala 50:57:@39743.4]
  wire [11:0] _T_87801; // @[Modules.scala 50:57:@39749.4]
  wire [10:0] _T_87802; // @[Modules.scala 50:57:@39750.4]
  wire [10:0] buffer_10_495; // @[Modules.scala 50:57:@39751.4]
  wire [11:0] _T_87804; // @[Modules.scala 50:57:@39753.4]
  wire [10:0] _T_87805; // @[Modules.scala 50:57:@39754.4]
  wire [10:0] buffer_10_496; // @[Modules.scala 50:57:@39755.4]
  wire [11:0] _T_87822; // @[Modules.scala 50:57:@39777.4]
  wire [10:0] _T_87823; // @[Modules.scala 50:57:@39778.4]
  wire [10:0] buffer_10_502; // @[Modules.scala 50:57:@39779.4]
  wire [11:0] _T_87831; // @[Modules.scala 50:57:@39789.4]
  wire [10:0] _T_87832; // @[Modules.scala 50:57:@39790.4]
  wire [10:0] buffer_10_505; // @[Modules.scala 50:57:@39791.4]
  wire [10:0] buffer_10_230; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87837; // @[Modules.scala 50:57:@39797.4]
  wire [10:0] _T_87838; // @[Modules.scala 50:57:@39798.4]
  wire [10:0] buffer_10_507; // @[Modules.scala 50:57:@39799.4]
  wire [11:0] _T_87843; // @[Modules.scala 50:57:@39805.4]
  wire [10:0] _T_87844; // @[Modules.scala 50:57:@39806.4]
  wire [10:0] buffer_10_509; // @[Modules.scala 50:57:@39807.4]
  wire [11:0] _T_87858; // @[Modules.scala 50:57:@39825.4]
  wire [10:0] _T_87859; // @[Modules.scala 50:57:@39826.4]
  wire [10:0] buffer_10_514; // @[Modules.scala 50:57:@39827.4]
  wire [11:0] _T_87861; // @[Modules.scala 50:57:@39829.4]
  wire [10:0] _T_87862; // @[Modules.scala 50:57:@39830.4]
  wire [10:0] buffer_10_515; // @[Modules.scala 50:57:@39831.4]
  wire [10:0] buffer_10_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87873; // @[Modules.scala 50:57:@39845.4]
  wire [10:0] _T_87874; // @[Modules.scala 50:57:@39846.4]
  wire [10:0] buffer_10_519; // @[Modules.scala 50:57:@39847.4]
  wire [11:0] _T_87876; // @[Modules.scala 50:57:@39849.4]
  wire [10:0] _T_87877; // @[Modules.scala 50:57:@39850.4]
  wire [10:0] buffer_10_520; // @[Modules.scala 50:57:@39851.4]
  wire [11:0] _T_87879; // @[Modules.scala 50:57:@39853.4]
  wire [10:0] _T_87880; // @[Modules.scala 50:57:@39854.4]
  wire [10:0] buffer_10_521; // @[Modules.scala 50:57:@39855.4]
  wire [11:0] _T_87897; // @[Modules.scala 50:57:@39877.4]
  wire [10:0] _T_87898; // @[Modules.scala 50:57:@39878.4]
  wire [10:0] buffer_10_527; // @[Modules.scala 50:57:@39879.4]
  wire [11:0] _T_87918; // @[Modules.scala 50:57:@39905.4]
  wire [10:0] _T_87919; // @[Modules.scala 50:57:@39906.4]
  wire [10:0] buffer_10_534; // @[Modules.scala 50:57:@39907.4]
  wire [11:0] _T_87927; // @[Modules.scala 50:57:@39917.4]
  wire [10:0] _T_87928; // @[Modules.scala 50:57:@39918.4]
  wire [10:0] buffer_10_537; // @[Modules.scala 50:57:@39919.4]
  wire [11:0] _T_87948; // @[Modules.scala 50:57:@39945.4]
  wire [10:0] _T_87949; // @[Modules.scala 50:57:@39946.4]
  wire [10:0] buffer_10_544; // @[Modules.scala 50:57:@39947.4]
  wire [11:0] _T_87951; // @[Modules.scala 50:57:@39949.4]
  wire [10:0] _T_87952; // @[Modules.scala 50:57:@39950.4]
  wire [10:0] buffer_10_545; // @[Modules.scala 50:57:@39951.4]
  wire [10:0] buffer_10_318; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87969; // @[Modules.scala 50:57:@39973.4]
  wire [10:0] _T_87970; // @[Modules.scala 50:57:@39974.4]
  wire [10:0] buffer_10_551; // @[Modules.scala 50:57:@39975.4]
  wire [11:0] _T_87972; // @[Modules.scala 50:57:@39977.4]
  wire [10:0] _T_87973; // @[Modules.scala 50:57:@39978.4]
  wire [10:0] buffer_10_552; // @[Modules.scala 50:57:@39979.4]
  wire [10:0] buffer_10_322; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_87975; // @[Modules.scala 50:57:@39981.4]
  wire [10:0] _T_87976; // @[Modules.scala 50:57:@39982.4]
  wire [10:0] buffer_10_553; // @[Modules.scala 50:57:@39983.4]
  wire [11:0] _T_87981; // @[Modules.scala 50:57:@39989.4]
  wire [10:0] _T_87982; // @[Modules.scala 50:57:@39990.4]
  wire [10:0] buffer_10_555; // @[Modules.scala 50:57:@39991.4]
  wire [11:0] _T_88005; // @[Modules.scala 50:57:@40021.4]
  wire [10:0] _T_88006; // @[Modules.scala 50:57:@40022.4]
  wire [10:0] buffer_10_563; // @[Modules.scala 50:57:@40023.4]
  wire [10:0] buffer_10_353; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_88020; // @[Modules.scala 50:57:@40041.4]
  wire [10:0] _T_88021; // @[Modules.scala 50:57:@40042.4]
  wire [10:0] buffer_10_568; // @[Modules.scala 50:57:@40043.4]
  wire [10:0] buffer_10_368; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_88044; // @[Modules.scala 50:57:@40073.4]
  wire [10:0] _T_88045; // @[Modules.scala 50:57:@40074.4]
  wire [10:0] buffer_10_576; // @[Modules.scala 50:57:@40075.4]
  wire [11:0] _T_88056; // @[Modules.scala 50:57:@40089.4]
  wire [10:0] _T_88057; // @[Modules.scala 50:57:@40090.4]
  wire [10:0] buffer_10_580; // @[Modules.scala 50:57:@40091.4]
  wire [11:0] _T_88059; // @[Modules.scala 50:57:@40093.4]
  wire [10:0] _T_88060; // @[Modules.scala 50:57:@40094.4]
  wire [10:0] buffer_10_581; // @[Modules.scala 50:57:@40095.4]
  wire [11:0] _T_88062; // @[Modules.scala 50:57:@40097.4]
  wire [10:0] _T_88063; // @[Modules.scala 50:57:@40098.4]
  wire [10:0] buffer_10_582; // @[Modules.scala 50:57:@40099.4]
  wire [11:0] _T_88077; // @[Modules.scala 50:57:@40117.4]
  wire [10:0] _T_88078; // @[Modules.scala 50:57:@40118.4]
  wire [10:0] buffer_10_587; // @[Modules.scala 50:57:@40119.4]
  wire [11:0] _T_88080; // @[Modules.scala 53:83:@40121.4]
  wire [10:0] _T_88081; // @[Modules.scala 53:83:@40122.4]
  wire [10:0] buffer_10_588; // @[Modules.scala 53:83:@40123.4]
  wire [11:0] _T_88083; // @[Modules.scala 53:83:@40125.4]
  wire [10:0] _T_88084; // @[Modules.scala 53:83:@40126.4]
  wire [10:0] buffer_10_589; // @[Modules.scala 53:83:@40127.4]
  wire [11:0] _T_88089; // @[Modules.scala 53:83:@40133.4]
  wire [10:0] _T_88090; // @[Modules.scala 53:83:@40134.4]
  wire [10:0] buffer_10_591; // @[Modules.scala 53:83:@40135.4]
  wire [11:0] _T_88098; // @[Modules.scala 53:83:@40145.4]
  wire [10:0] _T_88099; // @[Modules.scala 53:83:@40146.4]
  wire [10:0] buffer_10_594; // @[Modules.scala 53:83:@40147.4]
  wire [11:0] _T_88101; // @[Modules.scala 53:83:@40149.4]
  wire [10:0] _T_88102; // @[Modules.scala 53:83:@40150.4]
  wire [10:0] buffer_10_595; // @[Modules.scala 53:83:@40151.4]
  wire [11:0] _T_88110; // @[Modules.scala 53:83:@40161.4]
  wire [10:0] _T_88111; // @[Modules.scala 53:83:@40162.4]
  wire [10:0] buffer_10_598; // @[Modules.scala 53:83:@40163.4]
  wire [11:0] _T_88119; // @[Modules.scala 53:83:@40173.4]
  wire [10:0] _T_88120; // @[Modules.scala 53:83:@40174.4]
  wire [10:0] buffer_10_601; // @[Modules.scala 53:83:@40175.4]
  wire [11:0] _T_88122; // @[Modules.scala 53:83:@40177.4]
  wire [10:0] _T_88123; // @[Modules.scala 53:83:@40178.4]
  wire [10:0] buffer_10_602; // @[Modules.scala 53:83:@40179.4]
  wire [11:0] _T_88125; // @[Modules.scala 53:83:@40181.4]
  wire [10:0] _T_88126; // @[Modules.scala 53:83:@40182.4]
  wire [10:0] buffer_10_603; // @[Modules.scala 53:83:@40183.4]
  wire [11:0] _T_88128; // @[Modules.scala 53:83:@40185.4]
  wire [10:0] _T_88129; // @[Modules.scala 53:83:@40186.4]
  wire [10:0] buffer_10_604; // @[Modules.scala 53:83:@40187.4]
  wire [11:0] _T_88131; // @[Modules.scala 53:83:@40189.4]
  wire [10:0] _T_88132; // @[Modules.scala 53:83:@40190.4]
  wire [10:0] buffer_10_605; // @[Modules.scala 53:83:@40191.4]
  wire [11:0] _T_88134; // @[Modules.scala 53:83:@40193.4]
  wire [10:0] _T_88135; // @[Modules.scala 53:83:@40194.4]
  wire [10:0] buffer_10_606; // @[Modules.scala 53:83:@40195.4]
  wire [11:0] _T_88137; // @[Modules.scala 53:83:@40197.4]
  wire [10:0] _T_88138; // @[Modules.scala 53:83:@40198.4]
  wire [10:0] buffer_10_607; // @[Modules.scala 53:83:@40199.4]
  wire [11:0] _T_88140; // @[Modules.scala 53:83:@40201.4]
  wire [10:0] _T_88141; // @[Modules.scala 53:83:@40202.4]
  wire [10:0] buffer_10_608; // @[Modules.scala 53:83:@40203.4]
  wire [11:0] _T_88143; // @[Modules.scala 53:83:@40205.4]
  wire [10:0] _T_88144; // @[Modules.scala 53:83:@40206.4]
  wire [10:0] buffer_10_609; // @[Modules.scala 53:83:@40207.4]
  wire [11:0] _T_88146; // @[Modules.scala 53:83:@40209.4]
  wire [10:0] _T_88147; // @[Modules.scala 53:83:@40210.4]
  wire [10:0] buffer_10_610; // @[Modules.scala 53:83:@40211.4]
  wire [11:0] _T_88149; // @[Modules.scala 53:83:@40213.4]
  wire [10:0] _T_88150; // @[Modules.scala 53:83:@40214.4]
  wire [10:0] buffer_10_611; // @[Modules.scala 53:83:@40215.4]
  wire [11:0] _T_88152; // @[Modules.scala 53:83:@40217.4]
  wire [10:0] _T_88153; // @[Modules.scala 53:83:@40218.4]
  wire [10:0] buffer_10_612; // @[Modules.scala 53:83:@40219.4]
  wire [11:0] _T_88155; // @[Modules.scala 53:83:@40221.4]
  wire [10:0] _T_88156; // @[Modules.scala 53:83:@40222.4]
  wire [10:0] buffer_10_613; // @[Modules.scala 53:83:@40223.4]
  wire [11:0] _T_88158; // @[Modules.scala 53:83:@40225.4]
  wire [10:0] _T_88159; // @[Modules.scala 53:83:@40226.4]
  wire [10:0] buffer_10_614; // @[Modules.scala 53:83:@40227.4]
  wire [11:0] _T_88161; // @[Modules.scala 53:83:@40229.4]
  wire [10:0] _T_88162; // @[Modules.scala 53:83:@40230.4]
  wire [10:0] buffer_10_615; // @[Modules.scala 53:83:@40231.4]
  wire [11:0] _T_88164; // @[Modules.scala 53:83:@40233.4]
  wire [10:0] _T_88165; // @[Modules.scala 53:83:@40234.4]
  wire [10:0] buffer_10_616; // @[Modules.scala 53:83:@40235.4]
  wire [11:0] _T_88167; // @[Modules.scala 53:83:@40237.4]
  wire [10:0] _T_88168; // @[Modules.scala 53:83:@40238.4]
  wire [10:0] buffer_10_617; // @[Modules.scala 53:83:@40239.4]
  wire [11:0] _T_88173; // @[Modules.scala 53:83:@40245.4]
  wire [10:0] _T_88174; // @[Modules.scala 53:83:@40246.4]
  wire [10:0] buffer_10_619; // @[Modules.scala 53:83:@40247.4]
  wire [11:0] _T_88176; // @[Modules.scala 53:83:@40249.4]
  wire [10:0] _T_88177; // @[Modules.scala 53:83:@40250.4]
  wire [10:0] buffer_10_620; // @[Modules.scala 53:83:@40251.4]
  wire [11:0] _T_88185; // @[Modules.scala 53:83:@40261.4]
  wire [10:0] _T_88186; // @[Modules.scala 53:83:@40262.4]
  wire [10:0] buffer_10_623; // @[Modules.scala 53:83:@40263.4]
  wire [11:0] _T_88194; // @[Modules.scala 53:83:@40273.4]
  wire [10:0] _T_88195; // @[Modules.scala 53:83:@40274.4]
  wire [10:0] buffer_10_626; // @[Modules.scala 53:83:@40275.4]
  wire [11:0] _T_88200; // @[Modules.scala 53:83:@40281.4]
  wire [10:0] _T_88201; // @[Modules.scala 53:83:@40282.4]
  wire [10:0] buffer_10_628; // @[Modules.scala 53:83:@40283.4]
  wire [11:0] _T_88203; // @[Modules.scala 53:83:@40285.4]
  wire [10:0] _T_88204; // @[Modules.scala 53:83:@40286.4]
  wire [10:0] buffer_10_629; // @[Modules.scala 53:83:@40287.4]
  wire [11:0] _T_88212; // @[Modules.scala 53:83:@40297.4]
  wire [10:0] _T_88213; // @[Modules.scala 53:83:@40298.4]
  wire [10:0] buffer_10_632; // @[Modules.scala 53:83:@40299.4]
  wire [11:0] _T_88215; // @[Modules.scala 53:83:@40301.4]
  wire [10:0] _T_88216; // @[Modules.scala 53:83:@40302.4]
  wire [10:0] buffer_10_633; // @[Modules.scala 53:83:@40303.4]
  wire [11:0] _T_88221; // @[Modules.scala 53:83:@40309.4]
  wire [10:0] _T_88222; // @[Modules.scala 53:83:@40310.4]
  wire [10:0] buffer_10_635; // @[Modules.scala 53:83:@40311.4]
  wire [11:0] _T_88224; // @[Modules.scala 53:83:@40313.4]
  wire [10:0] _T_88225; // @[Modules.scala 53:83:@40314.4]
  wire [10:0] buffer_10_636; // @[Modules.scala 53:83:@40315.4]
  wire [11:0] _T_88227; // @[Modules.scala 53:83:@40317.4]
  wire [10:0] _T_88228; // @[Modules.scala 53:83:@40318.4]
  wire [10:0] buffer_10_637; // @[Modules.scala 53:83:@40319.4]
  wire [11:0] _T_88230; // @[Modules.scala 53:83:@40321.4]
  wire [10:0] _T_88231; // @[Modules.scala 53:83:@40322.4]
  wire [10:0] buffer_10_638; // @[Modules.scala 53:83:@40323.4]
  wire [11:0] _T_88233; // @[Modules.scala 53:83:@40325.4]
  wire [10:0] _T_88234; // @[Modules.scala 53:83:@40326.4]
  wire [10:0] buffer_10_639; // @[Modules.scala 53:83:@40327.4]
  wire [11:0] _T_88236; // @[Modules.scala 53:83:@40329.4]
  wire [10:0] _T_88237; // @[Modules.scala 53:83:@40330.4]
  wire [10:0] buffer_10_640; // @[Modules.scala 53:83:@40331.4]
  wire [11:0] _T_88239; // @[Modules.scala 53:83:@40333.4]
  wire [10:0] _T_88240; // @[Modules.scala 53:83:@40334.4]
  wire [10:0] buffer_10_641; // @[Modules.scala 53:83:@40335.4]
  wire [11:0] _T_88242; // @[Modules.scala 53:83:@40337.4]
  wire [10:0] _T_88243; // @[Modules.scala 53:83:@40338.4]
  wire [10:0] buffer_10_642; // @[Modules.scala 53:83:@40339.4]
  wire [11:0] _T_88245; // @[Modules.scala 53:83:@40341.4]
  wire [10:0] _T_88246; // @[Modules.scala 53:83:@40342.4]
  wire [10:0] buffer_10_643; // @[Modules.scala 53:83:@40343.4]
  wire [11:0] _T_88248; // @[Modules.scala 53:83:@40345.4]
  wire [10:0] _T_88249; // @[Modules.scala 53:83:@40346.4]
  wire [10:0] buffer_10_644; // @[Modules.scala 53:83:@40347.4]
  wire [11:0] _T_88251; // @[Modules.scala 53:83:@40349.4]
  wire [10:0] _T_88252; // @[Modules.scala 53:83:@40350.4]
  wire [10:0] buffer_10_645; // @[Modules.scala 53:83:@40351.4]
  wire [11:0] _T_88254; // @[Modules.scala 53:83:@40353.4]
  wire [10:0] _T_88255; // @[Modules.scala 53:83:@40354.4]
  wire [10:0] buffer_10_646; // @[Modules.scala 53:83:@40355.4]
  wire [11:0] _T_88260; // @[Modules.scala 53:83:@40361.4]
  wire [10:0] _T_88261; // @[Modules.scala 53:83:@40362.4]
  wire [10:0] buffer_10_648; // @[Modules.scala 53:83:@40363.4]
  wire [11:0] _T_88263; // @[Modules.scala 53:83:@40365.4]
  wire [10:0] _T_88264; // @[Modules.scala 53:83:@40366.4]
  wire [10:0] buffer_10_649; // @[Modules.scala 53:83:@40367.4]
  wire [11:0] _T_88269; // @[Modules.scala 53:83:@40373.4]
  wire [10:0] _T_88270; // @[Modules.scala 53:83:@40374.4]
  wire [10:0] buffer_10_651; // @[Modules.scala 53:83:@40375.4]
  wire [11:0] _T_88272; // @[Modules.scala 53:83:@40377.4]
  wire [10:0] _T_88273; // @[Modules.scala 53:83:@40378.4]
  wire [10:0] buffer_10_652; // @[Modules.scala 53:83:@40379.4]
  wire [11:0] _T_88275; // @[Modules.scala 53:83:@40381.4]
  wire [10:0] _T_88276; // @[Modules.scala 53:83:@40382.4]
  wire [10:0] buffer_10_653; // @[Modules.scala 53:83:@40383.4]
  wire [11:0] _T_88281; // @[Modules.scala 53:83:@40389.4]
  wire [10:0] _T_88282; // @[Modules.scala 53:83:@40390.4]
  wire [10:0] buffer_10_655; // @[Modules.scala 53:83:@40391.4]
  wire [11:0] _T_88284; // @[Modules.scala 53:83:@40393.4]
  wire [10:0] _T_88285; // @[Modules.scala 53:83:@40394.4]
  wire [10:0] buffer_10_656; // @[Modules.scala 53:83:@40395.4]
  wire [11:0] _T_88287; // @[Modules.scala 53:83:@40397.4]
  wire [10:0] _T_88288; // @[Modules.scala 53:83:@40398.4]
  wire [10:0] buffer_10_657; // @[Modules.scala 53:83:@40399.4]
  wire [11:0] _T_88290; // @[Modules.scala 53:83:@40401.4]
  wire [10:0] _T_88291; // @[Modules.scala 53:83:@40402.4]
  wire [10:0] buffer_10_658; // @[Modules.scala 53:83:@40403.4]
  wire [11:0] _T_88293; // @[Modules.scala 53:83:@40405.4]
  wire [10:0] _T_88294; // @[Modules.scala 53:83:@40406.4]
  wire [10:0] buffer_10_659; // @[Modules.scala 53:83:@40407.4]
  wire [11:0] _T_88296; // @[Modules.scala 53:83:@40409.4]
  wire [10:0] _T_88297; // @[Modules.scala 53:83:@40410.4]
  wire [10:0] buffer_10_660; // @[Modules.scala 53:83:@40411.4]
  wire [11:0] _T_88308; // @[Modules.scala 53:83:@40425.4]
  wire [10:0] _T_88309; // @[Modules.scala 53:83:@40426.4]
  wire [10:0] buffer_10_664; // @[Modules.scala 53:83:@40427.4]
  wire [11:0] _T_88314; // @[Modules.scala 53:83:@40433.4]
  wire [10:0] _T_88315; // @[Modules.scala 53:83:@40434.4]
  wire [10:0] buffer_10_666; // @[Modules.scala 53:83:@40435.4]
  wire [11:0] _T_88317; // @[Modules.scala 53:83:@40437.4]
  wire [10:0] _T_88318; // @[Modules.scala 53:83:@40438.4]
  wire [10:0] buffer_10_667; // @[Modules.scala 53:83:@40439.4]
  wire [11:0] _T_88320; // @[Modules.scala 53:83:@40441.4]
  wire [10:0] _T_88321; // @[Modules.scala 53:83:@40442.4]
  wire [10:0] buffer_10_668; // @[Modules.scala 53:83:@40443.4]
  wire [11:0] _T_88323; // @[Modules.scala 53:83:@40445.4]
  wire [10:0] _T_88324; // @[Modules.scala 53:83:@40446.4]
  wire [10:0] buffer_10_669; // @[Modules.scala 53:83:@40447.4]
  wire [11:0] _T_88335; // @[Modules.scala 53:83:@40461.4]
  wire [10:0] _T_88336; // @[Modules.scala 53:83:@40462.4]
  wire [10:0] buffer_10_673; // @[Modules.scala 53:83:@40463.4]
  wire [11:0] _T_88344; // @[Modules.scala 53:83:@40473.4]
  wire [10:0] _T_88345; // @[Modules.scala 53:83:@40474.4]
  wire [10:0] buffer_10_676; // @[Modules.scala 53:83:@40475.4]
  wire [11:0] _T_88350; // @[Modules.scala 53:83:@40481.4]
  wire [10:0] _T_88351; // @[Modules.scala 53:83:@40482.4]
  wire [10:0] buffer_10_678; // @[Modules.scala 53:83:@40483.4]
  wire [11:0] _T_88353; // @[Modules.scala 53:83:@40485.4]
  wire [10:0] _T_88354; // @[Modules.scala 53:83:@40486.4]
  wire [10:0] buffer_10_679; // @[Modules.scala 53:83:@40487.4]
  wire [11:0] _T_88356; // @[Modules.scala 53:83:@40489.4]
  wire [10:0] _T_88357; // @[Modules.scala 53:83:@40490.4]
  wire [10:0] buffer_10_680; // @[Modules.scala 53:83:@40491.4]
  wire [11:0] _T_88362; // @[Modules.scala 53:83:@40497.4]
  wire [10:0] _T_88363; // @[Modules.scala 53:83:@40498.4]
  wire [10:0] buffer_10_682; // @[Modules.scala 53:83:@40499.4]
  wire [11:0] _T_88365; // @[Modules.scala 53:83:@40501.4]
  wire [10:0] _T_88366; // @[Modules.scala 53:83:@40502.4]
  wire [10:0] buffer_10_683; // @[Modules.scala 53:83:@40503.4]
  wire [11:0] _T_88371; // @[Modules.scala 53:83:@40509.4]
  wire [10:0] _T_88372; // @[Modules.scala 53:83:@40510.4]
  wire [10:0] buffer_10_685; // @[Modules.scala 53:83:@40511.4]
  wire [11:0] _T_88374; // @[Modules.scala 56:109:@40513.4]
  wire [10:0] _T_88375; // @[Modules.scala 56:109:@40514.4]
  wire [10:0] buffer_10_686; // @[Modules.scala 56:109:@40515.4]
  wire [11:0] _T_88377; // @[Modules.scala 56:109:@40517.4]
  wire [10:0] _T_88378; // @[Modules.scala 56:109:@40518.4]
  wire [10:0] buffer_10_687; // @[Modules.scala 56:109:@40519.4]
  wire [11:0] _T_88383; // @[Modules.scala 56:109:@40525.4]
  wire [10:0] _T_88384; // @[Modules.scala 56:109:@40526.4]
  wire [10:0] buffer_10_689; // @[Modules.scala 56:109:@40527.4]
  wire [11:0] _T_88389; // @[Modules.scala 56:109:@40533.4]
  wire [10:0] _T_88390; // @[Modules.scala 56:109:@40534.4]
  wire [10:0] buffer_10_691; // @[Modules.scala 56:109:@40535.4]
  wire [11:0] _T_88392; // @[Modules.scala 56:109:@40537.4]
  wire [10:0] _T_88393; // @[Modules.scala 56:109:@40538.4]
  wire [10:0] buffer_10_692; // @[Modules.scala 56:109:@40539.4]
  wire [11:0] _T_88395; // @[Modules.scala 56:109:@40541.4]
  wire [10:0] _T_88396; // @[Modules.scala 56:109:@40542.4]
  wire [10:0] buffer_10_693; // @[Modules.scala 56:109:@40543.4]
  wire [11:0] _T_88398; // @[Modules.scala 56:109:@40545.4]
  wire [10:0] _T_88399; // @[Modules.scala 56:109:@40546.4]
  wire [10:0] buffer_10_694; // @[Modules.scala 56:109:@40547.4]
  wire [11:0] _T_88401; // @[Modules.scala 56:109:@40549.4]
  wire [10:0] _T_88402; // @[Modules.scala 56:109:@40550.4]
  wire [10:0] buffer_10_695; // @[Modules.scala 56:109:@40551.4]
  wire [11:0] _T_88404; // @[Modules.scala 56:109:@40553.4]
  wire [10:0] _T_88405; // @[Modules.scala 56:109:@40554.4]
  wire [10:0] buffer_10_696; // @[Modules.scala 56:109:@40555.4]
  wire [11:0] _T_88407; // @[Modules.scala 56:109:@40557.4]
  wire [10:0] _T_88408; // @[Modules.scala 56:109:@40558.4]
  wire [10:0] buffer_10_697; // @[Modules.scala 56:109:@40559.4]
  wire [11:0] _T_88410; // @[Modules.scala 56:109:@40561.4]
  wire [10:0] _T_88411; // @[Modules.scala 56:109:@40562.4]
  wire [10:0] buffer_10_698; // @[Modules.scala 56:109:@40563.4]
  wire [11:0] _T_88413; // @[Modules.scala 56:109:@40565.4]
  wire [10:0] _T_88414; // @[Modules.scala 56:109:@40566.4]
  wire [10:0] buffer_10_699; // @[Modules.scala 56:109:@40567.4]
  wire [11:0] _T_88416; // @[Modules.scala 56:109:@40569.4]
  wire [10:0] _T_88417; // @[Modules.scala 56:109:@40570.4]
  wire [10:0] buffer_10_700; // @[Modules.scala 56:109:@40571.4]
  wire [11:0] _T_88419; // @[Modules.scala 56:109:@40573.4]
  wire [10:0] _T_88420; // @[Modules.scala 56:109:@40574.4]
  wire [10:0] buffer_10_701; // @[Modules.scala 56:109:@40575.4]
  wire [11:0] _T_88422; // @[Modules.scala 56:109:@40577.4]
  wire [10:0] _T_88423; // @[Modules.scala 56:109:@40578.4]
  wire [10:0] buffer_10_702; // @[Modules.scala 56:109:@40579.4]
  wire [11:0] _T_88425; // @[Modules.scala 56:109:@40581.4]
  wire [10:0] _T_88426; // @[Modules.scala 56:109:@40582.4]
  wire [10:0] buffer_10_703; // @[Modules.scala 56:109:@40583.4]
  wire [11:0] _T_88428; // @[Modules.scala 56:109:@40585.4]
  wire [10:0] _T_88429; // @[Modules.scala 56:109:@40586.4]
  wire [10:0] buffer_10_704; // @[Modules.scala 56:109:@40587.4]
  wire [11:0] _T_88431; // @[Modules.scala 56:109:@40589.4]
  wire [10:0] _T_88432; // @[Modules.scala 56:109:@40590.4]
  wire [10:0] buffer_10_705; // @[Modules.scala 56:109:@40591.4]
  wire [11:0] _T_88434; // @[Modules.scala 56:109:@40593.4]
  wire [10:0] _T_88435; // @[Modules.scala 56:109:@40594.4]
  wire [10:0] buffer_10_706; // @[Modules.scala 56:109:@40595.4]
  wire [11:0] _T_88440; // @[Modules.scala 56:109:@40601.4]
  wire [10:0] _T_88441; // @[Modules.scala 56:109:@40602.4]
  wire [10:0] buffer_10_708; // @[Modules.scala 56:109:@40603.4]
  wire [11:0] _T_88443; // @[Modules.scala 56:109:@40605.4]
  wire [10:0] _T_88444; // @[Modules.scala 56:109:@40606.4]
  wire [10:0] buffer_10_709; // @[Modules.scala 56:109:@40607.4]
  wire [11:0] _T_88446; // @[Modules.scala 56:109:@40609.4]
  wire [10:0] _T_88447; // @[Modules.scala 56:109:@40610.4]
  wire [10:0] buffer_10_710; // @[Modules.scala 56:109:@40611.4]
  wire [11:0] _T_88449; // @[Modules.scala 56:109:@40613.4]
  wire [10:0] _T_88450; // @[Modules.scala 56:109:@40614.4]
  wire [10:0] buffer_10_711; // @[Modules.scala 56:109:@40615.4]
  wire [11:0] _T_88452; // @[Modules.scala 56:109:@40617.4]
  wire [10:0] _T_88453; // @[Modules.scala 56:109:@40618.4]
  wire [10:0] buffer_10_712; // @[Modules.scala 56:109:@40619.4]
  wire [11:0] _T_88455; // @[Modules.scala 56:109:@40621.4]
  wire [10:0] _T_88456; // @[Modules.scala 56:109:@40622.4]
  wire [10:0] buffer_10_713; // @[Modules.scala 56:109:@40623.4]
  wire [11:0] _T_88458; // @[Modules.scala 56:109:@40625.4]
  wire [10:0] _T_88459; // @[Modules.scala 56:109:@40626.4]
  wire [10:0] buffer_10_714; // @[Modules.scala 56:109:@40627.4]
  wire [11:0] _T_88461; // @[Modules.scala 56:109:@40629.4]
  wire [10:0] _T_88462; // @[Modules.scala 56:109:@40630.4]
  wire [10:0] buffer_10_715; // @[Modules.scala 56:109:@40631.4]
  wire [11:0] _T_88464; // @[Modules.scala 56:109:@40633.4]
  wire [10:0] _T_88465; // @[Modules.scala 56:109:@40634.4]
  wire [10:0] buffer_10_716; // @[Modules.scala 56:109:@40635.4]
  wire [11:0] _T_88467; // @[Modules.scala 56:109:@40637.4]
  wire [10:0] _T_88468; // @[Modules.scala 56:109:@40638.4]
  wire [10:0] buffer_10_717; // @[Modules.scala 56:109:@40639.4]
  wire [11:0] _T_88470; // @[Modules.scala 56:109:@40641.4]
  wire [10:0] _T_88471; // @[Modules.scala 56:109:@40642.4]
  wire [10:0] buffer_10_718; // @[Modules.scala 56:109:@40643.4]
  wire [11:0] _T_88473; // @[Modules.scala 56:109:@40645.4]
  wire [10:0] _T_88474; // @[Modules.scala 56:109:@40646.4]
  wire [10:0] buffer_10_719; // @[Modules.scala 56:109:@40647.4]
  wire [11:0] _T_88476; // @[Modules.scala 56:109:@40649.4]
  wire [10:0] _T_88477; // @[Modules.scala 56:109:@40650.4]
  wire [10:0] buffer_10_720; // @[Modules.scala 56:109:@40651.4]
  wire [11:0] _T_88479; // @[Modules.scala 56:109:@40653.4]
  wire [10:0] _T_88480; // @[Modules.scala 56:109:@40654.4]
  wire [10:0] buffer_10_721; // @[Modules.scala 56:109:@40655.4]
  wire [11:0] _T_88482; // @[Modules.scala 56:109:@40657.4]
  wire [10:0] _T_88483; // @[Modules.scala 56:109:@40658.4]
  wire [10:0] buffer_10_722; // @[Modules.scala 56:109:@40659.4]
  wire [11:0] _T_88485; // @[Modules.scala 56:109:@40661.4]
  wire [10:0] _T_88486; // @[Modules.scala 56:109:@40662.4]
  wire [10:0] buffer_10_723; // @[Modules.scala 56:109:@40663.4]
  wire [11:0] _T_88488; // @[Modules.scala 56:109:@40665.4]
  wire [10:0] _T_88489; // @[Modules.scala 56:109:@40666.4]
  wire [10:0] buffer_10_724; // @[Modules.scala 56:109:@40667.4]
  wire [11:0] _T_88491; // @[Modules.scala 56:109:@40669.4]
  wire [10:0] _T_88492; // @[Modules.scala 56:109:@40670.4]
  wire [10:0] buffer_10_725; // @[Modules.scala 56:109:@40671.4]
  wire [11:0] _T_88494; // @[Modules.scala 56:109:@40673.4]
  wire [10:0] _T_88495; // @[Modules.scala 56:109:@40674.4]
  wire [10:0] buffer_10_726; // @[Modules.scala 56:109:@40675.4]
  wire [11:0] _T_88497; // @[Modules.scala 56:109:@40677.4]
  wire [10:0] _T_88498; // @[Modules.scala 56:109:@40678.4]
  wire [10:0] buffer_10_727; // @[Modules.scala 56:109:@40679.4]
  wire [11:0] _T_88500; // @[Modules.scala 56:109:@40681.4]
  wire [10:0] _T_88501; // @[Modules.scala 56:109:@40682.4]
  wire [10:0] buffer_10_728; // @[Modules.scala 56:109:@40683.4]
  wire [11:0] _T_88503; // @[Modules.scala 56:109:@40685.4]
  wire [10:0] _T_88504; // @[Modules.scala 56:109:@40686.4]
  wire [10:0] buffer_10_729; // @[Modules.scala 56:109:@40687.4]
  wire [11:0] _T_88506; // @[Modules.scala 56:109:@40689.4]
  wire [10:0] _T_88507; // @[Modules.scala 56:109:@40690.4]
  wire [10:0] buffer_10_730; // @[Modules.scala 56:109:@40691.4]
  wire [11:0] _T_88509; // @[Modules.scala 56:109:@40693.4]
  wire [10:0] _T_88510; // @[Modules.scala 56:109:@40694.4]
  wire [10:0] buffer_10_731; // @[Modules.scala 56:109:@40695.4]
  wire [11:0] _T_88512; // @[Modules.scala 56:109:@40697.4]
  wire [10:0] _T_88513; // @[Modules.scala 56:109:@40698.4]
  wire [10:0] buffer_10_732; // @[Modules.scala 56:109:@40699.4]
  wire [11:0] _T_88515; // @[Modules.scala 56:109:@40701.4]
  wire [10:0] _T_88516; // @[Modules.scala 56:109:@40702.4]
  wire [10:0] buffer_10_733; // @[Modules.scala 56:109:@40703.4]
  wire [11:0] _T_88518; // @[Modules.scala 56:109:@40705.4]
  wire [10:0] _T_88519; // @[Modules.scala 56:109:@40706.4]
  wire [10:0] buffer_10_734; // @[Modules.scala 56:109:@40707.4]
  wire [11:0] _T_88521; // @[Modules.scala 63:156:@40710.4]
  wire [10:0] _T_88522; // @[Modules.scala 63:156:@40711.4]
  wire [10:0] buffer_10_736; // @[Modules.scala 63:156:@40712.4]
  wire [11:0] _T_88524; // @[Modules.scala 63:156:@40714.4]
  wire [10:0] _T_88525; // @[Modules.scala 63:156:@40715.4]
  wire [10:0] buffer_10_737; // @[Modules.scala 63:156:@40716.4]
  wire [11:0] _T_88527; // @[Modules.scala 63:156:@40718.4]
  wire [10:0] _T_88528; // @[Modules.scala 63:156:@40719.4]
  wire [10:0] buffer_10_738; // @[Modules.scala 63:156:@40720.4]
  wire [11:0] _T_88530; // @[Modules.scala 63:156:@40722.4]
  wire [10:0] _T_88531; // @[Modules.scala 63:156:@40723.4]
  wire [10:0] buffer_10_739; // @[Modules.scala 63:156:@40724.4]
  wire [11:0] _T_88533; // @[Modules.scala 63:156:@40726.4]
  wire [10:0] _T_88534; // @[Modules.scala 63:156:@40727.4]
  wire [10:0] buffer_10_740; // @[Modules.scala 63:156:@40728.4]
  wire [11:0] _T_88536; // @[Modules.scala 63:156:@40730.4]
  wire [10:0] _T_88537; // @[Modules.scala 63:156:@40731.4]
  wire [10:0] buffer_10_741; // @[Modules.scala 63:156:@40732.4]
  wire [11:0] _T_88539; // @[Modules.scala 63:156:@40734.4]
  wire [10:0] _T_88540; // @[Modules.scala 63:156:@40735.4]
  wire [10:0] buffer_10_742; // @[Modules.scala 63:156:@40736.4]
  wire [11:0] _T_88542; // @[Modules.scala 63:156:@40738.4]
  wire [10:0] _T_88543; // @[Modules.scala 63:156:@40739.4]
  wire [10:0] buffer_10_743; // @[Modules.scala 63:156:@40740.4]
  wire [11:0] _T_88545; // @[Modules.scala 63:156:@40742.4]
  wire [10:0] _T_88546; // @[Modules.scala 63:156:@40743.4]
  wire [10:0] buffer_10_744; // @[Modules.scala 63:156:@40744.4]
  wire [11:0] _T_88548; // @[Modules.scala 63:156:@40746.4]
  wire [10:0] _T_88549; // @[Modules.scala 63:156:@40747.4]
  wire [10:0] buffer_10_745; // @[Modules.scala 63:156:@40748.4]
  wire [11:0] _T_88551; // @[Modules.scala 63:156:@40750.4]
  wire [10:0] _T_88552; // @[Modules.scala 63:156:@40751.4]
  wire [10:0] buffer_10_746; // @[Modules.scala 63:156:@40752.4]
  wire [11:0] _T_88554; // @[Modules.scala 63:156:@40754.4]
  wire [10:0] _T_88555; // @[Modules.scala 63:156:@40755.4]
  wire [10:0] buffer_10_747; // @[Modules.scala 63:156:@40756.4]
  wire [11:0] _T_88557; // @[Modules.scala 63:156:@40758.4]
  wire [10:0] _T_88558; // @[Modules.scala 63:156:@40759.4]
  wire [10:0] buffer_10_748; // @[Modules.scala 63:156:@40760.4]
  wire [11:0] _T_88560; // @[Modules.scala 63:156:@40762.4]
  wire [10:0] _T_88561; // @[Modules.scala 63:156:@40763.4]
  wire [10:0] buffer_10_749; // @[Modules.scala 63:156:@40764.4]
  wire [11:0] _T_88563; // @[Modules.scala 63:156:@40766.4]
  wire [10:0] _T_88564; // @[Modules.scala 63:156:@40767.4]
  wire [10:0] buffer_10_750; // @[Modules.scala 63:156:@40768.4]
  wire [11:0] _T_88566; // @[Modules.scala 63:156:@40770.4]
  wire [10:0] _T_88567; // @[Modules.scala 63:156:@40771.4]
  wire [10:0] buffer_10_751; // @[Modules.scala 63:156:@40772.4]
  wire [11:0] _T_88569; // @[Modules.scala 63:156:@40774.4]
  wire [10:0] _T_88570; // @[Modules.scala 63:156:@40775.4]
  wire [10:0] buffer_10_752; // @[Modules.scala 63:156:@40776.4]
  wire [11:0] _T_88572; // @[Modules.scala 63:156:@40778.4]
  wire [10:0] _T_88573; // @[Modules.scala 63:156:@40779.4]
  wire [10:0] buffer_10_753; // @[Modules.scala 63:156:@40780.4]
  wire [11:0] _T_88575; // @[Modules.scala 63:156:@40782.4]
  wire [10:0] _T_88576; // @[Modules.scala 63:156:@40783.4]
  wire [10:0] buffer_10_754; // @[Modules.scala 63:156:@40784.4]
  wire [11:0] _T_88578; // @[Modules.scala 63:156:@40786.4]
  wire [10:0] _T_88579; // @[Modules.scala 63:156:@40787.4]
  wire [10:0] buffer_10_755; // @[Modules.scala 63:156:@40788.4]
  wire [11:0] _T_88581; // @[Modules.scala 63:156:@40790.4]
  wire [10:0] _T_88582; // @[Modules.scala 63:156:@40791.4]
  wire [10:0] buffer_10_756; // @[Modules.scala 63:156:@40792.4]
  wire [11:0] _T_88584; // @[Modules.scala 63:156:@40794.4]
  wire [10:0] _T_88585; // @[Modules.scala 63:156:@40795.4]
  wire [10:0] buffer_10_757; // @[Modules.scala 63:156:@40796.4]
  wire [11:0] _T_88587; // @[Modules.scala 63:156:@40798.4]
  wire [10:0] _T_88588; // @[Modules.scala 63:156:@40799.4]
  wire [10:0] buffer_10_758; // @[Modules.scala 63:156:@40800.4]
  wire [11:0] _T_88590; // @[Modules.scala 63:156:@40802.4]
  wire [10:0] _T_88591; // @[Modules.scala 63:156:@40803.4]
  wire [10:0] buffer_10_759; // @[Modules.scala 63:156:@40804.4]
  wire [11:0] _T_88593; // @[Modules.scala 63:156:@40806.4]
  wire [10:0] _T_88594; // @[Modules.scala 63:156:@40807.4]
  wire [10:0] buffer_10_760; // @[Modules.scala 63:156:@40808.4]
  wire [11:0] _T_88596; // @[Modules.scala 63:156:@40810.4]
  wire [10:0] _T_88597; // @[Modules.scala 63:156:@40811.4]
  wire [10:0] buffer_10_761; // @[Modules.scala 63:156:@40812.4]
  wire [11:0] _T_88599; // @[Modules.scala 63:156:@40814.4]
  wire [10:0] _T_88600; // @[Modules.scala 63:156:@40815.4]
  wire [10:0] buffer_10_762; // @[Modules.scala 63:156:@40816.4]
  wire [11:0] _T_88602; // @[Modules.scala 63:156:@40818.4]
  wire [10:0] _T_88603; // @[Modules.scala 63:156:@40819.4]
  wire [10:0] buffer_10_763; // @[Modules.scala 63:156:@40820.4]
  wire [11:0] _T_88605; // @[Modules.scala 63:156:@40822.4]
  wire [10:0] _T_88606; // @[Modules.scala 63:156:@40823.4]
  wire [10:0] buffer_10_764; // @[Modules.scala 63:156:@40824.4]
  wire [11:0] _T_88608; // @[Modules.scala 63:156:@40826.4]
  wire [10:0] _T_88609; // @[Modules.scala 63:156:@40827.4]
  wire [10:0] buffer_10_765; // @[Modules.scala 63:156:@40828.4]
  wire [11:0] _T_88611; // @[Modules.scala 63:156:@40830.4]
  wire [10:0] _T_88612; // @[Modules.scala 63:156:@40831.4]
  wire [10:0] buffer_10_766; // @[Modules.scala 63:156:@40832.4]
  wire [11:0] _T_88614; // @[Modules.scala 63:156:@40834.4]
  wire [10:0] _T_88615; // @[Modules.scala 63:156:@40835.4]
  wire [10:0] buffer_10_767; // @[Modules.scala 63:156:@40836.4]
  wire [11:0] _T_88617; // @[Modules.scala 63:156:@40838.4]
  wire [10:0] _T_88618; // @[Modules.scala 63:156:@40839.4]
  wire [10:0] buffer_10_768; // @[Modules.scala 63:156:@40840.4]
  wire [11:0] _T_88620; // @[Modules.scala 63:156:@40842.4]
  wire [10:0] _T_88621; // @[Modules.scala 63:156:@40843.4]
  wire [10:0] buffer_10_769; // @[Modules.scala 63:156:@40844.4]
  wire [11:0] _T_88623; // @[Modules.scala 63:156:@40846.4]
  wire [10:0] _T_88624; // @[Modules.scala 63:156:@40847.4]
  wire [10:0] buffer_10_770; // @[Modules.scala 63:156:@40848.4]
  wire [11:0] _T_88626; // @[Modules.scala 63:156:@40850.4]
  wire [10:0] _T_88627; // @[Modules.scala 63:156:@40851.4]
  wire [10:0] buffer_10_771; // @[Modules.scala 63:156:@40852.4]
  wire [11:0] _T_88629; // @[Modules.scala 63:156:@40854.4]
  wire [10:0] _T_88630; // @[Modules.scala 63:156:@40855.4]
  wire [10:0] buffer_10_772; // @[Modules.scala 63:156:@40856.4]
  wire [11:0] _T_88632; // @[Modules.scala 63:156:@40858.4]
  wire [10:0] _T_88633; // @[Modules.scala 63:156:@40859.4]
  wire [10:0] buffer_10_773; // @[Modules.scala 63:156:@40860.4]
  wire [11:0] _T_88635; // @[Modules.scala 63:156:@40862.4]
  wire [10:0] _T_88636; // @[Modules.scala 63:156:@40863.4]
  wire [10:0] buffer_10_774; // @[Modules.scala 63:156:@40864.4]
  wire [11:0] _T_88638; // @[Modules.scala 63:156:@40866.4]
  wire [10:0] _T_88639; // @[Modules.scala 63:156:@40867.4]
  wire [10:0] buffer_10_775; // @[Modules.scala 63:156:@40868.4]
  wire [11:0] _T_88641; // @[Modules.scala 63:156:@40870.4]
  wire [10:0] _T_88642; // @[Modules.scala 63:156:@40871.4]
  wire [10:0] buffer_10_776; // @[Modules.scala 63:156:@40872.4]
  wire [11:0] _T_88644; // @[Modules.scala 63:156:@40874.4]
  wire [10:0] _T_88645; // @[Modules.scala 63:156:@40875.4]
  wire [10:0] buffer_10_777; // @[Modules.scala 63:156:@40876.4]
  wire [11:0] _T_88647; // @[Modules.scala 63:156:@40878.4]
  wire [10:0] _T_88648; // @[Modules.scala 63:156:@40879.4]
  wire [10:0] buffer_10_778; // @[Modules.scala 63:156:@40880.4]
  wire [11:0] _T_88650; // @[Modules.scala 63:156:@40882.4]
  wire [10:0] _T_88651; // @[Modules.scala 63:156:@40883.4]
  wire [10:0] buffer_10_779; // @[Modules.scala 63:156:@40884.4]
  wire [11:0] _T_88653; // @[Modules.scala 63:156:@40886.4]
  wire [10:0] _T_88654; // @[Modules.scala 63:156:@40887.4]
  wire [10:0] buffer_10_780; // @[Modules.scala 63:156:@40888.4]
  wire [11:0] _T_88656; // @[Modules.scala 63:156:@40890.4]
  wire [10:0] _T_88657; // @[Modules.scala 63:156:@40891.4]
  wire [10:0] buffer_10_781; // @[Modules.scala 63:156:@40892.4]
  wire [11:0] _T_88659; // @[Modules.scala 63:156:@40894.4]
  wire [10:0] _T_88660; // @[Modules.scala 63:156:@40895.4]
  wire [10:0] buffer_10_782; // @[Modules.scala 63:156:@40896.4]
  wire [11:0] _T_88662; // @[Modules.scala 63:156:@40898.4]
  wire [10:0] _T_88663; // @[Modules.scala 63:156:@40899.4]
  wire [10:0] buffer_10_783; // @[Modules.scala 63:156:@40900.4]
  wire [5:0] _T_88750; // @[Modules.scala 43:47:@41000.4]
  wire [4:0] _T_88751; // @[Modules.scala 43:47:@41001.4]
  wire [4:0] _T_88752; // @[Modules.scala 43:47:@41002.4]
  wire [5:0] _T_88759; // @[Modules.scala 40:46:@41012.4]
  wire [4:0] _T_88760; // @[Modules.scala 40:46:@41013.4]
  wire [4:0] _T_88761; // @[Modules.scala 40:46:@41014.4]
  wire [5:0] _T_88766; // @[Modules.scala 43:47:@41019.4]
  wire [4:0] _T_88767; // @[Modules.scala 43:47:@41020.4]
  wire [4:0] _T_88768; // @[Modules.scala 43:47:@41021.4]
  wire [5:0] _T_88878; // @[Modules.scala 37:46:@41138.4]
  wire [4:0] _T_88879; // @[Modules.scala 37:46:@41139.4]
  wire [4:0] _T_88880; // @[Modules.scala 37:46:@41140.4]
  wire [5:0] _T_89147; // @[Modules.scala 43:47:@41422.4]
  wire [4:0] _T_89148; // @[Modules.scala 43:47:@41423.4]
  wire [4:0] _T_89149; // @[Modules.scala 43:47:@41424.4]
  wire [5:0] _T_89220; // @[Modules.scala 43:47:@41503.4]
  wire [4:0] _T_89221; // @[Modules.scala 43:47:@41504.4]
  wire [4:0] _T_89222; // @[Modules.scala 43:47:@41505.4]
  wire [5:0] _T_89245; // @[Modules.scala 40:46:@41534.4]
  wire [4:0] _T_89246; // @[Modules.scala 40:46:@41535.4]
  wire [4:0] _T_89247; // @[Modules.scala 40:46:@41536.4]
  wire [5:0] _T_89286; // @[Modules.scala 43:47:@41577.4]
  wire [4:0] _T_89287; // @[Modules.scala 43:47:@41578.4]
  wire [4:0] _T_89288; // @[Modules.scala 43:47:@41579.4]
  wire [5:0] _T_89366; // @[Modules.scala 43:47:@41665.4]
  wire [4:0] _T_89367; // @[Modules.scala 43:47:@41666.4]
  wire [4:0] _T_89368; // @[Modules.scala 43:47:@41667.4]
  wire [5:0] _T_89604; // @[Modules.scala 43:47:@41931.4]
  wire [4:0] _T_89605; // @[Modules.scala 43:47:@41932.4]
  wire [4:0] _T_89606; // @[Modules.scala 43:47:@41933.4]
  wire [5:0] _T_89611; // @[Modules.scala 43:47:@41938.4]
  wire [4:0] _T_89612; // @[Modules.scala 43:47:@41939.4]
  wire [4:0] _T_89613; // @[Modules.scala 43:47:@41940.4]
  wire [5:0] _T_89767; // @[Modules.scala 43:47:@42104.4]
  wire [4:0] _T_89768; // @[Modules.scala 43:47:@42105.4]
  wire [4:0] _T_89769; // @[Modules.scala 43:47:@42106.4]
  wire [5:0] _T_89780; // @[Modules.scala 40:46:@42119.4]
  wire [4:0] _T_89781; // @[Modules.scala 40:46:@42120.4]
  wire [4:0] _T_89782; // @[Modules.scala 40:46:@42121.4]
  wire [5:0] _T_89832; // @[Modules.scala 40:46:@42172.4]
  wire [4:0] _T_89833; // @[Modules.scala 40:46:@42173.4]
  wire [4:0] _T_89834; // @[Modules.scala 40:46:@42174.4]
  wire [5:0] _T_89894; // @[Modules.scala 43:47:@42236.4]
  wire [4:0] _T_89895; // @[Modules.scala 43:47:@42237.4]
  wire [4:0] _T_89896; // @[Modules.scala 43:47:@42238.4]
  wire [5:0] _T_89929; // @[Modules.scala 43:47:@42271.4]
  wire [4:0] _T_89930; // @[Modules.scala 43:47:@42272.4]
  wire [4:0] _T_89931; // @[Modules.scala 43:47:@42273.4]
  wire [5:0] _T_89980; // @[Modules.scala 43:47:@42325.4]
  wire [4:0] _T_89981; // @[Modules.scala 43:47:@42326.4]
  wire [4:0] _T_89982; // @[Modules.scala 43:47:@42327.4]
  wire [5:0] _T_90031; // @[Modules.scala 43:47:@42379.4]
  wire [4:0] _T_90032; // @[Modules.scala 43:47:@42380.4]
  wire [4:0] _T_90033; // @[Modules.scala 43:47:@42381.4]
  wire [5:0] _T_90168; // @[Modules.scala 40:46:@42522.4]
  wire [4:0] _T_90169; // @[Modules.scala 40:46:@42523.4]
  wire [4:0] _T_90170; // @[Modules.scala 40:46:@42524.4]
  wire [5:0] _T_90323; // @[Modules.scala 43:47:@42689.4]
  wire [4:0] _T_90324; // @[Modules.scala 43:47:@42690.4]
  wire [4:0] _T_90325; // @[Modules.scala 43:47:@42691.4]
  wire [5:0] _T_90592; // @[Modules.scala 43:47:@42980.4]
  wire [4:0] _T_90593; // @[Modules.scala 43:47:@42981.4]
  wire [4:0] _T_90594; // @[Modules.scala 43:47:@42982.4]
  wire [11:0] _T_90793; // @[Modules.scala 50:57:@43192.4]
  wire [10:0] _T_90794; // @[Modules.scala 50:57:@43193.4]
  wire [10:0] buffer_11_396; // @[Modules.scala 50:57:@43194.4]
  wire [11:0] _T_90796; // @[Modules.scala 50:57:@43196.4]
  wire [10:0] _T_90797; // @[Modules.scala 50:57:@43197.4]
  wire [10:0] buffer_11_397; // @[Modules.scala 50:57:@43198.4]
  wire [11:0] _T_90802; // @[Modules.scala 50:57:@43204.4]
  wire [10:0] _T_90803; // @[Modules.scala 50:57:@43205.4]
  wire [10:0] buffer_11_399; // @[Modules.scala 50:57:@43206.4]
  wire [10:0] buffer_11_19; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90808; // @[Modules.scala 50:57:@43212.4]
  wire [10:0] _T_90809; // @[Modules.scala 50:57:@43213.4]
  wire [10:0] buffer_11_401; // @[Modules.scala 50:57:@43214.4]
  wire [10:0] buffer_11_22; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_11_23; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90814; // @[Modules.scala 50:57:@43220.4]
  wire [10:0] _T_90815; // @[Modules.scala 50:57:@43221.4]
  wire [10:0] buffer_11_403; // @[Modules.scala 50:57:@43222.4]
  wire [11:0] _T_90820; // @[Modules.scala 50:57:@43228.4]
  wire [10:0] _T_90821; // @[Modules.scala 50:57:@43229.4]
  wire [10:0] buffer_11_405; // @[Modules.scala 50:57:@43230.4]
  wire [11:0] _T_90823; // @[Modules.scala 50:57:@43232.4]
  wire [10:0] _T_90824; // @[Modules.scala 50:57:@43233.4]
  wire [10:0] buffer_11_406; // @[Modules.scala 50:57:@43234.4]
  wire [11:0] _T_90832; // @[Modules.scala 50:57:@43244.4]
  wire [10:0] _T_90833; // @[Modules.scala 50:57:@43245.4]
  wire [10:0] buffer_11_409; // @[Modules.scala 50:57:@43246.4]
  wire [10:0] buffer_11_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90844; // @[Modules.scala 50:57:@43260.4]
  wire [10:0] _T_90845; // @[Modules.scala 50:57:@43261.4]
  wire [10:0] buffer_11_413; // @[Modules.scala 50:57:@43262.4]
  wire [11:0] _T_90847; // @[Modules.scala 50:57:@43264.4]
  wire [10:0] _T_90848; // @[Modules.scala 50:57:@43265.4]
  wire [10:0] buffer_11_414; // @[Modules.scala 50:57:@43266.4]
  wire [11:0] _T_90883; // @[Modules.scala 50:57:@43312.4]
  wire [10:0] _T_90884; // @[Modules.scala 50:57:@43313.4]
  wire [10:0] buffer_11_426; // @[Modules.scala 50:57:@43314.4]
  wire [11:0] _T_90886; // @[Modules.scala 50:57:@43316.4]
  wire [10:0] _T_90887; // @[Modules.scala 50:57:@43317.4]
  wire [10:0] buffer_11_427; // @[Modules.scala 50:57:@43318.4]
  wire [11:0] _T_90904; // @[Modules.scala 50:57:@43340.4]
  wire [10:0] _T_90905; // @[Modules.scala 50:57:@43341.4]
  wire [10:0] buffer_11_433; // @[Modules.scala 50:57:@43342.4]
  wire [10:0] buffer_11_90; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90916; // @[Modules.scala 50:57:@43356.4]
  wire [10:0] _T_90917; // @[Modules.scala 50:57:@43357.4]
  wire [10:0] buffer_11_437; // @[Modules.scala 50:57:@43358.4]
  wire [11:0] _T_90919; // @[Modules.scala 50:57:@43360.4]
  wire [10:0] _T_90920; // @[Modules.scala 50:57:@43361.4]
  wire [10:0] buffer_11_438; // @[Modules.scala 50:57:@43362.4]
  wire [11:0] _T_90922; // @[Modules.scala 50:57:@43364.4]
  wire [10:0] _T_90923; // @[Modules.scala 50:57:@43365.4]
  wire [10:0] buffer_11_439; // @[Modules.scala 50:57:@43366.4]
  wire [11:0] _T_90928; // @[Modules.scala 50:57:@43372.4]
  wire [10:0] _T_90929; // @[Modules.scala 50:57:@43373.4]
  wire [10:0] buffer_11_441; // @[Modules.scala 50:57:@43374.4]
  wire [10:0] buffer_11_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90937; // @[Modules.scala 50:57:@43384.4]
  wire [10:0] _T_90938; // @[Modules.scala 50:57:@43385.4]
  wire [10:0] buffer_11_444; // @[Modules.scala 50:57:@43386.4]
  wire [11:0] _T_90940; // @[Modules.scala 50:57:@43388.4]
  wire [10:0] _T_90941; // @[Modules.scala 50:57:@43389.4]
  wire [10:0] buffer_11_445; // @[Modules.scala 50:57:@43390.4]
  wire [10:0] buffer_11_112; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90949; // @[Modules.scala 50:57:@43400.4]
  wire [10:0] _T_90950; // @[Modules.scala 50:57:@43401.4]
  wire [10:0] buffer_11_448; // @[Modules.scala 50:57:@43402.4]
  wire [11:0] _T_90955; // @[Modules.scala 50:57:@43408.4]
  wire [10:0] _T_90956; // @[Modules.scala 50:57:@43409.4]
  wire [10:0] buffer_11_450; // @[Modules.scala 50:57:@43410.4]
  wire [10:0] buffer_11_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90958; // @[Modules.scala 50:57:@43412.4]
  wire [10:0] _T_90959; // @[Modules.scala 50:57:@43413.4]
  wire [10:0] buffer_11_451; // @[Modules.scala 50:57:@43414.4]
  wire [11:0] _T_90961; // @[Modules.scala 50:57:@43416.4]
  wire [10:0] _T_90962; // @[Modules.scala 50:57:@43417.4]
  wire [10:0] buffer_11_452; // @[Modules.scala 50:57:@43418.4]
  wire [11:0] _T_90964; // @[Modules.scala 50:57:@43420.4]
  wire [10:0] _T_90965; // @[Modules.scala 50:57:@43421.4]
  wire [10:0] buffer_11_453; // @[Modules.scala 50:57:@43422.4]
  wire [11:0] _T_90973; // @[Modules.scala 50:57:@43432.4]
  wire [10:0] _T_90974; // @[Modules.scala 50:57:@43433.4]
  wire [10:0] buffer_11_456; // @[Modules.scala 50:57:@43434.4]
  wire [11:0] _T_90979; // @[Modules.scala 50:57:@43440.4]
  wire [10:0] _T_90980; // @[Modules.scala 50:57:@43441.4]
  wire [10:0] buffer_11_458; // @[Modules.scala 50:57:@43442.4]
  wire [10:0] buffer_11_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_90982; // @[Modules.scala 50:57:@43444.4]
  wire [10:0] _T_90983; // @[Modules.scala 50:57:@43445.4]
  wire [10:0] buffer_11_459; // @[Modules.scala 50:57:@43446.4]
  wire [11:0] _T_90991; // @[Modules.scala 50:57:@43456.4]
  wire [10:0] _T_90992; // @[Modules.scala 50:57:@43457.4]
  wire [10:0] buffer_11_462; // @[Modules.scala 50:57:@43458.4]
  wire [11:0] _T_90994; // @[Modules.scala 50:57:@43460.4]
  wire [10:0] _T_90995; // @[Modules.scala 50:57:@43461.4]
  wire [10:0] buffer_11_463; // @[Modules.scala 50:57:@43462.4]
  wire [11:0] _T_91015; // @[Modules.scala 50:57:@43488.4]
  wire [10:0] _T_91016; // @[Modules.scala 50:57:@43489.4]
  wire [10:0] buffer_11_470; // @[Modules.scala 50:57:@43490.4]
  wire [11:0] _T_91021; // @[Modules.scala 50:57:@43496.4]
  wire [10:0] _T_91022; // @[Modules.scala 50:57:@43497.4]
  wire [10:0] buffer_11_472; // @[Modules.scala 50:57:@43498.4]
  wire [11:0] _T_91051; // @[Modules.scala 50:57:@43536.4]
  wire [10:0] _T_91052; // @[Modules.scala 50:57:@43537.4]
  wire [10:0] buffer_11_482; // @[Modules.scala 50:57:@43538.4]
  wire [10:0] buffer_11_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91057; // @[Modules.scala 50:57:@43544.4]
  wire [10:0] _T_91058; // @[Modules.scala 50:57:@43545.4]
  wire [10:0] buffer_11_484; // @[Modules.scala 50:57:@43546.4]
  wire [10:0] buffer_11_186; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91060; // @[Modules.scala 50:57:@43548.4]
  wire [10:0] _T_91061; // @[Modules.scala 50:57:@43549.4]
  wire [10:0] buffer_11_485; // @[Modules.scala 50:57:@43550.4]
  wire [11:0] _T_91072; // @[Modules.scala 50:57:@43564.4]
  wire [10:0] _T_91073; // @[Modules.scala 50:57:@43565.4]
  wire [10:0] buffer_11_489; // @[Modules.scala 50:57:@43566.4]
  wire [11:0] _T_91081; // @[Modules.scala 50:57:@43576.4]
  wire [10:0] _T_91082; // @[Modules.scala 50:57:@43577.4]
  wire [10:0] buffer_11_492; // @[Modules.scala 50:57:@43578.4]
  wire [11:0] _T_91087; // @[Modules.scala 50:57:@43584.4]
  wire [10:0] _T_91088; // @[Modules.scala 50:57:@43585.4]
  wire [10:0] buffer_11_494; // @[Modules.scala 50:57:@43586.4]
  wire [11:0] _T_91096; // @[Modules.scala 50:57:@43596.4]
  wire [10:0] _T_91097; // @[Modules.scala 50:57:@43597.4]
  wire [10:0] buffer_11_497; // @[Modules.scala 50:57:@43598.4]
  wire [10:0] buffer_11_214; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91102; // @[Modules.scala 50:57:@43604.4]
  wire [10:0] _T_91103; // @[Modules.scala 50:57:@43605.4]
  wire [10:0] buffer_11_499; // @[Modules.scala 50:57:@43606.4]
  wire [10:0] buffer_11_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91105; // @[Modules.scala 50:57:@43608.4]
  wire [10:0] _T_91106; // @[Modules.scala 50:57:@43609.4]
  wire [10:0] buffer_11_500; // @[Modules.scala 50:57:@43610.4]
  wire [10:0] buffer_11_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91117; // @[Modules.scala 50:57:@43624.4]
  wire [10:0] _T_91118; // @[Modules.scala 50:57:@43625.4]
  wire [10:0] buffer_11_504; // @[Modules.scala 50:57:@43626.4]
  wire [11:0] _T_91123; // @[Modules.scala 50:57:@43632.4]
  wire [10:0] _T_91124; // @[Modules.scala 50:57:@43633.4]
  wire [10:0] buffer_11_506; // @[Modules.scala 50:57:@43634.4]
  wire [10:0] buffer_11_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91132; // @[Modules.scala 50:57:@43644.4]
  wire [10:0] _T_91133; // @[Modules.scala 50:57:@43645.4]
  wire [10:0] buffer_11_509; // @[Modules.scala 50:57:@43646.4]
  wire [11:0] _T_91138; // @[Modules.scala 50:57:@43652.4]
  wire [10:0] _T_91139; // @[Modules.scala 50:57:@43653.4]
  wire [10:0] buffer_11_511; // @[Modules.scala 50:57:@43654.4]
  wire [10:0] buffer_11_240; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91141; // @[Modules.scala 50:57:@43656.4]
  wire [10:0] _T_91142; // @[Modules.scala 50:57:@43657.4]
  wire [10:0] buffer_11_512; // @[Modules.scala 50:57:@43658.4]
  wire [10:0] buffer_11_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91153; // @[Modules.scala 50:57:@43672.4]
  wire [10:0] _T_91154; // @[Modules.scala 50:57:@43673.4]
  wire [10:0] buffer_11_516; // @[Modules.scala 50:57:@43674.4]
  wire [11:0] _T_91165; // @[Modules.scala 50:57:@43688.4]
  wire [10:0] _T_91166; // @[Modules.scala 50:57:@43689.4]
  wire [10:0] buffer_11_520; // @[Modules.scala 50:57:@43690.4]
  wire [10:0] buffer_11_258; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91168; // @[Modules.scala 50:57:@43692.4]
  wire [10:0] _T_91169; // @[Modules.scala 50:57:@43693.4]
  wire [10:0] buffer_11_521; // @[Modules.scala 50:57:@43694.4]
  wire [11:0] _T_91174; // @[Modules.scala 50:57:@43700.4]
  wire [10:0] _T_91175; // @[Modules.scala 50:57:@43701.4]
  wire [10:0] buffer_11_523; // @[Modules.scala 50:57:@43702.4]
  wire [11:0] _T_91186; // @[Modules.scala 50:57:@43716.4]
  wire [10:0] _T_91187; // @[Modules.scala 50:57:@43717.4]
  wire [10:0] buffer_11_527; // @[Modules.scala 50:57:@43718.4]
  wire [11:0] _T_91189; // @[Modules.scala 50:57:@43720.4]
  wire [10:0] _T_91190; // @[Modules.scala 50:57:@43721.4]
  wire [10:0] buffer_11_528; // @[Modules.scala 50:57:@43722.4]
  wire [11:0] _T_91195; // @[Modules.scala 50:57:@43728.4]
  wire [10:0] _T_91196; // @[Modules.scala 50:57:@43729.4]
  wire [10:0] buffer_11_530; // @[Modules.scala 50:57:@43730.4]
  wire [10:0] buffer_11_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91201; // @[Modules.scala 50:57:@43736.4]
  wire [10:0] _T_91202; // @[Modules.scala 50:57:@43737.4]
  wire [10:0] buffer_11_532; // @[Modules.scala 50:57:@43738.4]
  wire [11:0] _T_91210; // @[Modules.scala 50:57:@43748.4]
  wire [10:0] _T_91211; // @[Modules.scala 50:57:@43749.4]
  wire [10:0] buffer_11_535; // @[Modules.scala 50:57:@43750.4]
  wire [11:0] _T_91216; // @[Modules.scala 50:57:@43756.4]
  wire [10:0] _T_91217; // @[Modules.scala 50:57:@43757.4]
  wire [10:0] buffer_11_537; // @[Modules.scala 50:57:@43758.4]
  wire [11:0] _T_91225; // @[Modules.scala 50:57:@43768.4]
  wire [10:0] _T_91226; // @[Modules.scala 50:57:@43769.4]
  wire [10:0] buffer_11_540; // @[Modules.scala 50:57:@43770.4]
  wire [11:0] _T_91234; // @[Modules.scala 50:57:@43780.4]
  wire [10:0] _T_91235; // @[Modules.scala 50:57:@43781.4]
  wire [10:0] buffer_11_543; // @[Modules.scala 50:57:@43782.4]
  wire [11:0] _T_91240; // @[Modules.scala 50:57:@43788.4]
  wire [10:0] _T_91241; // @[Modules.scala 50:57:@43789.4]
  wire [10:0] buffer_11_545; // @[Modules.scala 50:57:@43790.4]
  wire [10:0] buffer_11_310; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91246; // @[Modules.scala 50:57:@43796.4]
  wire [10:0] _T_91247; // @[Modules.scala 50:57:@43797.4]
  wire [10:0] buffer_11_547; // @[Modules.scala 50:57:@43798.4]
  wire [11:0] _T_91249; // @[Modules.scala 50:57:@43800.4]
  wire [10:0] _T_91250; // @[Modules.scala 50:57:@43801.4]
  wire [10:0] buffer_11_548; // @[Modules.scala 50:57:@43802.4]
  wire [11:0] _T_91261; // @[Modules.scala 50:57:@43816.4]
  wire [10:0] _T_91262; // @[Modules.scala 50:57:@43817.4]
  wire [10:0] buffer_11_552; // @[Modules.scala 50:57:@43818.4]
  wire [11:0] _T_91270; // @[Modules.scala 50:57:@43828.4]
  wire [10:0] _T_91271; // @[Modules.scala 50:57:@43829.4]
  wire [10:0] buffer_11_555; // @[Modules.scala 50:57:@43830.4]
  wire [11:0] _T_91285; // @[Modules.scala 50:57:@43848.4]
  wire [10:0] _T_91286; // @[Modules.scala 50:57:@43849.4]
  wire [10:0] buffer_11_560; // @[Modules.scala 50:57:@43850.4]
  wire [11:0] _T_91300; // @[Modules.scala 50:57:@43868.4]
  wire [10:0] _T_91301; // @[Modules.scala 50:57:@43869.4]
  wire [10:0] buffer_11_565; // @[Modules.scala 50:57:@43870.4]
  wire [11:0] _T_91303; // @[Modules.scala 50:57:@43872.4]
  wire [10:0] _T_91304; // @[Modules.scala 50:57:@43873.4]
  wire [10:0] buffer_11_566; // @[Modules.scala 50:57:@43874.4]
  wire [11:0] _T_91306; // @[Modules.scala 50:57:@43876.4]
  wire [10:0] _T_91307; // @[Modules.scala 50:57:@43877.4]
  wire [10:0] buffer_11_567; // @[Modules.scala 50:57:@43878.4]
  wire [10:0] buffer_11_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_91321; // @[Modules.scala 50:57:@43896.4]
  wire [10:0] _T_91322; // @[Modules.scala 50:57:@43897.4]
  wire [10:0] buffer_11_572; // @[Modules.scala 50:57:@43898.4]
  wire [11:0] _T_91348; // @[Modules.scala 50:57:@43932.4]
  wire [10:0] _T_91349; // @[Modules.scala 50:57:@43933.4]
  wire [10:0] buffer_11_581; // @[Modules.scala 50:57:@43934.4]
  wire [11:0] _T_91369; // @[Modules.scala 53:83:@43960.4]
  wire [10:0] _T_91370; // @[Modules.scala 53:83:@43961.4]
  wire [10:0] buffer_11_588; // @[Modules.scala 53:83:@43962.4]
  wire [11:0] _T_91372; // @[Modules.scala 53:83:@43964.4]
  wire [10:0] _T_91373; // @[Modules.scala 53:83:@43965.4]
  wire [10:0] buffer_11_589; // @[Modules.scala 53:83:@43966.4]
  wire [11:0] _T_91375; // @[Modules.scala 53:83:@43968.4]
  wire [10:0] _T_91376; // @[Modules.scala 53:83:@43969.4]
  wire [10:0] buffer_11_590; // @[Modules.scala 53:83:@43970.4]
  wire [11:0] _T_91378; // @[Modules.scala 53:83:@43972.4]
  wire [10:0] _T_91379; // @[Modules.scala 53:83:@43973.4]
  wire [10:0] buffer_11_591; // @[Modules.scala 53:83:@43974.4]
  wire [11:0] _T_91381; // @[Modules.scala 53:83:@43976.4]
  wire [10:0] _T_91382; // @[Modules.scala 53:83:@43977.4]
  wire [10:0] buffer_11_592; // @[Modules.scala 53:83:@43978.4]
  wire [11:0] _T_91384; // @[Modules.scala 53:83:@43980.4]
  wire [10:0] _T_91385; // @[Modules.scala 53:83:@43981.4]
  wire [10:0] buffer_11_593; // @[Modules.scala 53:83:@43982.4]
  wire [11:0] _T_91387; // @[Modules.scala 53:83:@43984.4]
  wire [10:0] _T_91388; // @[Modules.scala 53:83:@43985.4]
  wire [10:0] buffer_11_594; // @[Modules.scala 53:83:@43986.4]
  wire [11:0] _T_91390; // @[Modules.scala 53:83:@43988.4]
  wire [10:0] _T_91391; // @[Modules.scala 53:83:@43989.4]
  wire [10:0] buffer_11_595; // @[Modules.scala 53:83:@43990.4]
  wire [11:0] _T_91393; // @[Modules.scala 53:83:@43992.4]
  wire [10:0] _T_91394; // @[Modules.scala 53:83:@43993.4]
  wire [10:0] buffer_11_596; // @[Modules.scala 53:83:@43994.4]
  wire [11:0] _T_91399; // @[Modules.scala 53:83:@44000.4]
  wire [10:0] _T_91400; // @[Modules.scala 53:83:@44001.4]
  wire [10:0] buffer_11_598; // @[Modules.scala 53:83:@44002.4]
  wire [11:0] _T_91402; // @[Modules.scala 53:83:@44004.4]
  wire [10:0] _T_91403; // @[Modules.scala 53:83:@44005.4]
  wire [10:0] buffer_11_599; // @[Modules.scala 53:83:@44006.4]
  wire [11:0] _T_91414; // @[Modules.scala 53:83:@44020.4]
  wire [10:0] _T_91415; // @[Modules.scala 53:83:@44021.4]
  wire [10:0] buffer_11_603; // @[Modules.scala 53:83:@44022.4]
  wire [11:0] _T_91417; // @[Modules.scala 53:83:@44024.4]
  wire [10:0] _T_91418; // @[Modules.scala 53:83:@44025.4]
  wire [10:0] buffer_11_604; // @[Modules.scala 53:83:@44026.4]
  wire [11:0] _T_91420; // @[Modules.scala 53:83:@44028.4]
  wire [10:0] _T_91421; // @[Modules.scala 53:83:@44029.4]
  wire [10:0] buffer_11_605; // @[Modules.scala 53:83:@44030.4]
  wire [11:0] _T_91426; // @[Modules.scala 53:83:@44036.4]
  wire [10:0] _T_91427; // @[Modules.scala 53:83:@44037.4]
  wire [10:0] buffer_11_607; // @[Modules.scala 53:83:@44038.4]
  wire [11:0] _T_91429; // @[Modules.scala 53:83:@44040.4]
  wire [10:0] _T_91430; // @[Modules.scala 53:83:@44041.4]
  wire [10:0] buffer_11_608; // @[Modules.scala 53:83:@44042.4]
  wire [11:0] _T_91432; // @[Modules.scala 53:83:@44044.4]
  wire [10:0] _T_91433; // @[Modules.scala 53:83:@44045.4]
  wire [10:0] buffer_11_609; // @[Modules.scala 53:83:@44046.4]
  wire [11:0] _T_91435; // @[Modules.scala 53:83:@44048.4]
  wire [10:0] _T_91436; // @[Modules.scala 53:83:@44049.4]
  wire [10:0] buffer_11_610; // @[Modules.scala 53:83:@44050.4]
  wire [11:0] _T_91438; // @[Modules.scala 53:83:@44052.4]
  wire [10:0] _T_91439; // @[Modules.scala 53:83:@44053.4]
  wire [10:0] buffer_11_611; // @[Modules.scala 53:83:@44054.4]
  wire [11:0] _T_91441; // @[Modules.scala 53:83:@44056.4]
  wire [10:0] _T_91442; // @[Modules.scala 53:83:@44057.4]
  wire [10:0] buffer_11_612; // @[Modules.scala 53:83:@44058.4]
  wire [11:0] _T_91444; // @[Modules.scala 53:83:@44060.4]
  wire [10:0] _T_91445; // @[Modules.scala 53:83:@44061.4]
  wire [10:0] buffer_11_613; // @[Modules.scala 53:83:@44062.4]
  wire [11:0] _T_91447; // @[Modules.scala 53:83:@44064.4]
  wire [10:0] _T_91448; // @[Modules.scala 53:83:@44065.4]
  wire [10:0] buffer_11_614; // @[Modules.scala 53:83:@44066.4]
  wire [11:0] _T_91453; // @[Modules.scala 53:83:@44072.4]
  wire [10:0] _T_91454; // @[Modules.scala 53:83:@44073.4]
  wire [10:0] buffer_11_616; // @[Modules.scala 53:83:@44074.4]
  wire [11:0] _T_91456; // @[Modules.scala 53:83:@44076.4]
  wire [10:0] _T_91457; // @[Modules.scala 53:83:@44077.4]
  wire [10:0] buffer_11_617; // @[Modules.scala 53:83:@44078.4]
  wire [11:0] _T_91459; // @[Modules.scala 53:83:@44080.4]
  wire [10:0] _T_91460; // @[Modules.scala 53:83:@44081.4]
  wire [10:0] buffer_11_618; // @[Modules.scala 53:83:@44082.4]
  wire [11:0] _T_91462; // @[Modules.scala 53:83:@44084.4]
  wire [10:0] _T_91463; // @[Modules.scala 53:83:@44085.4]
  wire [10:0] buffer_11_619; // @[Modules.scala 53:83:@44086.4]
  wire [11:0] _T_91465; // @[Modules.scala 53:83:@44088.4]
  wire [10:0] _T_91466; // @[Modules.scala 53:83:@44089.4]
  wire [10:0] buffer_11_620; // @[Modules.scala 53:83:@44090.4]
  wire [11:0] _T_91468; // @[Modules.scala 53:83:@44092.4]
  wire [10:0] _T_91469; // @[Modules.scala 53:83:@44093.4]
  wire [10:0] buffer_11_621; // @[Modules.scala 53:83:@44094.4]
  wire [11:0] _T_91474; // @[Modules.scala 53:83:@44100.4]
  wire [10:0] _T_91475; // @[Modules.scala 53:83:@44101.4]
  wire [10:0] buffer_11_623; // @[Modules.scala 53:83:@44102.4]
  wire [11:0] _T_91477; // @[Modules.scala 53:83:@44104.4]
  wire [10:0] _T_91478; // @[Modules.scala 53:83:@44105.4]
  wire [10:0] buffer_11_624; // @[Modules.scala 53:83:@44106.4]
  wire [11:0] _T_91486; // @[Modules.scala 53:83:@44116.4]
  wire [10:0] _T_91487; // @[Modules.scala 53:83:@44117.4]
  wire [10:0] buffer_11_627; // @[Modules.scala 53:83:@44118.4]
  wire [11:0] _T_91489; // @[Modules.scala 53:83:@44120.4]
  wire [10:0] _T_91490; // @[Modules.scala 53:83:@44121.4]
  wire [10:0] buffer_11_628; // @[Modules.scala 53:83:@44122.4]
  wire [11:0] _T_91501; // @[Modules.scala 53:83:@44136.4]
  wire [10:0] _T_91502; // @[Modules.scala 53:83:@44137.4]
  wire [10:0] buffer_11_632; // @[Modules.scala 53:83:@44138.4]
  wire [11:0] _T_91504; // @[Modules.scala 53:83:@44140.4]
  wire [10:0] _T_91505; // @[Modules.scala 53:83:@44141.4]
  wire [10:0] buffer_11_633; // @[Modules.scala 53:83:@44142.4]
  wire [11:0] _T_91507; // @[Modules.scala 53:83:@44144.4]
  wire [10:0] _T_91508; // @[Modules.scala 53:83:@44145.4]
  wire [10:0] buffer_11_634; // @[Modules.scala 53:83:@44146.4]
  wire [11:0] _T_91510; // @[Modules.scala 53:83:@44148.4]
  wire [10:0] _T_91511; // @[Modules.scala 53:83:@44149.4]
  wire [10:0] buffer_11_635; // @[Modules.scala 53:83:@44150.4]
  wire [11:0] _T_91513; // @[Modules.scala 53:83:@44152.4]
  wire [10:0] _T_91514; // @[Modules.scala 53:83:@44153.4]
  wire [10:0] buffer_11_636; // @[Modules.scala 53:83:@44154.4]
  wire [11:0] _T_91519; // @[Modules.scala 53:83:@44160.4]
  wire [10:0] _T_91520; // @[Modules.scala 53:83:@44161.4]
  wire [10:0] buffer_11_638; // @[Modules.scala 53:83:@44162.4]
  wire [11:0] _T_91522; // @[Modules.scala 53:83:@44164.4]
  wire [10:0] _T_91523; // @[Modules.scala 53:83:@44165.4]
  wire [10:0] buffer_11_639; // @[Modules.scala 53:83:@44166.4]
  wire [11:0] _T_91525; // @[Modules.scala 53:83:@44168.4]
  wire [10:0] _T_91526; // @[Modules.scala 53:83:@44169.4]
  wire [10:0] buffer_11_640; // @[Modules.scala 53:83:@44170.4]
  wire [11:0] _T_91528; // @[Modules.scala 53:83:@44172.4]
  wire [10:0] _T_91529; // @[Modules.scala 53:83:@44173.4]
  wire [10:0] buffer_11_641; // @[Modules.scala 53:83:@44174.4]
  wire [11:0] _T_91531; // @[Modules.scala 53:83:@44176.4]
  wire [10:0] _T_91532; // @[Modules.scala 53:83:@44177.4]
  wire [10:0] buffer_11_642; // @[Modules.scala 53:83:@44178.4]
  wire [11:0] _T_91534; // @[Modules.scala 53:83:@44180.4]
  wire [10:0] _T_91535; // @[Modules.scala 53:83:@44181.4]
  wire [10:0] buffer_11_643; // @[Modules.scala 53:83:@44182.4]
  wire [11:0] _T_91537; // @[Modules.scala 53:83:@44184.4]
  wire [10:0] _T_91538; // @[Modules.scala 53:83:@44185.4]
  wire [10:0] buffer_11_644; // @[Modules.scala 53:83:@44186.4]
  wire [11:0] _T_91540; // @[Modules.scala 53:83:@44188.4]
  wire [10:0] _T_91541; // @[Modules.scala 53:83:@44189.4]
  wire [10:0] buffer_11_645; // @[Modules.scala 53:83:@44190.4]
  wire [11:0] _T_91543; // @[Modules.scala 53:83:@44192.4]
  wire [10:0] _T_91544; // @[Modules.scala 53:83:@44193.4]
  wire [10:0] buffer_11_646; // @[Modules.scala 53:83:@44194.4]
  wire [11:0] _T_91546; // @[Modules.scala 53:83:@44196.4]
  wire [10:0] _T_91547; // @[Modules.scala 53:83:@44197.4]
  wire [10:0] buffer_11_647; // @[Modules.scala 53:83:@44198.4]
  wire [11:0] _T_91549; // @[Modules.scala 53:83:@44200.4]
  wire [10:0] _T_91550; // @[Modules.scala 53:83:@44201.4]
  wire [10:0] buffer_11_648; // @[Modules.scala 53:83:@44202.4]
  wire [11:0] _T_91552; // @[Modules.scala 53:83:@44204.4]
  wire [10:0] _T_91553; // @[Modules.scala 53:83:@44205.4]
  wire [10:0] buffer_11_649; // @[Modules.scala 53:83:@44206.4]
  wire [11:0] _T_91555; // @[Modules.scala 53:83:@44208.4]
  wire [10:0] _T_91556; // @[Modules.scala 53:83:@44209.4]
  wire [10:0] buffer_11_650; // @[Modules.scala 53:83:@44210.4]
  wire [11:0] _T_91558; // @[Modules.scala 53:83:@44212.4]
  wire [10:0] _T_91559; // @[Modules.scala 53:83:@44213.4]
  wire [10:0] buffer_11_651; // @[Modules.scala 53:83:@44214.4]
  wire [11:0] _T_91561; // @[Modules.scala 53:83:@44216.4]
  wire [10:0] _T_91562; // @[Modules.scala 53:83:@44217.4]
  wire [10:0] buffer_11_652; // @[Modules.scala 53:83:@44218.4]
  wire [11:0] _T_91564; // @[Modules.scala 53:83:@44220.4]
  wire [10:0] _T_91565; // @[Modules.scala 53:83:@44221.4]
  wire [10:0] buffer_11_653; // @[Modules.scala 53:83:@44222.4]
  wire [11:0] _T_91570; // @[Modules.scala 53:83:@44228.4]
  wire [10:0] _T_91571; // @[Modules.scala 53:83:@44229.4]
  wire [10:0] buffer_11_655; // @[Modules.scala 53:83:@44230.4]
  wire [11:0] _T_91573; // @[Modules.scala 53:83:@44232.4]
  wire [10:0] _T_91574; // @[Modules.scala 53:83:@44233.4]
  wire [10:0] buffer_11_656; // @[Modules.scala 53:83:@44234.4]
  wire [11:0] _T_91576; // @[Modules.scala 53:83:@44236.4]
  wire [10:0] _T_91577; // @[Modules.scala 53:83:@44237.4]
  wire [10:0] buffer_11_657; // @[Modules.scala 53:83:@44238.4]
  wire [11:0] _T_91579; // @[Modules.scala 53:83:@44240.4]
  wire [10:0] _T_91580; // @[Modules.scala 53:83:@44241.4]
  wire [10:0] buffer_11_658; // @[Modules.scala 53:83:@44242.4]
  wire [11:0] _T_91582; // @[Modules.scala 53:83:@44244.4]
  wire [10:0] _T_91583; // @[Modules.scala 53:83:@44245.4]
  wire [10:0] buffer_11_659; // @[Modules.scala 53:83:@44246.4]
  wire [11:0] _T_91585; // @[Modules.scala 53:83:@44248.4]
  wire [10:0] _T_91586; // @[Modules.scala 53:83:@44249.4]
  wire [10:0] buffer_11_660; // @[Modules.scala 53:83:@44250.4]
  wire [11:0] _T_91588; // @[Modules.scala 53:83:@44252.4]
  wire [10:0] _T_91589; // @[Modules.scala 53:83:@44253.4]
  wire [10:0] buffer_11_661; // @[Modules.scala 53:83:@44254.4]
  wire [11:0] _T_91591; // @[Modules.scala 53:83:@44256.4]
  wire [10:0] _T_91592; // @[Modules.scala 53:83:@44257.4]
  wire [10:0] buffer_11_662; // @[Modules.scala 53:83:@44258.4]
  wire [11:0] _T_91594; // @[Modules.scala 53:83:@44260.4]
  wire [10:0] _T_91595; // @[Modules.scala 53:83:@44261.4]
  wire [10:0] buffer_11_663; // @[Modules.scala 53:83:@44262.4]
  wire [11:0] _T_91597; // @[Modules.scala 53:83:@44264.4]
  wire [10:0] _T_91598; // @[Modules.scala 53:83:@44265.4]
  wire [10:0] buffer_11_664; // @[Modules.scala 53:83:@44266.4]
  wire [11:0] _T_91600; // @[Modules.scala 53:83:@44268.4]
  wire [10:0] _T_91601; // @[Modules.scala 53:83:@44269.4]
  wire [10:0] buffer_11_665; // @[Modules.scala 53:83:@44270.4]
  wire [11:0] _T_91603; // @[Modules.scala 53:83:@44272.4]
  wire [10:0] _T_91604; // @[Modules.scala 53:83:@44273.4]
  wire [10:0] buffer_11_666; // @[Modules.scala 53:83:@44274.4]
  wire [11:0] _T_91609; // @[Modules.scala 53:83:@44280.4]
  wire [10:0] _T_91610; // @[Modules.scala 53:83:@44281.4]
  wire [10:0] buffer_11_668; // @[Modules.scala 53:83:@44282.4]
  wire [11:0] _T_91612; // @[Modules.scala 53:83:@44284.4]
  wire [10:0] _T_91613; // @[Modules.scala 53:83:@44285.4]
  wire [10:0] buffer_11_669; // @[Modules.scala 53:83:@44286.4]
  wire [11:0] _T_91615; // @[Modules.scala 53:83:@44288.4]
  wire [10:0] _T_91616; // @[Modules.scala 53:83:@44289.4]
  wire [10:0] buffer_11_670; // @[Modules.scala 53:83:@44290.4]
  wire [11:0] _T_91618; // @[Modules.scala 53:83:@44292.4]
  wire [10:0] _T_91619; // @[Modules.scala 53:83:@44293.4]
  wire [10:0] buffer_11_671; // @[Modules.scala 53:83:@44294.4]
  wire [11:0] _T_91621; // @[Modules.scala 53:83:@44296.4]
  wire [10:0] _T_91622; // @[Modules.scala 53:83:@44297.4]
  wire [10:0] buffer_11_672; // @[Modules.scala 53:83:@44298.4]
  wire [11:0] _T_91627; // @[Modules.scala 53:83:@44304.4]
  wire [10:0] _T_91628; // @[Modules.scala 53:83:@44305.4]
  wire [10:0] buffer_11_674; // @[Modules.scala 53:83:@44306.4]
  wire [11:0] _T_91630; // @[Modules.scala 53:83:@44308.4]
  wire [10:0] _T_91631; // @[Modules.scala 53:83:@44309.4]
  wire [10:0] buffer_11_675; // @[Modules.scala 53:83:@44310.4]
  wire [11:0] _T_91639; // @[Modules.scala 53:83:@44320.4]
  wire [10:0] _T_91640; // @[Modules.scala 53:83:@44321.4]
  wire [10:0] buffer_11_678; // @[Modules.scala 53:83:@44322.4]
  wire [11:0] _T_91651; // @[Modules.scala 53:83:@44336.4]
  wire [10:0] _T_91652; // @[Modules.scala 53:83:@44337.4]
  wire [10:0] buffer_11_682; // @[Modules.scala 53:83:@44338.4]
  wire [11:0] _T_91663; // @[Modules.scala 56:109:@44352.4]
  wire [10:0] _T_91664; // @[Modules.scala 56:109:@44353.4]
  wire [10:0] buffer_11_686; // @[Modules.scala 56:109:@44354.4]
  wire [11:0] _T_91666; // @[Modules.scala 56:109:@44356.4]
  wire [10:0] _T_91667; // @[Modules.scala 56:109:@44357.4]
  wire [10:0] buffer_11_687; // @[Modules.scala 56:109:@44358.4]
  wire [11:0] _T_91669; // @[Modules.scala 56:109:@44360.4]
  wire [10:0] _T_91670; // @[Modules.scala 56:109:@44361.4]
  wire [10:0] buffer_11_688; // @[Modules.scala 56:109:@44362.4]
  wire [11:0] _T_91672; // @[Modules.scala 56:109:@44364.4]
  wire [10:0] _T_91673; // @[Modules.scala 56:109:@44365.4]
  wire [10:0] buffer_11_689; // @[Modules.scala 56:109:@44366.4]
  wire [11:0] _T_91675; // @[Modules.scala 56:109:@44368.4]
  wire [10:0] _T_91676; // @[Modules.scala 56:109:@44369.4]
  wire [10:0] buffer_11_690; // @[Modules.scala 56:109:@44370.4]
  wire [11:0] _T_91678; // @[Modules.scala 56:109:@44372.4]
  wire [10:0] _T_91679; // @[Modules.scala 56:109:@44373.4]
  wire [10:0] buffer_11_691; // @[Modules.scala 56:109:@44374.4]
  wire [11:0] _T_91684; // @[Modules.scala 56:109:@44380.4]
  wire [10:0] _T_91685; // @[Modules.scala 56:109:@44381.4]
  wire [10:0] buffer_11_693; // @[Modules.scala 56:109:@44382.4]
  wire [11:0] _T_91687; // @[Modules.scala 56:109:@44384.4]
  wire [10:0] _T_91688; // @[Modules.scala 56:109:@44385.4]
  wire [10:0] buffer_11_694; // @[Modules.scala 56:109:@44386.4]
  wire [11:0] _T_91690; // @[Modules.scala 56:109:@44388.4]
  wire [10:0] _T_91691; // @[Modules.scala 56:109:@44389.4]
  wire [10:0] buffer_11_695; // @[Modules.scala 56:109:@44390.4]
  wire [11:0] _T_91693; // @[Modules.scala 56:109:@44392.4]
  wire [10:0] _T_91694; // @[Modules.scala 56:109:@44393.4]
  wire [10:0] buffer_11_696; // @[Modules.scala 56:109:@44394.4]
  wire [11:0] _T_91696; // @[Modules.scala 56:109:@44396.4]
  wire [10:0] _T_91697; // @[Modules.scala 56:109:@44397.4]
  wire [10:0] buffer_11_697; // @[Modules.scala 56:109:@44398.4]
  wire [11:0] _T_91699; // @[Modules.scala 56:109:@44400.4]
  wire [10:0] _T_91700; // @[Modules.scala 56:109:@44401.4]
  wire [10:0] buffer_11_698; // @[Modules.scala 56:109:@44402.4]
  wire [11:0] _T_91702; // @[Modules.scala 56:109:@44404.4]
  wire [10:0] _T_91703; // @[Modules.scala 56:109:@44405.4]
  wire [10:0] buffer_11_699; // @[Modules.scala 56:109:@44406.4]
  wire [11:0] _T_91705; // @[Modules.scala 56:109:@44408.4]
  wire [10:0] _T_91706; // @[Modules.scala 56:109:@44409.4]
  wire [10:0] buffer_11_700; // @[Modules.scala 56:109:@44410.4]
  wire [11:0] _T_91708; // @[Modules.scala 56:109:@44412.4]
  wire [10:0] _T_91709; // @[Modules.scala 56:109:@44413.4]
  wire [10:0] buffer_11_701; // @[Modules.scala 56:109:@44414.4]
  wire [11:0] _T_91711; // @[Modules.scala 56:109:@44416.4]
  wire [10:0] _T_91712; // @[Modules.scala 56:109:@44417.4]
  wire [10:0] buffer_11_702; // @[Modules.scala 56:109:@44418.4]
  wire [11:0] _T_91714; // @[Modules.scala 56:109:@44420.4]
  wire [10:0] _T_91715; // @[Modules.scala 56:109:@44421.4]
  wire [10:0] buffer_11_703; // @[Modules.scala 56:109:@44422.4]
  wire [11:0] _T_91717; // @[Modules.scala 56:109:@44424.4]
  wire [10:0] _T_91718; // @[Modules.scala 56:109:@44425.4]
  wire [10:0] buffer_11_704; // @[Modules.scala 56:109:@44426.4]
  wire [11:0] _T_91720; // @[Modules.scala 56:109:@44428.4]
  wire [10:0] _T_91721; // @[Modules.scala 56:109:@44429.4]
  wire [10:0] buffer_11_705; // @[Modules.scala 56:109:@44430.4]
  wire [11:0] _T_91723; // @[Modules.scala 56:109:@44432.4]
  wire [10:0] _T_91724; // @[Modules.scala 56:109:@44433.4]
  wire [10:0] buffer_11_706; // @[Modules.scala 56:109:@44434.4]
  wire [11:0] _T_91729; // @[Modules.scala 56:109:@44440.4]
  wire [10:0] _T_91730; // @[Modules.scala 56:109:@44441.4]
  wire [10:0] buffer_11_708; // @[Modules.scala 56:109:@44442.4]
  wire [11:0] _T_91732; // @[Modules.scala 56:109:@44444.4]
  wire [10:0] _T_91733; // @[Modules.scala 56:109:@44445.4]
  wire [10:0] buffer_11_709; // @[Modules.scala 56:109:@44446.4]
  wire [11:0] _T_91735; // @[Modules.scala 56:109:@44448.4]
  wire [10:0] _T_91736; // @[Modules.scala 56:109:@44449.4]
  wire [10:0] buffer_11_710; // @[Modules.scala 56:109:@44450.4]
  wire [11:0] _T_91738; // @[Modules.scala 56:109:@44452.4]
  wire [10:0] _T_91739; // @[Modules.scala 56:109:@44453.4]
  wire [10:0] buffer_11_711; // @[Modules.scala 56:109:@44454.4]
  wire [11:0] _T_91741; // @[Modules.scala 56:109:@44456.4]
  wire [10:0] _T_91742; // @[Modules.scala 56:109:@44457.4]
  wire [10:0] buffer_11_712; // @[Modules.scala 56:109:@44458.4]
  wire [11:0] _T_91744; // @[Modules.scala 56:109:@44460.4]
  wire [10:0] _T_91745; // @[Modules.scala 56:109:@44461.4]
  wire [10:0] buffer_11_713; // @[Modules.scala 56:109:@44462.4]
  wire [11:0] _T_91747; // @[Modules.scala 56:109:@44464.4]
  wire [10:0] _T_91748; // @[Modules.scala 56:109:@44465.4]
  wire [10:0] buffer_11_714; // @[Modules.scala 56:109:@44466.4]
  wire [11:0] _T_91750; // @[Modules.scala 56:109:@44468.4]
  wire [10:0] _T_91751; // @[Modules.scala 56:109:@44469.4]
  wire [10:0] buffer_11_715; // @[Modules.scala 56:109:@44470.4]
  wire [11:0] _T_91753; // @[Modules.scala 56:109:@44472.4]
  wire [10:0] _T_91754; // @[Modules.scala 56:109:@44473.4]
  wire [10:0] buffer_11_716; // @[Modules.scala 56:109:@44474.4]
  wire [11:0] _T_91756; // @[Modules.scala 56:109:@44476.4]
  wire [10:0] _T_91757; // @[Modules.scala 56:109:@44477.4]
  wire [10:0] buffer_11_717; // @[Modules.scala 56:109:@44478.4]
  wire [11:0] _T_91759; // @[Modules.scala 56:109:@44480.4]
  wire [10:0] _T_91760; // @[Modules.scala 56:109:@44481.4]
  wire [10:0] buffer_11_718; // @[Modules.scala 56:109:@44482.4]
  wire [11:0] _T_91762; // @[Modules.scala 56:109:@44484.4]
  wire [10:0] _T_91763; // @[Modules.scala 56:109:@44485.4]
  wire [10:0] buffer_11_719; // @[Modules.scala 56:109:@44486.4]
  wire [11:0] _T_91765; // @[Modules.scala 56:109:@44488.4]
  wire [10:0] _T_91766; // @[Modules.scala 56:109:@44489.4]
  wire [10:0] buffer_11_720; // @[Modules.scala 56:109:@44490.4]
  wire [11:0] _T_91768; // @[Modules.scala 56:109:@44492.4]
  wire [10:0] _T_91769; // @[Modules.scala 56:109:@44493.4]
  wire [10:0] buffer_11_721; // @[Modules.scala 56:109:@44494.4]
  wire [11:0] _T_91771; // @[Modules.scala 56:109:@44496.4]
  wire [10:0] _T_91772; // @[Modules.scala 56:109:@44497.4]
  wire [10:0] buffer_11_722; // @[Modules.scala 56:109:@44498.4]
  wire [11:0] _T_91774; // @[Modules.scala 56:109:@44500.4]
  wire [10:0] _T_91775; // @[Modules.scala 56:109:@44501.4]
  wire [10:0] buffer_11_723; // @[Modules.scala 56:109:@44502.4]
  wire [11:0] _T_91777; // @[Modules.scala 56:109:@44504.4]
  wire [10:0] _T_91778; // @[Modules.scala 56:109:@44505.4]
  wire [10:0] buffer_11_724; // @[Modules.scala 56:109:@44506.4]
  wire [11:0] _T_91780; // @[Modules.scala 56:109:@44508.4]
  wire [10:0] _T_91781; // @[Modules.scala 56:109:@44509.4]
  wire [10:0] buffer_11_725; // @[Modules.scala 56:109:@44510.4]
  wire [11:0] _T_91783; // @[Modules.scala 56:109:@44512.4]
  wire [10:0] _T_91784; // @[Modules.scala 56:109:@44513.4]
  wire [10:0] buffer_11_726; // @[Modules.scala 56:109:@44514.4]
  wire [11:0] _T_91786; // @[Modules.scala 56:109:@44516.4]
  wire [10:0] _T_91787; // @[Modules.scala 56:109:@44517.4]
  wire [10:0] buffer_11_727; // @[Modules.scala 56:109:@44518.4]
  wire [11:0] _T_91789; // @[Modules.scala 56:109:@44520.4]
  wire [10:0] _T_91790; // @[Modules.scala 56:109:@44521.4]
  wire [10:0] buffer_11_728; // @[Modules.scala 56:109:@44522.4]
  wire [11:0] _T_91792; // @[Modules.scala 56:109:@44524.4]
  wire [10:0] _T_91793; // @[Modules.scala 56:109:@44525.4]
  wire [10:0] buffer_11_729; // @[Modules.scala 56:109:@44526.4]
  wire [11:0] _T_91798; // @[Modules.scala 56:109:@44532.4]
  wire [10:0] _T_91799; // @[Modules.scala 56:109:@44533.4]
  wire [10:0] buffer_11_731; // @[Modules.scala 56:109:@44534.4]
  wire [11:0] _T_91804; // @[Modules.scala 56:109:@44540.4]
  wire [10:0] _T_91805; // @[Modules.scala 56:109:@44541.4]
  wire [10:0] buffer_11_733; // @[Modules.scala 56:109:@44542.4]
  wire [11:0] _T_91810; // @[Modules.scala 63:156:@44549.4]
  wire [10:0] _T_91811; // @[Modules.scala 63:156:@44550.4]
  wire [10:0] buffer_11_736; // @[Modules.scala 63:156:@44551.4]
  wire [11:0] _T_91813; // @[Modules.scala 63:156:@44553.4]
  wire [10:0] _T_91814; // @[Modules.scala 63:156:@44554.4]
  wire [10:0] buffer_11_737; // @[Modules.scala 63:156:@44555.4]
  wire [11:0] _T_91816; // @[Modules.scala 63:156:@44557.4]
  wire [10:0] _T_91817; // @[Modules.scala 63:156:@44558.4]
  wire [10:0] buffer_11_738; // @[Modules.scala 63:156:@44559.4]
  wire [11:0] _T_91819; // @[Modules.scala 63:156:@44561.4]
  wire [10:0] _T_91820; // @[Modules.scala 63:156:@44562.4]
  wire [10:0] buffer_11_739; // @[Modules.scala 63:156:@44563.4]
  wire [11:0] _T_91822; // @[Modules.scala 63:156:@44565.4]
  wire [10:0] _T_91823; // @[Modules.scala 63:156:@44566.4]
  wire [10:0] buffer_11_740; // @[Modules.scala 63:156:@44567.4]
  wire [11:0] _T_91825; // @[Modules.scala 63:156:@44569.4]
  wire [10:0] _T_91826; // @[Modules.scala 63:156:@44570.4]
  wire [10:0] buffer_11_741; // @[Modules.scala 63:156:@44571.4]
  wire [11:0] _T_91828; // @[Modules.scala 63:156:@44573.4]
  wire [10:0] _T_91829; // @[Modules.scala 63:156:@44574.4]
  wire [10:0] buffer_11_742; // @[Modules.scala 63:156:@44575.4]
  wire [11:0] _T_91831; // @[Modules.scala 63:156:@44577.4]
  wire [10:0] _T_91832; // @[Modules.scala 63:156:@44578.4]
  wire [10:0] buffer_11_743; // @[Modules.scala 63:156:@44579.4]
  wire [11:0] _T_91834; // @[Modules.scala 63:156:@44581.4]
  wire [10:0] _T_91835; // @[Modules.scala 63:156:@44582.4]
  wire [10:0] buffer_11_744; // @[Modules.scala 63:156:@44583.4]
  wire [11:0] _T_91837; // @[Modules.scala 63:156:@44585.4]
  wire [10:0] _T_91838; // @[Modules.scala 63:156:@44586.4]
  wire [10:0] buffer_11_745; // @[Modules.scala 63:156:@44587.4]
  wire [11:0] _T_91840; // @[Modules.scala 63:156:@44589.4]
  wire [10:0] _T_91841; // @[Modules.scala 63:156:@44590.4]
  wire [10:0] buffer_11_746; // @[Modules.scala 63:156:@44591.4]
  wire [11:0] _T_91843; // @[Modules.scala 63:156:@44593.4]
  wire [10:0] _T_91844; // @[Modules.scala 63:156:@44594.4]
  wire [10:0] buffer_11_747; // @[Modules.scala 63:156:@44595.4]
  wire [11:0] _T_91846; // @[Modules.scala 63:156:@44597.4]
  wire [10:0] _T_91847; // @[Modules.scala 63:156:@44598.4]
  wire [10:0] buffer_11_748; // @[Modules.scala 63:156:@44599.4]
  wire [11:0] _T_91849; // @[Modules.scala 63:156:@44601.4]
  wire [10:0] _T_91850; // @[Modules.scala 63:156:@44602.4]
  wire [10:0] buffer_11_749; // @[Modules.scala 63:156:@44603.4]
  wire [11:0] _T_91852; // @[Modules.scala 63:156:@44605.4]
  wire [10:0] _T_91853; // @[Modules.scala 63:156:@44606.4]
  wire [10:0] buffer_11_750; // @[Modules.scala 63:156:@44607.4]
  wire [11:0] _T_91855; // @[Modules.scala 63:156:@44609.4]
  wire [10:0] _T_91856; // @[Modules.scala 63:156:@44610.4]
  wire [10:0] buffer_11_751; // @[Modules.scala 63:156:@44611.4]
  wire [11:0] _T_91858; // @[Modules.scala 63:156:@44613.4]
  wire [10:0] _T_91859; // @[Modules.scala 63:156:@44614.4]
  wire [10:0] buffer_11_752; // @[Modules.scala 63:156:@44615.4]
  wire [11:0] _T_91861; // @[Modules.scala 63:156:@44617.4]
  wire [10:0] _T_91862; // @[Modules.scala 63:156:@44618.4]
  wire [10:0] buffer_11_753; // @[Modules.scala 63:156:@44619.4]
  wire [11:0] _T_91864; // @[Modules.scala 63:156:@44621.4]
  wire [10:0] _T_91865; // @[Modules.scala 63:156:@44622.4]
  wire [10:0] buffer_11_754; // @[Modules.scala 63:156:@44623.4]
  wire [11:0] _T_91867; // @[Modules.scala 63:156:@44625.4]
  wire [10:0] _T_91868; // @[Modules.scala 63:156:@44626.4]
  wire [10:0] buffer_11_755; // @[Modules.scala 63:156:@44627.4]
  wire [11:0] _T_91870; // @[Modules.scala 63:156:@44629.4]
  wire [10:0] _T_91871; // @[Modules.scala 63:156:@44630.4]
  wire [10:0] buffer_11_756; // @[Modules.scala 63:156:@44631.4]
  wire [11:0] _T_91873; // @[Modules.scala 63:156:@44633.4]
  wire [10:0] _T_91874; // @[Modules.scala 63:156:@44634.4]
  wire [10:0] buffer_11_757; // @[Modules.scala 63:156:@44635.4]
  wire [11:0] _T_91876; // @[Modules.scala 63:156:@44637.4]
  wire [10:0] _T_91877; // @[Modules.scala 63:156:@44638.4]
  wire [10:0] buffer_11_758; // @[Modules.scala 63:156:@44639.4]
  wire [11:0] _T_91879; // @[Modules.scala 63:156:@44641.4]
  wire [10:0] _T_91880; // @[Modules.scala 63:156:@44642.4]
  wire [10:0] buffer_11_759; // @[Modules.scala 63:156:@44643.4]
  wire [11:0] _T_91882; // @[Modules.scala 63:156:@44645.4]
  wire [10:0] _T_91883; // @[Modules.scala 63:156:@44646.4]
  wire [10:0] buffer_11_760; // @[Modules.scala 63:156:@44647.4]
  wire [11:0] _T_91885; // @[Modules.scala 63:156:@44649.4]
  wire [10:0] _T_91886; // @[Modules.scala 63:156:@44650.4]
  wire [10:0] buffer_11_761; // @[Modules.scala 63:156:@44651.4]
  wire [11:0] _T_91888; // @[Modules.scala 63:156:@44653.4]
  wire [10:0] _T_91889; // @[Modules.scala 63:156:@44654.4]
  wire [10:0] buffer_11_762; // @[Modules.scala 63:156:@44655.4]
  wire [11:0] _T_91891; // @[Modules.scala 63:156:@44657.4]
  wire [10:0] _T_91892; // @[Modules.scala 63:156:@44658.4]
  wire [10:0] buffer_11_763; // @[Modules.scala 63:156:@44659.4]
  wire [11:0] _T_91894; // @[Modules.scala 63:156:@44661.4]
  wire [10:0] _T_91895; // @[Modules.scala 63:156:@44662.4]
  wire [10:0] buffer_11_764; // @[Modules.scala 63:156:@44663.4]
  wire [11:0] _T_91897; // @[Modules.scala 63:156:@44665.4]
  wire [10:0] _T_91898; // @[Modules.scala 63:156:@44666.4]
  wire [10:0] buffer_11_765; // @[Modules.scala 63:156:@44667.4]
  wire [11:0] _T_91900; // @[Modules.scala 63:156:@44669.4]
  wire [10:0] _T_91901; // @[Modules.scala 63:156:@44670.4]
  wire [10:0] buffer_11_766; // @[Modules.scala 63:156:@44671.4]
  wire [11:0] _T_91903; // @[Modules.scala 63:156:@44673.4]
  wire [10:0] _T_91904; // @[Modules.scala 63:156:@44674.4]
  wire [10:0] buffer_11_767; // @[Modules.scala 63:156:@44675.4]
  wire [11:0] _T_91906; // @[Modules.scala 63:156:@44677.4]
  wire [10:0] _T_91907; // @[Modules.scala 63:156:@44678.4]
  wire [10:0] buffer_11_768; // @[Modules.scala 63:156:@44679.4]
  wire [11:0] _T_91909; // @[Modules.scala 63:156:@44681.4]
  wire [10:0] _T_91910; // @[Modules.scala 63:156:@44682.4]
  wire [10:0] buffer_11_769; // @[Modules.scala 63:156:@44683.4]
  wire [11:0] _T_91912; // @[Modules.scala 63:156:@44685.4]
  wire [10:0] _T_91913; // @[Modules.scala 63:156:@44686.4]
  wire [10:0] buffer_11_770; // @[Modules.scala 63:156:@44687.4]
  wire [11:0] _T_91915; // @[Modules.scala 63:156:@44689.4]
  wire [10:0] _T_91916; // @[Modules.scala 63:156:@44690.4]
  wire [10:0] buffer_11_771; // @[Modules.scala 63:156:@44691.4]
  wire [11:0] _T_91918; // @[Modules.scala 63:156:@44693.4]
  wire [10:0] _T_91919; // @[Modules.scala 63:156:@44694.4]
  wire [10:0] buffer_11_772; // @[Modules.scala 63:156:@44695.4]
  wire [11:0] _T_91921; // @[Modules.scala 63:156:@44697.4]
  wire [10:0] _T_91922; // @[Modules.scala 63:156:@44698.4]
  wire [10:0] buffer_11_773; // @[Modules.scala 63:156:@44699.4]
  wire [11:0] _T_91924; // @[Modules.scala 63:156:@44701.4]
  wire [10:0] _T_91925; // @[Modules.scala 63:156:@44702.4]
  wire [10:0] buffer_11_774; // @[Modules.scala 63:156:@44703.4]
  wire [11:0] _T_91927; // @[Modules.scala 63:156:@44705.4]
  wire [10:0] _T_91928; // @[Modules.scala 63:156:@44706.4]
  wire [10:0] buffer_11_775; // @[Modules.scala 63:156:@44707.4]
  wire [11:0] _T_91930; // @[Modules.scala 63:156:@44709.4]
  wire [10:0] _T_91931; // @[Modules.scala 63:156:@44710.4]
  wire [10:0] buffer_11_776; // @[Modules.scala 63:156:@44711.4]
  wire [11:0] _T_91933; // @[Modules.scala 63:156:@44713.4]
  wire [10:0] _T_91934; // @[Modules.scala 63:156:@44714.4]
  wire [10:0] buffer_11_777; // @[Modules.scala 63:156:@44715.4]
  wire [11:0] _T_91936; // @[Modules.scala 63:156:@44717.4]
  wire [10:0] _T_91937; // @[Modules.scala 63:156:@44718.4]
  wire [10:0] buffer_11_778; // @[Modules.scala 63:156:@44719.4]
  wire [11:0] _T_91939; // @[Modules.scala 63:156:@44721.4]
  wire [10:0] _T_91940; // @[Modules.scala 63:156:@44722.4]
  wire [10:0] buffer_11_779; // @[Modules.scala 63:156:@44723.4]
  wire [11:0] _T_91942; // @[Modules.scala 63:156:@44725.4]
  wire [10:0] _T_91943; // @[Modules.scala 63:156:@44726.4]
  wire [10:0] buffer_11_780; // @[Modules.scala 63:156:@44727.4]
  wire [11:0] _T_91945; // @[Modules.scala 63:156:@44729.4]
  wire [10:0] _T_91946; // @[Modules.scala 63:156:@44730.4]
  wire [10:0] buffer_11_781; // @[Modules.scala 63:156:@44731.4]
  wire [11:0] _T_91948; // @[Modules.scala 63:156:@44733.4]
  wire [10:0] _T_91949; // @[Modules.scala 63:156:@44734.4]
  wire [10:0] buffer_11_782; // @[Modules.scala 63:156:@44735.4]
  wire [11:0] _T_91951; // @[Modules.scala 63:156:@44737.4]
  wire [10:0] _T_91952; // @[Modules.scala 63:156:@44738.4]
  wire [10:0] buffer_11_783; // @[Modules.scala 63:156:@44739.4]
  wire [5:0] _T_91991; // @[Modules.scala 40:46:@44782.4]
  wire [4:0] _T_91992; // @[Modules.scala 40:46:@44783.4]
  wire [4:0] _T_91993; // @[Modules.scala 40:46:@44784.4]
  wire [5:0] _T_92493; // @[Modules.scala 40:46:@45344.4]
  wire [4:0] _T_92494; // @[Modules.scala 40:46:@45345.4]
  wire [4:0] _T_92495; // @[Modules.scala 40:46:@45346.4]
  wire [5:0] _T_92715; // @[Modules.scala 40:46:@45584.4]
  wire [4:0] _T_92716; // @[Modules.scala 40:46:@45585.4]
  wire [4:0] _T_92717; // @[Modules.scala 40:46:@45586.4]
  wire [5:0] _T_92771; // @[Modules.scala 43:47:@45640.4]
  wire [4:0] _T_92772; // @[Modules.scala 43:47:@45641.4]
  wire [4:0] _T_92773; // @[Modules.scala 43:47:@45642.4]
  wire [5:0] _T_92778; // @[Modules.scala 43:47:@45647.4]
  wire [4:0] _T_92779; // @[Modules.scala 43:47:@45648.4]
  wire [4:0] _T_92780; // @[Modules.scala 43:47:@45649.4]
  wire [5:0] _T_92784; // @[Modules.scala 40:46:@45655.4]
  wire [4:0] _T_92785; // @[Modules.scala 40:46:@45656.4]
  wire [4:0] _T_92786; // @[Modules.scala 40:46:@45657.4]
  wire [5:0] _T_93012; // @[Modules.scala 43:47:@45896.4]
  wire [4:0] _T_93013; // @[Modules.scala 43:47:@45897.4]
  wire [4:0] _T_93014; // @[Modules.scala 43:47:@45898.4]
  wire [5:0] _T_93144; // @[Modules.scala 40:46:@46051.4]
  wire [4:0] _T_93145; // @[Modules.scala 40:46:@46052.4]
  wire [4:0] _T_93146; // @[Modules.scala 40:46:@46053.4]
  wire [5:0] _T_93166; // @[Modules.scala 40:46:@46078.4]
  wire [4:0] _T_93167; // @[Modules.scala 40:46:@46079.4]
  wire [4:0] _T_93168; // @[Modules.scala 40:46:@46080.4]
  wire [5:0] _T_93173; // @[Modules.scala 43:47:@46085.4]
  wire [4:0] _T_93174; // @[Modules.scala 43:47:@46086.4]
  wire [4:0] _T_93175; // @[Modules.scala 43:47:@46087.4]
  wire [5:0] _T_93314; // @[Modules.scala 37:46:@46252.4]
  wire [4:0] _T_93315; // @[Modules.scala 37:46:@46253.4]
  wire [4:0] _T_93316; // @[Modules.scala 37:46:@46254.4]
  wire [5:0] _T_93346; // @[Modules.scala 43:47:@46290.4]
  wire [4:0] _T_93347; // @[Modules.scala 43:47:@46291.4]
  wire [4:0] _T_93348; // @[Modules.scala 43:47:@46292.4]
  wire [5:0] _T_93374; // @[Modules.scala 43:47:@46325.4]
  wire [4:0] _T_93375; // @[Modules.scala 43:47:@46326.4]
  wire [4:0] _T_93376; // @[Modules.scala 43:47:@46327.4]
  wire [5:0] _T_93425; // @[Modules.scala 43:47:@46386.4]
  wire [4:0] _T_93426; // @[Modules.scala 43:47:@46387.4]
  wire [4:0] _T_93427; // @[Modules.scala 43:47:@46388.4]
  wire [5:0] _T_93858; // @[Modules.scala 40:46:@46849.4]
  wire [4:0] _T_93859; // @[Modules.scala 40:46:@46850.4]
  wire [4:0] _T_93860; // @[Modules.scala 40:46:@46851.4]
  wire [11:0] _T_93878; // @[Modules.scala 50:57:@46871.4]
  wire [10:0] _T_93879; // @[Modules.scala 50:57:@46872.4]
  wire [10:0] buffer_12_392; // @[Modules.scala 50:57:@46873.4]
  wire [11:0] _T_93881; // @[Modules.scala 50:57:@46875.4]
  wire [10:0] _T_93882; // @[Modules.scala 50:57:@46876.4]
  wire [10:0] buffer_12_393; // @[Modules.scala 50:57:@46877.4]
  wire [10:0] buffer_12_7; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_93887; // @[Modules.scala 50:57:@46883.4]
  wire [10:0] _T_93888; // @[Modules.scala 50:57:@46884.4]
  wire [10:0] buffer_12_395; // @[Modules.scala 50:57:@46885.4]
  wire [11:0] _T_93890; // @[Modules.scala 50:57:@46887.4]
  wire [10:0] _T_93891; // @[Modules.scala 50:57:@46888.4]
  wire [10:0] buffer_12_396; // @[Modules.scala 50:57:@46889.4]
  wire [11:0] _T_93893; // @[Modules.scala 50:57:@46891.4]
  wire [10:0] _T_93894; // @[Modules.scala 50:57:@46892.4]
  wire [10:0] buffer_12_397; // @[Modules.scala 50:57:@46893.4]
  wire [11:0] _T_93896; // @[Modules.scala 50:57:@46895.4]
  wire [10:0] _T_93897; // @[Modules.scala 50:57:@46896.4]
  wire [10:0] buffer_12_398; // @[Modules.scala 50:57:@46897.4]
  wire [11:0] _T_93899; // @[Modules.scala 50:57:@46899.4]
  wire [10:0] _T_93900; // @[Modules.scala 50:57:@46900.4]
  wire [10:0] buffer_12_399; // @[Modules.scala 50:57:@46901.4]
  wire [11:0] _T_93959; // @[Modules.scala 50:57:@46979.4]
  wire [10:0] _T_93960; // @[Modules.scala 50:57:@46980.4]
  wire [10:0] buffer_12_419; // @[Modules.scala 50:57:@46981.4]
  wire [11:0] _T_93965; // @[Modules.scala 50:57:@46987.4]
  wire [10:0] _T_93966; // @[Modules.scala 50:57:@46988.4]
  wire [10:0] buffer_12_421; // @[Modules.scala 50:57:@46989.4]
  wire [11:0] _T_93971; // @[Modules.scala 50:57:@46995.4]
  wire [10:0] _T_93972; // @[Modules.scala 50:57:@46996.4]
  wire [10:0] buffer_12_423; // @[Modules.scala 50:57:@46997.4]
  wire [11:0] _T_93977; // @[Modules.scala 50:57:@47003.4]
  wire [10:0] _T_93978; // @[Modules.scala 50:57:@47004.4]
  wire [10:0] buffer_12_425; // @[Modules.scala 50:57:@47005.4]
  wire [11:0] _T_93980; // @[Modules.scala 50:57:@47007.4]
  wire [10:0] _T_93981; // @[Modules.scala 50:57:@47008.4]
  wire [10:0] buffer_12_426; // @[Modules.scala 50:57:@47009.4]
  wire [11:0] _T_93986; // @[Modules.scala 50:57:@47015.4]
  wire [10:0] _T_93987; // @[Modules.scala 50:57:@47016.4]
  wire [10:0] buffer_12_428; // @[Modules.scala 50:57:@47017.4]
  wire [11:0] _T_93989; // @[Modules.scala 50:57:@47019.4]
  wire [10:0] _T_93990; // @[Modules.scala 50:57:@47020.4]
  wire [10:0] buffer_12_429; // @[Modules.scala 50:57:@47021.4]
  wire [11:0] _T_93995; // @[Modules.scala 50:57:@47027.4]
  wire [10:0] _T_93996; // @[Modules.scala 50:57:@47028.4]
  wire [10:0] buffer_12_431; // @[Modules.scala 50:57:@47029.4]
  wire [11:0] _T_94001; // @[Modules.scala 50:57:@47035.4]
  wire [10:0] _T_94002; // @[Modules.scala 50:57:@47036.4]
  wire [10:0] buffer_12_433; // @[Modules.scala 50:57:@47037.4]
  wire [11:0] _T_94016; // @[Modules.scala 50:57:@47055.4]
  wire [10:0] _T_94017; // @[Modules.scala 50:57:@47056.4]
  wire [10:0] buffer_12_438; // @[Modules.scala 50:57:@47057.4]
  wire [11:0] _T_94028; // @[Modules.scala 50:57:@47071.4]
  wire [10:0] _T_94029; // @[Modules.scala 50:57:@47072.4]
  wire [10:0] buffer_12_442; // @[Modules.scala 50:57:@47073.4]
  wire [11:0] _T_94031; // @[Modules.scala 50:57:@47075.4]
  wire [10:0] _T_94032; // @[Modules.scala 50:57:@47076.4]
  wire [10:0] buffer_12_443; // @[Modules.scala 50:57:@47077.4]
  wire [11:0] _T_94037; // @[Modules.scala 50:57:@47083.4]
  wire [10:0] _T_94038; // @[Modules.scala 50:57:@47084.4]
  wire [10:0] buffer_12_445; // @[Modules.scala 50:57:@47085.4]
  wire [10:0] buffer_12_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94046; // @[Modules.scala 50:57:@47095.4]
  wire [10:0] _T_94047; // @[Modules.scala 50:57:@47096.4]
  wire [10:0] buffer_12_448; // @[Modules.scala 50:57:@47097.4]
  wire [11:0] _T_94052; // @[Modules.scala 50:57:@47103.4]
  wire [10:0] _T_94053; // @[Modules.scala 50:57:@47104.4]
  wire [10:0] buffer_12_450; // @[Modules.scala 50:57:@47105.4]
  wire [11:0] _T_94055; // @[Modules.scala 50:57:@47107.4]
  wire [10:0] _T_94056; // @[Modules.scala 50:57:@47108.4]
  wire [10:0] buffer_12_451; // @[Modules.scala 50:57:@47109.4]
  wire [11:0] _T_94067; // @[Modules.scala 50:57:@47123.4]
  wire [10:0] _T_94068; // @[Modules.scala 50:57:@47124.4]
  wire [10:0] buffer_12_455; // @[Modules.scala 50:57:@47125.4]
  wire [11:0] _T_94070; // @[Modules.scala 50:57:@47127.4]
  wire [10:0] _T_94071; // @[Modules.scala 50:57:@47128.4]
  wire [10:0] buffer_12_456; // @[Modules.scala 50:57:@47129.4]
  wire [11:0] _T_94073; // @[Modules.scala 50:57:@47131.4]
  wire [10:0] _T_94074; // @[Modules.scala 50:57:@47132.4]
  wire [10:0] buffer_12_457; // @[Modules.scala 50:57:@47133.4]
  wire [11:0] _T_94076; // @[Modules.scala 50:57:@47135.4]
  wire [10:0] _T_94077; // @[Modules.scala 50:57:@47136.4]
  wire [10:0] buffer_12_458; // @[Modules.scala 50:57:@47137.4]
  wire [11:0] _T_94079; // @[Modules.scala 50:57:@47139.4]
  wire [10:0] _T_94080; // @[Modules.scala 50:57:@47140.4]
  wire [10:0] buffer_12_459; // @[Modules.scala 50:57:@47141.4]
  wire [11:0] _T_94088; // @[Modules.scala 50:57:@47151.4]
  wire [10:0] _T_94089; // @[Modules.scala 50:57:@47152.4]
  wire [10:0] buffer_12_462; // @[Modules.scala 50:57:@47153.4]
  wire [11:0] _T_94100; // @[Modules.scala 50:57:@47167.4]
  wire [10:0] _T_94101; // @[Modules.scala 50:57:@47168.4]
  wire [10:0] buffer_12_466; // @[Modules.scala 50:57:@47169.4]
  wire [11:0] _T_94103; // @[Modules.scala 50:57:@47171.4]
  wire [10:0] _T_94104; // @[Modules.scala 50:57:@47172.4]
  wire [10:0] buffer_12_467; // @[Modules.scala 50:57:@47173.4]
  wire [10:0] buffer_12_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94109; // @[Modules.scala 50:57:@47179.4]
  wire [10:0] _T_94110; // @[Modules.scala 50:57:@47180.4]
  wire [10:0] buffer_12_469; // @[Modules.scala 50:57:@47181.4]
  wire [10:0] buffer_12_163; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94121; // @[Modules.scala 50:57:@47195.4]
  wire [10:0] _T_94122; // @[Modules.scala 50:57:@47196.4]
  wire [10:0] buffer_12_473; // @[Modules.scala 50:57:@47197.4]
  wire [10:0] buffer_12_164; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94124; // @[Modules.scala 50:57:@47199.4]
  wire [10:0] _T_94125; // @[Modules.scala 50:57:@47200.4]
  wire [10:0] buffer_12_474; // @[Modules.scala 50:57:@47201.4]
  wire [10:0] buffer_12_166; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94127; // @[Modules.scala 50:57:@47203.4]
  wire [10:0] _T_94128; // @[Modules.scala 50:57:@47204.4]
  wire [10:0] buffer_12_475; // @[Modules.scala 50:57:@47205.4]
  wire [11:0] _T_94130; // @[Modules.scala 50:57:@47207.4]
  wire [10:0] _T_94131; // @[Modules.scala 50:57:@47208.4]
  wire [10:0] buffer_12_476; // @[Modules.scala 50:57:@47209.4]
  wire [11:0] _T_94172; // @[Modules.scala 50:57:@47263.4]
  wire [10:0] _T_94173; // @[Modules.scala 50:57:@47264.4]
  wire [10:0] buffer_12_490; // @[Modules.scala 50:57:@47265.4]
  wire [11:0] _T_94175; // @[Modules.scala 50:57:@47267.4]
  wire [10:0] _T_94176; // @[Modules.scala 50:57:@47268.4]
  wire [10:0] buffer_12_491; // @[Modules.scala 50:57:@47269.4]
  wire [10:0] buffer_12_206; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94187; // @[Modules.scala 50:57:@47283.4]
  wire [10:0] _T_94188; // @[Modules.scala 50:57:@47284.4]
  wire [10:0] buffer_12_495; // @[Modules.scala 50:57:@47285.4]
  wire [11:0] _T_94193; // @[Modules.scala 50:57:@47291.4]
  wire [10:0] _T_94194; // @[Modules.scala 50:57:@47292.4]
  wire [10:0] buffer_12_497; // @[Modules.scala 50:57:@47293.4]
  wire [11:0] _T_94208; // @[Modules.scala 50:57:@47311.4]
  wire [10:0] _T_94209; // @[Modules.scala 50:57:@47312.4]
  wire [10:0] buffer_12_502; // @[Modules.scala 50:57:@47313.4]
  wire [11:0] _T_94223; // @[Modules.scala 50:57:@47331.4]
  wire [10:0] _T_94224; // @[Modules.scala 50:57:@47332.4]
  wire [10:0] buffer_12_507; // @[Modules.scala 50:57:@47333.4]
  wire [11:0] _T_94229; // @[Modules.scala 50:57:@47339.4]
  wire [10:0] _T_94230; // @[Modules.scala 50:57:@47340.4]
  wire [10:0] buffer_12_509; // @[Modules.scala 50:57:@47341.4]
  wire [10:0] buffer_12_238; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94235; // @[Modules.scala 50:57:@47347.4]
  wire [10:0] _T_94236; // @[Modules.scala 50:57:@47348.4]
  wire [10:0] buffer_12_511; // @[Modules.scala 50:57:@47349.4]
  wire [10:0] buffer_12_244; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_12_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94244; // @[Modules.scala 50:57:@47359.4]
  wire [10:0] _T_94245; // @[Modules.scala 50:57:@47360.4]
  wire [10:0] buffer_12_514; // @[Modules.scala 50:57:@47361.4]
  wire [11:0] _T_94256; // @[Modules.scala 50:57:@47375.4]
  wire [10:0] _T_94257; // @[Modules.scala 50:57:@47376.4]
  wire [10:0] buffer_12_518; // @[Modules.scala 50:57:@47377.4]
  wire [11:0] _T_94259; // @[Modules.scala 50:57:@47379.4]
  wire [10:0] _T_94260; // @[Modules.scala 50:57:@47380.4]
  wire [10:0] buffer_12_519; // @[Modules.scala 50:57:@47381.4]
  wire [11:0] _T_94265; // @[Modules.scala 50:57:@47387.4]
  wire [10:0] _T_94266; // @[Modules.scala 50:57:@47388.4]
  wire [10:0] buffer_12_521; // @[Modules.scala 50:57:@47389.4]
  wire [11:0] _T_94271; // @[Modules.scala 50:57:@47395.4]
  wire [10:0] _T_94272; // @[Modules.scala 50:57:@47396.4]
  wire [10:0] buffer_12_523; // @[Modules.scala 50:57:@47397.4]
  wire [11:0] _T_94277; // @[Modules.scala 50:57:@47403.4]
  wire [10:0] _T_94278; // @[Modules.scala 50:57:@47404.4]
  wire [10:0] buffer_12_525; // @[Modules.scala 50:57:@47405.4]
  wire [11:0] _T_94289; // @[Modules.scala 50:57:@47419.4]
  wire [10:0] _T_94290; // @[Modules.scala 50:57:@47420.4]
  wire [10:0] buffer_12_529; // @[Modules.scala 50:57:@47421.4]
  wire [10:0] buffer_12_280; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94298; // @[Modules.scala 50:57:@47431.4]
  wire [10:0] _T_94299; // @[Modules.scala 50:57:@47432.4]
  wire [10:0] buffer_12_532; // @[Modules.scala 50:57:@47433.4]
  wire [10:0] buffer_12_288; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94310; // @[Modules.scala 50:57:@47447.4]
  wire [10:0] _T_94311; // @[Modules.scala 50:57:@47448.4]
  wire [10:0] buffer_12_536; // @[Modules.scala 50:57:@47449.4]
  wire [11:0] _T_94319; // @[Modules.scala 50:57:@47459.4]
  wire [10:0] _T_94320; // @[Modules.scala 50:57:@47460.4]
  wire [10:0] buffer_12_539; // @[Modules.scala 50:57:@47461.4]
  wire [10:0] buffer_12_296; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94322; // @[Modules.scala 50:57:@47463.4]
  wire [10:0] _T_94323; // @[Modules.scala 50:57:@47464.4]
  wire [10:0] buffer_12_540; // @[Modules.scala 50:57:@47465.4]
  wire [11:0] _T_94325; // @[Modules.scala 50:57:@47467.4]
  wire [10:0] _T_94326; // @[Modules.scala 50:57:@47468.4]
  wire [10:0] buffer_12_541; // @[Modules.scala 50:57:@47469.4]
  wire [10:0] buffer_12_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94340; // @[Modules.scala 50:57:@47487.4]
  wire [10:0] _T_94341; // @[Modules.scala 50:57:@47488.4]
  wire [10:0] buffer_12_546; // @[Modules.scala 50:57:@47489.4]
  wire [11:0] _T_94361; // @[Modules.scala 50:57:@47515.4]
  wire [10:0] _T_94362; // @[Modules.scala 50:57:@47516.4]
  wire [10:0] buffer_12_553; // @[Modules.scala 50:57:@47517.4]
  wire [11:0] _T_94379; // @[Modules.scala 50:57:@47539.4]
  wire [10:0] _T_94380; // @[Modules.scala 50:57:@47540.4]
  wire [10:0] buffer_12_559; // @[Modules.scala 50:57:@47541.4]
  wire [11:0] _T_94388; // @[Modules.scala 50:57:@47551.4]
  wire [10:0] _T_94389; // @[Modules.scala 50:57:@47552.4]
  wire [10:0] buffer_12_562; // @[Modules.scala 50:57:@47553.4]
  wire [11:0] _T_94391; // @[Modules.scala 50:57:@47555.4]
  wire [10:0] _T_94392; // @[Modules.scala 50:57:@47556.4]
  wire [10:0] buffer_12_563; // @[Modules.scala 50:57:@47557.4]
  wire [11:0] _T_94400; // @[Modules.scala 50:57:@47567.4]
  wire [10:0] _T_94401; // @[Modules.scala 50:57:@47568.4]
  wire [10:0] buffer_12_566; // @[Modules.scala 50:57:@47569.4]
  wire [11:0] _T_94403; // @[Modules.scala 50:57:@47571.4]
  wire [10:0] _T_94404; // @[Modules.scala 50:57:@47572.4]
  wire [10:0] buffer_12_567; // @[Modules.scala 50:57:@47573.4]
  wire [11:0] _T_94424; // @[Modules.scala 50:57:@47599.4]
  wire [10:0] _T_94425; // @[Modules.scala 50:57:@47600.4]
  wire [10:0] buffer_12_574; // @[Modules.scala 50:57:@47601.4]
  wire [11:0] _T_94442; // @[Modules.scala 50:57:@47623.4]
  wire [10:0] _T_94443; // @[Modules.scala 50:57:@47624.4]
  wire [10:0] buffer_12_580; // @[Modules.scala 50:57:@47625.4]
  wire [11:0] _T_94445; // @[Modules.scala 50:57:@47627.4]
  wire [10:0] _T_94446; // @[Modules.scala 50:57:@47628.4]
  wire [10:0] buffer_12_581; // @[Modules.scala 50:57:@47629.4]
  wire [11:0] _T_94451; // @[Modules.scala 50:57:@47635.4]
  wire [10:0] _T_94452; // @[Modules.scala 50:57:@47636.4]
  wire [10:0] buffer_12_583; // @[Modules.scala 50:57:@47637.4]
  wire [10:0] buffer_12_388; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_94460; // @[Modules.scala 50:57:@47647.4]
  wire [10:0] _T_94461; // @[Modules.scala 50:57:@47648.4]
  wire [10:0] buffer_12_586; // @[Modules.scala 50:57:@47649.4]
  wire [11:0] _T_94466; // @[Modules.scala 53:83:@47655.4]
  wire [10:0] _T_94467; // @[Modules.scala 53:83:@47656.4]
  wire [10:0] buffer_12_588; // @[Modules.scala 53:83:@47657.4]
  wire [11:0] _T_94469; // @[Modules.scala 53:83:@47659.4]
  wire [10:0] _T_94470; // @[Modules.scala 53:83:@47660.4]
  wire [10:0] buffer_12_589; // @[Modules.scala 53:83:@47661.4]
  wire [11:0] _T_94472; // @[Modules.scala 53:83:@47663.4]
  wire [10:0] _T_94473; // @[Modules.scala 53:83:@47664.4]
  wire [10:0] buffer_12_590; // @[Modules.scala 53:83:@47665.4]
  wire [11:0] _T_94475; // @[Modules.scala 53:83:@47667.4]
  wire [10:0] _T_94476; // @[Modules.scala 53:83:@47668.4]
  wire [10:0] buffer_12_591; // @[Modules.scala 53:83:@47669.4]
  wire [11:0] _T_94487; // @[Modules.scala 53:83:@47683.4]
  wire [10:0] _T_94488; // @[Modules.scala 53:83:@47684.4]
  wire [10:0] buffer_12_595; // @[Modules.scala 53:83:@47685.4]
  wire [11:0] _T_94496; // @[Modules.scala 53:83:@47695.4]
  wire [10:0] _T_94497; // @[Modules.scala 53:83:@47696.4]
  wire [10:0] buffer_12_598; // @[Modules.scala 53:83:@47697.4]
  wire [11:0] _T_94505; // @[Modules.scala 53:83:@47707.4]
  wire [10:0] _T_94506; // @[Modules.scala 53:83:@47708.4]
  wire [10:0] buffer_12_601; // @[Modules.scala 53:83:@47709.4]
  wire [11:0] _T_94508; // @[Modules.scala 53:83:@47711.4]
  wire [10:0] _T_94509; // @[Modules.scala 53:83:@47712.4]
  wire [10:0] buffer_12_602; // @[Modules.scala 53:83:@47713.4]
  wire [11:0] _T_94511; // @[Modules.scala 53:83:@47715.4]
  wire [10:0] _T_94512; // @[Modules.scala 53:83:@47716.4]
  wire [10:0] buffer_12_603; // @[Modules.scala 53:83:@47717.4]
  wire [11:0] _T_94514; // @[Modules.scala 53:83:@47719.4]
  wire [10:0] _T_94515; // @[Modules.scala 53:83:@47720.4]
  wire [10:0] buffer_12_604; // @[Modules.scala 53:83:@47721.4]
  wire [11:0] _T_94517; // @[Modules.scala 53:83:@47723.4]
  wire [10:0] _T_94518; // @[Modules.scala 53:83:@47724.4]
  wire [10:0] buffer_12_605; // @[Modules.scala 53:83:@47725.4]
  wire [11:0] _T_94520; // @[Modules.scala 53:83:@47727.4]
  wire [10:0] _T_94521; // @[Modules.scala 53:83:@47728.4]
  wire [10:0] buffer_12_606; // @[Modules.scala 53:83:@47729.4]
  wire [11:0] _T_94523; // @[Modules.scala 53:83:@47731.4]
  wire [10:0] _T_94524; // @[Modules.scala 53:83:@47732.4]
  wire [10:0] buffer_12_607; // @[Modules.scala 53:83:@47733.4]
  wire [11:0] _T_94526; // @[Modules.scala 53:83:@47735.4]
  wire [10:0] _T_94527; // @[Modules.scala 53:83:@47736.4]
  wire [10:0] buffer_12_608; // @[Modules.scala 53:83:@47737.4]
  wire [11:0] _T_94532; // @[Modules.scala 53:83:@47743.4]
  wire [10:0] _T_94533; // @[Modules.scala 53:83:@47744.4]
  wire [10:0] buffer_12_610; // @[Modules.scala 53:83:@47745.4]
  wire [11:0] _T_94535; // @[Modules.scala 53:83:@47747.4]
  wire [10:0] _T_94536; // @[Modules.scala 53:83:@47748.4]
  wire [10:0] buffer_12_611; // @[Modules.scala 53:83:@47749.4]
  wire [11:0] _T_94541; // @[Modules.scala 53:83:@47755.4]
  wire [10:0] _T_94542; // @[Modules.scala 53:83:@47756.4]
  wire [10:0] buffer_12_613; // @[Modules.scala 53:83:@47757.4]
  wire [11:0] _T_94544; // @[Modules.scala 53:83:@47759.4]
  wire [10:0] _T_94545; // @[Modules.scala 53:83:@47760.4]
  wire [10:0] buffer_12_614; // @[Modules.scala 53:83:@47761.4]
  wire [11:0] _T_94550; // @[Modules.scala 53:83:@47767.4]
  wire [10:0] _T_94551; // @[Modules.scala 53:83:@47768.4]
  wire [10:0] buffer_12_616; // @[Modules.scala 53:83:@47769.4]
  wire [11:0] _T_94553; // @[Modules.scala 53:83:@47771.4]
  wire [10:0] _T_94554; // @[Modules.scala 53:83:@47772.4]
  wire [10:0] buffer_12_617; // @[Modules.scala 53:83:@47773.4]
  wire [11:0] _T_94556; // @[Modules.scala 53:83:@47775.4]
  wire [10:0] _T_94557; // @[Modules.scala 53:83:@47776.4]
  wire [10:0] buffer_12_618; // @[Modules.scala 53:83:@47777.4]
  wire [11:0] _T_94559; // @[Modules.scala 53:83:@47779.4]
  wire [10:0] _T_94560; // @[Modules.scala 53:83:@47780.4]
  wire [10:0] buffer_12_619; // @[Modules.scala 53:83:@47781.4]
  wire [11:0] _T_94562; // @[Modules.scala 53:83:@47783.4]
  wire [10:0] _T_94563; // @[Modules.scala 53:83:@47784.4]
  wire [10:0] buffer_12_620; // @[Modules.scala 53:83:@47785.4]
  wire [11:0] _T_94565; // @[Modules.scala 53:83:@47787.4]
  wire [10:0] _T_94566; // @[Modules.scala 53:83:@47788.4]
  wire [10:0] buffer_12_621; // @[Modules.scala 53:83:@47789.4]
  wire [11:0] _T_94571; // @[Modules.scala 53:83:@47795.4]
  wire [10:0] _T_94572; // @[Modules.scala 53:83:@47796.4]
  wire [10:0] buffer_12_623; // @[Modules.scala 53:83:@47797.4]
  wire [11:0] _T_94574; // @[Modules.scala 53:83:@47799.4]
  wire [10:0] _T_94575; // @[Modules.scala 53:83:@47800.4]
  wire [10:0] buffer_12_624; // @[Modules.scala 53:83:@47801.4]
  wire [11:0] _T_94577; // @[Modules.scala 53:83:@47803.4]
  wire [10:0] _T_94578; // @[Modules.scala 53:83:@47804.4]
  wire [10:0] buffer_12_625; // @[Modules.scala 53:83:@47805.4]
  wire [11:0] _T_94580; // @[Modules.scala 53:83:@47807.4]
  wire [10:0] _T_94581; // @[Modules.scala 53:83:@47808.4]
  wire [10:0] buffer_12_626; // @[Modules.scala 53:83:@47809.4]
  wire [11:0] _T_94586; // @[Modules.scala 53:83:@47815.4]
  wire [10:0] _T_94587; // @[Modules.scala 53:83:@47816.4]
  wire [10:0] buffer_12_628; // @[Modules.scala 53:83:@47817.4]
  wire [11:0] _T_94589; // @[Modules.scala 53:83:@47819.4]
  wire [10:0] _T_94590; // @[Modules.scala 53:83:@47820.4]
  wire [10:0] buffer_12_629; // @[Modules.scala 53:83:@47821.4]
  wire [11:0] _T_94592; // @[Modules.scala 53:83:@47823.4]
  wire [10:0] _T_94593; // @[Modules.scala 53:83:@47824.4]
  wire [10:0] buffer_12_630; // @[Modules.scala 53:83:@47825.4]
  wire [11:0] _T_94598; // @[Modules.scala 53:83:@47831.4]
  wire [10:0] _T_94599; // @[Modules.scala 53:83:@47832.4]
  wire [10:0] buffer_12_632; // @[Modules.scala 53:83:@47833.4]
  wire [11:0] _T_94601; // @[Modules.scala 53:83:@47835.4]
  wire [10:0] _T_94602; // @[Modules.scala 53:83:@47836.4]
  wire [10:0] buffer_12_633; // @[Modules.scala 53:83:@47837.4]
  wire [11:0] _T_94607; // @[Modules.scala 53:83:@47843.4]
  wire [10:0] _T_94608; // @[Modules.scala 53:83:@47844.4]
  wire [10:0] buffer_12_635; // @[Modules.scala 53:83:@47845.4]
  wire [11:0] _T_94610; // @[Modules.scala 53:83:@47847.4]
  wire [10:0] _T_94611; // @[Modules.scala 53:83:@47848.4]
  wire [10:0] buffer_12_636; // @[Modules.scala 53:83:@47849.4]
  wire [11:0] _T_94613; // @[Modules.scala 53:83:@47851.4]
  wire [10:0] _T_94614; // @[Modules.scala 53:83:@47852.4]
  wire [10:0] buffer_12_637; // @[Modules.scala 53:83:@47853.4]
  wire [11:0] _T_94616; // @[Modules.scala 53:83:@47855.4]
  wire [10:0] _T_94617; // @[Modules.scala 53:83:@47856.4]
  wire [10:0] buffer_12_638; // @[Modules.scala 53:83:@47857.4]
  wire [11:0] _T_94619; // @[Modules.scala 53:83:@47859.4]
  wire [10:0] _T_94620; // @[Modules.scala 53:83:@47860.4]
  wire [10:0] buffer_12_639; // @[Modules.scala 53:83:@47861.4]
  wire [11:0] _T_94622; // @[Modules.scala 53:83:@47863.4]
  wire [10:0] _T_94623; // @[Modules.scala 53:83:@47864.4]
  wire [10:0] buffer_12_640; // @[Modules.scala 53:83:@47865.4]
  wire [11:0] _T_94631; // @[Modules.scala 53:83:@47875.4]
  wire [10:0] _T_94632; // @[Modules.scala 53:83:@47876.4]
  wire [10:0] buffer_12_643; // @[Modules.scala 53:83:@47877.4]
  wire [11:0] _T_94637; // @[Modules.scala 53:83:@47883.4]
  wire [10:0] _T_94638; // @[Modules.scala 53:83:@47884.4]
  wire [10:0] buffer_12_645; // @[Modules.scala 53:83:@47885.4]
  wire [11:0] _T_94640; // @[Modules.scala 53:83:@47887.4]
  wire [10:0] _T_94641; // @[Modules.scala 53:83:@47888.4]
  wire [10:0] buffer_12_646; // @[Modules.scala 53:83:@47889.4]
  wire [11:0] _T_94643; // @[Modules.scala 53:83:@47891.4]
  wire [10:0] _T_94644; // @[Modules.scala 53:83:@47892.4]
  wire [10:0] buffer_12_647; // @[Modules.scala 53:83:@47893.4]
  wire [11:0] _T_94646; // @[Modules.scala 53:83:@47895.4]
  wire [10:0] _T_94647; // @[Modules.scala 53:83:@47896.4]
  wire [10:0] buffer_12_648; // @[Modules.scala 53:83:@47897.4]
  wire [11:0] _T_94649; // @[Modules.scala 53:83:@47899.4]
  wire [10:0] _T_94650; // @[Modules.scala 53:83:@47900.4]
  wire [10:0] buffer_12_649; // @[Modules.scala 53:83:@47901.4]
  wire [11:0] _T_94655; // @[Modules.scala 53:83:@47907.4]
  wire [10:0] _T_94656; // @[Modules.scala 53:83:@47908.4]
  wire [10:0] buffer_12_651; // @[Modules.scala 53:83:@47909.4]
  wire [11:0] _T_94658; // @[Modules.scala 53:83:@47911.4]
  wire [10:0] _T_94659; // @[Modules.scala 53:83:@47912.4]
  wire [10:0] buffer_12_652; // @[Modules.scala 53:83:@47913.4]
  wire [11:0] _T_94661; // @[Modules.scala 53:83:@47915.4]
  wire [10:0] _T_94662; // @[Modules.scala 53:83:@47916.4]
  wire [10:0] buffer_12_653; // @[Modules.scala 53:83:@47917.4]
  wire [11:0] _T_94664; // @[Modules.scala 53:83:@47919.4]
  wire [10:0] _T_94665; // @[Modules.scala 53:83:@47920.4]
  wire [10:0] buffer_12_654; // @[Modules.scala 53:83:@47921.4]
  wire [11:0] _T_94670; // @[Modules.scala 53:83:@47927.4]
  wire [10:0] _T_94671; // @[Modules.scala 53:83:@47928.4]
  wire [10:0] buffer_12_656; // @[Modules.scala 53:83:@47929.4]
  wire [11:0] _T_94676; // @[Modules.scala 53:83:@47935.4]
  wire [10:0] _T_94677; // @[Modules.scala 53:83:@47936.4]
  wire [10:0] buffer_12_658; // @[Modules.scala 53:83:@47937.4]
  wire [11:0] _T_94682; // @[Modules.scala 53:83:@47943.4]
  wire [10:0] _T_94683; // @[Modules.scala 53:83:@47944.4]
  wire [10:0] buffer_12_660; // @[Modules.scala 53:83:@47945.4]
  wire [11:0] _T_94685; // @[Modules.scala 53:83:@47947.4]
  wire [10:0] _T_94686; // @[Modules.scala 53:83:@47948.4]
  wire [10:0] buffer_12_661; // @[Modules.scala 53:83:@47949.4]
  wire [11:0] _T_94688; // @[Modules.scala 53:83:@47951.4]
  wire [10:0] _T_94689; // @[Modules.scala 53:83:@47952.4]
  wire [10:0] buffer_12_662; // @[Modules.scala 53:83:@47953.4]
  wire [11:0] _T_94694; // @[Modules.scala 53:83:@47959.4]
  wire [10:0] _T_94695; // @[Modules.scala 53:83:@47960.4]
  wire [10:0] buffer_12_664; // @[Modules.scala 53:83:@47961.4]
  wire [11:0] _T_94697; // @[Modules.scala 53:83:@47963.4]
  wire [10:0] _T_94698; // @[Modules.scala 53:83:@47964.4]
  wire [10:0] buffer_12_665; // @[Modules.scala 53:83:@47965.4]
  wire [11:0] _T_94700; // @[Modules.scala 53:83:@47967.4]
  wire [10:0] _T_94701; // @[Modules.scala 53:83:@47968.4]
  wire [10:0] buffer_12_666; // @[Modules.scala 53:83:@47969.4]
  wire [11:0] _T_94703; // @[Modules.scala 53:83:@47971.4]
  wire [10:0] _T_94704; // @[Modules.scala 53:83:@47972.4]
  wire [10:0] buffer_12_667; // @[Modules.scala 53:83:@47973.4]
  wire [11:0] _T_94706; // @[Modules.scala 53:83:@47975.4]
  wire [10:0] _T_94707; // @[Modules.scala 53:83:@47976.4]
  wire [10:0] buffer_12_668; // @[Modules.scala 53:83:@47977.4]
  wire [11:0] _T_94709; // @[Modules.scala 53:83:@47979.4]
  wire [10:0] _T_94710; // @[Modules.scala 53:83:@47980.4]
  wire [10:0] buffer_12_669; // @[Modules.scala 53:83:@47981.4]
  wire [11:0] _T_94715; // @[Modules.scala 53:83:@47987.4]
  wire [10:0] _T_94716; // @[Modules.scala 53:83:@47988.4]
  wire [10:0] buffer_12_671; // @[Modules.scala 53:83:@47989.4]
  wire [11:0] _T_94721; // @[Modules.scala 53:83:@47995.4]
  wire [10:0] _T_94722; // @[Modules.scala 53:83:@47996.4]
  wire [10:0] buffer_12_673; // @[Modules.scala 53:83:@47997.4]
  wire [11:0] _T_94727; // @[Modules.scala 53:83:@48003.4]
  wire [10:0] _T_94728; // @[Modules.scala 53:83:@48004.4]
  wire [10:0] buffer_12_675; // @[Modules.scala 53:83:@48005.4]
  wire [11:0] _T_94739; // @[Modules.scala 53:83:@48019.4]
  wire [10:0] _T_94740; // @[Modules.scala 53:83:@48020.4]
  wire [10:0] buffer_12_679; // @[Modules.scala 53:83:@48021.4]
  wire [11:0] _T_94748; // @[Modules.scala 53:83:@48031.4]
  wire [10:0] _T_94749; // @[Modules.scala 53:83:@48032.4]
  wire [10:0] buffer_12_682; // @[Modules.scala 53:83:@48033.4]
  wire [11:0] _T_94751; // @[Modules.scala 53:83:@48035.4]
  wire [10:0] _T_94752; // @[Modules.scala 53:83:@48036.4]
  wire [10:0] buffer_12_683; // @[Modules.scala 53:83:@48037.4]
  wire [11:0] _T_94757; // @[Modules.scala 53:83:@48043.4]
  wire [10:0] _T_94758; // @[Modules.scala 53:83:@48044.4]
  wire [10:0] buffer_12_685; // @[Modules.scala 53:83:@48045.4]
  wire [11:0] _T_94760; // @[Modules.scala 56:109:@48047.4]
  wire [10:0] _T_94761; // @[Modules.scala 56:109:@48048.4]
  wire [10:0] buffer_12_686; // @[Modules.scala 56:109:@48049.4]
  wire [11:0] _T_94763; // @[Modules.scala 56:109:@48051.4]
  wire [10:0] _T_94764; // @[Modules.scala 56:109:@48052.4]
  wire [10:0] buffer_12_687; // @[Modules.scala 56:109:@48053.4]
  wire [11:0] _T_94766; // @[Modules.scala 56:109:@48055.4]
  wire [10:0] _T_94767; // @[Modules.scala 56:109:@48056.4]
  wire [10:0] buffer_12_688; // @[Modules.scala 56:109:@48057.4]
  wire [11:0] _T_94769; // @[Modules.scala 56:109:@48059.4]
  wire [10:0] _T_94770; // @[Modules.scala 56:109:@48060.4]
  wire [10:0] buffer_12_689; // @[Modules.scala 56:109:@48061.4]
  wire [11:0] _T_94775; // @[Modules.scala 56:109:@48067.4]
  wire [10:0] _T_94776; // @[Modules.scala 56:109:@48068.4]
  wire [10:0] buffer_12_691; // @[Modules.scala 56:109:@48069.4]
  wire [11:0] _T_94778; // @[Modules.scala 56:109:@48071.4]
  wire [10:0] _T_94779; // @[Modules.scala 56:109:@48072.4]
  wire [10:0] buffer_12_692; // @[Modules.scala 56:109:@48073.4]
  wire [11:0] _T_94781; // @[Modules.scala 56:109:@48075.4]
  wire [10:0] _T_94782; // @[Modules.scala 56:109:@48076.4]
  wire [10:0] buffer_12_693; // @[Modules.scala 56:109:@48077.4]
  wire [11:0] _T_94784; // @[Modules.scala 56:109:@48079.4]
  wire [10:0] _T_94785; // @[Modules.scala 56:109:@48080.4]
  wire [10:0] buffer_12_694; // @[Modules.scala 56:109:@48081.4]
  wire [11:0] _T_94787; // @[Modules.scala 56:109:@48083.4]
  wire [10:0] _T_94788; // @[Modules.scala 56:109:@48084.4]
  wire [10:0] buffer_12_695; // @[Modules.scala 56:109:@48085.4]
  wire [11:0] _T_94790; // @[Modules.scala 56:109:@48087.4]
  wire [10:0] _T_94791; // @[Modules.scala 56:109:@48088.4]
  wire [10:0] buffer_12_696; // @[Modules.scala 56:109:@48089.4]
  wire [11:0] _T_94793; // @[Modules.scala 56:109:@48091.4]
  wire [10:0] _T_94794; // @[Modules.scala 56:109:@48092.4]
  wire [10:0] buffer_12_697; // @[Modules.scala 56:109:@48093.4]
  wire [11:0] _T_94796; // @[Modules.scala 56:109:@48095.4]
  wire [10:0] _T_94797; // @[Modules.scala 56:109:@48096.4]
  wire [10:0] buffer_12_698; // @[Modules.scala 56:109:@48097.4]
  wire [11:0] _T_94799; // @[Modules.scala 56:109:@48099.4]
  wire [10:0] _T_94800; // @[Modules.scala 56:109:@48100.4]
  wire [10:0] buffer_12_699; // @[Modules.scala 56:109:@48101.4]
  wire [11:0] _T_94802; // @[Modules.scala 56:109:@48103.4]
  wire [10:0] _T_94803; // @[Modules.scala 56:109:@48104.4]
  wire [10:0] buffer_12_700; // @[Modules.scala 56:109:@48105.4]
  wire [11:0] _T_94805; // @[Modules.scala 56:109:@48107.4]
  wire [10:0] _T_94806; // @[Modules.scala 56:109:@48108.4]
  wire [10:0] buffer_12_701; // @[Modules.scala 56:109:@48109.4]
  wire [11:0] _T_94808; // @[Modules.scala 56:109:@48111.4]
  wire [10:0] _T_94809; // @[Modules.scala 56:109:@48112.4]
  wire [10:0] buffer_12_702; // @[Modules.scala 56:109:@48113.4]
  wire [11:0] _T_94811; // @[Modules.scala 56:109:@48115.4]
  wire [10:0] _T_94812; // @[Modules.scala 56:109:@48116.4]
  wire [10:0] buffer_12_703; // @[Modules.scala 56:109:@48117.4]
  wire [11:0] _T_94814; // @[Modules.scala 56:109:@48119.4]
  wire [10:0] _T_94815; // @[Modules.scala 56:109:@48120.4]
  wire [10:0] buffer_12_704; // @[Modules.scala 56:109:@48121.4]
  wire [11:0] _T_94817; // @[Modules.scala 56:109:@48123.4]
  wire [10:0] _T_94818; // @[Modules.scala 56:109:@48124.4]
  wire [10:0] buffer_12_705; // @[Modules.scala 56:109:@48125.4]
  wire [11:0] _T_94820; // @[Modules.scala 56:109:@48127.4]
  wire [10:0] _T_94821; // @[Modules.scala 56:109:@48128.4]
  wire [10:0] buffer_12_706; // @[Modules.scala 56:109:@48129.4]
  wire [11:0] _T_94823; // @[Modules.scala 56:109:@48131.4]
  wire [10:0] _T_94824; // @[Modules.scala 56:109:@48132.4]
  wire [10:0] buffer_12_707; // @[Modules.scala 56:109:@48133.4]
  wire [11:0] _T_94826; // @[Modules.scala 56:109:@48135.4]
  wire [10:0] _T_94827; // @[Modules.scala 56:109:@48136.4]
  wire [10:0] buffer_12_708; // @[Modules.scala 56:109:@48137.4]
  wire [11:0] _T_94829; // @[Modules.scala 56:109:@48139.4]
  wire [10:0] _T_94830; // @[Modules.scala 56:109:@48140.4]
  wire [10:0] buffer_12_709; // @[Modules.scala 56:109:@48141.4]
  wire [11:0] _T_94832; // @[Modules.scala 56:109:@48143.4]
  wire [10:0] _T_94833; // @[Modules.scala 56:109:@48144.4]
  wire [10:0] buffer_12_710; // @[Modules.scala 56:109:@48145.4]
  wire [11:0] _T_94835; // @[Modules.scala 56:109:@48147.4]
  wire [10:0] _T_94836; // @[Modules.scala 56:109:@48148.4]
  wire [10:0] buffer_12_711; // @[Modules.scala 56:109:@48149.4]
  wire [11:0] _T_94838; // @[Modules.scala 56:109:@48151.4]
  wire [10:0] _T_94839; // @[Modules.scala 56:109:@48152.4]
  wire [10:0] buffer_12_712; // @[Modules.scala 56:109:@48153.4]
  wire [11:0] _T_94841; // @[Modules.scala 56:109:@48155.4]
  wire [10:0] _T_94842; // @[Modules.scala 56:109:@48156.4]
  wire [10:0] buffer_12_713; // @[Modules.scala 56:109:@48157.4]
  wire [11:0] _T_94844; // @[Modules.scala 56:109:@48159.4]
  wire [10:0] _T_94845; // @[Modules.scala 56:109:@48160.4]
  wire [10:0] buffer_12_714; // @[Modules.scala 56:109:@48161.4]
  wire [11:0] _T_94847; // @[Modules.scala 56:109:@48163.4]
  wire [10:0] _T_94848; // @[Modules.scala 56:109:@48164.4]
  wire [10:0] buffer_12_715; // @[Modules.scala 56:109:@48165.4]
  wire [11:0] _T_94850; // @[Modules.scala 56:109:@48167.4]
  wire [10:0] _T_94851; // @[Modules.scala 56:109:@48168.4]
  wire [10:0] buffer_12_716; // @[Modules.scala 56:109:@48169.4]
  wire [11:0] _T_94853; // @[Modules.scala 56:109:@48171.4]
  wire [10:0] _T_94854; // @[Modules.scala 56:109:@48172.4]
  wire [10:0] buffer_12_717; // @[Modules.scala 56:109:@48173.4]
  wire [11:0] _T_94856; // @[Modules.scala 56:109:@48175.4]
  wire [10:0] _T_94857; // @[Modules.scala 56:109:@48176.4]
  wire [10:0] buffer_12_718; // @[Modules.scala 56:109:@48177.4]
  wire [11:0] _T_94859; // @[Modules.scala 56:109:@48179.4]
  wire [10:0] _T_94860; // @[Modules.scala 56:109:@48180.4]
  wire [10:0] buffer_12_719; // @[Modules.scala 56:109:@48181.4]
  wire [11:0] _T_94862; // @[Modules.scala 56:109:@48183.4]
  wire [10:0] _T_94863; // @[Modules.scala 56:109:@48184.4]
  wire [10:0] buffer_12_720; // @[Modules.scala 56:109:@48185.4]
  wire [11:0] _T_94865; // @[Modules.scala 56:109:@48187.4]
  wire [10:0] _T_94866; // @[Modules.scala 56:109:@48188.4]
  wire [10:0] buffer_12_721; // @[Modules.scala 56:109:@48189.4]
  wire [11:0] _T_94868; // @[Modules.scala 56:109:@48191.4]
  wire [10:0] _T_94869; // @[Modules.scala 56:109:@48192.4]
  wire [10:0] buffer_12_722; // @[Modules.scala 56:109:@48193.4]
  wire [11:0] _T_94871; // @[Modules.scala 56:109:@48195.4]
  wire [10:0] _T_94872; // @[Modules.scala 56:109:@48196.4]
  wire [10:0] buffer_12_723; // @[Modules.scala 56:109:@48197.4]
  wire [11:0] _T_94874; // @[Modules.scala 56:109:@48199.4]
  wire [10:0] _T_94875; // @[Modules.scala 56:109:@48200.4]
  wire [10:0] buffer_12_724; // @[Modules.scala 56:109:@48201.4]
  wire [11:0] _T_94877; // @[Modules.scala 56:109:@48203.4]
  wire [10:0] _T_94878; // @[Modules.scala 56:109:@48204.4]
  wire [10:0] buffer_12_725; // @[Modules.scala 56:109:@48205.4]
  wire [11:0] _T_94880; // @[Modules.scala 56:109:@48207.4]
  wire [10:0] _T_94881; // @[Modules.scala 56:109:@48208.4]
  wire [10:0] buffer_12_726; // @[Modules.scala 56:109:@48209.4]
  wire [11:0] _T_94883; // @[Modules.scala 56:109:@48211.4]
  wire [10:0] _T_94884; // @[Modules.scala 56:109:@48212.4]
  wire [10:0] buffer_12_727; // @[Modules.scala 56:109:@48213.4]
  wire [11:0] _T_94886; // @[Modules.scala 56:109:@48215.4]
  wire [10:0] _T_94887; // @[Modules.scala 56:109:@48216.4]
  wire [10:0] buffer_12_728; // @[Modules.scala 56:109:@48217.4]
  wire [11:0] _T_94889; // @[Modules.scala 56:109:@48219.4]
  wire [10:0] _T_94890; // @[Modules.scala 56:109:@48220.4]
  wire [10:0] buffer_12_729; // @[Modules.scala 56:109:@48221.4]
  wire [11:0] _T_94895; // @[Modules.scala 56:109:@48227.4]
  wire [10:0] _T_94896; // @[Modules.scala 56:109:@48228.4]
  wire [10:0] buffer_12_731; // @[Modules.scala 56:109:@48229.4]
  wire [11:0] _T_94901; // @[Modules.scala 56:109:@48235.4]
  wire [10:0] _T_94902; // @[Modules.scala 56:109:@48236.4]
  wire [10:0] buffer_12_733; // @[Modules.scala 56:109:@48237.4]
  wire [11:0] _T_94904; // @[Modules.scala 56:109:@48239.4]
  wire [10:0] _T_94905; // @[Modules.scala 56:109:@48240.4]
  wire [10:0] buffer_12_734; // @[Modules.scala 56:109:@48241.4]
  wire [11:0] _T_94907; // @[Modules.scala 63:156:@48244.4]
  wire [10:0] _T_94908; // @[Modules.scala 63:156:@48245.4]
  wire [10:0] buffer_12_736; // @[Modules.scala 63:156:@48246.4]
  wire [11:0] _T_94910; // @[Modules.scala 63:156:@48248.4]
  wire [10:0] _T_94911; // @[Modules.scala 63:156:@48249.4]
  wire [10:0] buffer_12_737; // @[Modules.scala 63:156:@48250.4]
  wire [11:0] _T_94913; // @[Modules.scala 63:156:@48252.4]
  wire [10:0] _T_94914; // @[Modules.scala 63:156:@48253.4]
  wire [10:0] buffer_12_738; // @[Modules.scala 63:156:@48254.4]
  wire [11:0] _T_94916; // @[Modules.scala 63:156:@48256.4]
  wire [10:0] _T_94917; // @[Modules.scala 63:156:@48257.4]
  wire [10:0] buffer_12_739; // @[Modules.scala 63:156:@48258.4]
  wire [11:0] _T_94919; // @[Modules.scala 63:156:@48260.4]
  wire [10:0] _T_94920; // @[Modules.scala 63:156:@48261.4]
  wire [10:0] buffer_12_740; // @[Modules.scala 63:156:@48262.4]
  wire [11:0] _T_94922; // @[Modules.scala 63:156:@48264.4]
  wire [10:0] _T_94923; // @[Modules.scala 63:156:@48265.4]
  wire [10:0] buffer_12_741; // @[Modules.scala 63:156:@48266.4]
  wire [11:0] _T_94925; // @[Modules.scala 63:156:@48268.4]
  wire [10:0] _T_94926; // @[Modules.scala 63:156:@48269.4]
  wire [10:0] buffer_12_742; // @[Modules.scala 63:156:@48270.4]
  wire [11:0] _T_94928; // @[Modules.scala 63:156:@48272.4]
  wire [10:0] _T_94929; // @[Modules.scala 63:156:@48273.4]
  wire [10:0] buffer_12_743; // @[Modules.scala 63:156:@48274.4]
  wire [11:0] _T_94931; // @[Modules.scala 63:156:@48276.4]
  wire [10:0] _T_94932; // @[Modules.scala 63:156:@48277.4]
  wire [10:0] buffer_12_744; // @[Modules.scala 63:156:@48278.4]
  wire [11:0] _T_94934; // @[Modules.scala 63:156:@48280.4]
  wire [10:0] _T_94935; // @[Modules.scala 63:156:@48281.4]
  wire [10:0] buffer_12_745; // @[Modules.scala 63:156:@48282.4]
  wire [11:0] _T_94937; // @[Modules.scala 63:156:@48284.4]
  wire [10:0] _T_94938; // @[Modules.scala 63:156:@48285.4]
  wire [10:0] buffer_12_746; // @[Modules.scala 63:156:@48286.4]
  wire [11:0] _T_94940; // @[Modules.scala 63:156:@48288.4]
  wire [10:0] _T_94941; // @[Modules.scala 63:156:@48289.4]
  wire [10:0] buffer_12_747; // @[Modules.scala 63:156:@48290.4]
  wire [11:0] _T_94943; // @[Modules.scala 63:156:@48292.4]
  wire [10:0] _T_94944; // @[Modules.scala 63:156:@48293.4]
  wire [10:0] buffer_12_748; // @[Modules.scala 63:156:@48294.4]
  wire [11:0] _T_94946; // @[Modules.scala 63:156:@48296.4]
  wire [10:0] _T_94947; // @[Modules.scala 63:156:@48297.4]
  wire [10:0] buffer_12_749; // @[Modules.scala 63:156:@48298.4]
  wire [11:0] _T_94949; // @[Modules.scala 63:156:@48300.4]
  wire [10:0] _T_94950; // @[Modules.scala 63:156:@48301.4]
  wire [10:0] buffer_12_750; // @[Modules.scala 63:156:@48302.4]
  wire [11:0] _T_94952; // @[Modules.scala 63:156:@48304.4]
  wire [10:0] _T_94953; // @[Modules.scala 63:156:@48305.4]
  wire [10:0] buffer_12_751; // @[Modules.scala 63:156:@48306.4]
  wire [11:0] _T_94955; // @[Modules.scala 63:156:@48308.4]
  wire [10:0] _T_94956; // @[Modules.scala 63:156:@48309.4]
  wire [10:0] buffer_12_752; // @[Modules.scala 63:156:@48310.4]
  wire [11:0] _T_94958; // @[Modules.scala 63:156:@48312.4]
  wire [10:0] _T_94959; // @[Modules.scala 63:156:@48313.4]
  wire [10:0] buffer_12_753; // @[Modules.scala 63:156:@48314.4]
  wire [11:0] _T_94961; // @[Modules.scala 63:156:@48316.4]
  wire [10:0] _T_94962; // @[Modules.scala 63:156:@48317.4]
  wire [10:0] buffer_12_754; // @[Modules.scala 63:156:@48318.4]
  wire [11:0] _T_94964; // @[Modules.scala 63:156:@48320.4]
  wire [10:0] _T_94965; // @[Modules.scala 63:156:@48321.4]
  wire [10:0] buffer_12_755; // @[Modules.scala 63:156:@48322.4]
  wire [11:0] _T_94967; // @[Modules.scala 63:156:@48324.4]
  wire [10:0] _T_94968; // @[Modules.scala 63:156:@48325.4]
  wire [10:0] buffer_12_756; // @[Modules.scala 63:156:@48326.4]
  wire [11:0] _T_94970; // @[Modules.scala 63:156:@48328.4]
  wire [10:0] _T_94971; // @[Modules.scala 63:156:@48329.4]
  wire [10:0] buffer_12_757; // @[Modules.scala 63:156:@48330.4]
  wire [11:0] _T_94973; // @[Modules.scala 63:156:@48332.4]
  wire [10:0] _T_94974; // @[Modules.scala 63:156:@48333.4]
  wire [10:0] buffer_12_758; // @[Modules.scala 63:156:@48334.4]
  wire [11:0] _T_94976; // @[Modules.scala 63:156:@48336.4]
  wire [10:0] _T_94977; // @[Modules.scala 63:156:@48337.4]
  wire [10:0] buffer_12_759; // @[Modules.scala 63:156:@48338.4]
  wire [11:0] _T_94979; // @[Modules.scala 63:156:@48340.4]
  wire [10:0] _T_94980; // @[Modules.scala 63:156:@48341.4]
  wire [10:0] buffer_12_760; // @[Modules.scala 63:156:@48342.4]
  wire [11:0] _T_94982; // @[Modules.scala 63:156:@48344.4]
  wire [10:0] _T_94983; // @[Modules.scala 63:156:@48345.4]
  wire [10:0] buffer_12_761; // @[Modules.scala 63:156:@48346.4]
  wire [11:0] _T_94985; // @[Modules.scala 63:156:@48348.4]
  wire [10:0] _T_94986; // @[Modules.scala 63:156:@48349.4]
  wire [10:0] buffer_12_762; // @[Modules.scala 63:156:@48350.4]
  wire [11:0] _T_94988; // @[Modules.scala 63:156:@48352.4]
  wire [10:0] _T_94989; // @[Modules.scala 63:156:@48353.4]
  wire [10:0] buffer_12_763; // @[Modules.scala 63:156:@48354.4]
  wire [11:0] _T_94991; // @[Modules.scala 63:156:@48356.4]
  wire [10:0] _T_94992; // @[Modules.scala 63:156:@48357.4]
  wire [10:0] buffer_12_764; // @[Modules.scala 63:156:@48358.4]
  wire [11:0] _T_94994; // @[Modules.scala 63:156:@48360.4]
  wire [10:0] _T_94995; // @[Modules.scala 63:156:@48361.4]
  wire [10:0] buffer_12_765; // @[Modules.scala 63:156:@48362.4]
  wire [11:0] _T_94997; // @[Modules.scala 63:156:@48364.4]
  wire [10:0] _T_94998; // @[Modules.scala 63:156:@48365.4]
  wire [10:0] buffer_12_766; // @[Modules.scala 63:156:@48366.4]
  wire [11:0] _T_95000; // @[Modules.scala 63:156:@48368.4]
  wire [10:0] _T_95001; // @[Modules.scala 63:156:@48369.4]
  wire [10:0] buffer_12_767; // @[Modules.scala 63:156:@48370.4]
  wire [11:0] _T_95003; // @[Modules.scala 63:156:@48372.4]
  wire [10:0] _T_95004; // @[Modules.scala 63:156:@48373.4]
  wire [10:0] buffer_12_768; // @[Modules.scala 63:156:@48374.4]
  wire [11:0] _T_95006; // @[Modules.scala 63:156:@48376.4]
  wire [10:0] _T_95007; // @[Modules.scala 63:156:@48377.4]
  wire [10:0] buffer_12_769; // @[Modules.scala 63:156:@48378.4]
  wire [11:0] _T_95009; // @[Modules.scala 63:156:@48380.4]
  wire [10:0] _T_95010; // @[Modules.scala 63:156:@48381.4]
  wire [10:0] buffer_12_770; // @[Modules.scala 63:156:@48382.4]
  wire [11:0] _T_95012; // @[Modules.scala 63:156:@48384.4]
  wire [10:0] _T_95013; // @[Modules.scala 63:156:@48385.4]
  wire [10:0] buffer_12_771; // @[Modules.scala 63:156:@48386.4]
  wire [11:0] _T_95015; // @[Modules.scala 63:156:@48388.4]
  wire [10:0] _T_95016; // @[Modules.scala 63:156:@48389.4]
  wire [10:0] buffer_12_772; // @[Modules.scala 63:156:@48390.4]
  wire [11:0] _T_95018; // @[Modules.scala 63:156:@48392.4]
  wire [10:0] _T_95019; // @[Modules.scala 63:156:@48393.4]
  wire [10:0] buffer_12_773; // @[Modules.scala 63:156:@48394.4]
  wire [11:0] _T_95021; // @[Modules.scala 63:156:@48396.4]
  wire [10:0] _T_95022; // @[Modules.scala 63:156:@48397.4]
  wire [10:0] buffer_12_774; // @[Modules.scala 63:156:@48398.4]
  wire [11:0] _T_95024; // @[Modules.scala 63:156:@48400.4]
  wire [10:0] _T_95025; // @[Modules.scala 63:156:@48401.4]
  wire [10:0] buffer_12_775; // @[Modules.scala 63:156:@48402.4]
  wire [11:0] _T_95027; // @[Modules.scala 63:156:@48404.4]
  wire [10:0] _T_95028; // @[Modules.scala 63:156:@48405.4]
  wire [10:0] buffer_12_776; // @[Modules.scala 63:156:@48406.4]
  wire [11:0] _T_95030; // @[Modules.scala 63:156:@48408.4]
  wire [10:0] _T_95031; // @[Modules.scala 63:156:@48409.4]
  wire [10:0] buffer_12_777; // @[Modules.scala 63:156:@48410.4]
  wire [11:0] _T_95033; // @[Modules.scala 63:156:@48412.4]
  wire [10:0] _T_95034; // @[Modules.scala 63:156:@48413.4]
  wire [10:0] buffer_12_778; // @[Modules.scala 63:156:@48414.4]
  wire [11:0] _T_95036; // @[Modules.scala 63:156:@48416.4]
  wire [10:0] _T_95037; // @[Modules.scala 63:156:@48417.4]
  wire [10:0] buffer_12_779; // @[Modules.scala 63:156:@48418.4]
  wire [11:0] _T_95039; // @[Modules.scala 63:156:@48420.4]
  wire [10:0] _T_95040; // @[Modules.scala 63:156:@48421.4]
  wire [10:0] buffer_12_780; // @[Modules.scala 63:156:@48422.4]
  wire [11:0] _T_95042; // @[Modules.scala 63:156:@48424.4]
  wire [10:0] _T_95043; // @[Modules.scala 63:156:@48425.4]
  wire [10:0] buffer_12_781; // @[Modules.scala 63:156:@48426.4]
  wire [11:0] _T_95045; // @[Modules.scala 63:156:@48428.4]
  wire [10:0] _T_95046; // @[Modules.scala 63:156:@48429.4]
  wire [10:0] buffer_12_782; // @[Modules.scala 63:156:@48430.4]
  wire [11:0] _T_95048; // @[Modules.scala 63:156:@48432.4]
  wire [10:0] _T_95049; // @[Modules.scala 63:156:@48433.4]
  wire [10:0] buffer_12_783; // @[Modules.scala 63:156:@48434.4]
  wire [5:0] _T_95085; // @[Modules.scala 40:46:@48473.4]
  wire [4:0] _T_95086; // @[Modules.scala 40:46:@48474.4]
  wire [4:0] _T_95087; // @[Modules.scala 40:46:@48475.4]
  wire [5:0] _T_95149; // @[Modules.scala 40:46:@48542.4]
  wire [4:0] _T_95150; // @[Modules.scala 40:46:@48543.4]
  wire [4:0] _T_95151; // @[Modules.scala 40:46:@48544.4]
  wire [5:0] _T_95236; // @[Modules.scala 40:46:@48637.4]
  wire [4:0] _T_95237; // @[Modules.scala 40:46:@48638.4]
  wire [4:0] _T_95238; // @[Modules.scala 40:46:@48639.4]
  wire [5:0] _T_95255; // @[Modules.scala 40:46:@48660.4]
  wire [4:0] _T_95256; // @[Modules.scala 40:46:@48661.4]
  wire [4:0] _T_95257; // @[Modules.scala 40:46:@48662.4]
  wire [5:0] _T_95448; // @[Modules.scala 40:46:@48873.4]
  wire [4:0] _T_95449; // @[Modules.scala 40:46:@48874.4]
  wire [4:0] _T_95450; // @[Modules.scala 40:46:@48875.4]
  wire [5:0] _T_95482; // @[Modules.scala 40:46:@48909.4]
  wire [4:0] _T_95483; // @[Modules.scala 40:46:@48910.4]
  wire [4:0] _T_95484; // @[Modules.scala 40:46:@48911.4]
  wire [5:0] _T_95513; // @[Modules.scala 40:46:@48941.4]
  wire [4:0] _T_95514; // @[Modules.scala 40:46:@48942.4]
  wire [4:0] _T_95515; // @[Modules.scala 40:46:@48943.4]
  wire [5:0] _T_95530; // @[Modules.scala 43:47:@48959.4]
  wire [4:0] _T_95531; // @[Modules.scala 43:47:@48960.4]
  wire [4:0] _T_95532; // @[Modules.scala 43:47:@48961.4]
  wire [5:0] _T_95671; // @[Modules.scala 40:46:@49112.4]
  wire [4:0] _T_95672; // @[Modules.scala 40:46:@49113.4]
  wire [4:0] _T_95673; // @[Modules.scala 40:46:@49114.4]
  wire [5:0] _T_95747; // @[Modules.scala 40:46:@49190.4]
  wire [4:0] _T_95748; // @[Modules.scala 40:46:@49191.4]
  wire [4:0] _T_95749; // @[Modules.scala 40:46:@49192.4]
  wire [5:0] _T_95822; // @[Modules.scala 43:47:@49269.4]
  wire [4:0] _T_95823; // @[Modules.scala 43:47:@49270.4]
  wire [4:0] _T_95824; // @[Modules.scala 43:47:@49271.4]
  wire [5:0] _T_95889; // @[Modules.scala 40:46:@49342.4]
  wire [4:0] _T_95890; // @[Modules.scala 40:46:@49343.4]
  wire [4:0] _T_95891; // @[Modules.scala 40:46:@49344.4]
  wire [5:0] _T_95952; // @[Modules.scala 40:46:@49412.4]
  wire [4:0] _T_95953; // @[Modules.scala 40:46:@49413.4]
  wire [4:0] _T_95954; // @[Modules.scala 40:46:@49414.4]
  wire [5:0] _T_95959; // @[Modules.scala 43:47:@49419.4]
  wire [4:0] _T_95960; // @[Modules.scala 43:47:@49420.4]
  wire [4:0] _T_95961; // @[Modules.scala 43:47:@49421.4]
  wire [5:0] _T_95969; // @[Modules.scala 40:46:@49430.4]
  wire [4:0] _T_95970; // @[Modules.scala 40:46:@49431.4]
  wire [4:0] _T_95971; // @[Modules.scala 40:46:@49432.4]
  wire [5:0] _T_95983; // @[Modules.scala 43:47:@49444.4]
  wire [4:0] _T_95984; // @[Modules.scala 43:47:@49445.4]
  wire [4:0] _T_95985; // @[Modules.scala 43:47:@49446.4]
  wire [5:0] _T_96303; // @[Modules.scala 40:46:@49810.4]
  wire [4:0] _T_96304; // @[Modules.scala 40:46:@49811.4]
  wire [4:0] _T_96305; // @[Modules.scala 40:46:@49812.4]
  wire [5:0] _T_96378; // @[Modules.scala 40:46:@49896.4]
  wire [4:0] _T_96379; // @[Modules.scala 40:46:@49897.4]
  wire [4:0] _T_96380; // @[Modules.scala 40:46:@49898.4]
  wire [5:0] _T_96461; // @[Modules.scala 43:47:@49988.4]
  wire [4:0] _T_96462; // @[Modules.scala 43:47:@49989.4]
  wire [4:0] _T_96463; // @[Modules.scala 43:47:@49990.4]
  wire [5:0] _T_96602; // @[Modules.scala 40:46:@50141.4]
  wire [4:0] _T_96603; // @[Modules.scala 40:46:@50142.4]
  wire [4:0] _T_96604; // @[Modules.scala 40:46:@50143.4]
  wire [5:0] _T_96654; // @[Modules.scala 46:47:@50201.4]
  wire [4:0] _T_96655; // @[Modules.scala 46:47:@50202.4]
  wire [4:0] _T_96656; // @[Modules.scala 46:47:@50203.4]
  wire [5:0] _T_96706; // @[Modules.scala 43:47:@50254.4]
  wire [4:0] _T_96707; // @[Modules.scala 43:47:@50255.4]
  wire [4:0] _T_96708; // @[Modules.scala 43:47:@50256.4]
  wire [5:0] _T_97076; // @[Modules.scala 40:46:@50640.4]
  wire [4:0] _T_97077; // @[Modules.scala 40:46:@50641.4]
  wire [4:0] _T_97078; // @[Modules.scala 40:46:@50642.4]
  wire [11:0] _T_97079; // @[Modules.scala 50:57:@50644.4]
  wire [10:0] _T_97080; // @[Modules.scala 50:57:@50645.4]
  wire [10:0] buffer_13_392; // @[Modules.scala 50:57:@50646.4]
  wire [10:0] buffer_13_6; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97088; // @[Modules.scala 50:57:@50656.4]
  wire [10:0] _T_97089; // @[Modules.scala 50:57:@50657.4]
  wire [10:0] buffer_13_395; // @[Modules.scala 50:57:@50658.4]
  wire [11:0] _T_97097; // @[Modules.scala 50:57:@50668.4]
  wire [10:0] _T_97098; // @[Modules.scala 50:57:@50669.4]
  wire [10:0] buffer_13_398; // @[Modules.scala 50:57:@50670.4]
  wire [11:0] _T_97100; // @[Modules.scala 50:57:@50672.4]
  wire [10:0] _T_97101; // @[Modules.scala 50:57:@50673.4]
  wire [10:0] buffer_13_399; // @[Modules.scala 50:57:@50674.4]
  wire [10:0] buffer_13_18; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97106; // @[Modules.scala 50:57:@50680.4]
  wire [10:0] _T_97107; // @[Modules.scala 50:57:@50681.4]
  wire [10:0] buffer_13_401; // @[Modules.scala 50:57:@50682.4]
  wire [11:0] _T_97118; // @[Modules.scala 50:57:@50696.4]
  wire [10:0] _T_97119; // @[Modules.scala 50:57:@50697.4]
  wire [10:0] buffer_13_405; // @[Modules.scala 50:57:@50698.4]
  wire [10:0] buffer_13_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97130; // @[Modules.scala 50:57:@50712.4]
  wire [10:0] _T_97131; // @[Modules.scala 50:57:@50713.4]
  wire [10:0] buffer_13_409; // @[Modules.scala 50:57:@50714.4]
  wire [11:0] _T_97133; // @[Modules.scala 50:57:@50716.4]
  wire [10:0] _T_97134; // @[Modules.scala 50:57:@50717.4]
  wire [10:0] buffer_13_410; // @[Modules.scala 50:57:@50718.4]
  wire [10:0] buffer_13_40; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97139; // @[Modules.scala 50:57:@50724.4]
  wire [10:0] _T_97140; // @[Modules.scala 50:57:@50725.4]
  wire [10:0] buffer_13_412; // @[Modules.scala 50:57:@50726.4]
  wire [11:0] _T_97151; // @[Modules.scala 50:57:@50740.4]
  wire [10:0] _T_97152; // @[Modules.scala 50:57:@50741.4]
  wire [10:0] buffer_13_416; // @[Modules.scala 50:57:@50742.4]
  wire [11:0] _T_97169; // @[Modules.scala 50:57:@50764.4]
  wire [10:0] _T_97170; // @[Modules.scala 50:57:@50765.4]
  wire [10:0] buffer_13_422; // @[Modules.scala 50:57:@50766.4]
  wire [10:0] buffer_13_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97196; // @[Modules.scala 50:57:@50800.4]
  wire [10:0] _T_97197; // @[Modules.scala 50:57:@50801.4]
  wire [10:0] buffer_13_431; // @[Modules.scala 50:57:@50802.4]
  wire [11:0] _T_97199; // @[Modules.scala 50:57:@50804.4]
  wire [10:0] _T_97200; // @[Modules.scala 50:57:@50805.4]
  wire [10:0] buffer_13_432; // @[Modules.scala 50:57:@50806.4]
  wire [10:0] buffer_13_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97205; // @[Modules.scala 50:57:@50812.4]
  wire [10:0] _T_97206; // @[Modules.scala 50:57:@50813.4]
  wire [10:0] buffer_13_434; // @[Modules.scala 50:57:@50814.4]
  wire [10:0] buffer_13_90; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97214; // @[Modules.scala 50:57:@50824.4]
  wire [10:0] _T_97215; // @[Modules.scala 50:57:@50825.4]
  wire [10:0] buffer_13_437; // @[Modules.scala 50:57:@50826.4]
  wire [10:0] buffer_13_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97217; // @[Modules.scala 50:57:@50828.4]
  wire [10:0] _T_97218; // @[Modules.scala 50:57:@50829.4]
  wire [10:0] buffer_13_438; // @[Modules.scala 50:57:@50830.4]
  wire [11:0] _T_97220; // @[Modules.scala 50:57:@50832.4]
  wire [10:0] _T_97221; // @[Modules.scala 50:57:@50833.4]
  wire [10:0] buffer_13_439; // @[Modules.scala 50:57:@50834.4]
  wire [11:0] _T_97226; // @[Modules.scala 50:57:@50840.4]
  wire [10:0] _T_97227; // @[Modules.scala 50:57:@50841.4]
  wire [10:0] buffer_13_441; // @[Modules.scala 50:57:@50842.4]
  wire [11:0] _T_97229; // @[Modules.scala 50:57:@50844.4]
  wire [10:0] _T_97230; // @[Modules.scala 50:57:@50845.4]
  wire [10:0] buffer_13_442; // @[Modules.scala 50:57:@50846.4]
  wire [11:0] _T_97235; // @[Modules.scala 50:57:@50852.4]
  wire [10:0] _T_97236; // @[Modules.scala 50:57:@50853.4]
  wire [10:0] buffer_13_444; // @[Modules.scala 50:57:@50854.4]
  wire [11:0] _T_97247; // @[Modules.scala 50:57:@50868.4]
  wire [10:0] _T_97248; // @[Modules.scala 50:57:@50869.4]
  wire [10:0] buffer_13_448; // @[Modules.scala 50:57:@50870.4]
  wire [11:0] _T_97250; // @[Modules.scala 50:57:@50872.4]
  wire [10:0] _T_97251; // @[Modules.scala 50:57:@50873.4]
  wire [10:0] buffer_13_449; // @[Modules.scala 50:57:@50874.4]
  wire [10:0] buffer_13_120; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97259; // @[Modules.scala 50:57:@50884.4]
  wire [10:0] _T_97260; // @[Modules.scala 50:57:@50885.4]
  wire [10:0] buffer_13_452; // @[Modules.scala 50:57:@50886.4]
  wire [11:0] _T_97274; // @[Modules.scala 50:57:@50904.4]
  wire [10:0] _T_97275; // @[Modules.scala 50:57:@50905.4]
  wire [10:0] buffer_13_457; // @[Modules.scala 50:57:@50906.4]
  wire [10:0] buffer_13_132; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97277; // @[Modules.scala 50:57:@50908.4]
  wire [10:0] _T_97278; // @[Modules.scala 50:57:@50909.4]
  wire [10:0] buffer_13_458; // @[Modules.scala 50:57:@50910.4]
  wire [11:0] _T_97283; // @[Modules.scala 50:57:@50916.4]
  wire [10:0] _T_97284; // @[Modules.scala 50:57:@50917.4]
  wire [10:0] buffer_13_460; // @[Modules.scala 50:57:@50918.4]
  wire [10:0] buffer_13_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97295; // @[Modules.scala 50:57:@50932.4]
  wire [10:0] _T_97296; // @[Modules.scala 50:57:@50933.4]
  wire [10:0] buffer_13_464; // @[Modules.scala 50:57:@50934.4]
  wire [11:0] _T_97301; // @[Modules.scala 50:57:@50940.4]
  wire [10:0] _T_97302; // @[Modules.scala 50:57:@50941.4]
  wire [10:0] buffer_13_466; // @[Modules.scala 50:57:@50942.4]
  wire [11:0] _T_97304; // @[Modules.scala 50:57:@50944.4]
  wire [10:0] _T_97305; // @[Modules.scala 50:57:@50945.4]
  wire [10:0] buffer_13_467; // @[Modules.scala 50:57:@50946.4]
  wire [11:0] _T_97313; // @[Modules.scala 50:57:@50956.4]
  wire [10:0] _T_97314; // @[Modules.scala 50:57:@50957.4]
  wire [10:0] buffer_13_470; // @[Modules.scala 50:57:@50958.4]
  wire [10:0] buffer_13_158; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97316; // @[Modules.scala 50:57:@50960.4]
  wire [10:0] _T_97317; // @[Modules.scala 50:57:@50961.4]
  wire [10:0] buffer_13_471; // @[Modules.scala 50:57:@50962.4]
  wire [11:0] _T_97322; // @[Modules.scala 50:57:@50968.4]
  wire [10:0] _T_97323; // @[Modules.scala 50:57:@50969.4]
  wire [10:0] buffer_13_473; // @[Modules.scala 50:57:@50970.4]
  wire [11:0] _T_97331; // @[Modules.scala 50:57:@50980.4]
  wire [10:0] _T_97332; // @[Modules.scala 50:57:@50981.4]
  wire [10:0] buffer_13_476; // @[Modules.scala 50:57:@50982.4]
  wire [10:0] buffer_13_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97334; // @[Modules.scala 50:57:@50984.4]
  wire [10:0] _T_97335; // @[Modules.scala 50:57:@50985.4]
  wire [10:0] buffer_13_477; // @[Modules.scala 50:57:@50986.4]
  wire [10:0] buffer_13_172; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97337; // @[Modules.scala 50:57:@50988.4]
  wire [10:0] _T_97338; // @[Modules.scala 50:57:@50989.4]
  wire [10:0] buffer_13_478; // @[Modules.scala 50:57:@50990.4]
  wire [10:0] buffer_13_174; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97340; // @[Modules.scala 50:57:@50992.4]
  wire [10:0] _T_97341; // @[Modules.scala 50:57:@50993.4]
  wire [10:0] buffer_13_479; // @[Modules.scala 50:57:@50994.4]
  wire [10:0] buffer_13_176; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97343; // @[Modules.scala 50:57:@50996.4]
  wire [10:0] _T_97344; // @[Modules.scala 50:57:@50997.4]
  wire [10:0] buffer_13_480; // @[Modules.scala 50:57:@50998.4]
  wire [11:0] _T_97352; // @[Modules.scala 50:57:@51008.4]
  wire [10:0] _T_97353; // @[Modules.scala 50:57:@51009.4]
  wire [10:0] buffer_13_483; // @[Modules.scala 50:57:@51010.4]
  wire [11:0] _T_97358; // @[Modules.scala 50:57:@51016.4]
  wire [10:0] _T_97359; // @[Modules.scala 50:57:@51017.4]
  wire [10:0] buffer_13_485; // @[Modules.scala 50:57:@51018.4]
  wire [11:0] _T_97364; // @[Modules.scala 50:57:@51024.4]
  wire [10:0] _T_97365; // @[Modules.scala 50:57:@51025.4]
  wire [10:0] buffer_13_487; // @[Modules.scala 50:57:@51026.4]
  wire [11:0] _T_97367; // @[Modules.scala 50:57:@51028.4]
  wire [10:0] _T_97368; // @[Modules.scala 50:57:@51029.4]
  wire [10:0] buffer_13_488; // @[Modules.scala 50:57:@51030.4]
  wire [11:0] _T_97382; // @[Modules.scala 50:57:@51048.4]
  wire [10:0] _T_97383; // @[Modules.scala 50:57:@51049.4]
  wire [10:0] buffer_13_493; // @[Modules.scala 50:57:@51050.4]
  wire [11:0] _T_97385; // @[Modules.scala 50:57:@51052.4]
  wire [10:0] _T_97386; // @[Modules.scala 50:57:@51053.4]
  wire [10:0] buffer_13_494; // @[Modules.scala 50:57:@51054.4]
  wire [11:0] _T_97394; // @[Modules.scala 50:57:@51064.4]
  wire [10:0] _T_97395; // @[Modules.scala 50:57:@51065.4]
  wire [10:0] buffer_13_497; // @[Modules.scala 50:57:@51066.4]
  wire [11:0] _T_97415; // @[Modules.scala 50:57:@51092.4]
  wire [10:0] _T_97416; // @[Modules.scala 50:57:@51093.4]
  wire [10:0] buffer_13_504; // @[Modules.scala 50:57:@51094.4]
  wire [11:0] _T_97424; // @[Modules.scala 50:57:@51104.4]
  wire [10:0] _T_97425; // @[Modules.scala 50:57:@51105.4]
  wire [10:0] buffer_13_507; // @[Modules.scala 50:57:@51106.4]
  wire [11:0] _T_97427; // @[Modules.scala 50:57:@51108.4]
  wire [10:0] _T_97428; // @[Modules.scala 50:57:@51109.4]
  wire [10:0] buffer_13_508; // @[Modules.scala 50:57:@51110.4]
  wire [11:0] _T_97430; // @[Modules.scala 50:57:@51112.4]
  wire [10:0] _T_97431; // @[Modules.scala 50:57:@51113.4]
  wire [10:0] buffer_13_509; // @[Modules.scala 50:57:@51114.4]
  wire [11:0] _T_97439; // @[Modules.scala 50:57:@51124.4]
  wire [10:0] _T_97440; // @[Modules.scala 50:57:@51125.4]
  wire [10:0] buffer_13_512; // @[Modules.scala 50:57:@51126.4]
  wire [11:0] _T_97448; // @[Modules.scala 50:57:@51136.4]
  wire [10:0] _T_97449; // @[Modules.scala 50:57:@51137.4]
  wire [10:0] buffer_13_515; // @[Modules.scala 50:57:@51138.4]
  wire [10:0] buffer_13_248; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97451; // @[Modules.scala 50:57:@51140.4]
  wire [10:0] _T_97452; // @[Modules.scala 50:57:@51141.4]
  wire [10:0] buffer_13_516; // @[Modules.scala 50:57:@51142.4]
  wire [11:0] _T_97469; // @[Modules.scala 50:57:@51164.4]
  wire [10:0] _T_97470; // @[Modules.scala 50:57:@51165.4]
  wire [10:0] buffer_13_522; // @[Modules.scala 50:57:@51166.4]
  wire [11:0] _T_97472; // @[Modules.scala 50:57:@51168.4]
  wire [10:0] _T_97473; // @[Modules.scala 50:57:@51169.4]
  wire [10:0] buffer_13_523; // @[Modules.scala 50:57:@51170.4]
  wire [10:0] buffer_13_265; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97475; // @[Modules.scala 50:57:@51172.4]
  wire [10:0] _T_97476; // @[Modules.scala 50:57:@51173.4]
  wire [10:0] buffer_13_524; // @[Modules.scala 50:57:@51174.4]
  wire [11:0] _T_97481; // @[Modules.scala 50:57:@51180.4]
  wire [10:0] _T_97482; // @[Modules.scala 50:57:@51181.4]
  wire [10:0] buffer_13_526; // @[Modules.scala 50:57:@51182.4]
  wire [11:0] _T_97487; // @[Modules.scala 50:57:@51188.4]
  wire [10:0] _T_97488; // @[Modules.scala 50:57:@51189.4]
  wire [10:0] buffer_13_528; // @[Modules.scala 50:57:@51190.4]
  wire [11:0] _T_97499; // @[Modules.scala 50:57:@51204.4]
  wire [10:0] _T_97500; // @[Modules.scala 50:57:@51205.4]
  wire [10:0] buffer_13_532; // @[Modules.scala 50:57:@51206.4]
  wire [10:0] buffer_13_282; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97502; // @[Modules.scala 50:57:@51208.4]
  wire [10:0] _T_97503; // @[Modules.scala 50:57:@51209.4]
  wire [10:0] buffer_13_533; // @[Modules.scala 50:57:@51210.4]
  wire [11:0] _T_97514; // @[Modules.scala 50:57:@51224.4]
  wire [10:0] _T_97515; // @[Modules.scala 50:57:@51225.4]
  wire [10:0] buffer_13_537; // @[Modules.scala 50:57:@51226.4]
  wire [11:0] _T_97517; // @[Modules.scala 50:57:@51228.4]
  wire [10:0] _T_97518; // @[Modules.scala 50:57:@51229.4]
  wire [10:0] buffer_13_538; // @[Modules.scala 50:57:@51230.4]
  wire [11:0] _T_97523; // @[Modules.scala 50:57:@51236.4]
  wire [10:0] _T_97524; // @[Modules.scala 50:57:@51237.4]
  wire [10:0] buffer_13_540; // @[Modules.scala 50:57:@51238.4]
  wire [10:0] buffer_13_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97541; // @[Modules.scala 50:57:@51260.4]
  wire [10:0] _T_97542; // @[Modules.scala 50:57:@51261.4]
  wire [10:0] buffer_13_546; // @[Modules.scala 50:57:@51262.4]
  wire [11:0] _T_97544; // @[Modules.scala 50:57:@51264.4]
  wire [10:0] _T_97545; // @[Modules.scala 50:57:@51265.4]
  wire [10:0] buffer_13_547; // @[Modules.scala 50:57:@51266.4]
  wire [11:0] _T_97547; // @[Modules.scala 50:57:@51268.4]
  wire [10:0] _T_97548; // @[Modules.scala 50:57:@51269.4]
  wire [10:0] buffer_13_548; // @[Modules.scala 50:57:@51270.4]
  wire [11:0] _T_97550; // @[Modules.scala 50:57:@51272.4]
  wire [10:0] _T_97551; // @[Modules.scala 50:57:@51273.4]
  wire [10:0] buffer_13_549; // @[Modules.scala 50:57:@51274.4]
  wire [11:0] _T_97553; // @[Modules.scala 50:57:@51276.4]
  wire [10:0] _T_97554; // @[Modules.scala 50:57:@51277.4]
  wire [10:0] buffer_13_550; // @[Modules.scala 50:57:@51278.4]
  wire [10:0] buffer_13_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97559; // @[Modules.scala 50:57:@51284.4]
  wire [10:0] _T_97560; // @[Modules.scala 50:57:@51285.4]
  wire [10:0] buffer_13_552; // @[Modules.scala 50:57:@51286.4]
  wire [10:0] buffer_13_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97571; // @[Modules.scala 50:57:@51300.4]
  wire [10:0] _T_97572; // @[Modules.scala 50:57:@51301.4]
  wire [10:0] buffer_13_556; // @[Modules.scala 50:57:@51302.4]
  wire [11:0] _T_97583; // @[Modules.scala 50:57:@51316.4]
  wire [10:0] _T_97584; // @[Modules.scala 50:57:@51317.4]
  wire [10:0] buffer_13_560; // @[Modules.scala 50:57:@51318.4]
  wire [11:0] _T_97592; // @[Modules.scala 50:57:@51328.4]
  wire [10:0] _T_97593; // @[Modules.scala 50:57:@51329.4]
  wire [10:0] buffer_13_563; // @[Modules.scala 50:57:@51330.4]
  wire [11:0] _T_97604; // @[Modules.scala 50:57:@51344.4]
  wire [10:0] _T_97605; // @[Modules.scala 50:57:@51345.4]
  wire [10:0] buffer_13_567; // @[Modules.scala 50:57:@51346.4]
  wire [11:0] _T_97625; // @[Modules.scala 50:57:@51372.4]
  wire [10:0] _T_97626; // @[Modules.scala 50:57:@51373.4]
  wire [10:0] buffer_13_574; // @[Modules.scala 50:57:@51374.4]
  wire [11:0] _T_97646; // @[Modules.scala 50:57:@51400.4]
  wire [10:0] _T_97647; // @[Modules.scala 50:57:@51401.4]
  wire [10:0] buffer_13_581; // @[Modules.scala 50:57:@51402.4]
  wire [10:0] buffer_13_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_97664; // @[Modules.scala 50:57:@51424.4]
  wire [10:0] _T_97665; // @[Modules.scala 50:57:@51425.4]
  wire [10:0] buffer_13_587; // @[Modules.scala 50:57:@51426.4]
  wire [11:0] _T_97667; // @[Modules.scala 53:83:@51428.4]
  wire [10:0] _T_97668; // @[Modules.scala 53:83:@51429.4]
  wire [10:0] buffer_13_588; // @[Modules.scala 53:83:@51430.4]
  wire [11:0] _T_97670; // @[Modules.scala 53:83:@51432.4]
  wire [10:0] _T_97671; // @[Modules.scala 53:83:@51433.4]
  wire [10:0] buffer_13_589; // @[Modules.scala 53:83:@51434.4]
  wire [11:0] _T_97673; // @[Modules.scala 53:83:@51436.4]
  wire [10:0] _T_97674; // @[Modules.scala 53:83:@51437.4]
  wire [10:0] buffer_13_590; // @[Modules.scala 53:83:@51438.4]
  wire [11:0] _T_97676; // @[Modules.scala 53:83:@51440.4]
  wire [10:0] _T_97677; // @[Modules.scala 53:83:@51441.4]
  wire [10:0] buffer_13_591; // @[Modules.scala 53:83:@51442.4]
  wire [11:0] _T_97679; // @[Modules.scala 53:83:@51444.4]
  wire [10:0] _T_97680; // @[Modules.scala 53:83:@51445.4]
  wire [10:0] buffer_13_592; // @[Modules.scala 53:83:@51446.4]
  wire [11:0] _T_97682; // @[Modules.scala 53:83:@51448.4]
  wire [10:0] _T_97683; // @[Modules.scala 53:83:@51449.4]
  wire [10:0] buffer_13_593; // @[Modules.scala 53:83:@51450.4]
  wire [11:0] _T_97685; // @[Modules.scala 53:83:@51452.4]
  wire [10:0] _T_97686; // @[Modules.scala 53:83:@51453.4]
  wire [10:0] buffer_13_594; // @[Modules.scala 53:83:@51454.4]
  wire [11:0] _T_97688; // @[Modules.scala 53:83:@51456.4]
  wire [10:0] _T_97689; // @[Modules.scala 53:83:@51457.4]
  wire [10:0] buffer_13_595; // @[Modules.scala 53:83:@51458.4]
  wire [11:0] _T_97691; // @[Modules.scala 53:83:@51460.4]
  wire [10:0] _T_97692; // @[Modules.scala 53:83:@51461.4]
  wire [10:0] buffer_13_596; // @[Modules.scala 53:83:@51462.4]
  wire [11:0] _T_97694; // @[Modules.scala 53:83:@51464.4]
  wire [10:0] _T_97695; // @[Modules.scala 53:83:@51465.4]
  wire [10:0] buffer_13_597; // @[Modules.scala 53:83:@51466.4]
  wire [11:0] _T_97697; // @[Modules.scala 53:83:@51468.4]
  wire [10:0] _T_97698; // @[Modules.scala 53:83:@51469.4]
  wire [10:0] buffer_13_598; // @[Modules.scala 53:83:@51470.4]
  wire [11:0] _T_97703; // @[Modules.scala 53:83:@51476.4]
  wire [10:0] _T_97704; // @[Modules.scala 53:83:@51477.4]
  wire [10:0] buffer_13_600; // @[Modules.scala 53:83:@51478.4]
  wire [11:0] _T_97709; // @[Modules.scala 53:83:@51484.4]
  wire [10:0] _T_97710; // @[Modules.scala 53:83:@51485.4]
  wire [10:0] buffer_13_602; // @[Modules.scala 53:83:@51486.4]
  wire [11:0] _T_97712; // @[Modules.scala 53:83:@51488.4]
  wire [10:0] _T_97713; // @[Modules.scala 53:83:@51489.4]
  wire [10:0] buffer_13_603; // @[Modules.scala 53:83:@51490.4]
  wire [11:0] _T_97718; // @[Modules.scala 53:83:@51496.4]
  wire [10:0] _T_97719; // @[Modules.scala 53:83:@51497.4]
  wire [10:0] buffer_13_605; // @[Modules.scala 53:83:@51498.4]
  wire [11:0] _T_97721; // @[Modules.scala 53:83:@51500.4]
  wire [10:0] _T_97722; // @[Modules.scala 53:83:@51501.4]
  wire [10:0] buffer_13_606; // @[Modules.scala 53:83:@51502.4]
  wire [11:0] _T_97724; // @[Modules.scala 53:83:@51504.4]
  wire [10:0] _T_97725; // @[Modules.scala 53:83:@51505.4]
  wire [10:0] buffer_13_607; // @[Modules.scala 53:83:@51506.4]
  wire [11:0] _T_97727; // @[Modules.scala 53:83:@51508.4]
  wire [10:0] _T_97728; // @[Modules.scala 53:83:@51509.4]
  wire [10:0] buffer_13_608; // @[Modules.scala 53:83:@51510.4]
  wire [11:0] _T_97730; // @[Modules.scala 53:83:@51512.4]
  wire [10:0] _T_97731; // @[Modules.scala 53:83:@51513.4]
  wire [10:0] buffer_13_609; // @[Modules.scala 53:83:@51514.4]
  wire [11:0] _T_97733; // @[Modules.scala 53:83:@51516.4]
  wire [10:0] _T_97734; // @[Modules.scala 53:83:@51517.4]
  wire [10:0] buffer_13_610; // @[Modules.scala 53:83:@51518.4]
  wire [11:0] _T_97736; // @[Modules.scala 53:83:@51520.4]
  wire [10:0] _T_97737; // @[Modules.scala 53:83:@51521.4]
  wire [10:0] buffer_13_611; // @[Modules.scala 53:83:@51522.4]
  wire [11:0] _T_97739; // @[Modules.scala 53:83:@51524.4]
  wire [10:0] _T_97740; // @[Modules.scala 53:83:@51525.4]
  wire [10:0] buffer_13_612; // @[Modules.scala 53:83:@51526.4]
  wire [11:0] _T_97742; // @[Modules.scala 53:83:@51528.4]
  wire [10:0] _T_97743; // @[Modules.scala 53:83:@51529.4]
  wire [10:0] buffer_13_613; // @[Modules.scala 53:83:@51530.4]
  wire [11:0] _T_97745; // @[Modules.scala 53:83:@51532.4]
  wire [10:0] _T_97746; // @[Modules.scala 53:83:@51533.4]
  wire [10:0] buffer_13_614; // @[Modules.scala 53:83:@51534.4]
  wire [11:0] _T_97748; // @[Modules.scala 53:83:@51536.4]
  wire [10:0] _T_97749; // @[Modules.scala 53:83:@51537.4]
  wire [10:0] buffer_13_615; // @[Modules.scala 53:83:@51538.4]
  wire [11:0] _T_97751; // @[Modules.scala 53:83:@51540.4]
  wire [10:0] _T_97752; // @[Modules.scala 53:83:@51541.4]
  wire [10:0] buffer_13_616; // @[Modules.scala 53:83:@51542.4]
  wire [11:0] _T_97754; // @[Modules.scala 53:83:@51544.4]
  wire [10:0] _T_97755; // @[Modules.scala 53:83:@51545.4]
  wire [10:0] buffer_13_617; // @[Modules.scala 53:83:@51546.4]
  wire [11:0] _T_97757; // @[Modules.scala 53:83:@51548.4]
  wire [10:0] _T_97758; // @[Modules.scala 53:83:@51549.4]
  wire [10:0] buffer_13_618; // @[Modules.scala 53:83:@51550.4]
  wire [11:0] _T_97763; // @[Modules.scala 53:83:@51556.4]
  wire [10:0] _T_97764; // @[Modules.scala 53:83:@51557.4]
  wire [10:0] buffer_13_620; // @[Modules.scala 53:83:@51558.4]
  wire [11:0] _T_97766; // @[Modules.scala 53:83:@51560.4]
  wire [10:0] _T_97767; // @[Modules.scala 53:83:@51561.4]
  wire [10:0] buffer_13_621; // @[Modules.scala 53:83:@51562.4]
  wire [11:0] _T_97769; // @[Modules.scala 53:83:@51564.4]
  wire [10:0] _T_97770; // @[Modules.scala 53:83:@51565.4]
  wire [10:0] buffer_13_622; // @[Modules.scala 53:83:@51566.4]
  wire [11:0] _T_97772; // @[Modules.scala 53:83:@51568.4]
  wire [10:0] _T_97773; // @[Modules.scala 53:83:@51569.4]
  wire [10:0] buffer_13_623; // @[Modules.scala 53:83:@51570.4]
  wire [11:0] _T_97775; // @[Modules.scala 53:83:@51572.4]
  wire [10:0] _T_97776; // @[Modules.scala 53:83:@51573.4]
  wire [10:0] buffer_13_624; // @[Modules.scala 53:83:@51574.4]
  wire [11:0] _T_97778; // @[Modules.scala 53:83:@51576.4]
  wire [10:0] _T_97779; // @[Modules.scala 53:83:@51577.4]
  wire [10:0] buffer_13_625; // @[Modules.scala 53:83:@51578.4]
  wire [11:0] _T_97784; // @[Modules.scala 53:83:@51584.4]
  wire [10:0] _T_97785; // @[Modules.scala 53:83:@51585.4]
  wire [10:0] buffer_13_627; // @[Modules.scala 53:83:@51586.4]
  wire [11:0] _T_97787; // @[Modules.scala 53:83:@51588.4]
  wire [10:0] _T_97788; // @[Modules.scala 53:83:@51589.4]
  wire [10:0] buffer_13_628; // @[Modules.scala 53:83:@51590.4]
  wire [11:0] _T_97790; // @[Modules.scala 53:83:@51592.4]
  wire [10:0] _T_97791; // @[Modules.scala 53:83:@51593.4]
  wire [10:0] buffer_13_629; // @[Modules.scala 53:83:@51594.4]
  wire [11:0] _T_97793; // @[Modules.scala 53:83:@51596.4]
  wire [10:0] _T_97794; // @[Modules.scala 53:83:@51597.4]
  wire [10:0] buffer_13_630; // @[Modules.scala 53:83:@51598.4]
  wire [11:0] _T_97796; // @[Modules.scala 53:83:@51600.4]
  wire [10:0] _T_97797; // @[Modules.scala 53:83:@51601.4]
  wire [10:0] buffer_13_631; // @[Modules.scala 53:83:@51602.4]
  wire [11:0] _T_97799; // @[Modules.scala 53:83:@51604.4]
  wire [10:0] _T_97800; // @[Modules.scala 53:83:@51605.4]
  wire [10:0] buffer_13_632; // @[Modules.scala 53:83:@51606.4]
  wire [11:0] _T_97802; // @[Modules.scala 53:83:@51608.4]
  wire [10:0] _T_97803; // @[Modules.scala 53:83:@51609.4]
  wire [10:0] buffer_13_633; // @[Modules.scala 53:83:@51610.4]
  wire [11:0] _T_97805; // @[Modules.scala 53:83:@51612.4]
  wire [10:0] _T_97806; // @[Modules.scala 53:83:@51613.4]
  wire [10:0] buffer_13_634; // @[Modules.scala 53:83:@51614.4]
  wire [11:0] _T_97808; // @[Modules.scala 53:83:@51616.4]
  wire [10:0] _T_97809; // @[Modules.scala 53:83:@51617.4]
  wire [10:0] buffer_13_635; // @[Modules.scala 53:83:@51618.4]
  wire [11:0] _T_97811; // @[Modules.scala 53:83:@51620.4]
  wire [10:0] _T_97812; // @[Modules.scala 53:83:@51621.4]
  wire [10:0] buffer_13_636; // @[Modules.scala 53:83:@51622.4]
  wire [11:0] _T_97814; // @[Modules.scala 53:83:@51624.4]
  wire [10:0] _T_97815; // @[Modules.scala 53:83:@51625.4]
  wire [10:0] buffer_13_637; // @[Modules.scala 53:83:@51626.4]
  wire [11:0] _T_97817; // @[Modules.scala 53:83:@51628.4]
  wire [10:0] _T_97818; // @[Modules.scala 53:83:@51629.4]
  wire [10:0] buffer_13_638; // @[Modules.scala 53:83:@51630.4]
  wire [11:0] _T_97820; // @[Modules.scala 53:83:@51632.4]
  wire [10:0] _T_97821; // @[Modules.scala 53:83:@51633.4]
  wire [10:0] buffer_13_639; // @[Modules.scala 53:83:@51634.4]
  wire [11:0] _T_97823; // @[Modules.scala 53:83:@51636.4]
  wire [10:0] _T_97824; // @[Modules.scala 53:83:@51637.4]
  wire [10:0] buffer_13_640; // @[Modules.scala 53:83:@51638.4]
  wire [11:0] _T_97826; // @[Modules.scala 53:83:@51640.4]
  wire [10:0] _T_97827; // @[Modules.scala 53:83:@51641.4]
  wire [10:0] buffer_13_641; // @[Modules.scala 53:83:@51642.4]
  wire [11:0] _T_97829; // @[Modules.scala 53:83:@51644.4]
  wire [10:0] _T_97830; // @[Modules.scala 53:83:@51645.4]
  wire [10:0] buffer_13_642; // @[Modules.scala 53:83:@51646.4]
  wire [11:0] _T_97832; // @[Modules.scala 53:83:@51648.4]
  wire [10:0] _T_97833; // @[Modules.scala 53:83:@51649.4]
  wire [10:0] buffer_13_643; // @[Modules.scala 53:83:@51650.4]
  wire [11:0] _T_97835; // @[Modules.scala 53:83:@51652.4]
  wire [10:0] _T_97836; // @[Modules.scala 53:83:@51653.4]
  wire [10:0] buffer_13_644; // @[Modules.scala 53:83:@51654.4]
  wire [11:0] _T_97838; // @[Modules.scala 53:83:@51656.4]
  wire [10:0] _T_97839; // @[Modules.scala 53:83:@51657.4]
  wire [10:0] buffer_13_645; // @[Modules.scala 53:83:@51658.4]
  wire [11:0] _T_97841; // @[Modules.scala 53:83:@51660.4]
  wire [10:0] _T_97842; // @[Modules.scala 53:83:@51661.4]
  wire [10:0] buffer_13_646; // @[Modules.scala 53:83:@51662.4]
  wire [11:0] _T_97847; // @[Modules.scala 53:83:@51668.4]
  wire [10:0] _T_97848; // @[Modules.scala 53:83:@51669.4]
  wire [10:0] buffer_13_648; // @[Modules.scala 53:83:@51670.4]
  wire [11:0] _T_97850; // @[Modules.scala 53:83:@51672.4]
  wire [10:0] _T_97851; // @[Modules.scala 53:83:@51673.4]
  wire [10:0] buffer_13_649; // @[Modules.scala 53:83:@51674.4]
  wire [11:0] _T_97853; // @[Modules.scala 53:83:@51676.4]
  wire [10:0] _T_97854; // @[Modules.scala 53:83:@51677.4]
  wire [10:0] buffer_13_650; // @[Modules.scala 53:83:@51678.4]
  wire [11:0] _T_97862; // @[Modules.scala 53:83:@51688.4]
  wire [10:0] _T_97863; // @[Modules.scala 53:83:@51689.4]
  wire [10:0] buffer_13_653; // @[Modules.scala 53:83:@51690.4]
  wire [11:0] _T_97865; // @[Modules.scala 53:83:@51692.4]
  wire [10:0] _T_97866; // @[Modules.scala 53:83:@51693.4]
  wire [10:0] buffer_13_654; // @[Modules.scala 53:83:@51694.4]
  wire [11:0] _T_97868; // @[Modules.scala 53:83:@51696.4]
  wire [10:0] _T_97869; // @[Modules.scala 53:83:@51697.4]
  wire [10:0] buffer_13_655; // @[Modules.scala 53:83:@51698.4]
  wire [11:0] _T_97871; // @[Modules.scala 53:83:@51700.4]
  wire [10:0] _T_97872; // @[Modules.scala 53:83:@51701.4]
  wire [10:0] buffer_13_656; // @[Modules.scala 53:83:@51702.4]
  wire [11:0] _T_97877; // @[Modules.scala 53:83:@51708.4]
  wire [10:0] _T_97878; // @[Modules.scala 53:83:@51709.4]
  wire [10:0] buffer_13_658; // @[Modules.scala 53:83:@51710.4]
  wire [11:0] _T_97883; // @[Modules.scala 53:83:@51716.4]
  wire [10:0] _T_97884; // @[Modules.scala 53:83:@51717.4]
  wire [10:0] buffer_13_660; // @[Modules.scala 53:83:@51718.4]
  wire [11:0] _T_97886; // @[Modules.scala 53:83:@51720.4]
  wire [10:0] _T_97887; // @[Modules.scala 53:83:@51721.4]
  wire [10:0] buffer_13_661; // @[Modules.scala 53:83:@51722.4]
  wire [11:0] _T_97889; // @[Modules.scala 53:83:@51724.4]
  wire [10:0] _T_97890; // @[Modules.scala 53:83:@51725.4]
  wire [10:0] buffer_13_662; // @[Modules.scala 53:83:@51726.4]
  wire [11:0] _T_97898; // @[Modules.scala 53:83:@51736.4]
  wire [10:0] _T_97899; // @[Modules.scala 53:83:@51737.4]
  wire [10:0] buffer_13_665; // @[Modules.scala 53:83:@51738.4]
  wire [11:0] _T_97901; // @[Modules.scala 53:83:@51740.4]
  wire [10:0] _T_97902; // @[Modules.scala 53:83:@51741.4]
  wire [10:0] buffer_13_666; // @[Modules.scala 53:83:@51742.4]
  wire [11:0] _T_97904; // @[Modules.scala 53:83:@51744.4]
  wire [10:0] _T_97905; // @[Modules.scala 53:83:@51745.4]
  wire [10:0] buffer_13_667; // @[Modules.scala 53:83:@51746.4]
  wire [11:0] _T_97907; // @[Modules.scala 53:83:@51748.4]
  wire [10:0] _T_97908; // @[Modules.scala 53:83:@51749.4]
  wire [10:0] buffer_13_668; // @[Modules.scala 53:83:@51750.4]
  wire [11:0] _T_97913; // @[Modules.scala 53:83:@51756.4]
  wire [10:0] _T_97914; // @[Modules.scala 53:83:@51757.4]
  wire [10:0] buffer_13_670; // @[Modules.scala 53:83:@51758.4]
  wire [11:0] _T_97919; // @[Modules.scala 53:83:@51764.4]
  wire [10:0] _T_97920; // @[Modules.scala 53:83:@51765.4]
  wire [10:0] buffer_13_672; // @[Modules.scala 53:83:@51766.4]
  wire [11:0] _T_97922; // @[Modules.scala 53:83:@51768.4]
  wire [10:0] _T_97923; // @[Modules.scala 53:83:@51769.4]
  wire [10:0] buffer_13_673; // @[Modules.scala 53:83:@51770.4]
  wire [11:0] _T_97928; // @[Modules.scala 53:83:@51776.4]
  wire [10:0] _T_97929; // @[Modules.scala 53:83:@51777.4]
  wire [10:0] buffer_13_675; // @[Modules.scala 53:83:@51778.4]
  wire [11:0] _T_97937; // @[Modules.scala 53:83:@51788.4]
  wire [10:0] _T_97938; // @[Modules.scala 53:83:@51789.4]
  wire [10:0] buffer_13_678; // @[Modules.scala 53:83:@51790.4]
  wire [11:0] _T_97940; // @[Modules.scala 53:83:@51792.4]
  wire [10:0] _T_97941; // @[Modules.scala 53:83:@51793.4]
  wire [10:0] buffer_13_679; // @[Modules.scala 53:83:@51794.4]
  wire [11:0] _T_97949; // @[Modules.scala 53:83:@51804.4]
  wire [10:0] _T_97950; // @[Modules.scala 53:83:@51805.4]
  wire [10:0] buffer_13_682; // @[Modules.scala 53:83:@51806.4]
  wire [11:0] _T_97958; // @[Modules.scala 53:83:@51816.4]
  wire [10:0] _T_97959; // @[Modules.scala 53:83:@51817.4]
  wire [10:0] buffer_13_685; // @[Modules.scala 53:83:@51818.4]
  wire [11:0] _T_97961; // @[Modules.scala 56:109:@51820.4]
  wire [10:0] _T_97962; // @[Modules.scala 56:109:@51821.4]
  wire [10:0] buffer_13_686; // @[Modules.scala 56:109:@51822.4]
  wire [11:0] _T_97964; // @[Modules.scala 56:109:@51824.4]
  wire [10:0] _T_97965; // @[Modules.scala 56:109:@51825.4]
  wire [10:0] buffer_13_687; // @[Modules.scala 56:109:@51826.4]
  wire [11:0] _T_97967; // @[Modules.scala 56:109:@51828.4]
  wire [10:0] _T_97968; // @[Modules.scala 56:109:@51829.4]
  wire [10:0] buffer_13_688; // @[Modules.scala 56:109:@51830.4]
  wire [11:0] _T_97970; // @[Modules.scala 56:109:@51832.4]
  wire [10:0] _T_97971; // @[Modules.scala 56:109:@51833.4]
  wire [10:0] buffer_13_689; // @[Modules.scala 56:109:@51834.4]
  wire [11:0] _T_97973; // @[Modules.scala 56:109:@51836.4]
  wire [10:0] _T_97974; // @[Modules.scala 56:109:@51837.4]
  wire [10:0] buffer_13_690; // @[Modules.scala 56:109:@51838.4]
  wire [11:0] _T_97976; // @[Modules.scala 56:109:@51840.4]
  wire [10:0] _T_97977; // @[Modules.scala 56:109:@51841.4]
  wire [10:0] buffer_13_691; // @[Modules.scala 56:109:@51842.4]
  wire [11:0] _T_97979; // @[Modules.scala 56:109:@51844.4]
  wire [10:0] _T_97980; // @[Modules.scala 56:109:@51845.4]
  wire [10:0] buffer_13_692; // @[Modules.scala 56:109:@51846.4]
  wire [11:0] _T_97982; // @[Modules.scala 56:109:@51848.4]
  wire [10:0] _T_97983; // @[Modules.scala 56:109:@51849.4]
  wire [10:0] buffer_13_693; // @[Modules.scala 56:109:@51850.4]
  wire [11:0] _T_97985; // @[Modules.scala 56:109:@51852.4]
  wire [10:0] _T_97986; // @[Modules.scala 56:109:@51853.4]
  wire [10:0] buffer_13_694; // @[Modules.scala 56:109:@51854.4]
  wire [11:0] _T_97988; // @[Modules.scala 56:109:@51856.4]
  wire [10:0] _T_97989; // @[Modules.scala 56:109:@51857.4]
  wire [10:0] buffer_13_695; // @[Modules.scala 56:109:@51858.4]
  wire [11:0] _T_97991; // @[Modules.scala 56:109:@51860.4]
  wire [10:0] _T_97992; // @[Modules.scala 56:109:@51861.4]
  wire [10:0] buffer_13_696; // @[Modules.scala 56:109:@51862.4]
  wire [11:0] _T_97994; // @[Modules.scala 56:109:@51864.4]
  wire [10:0] _T_97995; // @[Modules.scala 56:109:@51865.4]
  wire [10:0] buffer_13_697; // @[Modules.scala 56:109:@51866.4]
  wire [11:0] _T_97997; // @[Modules.scala 56:109:@51868.4]
  wire [10:0] _T_97998; // @[Modules.scala 56:109:@51869.4]
  wire [10:0] buffer_13_698; // @[Modules.scala 56:109:@51870.4]
  wire [11:0] _T_98000; // @[Modules.scala 56:109:@51872.4]
  wire [10:0] _T_98001; // @[Modules.scala 56:109:@51873.4]
  wire [10:0] buffer_13_699; // @[Modules.scala 56:109:@51874.4]
  wire [11:0] _T_98003; // @[Modules.scala 56:109:@51876.4]
  wire [10:0] _T_98004; // @[Modules.scala 56:109:@51877.4]
  wire [10:0] buffer_13_700; // @[Modules.scala 56:109:@51878.4]
  wire [11:0] _T_98006; // @[Modules.scala 56:109:@51880.4]
  wire [10:0] _T_98007; // @[Modules.scala 56:109:@51881.4]
  wire [10:0] buffer_13_701; // @[Modules.scala 56:109:@51882.4]
  wire [11:0] _T_98009; // @[Modules.scala 56:109:@51884.4]
  wire [10:0] _T_98010; // @[Modules.scala 56:109:@51885.4]
  wire [10:0] buffer_13_702; // @[Modules.scala 56:109:@51886.4]
  wire [11:0] _T_98012; // @[Modules.scala 56:109:@51888.4]
  wire [10:0] _T_98013; // @[Modules.scala 56:109:@51889.4]
  wire [10:0] buffer_13_703; // @[Modules.scala 56:109:@51890.4]
  wire [11:0] _T_98015; // @[Modules.scala 56:109:@51892.4]
  wire [10:0] _T_98016; // @[Modules.scala 56:109:@51893.4]
  wire [10:0] buffer_13_704; // @[Modules.scala 56:109:@51894.4]
  wire [11:0] _T_98018; // @[Modules.scala 56:109:@51896.4]
  wire [10:0] _T_98019; // @[Modules.scala 56:109:@51897.4]
  wire [10:0] buffer_13_705; // @[Modules.scala 56:109:@51898.4]
  wire [11:0] _T_98021; // @[Modules.scala 56:109:@51900.4]
  wire [10:0] _T_98022; // @[Modules.scala 56:109:@51901.4]
  wire [10:0] buffer_13_706; // @[Modules.scala 56:109:@51902.4]
  wire [11:0] _T_98024; // @[Modules.scala 56:109:@51904.4]
  wire [10:0] _T_98025; // @[Modules.scala 56:109:@51905.4]
  wire [10:0] buffer_13_707; // @[Modules.scala 56:109:@51906.4]
  wire [11:0] _T_98027; // @[Modules.scala 56:109:@51908.4]
  wire [10:0] _T_98028; // @[Modules.scala 56:109:@51909.4]
  wire [10:0] buffer_13_708; // @[Modules.scala 56:109:@51910.4]
  wire [11:0] _T_98030; // @[Modules.scala 56:109:@51912.4]
  wire [10:0] _T_98031; // @[Modules.scala 56:109:@51913.4]
  wire [10:0] buffer_13_709; // @[Modules.scala 56:109:@51914.4]
  wire [11:0] _T_98033; // @[Modules.scala 56:109:@51916.4]
  wire [10:0] _T_98034; // @[Modules.scala 56:109:@51917.4]
  wire [10:0] buffer_13_710; // @[Modules.scala 56:109:@51918.4]
  wire [11:0] _T_98036; // @[Modules.scala 56:109:@51920.4]
  wire [10:0] _T_98037; // @[Modules.scala 56:109:@51921.4]
  wire [10:0] buffer_13_711; // @[Modules.scala 56:109:@51922.4]
  wire [11:0] _T_98039; // @[Modules.scala 56:109:@51924.4]
  wire [10:0] _T_98040; // @[Modules.scala 56:109:@51925.4]
  wire [10:0] buffer_13_712; // @[Modules.scala 56:109:@51926.4]
  wire [11:0] _T_98042; // @[Modules.scala 56:109:@51928.4]
  wire [10:0] _T_98043; // @[Modules.scala 56:109:@51929.4]
  wire [10:0] buffer_13_713; // @[Modules.scala 56:109:@51930.4]
  wire [11:0] _T_98045; // @[Modules.scala 56:109:@51932.4]
  wire [10:0] _T_98046; // @[Modules.scala 56:109:@51933.4]
  wire [10:0] buffer_13_714; // @[Modules.scala 56:109:@51934.4]
  wire [11:0] _T_98048; // @[Modules.scala 56:109:@51936.4]
  wire [10:0] _T_98049; // @[Modules.scala 56:109:@51937.4]
  wire [10:0] buffer_13_715; // @[Modules.scala 56:109:@51938.4]
  wire [11:0] _T_98051; // @[Modules.scala 56:109:@51940.4]
  wire [10:0] _T_98052; // @[Modules.scala 56:109:@51941.4]
  wire [10:0] buffer_13_716; // @[Modules.scala 56:109:@51942.4]
  wire [11:0] _T_98054; // @[Modules.scala 56:109:@51944.4]
  wire [10:0] _T_98055; // @[Modules.scala 56:109:@51945.4]
  wire [10:0] buffer_13_717; // @[Modules.scala 56:109:@51946.4]
  wire [11:0] _T_98057; // @[Modules.scala 56:109:@51948.4]
  wire [10:0] _T_98058; // @[Modules.scala 56:109:@51949.4]
  wire [10:0] buffer_13_718; // @[Modules.scala 56:109:@51950.4]
  wire [11:0] _T_98060; // @[Modules.scala 56:109:@51952.4]
  wire [10:0] _T_98061; // @[Modules.scala 56:109:@51953.4]
  wire [10:0] buffer_13_719; // @[Modules.scala 56:109:@51954.4]
  wire [11:0] _T_98063; // @[Modules.scala 56:109:@51956.4]
  wire [10:0] _T_98064; // @[Modules.scala 56:109:@51957.4]
  wire [10:0] buffer_13_720; // @[Modules.scala 56:109:@51958.4]
  wire [11:0] _T_98066; // @[Modules.scala 56:109:@51960.4]
  wire [10:0] _T_98067; // @[Modules.scala 56:109:@51961.4]
  wire [10:0] buffer_13_721; // @[Modules.scala 56:109:@51962.4]
  wire [11:0] _T_98069; // @[Modules.scala 56:109:@51964.4]
  wire [10:0] _T_98070; // @[Modules.scala 56:109:@51965.4]
  wire [10:0] buffer_13_722; // @[Modules.scala 56:109:@51966.4]
  wire [11:0] _T_98072; // @[Modules.scala 56:109:@51968.4]
  wire [10:0] _T_98073; // @[Modules.scala 56:109:@51969.4]
  wire [10:0] buffer_13_723; // @[Modules.scala 56:109:@51970.4]
  wire [11:0] _T_98075; // @[Modules.scala 56:109:@51972.4]
  wire [10:0] _T_98076; // @[Modules.scala 56:109:@51973.4]
  wire [10:0] buffer_13_724; // @[Modules.scala 56:109:@51974.4]
  wire [11:0] _T_98078; // @[Modules.scala 56:109:@51976.4]
  wire [10:0] _T_98079; // @[Modules.scala 56:109:@51977.4]
  wire [10:0] buffer_13_725; // @[Modules.scala 56:109:@51978.4]
  wire [11:0] _T_98081; // @[Modules.scala 56:109:@51980.4]
  wire [10:0] _T_98082; // @[Modules.scala 56:109:@51981.4]
  wire [10:0] buffer_13_726; // @[Modules.scala 56:109:@51982.4]
  wire [11:0] _T_98084; // @[Modules.scala 56:109:@51984.4]
  wire [10:0] _T_98085; // @[Modules.scala 56:109:@51985.4]
  wire [10:0] buffer_13_727; // @[Modules.scala 56:109:@51986.4]
  wire [11:0] _T_98087; // @[Modules.scala 56:109:@51988.4]
  wire [10:0] _T_98088; // @[Modules.scala 56:109:@51989.4]
  wire [10:0] buffer_13_728; // @[Modules.scala 56:109:@51990.4]
  wire [11:0] _T_98090; // @[Modules.scala 56:109:@51992.4]
  wire [10:0] _T_98091; // @[Modules.scala 56:109:@51993.4]
  wire [10:0] buffer_13_729; // @[Modules.scala 56:109:@51994.4]
  wire [11:0] _T_98096; // @[Modules.scala 56:109:@52000.4]
  wire [10:0] _T_98097; // @[Modules.scala 56:109:@52001.4]
  wire [10:0] buffer_13_731; // @[Modules.scala 56:109:@52002.4]
  wire [11:0] _T_98102; // @[Modules.scala 56:109:@52008.4]
  wire [10:0] _T_98103; // @[Modules.scala 56:109:@52009.4]
  wire [10:0] buffer_13_733; // @[Modules.scala 56:109:@52010.4]
  wire [11:0] _T_98105; // @[Modules.scala 56:109:@52012.4]
  wire [10:0] _T_98106; // @[Modules.scala 56:109:@52013.4]
  wire [10:0] buffer_13_734; // @[Modules.scala 56:109:@52014.4]
  wire [11:0] _T_98108; // @[Modules.scala 63:156:@52017.4]
  wire [10:0] _T_98109; // @[Modules.scala 63:156:@52018.4]
  wire [10:0] buffer_13_736; // @[Modules.scala 63:156:@52019.4]
  wire [11:0] _T_98111; // @[Modules.scala 63:156:@52021.4]
  wire [10:0] _T_98112; // @[Modules.scala 63:156:@52022.4]
  wire [10:0] buffer_13_737; // @[Modules.scala 63:156:@52023.4]
  wire [11:0] _T_98114; // @[Modules.scala 63:156:@52025.4]
  wire [10:0] _T_98115; // @[Modules.scala 63:156:@52026.4]
  wire [10:0] buffer_13_738; // @[Modules.scala 63:156:@52027.4]
  wire [11:0] _T_98117; // @[Modules.scala 63:156:@52029.4]
  wire [10:0] _T_98118; // @[Modules.scala 63:156:@52030.4]
  wire [10:0] buffer_13_739; // @[Modules.scala 63:156:@52031.4]
  wire [11:0] _T_98120; // @[Modules.scala 63:156:@52033.4]
  wire [10:0] _T_98121; // @[Modules.scala 63:156:@52034.4]
  wire [10:0] buffer_13_740; // @[Modules.scala 63:156:@52035.4]
  wire [11:0] _T_98123; // @[Modules.scala 63:156:@52037.4]
  wire [10:0] _T_98124; // @[Modules.scala 63:156:@52038.4]
  wire [10:0] buffer_13_741; // @[Modules.scala 63:156:@52039.4]
  wire [11:0] _T_98126; // @[Modules.scala 63:156:@52041.4]
  wire [10:0] _T_98127; // @[Modules.scala 63:156:@52042.4]
  wire [10:0] buffer_13_742; // @[Modules.scala 63:156:@52043.4]
  wire [11:0] _T_98129; // @[Modules.scala 63:156:@52045.4]
  wire [10:0] _T_98130; // @[Modules.scala 63:156:@52046.4]
  wire [10:0] buffer_13_743; // @[Modules.scala 63:156:@52047.4]
  wire [11:0] _T_98132; // @[Modules.scala 63:156:@52049.4]
  wire [10:0] _T_98133; // @[Modules.scala 63:156:@52050.4]
  wire [10:0] buffer_13_744; // @[Modules.scala 63:156:@52051.4]
  wire [11:0] _T_98135; // @[Modules.scala 63:156:@52053.4]
  wire [10:0] _T_98136; // @[Modules.scala 63:156:@52054.4]
  wire [10:0] buffer_13_745; // @[Modules.scala 63:156:@52055.4]
  wire [11:0] _T_98138; // @[Modules.scala 63:156:@52057.4]
  wire [10:0] _T_98139; // @[Modules.scala 63:156:@52058.4]
  wire [10:0] buffer_13_746; // @[Modules.scala 63:156:@52059.4]
  wire [11:0] _T_98141; // @[Modules.scala 63:156:@52061.4]
  wire [10:0] _T_98142; // @[Modules.scala 63:156:@52062.4]
  wire [10:0] buffer_13_747; // @[Modules.scala 63:156:@52063.4]
  wire [11:0] _T_98144; // @[Modules.scala 63:156:@52065.4]
  wire [10:0] _T_98145; // @[Modules.scala 63:156:@52066.4]
  wire [10:0] buffer_13_748; // @[Modules.scala 63:156:@52067.4]
  wire [11:0] _T_98147; // @[Modules.scala 63:156:@52069.4]
  wire [10:0] _T_98148; // @[Modules.scala 63:156:@52070.4]
  wire [10:0] buffer_13_749; // @[Modules.scala 63:156:@52071.4]
  wire [11:0] _T_98150; // @[Modules.scala 63:156:@52073.4]
  wire [10:0] _T_98151; // @[Modules.scala 63:156:@52074.4]
  wire [10:0] buffer_13_750; // @[Modules.scala 63:156:@52075.4]
  wire [11:0] _T_98153; // @[Modules.scala 63:156:@52077.4]
  wire [10:0] _T_98154; // @[Modules.scala 63:156:@52078.4]
  wire [10:0] buffer_13_751; // @[Modules.scala 63:156:@52079.4]
  wire [11:0] _T_98156; // @[Modules.scala 63:156:@52081.4]
  wire [10:0] _T_98157; // @[Modules.scala 63:156:@52082.4]
  wire [10:0] buffer_13_752; // @[Modules.scala 63:156:@52083.4]
  wire [11:0] _T_98159; // @[Modules.scala 63:156:@52085.4]
  wire [10:0] _T_98160; // @[Modules.scala 63:156:@52086.4]
  wire [10:0] buffer_13_753; // @[Modules.scala 63:156:@52087.4]
  wire [11:0] _T_98162; // @[Modules.scala 63:156:@52089.4]
  wire [10:0] _T_98163; // @[Modules.scala 63:156:@52090.4]
  wire [10:0] buffer_13_754; // @[Modules.scala 63:156:@52091.4]
  wire [11:0] _T_98165; // @[Modules.scala 63:156:@52093.4]
  wire [10:0] _T_98166; // @[Modules.scala 63:156:@52094.4]
  wire [10:0] buffer_13_755; // @[Modules.scala 63:156:@52095.4]
  wire [11:0] _T_98168; // @[Modules.scala 63:156:@52097.4]
  wire [10:0] _T_98169; // @[Modules.scala 63:156:@52098.4]
  wire [10:0] buffer_13_756; // @[Modules.scala 63:156:@52099.4]
  wire [11:0] _T_98171; // @[Modules.scala 63:156:@52101.4]
  wire [10:0] _T_98172; // @[Modules.scala 63:156:@52102.4]
  wire [10:0] buffer_13_757; // @[Modules.scala 63:156:@52103.4]
  wire [11:0] _T_98174; // @[Modules.scala 63:156:@52105.4]
  wire [10:0] _T_98175; // @[Modules.scala 63:156:@52106.4]
  wire [10:0] buffer_13_758; // @[Modules.scala 63:156:@52107.4]
  wire [11:0] _T_98177; // @[Modules.scala 63:156:@52109.4]
  wire [10:0] _T_98178; // @[Modules.scala 63:156:@52110.4]
  wire [10:0] buffer_13_759; // @[Modules.scala 63:156:@52111.4]
  wire [11:0] _T_98180; // @[Modules.scala 63:156:@52113.4]
  wire [10:0] _T_98181; // @[Modules.scala 63:156:@52114.4]
  wire [10:0] buffer_13_760; // @[Modules.scala 63:156:@52115.4]
  wire [11:0] _T_98183; // @[Modules.scala 63:156:@52117.4]
  wire [10:0] _T_98184; // @[Modules.scala 63:156:@52118.4]
  wire [10:0] buffer_13_761; // @[Modules.scala 63:156:@52119.4]
  wire [11:0] _T_98186; // @[Modules.scala 63:156:@52121.4]
  wire [10:0] _T_98187; // @[Modules.scala 63:156:@52122.4]
  wire [10:0] buffer_13_762; // @[Modules.scala 63:156:@52123.4]
  wire [11:0] _T_98189; // @[Modules.scala 63:156:@52125.4]
  wire [10:0] _T_98190; // @[Modules.scala 63:156:@52126.4]
  wire [10:0] buffer_13_763; // @[Modules.scala 63:156:@52127.4]
  wire [11:0] _T_98192; // @[Modules.scala 63:156:@52129.4]
  wire [10:0] _T_98193; // @[Modules.scala 63:156:@52130.4]
  wire [10:0] buffer_13_764; // @[Modules.scala 63:156:@52131.4]
  wire [11:0] _T_98195; // @[Modules.scala 63:156:@52133.4]
  wire [10:0] _T_98196; // @[Modules.scala 63:156:@52134.4]
  wire [10:0] buffer_13_765; // @[Modules.scala 63:156:@52135.4]
  wire [11:0] _T_98198; // @[Modules.scala 63:156:@52137.4]
  wire [10:0] _T_98199; // @[Modules.scala 63:156:@52138.4]
  wire [10:0] buffer_13_766; // @[Modules.scala 63:156:@52139.4]
  wire [11:0] _T_98201; // @[Modules.scala 63:156:@52141.4]
  wire [10:0] _T_98202; // @[Modules.scala 63:156:@52142.4]
  wire [10:0] buffer_13_767; // @[Modules.scala 63:156:@52143.4]
  wire [11:0] _T_98204; // @[Modules.scala 63:156:@52145.4]
  wire [10:0] _T_98205; // @[Modules.scala 63:156:@52146.4]
  wire [10:0] buffer_13_768; // @[Modules.scala 63:156:@52147.4]
  wire [11:0] _T_98207; // @[Modules.scala 63:156:@52149.4]
  wire [10:0] _T_98208; // @[Modules.scala 63:156:@52150.4]
  wire [10:0] buffer_13_769; // @[Modules.scala 63:156:@52151.4]
  wire [11:0] _T_98210; // @[Modules.scala 63:156:@52153.4]
  wire [10:0] _T_98211; // @[Modules.scala 63:156:@52154.4]
  wire [10:0] buffer_13_770; // @[Modules.scala 63:156:@52155.4]
  wire [11:0] _T_98213; // @[Modules.scala 63:156:@52157.4]
  wire [10:0] _T_98214; // @[Modules.scala 63:156:@52158.4]
  wire [10:0] buffer_13_771; // @[Modules.scala 63:156:@52159.4]
  wire [11:0] _T_98216; // @[Modules.scala 63:156:@52161.4]
  wire [10:0] _T_98217; // @[Modules.scala 63:156:@52162.4]
  wire [10:0] buffer_13_772; // @[Modules.scala 63:156:@52163.4]
  wire [11:0] _T_98219; // @[Modules.scala 63:156:@52165.4]
  wire [10:0] _T_98220; // @[Modules.scala 63:156:@52166.4]
  wire [10:0] buffer_13_773; // @[Modules.scala 63:156:@52167.4]
  wire [11:0] _T_98222; // @[Modules.scala 63:156:@52169.4]
  wire [10:0] _T_98223; // @[Modules.scala 63:156:@52170.4]
  wire [10:0] buffer_13_774; // @[Modules.scala 63:156:@52171.4]
  wire [11:0] _T_98225; // @[Modules.scala 63:156:@52173.4]
  wire [10:0] _T_98226; // @[Modules.scala 63:156:@52174.4]
  wire [10:0] buffer_13_775; // @[Modules.scala 63:156:@52175.4]
  wire [11:0] _T_98228; // @[Modules.scala 63:156:@52177.4]
  wire [10:0] _T_98229; // @[Modules.scala 63:156:@52178.4]
  wire [10:0] buffer_13_776; // @[Modules.scala 63:156:@52179.4]
  wire [11:0] _T_98231; // @[Modules.scala 63:156:@52181.4]
  wire [10:0] _T_98232; // @[Modules.scala 63:156:@52182.4]
  wire [10:0] buffer_13_777; // @[Modules.scala 63:156:@52183.4]
  wire [11:0] _T_98234; // @[Modules.scala 63:156:@52185.4]
  wire [10:0] _T_98235; // @[Modules.scala 63:156:@52186.4]
  wire [10:0] buffer_13_778; // @[Modules.scala 63:156:@52187.4]
  wire [11:0] _T_98237; // @[Modules.scala 63:156:@52189.4]
  wire [10:0] _T_98238; // @[Modules.scala 63:156:@52190.4]
  wire [10:0] buffer_13_779; // @[Modules.scala 63:156:@52191.4]
  wire [11:0] _T_98240; // @[Modules.scala 63:156:@52193.4]
  wire [10:0] _T_98241; // @[Modules.scala 63:156:@52194.4]
  wire [10:0] buffer_13_780; // @[Modules.scala 63:156:@52195.4]
  wire [11:0] _T_98243; // @[Modules.scala 63:156:@52197.4]
  wire [10:0] _T_98244; // @[Modules.scala 63:156:@52198.4]
  wire [10:0] buffer_13_781; // @[Modules.scala 63:156:@52199.4]
  wire [11:0] _T_98246; // @[Modules.scala 63:156:@52201.4]
  wire [10:0] _T_98247; // @[Modules.scala 63:156:@52202.4]
  wire [10:0] buffer_13_782; // @[Modules.scala 63:156:@52203.4]
  wire [11:0] _T_98249; // @[Modules.scala 63:156:@52205.4]
  wire [10:0] _T_98250; // @[Modules.scala 63:156:@52206.4]
  wire [10:0] buffer_13_783; // @[Modules.scala 63:156:@52207.4]
  wire [5:0] _T_98414; // @[Modules.scala 40:46:@52384.4]
  wire [4:0] _T_98415; // @[Modules.scala 40:46:@52385.4]
  wire [4:0] _T_98416; // @[Modules.scala 40:46:@52386.4]
  wire [5:0] _T_98499; // @[Modules.scala 43:47:@52474.4]
  wire [4:0] _T_98500; // @[Modules.scala 43:47:@52475.4]
  wire [4:0] _T_98501; // @[Modules.scala 43:47:@52476.4]
  wire [5:0] _T_98508; // @[Modules.scala 40:46:@52486.4]
  wire [4:0] _T_98509; // @[Modules.scala 40:46:@52487.4]
  wire [4:0] _T_98510; // @[Modules.scala 40:46:@52488.4]
  wire [5:0] _T_98630; // @[Modules.scala 46:47:@52616.4]
  wire [4:0] _T_98631; // @[Modules.scala 46:47:@52617.4]
  wire [4:0] _T_98632; // @[Modules.scala 46:47:@52618.4]
  wire [5:0] _T_98712; // @[Modules.scala 43:47:@52709.4]
  wire [4:0] _T_98713; // @[Modules.scala 43:47:@52710.4]
  wire [4:0] _T_98714; // @[Modules.scala 43:47:@52711.4]
  wire [5:0] _T_98934; // @[Modules.scala 43:47:@52956.4]
  wire [4:0] _T_98935; // @[Modules.scala 43:47:@52957.4]
  wire [4:0] _T_98936; // @[Modules.scala 43:47:@52958.4]
  wire [5:0] _T_99080; // @[Modules.scala 40:46:@53118.4]
  wire [4:0] _T_99081; // @[Modules.scala 40:46:@53119.4]
  wire [4:0] _T_99082; // @[Modules.scala 40:46:@53120.4]
  wire [5:0] _T_99127; // @[Modules.scala 40:46:@53169.4]
  wire [4:0] _T_99128; // @[Modules.scala 40:46:@53170.4]
  wire [4:0] _T_99129; // @[Modules.scala 40:46:@53171.4]
  wire [5:0] _T_99156; // @[Modules.scala 40:46:@53203.4]
  wire [4:0] _T_99157; // @[Modules.scala 40:46:@53204.4]
  wire [4:0] _T_99158; // @[Modules.scala 40:46:@53205.4]
  wire [5:0] _T_99349; // @[Modules.scala 40:46:@53409.4]
  wire [4:0] _T_99350; // @[Modules.scala 40:46:@53410.4]
  wire [4:0] _T_99351; // @[Modules.scala 40:46:@53411.4]
  wire [5:0] _T_99356; // @[Modules.scala 43:47:@53416.4]
  wire [4:0] _T_99357; // @[Modules.scala 43:47:@53417.4]
  wire [4:0] _T_99358; // @[Modules.scala 43:47:@53418.4]
  wire [5:0] _T_99640; // @[Modules.scala 40:46:@53748.4]
  wire [4:0] _T_99641; // @[Modules.scala 40:46:@53749.4]
  wire [4:0] _T_99642; // @[Modules.scala 40:46:@53750.4]
  wire [5:0] _T_99942; // @[Modules.scala 43:47:@54097.4]
  wire [4:0] _T_99943; // @[Modules.scala 43:47:@54098.4]
  wire [4:0] _T_99944; // @[Modules.scala 43:47:@54099.4]
  wire [5:0] _T_99973; // @[Modules.scala 43:47:@54136.4]
  wire [4:0] _T_99974; // @[Modules.scala 43:47:@54137.4]
  wire [4:0] _T_99975; // @[Modules.scala 43:47:@54138.4]
  wire [5:0] _T_99997; // @[Modules.scala 43:47:@54161.4]
  wire [4:0] _T_99998; // @[Modules.scala 43:47:@54162.4]
  wire [4:0] _T_99999; // @[Modules.scala 43:47:@54163.4]
  wire [5:0] _T_100000; // @[Modules.scala 40:46:@54165.4]
  wire [4:0] _T_100001; // @[Modules.scala 40:46:@54166.4]
  wire [4:0] _T_100002; // @[Modules.scala 40:46:@54167.4]
  wire [5:0] _T_100003; // @[Modules.scala 40:46:@54169.4]
  wire [4:0] _T_100004; // @[Modules.scala 40:46:@54170.4]
  wire [4:0] _T_100005; // @[Modules.scala 40:46:@54171.4]
  wire [11:0] _T_100116; // @[Modules.scala 50:57:@54294.4]
  wire [10:0] _T_100117; // @[Modules.scala 50:57:@54295.4]
  wire [10:0] buffer_14_392; // @[Modules.scala 50:57:@54296.4]
  wire [11:0] _T_100122; // @[Modules.scala 50:57:@54302.4]
  wire [10:0] _T_100123; // @[Modules.scala 50:57:@54303.4]
  wire [10:0] buffer_14_394; // @[Modules.scala 50:57:@54304.4]
  wire [11:0] _T_100137; // @[Modules.scala 50:57:@54322.4]
  wire [10:0] _T_100138; // @[Modules.scala 50:57:@54323.4]
  wire [10:0] buffer_14_399; // @[Modules.scala 50:57:@54324.4]
  wire [11:0] _T_100146; // @[Modules.scala 50:57:@54334.4]
  wire [10:0] _T_100147; // @[Modules.scala 50:57:@54335.4]
  wire [10:0] buffer_14_402; // @[Modules.scala 50:57:@54336.4]
  wire [11:0] _T_100155; // @[Modules.scala 50:57:@54346.4]
  wire [10:0] _T_100156; // @[Modules.scala 50:57:@54347.4]
  wire [10:0] buffer_14_405; // @[Modules.scala 50:57:@54348.4]
  wire [10:0] buffer_14_30; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100161; // @[Modules.scala 50:57:@54354.4]
  wire [10:0] _T_100162; // @[Modules.scala 50:57:@54355.4]
  wire [10:0] buffer_14_407; // @[Modules.scala 50:57:@54356.4]
  wire [11:0] _T_100179; // @[Modules.scala 50:57:@54378.4]
  wire [10:0] _T_100180; // @[Modules.scala 50:57:@54379.4]
  wire [10:0] buffer_14_413; // @[Modules.scala 50:57:@54380.4]
  wire [10:0] buffer_14_45; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100182; // @[Modules.scala 50:57:@54382.4]
  wire [10:0] _T_100183; // @[Modules.scala 50:57:@54383.4]
  wire [10:0] buffer_14_414; // @[Modules.scala 50:57:@54384.4]
  wire [10:0] buffer_14_48; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100188; // @[Modules.scala 50:57:@54390.4]
  wire [10:0] _T_100189; // @[Modules.scala 50:57:@54391.4]
  wire [10:0] buffer_14_416; // @[Modules.scala 50:57:@54392.4]
  wire [11:0] _T_100200; // @[Modules.scala 50:57:@54406.4]
  wire [10:0] _T_100201; // @[Modules.scala 50:57:@54407.4]
  wire [10:0] buffer_14_420; // @[Modules.scala 50:57:@54408.4]
  wire [11:0] _T_100209; // @[Modules.scala 50:57:@54418.4]
  wire [10:0] _T_100210; // @[Modules.scala 50:57:@54419.4]
  wire [10:0] buffer_14_423; // @[Modules.scala 50:57:@54420.4]
  wire [10:0] buffer_14_70; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100221; // @[Modules.scala 50:57:@54434.4]
  wire [10:0] _T_100222; // @[Modules.scala 50:57:@54435.4]
  wire [10:0] buffer_14_427; // @[Modules.scala 50:57:@54436.4]
  wire [10:0] buffer_14_88; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100248; // @[Modules.scala 50:57:@54470.4]
  wire [10:0] _T_100249; // @[Modules.scala 50:57:@54471.4]
  wire [10:0] buffer_14_436; // @[Modules.scala 50:57:@54472.4]
  wire [11:0] _T_100254; // @[Modules.scala 50:57:@54478.4]
  wire [10:0] _T_100255; // @[Modules.scala 50:57:@54479.4]
  wire [10:0] buffer_14_438; // @[Modules.scala 50:57:@54480.4]
  wire [11:0] _T_100257; // @[Modules.scala 50:57:@54482.4]
  wire [10:0] _T_100258; // @[Modules.scala 50:57:@54483.4]
  wire [10:0] buffer_14_439; // @[Modules.scala 50:57:@54484.4]
  wire [11:0] _T_100296; // @[Modules.scala 50:57:@54534.4]
  wire [10:0] _T_100297; // @[Modules.scala 50:57:@54535.4]
  wire [10:0] buffer_14_452; // @[Modules.scala 50:57:@54536.4]
  wire [10:0] buffer_14_134; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100317; // @[Modules.scala 50:57:@54562.4]
  wire [10:0] _T_100318; // @[Modules.scala 50:57:@54563.4]
  wire [10:0] buffer_14_459; // @[Modules.scala 50:57:@54564.4]
  wire [11:0] _T_100320; // @[Modules.scala 50:57:@54566.4]
  wire [10:0] _T_100321; // @[Modules.scala 50:57:@54567.4]
  wire [10:0] buffer_14_460; // @[Modules.scala 50:57:@54568.4]
  wire [11:0] _T_100323; // @[Modules.scala 50:57:@54570.4]
  wire [10:0] _T_100324; // @[Modules.scala 50:57:@54571.4]
  wire [10:0] buffer_14_461; // @[Modules.scala 50:57:@54572.4]
  wire [10:0] buffer_14_164; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100362; // @[Modules.scala 50:57:@54622.4]
  wire [10:0] _T_100363; // @[Modules.scala 50:57:@54623.4]
  wire [10:0] buffer_14_474; // @[Modules.scala 50:57:@54624.4]
  wire [11:0] _T_100371; // @[Modules.scala 50:57:@54634.4]
  wire [10:0] _T_100372; // @[Modules.scala 50:57:@54635.4]
  wire [10:0] buffer_14_477; // @[Modules.scala 50:57:@54636.4]
  wire [10:0] buffer_14_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100374; // @[Modules.scala 50:57:@54638.4]
  wire [10:0] _T_100375; // @[Modules.scala 50:57:@54639.4]
  wire [10:0] buffer_14_478; // @[Modules.scala 50:57:@54640.4]
  wire [10:0] buffer_14_180; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100386; // @[Modules.scala 50:57:@54654.4]
  wire [10:0] _T_100387; // @[Modules.scala 50:57:@54655.4]
  wire [10:0] buffer_14_482; // @[Modules.scala 50:57:@54656.4]
  wire [11:0] _T_100392; // @[Modules.scala 50:57:@54662.4]
  wire [10:0] _T_100393; // @[Modules.scala 50:57:@54663.4]
  wire [10:0] buffer_14_484; // @[Modules.scala 50:57:@54664.4]
  wire [11:0] _T_100395; // @[Modules.scala 50:57:@54666.4]
  wire [10:0] _T_100396; // @[Modules.scala 50:57:@54667.4]
  wire [10:0] buffer_14_485; // @[Modules.scala 50:57:@54668.4]
  wire [11:0] _T_100404; // @[Modules.scala 50:57:@54678.4]
  wire [10:0] _T_100405; // @[Modules.scala 50:57:@54679.4]
  wire [10:0] buffer_14_488; // @[Modules.scala 50:57:@54680.4]
  wire [11:0] _T_100428; // @[Modules.scala 50:57:@54710.4]
  wire [10:0] _T_100429; // @[Modules.scala 50:57:@54711.4]
  wire [10:0] buffer_14_496; // @[Modules.scala 50:57:@54712.4]
  wire [10:0] buffer_14_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100437; // @[Modules.scala 50:57:@54722.4]
  wire [10:0] _T_100438; // @[Modules.scala 50:57:@54723.4]
  wire [10:0] buffer_14_499; // @[Modules.scala 50:57:@54724.4]
  wire [10:0] buffer_14_216; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100440; // @[Modules.scala 50:57:@54726.4]
  wire [10:0] _T_100441; // @[Modules.scala 50:57:@54727.4]
  wire [10:0] buffer_14_500; // @[Modules.scala 50:57:@54728.4]
  wire [11:0] _T_100443; // @[Modules.scala 50:57:@54730.4]
  wire [10:0] _T_100444; // @[Modules.scala 50:57:@54731.4]
  wire [10:0] buffer_14_501; // @[Modules.scala 50:57:@54732.4]
  wire [11:0] _T_100464; // @[Modules.scala 50:57:@54758.4]
  wire [10:0] _T_100465; // @[Modules.scala 50:57:@54759.4]
  wire [10:0] buffer_14_508; // @[Modules.scala 50:57:@54760.4]
  wire [11:0] _T_100467; // @[Modules.scala 50:57:@54762.4]
  wire [10:0] _T_100468; // @[Modules.scala 50:57:@54763.4]
  wire [10:0] buffer_14_509; // @[Modules.scala 50:57:@54764.4]
  wire [11:0] _T_100470; // @[Modules.scala 50:57:@54766.4]
  wire [10:0] _T_100471; // @[Modules.scala 50:57:@54767.4]
  wire [10:0] buffer_14_510; // @[Modules.scala 50:57:@54768.4]
  wire [11:0] _T_100473; // @[Modules.scala 50:57:@54770.4]
  wire [10:0] _T_100474; // @[Modules.scala 50:57:@54771.4]
  wire [10:0] buffer_14_511; // @[Modules.scala 50:57:@54772.4]
  wire [11:0] _T_100482; // @[Modules.scala 50:57:@54782.4]
  wire [10:0] _T_100483; // @[Modules.scala 50:57:@54783.4]
  wire [10:0] buffer_14_514; // @[Modules.scala 50:57:@54784.4]
  wire [11:0] _T_100488; // @[Modules.scala 50:57:@54790.4]
  wire [10:0] _T_100489; // @[Modules.scala 50:57:@54791.4]
  wire [10:0] buffer_14_516; // @[Modules.scala 50:57:@54792.4]
  wire [11:0] _T_100494; // @[Modules.scala 50:57:@54798.4]
  wire [10:0] _T_100495; // @[Modules.scala 50:57:@54799.4]
  wire [10:0] buffer_14_518; // @[Modules.scala 50:57:@54800.4]
  wire [11:0] _T_100503; // @[Modules.scala 50:57:@54810.4]
  wire [10:0] _T_100504; // @[Modules.scala 50:57:@54811.4]
  wire [10:0] buffer_14_521; // @[Modules.scala 50:57:@54812.4]
  wire [11:0] _T_100515; // @[Modules.scala 50:57:@54826.4]
  wire [10:0] _T_100516; // @[Modules.scala 50:57:@54827.4]
  wire [10:0] buffer_14_525; // @[Modules.scala 50:57:@54828.4]
  wire [11:0] _T_100521; // @[Modules.scala 50:57:@54834.4]
  wire [10:0] _T_100522; // @[Modules.scala 50:57:@54835.4]
  wire [10:0] buffer_14_527; // @[Modules.scala 50:57:@54836.4]
  wire [11:0] _T_100536; // @[Modules.scala 50:57:@54854.4]
  wire [10:0] _T_100537; // @[Modules.scala 50:57:@54855.4]
  wire [10:0] buffer_14_532; // @[Modules.scala 50:57:@54856.4]
  wire [10:0] buffer_14_284; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100542; // @[Modules.scala 50:57:@54862.4]
  wire [10:0] _T_100543; // @[Modules.scala 50:57:@54863.4]
  wire [10:0] buffer_14_534; // @[Modules.scala 50:57:@54864.4]
  wire [11:0] _T_100548; // @[Modules.scala 50:57:@54870.4]
  wire [10:0] _T_100549; // @[Modules.scala 50:57:@54871.4]
  wire [10:0] buffer_14_536; // @[Modules.scala 50:57:@54872.4]
  wire [11:0] _T_100557; // @[Modules.scala 50:57:@54882.4]
  wire [10:0] _T_100558; // @[Modules.scala 50:57:@54883.4]
  wire [10:0] buffer_14_539; // @[Modules.scala 50:57:@54884.4]
  wire [11:0] _T_100569; // @[Modules.scala 50:57:@54898.4]
  wire [10:0] _T_100570; // @[Modules.scala 50:57:@54899.4]
  wire [10:0] buffer_14_543; // @[Modules.scala 50:57:@54900.4]
  wire [11:0] _T_100578; // @[Modules.scala 50:57:@54910.4]
  wire [10:0] _T_100579; // @[Modules.scala 50:57:@54911.4]
  wire [10:0] buffer_14_546; // @[Modules.scala 50:57:@54912.4]
  wire [11:0] _T_100581; // @[Modules.scala 50:57:@54914.4]
  wire [10:0] _T_100582; // @[Modules.scala 50:57:@54915.4]
  wire [10:0] buffer_14_547; // @[Modules.scala 50:57:@54916.4]
  wire [11:0] _T_100596; // @[Modules.scala 50:57:@54934.4]
  wire [10:0] _T_100597; // @[Modules.scala 50:57:@54935.4]
  wire [10:0] buffer_14_552; // @[Modules.scala 50:57:@54936.4]
  wire [11:0] _T_100605; // @[Modules.scala 50:57:@54946.4]
  wire [10:0] _T_100606; // @[Modules.scala 50:57:@54947.4]
  wire [10:0] buffer_14_555; // @[Modules.scala 50:57:@54948.4]
  wire [11:0] _T_100638; // @[Modules.scala 50:57:@54990.4]
  wire [10:0] _T_100639; // @[Modules.scala 50:57:@54991.4]
  wire [10:0] buffer_14_566; // @[Modules.scala 50:57:@54992.4]
  wire [11:0] _T_100644; // @[Modules.scala 50:57:@54998.4]
  wire [10:0] _T_100645; // @[Modules.scala 50:57:@54999.4]
  wire [10:0] buffer_14_568; // @[Modules.scala 50:57:@55000.4]
  wire [10:0] buffer_14_354; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100647; // @[Modules.scala 50:57:@55002.4]
  wire [10:0] _T_100648; // @[Modules.scala 50:57:@55003.4]
  wire [10:0] buffer_14_569; // @[Modules.scala 50:57:@55004.4]
  wire [11:0] _T_100650; // @[Modules.scala 50:57:@55006.4]
  wire [10:0] _T_100651; // @[Modules.scala 50:57:@55007.4]
  wire [10:0] buffer_14_570; // @[Modules.scala 50:57:@55008.4]
  wire [10:0] buffer_14_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100659; // @[Modules.scala 50:57:@55018.4]
  wire [10:0] _T_100660; // @[Modules.scala 50:57:@55019.4]
  wire [10:0] buffer_14_573; // @[Modules.scala 50:57:@55020.4]
  wire [11:0] _T_100662; // @[Modules.scala 50:57:@55022.4]
  wire [10:0] _T_100663; // @[Modules.scala 50:57:@55023.4]
  wire [10:0] buffer_14_574; // @[Modules.scala 50:57:@55024.4]
  wire [10:0] buffer_14_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100665; // @[Modules.scala 50:57:@55026.4]
  wire [10:0] _T_100666; // @[Modules.scala 50:57:@55027.4]
  wire [10:0] buffer_14_575; // @[Modules.scala 50:57:@55028.4]
  wire [10:0] buffer_14_368; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_14_369; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_100668; // @[Modules.scala 50:57:@55030.4]
  wire [10:0] _T_100669; // @[Modules.scala 50:57:@55031.4]
  wire [10:0] buffer_14_576; // @[Modules.scala 50:57:@55032.4]
  wire [11:0] _T_100671; // @[Modules.scala 50:57:@55034.4]
  wire [10:0] _T_100672; // @[Modules.scala 50:57:@55035.4]
  wire [10:0] buffer_14_577; // @[Modules.scala 50:57:@55036.4]
  wire [11:0] _T_100701; // @[Modules.scala 50:57:@55074.4]
  wire [10:0] _T_100702; // @[Modules.scala 50:57:@55075.4]
  wire [10:0] buffer_14_587; // @[Modules.scala 50:57:@55076.4]
  wire [11:0] _T_100704; // @[Modules.scala 53:83:@55078.4]
  wire [10:0] _T_100705; // @[Modules.scala 53:83:@55079.4]
  wire [10:0] buffer_14_588; // @[Modules.scala 53:83:@55080.4]
  wire [11:0] _T_100707; // @[Modules.scala 53:83:@55082.4]
  wire [10:0] _T_100708; // @[Modules.scala 53:83:@55083.4]
  wire [10:0] buffer_14_589; // @[Modules.scala 53:83:@55084.4]
  wire [11:0] _T_100710; // @[Modules.scala 53:83:@55086.4]
  wire [10:0] _T_100711; // @[Modules.scala 53:83:@55087.4]
  wire [10:0] buffer_14_590; // @[Modules.scala 53:83:@55088.4]
  wire [11:0] _T_100713; // @[Modules.scala 53:83:@55090.4]
  wire [10:0] _T_100714; // @[Modules.scala 53:83:@55091.4]
  wire [10:0] buffer_14_591; // @[Modules.scala 53:83:@55092.4]
  wire [11:0] _T_100716; // @[Modules.scala 53:83:@55094.4]
  wire [10:0] _T_100717; // @[Modules.scala 53:83:@55095.4]
  wire [10:0] buffer_14_592; // @[Modules.scala 53:83:@55096.4]
  wire [11:0] _T_100719; // @[Modules.scala 53:83:@55098.4]
  wire [10:0] _T_100720; // @[Modules.scala 53:83:@55099.4]
  wire [10:0] buffer_14_593; // @[Modules.scala 53:83:@55100.4]
  wire [11:0] _T_100722; // @[Modules.scala 53:83:@55102.4]
  wire [10:0] _T_100723; // @[Modules.scala 53:83:@55103.4]
  wire [10:0] buffer_14_594; // @[Modules.scala 53:83:@55104.4]
  wire [11:0] _T_100725; // @[Modules.scala 53:83:@55106.4]
  wire [10:0] _T_100726; // @[Modules.scala 53:83:@55107.4]
  wire [10:0] buffer_14_595; // @[Modules.scala 53:83:@55108.4]
  wire [11:0] _T_100734; // @[Modules.scala 53:83:@55118.4]
  wire [10:0] _T_100735; // @[Modules.scala 53:83:@55119.4]
  wire [10:0] buffer_14_598; // @[Modules.scala 53:83:@55120.4]
  wire [11:0] _T_100737; // @[Modules.scala 53:83:@55122.4]
  wire [10:0] _T_100738; // @[Modules.scala 53:83:@55123.4]
  wire [10:0] buffer_14_599; // @[Modules.scala 53:83:@55124.4]
  wire [11:0] _T_100740; // @[Modules.scala 53:83:@55126.4]
  wire [10:0] _T_100741; // @[Modules.scala 53:83:@55127.4]
  wire [10:0] buffer_14_600; // @[Modules.scala 53:83:@55128.4]
  wire [11:0] _T_100743; // @[Modules.scala 53:83:@55130.4]
  wire [10:0] _T_100744; // @[Modules.scala 53:83:@55131.4]
  wire [10:0] buffer_14_601; // @[Modules.scala 53:83:@55132.4]
  wire [11:0] _T_100746; // @[Modules.scala 53:83:@55134.4]
  wire [10:0] _T_100747; // @[Modules.scala 53:83:@55135.4]
  wire [10:0] buffer_14_602; // @[Modules.scala 53:83:@55136.4]
  wire [11:0] _T_100749; // @[Modules.scala 53:83:@55138.4]
  wire [10:0] _T_100750; // @[Modules.scala 53:83:@55139.4]
  wire [10:0] buffer_14_603; // @[Modules.scala 53:83:@55140.4]
  wire [11:0] _T_100752; // @[Modules.scala 53:83:@55142.4]
  wire [10:0] _T_100753; // @[Modules.scala 53:83:@55143.4]
  wire [10:0] buffer_14_604; // @[Modules.scala 53:83:@55144.4]
  wire [11:0] _T_100755; // @[Modules.scala 53:83:@55146.4]
  wire [10:0] _T_100756; // @[Modules.scala 53:83:@55147.4]
  wire [10:0] buffer_14_605; // @[Modules.scala 53:83:@55148.4]
  wire [11:0] _T_100758; // @[Modules.scala 53:83:@55150.4]
  wire [10:0] _T_100759; // @[Modules.scala 53:83:@55151.4]
  wire [10:0] buffer_14_606; // @[Modules.scala 53:83:@55152.4]
  wire [11:0] _T_100764; // @[Modules.scala 53:83:@55158.4]
  wire [10:0] _T_100765; // @[Modules.scala 53:83:@55159.4]
  wire [10:0] buffer_14_608; // @[Modules.scala 53:83:@55160.4]
  wire [11:0] _T_100767; // @[Modules.scala 53:83:@55162.4]
  wire [10:0] _T_100768; // @[Modules.scala 53:83:@55163.4]
  wire [10:0] buffer_14_609; // @[Modules.scala 53:83:@55164.4]
  wire [11:0] _T_100770; // @[Modules.scala 53:83:@55166.4]
  wire [10:0] _T_100771; // @[Modules.scala 53:83:@55167.4]
  wire [10:0] buffer_14_610; // @[Modules.scala 53:83:@55168.4]
  wire [11:0] _T_100773; // @[Modules.scala 53:83:@55170.4]
  wire [10:0] _T_100774; // @[Modules.scala 53:83:@55171.4]
  wire [10:0] buffer_14_611; // @[Modules.scala 53:83:@55172.4]
  wire [11:0] _T_100779; // @[Modules.scala 53:83:@55178.4]
  wire [10:0] _T_100780; // @[Modules.scala 53:83:@55179.4]
  wire [10:0] buffer_14_613; // @[Modules.scala 53:83:@55180.4]
  wire [11:0] _T_100782; // @[Modules.scala 53:83:@55182.4]
  wire [10:0] _T_100783; // @[Modules.scala 53:83:@55183.4]
  wire [10:0] buffer_14_614; // @[Modules.scala 53:83:@55184.4]
  wire [11:0] _T_100785; // @[Modules.scala 53:83:@55186.4]
  wire [10:0] _T_100786; // @[Modules.scala 53:83:@55187.4]
  wire [10:0] buffer_14_615; // @[Modules.scala 53:83:@55188.4]
  wire [11:0] _T_100791; // @[Modules.scala 53:83:@55194.4]
  wire [10:0] _T_100792; // @[Modules.scala 53:83:@55195.4]
  wire [10:0] buffer_14_617; // @[Modules.scala 53:83:@55196.4]
  wire [11:0] _T_100794; // @[Modules.scala 53:83:@55198.4]
  wire [10:0] _T_100795; // @[Modules.scala 53:83:@55199.4]
  wire [10:0] buffer_14_618; // @[Modules.scala 53:83:@55200.4]
  wire [11:0] _T_100803; // @[Modules.scala 53:83:@55210.4]
  wire [10:0] _T_100804; // @[Modules.scala 53:83:@55211.4]
  wire [10:0] buffer_14_621; // @[Modules.scala 53:83:@55212.4]
  wire [11:0] _T_100806; // @[Modules.scala 53:83:@55214.4]
  wire [10:0] _T_100807; // @[Modules.scala 53:83:@55215.4]
  wire [10:0] buffer_14_622; // @[Modules.scala 53:83:@55216.4]
  wire [11:0] _T_100812; // @[Modules.scala 53:83:@55222.4]
  wire [10:0] _T_100813; // @[Modules.scala 53:83:@55223.4]
  wire [10:0] buffer_14_624; // @[Modules.scala 53:83:@55224.4]
  wire [11:0] _T_100815; // @[Modules.scala 53:83:@55226.4]
  wire [10:0] _T_100816; // @[Modules.scala 53:83:@55227.4]
  wire [10:0] buffer_14_625; // @[Modules.scala 53:83:@55228.4]
  wire [11:0] _T_100824; // @[Modules.scala 53:83:@55238.4]
  wire [10:0] _T_100825; // @[Modules.scala 53:83:@55239.4]
  wire [10:0] buffer_14_628; // @[Modules.scala 53:83:@55240.4]
  wire [11:0] _T_100827; // @[Modules.scala 53:83:@55242.4]
  wire [10:0] _T_100828; // @[Modules.scala 53:83:@55243.4]
  wire [10:0] buffer_14_629; // @[Modules.scala 53:83:@55244.4]
  wire [11:0] _T_100830; // @[Modules.scala 53:83:@55246.4]
  wire [10:0] _T_100831; // @[Modules.scala 53:83:@55247.4]
  wire [10:0] buffer_14_630; // @[Modules.scala 53:83:@55248.4]
  wire [11:0] _T_100833; // @[Modules.scala 53:83:@55250.4]
  wire [10:0] _T_100834; // @[Modules.scala 53:83:@55251.4]
  wire [10:0] buffer_14_631; // @[Modules.scala 53:83:@55252.4]
  wire [11:0] _T_100839; // @[Modules.scala 53:83:@55258.4]
  wire [10:0] _T_100840; // @[Modules.scala 53:83:@55259.4]
  wire [10:0] buffer_14_633; // @[Modules.scala 53:83:@55260.4]
  wire [11:0] _T_100842; // @[Modules.scala 53:83:@55262.4]
  wire [10:0] _T_100843; // @[Modules.scala 53:83:@55263.4]
  wire [10:0] buffer_14_634; // @[Modules.scala 53:83:@55264.4]
  wire [11:0] _T_100845; // @[Modules.scala 53:83:@55266.4]
  wire [10:0] _T_100846; // @[Modules.scala 53:83:@55267.4]
  wire [10:0] buffer_14_635; // @[Modules.scala 53:83:@55268.4]
  wire [11:0] _T_100848; // @[Modules.scala 53:83:@55270.4]
  wire [10:0] _T_100849; // @[Modules.scala 53:83:@55271.4]
  wire [10:0] buffer_14_636; // @[Modules.scala 53:83:@55272.4]
  wire [11:0] _T_100851; // @[Modules.scala 53:83:@55274.4]
  wire [10:0] _T_100852; // @[Modules.scala 53:83:@55275.4]
  wire [10:0] buffer_14_637; // @[Modules.scala 53:83:@55276.4]
  wire [11:0] _T_100854; // @[Modules.scala 53:83:@55278.4]
  wire [10:0] _T_100855; // @[Modules.scala 53:83:@55279.4]
  wire [10:0] buffer_14_638; // @[Modules.scala 53:83:@55280.4]
  wire [11:0] _T_100857; // @[Modules.scala 53:83:@55282.4]
  wire [10:0] _T_100858; // @[Modules.scala 53:83:@55283.4]
  wire [10:0] buffer_14_639; // @[Modules.scala 53:83:@55284.4]
  wire [11:0] _T_100860; // @[Modules.scala 53:83:@55286.4]
  wire [10:0] _T_100861; // @[Modules.scala 53:83:@55287.4]
  wire [10:0] buffer_14_640; // @[Modules.scala 53:83:@55288.4]
  wire [11:0] _T_100863; // @[Modules.scala 53:83:@55290.4]
  wire [10:0] _T_100864; // @[Modules.scala 53:83:@55291.4]
  wire [10:0] buffer_14_641; // @[Modules.scala 53:83:@55292.4]
  wire [11:0] _T_100866; // @[Modules.scala 53:83:@55294.4]
  wire [10:0] _T_100867; // @[Modules.scala 53:83:@55295.4]
  wire [10:0] buffer_14_642; // @[Modules.scala 53:83:@55296.4]
  wire [11:0] _T_100869; // @[Modules.scala 53:83:@55298.4]
  wire [10:0] _T_100870; // @[Modules.scala 53:83:@55299.4]
  wire [10:0] buffer_14_643; // @[Modules.scala 53:83:@55300.4]
  wire [11:0] _T_100872; // @[Modules.scala 53:83:@55302.4]
  wire [10:0] _T_100873; // @[Modules.scala 53:83:@55303.4]
  wire [10:0] buffer_14_644; // @[Modules.scala 53:83:@55304.4]
  wire [11:0] _T_100878; // @[Modules.scala 53:83:@55310.4]
  wire [10:0] _T_100879; // @[Modules.scala 53:83:@55311.4]
  wire [10:0] buffer_14_646; // @[Modules.scala 53:83:@55312.4]
  wire [11:0] _T_100881; // @[Modules.scala 53:83:@55314.4]
  wire [10:0] _T_100882; // @[Modules.scala 53:83:@55315.4]
  wire [10:0] buffer_14_647; // @[Modules.scala 53:83:@55316.4]
  wire [11:0] _T_100887; // @[Modules.scala 53:83:@55322.4]
  wire [10:0] _T_100888; // @[Modules.scala 53:83:@55323.4]
  wire [10:0] buffer_14_649; // @[Modules.scala 53:83:@55324.4]
  wire [11:0] _T_100890; // @[Modules.scala 53:83:@55326.4]
  wire [10:0] _T_100891; // @[Modules.scala 53:83:@55327.4]
  wire [10:0] buffer_14_650; // @[Modules.scala 53:83:@55328.4]
  wire [11:0] _T_100893; // @[Modules.scala 53:83:@55330.4]
  wire [10:0] _T_100894; // @[Modules.scala 53:83:@55331.4]
  wire [10:0] buffer_14_651; // @[Modules.scala 53:83:@55332.4]
  wire [11:0] _T_100896; // @[Modules.scala 53:83:@55334.4]
  wire [10:0] _T_100897; // @[Modules.scala 53:83:@55335.4]
  wire [10:0] buffer_14_652; // @[Modules.scala 53:83:@55336.4]
  wire [11:0] _T_100899; // @[Modules.scala 53:83:@55338.4]
  wire [10:0] _T_100900; // @[Modules.scala 53:83:@55339.4]
  wire [10:0] buffer_14_653; // @[Modules.scala 53:83:@55340.4]
  wire [11:0] _T_100902; // @[Modules.scala 53:83:@55342.4]
  wire [10:0] _T_100903; // @[Modules.scala 53:83:@55343.4]
  wire [10:0] buffer_14_654; // @[Modules.scala 53:83:@55344.4]
  wire [11:0] _T_100905; // @[Modules.scala 53:83:@55346.4]
  wire [10:0] _T_100906; // @[Modules.scala 53:83:@55347.4]
  wire [10:0] buffer_14_655; // @[Modules.scala 53:83:@55348.4]
  wire [11:0] _T_100908; // @[Modules.scala 53:83:@55350.4]
  wire [10:0] _T_100909; // @[Modules.scala 53:83:@55351.4]
  wire [10:0] buffer_14_656; // @[Modules.scala 53:83:@55352.4]
  wire [11:0] _T_100914; // @[Modules.scala 53:83:@55358.4]
  wire [10:0] _T_100915; // @[Modules.scala 53:83:@55359.4]
  wire [10:0] buffer_14_658; // @[Modules.scala 53:83:@55360.4]
  wire [11:0] _T_100917; // @[Modules.scala 53:83:@55362.4]
  wire [10:0] _T_100918; // @[Modules.scala 53:83:@55363.4]
  wire [10:0] buffer_14_659; // @[Modules.scala 53:83:@55364.4]
  wire [11:0] _T_100920; // @[Modules.scala 53:83:@55366.4]
  wire [10:0] _T_100921; // @[Modules.scala 53:83:@55367.4]
  wire [10:0] buffer_14_660; // @[Modules.scala 53:83:@55368.4]
  wire [11:0] _T_100923; // @[Modules.scala 53:83:@55370.4]
  wire [10:0] _T_100924; // @[Modules.scala 53:83:@55371.4]
  wire [10:0] buffer_14_661; // @[Modules.scala 53:83:@55372.4]
  wire [11:0] _T_100926; // @[Modules.scala 53:83:@55374.4]
  wire [10:0] _T_100927; // @[Modules.scala 53:83:@55375.4]
  wire [10:0] buffer_14_662; // @[Modules.scala 53:83:@55376.4]
  wire [11:0] _T_100929; // @[Modules.scala 53:83:@55378.4]
  wire [10:0] _T_100930; // @[Modules.scala 53:83:@55379.4]
  wire [10:0] buffer_14_663; // @[Modules.scala 53:83:@55380.4]
  wire [11:0] _T_100935; // @[Modules.scala 53:83:@55386.4]
  wire [10:0] _T_100936; // @[Modules.scala 53:83:@55387.4]
  wire [10:0] buffer_14_665; // @[Modules.scala 53:83:@55388.4]
  wire [11:0] _T_100944; // @[Modules.scala 53:83:@55398.4]
  wire [10:0] _T_100945; // @[Modules.scala 53:83:@55399.4]
  wire [10:0] buffer_14_668; // @[Modules.scala 53:83:@55400.4]
  wire [11:0] _T_100947; // @[Modules.scala 53:83:@55402.4]
  wire [10:0] _T_100948; // @[Modules.scala 53:83:@55403.4]
  wire [10:0] buffer_14_669; // @[Modules.scala 53:83:@55404.4]
  wire [11:0] _T_100956; // @[Modules.scala 53:83:@55414.4]
  wire [10:0] _T_100957; // @[Modules.scala 53:83:@55415.4]
  wire [10:0] buffer_14_672; // @[Modules.scala 53:83:@55416.4]
  wire [11:0] _T_100959; // @[Modules.scala 53:83:@55418.4]
  wire [10:0] _T_100960; // @[Modules.scala 53:83:@55419.4]
  wire [10:0] buffer_14_673; // @[Modules.scala 53:83:@55420.4]
  wire [11:0] _T_100965; // @[Modules.scala 53:83:@55426.4]
  wire [10:0] _T_100966; // @[Modules.scala 53:83:@55427.4]
  wire [10:0] buffer_14_675; // @[Modules.scala 53:83:@55428.4]
  wire [11:0] _T_100968; // @[Modules.scala 53:83:@55430.4]
  wire [10:0] _T_100969; // @[Modules.scala 53:83:@55431.4]
  wire [10:0] buffer_14_676; // @[Modules.scala 53:83:@55432.4]
  wire [11:0] _T_100971; // @[Modules.scala 53:83:@55434.4]
  wire [10:0] _T_100972; // @[Modules.scala 53:83:@55435.4]
  wire [10:0] buffer_14_677; // @[Modules.scala 53:83:@55436.4]
  wire [11:0] _T_100974; // @[Modules.scala 53:83:@55438.4]
  wire [10:0] _T_100975; // @[Modules.scala 53:83:@55439.4]
  wire [10:0] buffer_14_678; // @[Modules.scala 53:83:@55440.4]
  wire [11:0] _T_100977; // @[Modules.scala 53:83:@55442.4]
  wire [10:0] _T_100978; // @[Modules.scala 53:83:@55443.4]
  wire [10:0] buffer_14_679; // @[Modules.scala 53:83:@55444.4]
  wire [11:0] _T_100980; // @[Modules.scala 53:83:@55446.4]
  wire [10:0] _T_100981; // @[Modules.scala 53:83:@55447.4]
  wire [10:0] buffer_14_680; // @[Modules.scala 53:83:@55448.4]
  wire [11:0] _T_100983; // @[Modules.scala 53:83:@55450.4]
  wire [10:0] _T_100984; // @[Modules.scala 53:83:@55451.4]
  wire [10:0] buffer_14_681; // @[Modules.scala 53:83:@55452.4]
  wire [11:0] _T_100986; // @[Modules.scala 53:83:@55454.4]
  wire [10:0] _T_100987; // @[Modules.scala 53:83:@55455.4]
  wire [10:0] buffer_14_682; // @[Modules.scala 53:83:@55456.4]
  wire [11:0] _T_100989; // @[Modules.scala 53:83:@55458.4]
  wire [10:0] _T_100990; // @[Modules.scala 53:83:@55459.4]
  wire [10:0] buffer_14_683; // @[Modules.scala 53:83:@55460.4]
  wire [11:0] _T_100995; // @[Modules.scala 53:83:@55466.4]
  wire [10:0] _T_100996; // @[Modules.scala 53:83:@55467.4]
  wire [10:0] buffer_14_685; // @[Modules.scala 53:83:@55468.4]
  wire [11:0] _T_100998; // @[Modules.scala 56:109:@55470.4]
  wire [10:0] _T_100999; // @[Modules.scala 56:109:@55471.4]
  wire [10:0] buffer_14_686; // @[Modules.scala 56:109:@55472.4]
  wire [11:0] _T_101001; // @[Modules.scala 56:109:@55474.4]
  wire [10:0] _T_101002; // @[Modules.scala 56:109:@55475.4]
  wire [10:0] buffer_14_687; // @[Modules.scala 56:109:@55476.4]
  wire [11:0] _T_101004; // @[Modules.scala 56:109:@55478.4]
  wire [10:0] _T_101005; // @[Modules.scala 56:109:@55479.4]
  wire [10:0] buffer_14_688; // @[Modules.scala 56:109:@55480.4]
  wire [11:0] _T_101007; // @[Modules.scala 56:109:@55482.4]
  wire [10:0] _T_101008; // @[Modules.scala 56:109:@55483.4]
  wire [10:0] buffer_14_689; // @[Modules.scala 56:109:@55484.4]
  wire [11:0] _T_101013; // @[Modules.scala 56:109:@55490.4]
  wire [10:0] _T_101014; // @[Modules.scala 56:109:@55491.4]
  wire [10:0] buffer_14_691; // @[Modules.scala 56:109:@55492.4]
  wire [11:0] _T_101016; // @[Modules.scala 56:109:@55494.4]
  wire [10:0] _T_101017; // @[Modules.scala 56:109:@55495.4]
  wire [10:0] buffer_14_692; // @[Modules.scala 56:109:@55496.4]
  wire [11:0] _T_101019; // @[Modules.scala 56:109:@55498.4]
  wire [10:0] _T_101020; // @[Modules.scala 56:109:@55499.4]
  wire [10:0] buffer_14_693; // @[Modules.scala 56:109:@55500.4]
  wire [11:0] _T_101022; // @[Modules.scala 56:109:@55502.4]
  wire [10:0] _T_101023; // @[Modules.scala 56:109:@55503.4]
  wire [10:0] buffer_14_694; // @[Modules.scala 56:109:@55504.4]
  wire [11:0] _T_101025; // @[Modules.scala 56:109:@55506.4]
  wire [10:0] _T_101026; // @[Modules.scala 56:109:@55507.4]
  wire [10:0] buffer_14_695; // @[Modules.scala 56:109:@55508.4]
  wire [11:0] _T_101028; // @[Modules.scala 56:109:@55510.4]
  wire [10:0] _T_101029; // @[Modules.scala 56:109:@55511.4]
  wire [10:0] buffer_14_696; // @[Modules.scala 56:109:@55512.4]
  wire [11:0] _T_101031; // @[Modules.scala 56:109:@55514.4]
  wire [10:0] _T_101032; // @[Modules.scala 56:109:@55515.4]
  wire [10:0] buffer_14_697; // @[Modules.scala 56:109:@55516.4]
  wire [11:0] _T_101034; // @[Modules.scala 56:109:@55518.4]
  wire [10:0] _T_101035; // @[Modules.scala 56:109:@55519.4]
  wire [10:0] buffer_14_698; // @[Modules.scala 56:109:@55520.4]
  wire [11:0] _T_101037; // @[Modules.scala 56:109:@55522.4]
  wire [10:0] _T_101038; // @[Modules.scala 56:109:@55523.4]
  wire [10:0] buffer_14_699; // @[Modules.scala 56:109:@55524.4]
  wire [11:0] _T_101040; // @[Modules.scala 56:109:@55526.4]
  wire [10:0] _T_101041; // @[Modules.scala 56:109:@55527.4]
  wire [10:0] buffer_14_700; // @[Modules.scala 56:109:@55528.4]
  wire [11:0] _T_101043; // @[Modules.scala 56:109:@55530.4]
  wire [10:0] _T_101044; // @[Modules.scala 56:109:@55531.4]
  wire [10:0] buffer_14_701; // @[Modules.scala 56:109:@55532.4]
  wire [11:0] _T_101046; // @[Modules.scala 56:109:@55534.4]
  wire [10:0] _T_101047; // @[Modules.scala 56:109:@55535.4]
  wire [10:0] buffer_14_702; // @[Modules.scala 56:109:@55536.4]
  wire [11:0] _T_101049; // @[Modules.scala 56:109:@55538.4]
  wire [10:0] _T_101050; // @[Modules.scala 56:109:@55539.4]
  wire [10:0] buffer_14_703; // @[Modules.scala 56:109:@55540.4]
  wire [11:0] _T_101052; // @[Modules.scala 56:109:@55542.4]
  wire [10:0] _T_101053; // @[Modules.scala 56:109:@55543.4]
  wire [10:0] buffer_14_704; // @[Modules.scala 56:109:@55544.4]
  wire [11:0] _T_101055; // @[Modules.scala 56:109:@55546.4]
  wire [10:0] _T_101056; // @[Modules.scala 56:109:@55547.4]
  wire [10:0] buffer_14_705; // @[Modules.scala 56:109:@55548.4]
  wire [11:0] _T_101058; // @[Modules.scala 56:109:@55550.4]
  wire [10:0] _T_101059; // @[Modules.scala 56:109:@55551.4]
  wire [10:0] buffer_14_706; // @[Modules.scala 56:109:@55552.4]
  wire [11:0] _T_101061; // @[Modules.scala 56:109:@55554.4]
  wire [10:0] _T_101062; // @[Modules.scala 56:109:@55555.4]
  wire [10:0] buffer_14_707; // @[Modules.scala 56:109:@55556.4]
  wire [11:0] _T_101064; // @[Modules.scala 56:109:@55558.4]
  wire [10:0] _T_101065; // @[Modules.scala 56:109:@55559.4]
  wire [10:0] buffer_14_708; // @[Modules.scala 56:109:@55560.4]
  wire [11:0] _T_101067; // @[Modules.scala 56:109:@55562.4]
  wire [10:0] _T_101068; // @[Modules.scala 56:109:@55563.4]
  wire [10:0] buffer_14_709; // @[Modules.scala 56:109:@55564.4]
  wire [11:0] _T_101070; // @[Modules.scala 56:109:@55566.4]
  wire [10:0] _T_101071; // @[Modules.scala 56:109:@55567.4]
  wire [10:0] buffer_14_710; // @[Modules.scala 56:109:@55568.4]
  wire [11:0] _T_101073; // @[Modules.scala 56:109:@55570.4]
  wire [10:0] _T_101074; // @[Modules.scala 56:109:@55571.4]
  wire [10:0] buffer_14_711; // @[Modules.scala 56:109:@55572.4]
  wire [11:0] _T_101076; // @[Modules.scala 56:109:@55574.4]
  wire [10:0] _T_101077; // @[Modules.scala 56:109:@55575.4]
  wire [10:0] buffer_14_712; // @[Modules.scala 56:109:@55576.4]
  wire [11:0] _T_101079; // @[Modules.scala 56:109:@55578.4]
  wire [10:0] _T_101080; // @[Modules.scala 56:109:@55579.4]
  wire [10:0] buffer_14_713; // @[Modules.scala 56:109:@55580.4]
  wire [11:0] _T_101082; // @[Modules.scala 56:109:@55582.4]
  wire [10:0] _T_101083; // @[Modules.scala 56:109:@55583.4]
  wire [10:0] buffer_14_714; // @[Modules.scala 56:109:@55584.4]
  wire [11:0] _T_101085; // @[Modules.scala 56:109:@55586.4]
  wire [10:0] _T_101086; // @[Modules.scala 56:109:@55587.4]
  wire [10:0] buffer_14_715; // @[Modules.scala 56:109:@55588.4]
  wire [11:0] _T_101088; // @[Modules.scala 56:109:@55590.4]
  wire [10:0] _T_101089; // @[Modules.scala 56:109:@55591.4]
  wire [10:0] buffer_14_716; // @[Modules.scala 56:109:@55592.4]
  wire [11:0] _T_101091; // @[Modules.scala 56:109:@55594.4]
  wire [10:0] _T_101092; // @[Modules.scala 56:109:@55595.4]
  wire [10:0] buffer_14_717; // @[Modules.scala 56:109:@55596.4]
  wire [11:0] _T_101094; // @[Modules.scala 56:109:@55598.4]
  wire [10:0] _T_101095; // @[Modules.scala 56:109:@55599.4]
  wire [10:0] buffer_14_718; // @[Modules.scala 56:109:@55600.4]
  wire [11:0] _T_101097; // @[Modules.scala 56:109:@55602.4]
  wire [10:0] _T_101098; // @[Modules.scala 56:109:@55603.4]
  wire [10:0] buffer_14_719; // @[Modules.scala 56:109:@55604.4]
  wire [11:0] _T_101100; // @[Modules.scala 56:109:@55606.4]
  wire [10:0] _T_101101; // @[Modules.scala 56:109:@55607.4]
  wire [10:0] buffer_14_720; // @[Modules.scala 56:109:@55608.4]
  wire [11:0] _T_101103; // @[Modules.scala 56:109:@55610.4]
  wire [10:0] _T_101104; // @[Modules.scala 56:109:@55611.4]
  wire [10:0] buffer_14_721; // @[Modules.scala 56:109:@55612.4]
  wire [11:0] _T_101106; // @[Modules.scala 56:109:@55614.4]
  wire [10:0] _T_101107; // @[Modules.scala 56:109:@55615.4]
  wire [10:0] buffer_14_722; // @[Modules.scala 56:109:@55616.4]
  wire [11:0] _T_101109; // @[Modules.scala 56:109:@55618.4]
  wire [10:0] _T_101110; // @[Modules.scala 56:109:@55619.4]
  wire [10:0] buffer_14_723; // @[Modules.scala 56:109:@55620.4]
  wire [11:0] _T_101112; // @[Modules.scala 56:109:@55622.4]
  wire [10:0] _T_101113; // @[Modules.scala 56:109:@55623.4]
  wire [10:0] buffer_14_724; // @[Modules.scala 56:109:@55624.4]
  wire [11:0] _T_101115; // @[Modules.scala 56:109:@55626.4]
  wire [10:0] _T_101116; // @[Modules.scala 56:109:@55627.4]
  wire [10:0] buffer_14_725; // @[Modules.scala 56:109:@55628.4]
  wire [11:0] _T_101118; // @[Modules.scala 56:109:@55630.4]
  wire [10:0] _T_101119; // @[Modules.scala 56:109:@55631.4]
  wire [10:0] buffer_14_726; // @[Modules.scala 56:109:@55632.4]
  wire [11:0] _T_101121; // @[Modules.scala 56:109:@55634.4]
  wire [10:0] _T_101122; // @[Modules.scala 56:109:@55635.4]
  wire [10:0] buffer_14_727; // @[Modules.scala 56:109:@55636.4]
  wire [11:0] _T_101124; // @[Modules.scala 56:109:@55638.4]
  wire [10:0] _T_101125; // @[Modules.scala 56:109:@55639.4]
  wire [10:0] buffer_14_728; // @[Modules.scala 56:109:@55640.4]
  wire [11:0] _T_101127; // @[Modules.scala 56:109:@55642.4]
  wire [10:0] _T_101128; // @[Modules.scala 56:109:@55643.4]
  wire [10:0] buffer_14_729; // @[Modules.scala 56:109:@55644.4]
  wire [11:0] _T_101130; // @[Modules.scala 56:109:@55646.4]
  wire [10:0] _T_101131; // @[Modules.scala 56:109:@55647.4]
  wire [10:0] buffer_14_730; // @[Modules.scala 56:109:@55648.4]
  wire [11:0] _T_101133; // @[Modules.scala 56:109:@55650.4]
  wire [10:0] _T_101134; // @[Modules.scala 56:109:@55651.4]
  wire [10:0] buffer_14_731; // @[Modules.scala 56:109:@55652.4]
  wire [11:0] _T_101136; // @[Modules.scala 56:109:@55654.4]
  wire [10:0] _T_101137; // @[Modules.scala 56:109:@55655.4]
  wire [10:0] buffer_14_732; // @[Modules.scala 56:109:@55656.4]
  wire [11:0] _T_101139; // @[Modules.scala 56:109:@55658.4]
  wire [10:0] _T_101140; // @[Modules.scala 56:109:@55659.4]
  wire [10:0] buffer_14_733; // @[Modules.scala 56:109:@55660.4]
  wire [11:0] _T_101142; // @[Modules.scala 56:109:@55662.4]
  wire [10:0] _T_101143; // @[Modules.scala 56:109:@55663.4]
  wire [10:0] buffer_14_734; // @[Modules.scala 56:109:@55664.4]
  wire [11:0] _T_101145; // @[Modules.scala 63:156:@55667.4]
  wire [10:0] _T_101146; // @[Modules.scala 63:156:@55668.4]
  wire [10:0] buffer_14_736; // @[Modules.scala 63:156:@55669.4]
  wire [11:0] _T_101148; // @[Modules.scala 63:156:@55671.4]
  wire [10:0] _T_101149; // @[Modules.scala 63:156:@55672.4]
  wire [10:0] buffer_14_737; // @[Modules.scala 63:156:@55673.4]
  wire [11:0] _T_101151; // @[Modules.scala 63:156:@55675.4]
  wire [10:0] _T_101152; // @[Modules.scala 63:156:@55676.4]
  wire [10:0] buffer_14_738; // @[Modules.scala 63:156:@55677.4]
  wire [11:0] _T_101154; // @[Modules.scala 63:156:@55679.4]
  wire [10:0] _T_101155; // @[Modules.scala 63:156:@55680.4]
  wire [10:0] buffer_14_739; // @[Modules.scala 63:156:@55681.4]
  wire [11:0] _T_101157; // @[Modules.scala 63:156:@55683.4]
  wire [10:0] _T_101158; // @[Modules.scala 63:156:@55684.4]
  wire [10:0] buffer_14_740; // @[Modules.scala 63:156:@55685.4]
  wire [11:0] _T_101160; // @[Modules.scala 63:156:@55687.4]
  wire [10:0] _T_101161; // @[Modules.scala 63:156:@55688.4]
  wire [10:0] buffer_14_741; // @[Modules.scala 63:156:@55689.4]
  wire [11:0] _T_101163; // @[Modules.scala 63:156:@55691.4]
  wire [10:0] _T_101164; // @[Modules.scala 63:156:@55692.4]
  wire [10:0] buffer_14_742; // @[Modules.scala 63:156:@55693.4]
  wire [11:0] _T_101166; // @[Modules.scala 63:156:@55695.4]
  wire [10:0] _T_101167; // @[Modules.scala 63:156:@55696.4]
  wire [10:0] buffer_14_743; // @[Modules.scala 63:156:@55697.4]
  wire [11:0] _T_101169; // @[Modules.scala 63:156:@55699.4]
  wire [10:0] _T_101170; // @[Modules.scala 63:156:@55700.4]
  wire [10:0] buffer_14_744; // @[Modules.scala 63:156:@55701.4]
  wire [11:0] _T_101172; // @[Modules.scala 63:156:@55703.4]
  wire [10:0] _T_101173; // @[Modules.scala 63:156:@55704.4]
  wire [10:0] buffer_14_745; // @[Modules.scala 63:156:@55705.4]
  wire [11:0] _T_101175; // @[Modules.scala 63:156:@55707.4]
  wire [10:0] _T_101176; // @[Modules.scala 63:156:@55708.4]
  wire [10:0] buffer_14_746; // @[Modules.scala 63:156:@55709.4]
  wire [11:0] _T_101178; // @[Modules.scala 63:156:@55711.4]
  wire [10:0] _T_101179; // @[Modules.scala 63:156:@55712.4]
  wire [10:0] buffer_14_747; // @[Modules.scala 63:156:@55713.4]
  wire [11:0] _T_101181; // @[Modules.scala 63:156:@55715.4]
  wire [10:0] _T_101182; // @[Modules.scala 63:156:@55716.4]
  wire [10:0] buffer_14_748; // @[Modules.scala 63:156:@55717.4]
  wire [11:0] _T_101184; // @[Modules.scala 63:156:@55719.4]
  wire [10:0] _T_101185; // @[Modules.scala 63:156:@55720.4]
  wire [10:0] buffer_14_749; // @[Modules.scala 63:156:@55721.4]
  wire [11:0] _T_101187; // @[Modules.scala 63:156:@55723.4]
  wire [10:0] _T_101188; // @[Modules.scala 63:156:@55724.4]
  wire [10:0] buffer_14_750; // @[Modules.scala 63:156:@55725.4]
  wire [11:0] _T_101190; // @[Modules.scala 63:156:@55727.4]
  wire [10:0] _T_101191; // @[Modules.scala 63:156:@55728.4]
  wire [10:0] buffer_14_751; // @[Modules.scala 63:156:@55729.4]
  wire [11:0] _T_101193; // @[Modules.scala 63:156:@55731.4]
  wire [10:0] _T_101194; // @[Modules.scala 63:156:@55732.4]
  wire [10:0] buffer_14_752; // @[Modules.scala 63:156:@55733.4]
  wire [11:0] _T_101196; // @[Modules.scala 63:156:@55735.4]
  wire [10:0] _T_101197; // @[Modules.scala 63:156:@55736.4]
  wire [10:0] buffer_14_753; // @[Modules.scala 63:156:@55737.4]
  wire [11:0] _T_101199; // @[Modules.scala 63:156:@55739.4]
  wire [10:0] _T_101200; // @[Modules.scala 63:156:@55740.4]
  wire [10:0] buffer_14_754; // @[Modules.scala 63:156:@55741.4]
  wire [11:0] _T_101202; // @[Modules.scala 63:156:@55743.4]
  wire [10:0] _T_101203; // @[Modules.scala 63:156:@55744.4]
  wire [10:0] buffer_14_755; // @[Modules.scala 63:156:@55745.4]
  wire [11:0] _T_101205; // @[Modules.scala 63:156:@55747.4]
  wire [10:0] _T_101206; // @[Modules.scala 63:156:@55748.4]
  wire [10:0] buffer_14_756; // @[Modules.scala 63:156:@55749.4]
  wire [11:0] _T_101208; // @[Modules.scala 63:156:@55751.4]
  wire [10:0] _T_101209; // @[Modules.scala 63:156:@55752.4]
  wire [10:0] buffer_14_757; // @[Modules.scala 63:156:@55753.4]
  wire [11:0] _T_101211; // @[Modules.scala 63:156:@55755.4]
  wire [10:0] _T_101212; // @[Modules.scala 63:156:@55756.4]
  wire [10:0] buffer_14_758; // @[Modules.scala 63:156:@55757.4]
  wire [11:0] _T_101214; // @[Modules.scala 63:156:@55759.4]
  wire [10:0] _T_101215; // @[Modules.scala 63:156:@55760.4]
  wire [10:0] buffer_14_759; // @[Modules.scala 63:156:@55761.4]
  wire [11:0] _T_101217; // @[Modules.scala 63:156:@55763.4]
  wire [10:0] _T_101218; // @[Modules.scala 63:156:@55764.4]
  wire [10:0] buffer_14_760; // @[Modules.scala 63:156:@55765.4]
  wire [11:0] _T_101220; // @[Modules.scala 63:156:@55767.4]
  wire [10:0] _T_101221; // @[Modules.scala 63:156:@55768.4]
  wire [10:0] buffer_14_761; // @[Modules.scala 63:156:@55769.4]
  wire [11:0] _T_101223; // @[Modules.scala 63:156:@55771.4]
  wire [10:0] _T_101224; // @[Modules.scala 63:156:@55772.4]
  wire [10:0] buffer_14_762; // @[Modules.scala 63:156:@55773.4]
  wire [11:0] _T_101226; // @[Modules.scala 63:156:@55775.4]
  wire [10:0] _T_101227; // @[Modules.scala 63:156:@55776.4]
  wire [10:0] buffer_14_763; // @[Modules.scala 63:156:@55777.4]
  wire [11:0] _T_101229; // @[Modules.scala 63:156:@55779.4]
  wire [10:0] _T_101230; // @[Modules.scala 63:156:@55780.4]
  wire [10:0] buffer_14_764; // @[Modules.scala 63:156:@55781.4]
  wire [11:0] _T_101232; // @[Modules.scala 63:156:@55783.4]
  wire [10:0] _T_101233; // @[Modules.scala 63:156:@55784.4]
  wire [10:0] buffer_14_765; // @[Modules.scala 63:156:@55785.4]
  wire [11:0] _T_101235; // @[Modules.scala 63:156:@55787.4]
  wire [10:0] _T_101236; // @[Modules.scala 63:156:@55788.4]
  wire [10:0] buffer_14_766; // @[Modules.scala 63:156:@55789.4]
  wire [11:0] _T_101238; // @[Modules.scala 63:156:@55791.4]
  wire [10:0] _T_101239; // @[Modules.scala 63:156:@55792.4]
  wire [10:0] buffer_14_767; // @[Modules.scala 63:156:@55793.4]
  wire [11:0] _T_101241; // @[Modules.scala 63:156:@55795.4]
  wire [10:0] _T_101242; // @[Modules.scala 63:156:@55796.4]
  wire [10:0] buffer_14_768; // @[Modules.scala 63:156:@55797.4]
  wire [11:0] _T_101244; // @[Modules.scala 63:156:@55799.4]
  wire [10:0] _T_101245; // @[Modules.scala 63:156:@55800.4]
  wire [10:0] buffer_14_769; // @[Modules.scala 63:156:@55801.4]
  wire [11:0] _T_101247; // @[Modules.scala 63:156:@55803.4]
  wire [10:0] _T_101248; // @[Modules.scala 63:156:@55804.4]
  wire [10:0] buffer_14_770; // @[Modules.scala 63:156:@55805.4]
  wire [11:0] _T_101250; // @[Modules.scala 63:156:@55807.4]
  wire [10:0] _T_101251; // @[Modules.scala 63:156:@55808.4]
  wire [10:0] buffer_14_771; // @[Modules.scala 63:156:@55809.4]
  wire [11:0] _T_101253; // @[Modules.scala 63:156:@55811.4]
  wire [10:0] _T_101254; // @[Modules.scala 63:156:@55812.4]
  wire [10:0] buffer_14_772; // @[Modules.scala 63:156:@55813.4]
  wire [11:0] _T_101256; // @[Modules.scala 63:156:@55815.4]
  wire [10:0] _T_101257; // @[Modules.scala 63:156:@55816.4]
  wire [10:0] buffer_14_773; // @[Modules.scala 63:156:@55817.4]
  wire [11:0] _T_101259; // @[Modules.scala 63:156:@55819.4]
  wire [10:0] _T_101260; // @[Modules.scala 63:156:@55820.4]
  wire [10:0] buffer_14_774; // @[Modules.scala 63:156:@55821.4]
  wire [11:0] _T_101262; // @[Modules.scala 63:156:@55823.4]
  wire [10:0] _T_101263; // @[Modules.scala 63:156:@55824.4]
  wire [10:0] buffer_14_775; // @[Modules.scala 63:156:@55825.4]
  wire [11:0] _T_101265; // @[Modules.scala 63:156:@55827.4]
  wire [10:0] _T_101266; // @[Modules.scala 63:156:@55828.4]
  wire [10:0] buffer_14_776; // @[Modules.scala 63:156:@55829.4]
  wire [11:0] _T_101268; // @[Modules.scala 63:156:@55831.4]
  wire [10:0] _T_101269; // @[Modules.scala 63:156:@55832.4]
  wire [10:0] buffer_14_777; // @[Modules.scala 63:156:@55833.4]
  wire [11:0] _T_101271; // @[Modules.scala 63:156:@55835.4]
  wire [10:0] _T_101272; // @[Modules.scala 63:156:@55836.4]
  wire [10:0] buffer_14_778; // @[Modules.scala 63:156:@55837.4]
  wire [11:0] _T_101274; // @[Modules.scala 63:156:@55839.4]
  wire [10:0] _T_101275; // @[Modules.scala 63:156:@55840.4]
  wire [10:0] buffer_14_779; // @[Modules.scala 63:156:@55841.4]
  wire [11:0] _T_101277; // @[Modules.scala 63:156:@55843.4]
  wire [10:0] _T_101278; // @[Modules.scala 63:156:@55844.4]
  wire [10:0] buffer_14_780; // @[Modules.scala 63:156:@55845.4]
  wire [11:0] _T_101280; // @[Modules.scala 63:156:@55847.4]
  wire [10:0] _T_101281; // @[Modules.scala 63:156:@55848.4]
  wire [10:0] buffer_14_781; // @[Modules.scala 63:156:@55849.4]
  wire [11:0] _T_101283; // @[Modules.scala 63:156:@55851.4]
  wire [10:0] _T_101284; // @[Modules.scala 63:156:@55852.4]
  wire [10:0] buffer_14_782; // @[Modules.scala 63:156:@55853.4]
  wire [11:0] _T_101286; // @[Modules.scala 63:156:@55855.4]
  wire [10:0] _T_101287; // @[Modules.scala 63:156:@55856.4]
  wire [10:0] buffer_14_783; // @[Modules.scala 63:156:@55857.4]
  wire [5:0] _T_101401; // @[Modules.scala 40:46:@55986.4]
  wire [4:0] _T_101402; // @[Modules.scala 40:46:@55987.4]
  wire [4:0] _T_101403; // @[Modules.scala 40:46:@55988.4]
  wire [5:0] _T_101459; // @[Modules.scala 43:47:@56054.4]
  wire [4:0] _T_101460; // @[Modules.scala 43:47:@56055.4]
  wire [4:0] _T_101461; // @[Modules.scala 43:47:@56056.4]
  wire [5:0] _T_101932; // @[Modules.scala 43:47:@56568.4]
  wire [4:0] _T_101933; // @[Modules.scala 43:47:@56569.4]
  wire [4:0] _T_101934; // @[Modules.scala 43:47:@56570.4]
  wire [5:0] _T_102198; // @[Modules.scala 37:46:@56862.4]
  wire [4:0] _T_102199; // @[Modules.scala 37:46:@56863.4]
  wire [4:0] _T_102200; // @[Modules.scala 37:46:@56864.4]
  wire [5:0] _T_102496; // @[Modules.scala 40:46:@57201.4]
  wire [4:0] _T_102497; // @[Modules.scala 40:46:@57202.4]
  wire [4:0] _T_102498; // @[Modules.scala 40:46:@57203.4]
  wire [5:0] _T_102670; // @[Modules.scala 40:46:@57398.4]
  wire [4:0] _T_102671; // @[Modules.scala 40:46:@57399.4]
  wire [4:0] _T_102672; // @[Modules.scala 40:46:@57400.4]
  wire [5:0] _T_102769; // @[Modules.scala 40:46:@57509.4]
  wire [4:0] _T_102770; // @[Modules.scala 40:46:@57510.4]
  wire [4:0] _T_102771; // @[Modules.scala 40:46:@57511.4]
  wire [5:0] _T_102935; // @[Modules.scala 43:47:@57686.4]
  wire [4:0] _T_102936; // @[Modules.scala 43:47:@57687.4]
  wire [4:0] _T_102937; // @[Modules.scala 43:47:@57688.4]
  wire [5:0] _T_103033; // @[Modules.scala 43:47:@57791.4]
  wire [4:0] _T_103034; // @[Modules.scala 43:47:@57792.4]
  wire [4:0] _T_103035; // @[Modules.scala 43:47:@57793.4]
  wire [5:0] _T_103087; // @[Modules.scala 43:47:@57849.4]
  wire [4:0] _T_103088; // @[Modules.scala 43:47:@57850.4]
  wire [4:0] _T_103089; // @[Modules.scala 43:47:@57851.4]
  wire [5:0] _T_103176; // @[Modules.scala 40:46:@57956.4]
  wire [4:0] _T_103177; // @[Modules.scala 40:46:@57957.4]
  wire [4:0] _T_103178; // @[Modules.scala 40:46:@57958.4]
  wire [11:0] _T_103198; // @[Modules.scala 50:57:@57983.4]
  wire [10:0] _T_103199; // @[Modules.scala 50:57:@57984.4]
  wire [10:0] buffer_15_395; // @[Modules.scala 50:57:@57985.4]
  wire [11:0] _T_103201; // @[Modules.scala 50:57:@57987.4]
  wire [10:0] _T_103202; // @[Modules.scala 50:57:@57988.4]
  wire [10:0] buffer_15_396; // @[Modules.scala 50:57:@57989.4]
  wire [11:0] _T_103204; // @[Modules.scala 50:57:@57991.4]
  wire [10:0] _T_103205; // @[Modules.scala 50:57:@57992.4]
  wire [10:0] buffer_15_397; // @[Modules.scala 50:57:@57993.4]
  wire [11:0] _T_103207; // @[Modules.scala 50:57:@57995.4]
  wire [10:0] _T_103208; // @[Modules.scala 50:57:@57996.4]
  wire [10:0] buffer_15_398; // @[Modules.scala 50:57:@57997.4]
  wire [11:0] _T_103216; // @[Modules.scala 50:57:@58007.4]
  wire [10:0] _T_103217; // @[Modules.scala 50:57:@58008.4]
  wire [10:0] buffer_15_401; // @[Modules.scala 50:57:@58009.4]
  wire [11:0] _T_103222; // @[Modules.scala 50:57:@58015.4]
  wire [10:0] _T_103223; // @[Modules.scala 50:57:@58016.4]
  wire [10:0] buffer_15_403; // @[Modules.scala 50:57:@58017.4]
  wire [10:0] buffer_15_24; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103225; // @[Modules.scala 50:57:@58019.4]
  wire [10:0] _T_103226; // @[Modules.scala 50:57:@58020.4]
  wire [10:0] buffer_15_404; // @[Modules.scala 50:57:@58021.4]
  wire [11:0] _T_103228; // @[Modules.scala 50:57:@58023.4]
  wire [10:0] _T_103229; // @[Modules.scala 50:57:@58024.4]
  wire [10:0] buffer_15_405; // @[Modules.scala 50:57:@58025.4]
  wire [10:0] buffer_15_38; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103246; // @[Modules.scala 50:57:@58047.4]
  wire [10:0] _T_103247; // @[Modules.scala 50:57:@58048.4]
  wire [10:0] buffer_15_411; // @[Modules.scala 50:57:@58049.4]
  wire [11:0] _T_103252; // @[Modules.scala 50:57:@58055.4]
  wire [10:0] _T_103253; // @[Modules.scala 50:57:@58056.4]
  wire [10:0] buffer_15_413; // @[Modules.scala 50:57:@58057.4]
  wire [11:0] _T_103255; // @[Modules.scala 50:57:@58059.4]
  wire [10:0] _T_103256; // @[Modules.scala 50:57:@58060.4]
  wire [10:0] buffer_15_414; // @[Modules.scala 50:57:@58061.4]
  wire [11:0] _T_103279; // @[Modules.scala 50:57:@58091.4]
  wire [10:0] _T_103280; // @[Modules.scala 50:57:@58092.4]
  wire [10:0] buffer_15_422; // @[Modules.scala 50:57:@58093.4]
  wire [11:0] _T_103285; // @[Modules.scala 50:57:@58099.4]
  wire [10:0] _T_103286; // @[Modules.scala 50:57:@58100.4]
  wire [10:0] buffer_15_424; // @[Modules.scala 50:57:@58101.4]
  wire [11:0] _T_103294; // @[Modules.scala 50:57:@58111.4]
  wire [10:0] _T_103295; // @[Modules.scala 50:57:@58112.4]
  wire [10:0] buffer_15_427; // @[Modules.scala 50:57:@58113.4]
  wire [11:0] _T_103303; // @[Modules.scala 50:57:@58123.4]
  wire [10:0] _T_103304; // @[Modules.scala 50:57:@58124.4]
  wire [10:0] buffer_15_430; // @[Modules.scala 50:57:@58125.4]
  wire [11:0] _T_103306; // @[Modules.scala 50:57:@58127.4]
  wire [10:0] _T_103307; // @[Modules.scala 50:57:@58128.4]
  wire [10:0] buffer_15_431; // @[Modules.scala 50:57:@58129.4]
  wire [11:0] _T_103312; // @[Modules.scala 50:57:@58135.4]
  wire [10:0] _T_103313; // @[Modules.scala 50:57:@58136.4]
  wire [10:0] buffer_15_433; // @[Modules.scala 50:57:@58137.4]
  wire [11:0] _T_103315; // @[Modules.scala 50:57:@58139.4]
  wire [10:0] _T_103316; // @[Modules.scala 50:57:@58140.4]
  wire [10:0] buffer_15_434; // @[Modules.scala 50:57:@58141.4]
  wire [11:0] _T_103318; // @[Modules.scala 50:57:@58143.4]
  wire [10:0] _T_103319; // @[Modules.scala 50:57:@58144.4]
  wire [10:0] buffer_15_435; // @[Modules.scala 50:57:@58145.4]
  wire [11:0] _T_103321; // @[Modules.scala 50:57:@58147.4]
  wire [10:0] _T_103322; // @[Modules.scala 50:57:@58148.4]
  wire [10:0] buffer_15_436; // @[Modules.scala 50:57:@58149.4]
  wire [11:0] _T_103336; // @[Modules.scala 50:57:@58167.4]
  wire [10:0] _T_103337; // @[Modules.scala 50:57:@58168.4]
  wire [10:0] buffer_15_441; // @[Modules.scala 50:57:@58169.4]
  wire [11:0] _T_103339; // @[Modules.scala 50:57:@58171.4]
  wire [10:0] _T_103340; // @[Modules.scala 50:57:@58172.4]
  wire [10:0] buffer_15_442; // @[Modules.scala 50:57:@58173.4]
  wire [11:0] _T_103348; // @[Modules.scala 50:57:@58183.4]
  wire [10:0] _T_103349; // @[Modules.scala 50:57:@58184.4]
  wire [10:0] buffer_15_445; // @[Modules.scala 50:57:@58185.4]
  wire [11:0] _T_103363; // @[Modules.scala 50:57:@58203.4]
  wire [10:0] _T_103364; // @[Modules.scala 50:57:@58204.4]
  wire [10:0] buffer_15_450; // @[Modules.scala 50:57:@58205.4]
  wire [10:0] buffer_15_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103381; // @[Modules.scala 50:57:@58227.4]
  wire [10:0] _T_103382; // @[Modules.scala 50:57:@58228.4]
  wire [10:0] buffer_15_456; // @[Modules.scala 50:57:@58229.4]
  wire [11:0] _T_103402; // @[Modules.scala 50:57:@58255.4]
  wire [10:0] _T_103403; // @[Modules.scala 50:57:@58256.4]
  wire [10:0] buffer_15_463; // @[Modules.scala 50:57:@58257.4]
  wire [11:0] _T_103414; // @[Modules.scala 50:57:@58271.4]
  wire [10:0] _T_103415; // @[Modules.scala 50:57:@58272.4]
  wire [10:0] buffer_15_467; // @[Modules.scala 50:57:@58273.4]
  wire [11:0] _T_103423; // @[Modules.scala 50:57:@58283.4]
  wire [10:0] _T_103424; // @[Modules.scala 50:57:@58284.4]
  wire [10:0] buffer_15_470; // @[Modules.scala 50:57:@58285.4]
  wire [11:0] _T_103426; // @[Modules.scala 50:57:@58287.4]
  wire [10:0] _T_103427; // @[Modules.scala 50:57:@58288.4]
  wire [10:0] buffer_15_471; // @[Modules.scala 50:57:@58289.4]
  wire [11:0] _T_103432; // @[Modules.scala 50:57:@58295.4]
  wire [10:0] _T_103433; // @[Modules.scala 50:57:@58296.4]
  wire [10:0] buffer_15_473; // @[Modules.scala 50:57:@58297.4]
  wire [11:0] _T_103441; // @[Modules.scala 50:57:@58307.4]
  wire [10:0] _T_103442; // @[Modules.scala 50:57:@58308.4]
  wire [10:0] buffer_15_476; // @[Modules.scala 50:57:@58309.4]
  wire [11:0] _T_103459; // @[Modules.scala 50:57:@58331.4]
  wire [10:0] _T_103460; // @[Modules.scala 50:57:@58332.4]
  wire [10:0] buffer_15_482; // @[Modules.scala 50:57:@58333.4]
  wire [10:0] buffer_15_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103462; // @[Modules.scala 50:57:@58335.4]
  wire [10:0] _T_103463; // @[Modules.scala 50:57:@58336.4]
  wire [10:0] buffer_15_483; // @[Modules.scala 50:57:@58337.4]
  wire [11:0] _T_103465; // @[Modules.scala 50:57:@58339.4]
  wire [10:0] _T_103466; // @[Modules.scala 50:57:@58340.4]
  wire [10:0] buffer_15_484; // @[Modules.scala 50:57:@58341.4]
  wire [11:0] _T_103495; // @[Modules.scala 50:57:@58379.4]
  wire [10:0] _T_103496; // @[Modules.scala 50:57:@58380.4]
  wire [10:0] buffer_15_494; // @[Modules.scala 50:57:@58381.4]
  wire [11:0] _T_103516; // @[Modules.scala 50:57:@58407.4]
  wire [10:0] _T_103517; // @[Modules.scala 50:57:@58408.4]
  wire [10:0] buffer_15_501; // @[Modules.scala 50:57:@58409.4]
  wire [11:0] _T_103531; // @[Modules.scala 50:57:@58427.4]
  wire [10:0] _T_103532; // @[Modules.scala 50:57:@58428.4]
  wire [10:0] buffer_15_506; // @[Modules.scala 50:57:@58429.4]
  wire [11:0] _T_103534; // @[Modules.scala 50:57:@58431.4]
  wire [10:0] _T_103535; // @[Modules.scala 50:57:@58432.4]
  wire [10:0] buffer_15_507; // @[Modules.scala 50:57:@58433.4]
  wire [11:0] _T_103558; // @[Modules.scala 50:57:@58463.4]
  wire [10:0] _T_103559; // @[Modules.scala 50:57:@58464.4]
  wire [10:0] buffer_15_515; // @[Modules.scala 50:57:@58465.4]
  wire [10:0] buffer_15_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103561; // @[Modules.scala 50:57:@58467.4]
  wire [10:0] _T_103562; // @[Modules.scala 50:57:@58468.4]
  wire [10:0] buffer_15_516; // @[Modules.scala 50:57:@58469.4]
  wire [11:0] _T_103582; // @[Modules.scala 50:57:@58495.4]
  wire [10:0] _T_103583; // @[Modules.scala 50:57:@58496.4]
  wire [10:0] buffer_15_523; // @[Modules.scala 50:57:@58497.4]
  wire [11:0] _T_103597; // @[Modules.scala 50:57:@58515.4]
  wire [10:0] _T_103598; // @[Modules.scala 50:57:@58516.4]
  wire [10:0] buffer_15_528; // @[Modules.scala 50:57:@58517.4]
  wire [11:0] _T_103600; // @[Modules.scala 50:57:@58519.4]
  wire [10:0] _T_103601; // @[Modules.scala 50:57:@58520.4]
  wire [10:0] buffer_15_529; // @[Modules.scala 50:57:@58521.4]
  wire [11:0] _T_103615; // @[Modules.scala 50:57:@58539.4]
  wire [10:0] _T_103616; // @[Modules.scala 50:57:@58540.4]
  wire [10:0] buffer_15_534; // @[Modules.scala 50:57:@58541.4]
  wire [10:0] buffer_15_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103618; // @[Modules.scala 50:57:@58543.4]
  wire [10:0] _T_103619; // @[Modules.scala 50:57:@58544.4]
  wire [10:0] buffer_15_535; // @[Modules.scala 50:57:@58545.4]
  wire [11:0] _T_103621; // @[Modules.scala 50:57:@58547.4]
  wire [10:0] _T_103622; // @[Modules.scala 50:57:@58548.4]
  wire [10:0] buffer_15_536; // @[Modules.scala 50:57:@58549.4]
  wire [11:0] _T_103630; // @[Modules.scala 50:57:@58559.4]
  wire [10:0] _T_103631; // @[Modules.scala 50:57:@58560.4]
  wire [10:0] buffer_15_539; // @[Modules.scala 50:57:@58561.4]
  wire [11:0] _T_103636; // @[Modules.scala 50:57:@58567.4]
  wire [10:0] _T_103637; // @[Modules.scala 50:57:@58568.4]
  wire [10:0] buffer_15_541; // @[Modules.scala 50:57:@58569.4]
  wire [11:0] _T_103639; // @[Modules.scala 50:57:@58571.4]
  wire [10:0] _T_103640; // @[Modules.scala 50:57:@58572.4]
  wire [10:0] buffer_15_542; // @[Modules.scala 50:57:@58573.4]
  wire [11:0] _T_103642; // @[Modules.scala 50:57:@58575.4]
  wire [10:0] _T_103643; // @[Modules.scala 50:57:@58576.4]
  wire [10:0] buffer_15_543; // @[Modules.scala 50:57:@58577.4]
  wire [11:0] _T_103645; // @[Modules.scala 50:57:@58579.4]
  wire [10:0] _T_103646; // @[Modules.scala 50:57:@58580.4]
  wire [10:0] buffer_15_544; // @[Modules.scala 50:57:@58581.4]
  wire [10:0] buffer_15_308; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103651; // @[Modules.scala 50:57:@58587.4]
  wire [10:0] _T_103652; // @[Modules.scala 50:57:@58588.4]
  wire [10:0] buffer_15_546; // @[Modules.scala 50:57:@58589.4]
  wire [11:0] _T_103654; // @[Modules.scala 50:57:@58591.4]
  wire [10:0] _T_103655; // @[Modules.scala 50:57:@58592.4]
  wire [10:0] buffer_15_547; // @[Modules.scala 50:57:@58593.4]
  wire [11:0] _T_103660; // @[Modules.scala 50:57:@58599.4]
  wire [10:0] _T_103661; // @[Modules.scala 50:57:@58600.4]
  wire [10:0] buffer_15_549; // @[Modules.scala 50:57:@58601.4]
  wire [11:0] _T_103669; // @[Modules.scala 50:57:@58611.4]
  wire [10:0] _T_103670; // @[Modules.scala 50:57:@58612.4]
  wire [10:0] buffer_15_552; // @[Modules.scala 50:57:@58613.4]
  wire [11:0] _T_103672; // @[Modules.scala 50:57:@58615.4]
  wire [10:0] _T_103673; // @[Modules.scala 50:57:@58616.4]
  wire [10:0] buffer_15_553; // @[Modules.scala 50:57:@58617.4]
  wire [11:0] _T_103675; // @[Modules.scala 50:57:@58619.4]
  wire [10:0] _T_103676; // @[Modules.scala 50:57:@58620.4]
  wire [10:0] buffer_15_554; // @[Modules.scala 50:57:@58621.4]
  wire [10:0] buffer_15_338; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103696; // @[Modules.scala 50:57:@58647.4]
  wire [10:0] _T_103697; // @[Modules.scala 50:57:@58648.4]
  wire [10:0] buffer_15_561; // @[Modules.scala 50:57:@58649.4]
  wire [11:0] _T_103699; // @[Modules.scala 50:57:@58651.4]
  wire [10:0] _T_103700; // @[Modules.scala 50:57:@58652.4]
  wire [10:0] buffer_15_562; // @[Modules.scala 50:57:@58653.4]
  wire [11:0] _T_103714; // @[Modules.scala 50:57:@58671.4]
  wire [10:0] _T_103715; // @[Modules.scala 50:57:@58672.4]
  wire [10:0] buffer_15_567; // @[Modules.scala 50:57:@58673.4]
  wire [11:0] _T_103717; // @[Modules.scala 50:57:@58675.4]
  wire [10:0] _T_103718; // @[Modules.scala 50:57:@58676.4]
  wire [10:0] buffer_15_568; // @[Modules.scala 50:57:@58677.4]
  wire [10:0] buffer_15_356; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103723; // @[Modules.scala 50:57:@58683.4]
  wire [10:0] _T_103724; // @[Modules.scala 50:57:@58684.4]
  wire [10:0] buffer_15_570; // @[Modules.scala 50:57:@58685.4]
  wire [10:0] buffer_15_366; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103738; // @[Modules.scala 50:57:@58703.4]
  wire [10:0] _T_103739; // @[Modules.scala 50:57:@58704.4]
  wire [10:0] buffer_15_575; // @[Modules.scala 50:57:@58705.4]
  wire [10:0] buffer_15_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_103771; // @[Modules.scala 50:57:@58747.4]
  wire [10:0] _T_103772; // @[Modules.scala 50:57:@58748.4]
  wire [10:0] buffer_15_586; // @[Modules.scala 50:57:@58749.4]
  wire [11:0] _T_103777; // @[Modules.scala 53:83:@58755.4]
  wire [10:0] _T_103778; // @[Modules.scala 53:83:@58756.4]
  wire [10:0] buffer_15_588; // @[Modules.scala 53:83:@58757.4]
  wire [11:0] _T_103780; // @[Modules.scala 53:83:@58759.4]
  wire [10:0] _T_103781; // @[Modules.scala 53:83:@58760.4]
  wire [10:0] buffer_15_589; // @[Modules.scala 53:83:@58761.4]
  wire [11:0] _T_103783; // @[Modules.scala 53:83:@58763.4]
  wire [10:0] _T_103784; // @[Modules.scala 53:83:@58764.4]
  wire [10:0] buffer_15_590; // @[Modules.scala 53:83:@58765.4]
  wire [11:0] _T_103786; // @[Modules.scala 53:83:@58767.4]
  wire [10:0] _T_103787; // @[Modules.scala 53:83:@58768.4]
  wire [10:0] buffer_15_591; // @[Modules.scala 53:83:@58769.4]
  wire [11:0] _T_103789; // @[Modules.scala 53:83:@58771.4]
  wire [10:0] _T_103790; // @[Modules.scala 53:83:@58772.4]
  wire [10:0] buffer_15_592; // @[Modules.scala 53:83:@58773.4]
  wire [11:0] _T_103792; // @[Modules.scala 53:83:@58775.4]
  wire [10:0] _T_103793; // @[Modules.scala 53:83:@58776.4]
  wire [10:0] buffer_15_593; // @[Modules.scala 53:83:@58777.4]
  wire [11:0] _T_103795; // @[Modules.scala 53:83:@58779.4]
  wire [10:0] _T_103796; // @[Modules.scala 53:83:@58780.4]
  wire [10:0] buffer_15_594; // @[Modules.scala 53:83:@58781.4]
  wire [11:0] _T_103798; // @[Modules.scala 53:83:@58783.4]
  wire [10:0] _T_103799; // @[Modules.scala 53:83:@58784.4]
  wire [10:0] buffer_15_595; // @[Modules.scala 53:83:@58785.4]
  wire [11:0] _T_103804; // @[Modules.scala 53:83:@58791.4]
  wire [10:0] _T_103805; // @[Modules.scala 53:83:@58792.4]
  wire [10:0] buffer_15_597; // @[Modules.scala 53:83:@58793.4]
  wire [11:0] _T_103807; // @[Modules.scala 53:83:@58795.4]
  wire [10:0] _T_103808; // @[Modules.scala 53:83:@58796.4]
  wire [10:0] buffer_15_598; // @[Modules.scala 53:83:@58797.4]
  wire [11:0] _T_103810; // @[Modules.scala 53:83:@58799.4]
  wire [10:0] _T_103811; // @[Modules.scala 53:83:@58800.4]
  wire [10:0] buffer_15_599; // @[Modules.scala 53:83:@58801.4]
  wire [11:0] _T_103819; // @[Modules.scala 53:83:@58811.4]
  wire [10:0] _T_103820; // @[Modules.scala 53:83:@58812.4]
  wire [10:0] buffer_15_602; // @[Modules.scala 53:83:@58813.4]
  wire [11:0] _T_103822; // @[Modules.scala 53:83:@58815.4]
  wire [10:0] _T_103823; // @[Modules.scala 53:83:@58816.4]
  wire [10:0] buffer_15_603; // @[Modules.scala 53:83:@58817.4]
  wire [11:0] _T_103825; // @[Modules.scala 53:83:@58819.4]
  wire [10:0] _T_103826; // @[Modules.scala 53:83:@58820.4]
  wire [10:0] buffer_15_604; // @[Modules.scala 53:83:@58821.4]
  wire [11:0] _T_103828; // @[Modules.scala 53:83:@58823.4]
  wire [10:0] _T_103829; // @[Modules.scala 53:83:@58824.4]
  wire [10:0] buffer_15_605; // @[Modules.scala 53:83:@58825.4]
  wire [11:0] _T_103831; // @[Modules.scala 53:83:@58827.4]
  wire [10:0] _T_103832; // @[Modules.scala 53:83:@58828.4]
  wire [10:0] buffer_15_606; // @[Modules.scala 53:83:@58829.4]
  wire [11:0] _T_103834; // @[Modules.scala 53:83:@58831.4]
  wire [10:0] _T_103835; // @[Modules.scala 53:83:@58832.4]
  wire [10:0] buffer_15_607; // @[Modules.scala 53:83:@58833.4]
  wire [11:0] _T_103837; // @[Modules.scala 53:83:@58835.4]
  wire [10:0] _T_103838; // @[Modules.scala 53:83:@58836.4]
  wire [10:0] buffer_15_608; // @[Modules.scala 53:83:@58837.4]
  wire [11:0] _T_103840; // @[Modules.scala 53:83:@58839.4]
  wire [10:0] _T_103841; // @[Modules.scala 53:83:@58840.4]
  wire [10:0] buffer_15_609; // @[Modules.scala 53:83:@58841.4]
  wire [11:0] _T_103843; // @[Modules.scala 53:83:@58843.4]
  wire [10:0] _T_103844; // @[Modules.scala 53:83:@58844.4]
  wire [10:0] buffer_15_610; // @[Modules.scala 53:83:@58845.4]
  wire [11:0] _T_103846; // @[Modules.scala 53:83:@58847.4]
  wire [10:0] _T_103847; // @[Modules.scala 53:83:@58848.4]
  wire [10:0] buffer_15_611; // @[Modules.scala 53:83:@58849.4]
  wire [11:0] _T_103849; // @[Modules.scala 53:83:@58851.4]
  wire [10:0] _T_103850; // @[Modules.scala 53:83:@58852.4]
  wire [10:0] buffer_15_612; // @[Modules.scala 53:83:@58853.4]
  wire [11:0] _T_103852; // @[Modules.scala 53:83:@58855.4]
  wire [10:0] _T_103853; // @[Modules.scala 53:83:@58856.4]
  wire [10:0] buffer_15_613; // @[Modules.scala 53:83:@58857.4]
  wire [11:0] _T_103855; // @[Modules.scala 53:83:@58859.4]
  wire [10:0] _T_103856; // @[Modules.scala 53:83:@58860.4]
  wire [10:0] buffer_15_614; // @[Modules.scala 53:83:@58861.4]
  wire [11:0] _T_103858; // @[Modules.scala 53:83:@58863.4]
  wire [10:0] _T_103859; // @[Modules.scala 53:83:@58864.4]
  wire [10:0] buffer_15_615; // @[Modules.scala 53:83:@58865.4]
  wire [11:0] _T_103861; // @[Modules.scala 53:83:@58867.4]
  wire [10:0] _T_103862; // @[Modules.scala 53:83:@58868.4]
  wire [10:0] buffer_15_616; // @[Modules.scala 53:83:@58869.4]
  wire [11:0] _T_103864; // @[Modules.scala 53:83:@58871.4]
  wire [10:0] _T_103865; // @[Modules.scala 53:83:@58872.4]
  wire [10:0] buffer_15_617; // @[Modules.scala 53:83:@58873.4]
  wire [11:0] _T_103867; // @[Modules.scala 53:83:@58875.4]
  wire [10:0] _T_103868; // @[Modules.scala 53:83:@58876.4]
  wire [10:0] buffer_15_618; // @[Modules.scala 53:83:@58877.4]
  wire [11:0] _T_103873; // @[Modules.scala 53:83:@58883.4]
  wire [10:0] _T_103874; // @[Modules.scala 53:83:@58884.4]
  wire [10:0] buffer_15_620; // @[Modules.scala 53:83:@58885.4]
  wire [11:0] _T_103876; // @[Modules.scala 53:83:@58887.4]
  wire [10:0] _T_103877; // @[Modules.scala 53:83:@58888.4]
  wire [10:0] buffer_15_621; // @[Modules.scala 53:83:@58889.4]
  wire [11:0] _T_103882; // @[Modules.scala 53:83:@58895.4]
  wire [10:0] _T_103883; // @[Modules.scala 53:83:@58896.4]
  wire [10:0] buffer_15_623; // @[Modules.scala 53:83:@58897.4]
  wire [11:0] _T_103888; // @[Modules.scala 53:83:@58903.4]
  wire [10:0] _T_103889; // @[Modules.scala 53:83:@58904.4]
  wire [10:0] buffer_15_625; // @[Modules.scala 53:83:@58905.4]
  wire [11:0] _T_103891; // @[Modules.scala 53:83:@58907.4]
  wire [10:0] _T_103892; // @[Modules.scala 53:83:@58908.4]
  wire [10:0] buffer_15_626; // @[Modules.scala 53:83:@58909.4]
  wire [11:0] _T_103894; // @[Modules.scala 53:83:@58911.4]
  wire [10:0] _T_103895; // @[Modules.scala 53:83:@58912.4]
  wire [10:0] buffer_15_627; // @[Modules.scala 53:83:@58913.4]
  wire [11:0] _T_103897; // @[Modules.scala 53:83:@58915.4]
  wire [10:0] _T_103898; // @[Modules.scala 53:83:@58916.4]
  wire [10:0] buffer_15_628; // @[Modules.scala 53:83:@58917.4]
  wire [11:0] _T_103900; // @[Modules.scala 53:83:@58919.4]
  wire [10:0] _T_103901; // @[Modules.scala 53:83:@58920.4]
  wire [10:0] buffer_15_629; // @[Modules.scala 53:83:@58921.4]
  wire [11:0] _T_103903; // @[Modules.scala 53:83:@58923.4]
  wire [10:0] _T_103904; // @[Modules.scala 53:83:@58924.4]
  wire [10:0] buffer_15_630; // @[Modules.scala 53:83:@58925.4]
  wire [11:0] _T_103909; // @[Modules.scala 53:83:@58931.4]
  wire [10:0] _T_103910; // @[Modules.scala 53:83:@58932.4]
  wire [10:0] buffer_15_632; // @[Modules.scala 53:83:@58933.4]
  wire [11:0] _T_103912; // @[Modules.scala 53:83:@58935.4]
  wire [10:0] _T_103913; // @[Modules.scala 53:83:@58936.4]
  wire [10:0] buffer_15_633; // @[Modules.scala 53:83:@58937.4]
  wire [11:0] _T_103915; // @[Modules.scala 53:83:@58939.4]
  wire [10:0] _T_103916; // @[Modules.scala 53:83:@58940.4]
  wire [10:0] buffer_15_634; // @[Modules.scala 53:83:@58941.4]
  wire [11:0] _T_103921; // @[Modules.scala 53:83:@58947.4]
  wire [10:0] _T_103922; // @[Modules.scala 53:83:@58948.4]
  wire [10:0] buffer_15_636; // @[Modules.scala 53:83:@58949.4]
  wire [11:0] _T_103927; // @[Modules.scala 53:83:@58955.4]
  wire [10:0] _T_103928; // @[Modules.scala 53:83:@58956.4]
  wire [10:0] buffer_15_638; // @[Modules.scala 53:83:@58957.4]
  wire [11:0] _T_103930; // @[Modules.scala 53:83:@58959.4]
  wire [10:0] _T_103931; // @[Modules.scala 53:83:@58960.4]
  wire [10:0] buffer_15_639; // @[Modules.scala 53:83:@58961.4]
  wire [11:0] _T_103933; // @[Modules.scala 53:83:@58963.4]
  wire [10:0] _T_103934; // @[Modules.scala 53:83:@58964.4]
  wire [10:0] buffer_15_640; // @[Modules.scala 53:83:@58965.4]
  wire [11:0] _T_103939; // @[Modules.scala 53:83:@58971.4]
  wire [10:0] _T_103940; // @[Modules.scala 53:83:@58972.4]
  wire [10:0] buffer_15_642; // @[Modules.scala 53:83:@58973.4]
  wire [11:0] _T_103942; // @[Modules.scala 53:83:@58975.4]
  wire [10:0] _T_103943; // @[Modules.scala 53:83:@58976.4]
  wire [10:0] buffer_15_643; // @[Modules.scala 53:83:@58977.4]
  wire [11:0] _T_103948; // @[Modules.scala 53:83:@58983.4]
  wire [10:0] _T_103949; // @[Modules.scala 53:83:@58984.4]
  wire [10:0] buffer_15_645; // @[Modules.scala 53:83:@58985.4]
  wire [11:0] _T_103951; // @[Modules.scala 53:83:@58987.4]
  wire [10:0] _T_103952; // @[Modules.scala 53:83:@58988.4]
  wire [10:0] buffer_15_646; // @[Modules.scala 53:83:@58989.4]
  wire [11:0] _T_103960; // @[Modules.scala 53:83:@58999.4]
  wire [10:0] _T_103961; // @[Modules.scala 53:83:@59000.4]
  wire [10:0] buffer_15_649; // @[Modules.scala 53:83:@59001.4]
  wire [11:0] _T_103963; // @[Modules.scala 53:83:@59003.4]
  wire [10:0] _T_103964; // @[Modules.scala 53:83:@59004.4]
  wire [10:0] buffer_15_650; // @[Modules.scala 53:83:@59005.4]
  wire [11:0] _T_103966; // @[Modules.scala 53:83:@59007.4]
  wire [10:0] _T_103967; // @[Modules.scala 53:83:@59008.4]
  wire [10:0] buffer_15_651; // @[Modules.scala 53:83:@59009.4]
  wire [11:0] _T_103969; // @[Modules.scala 53:83:@59011.4]
  wire [10:0] _T_103970; // @[Modules.scala 53:83:@59012.4]
  wire [10:0] buffer_15_652; // @[Modules.scala 53:83:@59013.4]
  wire [11:0] _T_103972; // @[Modules.scala 53:83:@59015.4]
  wire [10:0] _T_103973; // @[Modules.scala 53:83:@59016.4]
  wire [10:0] buffer_15_653; // @[Modules.scala 53:83:@59017.4]
  wire [11:0] _T_103978; // @[Modules.scala 53:83:@59023.4]
  wire [10:0] _T_103979; // @[Modules.scala 53:83:@59024.4]
  wire [10:0] buffer_15_655; // @[Modules.scala 53:83:@59025.4]
  wire [11:0] _T_103981; // @[Modules.scala 53:83:@59027.4]
  wire [10:0] _T_103982; // @[Modules.scala 53:83:@59028.4]
  wire [10:0] buffer_15_656; // @[Modules.scala 53:83:@59029.4]
  wire [11:0] _T_103990; // @[Modules.scala 53:83:@59039.4]
  wire [10:0] _T_103991; // @[Modules.scala 53:83:@59040.4]
  wire [10:0] buffer_15_659; // @[Modules.scala 53:83:@59041.4]
  wire [11:0] _T_103993; // @[Modules.scala 53:83:@59043.4]
  wire [10:0] _T_103994; // @[Modules.scala 53:83:@59044.4]
  wire [10:0] buffer_15_660; // @[Modules.scala 53:83:@59045.4]
  wire [11:0] _T_103996; // @[Modules.scala 53:83:@59047.4]
  wire [10:0] _T_103997; // @[Modules.scala 53:83:@59048.4]
  wire [10:0] buffer_15_661; // @[Modules.scala 53:83:@59049.4]
  wire [11:0] _T_103999; // @[Modules.scala 53:83:@59051.4]
  wire [10:0] _T_104000; // @[Modules.scala 53:83:@59052.4]
  wire [10:0] buffer_15_662; // @[Modules.scala 53:83:@59053.4]
  wire [11:0] _T_104002; // @[Modules.scala 53:83:@59055.4]
  wire [10:0] _T_104003; // @[Modules.scala 53:83:@59056.4]
  wire [10:0] buffer_15_663; // @[Modules.scala 53:83:@59057.4]
  wire [11:0] _T_104005; // @[Modules.scala 53:83:@59059.4]
  wire [10:0] _T_104006; // @[Modules.scala 53:83:@59060.4]
  wire [10:0] buffer_15_664; // @[Modules.scala 53:83:@59061.4]
  wire [11:0] _T_104008; // @[Modules.scala 53:83:@59063.4]
  wire [10:0] _T_104009; // @[Modules.scala 53:83:@59064.4]
  wire [10:0] buffer_15_665; // @[Modules.scala 53:83:@59065.4]
  wire [11:0] _T_104011; // @[Modules.scala 53:83:@59067.4]
  wire [10:0] _T_104012; // @[Modules.scala 53:83:@59068.4]
  wire [10:0] buffer_15_666; // @[Modules.scala 53:83:@59069.4]
  wire [11:0] _T_104017; // @[Modules.scala 53:83:@59075.4]
  wire [10:0] _T_104018; // @[Modules.scala 53:83:@59076.4]
  wire [10:0] buffer_15_668; // @[Modules.scala 53:83:@59077.4]
  wire [11:0] _T_104020; // @[Modules.scala 53:83:@59079.4]
  wire [10:0] _T_104021; // @[Modules.scala 53:83:@59080.4]
  wire [10:0] buffer_15_669; // @[Modules.scala 53:83:@59081.4]
  wire [11:0] _T_104026; // @[Modules.scala 53:83:@59087.4]
  wire [10:0] _T_104027; // @[Modules.scala 53:83:@59088.4]
  wire [10:0] buffer_15_671; // @[Modules.scala 53:83:@59089.4]
  wire [11:0] _T_104029; // @[Modules.scala 53:83:@59091.4]
  wire [10:0] _T_104030; // @[Modules.scala 53:83:@59092.4]
  wire [10:0] buffer_15_672; // @[Modules.scala 53:83:@59093.4]
  wire [11:0] _T_104032; // @[Modules.scala 53:83:@59095.4]
  wire [10:0] _T_104033; // @[Modules.scala 53:83:@59096.4]
  wire [10:0] buffer_15_673; // @[Modules.scala 53:83:@59097.4]
  wire [11:0] _T_104038; // @[Modules.scala 53:83:@59103.4]
  wire [10:0] _T_104039; // @[Modules.scala 53:83:@59104.4]
  wire [10:0] buffer_15_675; // @[Modules.scala 53:83:@59105.4]
  wire [11:0] _T_104041; // @[Modules.scala 53:83:@59107.4]
  wire [10:0] _T_104042; // @[Modules.scala 53:83:@59108.4]
  wire [10:0] buffer_15_676; // @[Modules.scala 53:83:@59109.4]
  wire [11:0] _T_104044; // @[Modules.scala 53:83:@59111.4]
  wire [10:0] _T_104045; // @[Modules.scala 53:83:@59112.4]
  wire [10:0] buffer_15_677; // @[Modules.scala 53:83:@59113.4]
  wire [11:0] _T_104050; // @[Modules.scala 53:83:@59119.4]
  wire [10:0] _T_104051; // @[Modules.scala 53:83:@59120.4]
  wire [10:0] buffer_15_679; // @[Modules.scala 53:83:@59121.4]
  wire [11:0] _T_104068; // @[Modules.scala 53:83:@59143.4]
  wire [10:0] _T_104069; // @[Modules.scala 53:83:@59144.4]
  wire [10:0] buffer_15_685; // @[Modules.scala 53:83:@59145.4]
  wire [11:0] _T_104071; // @[Modules.scala 56:109:@59147.4]
  wire [10:0] _T_104072; // @[Modules.scala 56:109:@59148.4]
  wire [10:0] buffer_15_686; // @[Modules.scala 56:109:@59149.4]
  wire [11:0] _T_104074; // @[Modules.scala 56:109:@59151.4]
  wire [10:0] _T_104075; // @[Modules.scala 56:109:@59152.4]
  wire [10:0] buffer_15_687; // @[Modules.scala 56:109:@59153.4]
  wire [11:0] _T_104077; // @[Modules.scala 56:109:@59155.4]
  wire [10:0] _T_104078; // @[Modules.scala 56:109:@59156.4]
  wire [10:0] buffer_15_688; // @[Modules.scala 56:109:@59157.4]
  wire [11:0] _T_104080; // @[Modules.scala 56:109:@59159.4]
  wire [10:0] _T_104081; // @[Modules.scala 56:109:@59160.4]
  wire [10:0] buffer_15_689; // @[Modules.scala 56:109:@59161.4]
  wire [11:0] _T_104083; // @[Modules.scala 56:109:@59163.4]
  wire [10:0] _T_104084; // @[Modules.scala 56:109:@59164.4]
  wire [10:0] buffer_15_690; // @[Modules.scala 56:109:@59165.4]
  wire [11:0] _T_104086; // @[Modules.scala 56:109:@59167.4]
  wire [10:0] _T_104087; // @[Modules.scala 56:109:@59168.4]
  wire [10:0] buffer_15_691; // @[Modules.scala 56:109:@59169.4]
  wire [11:0] _T_104092; // @[Modules.scala 56:109:@59175.4]
  wire [10:0] _T_104093; // @[Modules.scala 56:109:@59176.4]
  wire [10:0] buffer_15_693; // @[Modules.scala 56:109:@59177.4]
  wire [11:0] _T_104095; // @[Modules.scala 56:109:@59179.4]
  wire [10:0] _T_104096; // @[Modules.scala 56:109:@59180.4]
  wire [10:0] buffer_15_694; // @[Modules.scala 56:109:@59181.4]
  wire [11:0] _T_104098; // @[Modules.scala 56:109:@59183.4]
  wire [10:0] _T_104099; // @[Modules.scala 56:109:@59184.4]
  wire [10:0] buffer_15_695; // @[Modules.scala 56:109:@59185.4]
  wire [11:0] _T_104101; // @[Modules.scala 56:109:@59187.4]
  wire [10:0] _T_104102; // @[Modules.scala 56:109:@59188.4]
  wire [10:0] buffer_15_696; // @[Modules.scala 56:109:@59189.4]
  wire [11:0] _T_104104; // @[Modules.scala 56:109:@59191.4]
  wire [10:0] _T_104105; // @[Modules.scala 56:109:@59192.4]
  wire [10:0] buffer_15_697; // @[Modules.scala 56:109:@59193.4]
  wire [11:0] _T_104107; // @[Modules.scala 56:109:@59195.4]
  wire [10:0] _T_104108; // @[Modules.scala 56:109:@59196.4]
  wire [10:0] buffer_15_698; // @[Modules.scala 56:109:@59197.4]
  wire [11:0] _T_104110; // @[Modules.scala 56:109:@59199.4]
  wire [10:0] _T_104111; // @[Modules.scala 56:109:@59200.4]
  wire [10:0] buffer_15_699; // @[Modules.scala 56:109:@59201.4]
  wire [11:0] _T_104113; // @[Modules.scala 56:109:@59203.4]
  wire [10:0] _T_104114; // @[Modules.scala 56:109:@59204.4]
  wire [10:0] buffer_15_700; // @[Modules.scala 56:109:@59205.4]
  wire [11:0] _T_104116; // @[Modules.scala 56:109:@59207.4]
  wire [10:0] _T_104117; // @[Modules.scala 56:109:@59208.4]
  wire [10:0] buffer_15_701; // @[Modules.scala 56:109:@59209.4]
  wire [11:0] _T_104119; // @[Modules.scala 56:109:@59211.4]
  wire [10:0] _T_104120; // @[Modules.scala 56:109:@59212.4]
  wire [10:0] buffer_15_702; // @[Modules.scala 56:109:@59213.4]
  wire [11:0] _T_104122; // @[Modules.scala 56:109:@59215.4]
  wire [10:0] _T_104123; // @[Modules.scala 56:109:@59216.4]
  wire [10:0] buffer_15_703; // @[Modules.scala 56:109:@59217.4]
  wire [11:0] _T_104125; // @[Modules.scala 56:109:@59219.4]
  wire [10:0] _T_104126; // @[Modules.scala 56:109:@59220.4]
  wire [10:0] buffer_15_704; // @[Modules.scala 56:109:@59221.4]
  wire [11:0] _T_104128; // @[Modules.scala 56:109:@59223.4]
  wire [10:0] _T_104129; // @[Modules.scala 56:109:@59224.4]
  wire [10:0] buffer_15_705; // @[Modules.scala 56:109:@59225.4]
  wire [11:0] _T_104131; // @[Modules.scala 56:109:@59227.4]
  wire [10:0] _T_104132; // @[Modules.scala 56:109:@59228.4]
  wire [10:0] buffer_15_706; // @[Modules.scala 56:109:@59229.4]
  wire [11:0] _T_104134; // @[Modules.scala 56:109:@59231.4]
  wire [10:0] _T_104135; // @[Modules.scala 56:109:@59232.4]
  wire [10:0] buffer_15_707; // @[Modules.scala 56:109:@59233.4]
  wire [11:0] _T_104137; // @[Modules.scala 56:109:@59235.4]
  wire [10:0] _T_104138; // @[Modules.scala 56:109:@59236.4]
  wire [10:0] buffer_15_708; // @[Modules.scala 56:109:@59237.4]
  wire [11:0] _T_104140; // @[Modules.scala 56:109:@59239.4]
  wire [10:0] _T_104141; // @[Modules.scala 56:109:@59240.4]
  wire [10:0] buffer_15_709; // @[Modules.scala 56:109:@59241.4]
  wire [11:0] _T_104143; // @[Modules.scala 56:109:@59243.4]
  wire [10:0] _T_104144; // @[Modules.scala 56:109:@59244.4]
  wire [10:0] buffer_15_710; // @[Modules.scala 56:109:@59245.4]
  wire [11:0] _T_104146; // @[Modules.scala 56:109:@59247.4]
  wire [10:0] _T_104147; // @[Modules.scala 56:109:@59248.4]
  wire [10:0] buffer_15_711; // @[Modules.scala 56:109:@59249.4]
  wire [11:0] _T_104149; // @[Modules.scala 56:109:@59251.4]
  wire [10:0] _T_104150; // @[Modules.scala 56:109:@59252.4]
  wire [10:0] buffer_15_712; // @[Modules.scala 56:109:@59253.4]
  wire [11:0] _T_104152; // @[Modules.scala 56:109:@59255.4]
  wire [10:0] _T_104153; // @[Modules.scala 56:109:@59256.4]
  wire [10:0] buffer_15_713; // @[Modules.scala 56:109:@59257.4]
  wire [11:0] _T_104155; // @[Modules.scala 56:109:@59259.4]
  wire [10:0] _T_104156; // @[Modules.scala 56:109:@59260.4]
  wire [10:0] buffer_15_714; // @[Modules.scala 56:109:@59261.4]
  wire [11:0] _T_104158; // @[Modules.scala 56:109:@59263.4]
  wire [10:0] _T_104159; // @[Modules.scala 56:109:@59264.4]
  wire [10:0] buffer_15_715; // @[Modules.scala 56:109:@59265.4]
  wire [11:0] _T_104161; // @[Modules.scala 56:109:@59267.4]
  wire [10:0] _T_104162; // @[Modules.scala 56:109:@59268.4]
  wire [10:0] buffer_15_716; // @[Modules.scala 56:109:@59269.4]
  wire [11:0] _T_104164; // @[Modules.scala 56:109:@59271.4]
  wire [10:0] _T_104165; // @[Modules.scala 56:109:@59272.4]
  wire [10:0] buffer_15_717; // @[Modules.scala 56:109:@59273.4]
  wire [11:0] _T_104167; // @[Modules.scala 56:109:@59275.4]
  wire [10:0] _T_104168; // @[Modules.scala 56:109:@59276.4]
  wire [10:0] buffer_15_718; // @[Modules.scala 56:109:@59277.4]
  wire [11:0] _T_104170; // @[Modules.scala 56:109:@59279.4]
  wire [10:0] _T_104171; // @[Modules.scala 56:109:@59280.4]
  wire [10:0] buffer_15_719; // @[Modules.scala 56:109:@59281.4]
  wire [11:0] _T_104173; // @[Modules.scala 56:109:@59283.4]
  wire [10:0] _T_104174; // @[Modules.scala 56:109:@59284.4]
  wire [10:0] buffer_15_720; // @[Modules.scala 56:109:@59285.4]
  wire [11:0] _T_104176; // @[Modules.scala 56:109:@59287.4]
  wire [10:0] _T_104177; // @[Modules.scala 56:109:@59288.4]
  wire [10:0] buffer_15_721; // @[Modules.scala 56:109:@59289.4]
  wire [11:0] _T_104179; // @[Modules.scala 56:109:@59291.4]
  wire [10:0] _T_104180; // @[Modules.scala 56:109:@59292.4]
  wire [10:0] buffer_15_722; // @[Modules.scala 56:109:@59293.4]
  wire [11:0] _T_104182; // @[Modules.scala 56:109:@59295.4]
  wire [10:0] _T_104183; // @[Modules.scala 56:109:@59296.4]
  wire [10:0] buffer_15_723; // @[Modules.scala 56:109:@59297.4]
  wire [11:0] _T_104185; // @[Modules.scala 56:109:@59299.4]
  wire [10:0] _T_104186; // @[Modules.scala 56:109:@59300.4]
  wire [10:0] buffer_15_724; // @[Modules.scala 56:109:@59301.4]
  wire [11:0] _T_104188; // @[Modules.scala 56:109:@59303.4]
  wire [10:0] _T_104189; // @[Modules.scala 56:109:@59304.4]
  wire [10:0] buffer_15_725; // @[Modules.scala 56:109:@59305.4]
  wire [11:0] _T_104191; // @[Modules.scala 56:109:@59307.4]
  wire [10:0] _T_104192; // @[Modules.scala 56:109:@59308.4]
  wire [10:0] buffer_15_726; // @[Modules.scala 56:109:@59309.4]
  wire [11:0] _T_104194; // @[Modules.scala 56:109:@59311.4]
  wire [10:0] _T_104195; // @[Modules.scala 56:109:@59312.4]
  wire [10:0] buffer_15_727; // @[Modules.scala 56:109:@59313.4]
  wire [11:0] _T_104197; // @[Modules.scala 56:109:@59315.4]
  wire [10:0] _T_104198; // @[Modules.scala 56:109:@59316.4]
  wire [10:0] buffer_15_728; // @[Modules.scala 56:109:@59317.4]
  wire [11:0] _T_104200; // @[Modules.scala 56:109:@59319.4]
  wire [10:0] _T_104201; // @[Modules.scala 56:109:@59320.4]
  wire [10:0] buffer_15_729; // @[Modules.scala 56:109:@59321.4]
  wire [11:0] _T_104203; // @[Modules.scala 56:109:@59323.4]
  wire [10:0] _T_104204; // @[Modules.scala 56:109:@59324.4]
  wire [10:0] buffer_15_730; // @[Modules.scala 56:109:@59325.4]
  wire [11:0] _T_104206; // @[Modules.scala 56:109:@59327.4]
  wire [10:0] _T_104207; // @[Modules.scala 56:109:@59328.4]
  wire [10:0] buffer_15_731; // @[Modules.scala 56:109:@59329.4]
  wire [11:0] _T_104209; // @[Modules.scala 56:109:@59331.4]
  wire [10:0] _T_104210; // @[Modules.scala 56:109:@59332.4]
  wire [10:0] buffer_15_732; // @[Modules.scala 56:109:@59333.4]
  wire [11:0] _T_104212; // @[Modules.scala 56:109:@59335.4]
  wire [10:0] _T_104213; // @[Modules.scala 56:109:@59336.4]
  wire [10:0] buffer_15_733; // @[Modules.scala 56:109:@59337.4]
  wire [11:0] _T_104215; // @[Modules.scala 56:109:@59339.4]
  wire [10:0] _T_104216; // @[Modules.scala 56:109:@59340.4]
  wire [10:0] buffer_15_734; // @[Modules.scala 56:109:@59341.4]
  wire [11:0] _T_104218; // @[Modules.scala 63:156:@59344.4]
  wire [10:0] _T_104219; // @[Modules.scala 63:156:@59345.4]
  wire [10:0] buffer_15_736; // @[Modules.scala 63:156:@59346.4]
  wire [11:0] _T_104221; // @[Modules.scala 63:156:@59348.4]
  wire [10:0] _T_104222; // @[Modules.scala 63:156:@59349.4]
  wire [10:0] buffer_15_737; // @[Modules.scala 63:156:@59350.4]
  wire [11:0] _T_104224; // @[Modules.scala 63:156:@59352.4]
  wire [10:0] _T_104225; // @[Modules.scala 63:156:@59353.4]
  wire [10:0] buffer_15_738; // @[Modules.scala 63:156:@59354.4]
  wire [11:0] _T_104227; // @[Modules.scala 63:156:@59356.4]
  wire [10:0] _T_104228; // @[Modules.scala 63:156:@59357.4]
  wire [10:0] buffer_15_739; // @[Modules.scala 63:156:@59358.4]
  wire [11:0] _T_104230; // @[Modules.scala 63:156:@59360.4]
  wire [10:0] _T_104231; // @[Modules.scala 63:156:@59361.4]
  wire [10:0] buffer_15_740; // @[Modules.scala 63:156:@59362.4]
  wire [11:0] _T_104233; // @[Modules.scala 63:156:@59364.4]
  wire [10:0] _T_104234; // @[Modules.scala 63:156:@59365.4]
  wire [10:0] buffer_15_741; // @[Modules.scala 63:156:@59366.4]
  wire [11:0] _T_104236; // @[Modules.scala 63:156:@59368.4]
  wire [10:0] _T_104237; // @[Modules.scala 63:156:@59369.4]
  wire [10:0] buffer_15_742; // @[Modules.scala 63:156:@59370.4]
  wire [11:0] _T_104239; // @[Modules.scala 63:156:@59372.4]
  wire [10:0] _T_104240; // @[Modules.scala 63:156:@59373.4]
  wire [10:0] buffer_15_743; // @[Modules.scala 63:156:@59374.4]
  wire [11:0] _T_104242; // @[Modules.scala 63:156:@59376.4]
  wire [10:0] _T_104243; // @[Modules.scala 63:156:@59377.4]
  wire [10:0] buffer_15_744; // @[Modules.scala 63:156:@59378.4]
  wire [11:0] _T_104245; // @[Modules.scala 63:156:@59380.4]
  wire [10:0] _T_104246; // @[Modules.scala 63:156:@59381.4]
  wire [10:0] buffer_15_745; // @[Modules.scala 63:156:@59382.4]
  wire [11:0] _T_104248; // @[Modules.scala 63:156:@59384.4]
  wire [10:0] _T_104249; // @[Modules.scala 63:156:@59385.4]
  wire [10:0] buffer_15_746; // @[Modules.scala 63:156:@59386.4]
  wire [11:0] _T_104251; // @[Modules.scala 63:156:@59388.4]
  wire [10:0] _T_104252; // @[Modules.scala 63:156:@59389.4]
  wire [10:0] buffer_15_747; // @[Modules.scala 63:156:@59390.4]
  wire [11:0] _T_104254; // @[Modules.scala 63:156:@59392.4]
  wire [10:0] _T_104255; // @[Modules.scala 63:156:@59393.4]
  wire [10:0] buffer_15_748; // @[Modules.scala 63:156:@59394.4]
  wire [11:0] _T_104257; // @[Modules.scala 63:156:@59396.4]
  wire [10:0] _T_104258; // @[Modules.scala 63:156:@59397.4]
  wire [10:0] buffer_15_749; // @[Modules.scala 63:156:@59398.4]
  wire [11:0] _T_104260; // @[Modules.scala 63:156:@59400.4]
  wire [10:0] _T_104261; // @[Modules.scala 63:156:@59401.4]
  wire [10:0] buffer_15_750; // @[Modules.scala 63:156:@59402.4]
  wire [11:0] _T_104263; // @[Modules.scala 63:156:@59404.4]
  wire [10:0] _T_104264; // @[Modules.scala 63:156:@59405.4]
  wire [10:0] buffer_15_751; // @[Modules.scala 63:156:@59406.4]
  wire [11:0] _T_104266; // @[Modules.scala 63:156:@59408.4]
  wire [10:0] _T_104267; // @[Modules.scala 63:156:@59409.4]
  wire [10:0] buffer_15_752; // @[Modules.scala 63:156:@59410.4]
  wire [11:0] _T_104269; // @[Modules.scala 63:156:@59412.4]
  wire [10:0] _T_104270; // @[Modules.scala 63:156:@59413.4]
  wire [10:0] buffer_15_753; // @[Modules.scala 63:156:@59414.4]
  wire [11:0] _T_104272; // @[Modules.scala 63:156:@59416.4]
  wire [10:0] _T_104273; // @[Modules.scala 63:156:@59417.4]
  wire [10:0] buffer_15_754; // @[Modules.scala 63:156:@59418.4]
  wire [11:0] _T_104275; // @[Modules.scala 63:156:@59420.4]
  wire [10:0] _T_104276; // @[Modules.scala 63:156:@59421.4]
  wire [10:0] buffer_15_755; // @[Modules.scala 63:156:@59422.4]
  wire [11:0] _T_104278; // @[Modules.scala 63:156:@59424.4]
  wire [10:0] _T_104279; // @[Modules.scala 63:156:@59425.4]
  wire [10:0] buffer_15_756; // @[Modules.scala 63:156:@59426.4]
  wire [11:0] _T_104281; // @[Modules.scala 63:156:@59428.4]
  wire [10:0] _T_104282; // @[Modules.scala 63:156:@59429.4]
  wire [10:0] buffer_15_757; // @[Modules.scala 63:156:@59430.4]
  wire [11:0] _T_104284; // @[Modules.scala 63:156:@59432.4]
  wire [10:0] _T_104285; // @[Modules.scala 63:156:@59433.4]
  wire [10:0] buffer_15_758; // @[Modules.scala 63:156:@59434.4]
  wire [11:0] _T_104287; // @[Modules.scala 63:156:@59436.4]
  wire [10:0] _T_104288; // @[Modules.scala 63:156:@59437.4]
  wire [10:0] buffer_15_759; // @[Modules.scala 63:156:@59438.4]
  wire [11:0] _T_104290; // @[Modules.scala 63:156:@59440.4]
  wire [10:0] _T_104291; // @[Modules.scala 63:156:@59441.4]
  wire [10:0] buffer_15_760; // @[Modules.scala 63:156:@59442.4]
  wire [11:0] _T_104293; // @[Modules.scala 63:156:@59444.4]
  wire [10:0] _T_104294; // @[Modules.scala 63:156:@59445.4]
  wire [10:0] buffer_15_761; // @[Modules.scala 63:156:@59446.4]
  wire [11:0] _T_104296; // @[Modules.scala 63:156:@59448.4]
  wire [10:0] _T_104297; // @[Modules.scala 63:156:@59449.4]
  wire [10:0] buffer_15_762; // @[Modules.scala 63:156:@59450.4]
  wire [11:0] _T_104299; // @[Modules.scala 63:156:@59452.4]
  wire [10:0] _T_104300; // @[Modules.scala 63:156:@59453.4]
  wire [10:0] buffer_15_763; // @[Modules.scala 63:156:@59454.4]
  wire [11:0] _T_104302; // @[Modules.scala 63:156:@59456.4]
  wire [10:0] _T_104303; // @[Modules.scala 63:156:@59457.4]
  wire [10:0] buffer_15_764; // @[Modules.scala 63:156:@59458.4]
  wire [11:0] _T_104305; // @[Modules.scala 63:156:@59460.4]
  wire [10:0] _T_104306; // @[Modules.scala 63:156:@59461.4]
  wire [10:0] buffer_15_765; // @[Modules.scala 63:156:@59462.4]
  wire [11:0] _T_104308; // @[Modules.scala 63:156:@59464.4]
  wire [10:0] _T_104309; // @[Modules.scala 63:156:@59465.4]
  wire [10:0] buffer_15_766; // @[Modules.scala 63:156:@59466.4]
  wire [11:0] _T_104311; // @[Modules.scala 63:156:@59468.4]
  wire [10:0] _T_104312; // @[Modules.scala 63:156:@59469.4]
  wire [10:0] buffer_15_767; // @[Modules.scala 63:156:@59470.4]
  wire [11:0] _T_104314; // @[Modules.scala 63:156:@59472.4]
  wire [10:0] _T_104315; // @[Modules.scala 63:156:@59473.4]
  wire [10:0] buffer_15_768; // @[Modules.scala 63:156:@59474.4]
  wire [11:0] _T_104317; // @[Modules.scala 63:156:@59476.4]
  wire [10:0] _T_104318; // @[Modules.scala 63:156:@59477.4]
  wire [10:0] buffer_15_769; // @[Modules.scala 63:156:@59478.4]
  wire [11:0] _T_104320; // @[Modules.scala 63:156:@59480.4]
  wire [10:0] _T_104321; // @[Modules.scala 63:156:@59481.4]
  wire [10:0] buffer_15_770; // @[Modules.scala 63:156:@59482.4]
  wire [11:0] _T_104323; // @[Modules.scala 63:156:@59484.4]
  wire [10:0] _T_104324; // @[Modules.scala 63:156:@59485.4]
  wire [10:0] buffer_15_771; // @[Modules.scala 63:156:@59486.4]
  wire [11:0] _T_104326; // @[Modules.scala 63:156:@59488.4]
  wire [10:0] _T_104327; // @[Modules.scala 63:156:@59489.4]
  wire [10:0] buffer_15_772; // @[Modules.scala 63:156:@59490.4]
  wire [11:0] _T_104329; // @[Modules.scala 63:156:@59492.4]
  wire [10:0] _T_104330; // @[Modules.scala 63:156:@59493.4]
  wire [10:0] buffer_15_773; // @[Modules.scala 63:156:@59494.4]
  wire [11:0] _T_104332; // @[Modules.scala 63:156:@59496.4]
  wire [10:0] _T_104333; // @[Modules.scala 63:156:@59497.4]
  wire [10:0] buffer_15_774; // @[Modules.scala 63:156:@59498.4]
  wire [11:0] _T_104335; // @[Modules.scala 63:156:@59500.4]
  wire [10:0] _T_104336; // @[Modules.scala 63:156:@59501.4]
  wire [10:0] buffer_15_775; // @[Modules.scala 63:156:@59502.4]
  wire [11:0] _T_104338; // @[Modules.scala 63:156:@59504.4]
  wire [10:0] _T_104339; // @[Modules.scala 63:156:@59505.4]
  wire [10:0] buffer_15_776; // @[Modules.scala 63:156:@59506.4]
  wire [11:0] _T_104341; // @[Modules.scala 63:156:@59508.4]
  wire [10:0] _T_104342; // @[Modules.scala 63:156:@59509.4]
  wire [10:0] buffer_15_777; // @[Modules.scala 63:156:@59510.4]
  wire [11:0] _T_104344; // @[Modules.scala 63:156:@59512.4]
  wire [10:0] _T_104345; // @[Modules.scala 63:156:@59513.4]
  wire [10:0] buffer_15_778; // @[Modules.scala 63:156:@59514.4]
  wire [11:0] _T_104347; // @[Modules.scala 63:156:@59516.4]
  wire [10:0] _T_104348; // @[Modules.scala 63:156:@59517.4]
  wire [10:0] buffer_15_779; // @[Modules.scala 63:156:@59518.4]
  wire [11:0] _T_104350; // @[Modules.scala 63:156:@59520.4]
  wire [10:0] _T_104351; // @[Modules.scala 63:156:@59521.4]
  wire [10:0] buffer_15_780; // @[Modules.scala 63:156:@59522.4]
  wire [11:0] _T_104353; // @[Modules.scala 63:156:@59524.4]
  wire [10:0] _T_104354; // @[Modules.scala 63:156:@59525.4]
  wire [10:0] buffer_15_781; // @[Modules.scala 63:156:@59526.4]
  wire [11:0] _T_104356; // @[Modules.scala 63:156:@59528.4]
  wire [10:0] _T_104357; // @[Modules.scala 63:156:@59529.4]
  wire [10:0] buffer_15_782; // @[Modules.scala 63:156:@59530.4]
  wire [11:0] _T_104359; // @[Modules.scala 63:156:@59532.4]
  wire [10:0] _T_104360; // @[Modules.scala 63:156:@59533.4]
  wire [10:0] buffer_15_783; // @[Modules.scala 63:156:@59534.4]
  assign _T_54267 = $signed(5'sh0) - $signed(io_in_0); // @[Modules.scala 43:37:@9.4]
  assign _T_54268 = _T_54267[4:0]; // @[Modules.scala 43:37:@10.4]
  assign _T_54269 = $signed(_T_54268); // @[Modules.scala 43:37:@11.4]
  assign _T_54270 = $signed(_T_54269) + $signed(io_in_1); // @[Modules.scala 43:47:@12.4]
  assign _T_54271 = _T_54270[4:0]; // @[Modules.scala 43:47:@13.4]
  assign _T_54272 = $signed(_T_54271); // @[Modules.scala 43:47:@14.4]
  assign _T_54274 = $signed(5'sh0) - $signed(io_in_2); // @[Modules.scala 46:37:@16.4]
  assign _T_54275 = _T_54274[4:0]; // @[Modules.scala 46:37:@17.4]
  assign _T_54276 = $signed(_T_54275); // @[Modules.scala 46:37:@18.4]
  assign _T_54277 = $signed(_T_54276) - $signed(io_in_3); // @[Modules.scala 46:47:@19.4]
  assign _T_54278 = _T_54277[4:0]; // @[Modules.scala 46:47:@20.4]
  assign _T_54279 = $signed(_T_54278); // @[Modules.scala 46:47:@21.4]
  assign _T_54281 = $signed(5'sh0) - $signed(io_in_4); // @[Modules.scala 43:37:@23.4]
  assign _T_54282 = _T_54281[4:0]; // @[Modules.scala 43:37:@24.4]
  assign _T_54283 = $signed(_T_54282); // @[Modules.scala 43:37:@25.4]
  assign _T_54284 = $signed(_T_54283) + $signed(io_in_5); // @[Modules.scala 43:47:@26.4]
  assign _T_54285 = _T_54284[4:0]; // @[Modules.scala 43:47:@27.4]
  assign _T_54286 = $signed(_T_54285); // @[Modules.scala 43:47:@28.4]
  assign _T_54288 = $signed(5'sh0) - $signed(io_in_6); // @[Modules.scala 43:37:@30.4]
  assign _T_54289 = _T_54288[4:0]; // @[Modules.scala 43:37:@31.4]
  assign _T_54290 = $signed(_T_54289); // @[Modules.scala 43:37:@32.4]
  assign _T_54291 = $signed(_T_54290) + $signed(io_in_7); // @[Modules.scala 43:47:@33.4]
  assign _T_54292 = _T_54291[4:0]; // @[Modules.scala 43:47:@34.4]
  assign _T_54293 = $signed(_T_54292); // @[Modules.scala 43:47:@35.4]
  assign _T_54295 = $signed(5'sh0) - $signed(io_in_8); // @[Modules.scala 43:37:@37.4]
  assign _T_54296 = _T_54295[4:0]; // @[Modules.scala 43:37:@38.4]
  assign _T_54297 = $signed(_T_54296); // @[Modules.scala 43:37:@39.4]
  assign _T_54298 = $signed(_T_54297) + $signed(io_in_9); // @[Modules.scala 43:47:@40.4]
  assign _T_54299 = _T_54298[4:0]; // @[Modules.scala 43:47:@41.4]
  assign _T_54300 = $signed(_T_54299); // @[Modules.scala 43:47:@42.4]
  assign _T_54302 = $signed(5'sh0) - $signed(io_in_10); // @[Modules.scala 46:37:@44.4]
  assign _T_54303 = _T_54302[4:0]; // @[Modules.scala 46:37:@45.4]
  assign _T_54304 = $signed(_T_54303); // @[Modules.scala 46:37:@46.4]
  assign _T_54305 = $signed(_T_54304) - $signed(io_in_11); // @[Modules.scala 46:47:@47.4]
  assign _T_54306 = _T_54305[4:0]; // @[Modules.scala 46:47:@48.4]
  assign _T_54307 = $signed(_T_54306); // @[Modules.scala 46:47:@49.4]
  assign _T_54309 = $signed(5'sh0) - $signed(io_in_12); // @[Modules.scala 46:37:@51.4]
  assign _T_54310 = _T_54309[4:0]; // @[Modules.scala 46:37:@52.4]
  assign _T_54311 = $signed(_T_54310); // @[Modules.scala 46:37:@53.4]
  assign _T_54312 = $signed(_T_54311) - $signed(io_in_13); // @[Modules.scala 46:47:@54.4]
  assign _T_54313 = _T_54312[4:0]; // @[Modules.scala 46:47:@55.4]
  assign _T_54314 = $signed(_T_54313); // @[Modules.scala 46:47:@56.4]
  assign _T_54316 = $signed(5'sh0) - $signed(io_in_14); // @[Modules.scala 46:37:@58.4]
  assign _T_54317 = _T_54316[4:0]; // @[Modules.scala 46:37:@59.4]
  assign _T_54318 = $signed(_T_54317); // @[Modules.scala 46:37:@60.4]
  assign _T_54319 = $signed(_T_54318) - $signed(io_in_15); // @[Modules.scala 46:47:@61.4]
  assign _T_54320 = _T_54319[4:0]; // @[Modules.scala 46:47:@62.4]
  assign _T_54321 = $signed(_T_54320); // @[Modules.scala 46:47:@63.4]
  assign _T_54322 = $signed(io_in_16) + $signed(io_in_17); // @[Modules.scala 37:46:@65.4]
  assign _T_54323 = _T_54322[4:0]; // @[Modules.scala 37:46:@66.4]
  assign _T_54324 = $signed(_T_54323); // @[Modules.scala 37:46:@67.4]
  assign _T_54326 = $signed(5'sh0) - $signed(io_in_18); // @[Modules.scala 46:37:@69.4]
  assign _T_54327 = _T_54326[4:0]; // @[Modules.scala 46:37:@70.4]
  assign _T_54328 = $signed(_T_54327); // @[Modules.scala 46:37:@71.4]
  assign _T_54329 = $signed(_T_54328) - $signed(io_in_19); // @[Modules.scala 46:47:@72.4]
  assign _T_54330 = _T_54329[4:0]; // @[Modules.scala 46:47:@73.4]
  assign _T_54331 = $signed(_T_54330); // @[Modules.scala 46:47:@74.4]
  assign _T_54332 = $signed(io_in_20) + $signed(io_in_21); // @[Modules.scala 37:46:@76.4]
  assign _T_54333 = _T_54332[4:0]; // @[Modules.scala 37:46:@77.4]
  assign _T_54334 = $signed(_T_54333); // @[Modules.scala 37:46:@78.4]
  assign _T_54336 = $signed(5'sh0) - $signed(io_in_22); // @[Modules.scala 43:37:@80.4]
  assign _T_54337 = _T_54336[4:0]; // @[Modules.scala 43:37:@81.4]
  assign _T_54338 = $signed(_T_54337); // @[Modules.scala 43:37:@82.4]
  assign _T_54339 = $signed(_T_54338) + $signed(io_in_23); // @[Modules.scala 43:47:@83.4]
  assign _T_54340 = _T_54339[4:0]; // @[Modules.scala 43:47:@84.4]
  assign _T_54341 = $signed(_T_54340); // @[Modules.scala 43:47:@85.4]
  assign _T_54343 = $signed(5'sh0) - $signed(io_in_24); // @[Modules.scala 43:37:@87.4]
  assign _T_54344 = _T_54343[4:0]; // @[Modules.scala 43:37:@88.4]
  assign _T_54345 = $signed(_T_54344); // @[Modules.scala 43:37:@89.4]
  assign _T_54346 = $signed(_T_54345) + $signed(io_in_25); // @[Modules.scala 43:47:@90.4]
  assign _T_54347 = _T_54346[4:0]; // @[Modules.scala 43:47:@91.4]
  assign _T_54348 = $signed(_T_54347); // @[Modules.scala 43:47:@92.4]
  assign _T_54349 = $signed(io_in_26) - $signed(io_in_27); // @[Modules.scala 40:46:@94.4]
  assign _T_54350 = _T_54349[4:0]; // @[Modules.scala 40:46:@95.4]
  assign _T_54351 = $signed(_T_54350); // @[Modules.scala 40:46:@96.4]
  assign _T_54353 = $signed(5'sh0) - $signed(io_in_28); // @[Modules.scala 46:37:@98.4]
  assign _T_54354 = _T_54353[4:0]; // @[Modules.scala 46:37:@99.4]
  assign _T_54355 = $signed(_T_54354); // @[Modules.scala 46:37:@100.4]
  assign _T_54356 = $signed(_T_54355) - $signed(io_in_29); // @[Modules.scala 46:47:@101.4]
  assign _T_54357 = _T_54356[4:0]; // @[Modules.scala 46:47:@102.4]
  assign _T_54358 = $signed(_T_54357); // @[Modules.scala 46:47:@103.4]
  assign _T_54360 = $signed(5'sh0) - $signed(io_in_30); // @[Modules.scala 43:37:@105.4]
  assign _T_54361 = _T_54360[4:0]; // @[Modules.scala 43:37:@106.4]
  assign _T_54362 = $signed(_T_54361); // @[Modules.scala 43:37:@107.4]
  assign _T_54363 = $signed(_T_54362) + $signed(io_in_31); // @[Modules.scala 43:47:@108.4]
  assign _T_54364 = _T_54363[4:0]; // @[Modules.scala 43:47:@109.4]
  assign _T_54365 = $signed(_T_54364); // @[Modules.scala 43:47:@110.4]
  assign _T_54366 = $signed(io_in_32) + $signed(io_in_33); // @[Modules.scala 37:46:@112.4]
  assign _T_54367 = _T_54366[4:0]; // @[Modules.scala 37:46:@113.4]
  assign _T_54368 = $signed(_T_54367); // @[Modules.scala 37:46:@114.4]
  assign _T_54370 = $signed(5'sh0) - $signed(io_in_34); // @[Modules.scala 46:37:@116.4]
  assign _T_54371 = _T_54370[4:0]; // @[Modules.scala 46:37:@117.4]
  assign _T_54372 = $signed(_T_54371); // @[Modules.scala 46:37:@118.4]
  assign _T_54373 = $signed(_T_54372) - $signed(io_in_35); // @[Modules.scala 46:47:@119.4]
  assign _T_54374 = _T_54373[4:0]; // @[Modules.scala 46:47:@120.4]
  assign _T_54375 = $signed(_T_54374); // @[Modules.scala 46:47:@121.4]
  assign _T_54377 = $signed(5'sh0) - $signed(io_in_36); // @[Modules.scala 46:37:@123.4]
  assign _T_54378 = _T_54377[4:0]; // @[Modules.scala 46:37:@124.4]
  assign _T_54379 = $signed(_T_54378); // @[Modules.scala 46:37:@125.4]
  assign _T_54380 = $signed(_T_54379) - $signed(io_in_37); // @[Modules.scala 46:47:@126.4]
  assign _T_54381 = _T_54380[4:0]; // @[Modules.scala 46:47:@127.4]
  assign _T_54382 = $signed(_T_54381); // @[Modules.scala 46:47:@128.4]
  assign _T_54384 = $signed(5'sh0) - $signed(io_in_38); // @[Modules.scala 46:37:@130.4]
  assign _T_54385 = _T_54384[4:0]; // @[Modules.scala 46:37:@131.4]
  assign _T_54386 = $signed(_T_54385); // @[Modules.scala 46:37:@132.4]
  assign _T_54387 = $signed(_T_54386) - $signed(io_in_39); // @[Modules.scala 46:47:@133.4]
  assign _T_54388 = _T_54387[4:0]; // @[Modules.scala 46:47:@134.4]
  assign _T_54389 = $signed(_T_54388); // @[Modules.scala 46:47:@135.4]
  assign _T_54391 = $signed(5'sh0) - $signed(io_in_40); // @[Modules.scala 46:37:@137.4]
  assign _T_54392 = _T_54391[4:0]; // @[Modules.scala 46:37:@138.4]
  assign _T_54393 = $signed(_T_54392); // @[Modules.scala 46:37:@139.4]
  assign _T_54394 = $signed(_T_54393) - $signed(io_in_41); // @[Modules.scala 46:47:@140.4]
  assign _T_54395 = _T_54394[4:0]; // @[Modules.scala 46:47:@141.4]
  assign _T_54396 = $signed(_T_54395); // @[Modules.scala 46:47:@142.4]
  assign _T_54398 = $signed(5'sh0) - $signed(io_in_42); // @[Modules.scala 46:37:@144.4]
  assign _T_54399 = _T_54398[4:0]; // @[Modules.scala 46:37:@145.4]
  assign _T_54400 = $signed(_T_54399); // @[Modules.scala 46:37:@146.4]
  assign _T_54401 = $signed(_T_54400) - $signed(io_in_43); // @[Modules.scala 46:47:@147.4]
  assign _T_54402 = _T_54401[4:0]; // @[Modules.scala 46:47:@148.4]
  assign _T_54403 = $signed(_T_54402); // @[Modules.scala 46:47:@149.4]
  assign _T_54405 = $signed(5'sh0) - $signed(io_in_44); // @[Modules.scala 46:37:@151.4]
  assign _T_54406 = _T_54405[4:0]; // @[Modules.scala 46:37:@152.4]
  assign _T_54407 = $signed(_T_54406); // @[Modules.scala 46:37:@153.4]
  assign _T_54408 = $signed(_T_54407) - $signed(io_in_45); // @[Modules.scala 46:47:@154.4]
  assign _T_54409 = _T_54408[4:0]; // @[Modules.scala 46:47:@155.4]
  assign _T_54410 = $signed(_T_54409); // @[Modules.scala 46:47:@156.4]
  assign _T_54412 = $signed(5'sh0) - $signed(io_in_46); // @[Modules.scala 46:37:@158.4]
  assign _T_54413 = _T_54412[4:0]; // @[Modules.scala 46:37:@159.4]
  assign _T_54414 = $signed(_T_54413); // @[Modules.scala 46:37:@160.4]
  assign _T_54415 = $signed(_T_54414) - $signed(io_in_47); // @[Modules.scala 46:47:@161.4]
  assign _T_54416 = _T_54415[4:0]; // @[Modules.scala 46:47:@162.4]
  assign _T_54417 = $signed(_T_54416); // @[Modules.scala 46:47:@163.4]
  assign _T_54419 = $signed(5'sh0) - $signed(io_in_48); // @[Modules.scala 46:37:@165.4]
  assign _T_54420 = _T_54419[4:0]; // @[Modules.scala 46:37:@166.4]
  assign _T_54421 = $signed(_T_54420); // @[Modules.scala 46:37:@167.4]
  assign _T_54422 = $signed(_T_54421) - $signed(io_in_49); // @[Modules.scala 46:47:@168.4]
  assign _T_54423 = _T_54422[4:0]; // @[Modules.scala 46:47:@169.4]
  assign _T_54424 = $signed(_T_54423); // @[Modules.scala 46:47:@170.4]
  assign _T_54426 = $signed(5'sh0) - $signed(io_in_50); // @[Modules.scala 46:37:@172.4]
  assign _T_54427 = _T_54426[4:0]; // @[Modules.scala 46:37:@173.4]
  assign _T_54428 = $signed(_T_54427); // @[Modules.scala 46:37:@174.4]
  assign _T_54429 = $signed(_T_54428) - $signed(io_in_51); // @[Modules.scala 46:47:@175.4]
  assign _T_54430 = _T_54429[4:0]; // @[Modules.scala 46:47:@176.4]
  assign _T_54431 = $signed(_T_54430); // @[Modules.scala 46:47:@177.4]
  assign _T_54432 = $signed(io_in_52) + $signed(io_in_53); // @[Modules.scala 37:46:@179.4]
  assign _T_54433 = _T_54432[4:0]; // @[Modules.scala 37:46:@180.4]
  assign _T_54434 = $signed(_T_54433); // @[Modules.scala 37:46:@181.4]
  assign _T_54435 = $signed(io_in_54) - $signed(io_in_55); // @[Modules.scala 40:46:@183.4]
  assign _T_54436 = _T_54435[4:0]; // @[Modules.scala 40:46:@184.4]
  assign _T_54437 = $signed(_T_54436); // @[Modules.scala 40:46:@185.4]
  assign _T_54438 = $signed(io_in_56) - $signed(io_in_57); // @[Modules.scala 40:46:@187.4]
  assign _T_54439 = _T_54438[4:0]; // @[Modules.scala 40:46:@188.4]
  assign _T_54440 = $signed(_T_54439); // @[Modules.scala 40:46:@189.4]
  assign _T_54442 = $signed(5'sh0) - $signed(io_in_58); // @[Modules.scala 46:37:@191.4]
  assign _T_54443 = _T_54442[4:0]; // @[Modules.scala 46:37:@192.4]
  assign _T_54444 = $signed(_T_54443); // @[Modules.scala 46:37:@193.4]
  assign _T_54445 = $signed(_T_54444) - $signed(io_in_59); // @[Modules.scala 46:47:@194.4]
  assign _T_54446 = _T_54445[4:0]; // @[Modules.scala 46:47:@195.4]
  assign _T_54447 = $signed(_T_54446); // @[Modules.scala 46:47:@196.4]
  assign _T_54449 = $signed(5'sh0) - $signed(io_in_60); // @[Modules.scala 46:37:@198.4]
  assign _T_54450 = _T_54449[4:0]; // @[Modules.scala 46:37:@199.4]
  assign _T_54451 = $signed(_T_54450); // @[Modules.scala 46:37:@200.4]
  assign _T_54452 = $signed(_T_54451) - $signed(io_in_61); // @[Modules.scala 46:47:@201.4]
  assign _T_54453 = _T_54452[4:0]; // @[Modules.scala 46:47:@202.4]
  assign _T_54454 = $signed(_T_54453); // @[Modules.scala 46:47:@203.4]
  assign _T_54456 = $signed(5'sh0) - $signed(io_in_62); // @[Modules.scala 46:37:@205.4]
  assign _T_54457 = _T_54456[4:0]; // @[Modules.scala 46:37:@206.4]
  assign _T_54458 = $signed(_T_54457); // @[Modules.scala 46:37:@207.4]
  assign _T_54459 = $signed(_T_54458) - $signed(io_in_63); // @[Modules.scala 46:47:@208.4]
  assign _T_54460 = _T_54459[4:0]; // @[Modules.scala 46:47:@209.4]
  assign _T_54461 = $signed(_T_54460); // @[Modules.scala 46:47:@210.4]
  assign _T_54463 = $signed(5'sh0) - $signed(io_in_64); // @[Modules.scala 43:37:@212.4]
  assign _T_54464 = _T_54463[4:0]; // @[Modules.scala 43:37:@213.4]
  assign _T_54465 = $signed(_T_54464); // @[Modules.scala 43:37:@214.4]
  assign _T_54466 = $signed(_T_54465) + $signed(io_in_65); // @[Modules.scala 43:47:@215.4]
  assign _T_54467 = _T_54466[4:0]; // @[Modules.scala 43:47:@216.4]
  assign _T_54468 = $signed(_T_54467); // @[Modules.scala 43:47:@217.4]
  assign _T_54470 = $signed(5'sh0) - $signed(io_in_66); // @[Modules.scala 46:37:@219.4]
  assign _T_54471 = _T_54470[4:0]; // @[Modules.scala 46:37:@220.4]
  assign _T_54472 = $signed(_T_54471); // @[Modules.scala 46:37:@221.4]
  assign _T_54473 = $signed(_T_54472) - $signed(io_in_67); // @[Modules.scala 46:47:@222.4]
  assign _T_54474 = _T_54473[4:0]; // @[Modules.scala 46:47:@223.4]
  assign _T_54475 = $signed(_T_54474); // @[Modules.scala 46:47:@224.4]
  assign _T_54477 = $signed(5'sh0) - $signed(io_in_68); // @[Modules.scala 46:37:@226.4]
  assign _T_54478 = _T_54477[4:0]; // @[Modules.scala 46:37:@227.4]
  assign _T_54479 = $signed(_T_54478); // @[Modules.scala 46:37:@228.4]
  assign _T_54480 = $signed(_T_54479) - $signed(io_in_69); // @[Modules.scala 46:47:@229.4]
  assign _T_54481 = _T_54480[4:0]; // @[Modules.scala 46:47:@230.4]
  assign _T_54482 = $signed(_T_54481); // @[Modules.scala 46:47:@231.4]
  assign _T_54484 = $signed(5'sh0) - $signed(io_in_70); // @[Modules.scala 46:37:@233.4]
  assign _T_54485 = _T_54484[4:0]; // @[Modules.scala 46:37:@234.4]
  assign _T_54486 = $signed(_T_54485); // @[Modules.scala 46:37:@235.4]
  assign _T_54487 = $signed(_T_54486) - $signed(io_in_71); // @[Modules.scala 46:47:@236.4]
  assign _T_54488 = _T_54487[4:0]; // @[Modules.scala 46:47:@237.4]
  assign _T_54489 = $signed(_T_54488); // @[Modules.scala 46:47:@238.4]
  assign _T_54491 = $signed(5'sh0) - $signed(io_in_72); // @[Modules.scala 46:37:@240.4]
  assign _T_54492 = _T_54491[4:0]; // @[Modules.scala 46:37:@241.4]
  assign _T_54493 = $signed(_T_54492); // @[Modules.scala 46:37:@242.4]
  assign _T_54494 = $signed(_T_54493) - $signed(io_in_73); // @[Modules.scala 46:47:@243.4]
  assign _T_54495 = _T_54494[4:0]; // @[Modules.scala 46:47:@244.4]
  assign _T_54496 = $signed(_T_54495); // @[Modules.scala 46:47:@245.4]
  assign _T_54498 = $signed(5'sh0) - $signed(io_in_74); // @[Modules.scala 43:37:@247.4]
  assign _T_54499 = _T_54498[4:0]; // @[Modules.scala 43:37:@248.4]
  assign _T_54500 = $signed(_T_54499); // @[Modules.scala 43:37:@249.4]
  assign _T_54501 = $signed(_T_54500) + $signed(io_in_75); // @[Modules.scala 43:47:@250.4]
  assign _T_54502 = _T_54501[4:0]; // @[Modules.scala 43:47:@251.4]
  assign _T_54503 = $signed(_T_54502); // @[Modules.scala 43:47:@252.4]
  assign _T_54504 = $signed(io_in_76) - $signed(io_in_77); // @[Modules.scala 40:46:@254.4]
  assign _T_54505 = _T_54504[4:0]; // @[Modules.scala 40:46:@255.4]
  assign _T_54506 = $signed(_T_54505); // @[Modules.scala 40:46:@256.4]
  assign _T_54507 = $signed(io_in_78) + $signed(io_in_79); // @[Modules.scala 37:46:@258.4]
  assign _T_54508 = _T_54507[4:0]; // @[Modules.scala 37:46:@259.4]
  assign _T_54509 = $signed(_T_54508); // @[Modules.scala 37:46:@260.4]
  assign _T_54511 = $signed(5'sh0) - $signed(io_in_80); // @[Modules.scala 46:37:@262.4]
  assign _T_54512 = _T_54511[4:0]; // @[Modules.scala 46:37:@263.4]
  assign _T_54513 = $signed(_T_54512); // @[Modules.scala 46:37:@264.4]
  assign _T_54514 = $signed(_T_54513) - $signed(io_in_81); // @[Modules.scala 46:47:@265.4]
  assign _T_54515 = _T_54514[4:0]; // @[Modules.scala 46:47:@266.4]
  assign _T_54516 = $signed(_T_54515); // @[Modules.scala 46:47:@267.4]
  assign _T_54517 = $signed(io_in_82) - $signed(io_in_83); // @[Modules.scala 40:46:@269.4]
  assign _T_54518 = _T_54517[4:0]; // @[Modules.scala 40:46:@270.4]
  assign _T_54519 = $signed(_T_54518); // @[Modules.scala 40:46:@271.4]
  assign _T_54520 = $signed(io_in_84) - $signed(io_in_85); // @[Modules.scala 40:46:@273.4]
  assign _T_54521 = _T_54520[4:0]; // @[Modules.scala 40:46:@274.4]
  assign _T_54522 = $signed(_T_54521); // @[Modules.scala 40:46:@275.4]
  assign _T_54524 = $signed(5'sh0) - $signed(io_in_86); // @[Modules.scala 46:37:@277.4]
  assign _T_54525 = _T_54524[4:0]; // @[Modules.scala 46:37:@278.4]
  assign _T_54526 = $signed(_T_54525); // @[Modules.scala 46:37:@279.4]
  assign _T_54527 = $signed(_T_54526) - $signed(io_in_87); // @[Modules.scala 46:47:@280.4]
  assign _T_54528 = _T_54527[4:0]; // @[Modules.scala 46:47:@281.4]
  assign _T_54529 = $signed(_T_54528); // @[Modules.scala 46:47:@282.4]
  assign _T_54530 = $signed(io_in_88) + $signed(io_in_89); // @[Modules.scala 37:46:@284.4]
  assign _T_54531 = _T_54530[4:0]; // @[Modules.scala 37:46:@285.4]
  assign _T_54532 = $signed(_T_54531); // @[Modules.scala 37:46:@286.4]
  assign _T_54533 = $signed(io_in_90) + $signed(io_in_91); // @[Modules.scala 37:46:@288.4]
  assign _T_54534 = _T_54533[4:0]; // @[Modules.scala 37:46:@289.4]
  assign _T_54535 = $signed(_T_54534); // @[Modules.scala 37:46:@290.4]
  assign _T_54537 = $signed(5'sh0) - $signed(io_in_92); // @[Modules.scala 43:37:@292.4]
  assign _T_54538 = _T_54537[4:0]; // @[Modules.scala 43:37:@293.4]
  assign _T_54539 = $signed(_T_54538); // @[Modules.scala 43:37:@294.4]
  assign _T_54540 = $signed(_T_54539) + $signed(io_in_93); // @[Modules.scala 43:47:@295.4]
  assign _T_54541 = _T_54540[4:0]; // @[Modules.scala 43:47:@296.4]
  assign _T_54542 = $signed(_T_54541); // @[Modules.scala 43:47:@297.4]
  assign _T_54543 = $signed(io_in_94) + $signed(io_in_95); // @[Modules.scala 37:46:@299.4]
  assign _T_54544 = _T_54543[4:0]; // @[Modules.scala 37:46:@300.4]
  assign _T_54545 = $signed(_T_54544); // @[Modules.scala 37:46:@301.4]
  assign _T_54547 = $signed(5'sh0) - $signed(io_in_96); // @[Modules.scala 43:37:@303.4]
  assign _T_54548 = _T_54547[4:0]; // @[Modules.scala 43:37:@304.4]
  assign _T_54549 = $signed(_T_54548); // @[Modules.scala 43:37:@305.4]
  assign _T_54550 = $signed(_T_54549) + $signed(io_in_97); // @[Modules.scala 43:47:@306.4]
  assign _T_54551 = _T_54550[4:0]; // @[Modules.scala 43:47:@307.4]
  assign _T_54552 = $signed(_T_54551); // @[Modules.scala 43:47:@308.4]
  assign _T_54553 = $signed(io_in_98) + $signed(io_in_99); // @[Modules.scala 37:46:@310.4]
  assign _T_54554 = _T_54553[4:0]; // @[Modules.scala 37:46:@311.4]
  assign _T_54555 = $signed(_T_54554); // @[Modules.scala 37:46:@312.4]
  assign _T_54556 = $signed(io_in_100) + $signed(io_in_101); // @[Modules.scala 37:46:@314.4]
  assign _T_54557 = _T_54556[4:0]; // @[Modules.scala 37:46:@315.4]
  assign _T_54558 = $signed(_T_54557); // @[Modules.scala 37:46:@316.4]
  assign _T_54559 = $signed(io_in_102) + $signed(io_in_103); // @[Modules.scala 37:46:@318.4]
  assign _T_54560 = _T_54559[4:0]; // @[Modules.scala 37:46:@319.4]
  assign _T_54561 = $signed(_T_54560); // @[Modules.scala 37:46:@320.4]
  assign _T_54562 = $signed(io_in_104) + $signed(io_in_105); // @[Modules.scala 37:46:@322.4]
  assign _T_54563 = _T_54562[4:0]; // @[Modules.scala 37:46:@323.4]
  assign _T_54564 = $signed(_T_54563); // @[Modules.scala 37:46:@324.4]
  assign _T_54565 = $signed(io_in_106) + $signed(io_in_107); // @[Modules.scala 37:46:@326.4]
  assign _T_54566 = _T_54565[4:0]; // @[Modules.scala 37:46:@327.4]
  assign _T_54567 = $signed(_T_54566); // @[Modules.scala 37:46:@328.4]
  assign _T_54568 = $signed(io_in_108) - $signed(io_in_109); // @[Modules.scala 40:46:@330.4]
  assign _T_54569 = _T_54568[4:0]; // @[Modules.scala 40:46:@331.4]
  assign _T_54570 = $signed(_T_54569); // @[Modules.scala 40:46:@332.4]
  assign _T_54571 = $signed(io_in_110) + $signed(io_in_111); // @[Modules.scala 37:46:@334.4]
  assign _T_54572 = _T_54571[4:0]; // @[Modules.scala 37:46:@335.4]
  assign _T_54573 = $signed(_T_54572); // @[Modules.scala 37:46:@336.4]
  assign _T_54575 = $signed(5'sh0) - $signed(io_in_112); // @[Modules.scala 43:37:@338.4]
  assign _T_54576 = _T_54575[4:0]; // @[Modules.scala 43:37:@339.4]
  assign _T_54577 = $signed(_T_54576); // @[Modules.scala 43:37:@340.4]
  assign _T_54578 = $signed(_T_54577) + $signed(io_in_113); // @[Modules.scala 43:47:@341.4]
  assign _T_54579 = _T_54578[4:0]; // @[Modules.scala 43:47:@342.4]
  assign _T_54580 = $signed(_T_54579); // @[Modules.scala 43:47:@343.4]
  assign _T_54582 = $signed(5'sh0) - $signed(io_in_114); // @[Modules.scala 46:37:@345.4]
  assign _T_54583 = _T_54582[4:0]; // @[Modules.scala 46:37:@346.4]
  assign _T_54584 = $signed(_T_54583); // @[Modules.scala 46:37:@347.4]
  assign _T_54585 = $signed(_T_54584) - $signed(io_in_115); // @[Modules.scala 46:47:@348.4]
  assign _T_54586 = _T_54585[4:0]; // @[Modules.scala 46:47:@349.4]
  assign _T_54587 = $signed(_T_54586); // @[Modules.scala 46:47:@350.4]
  assign _T_54588 = $signed(io_in_116) - $signed(io_in_117); // @[Modules.scala 40:46:@352.4]
  assign _T_54589 = _T_54588[4:0]; // @[Modules.scala 40:46:@353.4]
  assign _T_54590 = $signed(_T_54589); // @[Modules.scala 40:46:@354.4]
  assign _T_54591 = $signed(io_in_118) + $signed(io_in_119); // @[Modules.scala 37:46:@356.4]
  assign _T_54592 = _T_54591[4:0]; // @[Modules.scala 37:46:@357.4]
  assign _T_54593 = $signed(_T_54592); // @[Modules.scala 37:46:@358.4]
  assign _T_54595 = $signed(5'sh0) - $signed(io_in_120); // @[Modules.scala 46:37:@360.4]
  assign _T_54596 = _T_54595[4:0]; // @[Modules.scala 46:37:@361.4]
  assign _T_54597 = $signed(_T_54596); // @[Modules.scala 46:37:@362.4]
  assign _T_54598 = $signed(_T_54597) - $signed(io_in_121); // @[Modules.scala 46:47:@363.4]
  assign _T_54599 = _T_54598[4:0]; // @[Modules.scala 46:47:@364.4]
  assign _T_54600 = $signed(_T_54599); // @[Modules.scala 46:47:@365.4]
  assign _T_54602 = $signed(5'sh0) - $signed(io_in_122); // @[Modules.scala 46:37:@367.4]
  assign _T_54603 = _T_54602[4:0]; // @[Modules.scala 46:37:@368.4]
  assign _T_54604 = $signed(_T_54603); // @[Modules.scala 46:37:@369.4]
  assign _T_54605 = $signed(_T_54604) - $signed(io_in_123); // @[Modules.scala 46:47:@370.4]
  assign _T_54606 = _T_54605[4:0]; // @[Modules.scala 46:47:@371.4]
  assign _T_54607 = $signed(_T_54606); // @[Modules.scala 46:47:@372.4]
  assign _T_54609 = $signed(5'sh0) - $signed(io_in_124); // @[Modules.scala 46:37:@374.4]
  assign _T_54610 = _T_54609[4:0]; // @[Modules.scala 46:37:@375.4]
  assign _T_54611 = $signed(_T_54610); // @[Modules.scala 46:37:@376.4]
  assign _T_54612 = $signed(_T_54611) - $signed(io_in_125); // @[Modules.scala 46:47:@377.4]
  assign _T_54613 = _T_54612[4:0]; // @[Modules.scala 46:47:@378.4]
  assign _T_54614 = $signed(_T_54613); // @[Modules.scala 46:47:@379.4]
  assign _T_54616 = $signed(5'sh0) - $signed(io_in_126); // @[Modules.scala 46:37:@381.4]
  assign _T_54617 = _T_54616[4:0]; // @[Modules.scala 46:37:@382.4]
  assign _T_54618 = $signed(_T_54617); // @[Modules.scala 46:37:@383.4]
  assign _T_54619 = $signed(_T_54618) - $signed(io_in_127); // @[Modules.scala 46:47:@384.4]
  assign _T_54620 = _T_54619[4:0]; // @[Modules.scala 46:47:@385.4]
  assign _T_54621 = $signed(_T_54620); // @[Modules.scala 46:47:@386.4]
  assign _T_54623 = $signed(5'sh0) - $signed(io_in_128); // @[Modules.scala 43:37:@388.4]
  assign _T_54624 = _T_54623[4:0]; // @[Modules.scala 43:37:@389.4]
  assign _T_54625 = $signed(_T_54624); // @[Modules.scala 43:37:@390.4]
  assign _T_54626 = $signed(_T_54625) + $signed(io_in_129); // @[Modules.scala 43:47:@391.4]
  assign _T_54627 = _T_54626[4:0]; // @[Modules.scala 43:47:@392.4]
  assign _T_54628 = $signed(_T_54627); // @[Modules.scala 43:47:@393.4]
  assign _T_54630 = $signed(5'sh0) - $signed(io_in_130); // @[Modules.scala 43:37:@395.4]
  assign _T_54631 = _T_54630[4:0]; // @[Modules.scala 43:37:@396.4]
  assign _T_54632 = $signed(_T_54631); // @[Modules.scala 43:37:@397.4]
  assign _T_54633 = $signed(_T_54632) + $signed(io_in_131); // @[Modules.scala 43:47:@398.4]
  assign _T_54634 = _T_54633[4:0]; // @[Modules.scala 43:47:@399.4]
  assign _T_54635 = $signed(_T_54634); // @[Modules.scala 43:47:@400.4]
  assign _T_54636 = $signed(io_in_132) + $signed(io_in_133); // @[Modules.scala 37:46:@402.4]
  assign _T_54637 = _T_54636[4:0]; // @[Modules.scala 37:46:@403.4]
  assign _T_54638 = $signed(_T_54637); // @[Modules.scala 37:46:@404.4]
  assign _T_54639 = $signed(io_in_134) + $signed(io_in_135); // @[Modules.scala 37:46:@406.4]
  assign _T_54640 = _T_54639[4:0]; // @[Modules.scala 37:46:@407.4]
  assign _T_54641 = $signed(_T_54640); // @[Modules.scala 37:46:@408.4]
  assign _T_54642 = $signed(io_in_136) - $signed(io_in_137); // @[Modules.scala 40:46:@410.4]
  assign _T_54643 = _T_54642[4:0]; // @[Modules.scala 40:46:@411.4]
  assign _T_54644 = $signed(_T_54643); // @[Modules.scala 40:46:@412.4]
  assign _T_54646 = $signed(5'sh0) - $signed(io_in_138); // @[Modules.scala 46:37:@414.4]
  assign _T_54647 = _T_54646[4:0]; // @[Modules.scala 46:37:@415.4]
  assign _T_54648 = $signed(_T_54647); // @[Modules.scala 46:37:@416.4]
  assign _T_54649 = $signed(_T_54648) - $signed(io_in_139); // @[Modules.scala 46:47:@417.4]
  assign _T_54650 = _T_54649[4:0]; // @[Modules.scala 46:47:@418.4]
  assign _T_54651 = $signed(_T_54650); // @[Modules.scala 46:47:@419.4]
  assign _T_54652 = $signed(io_in_140) + $signed(io_in_141); // @[Modules.scala 37:46:@421.4]
  assign _T_54653 = _T_54652[4:0]; // @[Modules.scala 37:46:@422.4]
  assign _T_54654 = $signed(_T_54653); // @[Modules.scala 37:46:@423.4]
  assign _T_54656 = $signed(5'sh0) - $signed(io_in_142); // @[Modules.scala 46:37:@425.4]
  assign _T_54657 = _T_54656[4:0]; // @[Modules.scala 46:37:@426.4]
  assign _T_54658 = $signed(_T_54657); // @[Modules.scala 46:37:@427.4]
  assign _T_54659 = $signed(_T_54658) - $signed(io_in_143); // @[Modules.scala 46:47:@428.4]
  assign _T_54660 = _T_54659[4:0]; // @[Modules.scala 46:47:@429.4]
  assign _T_54661 = $signed(_T_54660); // @[Modules.scala 46:47:@430.4]
  assign _T_54662 = $signed(io_in_144) - $signed(io_in_145); // @[Modules.scala 40:46:@432.4]
  assign _T_54663 = _T_54662[4:0]; // @[Modules.scala 40:46:@433.4]
  assign _T_54664 = $signed(_T_54663); // @[Modules.scala 40:46:@434.4]
  assign _T_54665 = $signed(io_in_146) + $signed(io_in_147); // @[Modules.scala 37:46:@436.4]
  assign _T_54666 = _T_54665[4:0]; // @[Modules.scala 37:46:@437.4]
  assign _T_54667 = $signed(_T_54666); // @[Modules.scala 37:46:@438.4]
  assign _T_54668 = $signed(io_in_148) + $signed(io_in_149); // @[Modules.scala 37:46:@440.4]
  assign _T_54669 = _T_54668[4:0]; // @[Modules.scala 37:46:@441.4]
  assign _T_54670 = $signed(_T_54669); // @[Modules.scala 37:46:@442.4]
  assign _T_54672 = $signed(5'sh0) - $signed(io_in_150); // @[Modules.scala 46:37:@444.4]
  assign _T_54673 = _T_54672[4:0]; // @[Modules.scala 46:37:@445.4]
  assign _T_54674 = $signed(_T_54673); // @[Modules.scala 46:37:@446.4]
  assign _T_54675 = $signed(_T_54674) - $signed(io_in_151); // @[Modules.scala 46:47:@447.4]
  assign _T_54676 = _T_54675[4:0]; // @[Modules.scala 46:47:@448.4]
  assign _T_54677 = $signed(_T_54676); // @[Modules.scala 46:47:@449.4]
  assign _T_54679 = $signed(5'sh0) - $signed(io_in_152); // @[Modules.scala 46:37:@451.4]
  assign _T_54680 = _T_54679[4:0]; // @[Modules.scala 46:37:@452.4]
  assign _T_54681 = $signed(_T_54680); // @[Modules.scala 46:37:@453.4]
  assign _T_54682 = $signed(_T_54681) - $signed(io_in_153); // @[Modules.scala 46:47:@454.4]
  assign _T_54683 = _T_54682[4:0]; // @[Modules.scala 46:47:@455.4]
  assign _T_54684 = $signed(_T_54683); // @[Modules.scala 46:47:@456.4]
  assign _T_54686 = $signed(5'sh0) - $signed(io_in_154); // @[Modules.scala 46:37:@458.4]
  assign _T_54687 = _T_54686[4:0]; // @[Modules.scala 46:37:@459.4]
  assign _T_54688 = $signed(_T_54687); // @[Modules.scala 46:37:@460.4]
  assign _T_54689 = $signed(_T_54688) - $signed(io_in_155); // @[Modules.scala 46:47:@461.4]
  assign _T_54690 = _T_54689[4:0]; // @[Modules.scala 46:47:@462.4]
  assign _T_54691 = $signed(_T_54690); // @[Modules.scala 46:47:@463.4]
  assign _T_54693 = $signed(5'sh0) - $signed(io_in_156); // @[Modules.scala 46:37:@465.4]
  assign _T_54694 = _T_54693[4:0]; // @[Modules.scala 46:37:@466.4]
  assign _T_54695 = $signed(_T_54694); // @[Modules.scala 46:37:@467.4]
  assign _T_54696 = $signed(_T_54695) - $signed(io_in_157); // @[Modules.scala 46:47:@468.4]
  assign _T_54697 = _T_54696[4:0]; // @[Modules.scala 46:47:@469.4]
  assign _T_54698 = $signed(_T_54697); // @[Modules.scala 46:47:@470.4]
  assign _T_54700 = $signed(5'sh0) - $signed(io_in_158); // @[Modules.scala 46:37:@472.4]
  assign _T_54701 = _T_54700[4:0]; // @[Modules.scala 46:37:@473.4]
  assign _T_54702 = $signed(_T_54701); // @[Modules.scala 46:37:@474.4]
  assign _T_54703 = $signed(_T_54702) - $signed(io_in_159); // @[Modules.scala 46:47:@475.4]
  assign _T_54704 = _T_54703[4:0]; // @[Modules.scala 46:47:@476.4]
  assign _T_54705 = $signed(_T_54704); // @[Modules.scala 46:47:@477.4]
  assign _T_54707 = $signed(5'sh0) - $signed(io_in_160); // @[Modules.scala 46:37:@479.4]
  assign _T_54708 = _T_54707[4:0]; // @[Modules.scala 46:37:@480.4]
  assign _T_54709 = $signed(_T_54708); // @[Modules.scala 46:37:@481.4]
  assign _T_54710 = $signed(_T_54709) - $signed(io_in_161); // @[Modules.scala 46:47:@482.4]
  assign _T_54711 = _T_54710[4:0]; // @[Modules.scala 46:47:@483.4]
  assign _T_54712 = $signed(_T_54711); // @[Modules.scala 46:47:@484.4]
  assign _T_54713 = $signed(io_in_162) + $signed(io_in_163); // @[Modules.scala 37:46:@486.4]
  assign _T_54714 = _T_54713[4:0]; // @[Modules.scala 37:46:@487.4]
  assign _T_54715 = $signed(_T_54714); // @[Modules.scala 37:46:@488.4]
  assign _T_54716 = $signed(io_in_164) - $signed(io_in_165); // @[Modules.scala 40:46:@490.4]
  assign _T_54717 = _T_54716[4:0]; // @[Modules.scala 40:46:@491.4]
  assign _T_54718 = $signed(_T_54717); // @[Modules.scala 40:46:@492.4]
  assign _T_54720 = $signed(5'sh0) - $signed(io_in_166); // @[Modules.scala 43:37:@494.4]
  assign _T_54721 = _T_54720[4:0]; // @[Modules.scala 43:37:@495.4]
  assign _T_54722 = $signed(_T_54721); // @[Modules.scala 43:37:@496.4]
  assign _T_54723 = $signed(_T_54722) + $signed(io_in_167); // @[Modules.scala 43:47:@497.4]
  assign _T_54724 = _T_54723[4:0]; // @[Modules.scala 43:47:@498.4]
  assign _T_54725 = $signed(_T_54724); // @[Modules.scala 43:47:@499.4]
  assign _T_54727 = $signed(5'sh0) - $signed(io_in_168); // @[Modules.scala 46:37:@501.4]
  assign _T_54728 = _T_54727[4:0]; // @[Modules.scala 46:37:@502.4]
  assign _T_54729 = $signed(_T_54728); // @[Modules.scala 46:37:@503.4]
  assign _T_54730 = $signed(_T_54729) - $signed(io_in_169); // @[Modules.scala 46:47:@504.4]
  assign _T_54731 = _T_54730[4:0]; // @[Modules.scala 46:47:@505.4]
  assign _T_54732 = $signed(_T_54731); // @[Modules.scala 46:47:@506.4]
  assign _T_54734 = $signed(5'sh0) - $signed(io_in_170); // @[Modules.scala 46:37:@508.4]
  assign _T_54735 = _T_54734[4:0]; // @[Modules.scala 46:37:@509.4]
  assign _T_54736 = $signed(_T_54735); // @[Modules.scala 46:37:@510.4]
  assign _T_54737 = $signed(_T_54736) - $signed(io_in_171); // @[Modules.scala 46:47:@511.4]
  assign _T_54738 = _T_54737[4:0]; // @[Modules.scala 46:47:@512.4]
  assign _T_54739 = $signed(_T_54738); // @[Modules.scala 46:47:@513.4]
  assign _T_54740 = $signed(io_in_172) - $signed(io_in_173); // @[Modules.scala 40:46:@515.4]
  assign _T_54741 = _T_54740[4:0]; // @[Modules.scala 40:46:@516.4]
  assign _T_54742 = $signed(_T_54741); // @[Modules.scala 40:46:@517.4]
  assign _T_54744 = $signed(5'sh0) - $signed(io_in_174); // @[Modules.scala 46:37:@519.4]
  assign _T_54745 = _T_54744[4:0]; // @[Modules.scala 46:37:@520.4]
  assign _T_54746 = $signed(_T_54745); // @[Modules.scala 46:37:@521.4]
  assign _T_54747 = $signed(_T_54746) - $signed(io_in_175); // @[Modules.scala 46:47:@522.4]
  assign _T_54748 = _T_54747[4:0]; // @[Modules.scala 46:47:@523.4]
  assign _T_54749 = $signed(_T_54748); // @[Modules.scala 46:47:@524.4]
  assign _T_54751 = $signed(5'sh0) - $signed(io_in_176); // @[Modules.scala 46:37:@526.4]
  assign _T_54752 = _T_54751[4:0]; // @[Modules.scala 46:37:@527.4]
  assign _T_54753 = $signed(_T_54752); // @[Modules.scala 46:37:@528.4]
  assign _T_54754 = $signed(_T_54753) - $signed(io_in_177); // @[Modules.scala 46:47:@529.4]
  assign _T_54755 = _T_54754[4:0]; // @[Modules.scala 46:47:@530.4]
  assign _T_54756 = $signed(_T_54755); // @[Modules.scala 46:47:@531.4]
  assign _T_54758 = $signed(5'sh0) - $signed(io_in_178); // @[Modules.scala 46:37:@533.4]
  assign _T_54759 = _T_54758[4:0]; // @[Modules.scala 46:37:@534.4]
  assign _T_54760 = $signed(_T_54759); // @[Modules.scala 46:37:@535.4]
  assign _T_54761 = $signed(_T_54760) - $signed(io_in_179); // @[Modules.scala 46:47:@536.4]
  assign _T_54762 = _T_54761[4:0]; // @[Modules.scala 46:47:@537.4]
  assign _T_54763 = $signed(_T_54762); // @[Modules.scala 46:47:@538.4]
  assign _T_54765 = $signed(5'sh0) - $signed(io_in_180); // @[Modules.scala 46:37:@540.4]
  assign _T_54766 = _T_54765[4:0]; // @[Modules.scala 46:37:@541.4]
  assign _T_54767 = $signed(_T_54766); // @[Modules.scala 46:37:@542.4]
  assign _T_54768 = $signed(_T_54767) - $signed(io_in_181); // @[Modules.scala 46:47:@543.4]
  assign _T_54769 = _T_54768[4:0]; // @[Modules.scala 46:47:@544.4]
  assign _T_54770 = $signed(_T_54769); // @[Modules.scala 46:47:@545.4]
  assign _T_54772 = $signed(5'sh0) - $signed(io_in_182); // @[Modules.scala 46:37:@547.4]
  assign _T_54773 = _T_54772[4:0]; // @[Modules.scala 46:37:@548.4]
  assign _T_54774 = $signed(_T_54773); // @[Modules.scala 46:37:@549.4]
  assign _T_54775 = $signed(_T_54774) - $signed(io_in_183); // @[Modules.scala 46:47:@550.4]
  assign _T_54776 = _T_54775[4:0]; // @[Modules.scala 46:47:@551.4]
  assign _T_54777 = $signed(_T_54776); // @[Modules.scala 46:47:@552.4]
  assign _T_54779 = $signed(5'sh0) - $signed(io_in_184); // @[Modules.scala 46:37:@554.4]
  assign _T_54780 = _T_54779[4:0]; // @[Modules.scala 46:37:@555.4]
  assign _T_54781 = $signed(_T_54780); // @[Modules.scala 46:37:@556.4]
  assign _T_54782 = $signed(_T_54781) - $signed(io_in_185); // @[Modules.scala 46:47:@557.4]
  assign _T_54783 = _T_54782[4:0]; // @[Modules.scala 46:47:@558.4]
  assign _T_54784 = $signed(_T_54783); // @[Modules.scala 46:47:@559.4]
  assign _T_54785 = $signed(io_in_186) + $signed(io_in_187); // @[Modules.scala 37:46:@561.4]
  assign _T_54786 = _T_54785[4:0]; // @[Modules.scala 37:46:@562.4]
  assign _T_54787 = $signed(_T_54786); // @[Modules.scala 37:46:@563.4]
  assign _T_54789 = $signed(5'sh0) - $signed(io_in_188); // @[Modules.scala 46:37:@565.4]
  assign _T_54790 = _T_54789[4:0]; // @[Modules.scala 46:37:@566.4]
  assign _T_54791 = $signed(_T_54790); // @[Modules.scala 46:37:@567.4]
  assign _T_54792 = $signed(_T_54791) - $signed(io_in_189); // @[Modules.scala 46:47:@568.4]
  assign _T_54793 = _T_54792[4:0]; // @[Modules.scala 46:47:@569.4]
  assign _T_54794 = $signed(_T_54793); // @[Modules.scala 46:47:@570.4]
  assign _T_54795 = $signed(io_in_190) - $signed(io_in_191); // @[Modules.scala 40:46:@572.4]
  assign _T_54796 = _T_54795[4:0]; // @[Modules.scala 40:46:@573.4]
  assign _T_54797 = $signed(_T_54796); // @[Modules.scala 40:46:@574.4]
  assign _T_54799 = $signed(5'sh0) - $signed(io_in_192); // @[Modules.scala 46:37:@576.4]
  assign _T_54800 = _T_54799[4:0]; // @[Modules.scala 46:37:@577.4]
  assign _T_54801 = $signed(_T_54800); // @[Modules.scala 46:37:@578.4]
  assign _T_54802 = $signed(_T_54801) - $signed(io_in_193); // @[Modules.scala 46:47:@579.4]
  assign _T_54803 = _T_54802[4:0]; // @[Modules.scala 46:47:@580.4]
  assign _T_54804 = $signed(_T_54803); // @[Modules.scala 46:47:@581.4]
  assign _T_54806 = $signed(5'sh0) - $signed(io_in_194); // @[Modules.scala 46:37:@583.4]
  assign _T_54807 = _T_54806[4:0]; // @[Modules.scala 46:37:@584.4]
  assign _T_54808 = $signed(_T_54807); // @[Modules.scala 46:37:@585.4]
  assign _T_54809 = $signed(_T_54808) - $signed(io_in_195); // @[Modules.scala 46:47:@586.4]
  assign _T_54810 = _T_54809[4:0]; // @[Modules.scala 46:47:@587.4]
  assign _T_54811 = $signed(_T_54810); // @[Modules.scala 46:47:@588.4]
  assign _T_54812 = $signed(io_in_196) - $signed(io_in_197); // @[Modules.scala 40:46:@590.4]
  assign _T_54813 = _T_54812[4:0]; // @[Modules.scala 40:46:@591.4]
  assign _T_54814 = $signed(_T_54813); // @[Modules.scala 40:46:@592.4]
  assign _T_54815 = $signed(io_in_198) - $signed(io_in_199); // @[Modules.scala 40:46:@594.4]
  assign _T_54816 = _T_54815[4:0]; // @[Modules.scala 40:46:@595.4]
  assign _T_54817 = $signed(_T_54816); // @[Modules.scala 40:46:@596.4]
  assign _T_54819 = $signed(5'sh0) - $signed(io_in_200); // @[Modules.scala 46:37:@598.4]
  assign _T_54820 = _T_54819[4:0]; // @[Modules.scala 46:37:@599.4]
  assign _T_54821 = $signed(_T_54820); // @[Modules.scala 46:37:@600.4]
  assign _T_54822 = $signed(_T_54821) - $signed(io_in_201); // @[Modules.scala 46:47:@601.4]
  assign _T_54823 = _T_54822[4:0]; // @[Modules.scala 46:47:@602.4]
  assign _T_54824 = $signed(_T_54823); // @[Modules.scala 46:47:@603.4]
  assign _T_54826 = $signed(5'sh0) - $signed(io_in_202); // @[Modules.scala 46:37:@605.4]
  assign _T_54827 = _T_54826[4:0]; // @[Modules.scala 46:37:@606.4]
  assign _T_54828 = $signed(_T_54827); // @[Modules.scala 46:37:@607.4]
  assign _T_54829 = $signed(_T_54828) - $signed(io_in_203); // @[Modules.scala 46:47:@608.4]
  assign _T_54830 = _T_54829[4:0]; // @[Modules.scala 46:47:@609.4]
  assign _T_54831 = $signed(_T_54830); // @[Modules.scala 46:47:@610.4]
  assign _T_54833 = $signed(5'sh0) - $signed(io_in_204); // @[Modules.scala 46:37:@612.4]
  assign _T_54834 = _T_54833[4:0]; // @[Modules.scala 46:37:@613.4]
  assign _T_54835 = $signed(_T_54834); // @[Modules.scala 46:37:@614.4]
  assign _T_54836 = $signed(_T_54835) - $signed(io_in_205); // @[Modules.scala 46:47:@615.4]
  assign _T_54837 = _T_54836[4:0]; // @[Modules.scala 46:47:@616.4]
  assign _T_54838 = $signed(_T_54837); // @[Modules.scala 46:47:@617.4]
  assign _T_54840 = $signed(5'sh0) - $signed(io_in_206); // @[Modules.scala 43:37:@619.4]
  assign _T_54841 = _T_54840[4:0]; // @[Modules.scala 43:37:@620.4]
  assign _T_54842 = $signed(_T_54841); // @[Modules.scala 43:37:@621.4]
  assign _T_54843 = $signed(_T_54842) + $signed(io_in_207); // @[Modules.scala 43:47:@622.4]
  assign _T_54844 = _T_54843[4:0]; // @[Modules.scala 43:47:@623.4]
  assign _T_54845 = $signed(_T_54844); // @[Modules.scala 43:47:@624.4]
  assign _T_54847 = $signed(5'sh0) - $signed(io_in_208); // @[Modules.scala 43:37:@626.4]
  assign _T_54848 = _T_54847[4:0]; // @[Modules.scala 43:37:@627.4]
  assign _T_54849 = $signed(_T_54848); // @[Modules.scala 43:37:@628.4]
  assign _T_54850 = $signed(_T_54849) + $signed(io_in_209); // @[Modules.scala 43:47:@629.4]
  assign _T_54851 = _T_54850[4:0]; // @[Modules.scala 43:47:@630.4]
  assign _T_54852 = $signed(_T_54851); // @[Modules.scala 43:47:@631.4]
  assign _T_54853 = $signed(io_in_210) + $signed(io_in_211); // @[Modules.scala 37:46:@633.4]
  assign _T_54854 = _T_54853[4:0]; // @[Modules.scala 37:46:@634.4]
  assign _T_54855 = $signed(_T_54854); // @[Modules.scala 37:46:@635.4]
  assign _T_54856 = $signed(io_in_212) - $signed(io_in_213); // @[Modules.scala 40:46:@637.4]
  assign _T_54857 = _T_54856[4:0]; // @[Modules.scala 40:46:@638.4]
  assign _T_54858 = $signed(_T_54857); // @[Modules.scala 40:46:@639.4]
  assign _T_54860 = $signed(5'sh0) - $signed(io_in_214); // @[Modules.scala 46:37:@641.4]
  assign _T_54861 = _T_54860[4:0]; // @[Modules.scala 46:37:@642.4]
  assign _T_54862 = $signed(_T_54861); // @[Modules.scala 46:37:@643.4]
  assign _T_54863 = $signed(_T_54862) - $signed(io_in_215); // @[Modules.scala 46:47:@644.4]
  assign _T_54864 = _T_54863[4:0]; // @[Modules.scala 46:47:@645.4]
  assign _T_54865 = $signed(_T_54864); // @[Modules.scala 46:47:@646.4]
  assign _T_54867 = $signed(5'sh0) - $signed(io_in_216); // @[Modules.scala 46:37:@648.4]
  assign _T_54868 = _T_54867[4:0]; // @[Modules.scala 46:37:@649.4]
  assign _T_54869 = $signed(_T_54868); // @[Modules.scala 46:37:@650.4]
  assign _T_54870 = $signed(_T_54869) - $signed(io_in_217); // @[Modules.scala 46:47:@651.4]
  assign _T_54871 = _T_54870[4:0]; // @[Modules.scala 46:47:@652.4]
  assign _T_54872 = $signed(_T_54871); // @[Modules.scala 46:47:@653.4]
  assign _T_54874 = $signed(5'sh0) - $signed(io_in_218); // @[Modules.scala 46:37:@655.4]
  assign _T_54875 = _T_54874[4:0]; // @[Modules.scala 46:37:@656.4]
  assign _T_54876 = $signed(_T_54875); // @[Modules.scala 46:37:@657.4]
  assign _T_54877 = $signed(_T_54876) - $signed(io_in_219); // @[Modules.scala 46:47:@658.4]
  assign _T_54878 = _T_54877[4:0]; // @[Modules.scala 46:47:@659.4]
  assign _T_54879 = $signed(_T_54878); // @[Modules.scala 46:47:@660.4]
  assign _T_54881 = $signed(5'sh0) - $signed(io_in_220); // @[Modules.scala 46:37:@662.4]
  assign _T_54882 = _T_54881[4:0]; // @[Modules.scala 46:37:@663.4]
  assign _T_54883 = $signed(_T_54882); // @[Modules.scala 46:37:@664.4]
  assign _T_54884 = $signed(_T_54883) - $signed(io_in_221); // @[Modules.scala 46:47:@665.4]
  assign _T_54885 = _T_54884[4:0]; // @[Modules.scala 46:47:@666.4]
  assign _T_54886 = $signed(_T_54885); // @[Modules.scala 46:47:@667.4]
  assign _T_54888 = $signed(5'sh0) - $signed(io_in_222); // @[Modules.scala 46:37:@669.4]
  assign _T_54889 = _T_54888[4:0]; // @[Modules.scala 46:37:@670.4]
  assign _T_54890 = $signed(_T_54889); // @[Modules.scala 46:37:@671.4]
  assign _T_54891 = $signed(_T_54890) - $signed(io_in_223); // @[Modules.scala 46:47:@672.4]
  assign _T_54892 = _T_54891[4:0]; // @[Modules.scala 46:47:@673.4]
  assign _T_54893 = $signed(_T_54892); // @[Modules.scala 46:47:@674.4]
  assign _T_54895 = $signed(5'sh0) - $signed(io_in_224); // @[Modules.scala 46:37:@676.4]
  assign _T_54896 = _T_54895[4:0]; // @[Modules.scala 46:37:@677.4]
  assign _T_54897 = $signed(_T_54896); // @[Modules.scala 46:37:@678.4]
  assign _T_54898 = $signed(_T_54897) - $signed(io_in_225); // @[Modules.scala 46:47:@679.4]
  assign _T_54899 = _T_54898[4:0]; // @[Modules.scala 46:47:@680.4]
  assign _T_54900 = $signed(_T_54899); // @[Modules.scala 46:47:@681.4]
  assign _T_54902 = $signed(5'sh0) - $signed(io_in_226); // @[Modules.scala 46:37:@683.4]
  assign _T_54903 = _T_54902[4:0]; // @[Modules.scala 46:37:@684.4]
  assign _T_54904 = $signed(_T_54903); // @[Modules.scala 46:37:@685.4]
  assign _T_54905 = $signed(_T_54904) - $signed(io_in_227); // @[Modules.scala 46:47:@686.4]
  assign _T_54906 = _T_54905[4:0]; // @[Modules.scala 46:47:@687.4]
  assign _T_54907 = $signed(_T_54906); // @[Modules.scala 46:47:@688.4]
  assign _T_54909 = $signed(5'sh0) - $signed(io_in_228); // @[Modules.scala 46:37:@690.4]
  assign _T_54910 = _T_54909[4:0]; // @[Modules.scala 46:37:@691.4]
  assign _T_54911 = $signed(_T_54910); // @[Modules.scala 46:37:@692.4]
  assign _T_54912 = $signed(_T_54911) - $signed(io_in_229); // @[Modules.scala 46:47:@693.4]
  assign _T_54913 = _T_54912[4:0]; // @[Modules.scala 46:47:@694.4]
  assign _T_54914 = $signed(_T_54913); // @[Modules.scala 46:47:@695.4]
  assign _T_54916 = $signed(5'sh0) - $signed(io_in_230); // @[Modules.scala 46:37:@697.4]
  assign _T_54917 = _T_54916[4:0]; // @[Modules.scala 46:37:@698.4]
  assign _T_54918 = $signed(_T_54917); // @[Modules.scala 46:37:@699.4]
  assign _T_54919 = $signed(_T_54918) - $signed(io_in_231); // @[Modules.scala 46:47:@700.4]
  assign _T_54920 = _T_54919[4:0]; // @[Modules.scala 46:47:@701.4]
  assign _T_54921 = $signed(_T_54920); // @[Modules.scala 46:47:@702.4]
  assign _T_54923 = $signed(5'sh0) - $signed(io_in_232); // @[Modules.scala 46:37:@704.4]
  assign _T_54924 = _T_54923[4:0]; // @[Modules.scala 46:37:@705.4]
  assign _T_54925 = $signed(_T_54924); // @[Modules.scala 46:37:@706.4]
  assign _T_54926 = $signed(_T_54925) - $signed(io_in_233); // @[Modules.scala 46:47:@707.4]
  assign _T_54927 = _T_54926[4:0]; // @[Modules.scala 46:47:@708.4]
  assign _T_54928 = $signed(_T_54927); // @[Modules.scala 46:47:@709.4]
  assign _T_54930 = $signed(5'sh0) - $signed(io_in_234); // @[Modules.scala 46:37:@711.4]
  assign _T_54931 = _T_54930[4:0]; // @[Modules.scala 46:37:@712.4]
  assign _T_54932 = $signed(_T_54931); // @[Modules.scala 46:37:@713.4]
  assign _T_54933 = $signed(_T_54932) - $signed(io_in_235); // @[Modules.scala 46:47:@714.4]
  assign _T_54934 = _T_54933[4:0]; // @[Modules.scala 46:47:@715.4]
  assign _T_54935 = $signed(_T_54934); // @[Modules.scala 46:47:@716.4]
  assign _T_54937 = $signed(5'sh0) - $signed(io_in_236); // @[Modules.scala 43:37:@718.4]
  assign _T_54938 = _T_54937[4:0]; // @[Modules.scala 43:37:@719.4]
  assign _T_54939 = $signed(_T_54938); // @[Modules.scala 43:37:@720.4]
  assign _T_54940 = $signed(_T_54939) + $signed(io_in_237); // @[Modules.scala 43:47:@721.4]
  assign _T_54941 = _T_54940[4:0]; // @[Modules.scala 43:47:@722.4]
  assign _T_54942 = $signed(_T_54941); // @[Modules.scala 43:47:@723.4]
  assign _T_54944 = $signed(5'sh0) - $signed(io_in_238); // @[Modules.scala 46:37:@725.4]
  assign _T_54945 = _T_54944[4:0]; // @[Modules.scala 46:37:@726.4]
  assign _T_54946 = $signed(_T_54945); // @[Modules.scala 46:37:@727.4]
  assign _T_54947 = $signed(_T_54946) - $signed(io_in_239); // @[Modules.scala 46:47:@728.4]
  assign _T_54948 = _T_54947[4:0]; // @[Modules.scala 46:47:@729.4]
  assign _T_54949 = $signed(_T_54948); // @[Modules.scala 46:47:@730.4]
  assign _T_54951 = $signed(5'sh0) - $signed(io_in_240); // @[Modules.scala 46:37:@732.4]
  assign _T_54952 = _T_54951[4:0]; // @[Modules.scala 46:37:@733.4]
  assign _T_54953 = $signed(_T_54952); // @[Modules.scala 46:37:@734.4]
  assign _T_54954 = $signed(_T_54953) - $signed(io_in_241); // @[Modules.scala 46:47:@735.4]
  assign _T_54955 = _T_54954[4:0]; // @[Modules.scala 46:47:@736.4]
  assign _T_54956 = $signed(_T_54955); // @[Modules.scala 46:47:@737.4]
  assign _T_54958 = $signed(5'sh0) - $signed(io_in_242); // @[Modules.scala 46:37:@739.4]
  assign _T_54959 = _T_54958[4:0]; // @[Modules.scala 46:37:@740.4]
  assign _T_54960 = $signed(_T_54959); // @[Modules.scala 46:37:@741.4]
  assign _T_54961 = $signed(_T_54960) - $signed(io_in_243); // @[Modules.scala 46:47:@742.4]
  assign _T_54962 = _T_54961[4:0]; // @[Modules.scala 46:47:@743.4]
  assign _T_54963 = $signed(_T_54962); // @[Modules.scala 46:47:@744.4]
  assign _T_54965 = $signed(5'sh0) - $signed(io_in_244); // @[Modules.scala 46:37:@746.4]
  assign _T_54966 = _T_54965[4:0]; // @[Modules.scala 46:37:@747.4]
  assign _T_54967 = $signed(_T_54966); // @[Modules.scala 46:37:@748.4]
  assign _T_54968 = $signed(_T_54967) - $signed(io_in_245); // @[Modules.scala 46:47:@749.4]
  assign _T_54969 = _T_54968[4:0]; // @[Modules.scala 46:47:@750.4]
  assign _T_54970 = $signed(_T_54969); // @[Modules.scala 46:47:@751.4]
  assign _T_54972 = $signed(5'sh0) - $signed(io_in_246); // @[Modules.scala 46:37:@753.4]
  assign _T_54973 = _T_54972[4:0]; // @[Modules.scala 46:37:@754.4]
  assign _T_54974 = $signed(_T_54973); // @[Modules.scala 46:37:@755.4]
  assign _T_54975 = $signed(_T_54974) - $signed(io_in_247); // @[Modules.scala 46:47:@756.4]
  assign _T_54976 = _T_54975[4:0]; // @[Modules.scala 46:47:@757.4]
  assign _T_54977 = $signed(_T_54976); // @[Modules.scala 46:47:@758.4]
  assign _T_54979 = $signed(5'sh0) - $signed(io_in_248); // @[Modules.scala 46:37:@760.4]
  assign _T_54980 = _T_54979[4:0]; // @[Modules.scala 46:37:@761.4]
  assign _T_54981 = $signed(_T_54980); // @[Modules.scala 46:37:@762.4]
  assign _T_54982 = $signed(_T_54981) - $signed(io_in_249); // @[Modules.scala 46:47:@763.4]
  assign _T_54983 = _T_54982[4:0]; // @[Modules.scala 46:47:@764.4]
  assign _T_54984 = $signed(_T_54983); // @[Modules.scala 46:47:@765.4]
  assign _T_54986 = $signed(5'sh0) - $signed(io_in_250); // @[Modules.scala 46:37:@767.4]
  assign _T_54987 = _T_54986[4:0]; // @[Modules.scala 46:37:@768.4]
  assign _T_54988 = $signed(_T_54987); // @[Modules.scala 46:37:@769.4]
  assign _T_54989 = $signed(_T_54988) - $signed(io_in_251); // @[Modules.scala 46:47:@770.4]
  assign _T_54990 = _T_54989[4:0]; // @[Modules.scala 46:47:@771.4]
  assign _T_54991 = $signed(_T_54990); // @[Modules.scala 46:47:@772.4]
  assign _T_54993 = $signed(5'sh0) - $signed(io_in_252); // @[Modules.scala 46:37:@774.4]
  assign _T_54994 = _T_54993[4:0]; // @[Modules.scala 46:37:@775.4]
  assign _T_54995 = $signed(_T_54994); // @[Modules.scala 46:37:@776.4]
  assign _T_54996 = $signed(_T_54995) - $signed(io_in_253); // @[Modules.scala 46:47:@777.4]
  assign _T_54997 = _T_54996[4:0]; // @[Modules.scala 46:47:@778.4]
  assign _T_54998 = $signed(_T_54997); // @[Modules.scala 46:47:@779.4]
  assign _T_55000 = $signed(5'sh0) - $signed(io_in_254); // @[Modules.scala 46:37:@781.4]
  assign _T_55001 = _T_55000[4:0]; // @[Modules.scala 46:37:@782.4]
  assign _T_55002 = $signed(_T_55001); // @[Modules.scala 46:37:@783.4]
  assign _T_55003 = $signed(_T_55002) - $signed(io_in_255); // @[Modules.scala 46:47:@784.4]
  assign _T_55004 = _T_55003[4:0]; // @[Modules.scala 46:47:@785.4]
  assign _T_55005 = $signed(_T_55004); // @[Modules.scala 46:47:@786.4]
  assign _T_55007 = $signed(5'sh0) - $signed(io_in_256); // @[Modules.scala 46:37:@788.4]
  assign _T_55008 = _T_55007[4:0]; // @[Modules.scala 46:37:@789.4]
  assign _T_55009 = $signed(_T_55008); // @[Modules.scala 46:37:@790.4]
  assign _T_55010 = $signed(_T_55009) - $signed(io_in_257); // @[Modules.scala 46:47:@791.4]
  assign _T_55011 = _T_55010[4:0]; // @[Modules.scala 46:47:@792.4]
  assign _T_55012 = $signed(_T_55011); // @[Modules.scala 46:47:@793.4]
  assign _T_55014 = $signed(5'sh0) - $signed(io_in_258); // @[Modules.scala 46:37:@795.4]
  assign _T_55015 = _T_55014[4:0]; // @[Modules.scala 46:37:@796.4]
  assign _T_55016 = $signed(_T_55015); // @[Modules.scala 46:37:@797.4]
  assign _T_55017 = $signed(_T_55016) - $signed(io_in_259); // @[Modules.scala 46:47:@798.4]
  assign _T_55018 = _T_55017[4:0]; // @[Modules.scala 46:47:@799.4]
  assign _T_55019 = $signed(_T_55018); // @[Modules.scala 46:47:@800.4]
  assign _T_55021 = $signed(5'sh0) - $signed(io_in_260); // @[Modules.scala 46:37:@802.4]
  assign _T_55022 = _T_55021[4:0]; // @[Modules.scala 46:37:@803.4]
  assign _T_55023 = $signed(_T_55022); // @[Modules.scala 46:37:@804.4]
  assign _T_55024 = $signed(_T_55023) - $signed(io_in_261); // @[Modules.scala 46:47:@805.4]
  assign _T_55025 = _T_55024[4:0]; // @[Modules.scala 46:47:@806.4]
  assign _T_55026 = $signed(_T_55025); // @[Modules.scala 46:47:@807.4]
  assign _T_55027 = $signed(io_in_262) - $signed(io_in_263); // @[Modules.scala 40:46:@809.4]
  assign _T_55028 = _T_55027[4:0]; // @[Modules.scala 40:46:@810.4]
  assign _T_55029 = $signed(_T_55028); // @[Modules.scala 40:46:@811.4]
  assign _T_55031 = $signed(5'sh0) - $signed(io_in_264); // @[Modules.scala 46:37:@813.4]
  assign _T_55032 = _T_55031[4:0]; // @[Modules.scala 46:37:@814.4]
  assign _T_55033 = $signed(_T_55032); // @[Modules.scala 46:37:@815.4]
  assign _T_55034 = $signed(_T_55033) - $signed(io_in_265); // @[Modules.scala 46:47:@816.4]
  assign _T_55035 = _T_55034[4:0]; // @[Modules.scala 46:47:@817.4]
  assign _T_55036 = $signed(_T_55035); // @[Modules.scala 46:47:@818.4]
  assign _T_55038 = $signed(5'sh0) - $signed(io_in_266); // @[Modules.scala 46:37:@820.4]
  assign _T_55039 = _T_55038[4:0]; // @[Modules.scala 46:37:@821.4]
  assign _T_55040 = $signed(_T_55039); // @[Modules.scala 46:37:@822.4]
  assign _T_55041 = $signed(_T_55040) - $signed(io_in_267); // @[Modules.scala 46:47:@823.4]
  assign _T_55042 = _T_55041[4:0]; // @[Modules.scala 46:47:@824.4]
  assign _T_55043 = $signed(_T_55042); // @[Modules.scala 46:47:@825.4]
  assign _T_55045 = $signed(5'sh0) - $signed(io_in_268); // @[Modules.scala 46:37:@827.4]
  assign _T_55046 = _T_55045[4:0]; // @[Modules.scala 46:37:@828.4]
  assign _T_55047 = $signed(_T_55046); // @[Modules.scala 46:37:@829.4]
  assign _T_55048 = $signed(_T_55047) - $signed(io_in_269); // @[Modules.scala 46:47:@830.4]
  assign _T_55049 = _T_55048[4:0]; // @[Modules.scala 46:47:@831.4]
  assign _T_55050 = $signed(_T_55049); // @[Modules.scala 46:47:@832.4]
  assign _T_55052 = $signed(5'sh0) - $signed(io_in_270); // @[Modules.scala 46:37:@834.4]
  assign _T_55053 = _T_55052[4:0]; // @[Modules.scala 46:37:@835.4]
  assign _T_55054 = $signed(_T_55053); // @[Modules.scala 46:37:@836.4]
  assign _T_55055 = $signed(_T_55054) - $signed(io_in_271); // @[Modules.scala 46:47:@837.4]
  assign _T_55056 = _T_55055[4:0]; // @[Modules.scala 46:47:@838.4]
  assign _T_55057 = $signed(_T_55056); // @[Modules.scala 46:47:@839.4]
  assign _T_55059 = $signed(5'sh0) - $signed(io_in_272); // @[Modules.scala 46:37:@841.4]
  assign _T_55060 = _T_55059[4:0]; // @[Modules.scala 46:37:@842.4]
  assign _T_55061 = $signed(_T_55060); // @[Modules.scala 46:37:@843.4]
  assign _T_55062 = $signed(_T_55061) - $signed(io_in_273); // @[Modules.scala 46:47:@844.4]
  assign _T_55063 = _T_55062[4:0]; // @[Modules.scala 46:47:@845.4]
  assign _T_55064 = $signed(_T_55063); // @[Modules.scala 46:47:@846.4]
  assign _T_55066 = $signed(5'sh0) - $signed(io_in_274); // @[Modules.scala 46:37:@848.4]
  assign _T_55067 = _T_55066[4:0]; // @[Modules.scala 46:37:@849.4]
  assign _T_55068 = $signed(_T_55067); // @[Modules.scala 46:37:@850.4]
  assign _T_55069 = $signed(_T_55068) - $signed(io_in_275); // @[Modules.scala 46:47:@851.4]
  assign _T_55070 = _T_55069[4:0]; // @[Modules.scala 46:47:@852.4]
  assign _T_55071 = $signed(_T_55070); // @[Modules.scala 46:47:@853.4]
  assign _T_55073 = $signed(5'sh0) - $signed(io_in_276); // @[Modules.scala 46:37:@855.4]
  assign _T_55074 = _T_55073[4:0]; // @[Modules.scala 46:37:@856.4]
  assign _T_55075 = $signed(_T_55074); // @[Modules.scala 46:37:@857.4]
  assign _T_55076 = $signed(_T_55075) - $signed(io_in_277); // @[Modules.scala 46:47:@858.4]
  assign _T_55077 = _T_55076[4:0]; // @[Modules.scala 46:47:@859.4]
  assign _T_55078 = $signed(_T_55077); // @[Modules.scala 46:47:@860.4]
  assign _T_55080 = $signed(5'sh0) - $signed(io_in_278); // @[Modules.scala 46:37:@862.4]
  assign _T_55081 = _T_55080[4:0]; // @[Modules.scala 46:37:@863.4]
  assign _T_55082 = $signed(_T_55081); // @[Modules.scala 46:37:@864.4]
  assign _T_55083 = $signed(_T_55082) - $signed(io_in_279); // @[Modules.scala 46:47:@865.4]
  assign _T_55084 = _T_55083[4:0]; // @[Modules.scala 46:47:@866.4]
  assign _T_55085 = $signed(_T_55084); // @[Modules.scala 46:47:@867.4]
  assign _T_55087 = $signed(5'sh0) - $signed(io_in_280); // @[Modules.scala 46:37:@869.4]
  assign _T_55088 = _T_55087[4:0]; // @[Modules.scala 46:37:@870.4]
  assign _T_55089 = $signed(_T_55088); // @[Modules.scala 46:37:@871.4]
  assign _T_55090 = $signed(_T_55089) - $signed(io_in_281); // @[Modules.scala 46:47:@872.4]
  assign _T_55091 = _T_55090[4:0]; // @[Modules.scala 46:47:@873.4]
  assign _T_55092 = $signed(_T_55091); // @[Modules.scala 46:47:@874.4]
  assign _T_55094 = $signed(5'sh0) - $signed(io_in_282); // @[Modules.scala 46:37:@876.4]
  assign _T_55095 = _T_55094[4:0]; // @[Modules.scala 46:37:@877.4]
  assign _T_55096 = $signed(_T_55095); // @[Modules.scala 46:37:@878.4]
  assign _T_55097 = $signed(_T_55096) - $signed(io_in_283); // @[Modules.scala 46:47:@879.4]
  assign _T_55098 = _T_55097[4:0]; // @[Modules.scala 46:47:@880.4]
  assign _T_55099 = $signed(_T_55098); // @[Modules.scala 46:47:@881.4]
  assign _T_55101 = $signed(5'sh0) - $signed(io_in_284); // @[Modules.scala 46:37:@883.4]
  assign _T_55102 = _T_55101[4:0]; // @[Modules.scala 46:37:@884.4]
  assign _T_55103 = $signed(_T_55102); // @[Modules.scala 46:37:@885.4]
  assign _T_55104 = $signed(_T_55103) - $signed(io_in_285); // @[Modules.scala 46:47:@886.4]
  assign _T_55105 = _T_55104[4:0]; // @[Modules.scala 46:47:@887.4]
  assign _T_55106 = $signed(_T_55105); // @[Modules.scala 46:47:@888.4]
  assign _T_55108 = $signed(5'sh0) - $signed(io_in_286); // @[Modules.scala 46:37:@890.4]
  assign _T_55109 = _T_55108[4:0]; // @[Modules.scala 46:37:@891.4]
  assign _T_55110 = $signed(_T_55109); // @[Modules.scala 46:37:@892.4]
  assign _T_55111 = $signed(_T_55110) - $signed(io_in_287); // @[Modules.scala 46:47:@893.4]
  assign _T_55112 = _T_55111[4:0]; // @[Modules.scala 46:47:@894.4]
  assign _T_55113 = $signed(_T_55112); // @[Modules.scala 46:47:@895.4]
  assign _T_55115 = $signed(5'sh0) - $signed(io_in_288); // @[Modules.scala 43:37:@897.4]
  assign _T_55116 = _T_55115[4:0]; // @[Modules.scala 43:37:@898.4]
  assign _T_55117 = $signed(_T_55116); // @[Modules.scala 43:37:@899.4]
  assign _T_55118 = $signed(_T_55117) + $signed(io_in_289); // @[Modules.scala 43:47:@900.4]
  assign _T_55119 = _T_55118[4:0]; // @[Modules.scala 43:47:@901.4]
  assign _T_55120 = $signed(_T_55119); // @[Modules.scala 43:47:@902.4]
  assign _T_55122 = $signed(5'sh0) - $signed(io_in_290); // @[Modules.scala 46:37:@904.4]
  assign _T_55123 = _T_55122[4:0]; // @[Modules.scala 46:37:@905.4]
  assign _T_55124 = $signed(_T_55123); // @[Modules.scala 46:37:@906.4]
  assign _T_55125 = $signed(_T_55124) - $signed(io_in_291); // @[Modules.scala 46:47:@907.4]
  assign _T_55126 = _T_55125[4:0]; // @[Modules.scala 46:47:@908.4]
  assign _T_55127 = $signed(_T_55126); // @[Modules.scala 46:47:@909.4]
  assign _T_55129 = $signed(5'sh0) - $signed(io_in_292); // @[Modules.scala 46:37:@911.4]
  assign _T_55130 = _T_55129[4:0]; // @[Modules.scala 46:37:@912.4]
  assign _T_55131 = $signed(_T_55130); // @[Modules.scala 46:37:@913.4]
  assign _T_55132 = $signed(_T_55131) - $signed(io_in_293); // @[Modules.scala 46:47:@914.4]
  assign _T_55133 = _T_55132[4:0]; // @[Modules.scala 46:47:@915.4]
  assign _T_55134 = $signed(_T_55133); // @[Modules.scala 46:47:@916.4]
  assign _T_55136 = $signed(5'sh0) - $signed(io_in_294); // @[Modules.scala 46:37:@918.4]
  assign _T_55137 = _T_55136[4:0]; // @[Modules.scala 46:37:@919.4]
  assign _T_55138 = $signed(_T_55137); // @[Modules.scala 46:37:@920.4]
  assign _T_55139 = $signed(_T_55138) - $signed(io_in_295); // @[Modules.scala 46:47:@921.4]
  assign _T_55140 = _T_55139[4:0]; // @[Modules.scala 46:47:@922.4]
  assign _T_55141 = $signed(_T_55140); // @[Modules.scala 46:47:@923.4]
  assign _T_55143 = $signed(5'sh0) - $signed(io_in_296); // @[Modules.scala 46:37:@925.4]
  assign _T_55144 = _T_55143[4:0]; // @[Modules.scala 46:37:@926.4]
  assign _T_55145 = $signed(_T_55144); // @[Modules.scala 46:37:@927.4]
  assign _T_55146 = $signed(_T_55145) - $signed(io_in_297); // @[Modules.scala 46:47:@928.4]
  assign _T_55147 = _T_55146[4:0]; // @[Modules.scala 46:47:@929.4]
  assign _T_55148 = $signed(_T_55147); // @[Modules.scala 46:47:@930.4]
  assign _T_55150 = $signed(5'sh0) - $signed(io_in_298); // @[Modules.scala 46:37:@932.4]
  assign _T_55151 = _T_55150[4:0]; // @[Modules.scala 46:37:@933.4]
  assign _T_55152 = $signed(_T_55151); // @[Modules.scala 46:37:@934.4]
  assign _T_55153 = $signed(_T_55152) - $signed(io_in_299); // @[Modules.scala 46:47:@935.4]
  assign _T_55154 = _T_55153[4:0]; // @[Modules.scala 46:47:@936.4]
  assign _T_55155 = $signed(_T_55154); // @[Modules.scala 46:47:@937.4]
  assign _T_55157 = $signed(5'sh0) - $signed(io_in_300); // @[Modules.scala 46:37:@939.4]
  assign _T_55158 = _T_55157[4:0]; // @[Modules.scala 46:37:@940.4]
  assign _T_55159 = $signed(_T_55158); // @[Modules.scala 46:37:@941.4]
  assign _T_55160 = $signed(_T_55159) - $signed(io_in_301); // @[Modules.scala 46:47:@942.4]
  assign _T_55161 = _T_55160[4:0]; // @[Modules.scala 46:47:@943.4]
  assign _T_55162 = $signed(_T_55161); // @[Modules.scala 46:47:@944.4]
  assign _T_55164 = $signed(5'sh0) - $signed(io_in_302); // @[Modules.scala 46:37:@946.4]
  assign _T_55165 = _T_55164[4:0]; // @[Modules.scala 46:37:@947.4]
  assign _T_55166 = $signed(_T_55165); // @[Modules.scala 46:37:@948.4]
  assign _T_55167 = $signed(_T_55166) - $signed(io_in_303); // @[Modules.scala 46:47:@949.4]
  assign _T_55168 = _T_55167[4:0]; // @[Modules.scala 46:47:@950.4]
  assign _T_55169 = $signed(_T_55168); // @[Modules.scala 46:47:@951.4]
  assign _T_55171 = $signed(5'sh0) - $signed(io_in_304); // @[Modules.scala 46:37:@953.4]
  assign _T_55172 = _T_55171[4:0]; // @[Modules.scala 46:37:@954.4]
  assign _T_55173 = $signed(_T_55172); // @[Modules.scala 46:37:@955.4]
  assign _T_55174 = $signed(_T_55173) - $signed(io_in_305); // @[Modules.scala 46:47:@956.4]
  assign _T_55175 = _T_55174[4:0]; // @[Modules.scala 46:47:@957.4]
  assign _T_55176 = $signed(_T_55175); // @[Modules.scala 46:47:@958.4]
  assign _T_55178 = $signed(5'sh0) - $signed(io_in_306); // @[Modules.scala 46:37:@960.4]
  assign _T_55179 = _T_55178[4:0]; // @[Modules.scala 46:37:@961.4]
  assign _T_55180 = $signed(_T_55179); // @[Modules.scala 46:37:@962.4]
  assign _T_55181 = $signed(_T_55180) - $signed(io_in_307); // @[Modules.scala 46:47:@963.4]
  assign _T_55182 = _T_55181[4:0]; // @[Modules.scala 46:47:@964.4]
  assign _T_55183 = $signed(_T_55182); // @[Modules.scala 46:47:@965.4]
  assign _T_55185 = $signed(5'sh0) - $signed(io_in_308); // @[Modules.scala 46:37:@967.4]
  assign _T_55186 = _T_55185[4:0]; // @[Modules.scala 46:37:@968.4]
  assign _T_55187 = $signed(_T_55186); // @[Modules.scala 46:37:@969.4]
  assign _T_55188 = $signed(_T_55187) - $signed(io_in_309); // @[Modules.scala 46:47:@970.4]
  assign _T_55189 = _T_55188[4:0]; // @[Modules.scala 46:47:@971.4]
  assign _T_55190 = $signed(_T_55189); // @[Modules.scala 46:47:@972.4]
  assign _T_55192 = $signed(5'sh0) - $signed(io_in_310); // @[Modules.scala 46:37:@974.4]
  assign _T_55193 = _T_55192[4:0]; // @[Modules.scala 46:37:@975.4]
  assign _T_55194 = $signed(_T_55193); // @[Modules.scala 46:37:@976.4]
  assign _T_55195 = $signed(_T_55194) - $signed(io_in_311); // @[Modules.scala 46:47:@977.4]
  assign _T_55196 = _T_55195[4:0]; // @[Modules.scala 46:47:@978.4]
  assign _T_55197 = $signed(_T_55196); // @[Modules.scala 46:47:@979.4]
  assign _T_55199 = $signed(5'sh0) - $signed(io_in_312); // @[Modules.scala 46:37:@981.4]
  assign _T_55200 = _T_55199[4:0]; // @[Modules.scala 46:37:@982.4]
  assign _T_55201 = $signed(_T_55200); // @[Modules.scala 46:37:@983.4]
  assign _T_55202 = $signed(_T_55201) - $signed(io_in_313); // @[Modules.scala 46:47:@984.4]
  assign _T_55203 = _T_55202[4:0]; // @[Modules.scala 46:47:@985.4]
  assign _T_55204 = $signed(_T_55203); // @[Modules.scala 46:47:@986.4]
  assign _T_55206 = $signed(5'sh0) - $signed(io_in_314); // @[Modules.scala 43:37:@988.4]
  assign _T_55207 = _T_55206[4:0]; // @[Modules.scala 43:37:@989.4]
  assign _T_55208 = $signed(_T_55207); // @[Modules.scala 43:37:@990.4]
  assign _T_55209 = $signed(_T_55208) + $signed(io_in_315); // @[Modules.scala 43:47:@991.4]
  assign _T_55210 = _T_55209[4:0]; // @[Modules.scala 43:47:@992.4]
  assign _T_55211 = $signed(_T_55210); // @[Modules.scala 43:47:@993.4]
  assign _T_55212 = $signed(io_in_316) + $signed(io_in_317); // @[Modules.scala 37:46:@995.4]
  assign _T_55213 = _T_55212[4:0]; // @[Modules.scala 37:46:@996.4]
  assign _T_55214 = $signed(_T_55213); // @[Modules.scala 37:46:@997.4]
  assign _T_55215 = $signed(io_in_318) + $signed(io_in_319); // @[Modules.scala 37:46:@999.4]
  assign _T_55216 = _T_55215[4:0]; // @[Modules.scala 37:46:@1000.4]
  assign _T_55217 = $signed(_T_55216); // @[Modules.scala 37:46:@1001.4]
  assign _T_55219 = $signed(5'sh0) - $signed(io_in_320); // @[Modules.scala 46:37:@1003.4]
  assign _T_55220 = _T_55219[4:0]; // @[Modules.scala 46:37:@1004.4]
  assign _T_55221 = $signed(_T_55220); // @[Modules.scala 46:37:@1005.4]
  assign _T_55222 = $signed(_T_55221) - $signed(io_in_321); // @[Modules.scala 46:47:@1006.4]
  assign _T_55223 = _T_55222[4:0]; // @[Modules.scala 46:47:@1007.4]
  assign _T_55224 = $signed(_T_55223); // @[Modules.scala 46:47:@1008.4]
  assign _T_55226 = $signed(5'sh0) - $signed(io_in_322); // @[Modules.scala 46:37:@1010.4]
  assign _T_55227 = _T_55226[4:0]; // @[Modules.scala 46:37:@1011.4]
  assign _T_55228 = $signed(_T_55227); // @[Modules.scala 46:37:@1012.4]
  assign _T_55229 = $signed(_T_55228) - $signed(io_in_323); // @[Modules.scala 46:47:@1013.4]
  assign _T_55230 = _T_55229[4:0]; // @[Modules.scala 46:47:@1014.4]
  assign _T_55231 = $signed(_T_55230); // @[Modules.scala 46:47:@1015.4]
  assign _T_55233 = $signed(5'sh0) - $signed(io_in_324); // @[Modules.scala 43:37:@1017.4]
  assign _T_55234 = _T_55233[4:0]; // @[Modules.scala 43:37:@1018.4]
  assign _T_55235 = $signed(_T_55234); // @[Modules.scala 43:37:@1019.4]
  assign _T_55236 = $signed(_T_55235) + $signed(io_in_325); // @[Modules.scala 43:47:@1020.4]
  assign _T_55237 = _T_55236[4:0]; // @[Modules.scala 43:47:@1021.4]
  assign _T_55238 = $signed(_T_55237); // @[Modules.scala 43:47:@1022.4]
  assign _T_55240 = $signed(5'sh0) - $signed(io_in_326); // @[Modules.scala 46:37:@1024.4]
  assign _T_55241 = _T_55240[4:0]; // @[Modules.scala 46:37:@1025.4]
  assign _T_55242 = $signed(_T_55241); // @[Modules.scala 46:37:@1026.4]
  assign _T_55243 = $signed(_T_55242) - $signed(io_in_327); // @[Modules.scala 46:47:@1027.4]
  assign _T_55244 = _T_55243[4:0]; // @[Modules.scala 46:47:@1028.4]
  assign _T_55245 = $signed(_T_55244); // @[Modules.scala 46:47:@1029.4]
  assign _T_55246 = $signed(io_in_328) + $signed(io_in_329); // @[Modules.scala 37:46:@1031.4]
  assign _T_55247 = _T_55246[4:0]; // @[Modules.scala 37:46:@1032.4]
  assign _T_55248 = $signed(_T_55247); // @[Modules.scala 37:46:@1033.4]
  assign _T_55250 = $signed(5'sh0) - $signed(io_in_330); // @[Modules.scala 46:37:@1035.4]
  assign _T_55251 = _T_55250[4:0]; // @[Modules.scala 46:37:@1036.4]
  assign _T_55252 = $signed(_T_55251); // @[Modules.scala 46:37:@1037.4]
  assign _T_55253 = $signed(_T_55252) - $signed(io_in_331); // @[Modules.scala 46:47:@1038.4]
  assign _T_55254 = _T_55253[4:0]; // @[Modules.scala 46:47:@1039.4]
  assign _T_55255 = $signed(_T_55254); // @[Modules.scala 46:47:@1040.4]
  assign _T_55257 = $signed(5'sh0) - $signed(io_in_332); // @[Modules.scala 46:37:@1042.4]
  assign _T_55258 = _T_55257[4:0]; // @[Modules.scala 46:37:@1043.4]
  assign _T_55259 = $signed(_T_55258); // @[Modules.scala 46:37:@1044.4]
  assign _T_55260 = $signed(_T_55259) - $signed(io_in_333); // @[Modules.scala 46:47:@1045.4]
  assign _T_55261 = _T_55260[4:0]; // @[Modules.scala 46:47:@1046.4]
  assign _T_55262 = $signed(_T_55261); // @[Modules.scala 46:47:@1047.4]
  assign _T_55264 = $signed(5'sh0) - $signed(io_in_334); // @[Modules.scala 43:37:@1049.4]
  assign _T_55265 = _T_55264[4:0]; // @[Modules.scala 43:37:@1050.4]
  assign _T_55266 = $signed(_T_55265); // @[Modules.scala 43:37:@1051.4]
  assign _T_55267 = $signed(_T_55266) + $signed(io_in_335); // @[Modules.scala 43:47:@1052.4]
  assign _T_55268 = _T_55267[4:0]; // @[Modules.scala 43:47:@1053.4]
  assign _T_55269 = $signed(_T_55268); // @[Modules.scala 43:47:@1054.4]
  assign _T_55270 = $signed(io_in_336) - $signed(io_in_337); // @[Modules.scala 40:46:@1056.4]
  assign _T_55271 = _T_55270[4:0]; // @[Modules.scala 40:46:@1057.4]
  assign _T_55272 = $signed(_T_55271); // @[Modules.scala 40:46:@1058.4]
  assign _T_55274 = $signed(5'sh0) - $signed(io_in_338); // @[Modules.scala 46:37:@1060.4]
  assign _T_55275 = _T_55274[4:0]; // @[Modules.scala 46:37:@1061.4]
  assign _T_55276 = $signed(_T_55275); // @[Modules.scala 46:37:@1062.4]
  assign _T_55277 = $signed(_T_55276) - $signed(io_in_339); // @[Modules.scala 46:47:@1063.4]
  assign _T_55278 = _T_55277[4:0]; // @[Modules.scala 46:47:@1064.4]
  assign _T_55279 = $signed(_T_55278); // @[Modules.scala 46:47:@1065.4]
  assign _T_55281 = $signed(5'sh0) - $signed(io_in_340); // @[Modules.scala 43:37:@1067.4]
  assign _T_55282 = _T_55281[4:0]; // @[Modules.scala 43:37:@1068.4]
  assign _T_55283 = $signed(_T_55282); // @[Modules.scala 43:37:@1069.4]
  assign _T_55284 = $signed(_T_55283) + $signed(io_in_341); // @[Modules.scala 43:47:@1070.4]
  assign _T_55285 = _T_55284[4:0]; // @[Modules.scala 43:47:@1071.4]
  assign _T_55286 = $signed(_T_55285); // @[Modules.scala 43:47:@1072.4]
  assign _T_55287 = $signed(io_in_342) + $signed(io_in_343); // @[Modules.scala 37:46:@1074.4]
  assign _T_55288 = _T_55287[4:0]; // @[Modules.scala 37:46:@1075.4]
  assign _T_55289 = $signed(_T_55288); // @[Modules.scala 37:46:@1076.4]
  assign _T_55290 = $signed(io_in_344) + $signed(io_in_345); // @[Modules.scala 37:46:@1078.4]
  assign _T_55291 = _T_55290[4:0]; // @[Modules.scala 37:46:@1079.4]
  assign _T_55292 = $signed(_T_55291); // @[Modules.scala 37:46:@1080.4]
  assign _T_55293 = $signed(io_in_346) + $signed(io_in_347); // @[Modules.scala 37:46:@1082.4]
  assign _T_55294 = _T_55293[4:0]; // @[Modules.scala 37:46:@1083.4]
  assign _T_55295 = $signed(_T_55294); // @[Modules.scala 37:46:@1084.4]
  assign _T_55296 = $signed(io_in_348) + $signed(io_in_349); // @[Modules.scala 37:46:@1086.4]
  assign _T_55297 = _T_55296[4:0]; // @[Modules.scala 37:46:@1087.4]
  assign _T_55298 = $signed(_T_55297); // @[Modules.scala 37:46:@1088.4]
  assign _T_55299 = $signed(io_in_350) + $signed(io_in_351); // @[Modules.scala 37:46:@1090.4]
  assign _T_55300 = _T_55299[4:0]; // @[Modules.scala 37:46:@1091.4]
  assign _T_55301 = $signed(_T_55300); // @[Modules.scala 37:46:@1092.4]
  assign _T_55302 = $signed(io_in_352) + $signed(io_in_353); // @[Modules.scala 37:46:@1094.4]
  assign _T_55303 = _T_55302[4:0]; // @[Modules.scala 37:46:@1095.4]
  assign _T_55304 = $signed(_T_55303); // @[Modules.scala 37:46:@1096.4]
  assign _T_55305 = $signed(io_in_354) + $signed(io_in_355); // @[Modules.scala 37:46:@1098.4]
  assign _T_55306 = _T_55305[4:0]; // @[Modules.scala 37:46:@1099.4]
  assign _T_55307 = $signed(_T_55306); // @[Modules.scala 37:46:@1100.4]
  assign _T_55308 = $signed(io_in_356) + $signed(io_in_357); // @[Modules.scala 37:46:@1102.4]
  assign _T_55309 = _T_55308[4:0]; // @[Modules.scala 37:46:@1103.4]
  assign _T_55310 = $signed(_T_55309); // @[Modules.scala 37:46:@1104.4]
  assign _T_55311 = $signed(io_in_358) + $signed(io_in_359); // @[Modules.scala 37:46:@1106.4]
  assign _T_55312 = _T_55311[4:0]; // @[Modules.scala 37:46:@1107.4]
  assign _T_55313 = $signed(_T_55312); // @[Modules.scala 37:46:@1108.4]
  assign _T_55315 = $signed(5'sh0) - $signed(io_in_360); // @[Modules.scala 46:37:@1110.4]
  assign _T_55316 = _T_55315[4:0]; // @[Modules.scala 46:37:@1111.4]
  assign _T_55317 = $signed(_T_55316); // @[Modules.scala 46:37:@1112.4]
  assign _T_55318 = $signed(_T_55317) - $signed(io_in_361); // @[Modules.scala 46:47:@1113.4]
  assign _T_55319 = _T_55318[4:0]; // @[Modules.scala 46:47:@1114.4]
  assign _T_55320 = $signed(_T_55319); // @[Modules.scala 46:47:@1115.4]
  assign _T_55322 = $signed(5'sh0) - $signed(io_in_362); // @[Modules.scala 43:37:@1117.4]
  assign _T_55323 = _T_55322[4:0]; // @[Modules.scala 43:37:@1118.4]
  assign _T_55324 = $signed(_T_55323); // @[Modules.scala 43:37:@1119.4]
  assign _T_55325 = $signed(_T_55324) + $signed(io_in_363); // @[Modules.scala 43:47:@1120.4]
  assign _T_55326 = _T_55325[4:0]; // @[Modules.scala 43:47:@1121.4]
  assign _T_55327 = $signed(_T_55326); // @[Modules.scala 43:47:@1122.4]
  assign _T_55329 = $signed(5'sh0) - $signed(io_in_364); // @[Modules.scala 46:37:@1124.4]
  assign _T_55330 = _T_55329[4:0]; // @[Modules.scala 46:37:@1125.4]
  assign _T_55331 = $signed(_T_55330); // @[Modules.scala 46:37:@1126.4]
  assign _T_55332 = $signed(_T_55331) - $signed(io_in_365); // @[Modules.scala 46:47:@1127.4]
  assign _T_55333 = _T_55332[4:0]; // @[Modules.scala 46:47:@1128.4]
  assign _T_55334 = $signed(_T_55333); // @[Modules.scala 46:47:@1129.4]
  assign _T_55336 = $signed(5'sh0) - $signed(io_in_366); // @[Modules.scala 46:37:@1131.4]
  assign _T_55337 = _T_55336[4:0]; // @[Modules.scala 46:37:@1132.4]
  assign _T_55338 = $signed(_T_55337); // @[Modules.scala 46:37:@1133.4]
  assign _T_55339 = $signed(_T_55338) - $signed(io_in_367); // @[Modules.scala 46:47:@1134.4]
  assign _T_55340 = _T_55339[4:0]; // @[Modules.scala 46:47:@1135.4]
  assign _T_55341 = $signed(_T_55340); // @[Modules.scala 46:47:@1136.4]
  assign _T_55342 = $signed(io_in_368) + $signed(io_in_369); // @[Modules.scala 37:46:@1138.4]
  assign _T_55343 = _T_55342[4:0]; // @[Modules.scala 37:46:@1139.4]
  assign _T_55344 = $signed(_T_55343); // @[Modules.scala 37:46:@1140.4]
  assign _T_55345 = $signed(io_in_370) + $signed(io_in_371); // @[Modules.scala 37:46:@1142.4]
  assign _T_55346 = _T_55345[4:0]; // @[Modules.scala 37:46:@1143.4]
  assign _T_55347 = $signed(_T_55346); // @[Modules.scala 37:46:@1144.4]
  assign _T_55348 = $signed(io_in_372) + $signed(io_in_373); // @[Modules.scala 37:46:@1146.4]
  assign _T_55349 = _T_55348[4:0]; // @[Modules.scala 37:46:@1147.4]
  assign _T_55350 = $signed(_T_55349); // @[Modules.scala 37:46:@1148.4]
  assign _T_55351 = $signed(io_in_374) + $signed(io_in_375); // @[Modules.scala 37:46:@1150.4]
  assign _T_55352 = _T_55351[4:0]; // @[Modules.scala 37:46:@1151.4]
  assign _T_55353 = $signed(_T_55352); // @[Modules.scala 37:46:@1152.4]
  assign _T_55354 = $signed(io_in_376) + $signed(io_in_377); // @[Modules.scala 37:46:@1154.4]
  assign _T_55355 = _T_55354[4:0]; // @[Modules.scala 37:46:@1155.4]
  assign _T_55356 = $signed(_T_55355); // @[Modules.scala 37:46:@1156.4]
  assign _T_55357 = $signed(io_in_378) + $signed(io_in_379); // @[Modules.scala 37:46:@1158.4]
  assign _T_55358 = _T_55357[4:0]; // @[Modules.scala 37:46:@1159.4]
  assign _T_55359 = $signed(_T_55358); // @[Modules.scala 37:46:@1160.4]
  assign _T_55360 = $signed(io_in_380) + $signed(io_in_381); // @[Modules.scala 37:46:@1162.4]
  assign _T_55361 = _T_55360[4:0]; // @[Modules.scala 37:46:@1163.4]
  assign _T_55362 = $signed(_T_55361); // @[Modules.scala 37:46:@1164.4]
  assign _T_55363 = $signed(io_in_382) + $signed(io_in_383); // @[Modules.scala 37:46:@1166.4]
  assign _T_55364 = _T_55363[4:0]; // @[Modules.scala 37:46:@1167.4]
  assign _T_55365 = $signed(_T_55364); // @[Modules.scala 37:46:@1168.4]
  assign _T_55367 = $signed(5'sh0) - $signed(io_in_384); // @[Modules.scala 43:37:@1170.4]
  assign _T_55368 = _T_55367[4:0]; // @[Modules.scala 43:37:@1171.4]
  assign _T_55369 = $signed(_T_55368); // @[Modules.scala 43:37:@1172.4]
  assign _T_55370 = $signed(_T_55369) + $signed(io_in_385); // @[Modules.scala 43:47:@1173.4]
  assign _T_55371 = _T_55370[4:0]; // @[Modules.scala 43:47:@1174.4]
  assign _T_55372 = $signed(_T_55371); // @[Modules.scala 43:47:@1175.4]
  assign _T_55373 = $signed(io_in_386) + $signed(io_in_387); // @[Modules.scala 37:46:@1177.4]
  assign _T_55374 = _T_55373[4:0]; // @[Modules.scala 37:46:@1178.4]
  assign _T_55375 = $signed(_T_55374); // @[Modules.scala 37:46:@1179.4]
  assign _T_55376 = $signed(io_in_388) - $signed(io_in_389); // @[Modules.scala 40:46:@1181.4]
  assign _T_55377 = _T_55376[4:0]; // @[Modules.scala 40:46:@1182.4]
  assign _T_55378 = $signed(_T_55377); // @[Modules.scala 40:46:@1183.4]
  assign _T_55380 = $signed(5'sh0) - $signed(io_in_390); // @[Modules.scala 43:37:@1185.4]
  assign _T_55381 = _T_55380[4:0]; // @[Modules.scala 43:37:@1186.4]
  assign _T_55382 = $signed(_T_55381); // @[Modules.scala 43:37:@1187.4]
  assign _T_55383 = $signed(_T_55382) + $signed(io_in_391); // @[Modules.scala 43:47:@1188.4]
  assign _T_55384 = _T_55383[4:0]; // @[Modules.scala 43:47:@1189.4]
  assign _T_55385 = $signed(_T_55384); // @[Modules.scala 43:47:@1190.4]
  assign _T_55387 = $signed(5'sh0) - $signed(io_in_392); // @[Modules.scala 46:37:@1192.4]
  assign _T_55388 = _T_55387[4:0]; // @[Modules.scala 46:37:@1193.4]
  assign _T_55389 = $signed(_T_55388); // @[Modules.scala 46:37:@1194.4]
  assign _T_55390 = $signed(_T_55389) - $signed(io_in_393); // @[Modules.scala 46:47:@1195.4]
  assign _T_55391 = _T_55390[4:0]; // @[Modules.scala 46:47:@1196.4]
  assign _T_55392 = $signed(_T_55391); // @[Modules.scala 46:47:@1197.4]
  assign _T_55394 = $signed(5'sh0) - $signed(io_in_394); // @[Modules.scala 46:37:@1199.4]
  assign _T_55395 = _T_55394[4:0]; // @[Modules.scala 46:37:@1200.4]
  assign _T_55396 = $signed(_T_55395); // @[Modules.scala 46:37:@1201.4]
  assign _T_55397 = $signed(_T_55396) - $signed(io_in_395); // @[Modules.scala 46:47:@1202.4]
  assign _T_55398 = _T_55397[4:0]; // @[Modules.scala 46:47:@1203.4]
  assign _T_55399 = $signed(_T_55398); // @[Modules.scala 46:47:@1204.4]
  assign _T_55400 = $signed(io_in_396) + $signed(io_in_397); // @[Modules.scala 37:46:@1206.4]
  assign _T_55401 = _T_55400[4:0]; // @[Modules.scala 37:46:@1207.4]
  assign _T_55402 = $signed(_T_55401); // @[Modules.scala 37:46:@1208.4]
  assign _T_55403 = $signed(io_in_398) + $signed(io_in_399); // @[Modules.scala 37:46:@1210.4]
  assign _T_55404 = _T_55403[4:0]; // @[Modules.scala 37:46:@1211.4]
  assign _T_55405 = $signed(_T_55404); // @[Modules.scala 37:46:@1212.4]
  assign _T_55406 = $signed(io_in_400) + $signed(io_in_401); // @[Modules.scala 37:46:@1214.4]
  assign _T_55407 = _T_55406[4:0]; // @[Modules.scala 37:46:@1215.4]
  assign _T_55408 = $signed(_T_55407); // @[Modules.scala 37:46:@1216.4]
  assign _T_55409 = $signed(io_in_402) + $signed(io_in_403); // @[Modules.scala 37:46:@1218.4]
  assign _T_55410 = _T_55409[4:0]; // @[Modules.scala 37:46:@1219.4]
  assign _T_55411 = $signed(_T_55410); // @[Modules.scala 37:46:@1220.4]
  assign _T_55412 = $signed(io_in_404) + $signed(io_in_405); // @[Modules.scala 37:46:@1222.4]
  assign _T_55413 = _T_55412[4:0]; // @[Modules.scala 37:46:@1223.4]
  assign _T_55414 = $signed(_T_55413); // @[Modules.scala 37:46:@1224.4]
  assign _T_55415 = $signed(io_in_406) + $signed(io_in_407); // @[Modules.scala 37:46:@1226.4]
  assign _T_55416 = _T_55415[4:0]; // @[Modules.scala 37:46:@1227.4]
  assign _T_55417 = $signed(_T_55416); // @[Modules.scala 37:46:@1228.4]
  assign _T_55418 = $signed(io_in_408) + $signed(io_in_409); // @[Modules.scala 37:46:@1230.4]
  assign _T_55419 = _T_55418[4:0]; // @[Modules.scala 37:46:@1231.4]
  assign _T_55420 = $signed(_T_55419); // @[Modules.scala 37:46:@1232.4]
  assign _T_55421 = $signed(io_in_410) + $signed(io_in_411); // @[Modules.scala 37:46:@1234.4]
  assign _T_55422 = _T_55421[4:0]; // @[Modules.scala 37:46:@1235.4]
  assign _T_55423 = $signed(_T_55422); // @[Modules.scala 37:46:@1236.4]
  assign _T_55424 = $signed(io_in_412) + $signed(io_in_413); // @[Modules.scala 37:46:@1238.4]
  assign _T_55425 = _T_55424[4:0]; // @[Modules.scala 37:46:@1239.4]
  assign _T_55426 = $signed(_T_55425); // @[Modules.scala 37:46:@1240.4]
  assign _T_55427 = $signed(io_in_414) + $signed(io_in_415); // @[Modules.scala 37:46:@1242.4]
  assign _T_55428 = _T_55427[4:0]; // @[Modules.scala 37:46:@1243.4]
  assign _T_55429 = $signed(_T_55428); // @[Modules.scala 37:46:@1244.4]
  assign _T_55430 = $signed(io_in_416) - $signed(io_in_417); // @[Modules.scala 40:46:@1246.4]
  assign _T_55431 = _T_55430[4:0]; // @[Modules.scala 40:46:@1247.4]
  assign _T_55432 = $signed(_T_55431); // @[Modules.scala 40:46:@1248.4]
  assign _T_55434 = $signed(5'sh0) - $signed(io_in_418); // @[Modules.scala 43:37:@1250.4]
  assign _T_55435 = _T_55434[4:0]; // @[Modules.scala 43:37:@1251.4]
  assign _T_55436 = $signed(_T_55435); // @[Modules.scala 43:37:@1252.4]
  assign _T_55437 = $signed(_T_55436) + $signed(io_in_419); // @[Modules.scala 43:47:@1253.4]
  assign _T_55438 = _T_55437[4:0]; // @[Modules.scala 43:47:@1254.4]
  assign _T_55439 = $signed(_T_55438); // @[Modules.scala 43:47:@1255.4]
  assign _T_55441 = $signed(5'sh0) - $signed(io_in_420); // @[Modules.scala 43:37:@1257.4]
  assign _T_55442 = _T_55441[4:0]; // @[Modules.scala 43:37:@1258.4]
  assign _T_55443 = $signed(_T_55442); // @[Modules.scala 43:37:@1259.4]
  assign _T_55444 = $signed(_T_55443) + $signed(io_in_421); // @[Modules.scala 43:47:@1260.4]
  assign _T_55445 = _T_55444[4:0]; // @[Modules.scala 43:47:@1261.4]
  assign _T_55446 = $signed(_T_55445); // @[Modules.scala 43:47:@1262.4]
  assign _T_55448 = $signed(5'sh0) - $signed(io_in_422); // @[Modules.scala 46:37:@1264.4]
  assign _T_55449 = _T_55448[4:0]; // @[Modules.scala 46:37:@1265.4]
  assign _T_55450 = $signed(_T_55449); // @[Modules.scala 46:37:@1266.4]
  assign _T_55451 = $signed(_T_55450) - $signed(io_in_423); // @[Modules.scala 46:47:@1267.4]
  assign _T_55452 = _T_55451[4:0]; // @[Modules.scala 46:47:@1268.4]
  assign _T_55453 = $signed(_T_55452); // @[Modules.scala 46:47:@1269.4]
  assign _T_55455 = $signed(5'sh0) - $signed(io_in_424); // @[Modules.scala 43:37:@1271.4]
  assign _T_55456 = _T_55455[4:0]; // @[Modules.scala 43:37:@1272.4]
  assign _T_55457 = $signed(_T_55456); // @[Modules.scala 43:37:@1273.4]
  assign _T_55458 = $signed(_T_55457) + $signed(io_in_425); // @[Modules.scala 43:47:@1274.4]
  assign _T_55459 = _T_55458[4:0]; // @[Modules.scala 43:47:@1275.4]
  assign _T_55460 = $signed(_T_55459); // @[Modules.scala 43:47:@1276.4]
  assign _T_55461 = $signed(io_in_426) + $signed(io_in_427); // @[Modules.scala 37:46:@1278.4]
  assign _T_55462 = _T_55461[4:0]; // @[Modules.scala 37:46:@1279.4]
  assign _T_55463 = $signed(_T_55462); // @[Modules.scala 37:46:@1280.4]
  assign _T_55464 = $signed(io_in_428) + $signed(io_in_429); // @[Modules.scala 37:46:@1282.4]
  assign _T_55465 = _T_55464[4:0]; // @[Modules.scala 37:46:@1283.4]
  assign _T_55466 = $signed(_T_55465); // @[Modules.scala 37:46:@1284.4]
  assign _T_55467 = $signed(io_in_430) + $signed(io_in_431); // @[Modules.scala 37:46:@1286.4]
  assign _T_55468 = _T_55467[4:0]; // @[Modules.scala 37:46:@1287.4]
  assign _T_55469 = $signed(_T_55468); // @[Modules.scala 37:46:@1288.4]
  assign _T_55470 = $signed(io_in_432) + $signed(io_in_433); // @[Modules.scala 37:46:@1290.4]
  assign _T_55471 = _T_55470[4:0]; // @[Modules.scala 37:46:@1291.4]
  assign _T_55472 = $signed(_T_55471); // @[Modules.scala 37:46:@1292.4]
  assign _T_55473 = $signed(io_in_434) + $signed(io_in_435); // @[Modules.scala 37:46:@1294.4]
  assign _T_55474 = _T_55473[4:0]; // @[Modules.scala 37:46:@1295.4]
  assign _T_55475 = $signed(_T_55474); // @[Modules.scala 37:46:@1296.4]
  assign _T_55476 = $signed(io_in_436) + $signed(io_in_437); // @[Modules.scala 37:46:@1298.4]
  assign _T_55477 = _T_55476[4:0]; // @[Modules.scala 37:46:@1299.4]
  assign _T_55478 = $signed(_T_55477); // @[Modules.scala 37:46:@1300.4]
  assign _T_55479 = $signed(io_in_438) - $signed(io_in_439); // @[Modules.scala 40:46:@1302.4]
  assign _T_55480 = _T_55479[4:0]; // @[Modules.scala 40:46:@1303.4]
  assign _T_55481 = $signed(_T_55480); // @[Modules.scala 40:46:@1304.4]
  assign _T_55482 = $signed(io_in_440) - $signed(io_in_441); // @[Modules.scala 40:46:@1306.4]
  assign _T_55483 = _T_55482[4:0]; // @[Modules.scala 40:46:@1307.4]
  assign _T_55484 = $signed(_T_55483); // @[Modules.scala 40:46:@1308.4]
  assign _T_55486 = $signed(5'sh0) - $signed(io_in_442); // @[Modules.scala 43:37:@1310.4]
  assign _T_55487 = _T_55486[4:0]; // @[Modules.scala 43:37:@1311.4]
  assign _T_55488 = $signed(_T_55487); // @[Modules.scala 43:37:@1312.4]
  assign _T_55489 = $signed(_T_55488) + $signed(io_in_443); // @[Modules.scala 43:47:@1313.4]
  assign _T_55490 = _T_55489[4:0]; // @[Modules.scala 43:47:@1314.4]
  assign _T_55491 = $signed(_T_55490); // @[Modules.scala 43:47:@1315.4]
  assign _T_55493 = $signed(5'sh0) - $signed(io_in_444); // @[Modules.scala 46:37:@1317.4]
  assign _T_55494 = _T_55493[4:0]; // @[Modules.scala 46:37:@1318.4]
  assign _T_55495 = $signed(_T_55494); // @[Modules.scala 46:37:@1319.4]
  assign _T_55496 = $signed(_T_55495) - $signed(io_in_445); // @[Modules.scala 46:47:@1320.4]
  assign _T_55497 = _T_55496[4:0]; // @[Modules.scala 46:47:@1321.4]
  assign _T_55498 = $signed(_T_55497); // @[Modules.scala 46:47:@1322.4]
  assign _T_55500 = $signed(5'sh0) - $signed(io_in_446); // @[Modules.scala 46:37:@1324.4]
  assign _T_55501 = _T_55500[4:0]; // @[Modules.scala 46:37:@1325.4]
  assign _T_55502 = $signed(_T_55501); // @[Modules.scala 46:37:@1326.4]
  assign _T_55503 = $signed(_T_55502) - $signed(io_in_447); // @[Modules.scala 46:47:@1327.4]
  assign _T_55504 = _T_55503[4:0]; // @[Modules.scala 46:47:@1328.4]
  assign _T_55505 = $signed(_T_55504); // @[Modules.scala 46:47:@1329.4]
  assign _T_55506 = $signed(io_in_448) + $signed(io_in_449); // @[Modules.scala 37:46:@1331.4]
  assign _T_55507 = _T_55506[4:0]; // @[Modules.scala 37:46:@1332.4]
  assign _T_55508 = $signed(_T_55507); // @[Modules.scala 37:46:@1333.4]
  assign _T_55510 = $signed(5'sh0) - $signed(io_in_450); // @[Modules.scala 46:37:@1335.4]
  assign _T_55511 = _T_55510[4:0]; // @[Modules.scala 46:37:@1336.4]
  assign _T_55512 = $signed(_T_55511); // @[Modules.scala 46:37:@1337.4]
  assign _T_55513 = $signed(_T_55512) - $signed(io_in_451); // @[Modules.scala 46:47:@1338.4]
  assign _T_55514 = _T_55513[4:0]; // @[Modules.scala 46:47:@1339.4]
  assign _T_55515 = $signed(_T_55514); // @[Modules.scala 46:47:@1340.4]
  assign _T_55517 = $signed(5'sh0) - $signed(io_in_452); // @[Modules.scala 43:37:@1342.4]
  assign _T_55518 = _T_55517[4:0]; // @[Modules.scala 43:37:@1343.4]
  assign _T_55519 = $signed(_T_55518); // @[Modules.scala 43:37:@1344.4]
  assign _T_55520 = $signed(_T_55519) + $signed(io_in_453); // @[Modules.scala 43:47:@1345.4]
  assign _T_55521 = _T_55520[4:0]; // @[Modules.scala 43:47:@1346.4]
  assign _T_55522 = $signed(_T_55521); // @[Modules.scala 43:47:@1347.4]
  assign _T_55523 = $signed(io_in_454) + $signed(io_in_455); // @[Modules.scala 37:46:@1349.4]
  assign _T_55524 = _T_55523[4:0]; // @[Modules.scala 37:46:@1350.4]
  assign _T_55525 = $signed(_T_55524); // @[Modules.scala 37:46:@1351.4]
  assign _T_55526 = $signed(io_in_456) + $signed(io_in_457); // @[Modules.scala 37:46:@1353.4]
  assign _T_55527 = _T_55526[4:0]; // @[Modules.scala 37:46:@1354.4]
  assign _T_55528 = $signed(_T_55527); // @[Modules.scala 37:46:@1355.4]
  assign _T_55529 = $signed(io_in_458) + $signed(io_in_459); // @[Modules.scala 37:46:@1357.4]
  assign _T_55530 = _T_55529[4:0]; // @[Modules.scala 37:46:@1358.4]
  assign _T_55531 = $signed(_T_55530); // @[Modules.scala 37:46:@1359.4]
  assign _T_55532 = $signed(io_in_460) - $signed(io_in_461); // @[Modules.scala 40:46:@1361.4]
  assign _T_55533 = _T_55532[4:0]; // @[Modules.scala 40:46:@1362.4]
  assign _T_55534 = $signed(_T_55533); // @[Modules.scala 40:46:@1363.4]
  assign _T_55535 = $signed(io_in_462) + $signed(io_in_463); // @[Modules.scala 37:46:@1365.4]
  assign _T_55536 = _T_55535[4:0]; // @[Modules.scala 37:46:@1366.4]
  assign _T_55537 = $signed(_T_55536); // @[Modules.scala 37:46:@1367.4]
  assign _T_55538 = $signed(io_in_464) + $signed(io_in_465); // @[Modules.scala 37:46:@1369.4]
  assign _T_55539 = _T_55538[4:0]; // @[Modules.scala 37:46:@1370.4]
  assign _T_55540 = $signed(_T_55539); // @[Modules.scala 37:46:@1371.4]
  assign _T_55541 = $signed(io_in_466) + $signed(io_in_467); // @[Modules.scala 37:46:@1373.4]
  assign _T_55542 = _T_55541[4:0]; // @[Modules.scala 37:46:@1374.4]
  assign _T_55543 = $signed(_T_55542); // @[Modules.scala 37:46:@1375.4]
  assign _T_55544 = $signed(io_in_468) - $signed(io_in_469); // @[Modules.scala 40:46:@1377.4]
  assign _T_55545 = _T_55544[4:0]; // @[Modules.scala 40:46:@1378.4]
  assign _T_55546 = $signed(_T_55545); // @[Modules.scala 40:46:@1379.4]
  assign _T_55548 = $signed(5'sh0) - $signed(io_in_470); // @[Modules.scala 46:37:@1381.4]
  assign _T_55549 = _T_55548[4:0]; // @[Modules.scala 46:37:@1382.4]
  assign _T_55550 = $signed(_T_55549); // @[Modules.scala 46:37:@1383.4]
  assign _T_55551 = $signed(_T_55550) - $signed(io_in_471); // @[Modules.scala 46:47:@1384.4]
  assign _T_55552 = _T_55551[4:0]; // @[Modules.scala 46:47:@1385.4]
  assign _T_55553 = $signed(_T_55552); // @[Modules.scala 46:47:@1386.4]
  assign _T_55555 = $signed(5'sh0) - $signed(io_in_472); // @[Modules.scala 46:37:@1388.4]
  assign _T_55556 = _T_55555[4:0]; // @[Modules.scala 46:37:@1389.4]
  assign _T_55557 = $signed(_T_55556); // @[Modules.scala 46:37:@1390.4]
  assign _T_55558 = $signed(_T_55557) - $signed(io_in_473); // @[Modules.scala 46:47:@1391.4]
  assign _T_55559 = _T_55558[4:0]; // @[Modules.scala 46:47:@1392.4]
  assign _T_55560 = $signed(_T_55559); // @[Modules.scala 46:47:@1393.4]
  assign _T_55562 = $signed(5'sh0) - $signed(io_in_474); // @[Modules.scala 46:37:@1395.4]
  assign _T_55563 = _T_55562[4:0]; // @[Modules.scala 46:37:@1396.4]
  assign _T_55564 = $signed(_T_55563); // @[Modules.scala 46:37:@1397.4]
  assign _T_55565 = $signed(_T_55564) - $signed(io_in_475); // @[Modules.scala 46:47:@1398.4]
  assign _T_55566 = _T_55565[4:0]; // @[Modules.scala 46:47:@1399.4]
  assign _T_55567 = $signed(_T_55566); // @[Modules.scala 46:47:@1400.4]
  assign _T_55569 = $signed(5'sh0) - $signed(io_in_476); // @[Modules.scala 46:37:@1402.4]
  assign _T_55570 = _T_55569[4:0]; // @[Modules.scala 46:37:@1403.4]
  assign _T_55571 = $signed(_T_55570); // @[Modules.scala 46:37:@1404.4]
  assign _T_55572 = $signed(_T_55571) - $signed(io_in_477); // @[Modules.scala 46:47:@1405.4]
  assign _T_55573 = _T_55572[4:0]; // @[Modules.scala 46:47:@1406.4]
  assign _T_55574 = $signed(_T_55573); // @[Modules.scala 46:47:@1407.4]
  assign _T_55575 = $signed(io_in_478) - $signed(io_in_479); // @[Modules.scala 40:46:@1409.4]
  assign _T_55576 = _T_55575[4:0]; // @[Modules.scala 40:46:@1410.4]
  assign _T_55577 = $signed(_T_55576); // @[Modules.scala 40:46:@1411.4]
  assign _T_55579 = $signed(5'sh0) - $signed(io_in_480); // @[Modules.scala 46:37:@1413.4]
  assign _T_55580 = _T_55579[4:0]; // @[Modules.scala 46:37:@1414.4]
  assign _T_55581 = $signed(_T_55580); // @[Modules.scala 46:37:@1415.4]
  assign _T_55582 = $signed(_T_55581) - $signed(io_in_481); // @[Modules.scala 46:47:@1416.4]
  assign _T_55583 = _T_55582[4:0]; // @[Modules.scala 46:47:@1417.4]
  assign _T_55584 = $signed(_T_55583); // @[Modules.scala 46:47:@1418.4]
  assign _T_55585 = $signed(io_in_482) + $signed(io_in_483); // @[Modules.scala 37:46:@1420.4]
  assign _T_55586 = _T_55585[4:0]; // @[Modules.scala 37:46:@1421.4]
  assign _T_55587 = $signed(_T_55586); // @[Modules.scala 37:46:@1422.4]
  assign _T_55588 = $signed(io_in_484) + $signed(io_in_485); // @[Modules.scala 37:46:@1424.4]
  assign _T_55589 = _T_55588[4:0]; // @[Modules.scala 37:46:@1425.4]
  assign _T_55590 = $signed(_T_55589); // @[Modules.scala 37:46:@1426.4]
  assign _T_55591 = $signed(io_in_486) + $signed(io_in_487); // @[Modules.scala 37:46:@1428.4]
  assign _T_55592 = _T_55591[4:0]; // @[Modules.scala 37:46:@1429.4]
  assign _T_55593 = $signed(_T_55592); // @[Modules.scala 37:46:@1430.4]
  assign _T_55595 = $signed(5'sh0) - $signed(io_in_488); // @[Modules.scala 43:37:@1432.4]
  assign _T_55596 = _T_55595[4:0]; // @[Modules.scala 43:37:@1433.4]
  assign _T_55597 = $signed(_T_55596); // @[Modules.scala 43:37:@1434.4]
  assign _T_55598 = $signed(_T_55597) + $signed(io_in_489); // @[Modules.scala 43:47:@1435.4]
  assign _T_55599 = _T_55598[4:0]; // @[Modules.scala 43:47:@1436.4]
  assign _T_55600 = $signed(_T_55599); // @[Modules.scala 43:47:@1437.4]
  assign _T_55601 = $signed(io_in_490) + $signed(io_in_491); // @[Modules.scala 37:46:@1439.4]
  assign _T_55602 = _T_55601[4:0]; // @[Modules.scala 37:46:@1440.4]
  assign _T_55603 = $signed(_T_55602); // @[Modules.scala 37:46:@1441.4]
  assign _T_55604 = $signed(io_in_492) - $signed(io_in_493); // @[Modules.scala 40:46:@1443.4]
  assign _T_55605 = _T_55604[4:0]; // @[Modules.scala 40:46:@1444.4]
  assign _T_55606 = $signed(_T_55605); // @[Modules.scala 40:46:@1445.4]
  assign _T_55607 = $signed(io_in_494) - $signed(io_in_495); // @[Modules.scala 40:46:@1447.4]
  assign _T_55608 = _T_55607[4:0]; // @[Modules.scala 40:46:@1448.4]
  assign _T_55609 = $signed(_T_55608); // @[Modules.scala 40:46:@1449.4]
  assign _T_55611 = $signed(5'sh0) - $signed(io_in_496); // @[Modules.scala 46:37:@1451.4]
  assign _T_55612 = _T_55611[4:0]; // @[Modules.scala 46:37:@1452.4]
  assign _T_55613 = $signed(_T_55612); // @[Modules.scala 46:37:@1453.4]
  assign _T_55614 = $signed(_T_55613) - $signed(io_in_497); // @[Modules.scala 46:47:@1454.4]
  assign _T_55615 = _T_55614[4:0]; // @[Modules.scala 46:47:@1455.4]
  assign _T_55616 = $signed(_T_55615); // @[Modules.scala 46:47:@1456.4]
  assign _T_55617 = $signed(io_in_498) + $signed(io_in_499); // @[Modules.scala 37:46:@1458.4]
  assign _T_55618 = _T_55617[4:0]; // @[Modules.scala 37:46:@1459.4]
  assign _T_55619 = $signed(_T_55618); // @[Modules.scala 37:46:@1460.4]
  assign _T_55621 = $signed(5'sh0) - $signed(io_in_500); // @[Modules.scala 46:37:@1462.4]
  assign _T_55622 = _T_55621[4:0]; // @[Modules.scala 46:37:@1463.4]
  assign _T_55623 = $signed(_T_55622); // @[Modules.scala 46:37:@1464.4]
  assign _T_55624 = $signed(_T_55623) - $signed(io_in_501); // @[Modules.scala 46:47:@1465.4]
  assign _T_55625 = _T_55624[4:0]; // @[Modules.scala 46:47:@1466.4]
  assign _T_55626 = $signed(_T_55625); // @[Modules.scala 46:47:@1467.4]
  assign _T_55628 = $signed(5'sh0) - $signed(io_in_502); // @[Modules.scala 46:37:@1469.4]
  assign _T_55629 = _T_55628[4:0]; // @[Modules.scala 46:37:@1470.4]
  assign _T_55630 = $signed(_T_55629); // @[Modules.scala 46:37:@1471.4]
  assign _T_55631 = $signed(_T_55630) - $signed(io_in_503); // @[Modules.scala 46:47:@1472.4]
  assign _T_55632 = _T_55631[4:0]; // @[Modules.scala 46:47:@1473.4]
  assign _T_55633 = $signed(_T_55632); // @[Modules.scala 46:47:@1474.4]
  assign _T_55635 = $signed(5'sh0) - $signed(io_in_504); // @[Modules.scala 46:37:@1476.4]
  assign _T_55636 = _T_55635[4:0]; // @[Modules.scala 46:37:@1477.4]
  assign _T_55637 = $signed(_T_55636); // @[Modules.scala 46:37:@1478.4]
  assign _T_55638 = $signed(_T_55637) - $signed(io_in_505); // @[Modules.scala 46:47:@1479.4]
  assign _T_55639 = _T_55638[4:0]; // @[Modules.scala 46:47:@1480.4]
  assign _T_55640 = $signed(_T_55639); // @[Modules.scala 46:47:@1481.4]
  assign _T_55642 = $signed(5'sh0) - $signed(io_in_506); // @[Modules.scala 43:37:@1483.4]
  assign _T_55643 = _T_55642[4:0]; // @[Modules.scala 43:37:@1484.4]
  assign _T_55644 = $signed(_T_55643); // @[Modules.scala 43:37:@1485.4]
  assign _T_55645 = $signed(_T_55644) + $signed(io_in_507); // @[Modules.scala 43:47:@1486.4]
  assign _T_55646 = _T_55645[4:0]; // @[Modules.scala 43:47:@1487.4]
  assign _T_55647 = $signed(_T_55646); // @[Modules.scala 43:47:@1488.4]
  assign _T_55649 = $signed(5'sh0) - $signed(io_in_508); // @[Modules.scala 46:37:@1490.4]
  assign _T_55650 = _T_55649[4:0]; // @[Modules.scala 46:37:@1491.4]
  assign _T_55651 = $signed(_T_55650); // @[Modules.scala 46:37:@1492.4]
  assign _T_55652 = $signed(_T_55651) - $signed(io_in_509); // @[Modules.scala 46:47:@1493.4]
  assign _T_55653 = _T_55652[4:0]; // @[Modules.scala 46:47:@1494.4]
  assign _T_55654 = $signed(_T_55653); // @[Modules.scala 46:47:@1495.4]
  assign _T_55656 = $signed(5'sh0) - $signed(io_in_510); // @[Modules.scala 46:37:@1497.4]
  assign _T_55657 = _T_55656[4:0]; // @[Modules.scala 46:37:@1498.4]
  assign _T_55658 = $signed(_T_55657); // @[Modules.scala 46:37:@1499.4]
  assign _T_55659 = $signed(_T_55658) - $signed(io_in_511); // @[Modules.scala 46:47:@1500.4]
  assign _T_55660 = _T_55659[4:0]; // @[Modules.scala 46:47:@1501.4]
  assign _T_55661 = $signed(_T_55660); // @[Modules.scala 46:47:@1502.4]
  assign _T_55662 = $signed(io_in_512) + $signed(io_in_513); // @[Modules.scala 37:46:@1504.4]
  assign _T_55663 = _T_55662[4:0]; // @[Modules.scala 37:46:@1505.4]
  assign _T_55664 = $signed(_T_55663); // @[Modules.scala 37:46:@1506.4]
  assign _T_55665 = $signed(io_in_514) + $signed(io_in_515); // @[Modules.scala 37:46:@1508.4]
  assign _T_55666 = _T_55665[4:0]; // @[Modules.scala 37:46:@1509.4]
  assign _T_55667 = $signed(_T_55666); // @[Modules.scala 37:46:@1510.4]
  assign _T_55668 = $signed(io_in_516) - $signed(io_in_517); // @[Modules.scala 40:46:@1512.4]
  assign _T_55669 = _T_55668[4:0]; // @[Modules.scala 40:46:@1513.4]
  assign _T_55670 = $signed(_T_55669); // @[Modules.scala 40:46:@1514.4]
  assign _T_55671 = $signed(io_in_518) + $signed(io_in_519); // @[Modules.scala 37:46:@1516.4]
  assign _T_55672 = _T_55671[4:0]; // @[Modules.scala 37:46:@1517.4]
  assign _T_55673 = $signed(_T_55672); // @[Modules.scala 37:46:@1518.4]
  assign _T_55675 = $signed(5'sh0) - $signed(io_in_520); // @[Modules.scala 43:37:@1520.4]
  assign _T_55676 = _T_55675[4:0]; // @[Modules.scala 43:37:@1521.4]
  assign _T_55677 = $signed(_T_55676); // @[Modules.scala 43:37:@1522.4]
  assign _T_55678 = $signed(_T_55677) + $signed(io_in_521); // @[Modules.scala 43:47:@1523.4]
  assign _T_55679 = _T_55678[4:0]; // @[Modules.scala 43:47:@1524.4]
  assign _T_55680 = $signed(_T_55679); // @[Modules.scala 43:47:@1525.4]
  assign _T_55682 = $signed(5'sh0) - $signed(io_in_522); // @[Modules.scala 43:37:@1527.4]
  assign _T_55683 = _T_55682[4:0]; // @[Modules.scala 43:37:@1528.4]
  assign _T_55684 = $signed(_T_55683); // @[Modules.scala 43:37:@1529.4]
  assign _T_55685 = $signed(_T_55684) + $signed(io_in_523); // @[Modules.scala 43:47:@1530.4]
  assign _T_55686 = _T_55685[4:0]; // @[Modules.scala 43:47:@1531.4]
  assign _T_55687 = $signed(_T_55686); // @[Modules.scala 43:47:@1532.4]
  assign _T_55689 = $signed(5'sh0) - $signed(io_in_524); // @[Modules.scala 43:37:@1534.4]
  assign _T_55690 = _T_55689[4:0]; // @[Modules.scala 43:37:@1535.4]
  assign _T_55691 = $signed(_T_55690); // @[Modules.scala 43:37:@1536.4]
  assign _T_55692 = $signed(_T_55691) + $signed(io_in_525); // @[Modules.scala 43:47:@1537.4]
  assign _T_55693 = _T_55692[4:0]; // @[Modules.scala 43:47:@1538.4]
  assign _T_55694 = $signed(_T_55693); // @[Modules.scala 43:47:@1539.4]
  assign _T_55695 = $signed(io_in_526) + $signed(io_in_527); // @[Modules.scala 37:46:@1541.4]
  assign _T_55696 = _T_55695[4:0]; // @[Modules.scala 37:46:@1542.4]
  assign _T_55697 = $signed(_T_55696); // @[Modules.scala 37:46:@1543.4]
  assign _T_55698 = $signed(io_in_528) + $signed(io_in_529); // @[Modules.scala 37:46:@1545.4]
  assign _T_55699 = _T_55698[4:0]; // @[Modules.scala 37:46:@1546.4]
  assign _T_55700 = $signed(_T_55699); // @[Modules.scala 37:46:@1547.4]
  assign _T_55702 = $signed(5'sh0) - $signed(io_in_530); // @[Modules.scala 46:37:@1549.4]
  assign _T_55703 = _T_55702[4:0]; // @[Modules.scala 46:37:@1550.4]
  assign _T_55704 = $signed(_T_55703); // @[Modules.scala 46:37:@1551.4]
  assign _T_55705 = $signed(_T_55704) - $signed(io_in_531); // @[Modules.scala 46:47:@1552.4]
  assign _T_55706 = _T_55705[4:0]; // @[Modules.scala 46:47:@1553.4]
  assign _T_55707 = $signed(_T_55706); // @[Modules.scala 46:47:@1554.4]
  assign _T_55708 = $signed(io_in_532) - $signed(io_in_533); // @[Modules.scala 40:46:@1556.4]
  assign _T_55709 = _T_55708[4:0]; // @[Modules.scala 40:46:@1557.4]
  assign _T_55710 = $signed(_T_55709); // @[Modules.scala 40:46:@1558.4]
  assign _T_55712 = $signed(5'sh0) - $signed(io_in_534); // @[Modules.scala 43:37:@1560.4]
  assign _T_55713 = _T_55712[4:0]; // @[Modules.scala 43:37:@1561.4]
  assign _T_55714 = $signed(_T_55713); // @[Modules.scala 43:37:@1562.4]
  assign _T_55715 = $signed(_T_55714) + $signed(io_in_535); // @[Modules.scala 43:47:@1563.4]
  assign _T_55716 = _T_55715[4:0]; // @[Modules.scala 43:47:@1564.4]
  assign _T_55717 = $signed(_T_55716); // @[Modules.scala 43:47:@1565.4]
  assign _T_55719 = $signed(5'sh0) - $signed(io_in_536); // @[Modules.scala 46:37:@1567.4]
  assign _T_55720 = _T_55719[4:0]; // @[Modules.scala 46:37:@1568.4]
  assign _T_55721 = $signed(_T_55720); // @[Modules.scala 46:37:@1569.4]
  assign _T_55722 = $signed(_T_55721) - $signed(io_in_537); // @[Modules.scala 46:47:@1570.4]
  assign _T_55723 = _T_55722[4:0]; // @[Modules.scala 46:47:@1571.4]
  assign _T_55724 = $signed(_T_55723); // @[Modules.scala 46:47:@1572.4]
  assign _T_55726 = $signed(5'sh0) - $signed(io_in_538); // @[Modules.scala 46:37:@1574.4]
  assign _T_55727 = _T_55726[4:0]; // @[Modules.scala 46:37:@1575.4]
  assign _T_55728 = $signed(_T_55727); // @[Modules.scala 46:37:@1576.4]
  assign _T_55729 = $signed(_T_55728) - $signed(io_in_539); // @[Modules.scala 46:47:@1577.4]
  assign _T_55730 = _T_55729[4:0]; // @[Modules.scala 46:47:@1578.4]
  assign _T_55731 = $signed(_T_55730); // @[Modules.scala 46:47:@1579.4]
  assign _T_55733 = $signed(5'sh0) - $signed(io_in_540); // @[Modules.scala 46:37:@1581.4]
  assign _T_55734 = _T_55733[4:0]; // @[Modules.scala 46:37:@1582.4]
  assign _T_55735 = $signed(_T_55734); // @[Modules.scala 46:37:@1583.4]
  assign _T_55736 = $signed(_T_55735) - $signed(io_in_541); // @[Modules.scala 46:47:@1584.4]
  assign _T_55737 = _T_55736[4:0]; // @[Modules.scala 46:47:@1585.4]
  assign _T_55738 = $signed(_T_55737); // @[Modules.scala 46:47:@1586.4]
  assign _T_55740 = $signed(5'sh0) - $signed(io_in_542); // @[Modules.scala 43:37:@1588.4]
  assign _T_55741 = _T_55740[4:0]; // @[Modules.scala 43:37:@1589.4]
  assign _T_55742 = $signed(_T_55741); // @[Modules.scala 43:37:@1590.4]
  assign _T_55743 = $signed(_T_55742) + $signed(io_in_543); // @[Modules.scala 43:47:@1591.4]
  assign _T_55744 = _T_55743[4:0]; // @[Modules.scala 43:47:@1592.4]
  assign _T_55745 = $signed(_T_55744); // @[Modules.scala 43:47:@1593.4]
  assign _T_55747 = $signed(5'sh0) - $signed(io_in_544); // @[Modules.scala 46:37:@1595.4]
  assign _T_55748 = _T_55747[4:0]; // @[Modules.scala 46:37:@1596.4]
  assign _T_55749 = $signed(_T_55748); // @[Modules.scala 46:37:@1597.4]
  assign _T_55750 = $signed(_T_55749) - $signed(io_in_545); // @[Modules.scala 46:47:@1598.4]
  assign _T_55751 = _T_55750[4:0]; // @[Modules.scala 46:47:@1599.4]
  assign _T_55752 = $signed(_T_55751); // @[Modules.scala 46:47:@1600.4]
  assign _T_55754 = $signed(5'sh0) - $signed(io_in_546); // @[Modules.scala 46:37:@1602.4]
  assign _T_55755 = _T_55754[4:0]; // @[Modules.scala 46:37:@1603.4]
  assign _T_55756 = $signed(_T_55755); // @[Modules.scala 46:37:@1604.4]
  assign _T_55757 = $signed(_T_55756) - $signed(io_in_547); // @[Modules.scala 46:47:@1605.4]
  assign _T_55758 = _T_55757[4:0]; // @[Modules.scala 46:47:@1606.4]
  assign _T_55759 = $signed(_T_55758); // @[Modules.scala 46:47:@1607.4]
  assign _T_55761 = $signed(5'sh0) - $signed(io_in_548); // @[Modules.scala 46:37:@1609.4]
  assign _T_55762 = _T_55761[4:0]; // @[Modules.scala 46:37:@1610.4]
  assign _T_55763 = $signed(_T_55762); // @[Modules.scala 46:37:@1611.4]
  assign _T_55764 = $signed(_T_55763) - $signed(io_in_549); // @[Modules.scala 46:47:@1612.4]
  assign _T_55765 = _T_55764[4:0]; // @[Modules.scala 46:47:@1613.4]
  assign _T_55766 = $signed(_T_55765); // @[Modules.scala 46:47:@1614.4]
  assign _T_55767 = $signed(io_in_550) - $signed(io_in_551); // @[Modules.scala 40:46:@1616.4]
  assign _T_55768 = _T_55767[4:0]; // @[Modules.scala 40:46:@1617.4]
  assign _T_55769 = $signed(_T_55768); // @[Modules.scala 40:46:@1618.4]
  assign _T_55770 = $signed(io_in_552) - $signed(io_in_553); // @[Modules.scala 40:46:@1620.4]
  assign _T_55771 = _T_55770[4:0]; // @[Modules.scala 40:46:@1621.4]
  assign _T_55772 = $signed(_T_55771); // @[Modules.scala 40:46:@1622.4]
  assign _T_55774 = $signed(5'sh0) - $signed(io_in_554); // @[Modules.scala 46:37:@1624.4]
  assign _T_55775 = _T_55774[4:0]; // @[Modules.scala 46:37:@1625.4]
  assign _T_55776 = $signed(_T_55775); // @[Modules.scala 46:37:@1626.4]
  assign _T_55777 = $signed(_T_55776) - $signed(io_in_555); // @[Modules.scala 46:47:@1627.4]
  assign _T_55778 = _T_55777[4:0]; // @[Modules.scala 46:47:@1628.4]
  assign _T_55779 = $signed(_T_55778); // @[Modules.scala 46:47:@1629.4]
  assign _T_55780 = $signed(io_in_556) - $signed(io_in_557); // @[Modules.scala 40:46:@1631.4]
  assign _T_55781 = _T_55780[4:0]; // @[Modules.scala 40:46:@1632.4]
  assign _T_55782 = $signed(_T_55781); // @[Modules.scala 40:46:@1633.4]
  assign _T_55784 = $signed(5'sh0) - $signed(io_in_558); // @[Modules.scala 43:37:@1635.4]
  assign _T_55785 = _T_55784[4:0]; // @[Modules.scala 43:37:@1636.4]
  assign _T_55786 = $signed(_T_55785); // @[Modules.scala 43:37:@1637.4]
  assign _T_55787 = $signed(_T_55786) + $signed(io_in_559); // @[Modules.scala 43:47:@1638.4]
  assign _T_55788 = _T_55787[4:0]; // @[Modules.scala 43:47:@1639.4]
  assign _T_55789 = $signed(_T_55788); // @[Modules.scala 43:47:@1640.4]
  assign _T_55791 = $signed(5'sh0) - $signed(io_in_560); // @[Modules.scala 46:37:@1642.4]
  assign _T_55792 = _T_55791[4:0]; // @[Modules.scala 46:37:@1643.4]
  assign _T_55793 = $signed(_T_55792); // @[Modules.scala 46:37:@1644.4]
  assign _T_55794 = $signed(_T_55793) - $signed(io_in_561); // @[Modules.scala 46:47:@1645.4]
  assign _T_55795 = _T_55794[4:0]; // @[Modules.scala 46:47:@1646.4]
  assign _T_55796 = $signed(_T_55795); // @[Modules.scala 46:47:@1647.4]
  assign _T_55798 = $signed(5'sh0) - $signed(io_in_562); // @[Modules.scala 46:37:@1649.4]
  assign _T_55799 = _T_55798[4:0]; // @[Modules.scala 46:37:@1650.4]
  assign _T_55800 = $signed(_T_55799); // @[Modules.scala 46:37:@1651.4]
  assign _T_55801 = $signed(_T_55800) - $signed(io_in_563); // @[Modules.scala 46:47:@1652.4]
  assign _T_55802 = _T_55801[4:0]; // @[Modules.scala 46:47:@1653.4]
  assign _T_55803 = $signed(_T_55802); // @[Modules.scala 46:47:@1654.4]
  assign _T_55805 = $signed(5'sh0) - $signed(io_in_564); // @[Modules.scala 46:37:@1656.4]
  assign _T_55806 = _T_55805[4:0]; // @[Modules.scala 46:37:@1657.4]
  assign _T_55807 = $signed(_T_55806); // @[Modules.scala 46:37:@1658.4]
  assign _T_55808 = $signed(_T_55807) - $signed(io_in_565); // @[Modules.scala 46:47:@1659.4]
  assign _T_55809 = _T_55808[4:0]; // @[Modules.scala 46:47:@1660.4]
  assign _T_55810 = $signed(_T_55809); // @[Modules.scala 46:47:@1661.4]
  assign _T_55812 = $signed(5'sh0) - $signed(io_in_566); // @[Modules.scala 46:37:@1663.4]
  assign _T_55813 = _T_55812[4:0]; // @[Modules.scala 46:37:@1664.4]
  assign _T_55814 = $signed(_T_55813); // @[Modules.scala 46:37:@1665.4]
  assign _T_55815 = $signed(_T_55814) - $signed(io_in_567); // @[Modules.scala 46:47:@1666.4]
  assign _T_55816 = _T_55815[4:0]; // @[Modules.scala 46:47:@1667.4]
  assign _T_55817 = $signed(_T_55816); // @[Modules.scala 46:47:@1668.4]
  assign _T_55819 = $signed(5'sh0) - $signed(io_in_568); // @[Modules.scala 46:37:@1670.4]
  assign _T_55820 = _T_55819[4:0]; // @[Modules.scala 46:37:@1671.4]
  assign _T_55821 = $signed(_T_55820); // @[Modules.scala 46:37:@1672.4]
  assign _T_55822 = $signed(_T_55821) - $signed(io_in_569); // @[Modules.scala 46:47:@1673.4]
  assign _T_55823 = _T_55822[4:0]; // @[Modules.scala 46:47:@1674.4]
  assign _T_55824 = $signed(_T_55823); // @[Modules.scala 46:47:@1675.4]
  assign _T_55826 = $signed(5'sh0) - $signed(io_in_570); // @[Modules.scala 43:37:@1677.4]
  assign _T_55827 = _T_55826[4:0]; // @[Modules.scala 43:37:@1678.4]
  assign _T_55828 = $signed(_T_55827); // @[Modules.scala 43:37:@1679.4]
  assign _T_55829 = $signed(_T_55828) + $signed(io_in_571); // @[Modules.scala 43:47:@1680.4]
  assign _T_55830 = _T_55829[4:0]; // @[Modules.scala 43:47:@1681.4]
  assign _T_55831 = $signed(_T_55830); // @[Modules.scala 43:47:@1682.4]
  assign _T_55833 = $signed(5'sh0) - $signed(io_in_572); // @[Modules.scala 43:37:@1684.4]
  assign _T_55834 = _T_55833[4:0]; // @[Modules.scala 43:37:@1685.4]
  assign _T_55835 = $signed(_T_55834); // @[Modules.scala 43:37:@1686.4]
  assign _T_55836 = $signed(_T_55835) + $signed(io_in_573); // @[Modules.scala 43:47:@1687.4]
  assign _T_55837 = _T_55836[4:0]; // @[Modules.scala 43:47:@1688.4]
  assign _T_55838 = $signed(_T_55837); // @[Modules.scala 43:47:@1689.4]
  assign _T_55840 = $signed(5'sh0) - $signed(io_in_574); // @[Modules.scala 43:37:@1691.4]
  assign _T_55841 = _T_55840[4:0]; // @[Modules.scala 43:37:@1692.4]
  assign _T_55842 = $signed(_T_55841); // @[Modules.scala 43:37:@1693.4]
  assign _T_55843 = $signed(_T_55842) + $signed(io_in_575); // @[Modules.scala 43:47:@1694.4]
  assign _T_55844 = _T_55843[4:0]; // @[Modules.scala 43:47:@1695.4]
  assign _T_55845 = $signed(_T_55844); // @[Modules.scala 43:47:@1696.4]
  assign _T_55846 = $signed(io_in_576) + $signed(io_in_577); // @[Modules.scala 37:46:@1698.4]
  assign _T_55847 = _T_55846[4:0]; // @[Modules.scala 37:46:@1699.4]
  assign _T_55848 = $signed(_T_55847); // @[Modules.scala 37:46:@1700.4]
  assign _T_55849 = $signed(io_in_578) - $signed(io_in_579); // @[Modules.scala 40:46:@1702.4]
  assign _T_55850 = _T_55849[4:0]; // @[Modules.scala 40:46:@1703.4]
  assign _T_55851 = $signed(_T_55850); // @[Modules.scala 40:46:@1704.4]
  assign _T_55852 = $signed(io_in_580) - $signed(io_in_581); // @[Modules.scala 40:46:@1706.4]
  assign _T_55853 = _T_55852[4:0]; // @[Modules.scala 40:46:@1707.4]
  assign _T_55854 = $signed(_T_55853); // @[Modules.scala 40:46:@1708.4]
  assign _T_55856 = $signed(5'sh0) - $signed(io_in_582); // @[Modules.scala 46:37:@1710.4]
  assign _T_55857 = _T_55856[4:0]; // @[Modules.scala 46:37:@1711.4]
  assign _T_55858 = $signed(_T_55857); // @[Modules.scala 46:37:@1712.4]
  assign _T_55859 = $signed(_T_55858) - $signed(io_in_583); // @[Modules.scala 46:47:@1713.4]
  assign _T_55860 = _T_55859[4:0]; // @[Modules.scala 46:47:@1714.4]
  assign _T_55861 = $signed(_T_55860); // @[Modules.scala 46:47:@1715.4]
  assign _T_55862 = $signed(io_in_584) + $signed(io_in_585); // @[Modules.scala 37:46:@1717.4]
  assign _T_55863 = _T_55862[4:0]; // @[Modules.scala 37:46:@1718.4]
  assign _T_55864 = $signed(_T_55863); // @[Modules.scala 37:46:@1719.4]
  assign _T_55866 = $signed(5'sh0) - $signed(io_in_586); // @[Modules.scala 43:37:@1721.4]
  assign _T_55867 = _T_55866[4:0]; // @[Modules.scala 43:37:@1722.4]
  assign _T_55868 = $signed(_T_55867); // @[Modules.scala 43:37:@1723.4]
  assign _T_55869 = $signed(_T_55868) + $signed(io_in_587); // @[Modules.scala 43:47:@1724.4]
  assign _T_55870 = _T_55869[4:0]; // @[Modules.scala 43:47:@1725.4]
  assign _T_55871 = $signed(_T_55870); // @[Modules.scala 43:47:@1726.4]
  assign _T_55873 = $signed(5'sh0) - $signed(io_in_588); // @[Modules.scala 43:37:@1728.4]
  assign _T_55874 = _T_55873[4:0]; // @[Modules.scala 43:37:@1729.4]
  assign _T_55875 = $signed(_T_55874); // @[Modules.scala 43:37:@1730.4]
  assign _T_55876 = $signed(_T_55875) + $signed(io_in_589); // @[Modules.scala 43:47:@1731.4]
  assign _T_55877 = _T_55876[4:0]; // @[Modules.scala 43:47:@1732.4]
  assign _T_55878 = $signed(_T_55877); // @[Modules.scala 43:47:@1733.4]
  assign _T_55880 = $signed(5'sh0) - $signed(io_in_590); // @[Modules.scala 46:37:@1735.4]
  assign _T_55881 = _T_55880[4:0]; // @[Modules.scala 46:37:@1736.4]
  assign _T_55882 = $signed(_T_55881); // @[Modules.scala 46:37:@1737.4]
  assign _T_55883 = $signed(_T_55882) - $signed(io_in_591); // @[Modules.scala 46:47:@1738.4]
  assign _T_55884 = _T_55883[4:0]; // @[Modules.scala 46:47:@1739.4]
  assign _T_55885 = $signed(_T_55884); // @[Modules.scala 46:47:@1740.4]
  assign _T_55887 = $signed(5'sh0) - $signed(io_in_592); // @[Modules.scala 46:37:@1742.4]
  assign _T_55888 = _T_55887[4:0]; // @[Modules.scala 46:37:@1743.4]
  assign _T_55889 = $signed(_T_55888); // @[Modules.scala 46:37:@1744.4]
  assign _T_55890 = $signed(_T_55889) - $signed(io_in_593); // @[Modules.scala 46:47:@1745.4]
  assign _T_55891 = _T_55890[4:0]; // @[Modules.scala 46:47:@1746.4]
  assign _T_55892 = $signed(_T_55891); // @[Modules.scala 46:47:@1747.4]
  assign _T_55894 = $signed(5'sh0) - $signed(io_in_594); // @[Modules.scala 46:37:@1749.4]
  assign _T_55895 = _T_55894[4:0]; // @[Modules.scala 46:37:@1750.4]
  assign _T_55896 = $signed(_T_55895); // @[Modules.scala 46:37:@1751.4]
  assign _T_55897 = $signed(_T_55896) - $signed(io_in_595); // @[Modules.scala 46:47:@1752.4]
  assign _T_55898 = _T_55897[4:0]; // @[Modules.scala 46:47:@1753.4]
  assign _T_55899 = $signed(_T_55898); // @[Modules.scala 46:47:@1754.4]
  assign _T_55901 = $signed(5'sh0) - $signed(io_in_596); // @[Modules.scala 46:37:@1756.4]
  assign _T_55902 = _T_55901[4:0]; // @[Modules.scala 46:37:@1757.4]
  assign _T_55903 = $signed(_T_55902); // @[Modules.scala 46:37:@1758.4]
  assign _T_55904 = $signed(_T_55903) - $signed(io_in_597); // @[Modules.scala 46:47:@1759.4]
  assign _T_55905 = _T_55904[4:0]; // @[Modules.scala 46:47:@1760.4]
  assign _T_55906 = $signed(_T_55905); // @[Modules.scala 46:47:@1761.4]
  assign _T_55908 = $signed(5'sh0) - $signed(io_in_598); // @[Modules.scala 46:37:@1763.4]
  assign _T_55909 = _T_55908[4:0]; // @[Modules.scala 46:37:@1764.4]
  assign _T_55910 = $signed(_T_55909); // @[Modules.scala 46:37:@1765.4]
  assign _T_55911 = $signed(_T_55910) - $signed(io_in_599); // @[Modules.scala 46:47:@1766.4]
  assign _T_55912 = _T_55911[4:0]; // @[Modules.scala 46:47:@1767.4]
  assign _T_55913 = $signed(_T_55912); // @[Modules.scala 46:47:@1768.4]
  assign _T_55914 = $signed(io_in_600) + $signed(io_in_601); // @[Modules.scala 37:46:@1770.4]
  assign _T_55915 = _T_55914[4:0]; // @[Modules.scala 37:46:@1771.4]
  assign _T_55916 = $signed(_T_55915); // @[Modules.scala 37:46:@1772.4]
  assign _T_55917 = $signed(io_in_602) - $signed(io_in_603); // @[Modules.scala 40:46:@1774.4]
  assign _T_55918 = _T_55917[4:0]; // @[Modules.scala 40:46:@1775.4]
  assign _T_55919 = $signed(_T_55918); // @[Modules.scala 40:46:@1776.4]
  assign _T_55920 = $signed(io_in_604) + $signed(io_in_605); // @[Modules.scala 37:46:@1778.4]
  assign _T_55921 = _T_55920[4:0]; // @[Modules.scala 37:46:@1779.4]
  assign _T_55922 = $signed(_T_55921); // @[Modules.scala 37:46:@1780.4]
  assign _T_55923 = $signed(io_in_606) + $signed(io_in_607); // @[Modules.scala 37:46:@1782.4]
  assign _T_55924 = _T_55923[4:0]; // @[Modules.scala 37:46:@1783.4]
  assign _T_55925 = $signed(_T_55924); // @[Modules.scala 37:46:@1784.4]
  assign _T_55927 = $signed(5'sh0) - $signed(io_in_608); // @[Modules.scala 46:37:@1786.4]
  assign _T_55928 = _T_55927[4:0]; // @[Modules.scala 46:37:@1787.4]
  assign _T_55929 = $signed(_T_55928); // @[Modules.scala 46:37:@1788.4]
  assign _T_55930 = $signed(_T_55929) - $signed(io_in_609); // @[Modules.scala 46:47:@1789.4]
  assign _T_55931 = _T_55930[4:0]; // @[Modules.scala 46:47:@1790.4]
  assign _T_55932 = $signed(_T_55931); // @[Modules.scala 46:47:@1791.4]
  assign _T_55934 = $signed(5'sh0) - $signed(io_in_610); // @[Modules.scala 46:37:@1793.4]
  assign _T_55935 = _T_55934[4:0]; // @[Modules.scala 46:37:@1794.4]
  assign _T_55936 = $signed(_T_55935); // @[Modules.scala 46:37:@1795.4]
  assign _T_55937 = $signed(_T_55936) - $signed(io_in_611); // @[Modules.scala 46:47:@1796.4]
  assign _T_55938 = _T_55937[4:0]; // @[Modules.scala 46:47:@1797.4]
  assign _T_55939 = $signed(_T_55938); // @[Modules.scala 46:47:@1798.4]
  assign _T_55940 = $signed(io_in_612) + $signed(io_in_613); // @[Modules.scala 37:46:@1800.4]
  assign _T_55941 = _T_55940[4:0]; // @[Modules.scala 37:46:@1801.4]
  assign _T_55942 = $signed(_T_55941); // @[Modules.scala 37:46:@1802.4]
  assign _T_55944 = $signed(5'sh0) - $signed(io_in_614); // @[Modules.scala 43:37:@1804.4]
  assign _T_55945 = _T_55944[4:0]; // @[Modules.scala 43:37:@1805.4]
  assign _T_55946 = $signed(_T_55945); // @[Modules.scala 43:37:@1806.4]
  assign _T_55947 = $signed(_T_55946) + $signed(io_in_615); // @[Modules.scala 43:47:@1807.4]
  assign _T_55948 = _T_55947[4:0]; // @[Modules.scala 43:47:@1808.4]
  assign _T_55949 = $signed(_T_55948); // @[Modules.scala 43:47:@1809.4]
  assign _T_55951 = $signed(5'sh0) - $signed(io_in_616); // @[Modules.scala 43:37:@1811.4]
  assign _T_55952 = _T_55951[4:0]; // @[Modules.scala 43:37:@1812.4]
  assign _T_55953 = $signed(_T_55952); // @[Modules.scala 43:37:@1813.4]
  assign _T_55954 = $signed(_T_55953) + $signed(io_in_617); // @[Modules.scala 43:47:@1814.4]
  assign _T_55955 = _T_55954[4:0]; // @[Modules.scala 43:47:@1815.4]
  assign _T_55956 = $signed(_T_55955); // @[Modules.scala 43:47:@1816.4]
  assign _T_55957 = $signed(io_in_618) + $signed(io_in_619); // @[Modules.scala 37:46:@1818.4]
  assign _T_55958 = _T_55957[4:0]; // @[Modules.scala 37:46:@1819.4]
  assign _T_55959 = $signed(_T_55958); // @[Modules.scala 37:46:@1820.4]
  assign _T_55961 = $signed(5'sh0) - $signed(io_in_620); // @[Modules.scala 46:37:@1822.4]
  assign _T_55962 = _T_55961[4:0]; // @[Modules.scala 46:37:@1823.4]
  assign _T_55963 = $signed(_T_55962); // @[Modules.scala 46:37:@1824.4]
  assign _T_55964 = $signed(_T_55963) - $signed(io_in_621); // @[Modules.scala 46:47:@1825.4]
  assign _T_55965 = _T_55964[4:0]; // @[Modules.scala 46:47:@1826.4]
  assign _T_55966 = $signed(_T_55965); // @[Modules.scala 46:47:@1827.4]
  assign _T_55968 = $signed(5'sh0) - $signed(io_in_622); // @[Modules.scala 46:37:@1829.4]
  assign _T_55969 = _T_55968[4:0]; // @[Modules.scala 46:37:@1830.4]
  assign _T_55970 = $signed(_T_55969); // @[Modules.scala 46:37:@1831.4]
  assign _T_55971 = $signed(_T_55970) - $signed(io_in_623); // @[Modules.scala 46:47:@1832.4]
  assign _T_55972 = _T_55971[4:0]; // @[Modules.scala 46:47:@1833.4]
  assign _T_55973 = $signed(_T_55972); // @[Modules.scala 46:47:@1834.4]
  assign _T_55975 = $signed(5'sh0) - $signed(io_in_624); // @[Modules.scala 46:37:@1836.4]
  assign _T_55976 = _T_55975[4:0]; // @[Modules.scala 46:37:@1837.4]
  assign _T_55977 = $signed(_T_55976); // @[Modules.scala 46:37:@1838.4]
  assign _T_55978 = $signed(_T_55977) - $signed(io_in_625); // @[Modules.scala 46:47:@1839.4]
  assign _T_55979 = _T_55978[4:0]; // @[Modules.scala 46:47:@1840.4]
  assign _T_55980 = $signed(_T_55979); // @[Modules.scala 46:47:@1841.4]
  assign _T_55982 = $signed(5'sh0) - $signed(io_in_626); // @[Modules.scala 46:37:@1843.4]
  assign _T_55983 = _T_55982[4:0]; // @[Modules.scala 46:37:@1844.4]
  assign _T_55984 = $signed(_T_55983); // @[Modules.scala 46:37:@1845.4]
  assign _T_55985 = $signed(_T_55984) - $signed(io_in_627); // @[Modules.scala 46:47:@1846.4]
  assign _T_55986 = _T_55985[4:0]; // @[Modules.scala 46:47:@1847.4]
  assign _T_55987 = $signed(_T_55986); // @[Modules.scala 46:47:@1848.4]
  assign _T_55989 = $signed(5'sh0) - $signed(io_in_628); // @[Modules.scala 46:37:@1850.4]
  assign _T_55990 = _T_55989[4:0]; // @[Modules.scala 46:37:@1851.4]
  assign _T_55991 = $signed(_T_55990); // @[Modules.scala 46:37:@1852.4]
  assign _T_55992 = $signed(_T_55991) - $signed(io_in_629); // @[Modules.scala 46:47:@1853.4]
  assign _T_55993 = _T_55992[4:0]; // @[Modules.scala 46:47:@1854.4]
  assign _T_55994 = $signed(_T_55993); // @[Modules.scala 46:47:@1855.4]
  assign _T_55996 = $signed(5'sh0) - $signed(io_in_630); // @[Modules.scala 46:37:@1857.4]
  assign _T_55997 = _T_55996[4:0]; // @[Modules.scala 46:37:@1858.4]
  assign _T_55998 = $signed(_T_55997); // @[Modules.scala 46:37:@1859.4]
  assign _T_55999 = $signed(_T_55998) - $signed(io_in_631); // @[Modules.scala 46:47:@1860.4]
  assign _T_56000 = _T_55999[4:0]; // @[Modules.scala 46:47:@1861.4]
  assign _T_56001 = $signed(_T_56000); // @[Modules.scala 46:47:@1862.4]
  assign _T_56003 = $signed(5'sh0) - $signed(io_in_632); // @[Modules.scala 46:37:@1864.4]
  assign _T_56004 = _T_56003[4:0]; // @[Modules.scala 46:37:@1865.4]
  assign _T_56005 = $signed(_T_56004); // @[Modules.scala 46:37:@1866.4]
  assign _T_56006 = $signed(_T_56005) - $signed(io_in_633); // @[Modules.scala 46:47:@1867.4]
  assign _T_56007 = _T_56006[4:0]; // @[Modules.scala 46:47:@1868.4]
  assign _T_56008 = $signed(_T_56007); // @[Modules.scala 46:47:@1869.4]
  assign _T_56010 = $signed(5'sh0) - $signed(io_in_634); // @[Modules.scala 46:37:@1871.4]
  assign _T_56011 = _T_56010[4:0]; // @[Modules.scala 46:37:@1872.4]
  assign _T_56012 = $signed(_T_56011); // @[Modules.scala 46:37:@1873.4]
  assign _T_56013 = $signed(_T_56012) - $signed(io_in_635); // @[Modules.scala 46:47:@1874.4]
  assign _T_56014 = _T_56013[4:0]; // @[Modules.scala 46:47:@1875.4]
  assign _T_56015 = $signed(_T_56014); // @[Modules.scala 46:47:@1876.4]
  assign _T_56017 = $signed(5'sh0) - $signed(io_in_636); // @[Modules.scala 46:37:@1878.4]
  assign _T_56018 = _T_56017[4:0]; // @[Modules.scala 46:37:@1879.4]
  assign _T_56019 = $signed(_T_56018); // @[Modules.scala 46:37:@1880.4]
  assign _T_56020 = $signed(_T_56019) - $signed(io_in_637); // @[Modules.scala 46:47:@1881.4]
  assign _T_56021 = _T_56020[4:0]; // @[Modules.scala 46:47:@1882.4]
  assign _T_56022 = $signed(_T_56021); // @[Modules.scala 46:47:@1883.4]
  assign _T_56024 = $signed(5'sh0) - $signed(io_in_638); // @[Modules.scala 43:37:@1885.4]
  assign _T_56025 = _T_56024[4:0]; // @[Modules.scala 43:37:@1886.4]
  assign _T_56026 = $signed(_T_56025); // @[Modules.scala 43:37:@1887.4]
  assign _T_56027 = $signed(_T_56026) + $signed(io_in_639); // @[Modules.scala 43:47:@1888.4]
  assign _T_56028 = _T_56027[4:0]; // @[Modules.scala 43:47:@1889.4]
  assign _T_56029 = $signed(_T_56028); // @[Modules.scala 43:47:@1890.4]
  assign _T_56030 = $signed(io_in_640) + $signed(io_in_641); // @[Modules.scala 37:46:@1892.4]
  assign _T_56031 = _T_56030[4:0]; // @[Modules.scala 37:46:@1893.4]
  assign _T_56032 = $signed(_T_56031); // @[Modules.scala 37:46:@1894.4]
  assign _T_56034 = $signed(5'sh0) - $signed(io_in_642); // @[Modules.scala 43:37:@1896.4]
  assign _T_56035 = _T_56034[4:0]; // @[Modules.scala 43:37:@1897.4]
  assign _T_56036 = $signed(_T_56035); // @[Modules.scala 43:37:@1898.4]
  assign _T_56037 = $signed(_T_56036) + $signed(io_in_643); // @[Modules.scala 43:47:@1899.4]
  assign _T_56038 = _T_56037[4:0]; // @[Modules.scala 43:47:@1900.4]
  assign _T_56039 = $signed(_T_56038); // @[Modules.scala 43:47:@1901.4]
  assign _T_56041 = $signed(5'sh0) - $signed(io_in_644); // @[Modules.scala 43:37:@1903.4]
  assign _T_56042 = _T_56041[4:0]; // @[Modules.scala 43:37:@1904.4]
  assign _T_56043 = $signed(_T_56042); // @[Modules.scala 43:37:@1905.4]
  assign _T_56044 = $signed(_T_56043) + $signed(io_in_645); // @[Modules.scala 43:47:@1906.4]
  assign _T_56045 = _T_56044[4:0]; // @[Modules.scala 43:47:@1907.4]
  assign _T_56046 = $signed(_T_56045); // @[Modules.scala 43:47:@1908.4]
  assign _T_56047 = $signed(io_in_646) + $signed(io_in_647); // @[Modules.scala 37:46:@1910.4]
  assign _T_56048 = _T_56047[4:0]; // @[Modules.scala 37:46:@1911.4]
  assign _T_56049 = $signed(_T_56048); // @[Modules.scala 37:46:@1912.4]
  assign _T_56051 = $signed(5'sh0) - $signed(io_in_648); // @[Modules.scala 46:37:@1914.4]
  assign _T_56052 = _T_56051[4:0]; // @[Modules.scala 46:37:@1915.4]
  assign _T_56053 = $signed(_T_56052); // @[Modules.scala 46:37:@1916.4]
  assign _T_56054 = $signed(_T_56053) - $signed(io_in_649); // @[Modules.scala 46:47:@1917.4]
  assign _T_56055 = _T_56054[4:0]; // @[Modules.scala 46:47:@1918.4]
  assign _T_56056 = $signed(_T_56055); // @[Modules.scala 46:47:@1919.4]
  assign _T_56058 = $signed(5'sh0) - $signed(io_in_650); // @[Modules.scala 46:37:@1921.4]
  assign _T_56059 = _T_56058[4:0]; // @[Modules.scala 46:37:@1922.4]
  assign _T_56060 = $signed(_T_56059); // @[Modules.scala 46:37:@1923.4]
  assign _T_56061 = $signed(_T_56060) - $signed(io_in_651); // @[Modules.scala 46:47:@1924.4]
  assign _T_56062 = _T_56061[4:0]; // @[Modules.scala 46:47:@1925.4]
  assign _T_56063 = $signed(_T_56062); // @[Modules.scala 46:47:@1926.4]
  assign _T_56065 = $signed(5'sh0) - $signed(io_in_652); // @[Modules.scala 46:37:@1928.4]
  assign _T_56066 = _T_56065[4:0]; // @[Modules.scala 46:37:@1929.4]
  assign _T_56067 = $signed(_T_56066); // @[Modules.scala 46:37:@1930.4]
  assign _T_56068 = $signed(_T_56067) - $signed(io_in_653); // @[Modules.scala 46:47:@1931.4]
  assign _T_56069 = _T_56068[4:0]; // @[Modules.scala 46:47:@1932.4]
  assign _T_56070 = $signed(_T_56069); // @[Modules.scala 46:47:@1933.4]
  assign _T_56072 = $signed(5'sh0) - $signed(io_in_654); // @[Modules.scala 46:37:@1935.4]
  assign _T_56073 = _T_56072[4:0]; // @[Modules.scala 46:37:@1936.4]
  assign _T_56074 = $signed(_T_56073); // @[Modules.scala 46:37:@1937.4]
  assign _T_56075 = $signed(_T_56074) - $signed(io_in_655); // @[Modules.scala 46:47:@1938.4]
  assign _T_56076 = _T_56075[4:0]; // @[Modules.scala 46:47:@1939.4]
  assign _T_56077 = $signed(_T_56076); // @[Modules.scala 46:47:@1940.4]
  assign _T_56079 = $signed(5'sh0) - $signed(io_in_656); // @[Modules.scala 46:37:@1942.4]
  assign _T_56080 = _T_56079[4:0]; // @[Modules.scala 46:37:@1943.4]
  assign _T_56081 = $signed(_T_56080); // @[Modules.scala 46:37:@1944.4]
  assign _T_56082 = $signed(_T_56081) - $signed(io_in_657); // @[Modules.scala 46:47:@1945.4]
  assign _T_56083 = _T_56082[4:0]; // @[Modules.scala 46:47:@1946.4]
  assign _T_56084 = $signed(_T_56083); // @[Modules.scala 46:47:@1947.4]
  assign _T_56086 = $signed(5'sh0) - $signed(io_in_658); // @[Modules.scala 46:37:@1949.4]
  assign _T_56087 = _T_56086[4:0]; // @[Modules.scala 46:37:@1950.4]
  assign _T_56088 = $signed(_T_56087); // @[Modules.scala 46:37:@1951.4]
  assign _T_56089 = $signed(_T_56088) - $signed(io_in_659); // @[Modules.scala 46:47:@1952.4]
  assign _T_56090 = _T_56089[4:0]; // @[Modules.scala 46:47:@1953.4]
  assign _T_56091 = $signed(_T_56090); // @[Modules.scala 46:47:@1954.4]
  assign _T_56093 = $signed(5'sh0) - $signed(io_in_660); // @[Modules.scala 46:37:@1956.4]
  assign _T_56094 = _T_56093[4:0]; // @[Modules.scala 46:37:@1957.4]
  assign _T_56095 = $signed(_T_56094); // @[Modules.scala 46:37:@1958.4]
  assign _T_56096 = $signed(_T_56095) - $signed(io_in_661); // @[Modules.scala 46:47:@1959.4]
  assign _T_56097 = _T_56096[4:0]; // @[Modules.scala 46:47:@1960.4]
  assign _T_56098 = $signed(_T_56097); // @[Modules.scala 46:47:@1961.4]
  assign _T_56100 = $signed(5'sh0) - $signed(io_in_662); // @[Modules.scala 43:37:@1963.4]
  assign _T_56101 = _T_56100[4:0]; // @[Modules.scala 43:37:@1964.4]
  assign _T_56102 = $signed(_T_56101); // @[Modules.scala 43:37:@1965.4]
  assign _T_56103 = $signed(_T_56102) + $signed(io_in_663); // @[Modules.scala 43:47:@1966.4]
  assign _T_56104 = _T_56103[4:0]; // @[Modules.scala 43:47:@1967.4]
  assign _T_56105 = $signed(_T_56104); // @[Modules.scala 43:47:@1968.4]
  assign _T_56106 = $signed(io_in_664) + $signed(io_in_665); // @[Modules.scala 37:46:@1970.4]
  assign _T_56107 = _T_56106[4:0]; // @[Modules.scala 37:46:@1971.4]
  assign _T_56108 = $signed(_T_56107); // @[Modules.scala 37:46:@1972.4]
  assign _T_56109 = $signed(io_in_666) + $signed(io_in_667); // @[Modules.scala 37:46:@1974.4]
  assign _T_56110 = _T_56109[4:0]; // @[Modules.scala 37:46:@1975.4]
  assign _T_56111 = $signed(_T_56110); // @[Modules.scala 37:46:@1976.4]
  assign _T_56112 = $signed(io_in_668) + $signed(io_in_669); // @[Modules.scala 37:46:@1978.4]
  assign _T_56113 = _T_56112[4:0]; // @[Modules.scala 37:46:@1979.4]
  assign _T_56114 = $signed(_T_56113); // @[Modules.scala 37:46:@1980.4]
  assign _T_56116 = $signed(5'sh0) - $signed(io_in_670); // @[Modules.scala 46:37:@1982.4]
  assign _T_56117 = _T_56116[4:0]; // @[Modules.scala 46:37:@1983.4]
  assign _T_56118 = $signed(_T_56117); // @[Modules.scala 46:37:@1984.4]
  assign _T_56119 = $signed(_T_56118) - $signed(io_in_671); // @[Modules.scala 46:47:@1985.4]
  assign _T_56120 = _T_56119[4:0]; // @[Modules.scala 46:47:@1986.4]
  assign _T_56121 = $signed(_T_56120); // @[Modules.scala 46:47:@1987.4]
  assign _T_56123 = $signed(5'sh0) - $signed(io_in_672); // @[Modules.scala 43:37:@1989.4]
  assign _T_56124 = _T_56123[4:0]; // @[Modules.scala 43:37:@1990.4]
  assign _T_56125 = $signed(_T_56124); // @[Modules.scala 43:37:@1991.4]
  assign _T_56126 = $signed(_T_56125) + $signed(io_in_673); // @[Modules.scala 43:47:@1992.4]
  assign _T_56127 = _T_56126[4:0]; // @[Modules.scala 43:47:@1993.4]
  assign _T_56128 = $signed(_T_56127); // @[Modules.scala 43:47:@1994.4]
  assign _T_56129 = $signed(io_in_674) - $signed(io_in_675); // @[Modules.scala 40:46:@1996.4]
  assign _T_56130 = _T_56129[4:0]; // @[Modules.scala 40:46:@1997.4]
  assign _T_56131 = $signed(_T_56130); // @[Modules.scala 40:46:@1998.4]
  assign _T_56132 = $signed(io_in_676) + $signed(io_in_677); // @[Modules.scala 37:46:@2000.4]
  assign _T_56133 = _T_56132[4:0]; // @[Modules.scala 37:46:@2001.4]
  assign _T_56134 = $signed(_T_56133); // @[Modules.scala 37:46:@2002.4]
  assign _T_56135 = $signed(io_in_678) + $signed(io_in_679); // @[Modules.scala 37:46:@2004.4]
  assign _T_56136 = _T_56135[4:0]; // @[Modules.scala 37:46:@2005.4]
  assign _T_56137 = $signed(_T_56136); // @[Modules.scala 37:46:@2006.4]
  assign _T_56138 = $signed(io_in_680) + $signed(io_in_681); // @[Modules.scala 37:46:@2008.4]
  assign _T_56139 = _T_56138[4:0]; // @[Modules.scala 37:46:@2009.4]
  assign _T_56140 = $signed(_T_56139); // @[Modules.scala 37:46:@2010.4]
  assign _T_56141 = $signed(io_in_682) - $signed(io_in_683); // @[Modules.scala 40:46:@2012.4]
  assign _T_56142 = _T_56141[4:0]; // @[Modules.scala 40:46:@2013.4]
  assign _T_56143 = $signed(_T_56142); // @[Modules.scala 40:46:@2014.4]
  assign _T_56145 = $signed(5'sh0) - $signed(io_in_684); // @[Modules.scala 46:37:@2016.4]
  assign _T_56146 = _T_56145[4:0]; // @[Modules.scala 46:37:@2017.4]
  assign _T_56147 = $signed(_T_56146); // @[Modules.scala 46:37:@2018.4]
  assign _T_56148 = $signed(_T_56147) - $signed(io_in_685); // @[Modules.scala 46:47:@2019.4]
  assign _T_56149 = _T_56148[4:0]; // @[Modules.scala 46:47:@2020.4]
  assign _T_56150 = $signed(_T_56149); // @[Modules.scala 46:47:@2021.4]
  assign _T_56152 = $signed(5'sh0) - $signed(io_in_686); // @[Modules.scala 46:37:@2023.4]
  assign _T_56153 = _T_56152[4:0]; // @[Modules.scala 46:37:@2024.4]
  assign _T_56154 = $signed(_T_56153); // @[Modules.scala 46:37:@2025.4]
  assign _T_56155 = $signed(_T_56154) - $signed(io_in_687); // @[Modules.scala 46:47:@2026.4]
  assign _T_56156 = _T_56155[4:0]; // @[Modules.scala 46:47:@2027.4]
  assign _T_56157 = $signed(_T_56156); // @[Modules.scala 46:47:@2028.4]
  assign _T_56158 = $signed(io_in_688) + $signed(io_in_689); // @[Modules.scala 37:46:@2030.4]
  assign _T_56159 = _T_56158[4:0]; // @[Modules.scala 37:46:@2031.4]
  assign _T_56160 = $signed(_T_56159); // @[Modules.scala 37:46:@2032.4]
  assign _T_56161 = $signed(io_in_690) + $signed(io_in_691); // @[Modules.scala 37:46:@2034.4]
  assign _T_56162 = _T_56161[4:0]; // @[Modules.scala 37:46:@2035.4]
  assign _T_56163 = $signed(_T_56162); // @[Modules.scala 37:46:@2036.4]
  assign _T_56164 = $signed(io_in_692) + $signed(io_in_693); // @[Modules.scala 37:46:@2038.4]
  assign _T_56165 = _T_56164[4:0]; // @[Modules.scala 37:46:@2039.4]
  assign _T_56166 = $signed(_T_56165); // @[Modules.scala 37:46:@2040.4]
  assign _T_56167 = $signed(io_in_694) + $signed(io_in_695); // @[Modules.scala 37:46:@2042.4]
  assign _T_56168 = _T_56167[4:0]; // @[Modules.scala 37:46:@2043.4]
  assign _T_56169 = $signed(_T_56168); // @[Modules.scala 37:46:@2044.4]
  assign _T_56170 = $signed(io_in_696) + $signed(io_in_697); // @[Modules.scala 37:46:@2046.4]
  assign _T_56171 = _T_56170[4:0]; // @[Modules.scala 37:46:@2047.4]
  assign _T_56172 = $signed(_T_56171); // @[Modules.scala 37:46:@2048.4]
  assign _T_56174 = $signed(5'sh0) - $signed(io_in_698); // @[Modules.scala 43:37:@2050.4]
  assign _T_56175 = _T_56174[4:0]; // @[Modules.scala 43:37:@2051.4]
  assign _T_56176 = $signed(_T_56175); // @[Modules.scala 43:37:@2052.4]
  assign _T_56177 = $signed(_T_56176) + $signed(io_in_699); // @[Modules.scala 43:47:@2053.4]
  assign _T_56178 = _T_56177[4:0]; // @[Modules.scala 43:47:@2054.4]
  assign _T_56179 = $signed(_T_56178); // @[Modules.scala 43:47:@2055.4]
  assign _T_56181 = $signed(5'sh0) - $signed(io_in_700); // @[Modules.scala 43:37:@2057.4]
  assign _T_56182 = _T_56181[4:0]; // @[Modules.scala 43:37:@2058.4]
  assign _T_56183 = $signed(_T_56182); // @[Modules.scala 43:37:@2059.4]
  assign _T_56184 = $signed(_T_56183) + $signed(io_in_701); // @[Modules.scala 43:47:@2060.4]
  assign _T_56185 = _T_56184[4:0]; // @[Modules.scala 43:47:@2061.4]
  assign _T_56186 = $signed(_T_56185); // @[Modules.scala 43:47:@2062.4]
  assign _T_56187 = $signed(io_in_702) - $signed(io_in_703); // @[Modules.scala 40:46:@2064.4]
  assign _T_56188 = _T_56187[4:0]; // @[Modules.scala 40:46:@2065.4]
  assign _T_56189 = $signed(_T_56188); // @[Modules.scala 40:46:@2066.4]
  assign _T_56190 = $signed(io_in_704) + $signed(io_in_705); // @[Modules.scala 37:46:@2068.4]
  assign _T_56191 = _T_56190[4:0]; // @[Modules.scala 37:46:@2069.4]
  assign _T_56192 = $signed(_T_56191); // @[Modules.scala 37:46:@2070.4]
  assign _T_56193 = $signed(io_in_706) + $signed(io_in_707); // @[Modules.scala 37:46:@2072.4]
  assign _T_56194 = _T_56193[4:0]; // @[Modules.scala 37:46:@2073.4]
  assign _T_56195 = $signed(_T_56194); // @[Modules.scala 37:46:@2074.4]
  assign _T_56196 = $signed(io_in_708) + $signed(io_in_709); // @[Modules.scala 37:46:@2076.4]
  assign _T_56197 = _T_56196[4:0]; // @[Modules.scala 37:46:@2077.4]
  assign _T_56198 = $signed(_T_56197); // @[Modules.scala 37:46:@2078.4]
  assign _T_56199 = $signed(io_in_710) - $signed(io_in_711); // @[Modules.scala 40:46:@2080.4]
  assign _T_56200 = _T_56199[4:0]; // @[Modules.scala 40:46:@2081.4]
  assign _T_56201 = $signed(_T_56200); // @[Modules.scala 40:46:@2082.4]
  assign _T_56202 = $signed(io_in_712) + $signed(io_in_713); // @[Modules.scala 37:46:@2084.4]
  assign _T_56203 = _T_56202[4:0]; // @[Modules.scala 37:46:@2085.4]
  assign _T_56204 = $signed(_T_56203); // @[Modules.scala 37:46:@2086.4]
  assign _T_56205 = $signed(io_in_714) + $signed(io_in_715); // @[Modules.scala 37:46:@2088.4]
  assign _T_56206 = _T_56205[4:0]; // @[Modules.scala 37:46:@2089.4]
  assign _T_56207 = $signed(_T_56206); // @[Modules.scala 37:46:@2090.4]
  assign _T_56208 = $signed(io_in_716) + $signed(io_in_717); // @[Modules.scala 37:46:@2092.4]
  assign _T_56209 = _T_56208[4:0]; // @[Modules.scala 37:46:@2093.4]
  assign _T_56210 = $signed(_T_56209); // @[Modules.scala 37:46:@2094.4]
  assign _T_56211 = $signed(io_in_718) + $signed(io_in_719); // @[Modules.scala 37:46:@2096.4]
  assign _T_56212 = _T_56211[4:0]; // @[Modules.scala 37:46:@2097.4]
  assign _T_56213 = $signed(_T_56212); // @[Modules.scala 37:46:@2098.4]
  assign _T_56214 = $signed(io_in_720) + $signed(io_in_721); // @[Modules.scala 37:46:@2100.4]
  assign _T_56215 = _T_56214[4:0]; // @[Modules.scala 37:46:@2101.4]
  assign _T_56216 = $signed(_T_56215); // @[Modules.scala 37:46:@2102.4]
  assign _T_56217 = $signed(io_in_722) + $signed(io_in_723); // @[Modules.scala 37:46:@2104.4]
  assign _T_56218 = _T_56217[4:0]; // @[Modules.scala 37:46:@2105.4]
  assign _T_56219 = $signed(_T_56218); // @[Modules.scala 37:46:@2106.4]
  assign _T_56220 = $signed(io_in_724) - $signed(io_in_725); // @[Modules.scala 40:46:@2108.4]
  assign _T_56221 = _T_56220[4:0]; // @[Modules.scala 40:46:@2109.4]
  assign _T_56222 = $signed(_T_56221); // @[Modules.scala 40:46:@2110.4]
  assign _T_56224 = $signed(5'sh0) - $signed(io_in_726); // @[Modules.scala 46:37:@2112.4]
  assign _T_56225 = _T_56224[4:0]; // @[Modules.scala 46:37:@2113.4]
  assign _T_56226 = $signed(_T_56225); // @[Modules.scala 46:37:@2114.4]
  assign _T_56227 = $signed(_T_56226) - $signed(io_in_727); // @[Modules.scala 46:47:@2115.4]
  assign _T_56228 = _T_56227[4:0]; // @[Modules.scala 46:47:@2116.4]
  assign _T_56229 = $signed(_T_56228); // @[Modules.scala 46:47:@2117.4]
  assign _T_56230 = $signed(io_in_728) - $signed(io_in_729); // @[Modules.scala 40:46:@2119.4]
  assign _T_56231 = _T_56230[4:0]; // @[Modules.scala 40:46:@2120.4]
  assign _T_56232 = $signed(_T_56231); // @[Modules.scala 40:46:@2121.4]
  assign _T_56234 = $signed(5'sh0) - $signed(io_in_730); // @[Modules.scala 43:37:@2123.4]
  assign _T_56235 = _T_56234[4:0]; // @[Modules.scala 43:37:@2124.4]
  assign _T_56236 = $signed(_T_56235); // @[Modules.scala 43:37:@2125.4]
  assign _T_56237 = $signed(_T_56236) + $signed(io_in_731); // @[Modules.scala 43:47:@2126.4]
  assign _T_56238 = _T_56237[4:0]; // @[Modules.scala 43:47:@2127.4]
  assign _T_56239 = $signed(_T_56238); // @[Modules.scala 43:47:@2128.4]
  assign _T_56240 = $signed(io_in_732) + $signed(io_in_733); // @[Modules.scala 37:46:@2130.4]
  assign _T_56241 = _T_56240[4:0]; // @[Modules.scala 37:46:@2131.4]
  assign _T_56242 = $signed(_T_56241); // @[Modules.scala 37:46:@2132.4]
  assign _T_56243 = $signed(io_in_734) + $signed(io_in_735); // @[Modules.scala 37:46:@2134.4]
  assign _T_56244 = _T_56243[4:0]; // @[Modules.scala 37:46:@2135.4]
  assign _T_56245 = $signed(_T_56244); // @[Modules.scala 37:46:@2136.4]
  assign _T_56247 = $signed(5'sh0) - $signed(io_in_736); // @[Modules.scala 46:37:@2138.4]
  assign _T_56248 = _T_56247[4:0]; // @[Modules.scala 46:37:@2139.4]
  assign _T_56249 = $signed(_T_56248); // @[Modules.scala 46:37:@2140.4]
  assign _T_56250 = $signed(_T_56249) - $signed(io_in_737); // @[Modules.scala 46:47:@2141.4]
  assign _T_56251 = _T_56250[4:0]; // @[Modules.scala 46:47:@2142.4]
  assign _T_56252 = $signed(_T_56251); // @[Modules.scala 46:47:@2143.4]
  assign _T_56254 = $signed(5'sh0) - $signed(io_in_738); // @[Modules.scala 46:37:@2145.4]
  assign _T_56255 = _T_56254[4:0]; // @[Modules.scala 46:37:@2146.4]
  assign _T_56256 = $signed(_T_56255); // @[Modules.scala 46:37:@2147.4]
  assign _T_56257 = $signed(_T_56256) - $signed(io_in_739); // @[Modules.scala 46:47:@2148.4]
  assign _T_56258 = _T_56257[4:0]; // @[Modules.scala 46:47:@2149.4]
  assign _T_56259 = $signed(_T_56258); // @[Modules.scala 46:47:@2150.4]
  assign _T_56260 = $signed(io_in_740) - $signed(io_in_741); // @[Modules.scala 40:46:@2152.4]
  assign _T_56261 = _T_56260[4:0]; // @[Modules.scala 40:46:@2153.4]
  assign _T_56262 = $signed(_T_56261); // @[Modules.scala 40:46:@2154.4]
  assign _T_56263 = $signed(io_in_742) - $signed(io_in_743); // @[Modules.scala 40:46:@2156.4]
  assign _T_56264 = _T_56263[4:0]; // @[Modules.scala 40:46:@2157.4]
  assign _T_56265 = $signed(_T_56264); // @[Modules.scala 40:46:@2158.4]
  assign _T_56267 = $signed(5'sh0) - $signed(io_in_744); // @[Modules.scala 46:37:@2160.4]
  assign _T_56268 = _T_56267[4:0]; // @[Modules.scala 46:37:@2161.4]
  assign _T_56269 = $signed(_T_56268); // @[Modules.scala 46:37:@2162.4]
  assign _T_56270 = $signed(_T_56269) - $signed(io_in_745); // @[Modules.scala 46:47:@2163.4]
  assign _T_56271 = _T_56270[4:0]; // @[Modules.scala 46:47:@2164.4]
  assign _T_56272 = $signed(_T_56271); // @[Modules.scala 46:47:@2165.4]
  assign _T_56274 = $signed(5'sh0) - $signed(io_in_746); // @[Modules.scala 46:37:@2167.4]
  assign _T_56275 = _T_56274[4:0]; // @[Modules.scala 46:37:@2168.4]
  assign _T_56276 = $signed(_T_56275); // @[Modules.scala 46:37:@2169.4]
  assign _T_56277 = $signed(_T_56276) - $signed(io_in_747); // @[Modules.scala 46:47:@2170.4]
  assign _T_56278 = _T_56277[4:0]; // @[Modules.scala 46:47:@2171.4]
  assign _T_56279 = $signed(_T_56278); // @[Modules.scala 46:47:@2172.4]
  assign _T_56280 = $signed(io_in_748) + $signed(io_in_749); // @[Modules.scala 37:46:@2174.4]
  assign _T_56281 = _T_56280[4:0]; // @[Modules.scala 37:46:@2175.4]
  assign _T_56282 = $signed(_T_56281); // @[Modules.scala 37:46:@2176.4]
  assign _T_56283 = $signed(io_in_750) - $signed(io_in_751); // @[Modules.scala 40:46:@2178.4]
  assign _T_56284 = _T_56283[4:0]; // @[Modules.scala 40:46:@2179.4]
  assign _T_56285 = $signed(_T_56284); // @[Modules.scala 40:46:@2180.4]
  assign _T_56286 = $signed(io_in_752) + $signed(io_in_753); // @[Modules.scala 37:46:@2182.4]
  assign _T_56287 = _T_56286[4:0]; // @[Modules.scala 37:46:@2183.4]
  assign _T_56288 = $signed(_T_56287); // @[Modules.scala 37:46:@2184.4]
  assign _T_56289 = $signed(io_in_754) + $signed(io_in_755); // @[Modules.scala 37:46:@2186.4]
  assign _T_56290 = _T_56289[4:0]; // @[Modules.scala 37:46:@2187.4]
  assign _T_56291 = $signed(_T_56290); // @[Modules.scala 37:46:@2188.4]
  assign _T_56293 = $signed(5'sh0) - $signed(io_in_756); // @[Modules.scala 43:37:@2190.4]
  assign _T_56294 = _T_56293[4:0]; // @[Modules.scala 43:37:@2191.4]
  assign _T_56295 = $signed(_T_56294); // @[Modules.scala 43:37:@2192.4]
  assign _T_56296 = $signed(_T_56295) + $signed(io_in_757); // @[Modules.scala 43:47:@2193.4]
  assign _T_56297 = _T_56296[4:0]; // @[Modules.scala 43:47:@2194.4]
  assign _T_56298 = $signed(_T_56297); // @[Modules.scala 43:47:@2195.4]
  assign _T_56300 = $signed(5'sh0) - $signed(io_in_758); // @[Modules.scala 46:37:@2197.4]
  assign _T_56301 = _T_56300[4:0]; // @[Modules.scala 46:37:@2198.4]
  assign _T_56302 = $signed(_T_56301); // @[Modules.scala 46:37:@2199.4]
  assign _T_56303 = $signed(_T_56302) - $signed(io_in_759); // @[Modules.scala 46:47:@2200.4]
  assign _T_56304 = _T_56303[4:0]; // @[Modules.scala 46:47:@2201.4]
  assign _T_56305 = $signed(_T_56304); // @[Modules.scala 46:47:@2202.4]
  assign _T_56306 = $signed(io_in_760) - $signed(io_in_761); // @[Modules.scala 40:46:@2204.4]
  assign _T_56307 = _T_56306[4:0]; // @[Modules.scala 40:46:@2205.4]
  assign _T_56308 = $signed(_T_56307); // @[Modules.scala 40:46:@2206.4]
  assign _T_56310 = $signed(5'sh0) - $signed(io_in_762); // @[Modules.scala 46:37:@2208.4]
  assign _T_56311 = _T_56310[4:0]; // @[Modules.scala 46:37:@2209.4]
  assign _T_56312 = $signed(_T_56311); // @[Modules.scala 46:37:@2210.4]
  assign _T_56313 = $signed(_T_56312) - $signed(io_in_763); // @[Modules.scala 46:47:@2211.4]
  assign _T_56314 = _T_56313[4:0]; // @[Modules.scala 46:47:@2212.4]
  assign _T_56315 = $signed(_T_56314); // @[Modules.scala 46:47:@2213.4]
  assign _T_56317 = $signed(5'sh0) - $signed(io_in_764); // @[Modules.scala 46:37:@2215.4]
  assign _T_56318 = _T_56317[4:0]; // @[Modules.scala 46:37:@2216.4]
  assign _T_56319 = $signed(_T_56318); // @[Modules.scala 46:37:@2217.4]
  assign _T_56320 = $signed(_T_56319) - $signed(io_in_765); // @[Modules.scala 46:47:@2218.4]
  assign _T_56321 = _T_56320[4:0]; // @[Modules.scala 46:47:@2219.4]
  assign _T_56322 = $signed(_T_56321); // @[Modules.scala 46:47:@2220.4]
  assign _T_56324 = $signed(5'sh0) - $signed(io_in_766); // @[Modules.scala 46:37:@2222.4]
  assign _T_56325 = _T_56324[4:0]; // @[Modules.scala 46:37:@2223.4]
  assign _T_56326 = $signed(_T_56325); // @[Modules.scala 46:37:@2224.4]
  assign _T_56327 = $signed(_T_56326) - $signed(io_in_767); // @[Modules.scala 46:47:@2225.4]
  assign _T_56328 = _T_56327[4:0]; // @[Modules.scala 46:47:@2226.4]
  assign _T_56329 = $signed(_T_56328); // @[Modules.scala 46:47:@2227.4]
  assign _T_56330 = $signed(io_in_768) - $signed(io_in_769); // @[Modules.scala 40:46:@2229.4]
  assign _T_56331 = _T_56330[4:0]; // @[Modules.scala 40:46:@2230.4]
  assign _T_56332 = $signed(_T_56331); // @[Modules.scala 40:46:@2231.4]
  assign _T_56334 = $signed(5'sh0) - $signed(io_in_770); // @[Modules.scala 43:37:@2233.4]
  assign _T_56335 = _T_56334[4:0]; // @[Modules.scala 43:37:@2234.4]
  assign _T_56336 = $signed(_T_56335); // @[Modules.scala 43:37:@2235.4]
  assign _T_56337 = $signed(_T_56336) + $signed(io_in_771); // @[Modules.scala 43:47:@2236.4]
  assign _T_56338 = _T_56337[4:0]; // @[Modules.scala 43:47:@2237.4]
  assign _T_56339 = $signed(_T_56338); // @[Modules.scala 43:47:@2238.4]
  assign _T_56341 = $signed(5'sh0) - $signed(io_in_772); // @[Modules.scala 46:37:@2240.4]
  assign _T_56342 = _T_56341[4:0]; // @[Modules.scala 46:37:@2241.4]
  assign _T_56343 = $signed(_T_56342); // @[Modules.scala 46:37:@2242.4]
  assign _T_56344 = $signed(_T_56343) - $signed(io_in_773); // @[Modules.scala 46:47:@2243.4]
  assign _T_56345 = _T_56344[4:0]; // @[Modules.scala 46:47:@2244.4]
  assign _T_56346 = $signed(_T_56345); // @[Modules.scala 46:47:@2245.4]
  assign _T_56348 = $signed(5'sh0) - $signed(io_in_774); // @[Modules.scala 46:37:@2247.4]
  assign _T_56349 = _T_56348[4:0]; // @[Modules.scala 46:37:@2248.4]
  assign _T_56350 = $signed(_T_56349); // @[Modules.scala 46:37:@2249.4]
  assign _T_56351 = $signed(_T_56350) - $signed(io_in_775); // @[Modules.scala 46:47:@2250.4]
  assign _T_56352 = _T_56351[4:0]; // @[Modules.scala 46:47:@2251.4]
  assign _T_56353 = $signed(_T_56352); // @[Modules.scala 46:47:@2252.4]
  assign _T_56354 = $signed(io_in_776) + $signed(io_in_777); // @[Modules.scala 37:46:@2254.4]
  assign _T_56355 = _T_56354[4:0]; // @[Modules.scala 37:46:@2255.4]
  assign _T_56356 = $signed(_T_56355); // @[Modules.scala 37:46:@2256.4]
  assign _T_56358 = $signed(5'sh0) - $signed(io_in_778); // @[Modules.scala 46:37:@2258.4]
  assign _T_56359 = _T_56358[4:0]; // @[Modules.scala 46:37:@2259.4]
  assign _T_56360 = $signed(_T_56359); // @[Modules.scala 46:37:@2260.4]
  assign _T_56361 = $signed(_T_56360) - $signed(io_in_779); // @[Modules.scala 46:47:@2261.4]
  assign _T_56362 = _T_56361[4:0]; // @[Modules.scala 46:47:@2262.4]
  assign _T_56363 = $signed(_T_56362); // @[Modules.scala 46:47:@2263.4]
  assign _T_56365 = $signed(5'sh0) - $signed(io_in_780); // @[Modules.scala 43:37:@2265.4]
  assign _T_56366 = _T_56365[4:0]; // @[Modules.scala 43:37:@2266.4]
  assign _T_56367 = $signed(_T_56366); // @[Modules.scala 43:37:@2267.4]
  assign _T_56368 = $signed(_T_56367) + $signed(io_in_781); // @[Modules.scala 43:47:@2268.4]
  assign _T_56369 = _T_56368[4:0]; // @[Modules.scala 43:47:@2269.4]
  assign _T_56370 = $signed(_T_56369); // @[Modules.scala 43:47:@2270.4]
  assign _T_56371 = $signed(io_in_782) + $signed(io_in_783); // @[Modules.scala 37:46:@2272.4]
  assign _T_56372 = _T_56371[4:0]; // @[Modules.scala 37:46:@2273.4]
  assign _T_56373 = $signed(_T_56372); // @[Modules.scala 37:46:@2274.4]
  assign buffer_0_0 = {{6{_T_54272[4]}},_T_54272}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_1 = {{6{_T_54279[4]}},_T_54279}; // @[Modules.scala 32:22:@8.4]
  assign _T_56374 = $signed(buffer_0_0) + $signed(buffer_0_1); // @[Modules.scala 50:57:@2276.4]
  assign _T_56375 = _T_56374[10:0]; // @[Modules.scala 50:57:@2277.4]
  assign buffer_0_392 = $signed(_T_56375); // @[Modules.scala 50:57:@2278.4]
  assign buffer_0_2 = {{6{_T_54286[4]}},_T_54286}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_3 = {{6{_T_54293[4]}},_T_54293}; // @[Modules.scala 32:22:@8.4]
  assign _T_56377 = $signed(buffer_0_2) + $signed(buffer_0_3); // @[Modules.scala 50:57:@2280.4]
  assign _T_56378 = _T_56377[10:0]; // @[Modules.scala 50:57:@2281.4]
  assign buffer_0_393 = $signed(_T_56378); // @[Modules.scala 50:57:@2282.4]
  assign buffer_0_4 = {{6{_T_54300[4]}},_T_54300}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_5 = {{6{_T_54307[4]}},_T_54307}; // @[Modules.scala 32:22:@8.4]
  assign _T_56380 = $signed(buffer_0_4) + $signed(buffer_0_5); // @[Modules.scala 50:57:@2284.4]
  assign _T_56381 = _T_56380[10:0]; // @[Modules.scala 50:57:@2285.4]
  assign buffer_0_394 = $signed(_T_56381); // @[Modules.scala 50:57:@2286.4]
  assign buffer_0_6 = {{6{_T_54314[4]}},_T_54314}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_7 = {{6{_T_54321[4]}},_T_54321}; // @[Modules.scala 32:22:@8.4]
  assign _T_56383 = $signed(buffer_0_6) + $signed(buffer_0_7); // @[Modules.scala 50:57:@2288.4]
  assign _T_56384 = _T_56383[10:0]; // @[Modules.scala 50:57:@2289.4]
  assign buffer_0_395 = $signed(_T_56384); // @[Modules.scala 50:57:@2290.4]
  assign buffer_0_8 = {{6{_T_54324[4]}},_T_54324}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_9 = {{6{_T_54331[4]}},_T_54331}; // @[Modules.scala 32:22:@8.4]
  assign _T_56386 = $signed(buffer_0_8) + $signed(buffer_0_9); // @[Modules.scala 50:57:@2292.4]
  assign _T_56387 = _T_56386[10:0]; // @[Modules.scala 50:57:@2293.4]
  assign buffer_0_396 = $signed(_T_56387); // @[Modules.scala 50:57:@2294.4]
  assign buffer_0_10 = {{6{_T_54334[4]}},_T_54334}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_11 = {{6{_T_54341[4]}},_T_54341}; // @[Modules.scala 32:22:@8.4]
  assign _T_56389 = $signed(buffer_0_10) + $signed(buffer_0_11); // @[Modules.scala 50:57:@2296.4]
  assign _T_56390 = _T_56389[10:0]; // @[Modules.scala 50:57:@2297.4]
  assign buffer_0_397 = $signed(_T_56390); // @[Modules.scala 50:57:@2298.4]
  assign buffer_0_12 = {{6{_T_54348[4]}},_T_54348}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_13 = {{6{_T_54351[4]}},_T_54351}; // @[Modules.scala 32:22:@8.4]
  assign _T_56392 = $signed(buffer_0_12) + $signed(buffer_0_13); // @[Modules.scala 50:57:@2300.4]
  assign _T_56393 = _T_56392[10:0]; // @[Modules.scala 50:57:@2301.4]
  assign buffer_0_398 = $signed(_T_56393); // @[Modules.scala 50:57:@2302.4]
  assign buffer_0_14 = {{6{_T_54358[4]}},_T_54358}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_15 = {{6{_T_54365[4]}},_T_54365}; // @[Modules.scala 32:22:@8.4]
  assign _T_56395 = $signed(buffer_0_14) + $signed(buffer_0_15); // @[Modules.scala 50:57:@2304.4]
  assign _T_56396 = _T_56395[10:0]; // @[Modules.scala 50:57:@2305.4]
  assign buffer_0_399 = $signed(_T_56396); // @[Modules.scala 50:57:@2306.4]
  assign buffer_0_16 = {{6{_T_54368[4]}},_T_54368}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_17 = {{6{_T_54375[4]}},_T_54375}; // @[Modules.scala 32:22:@8.4]
  assign _T_56398 = $signed(buffer_0_16) + $signed(buffer_0_17); // @[Modules.scala 50:57:@2308.4]
  assign _T_56399 = _T_56398[10:0]; // @[Modules.scala 50:57:@2309.4]
  assign buffer_0_400 = $signed(_T_56399); // @[Modules.scala 50:57:@2310.4]
  assign buffer_0_18 = {{6{_T_54382[4]}},_T_54382}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_19 = {{6{_T_54389[4]}},_T_54389}; // @[Modules.scala 32:22:@8.4]
  assign _T_56401 = $signed(buffer_0_18) + $signed(buffer_0_19); // @[Modules.scala 50:57:@2312.4]
  assign _T_56402 = _T_56401[10:0]; // @[Modules.scala 50:57:@2313.4]
  assign buffer_0_401 = $signed(_T_56402); // @[Modules.scala 50:57:@2314.4]
  assign buffer_0_20 = {{6{_T_54396[4]}},_T_54396}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_21 = {{6{_T_54403[4]}},_T_54403}; // @[Modules.scala 32:22:@8.4]
  assign _T_56404 = $signed(buffer_0_20) + $signed(buffer_0_21); // @[Modules.scala 50:57:@2316.4]
  assign _T_56405 = _T_56404[10:0]; // @[Modules.scala 50:57:@2317.4]
  assign buffer_0_402 = $signed(_T_56405); // @[Modules.scala 50:57:@2318.4]
  assign buffer_0_22 = {{6{_T_54410[4]}},_T_54410}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_23 = {{6{_T_54417[4]}},_T_54417}; // @[Modules.scala 32:22:@8.4]
  assign _T_56407 = $signed(buffer_0_22) + $signed(buffer_0_23); // @[Modules.scala 50:57:@2320.4]
  assign _T_56408 = _T_56407[10:0]; // @[Modules.scala 50:57:@2321.4]
  assign buffer_0_403 = $signed(_T_56408); // @[Modules.scala 50:57:@2322.4]
  assign buffer_0_24 = {{6{_T_54424[4]}},_T_54424}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_25 = {{6{_T_54431[4]}},_T_54431}; // @[Modules.scala 32:22:@8.4]
  assign _T_56410 = $signed(buffer_0_24) + $signed(buffer_0_25); // @[Modules.scala 50:57:@2324.4]
  assign _T_56411 = _T_56410[10:0]; // @[Modules.scala 50:57:@2325.4]
  assign buffer_0_404 = $signed(_T_56411); // @[Modules.scala 50:57:@2326.4]
  assign buffer_0_26 = {{6{_T_54434[4]}},_T_54434}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_27 = {{6{_T_54437[4]}},_T_54437}; // @[Modules.scala 32:22:@8.4]
  assign _T_56413 = $signed(buffer_0_26) + $signed(buffer_0_27); // @[Modules.scala 50:57:@2328.4]
  assign _T_56414 = _T_56413[10:0]; // @[Modules.scala 50:57:@2329.4]
  assign buffer_0_405 = $signed(_T_56414); // @[Modules.scala 50:57:@2330.4]
  assign buffer_0_28 = {{6{_T_54440[4]}},_T_54440}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_29 = {{6{_T_54447[4]}},_T_54447}; // @[Modules.scala 32:22:@8.4]
  assign _T_56416 = $signed(buffer_0_28) + $signed(buffer_0_29); // @[Modules.scala 50:57:@2332.4]
  assign _T_56417 = _T_56416[10:0]; // @[Modules.scala 50:57:@2333.4]
  assign buffer_0_406 = $signed(_T_56417); // @[Modules.scala 50:57:@2334.4]
  assign buffer_0_30 = {{6{_T_54454[4]}},_T_54454}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_31 = {{6{_T_54461[4]}},_T_54461}; // @[Modules.scala 32:22:@8.4]
  assign _T_56419 = $signed(buffer_0_30) + $signed(buffer_0_31); // @[Modules.scala 50:57:@2336.4]
  assign _T_56420 = _T_56419[10:0]; // @[Modules.scala 50:57:@2337.4]
  assign buffer_0_407 = $signed(_T_56420); // @[Modules.scala 50:57:@2338.4]
  assign buffer_0_32 = {{6{_T_54468[4]}},_T_54468}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_33 = {{6{_T_54475[4]}},_T_54475}; // @[Modules.scala 32:22:@8.4]
  assign _T_56422 = $signed(buffer_0_32) + $signed(buffer_0_33); // @[Modules.scala 50:57:@2340.4]
  assign _T_56423 = _T_56422[10:0]; // @[Modules.scala 50:57:@2341.4]
  assign buffer_0_408 = $signed(_T_56423); // @[Modules.scala 50:57:@2342.4]
  assign buffer_0_34 = {{6{_T_54482[4]}},_T_54482}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_35 = {{6{_T_54489[4]}},_T_54489}; // @[Modules.scala 32:22:@8.4]
  assign _T_56425 = $signed(buffer_0_34) + $signed(buffer_0_35); // @[Modules.scala 50:57:@2344.4]
  assign _T_56426 = _T_56425[10:0]; // @[Modules.scala 50:57:@2345.4]
  assign buffer_0_409 = $signed(_T_56426); // @[Modules.scala 50:57:@2346.4]
  assign buffer_0_36 = {{6{_T_54496[4]}},_T_54496}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_37 = {{6{_T_54503[4]}},_T_54503}; // @[Modules.scala 32:22:@8.4]
  assign _T_56428 = $signed(buffer_0_36) + $signed(buffer_0_37); // @[Modules.scala 50:57:@2348.4]
  assign _T_56429 = _T_56428[10:0]; // @[Modules.scala 50:57:@2349.4]
  assign buffer_0_410 = $signed(_T_56429); // @[Modules.scala 50:57:@2350.4]
  assign buffer_0_38 = {{6{_T_54506[4]}},_T_54506}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_39 = {{6{_T_54509[4]}},_T_54509}; // @[Modules.scala 32:22:@8.4]
  assign _T_56431 = $signed(buffer_0_38) + $signed(buffer_0_39); // @[Modules.scala 50:57:@2352.4]
  assign _T_56432 = _T_56431[10:0]; // @[Modules.scala 50:57:@2353.4]
  assign buffer_0_411 = $signed(_T_56432); // @[Modules.scala 50:57:@2354.4]
  assign buffer_0_40 = {{6{_T_54516[4]}},_T_54516}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_41 = {{6{_T_54519[4]}},_T_54519}; // @[Modules.scala 32:22:@8.4]
  assign _T_56434 = $signed(buffer_0_40) + $signed(buffer_0_41); // @[Modules.scala 50:57:@2356.4]
  assign _T_56435 = _T_56434[10:0]; // @[Modules.scala 50:57:@2357.4]
  assign buffer_0_412 = $signed(_T_56435); // @[Modules.scala 50:57:@2358.4]
  assign buffer_0_42 = {{6{_T_54522[4]}},_T_54522}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_43 = {{6{_T_54529[4]}},_T_54529}; // @[Modules.scala 32:22:@8.4]
  assign _T_56437 = $signed(buffer_0_42) + $signed(buffer_0_43); // @[Modules.scala 50:57:@2360.4]
  assign _T_56438 = _T_56437[10:0]; // @[Modules.scala 50:57:@2361.4]
  assign buffer_0_413 = $signed(_T_56438); // @[Modules.scala 50:57:@2362.4]
  assign buffer_0_44 = {{6{_T_54532[4]}},_T_54532}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_45 = {{6{_T_54535[4]}},_T_54535}; // @[Modules.scala 32:22:@8.4]
  assign _T_56440 = $signed(buffer_0_44) + $signed(buffer_0_45); // @[Modules.scala 50:57:@2364.4]
  assign _T_56441 = _T_56440[10:0]; // @[Modules.scala 50:57:@2365.4]
  assign buffer_0_414 = $signed(_T_56441); // @[Modules.scala 50:57:@2366.4]
  assign buffer_0_46 = {{6{_T_54542[4]}},_T_54542}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_47 = {{6{_T_54545[4]}},_T_54545}; // @[Modules.scala 32:22:@8.4]
  assign _T_56443 = $signed(buffer_0_46) + $signed(buffer_0_47); // @[Modules.scala 50:57:@2368.4]
  assign _T_56444 = _T_56443[10:0]; // @[Modules.scala 50:57:@2369.4]
  assign buffer_0_415 = $signed(_T_56444); // @[Modules.scala 50:57:@2370.4]
  assign buffer_0_48 = {{6{_T_54552[4]}},_T_54552}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_49 = {{6{_T_54555[4]}},_T_54555}; // @[Modules.scala 32:22:@8.4]
  assign _T_56446 = $signed(buffer_0_48) + $signed(buffer_0_49); // @[Modules.scala 50:57:@2372.4]
  assign _T_56447 = _T_56446[10:0]; // @[Modules.scala 50:57:@2373.4]
  assign buffer_0_416 = $signed(_T_56447); // @[Modules.scala 50:57:@2374.4]
  assign buffer_0_50 = {{6{_T_54558[4]}},_T_54558}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_51 = {{6{_T_54561[4]}},_T_54561}; // @[Modules.scala 32:22:@8.4]
  assign _T_56449 = $signed(buffer_0_50) + $signed(buffer_0_51); // @[Modules.scala 50:57:@2376.4]
  assign _T_56450 = _T_56449[10:0]; // @[Modules.scala 50:57:@2377.4]
  assign buffer_0_417 = $signed(_T_56450); // @[Modules.scala 50:57:@2378.4]
  assign buffer_0_52 = {{6{_T_54564[4]}},_T_54564}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_53 = {{6{_T_54567[4]}},_T_54567}; // @[Modules.scala 32:22:@8.4]
  assign _T_56452 = $signed(buffer_0_52) + $signed(buffer_0_53); // @[Modules.scala 50:57:@2380.4]
  assign _T_56453 = _T_56452[10:0]; // @[Modules.scala 50:57:@2381.4]
  assign buffer_0_418 = $signed(_T_56453); // @[Modules.scala 50:57:@2382.4]
  assign buffer_0_54 = {{6{_T_54570[4]}},_T_54570}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_55 = {{6{_T_54573[4]}},_T_54573}; // @[Modules.scala 32:22:@8.4]
  assign _T_56455 = $signed(buffer_0_54) + $signed(buffer_0_55); // @[Modules.scala 50:57:@2384.4]
  assign _T_56456 = _T_56455[10:0]; // @[Modules.scala 50:57:@2385.4]
  assign buffer_0_419 = $signed(_T_56456); // @[Modules.scala 50:57:@2386.4]
  assign buffer_0_56 = {{6{_T_54580[4]}},_T_54580}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_57 = {{6{_T_54587[4]}},_T_54587}; // @[Modules.scala 32:22:@8.4]
  assign _T_56458 = $signed(buffer_0_56) + $signed(buffer_0_57); // @[Modules.scala 50:57:@2388.4]
  assign _T_56459 = _T_56458[10:0]; // @[Modules.scala 50:57:@2389.4]
  assign buffer_0_420 = $signed(_T_56459); // @[Modules.scala 50:57:@2390.4]
  assign buffer_0_58 = {{6{_T_54590[4]}},_T_54590}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_59 = {{6{_T_54593[4]}},_T_54593}; // @[Modules.scala 32:22:@8.4]
  assign _T_56461 = $signed(buffer_0_58) + $signed(buffer_0_59); // @[Modules.scala 50:57:@2392.4]
  assign _T_56462 = _T_56461[10:0]; // @[Modules.scala 50:57:@2393.4]
  assign buffer_0_421 = $signed(_T_56462); // @[Modules.scala 50:57:@2394.4]
  assign buffer_0_60 = {{6{_T_54600[4]}},_T_54600}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_61 = {{6{_T_54607[4]}},_T_54607}; // @[Modules.scala 32:22:@8.4]
  assign _T_56464 = $signed(buffer_0_60) + $signed(buffer_0_61); // @[Modules.scala 50:57:@2396.4]
  assign _T_56465 = _T_56464[10:0]; // @[Modules.scala 50:57:@2397.4]
  assign buffer_0_422 = $signed(_T_56465); // @[Modules.scala 50:57:@2398.4]
  assign buffer_0_62 = {{6{_T_54614[4]}},_T_54614}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_63 = {{6{_T_54621[4]}},_T_54621}; // @[Modules.scala 32:22:@8.4]
  assign _T_56467 = $signed(buffer_0_62) + $signed(buffer_0_63); // @[Modules.scala 50:57:@2400.4]
  assign _T_56468 = _T_56467[10:0]; // @[Modules.scala 50:57:@2401.4]
  assign buffer_0_423 = $signed(_T_56468); // @[Modules.scala 50:57:@2402.4]
  assign buffer_0_64 = {{6{_T_54628[4]}},_T_54628}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_65 = {{6{_T_54635[4]}},_T_54635}; // @[Modules.scala 32:22:@8.4]
  assign _T_56470 = $signed(buffer_0_64) + $signed(buffer_0_65); // @[Modules.scala 50:57:@2404.4]
  assign _T_56471 = _T_56470[10:0]; // @[Modules.scala 50:57:@2405.4]
  assign buffer_0_424 = $signed(_T_56471); // @[Modules.scala 50:57:@2406.4]
  assign buffer_0_66 = {{6{_T_54638[4]}},_T_54638}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_67 = {{6{_T_54641[4]}},_T_54641}; // @[Modules.scala 32:22:@8.4]
  assign _T_56473 = $signed(buffer_0_66) + $signed(buffer_0_67); // @[Modules.scala 50:57:@2408.4]
  assign _T_56474 = _T_56473[10:0]; // @[Modules.scala 50:57:@2409.4]
  assign buffer_0_425 = $signed(_T_56474); // @[Modules.scala 50:57:@2410.4]
  assign buffer_0_68 = {{6{_T_54644[4]}},_T_54644}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_69 = {{6{_T_54651[4]}},_T_54651}; // @[Modules.scala 32:22:@8.4]
  assign _T_56476 = $signed(buffer_0_68) + $signed(buffer_0_69); // @[Modules.scala 50:57:@2412.4]
  assign _T_56477 = _T_56476[10:0]; // @[Modules.scala 50:57:@2413.4]
  assign buffer_0_426 = $signed(_T_56477); // @[Modules.scala 50:57:@2414.4]
  assign buffer_0_70 = {{6{_T_54654[4]}},_T_54654}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_71 = {{6{_T_54661[4]}},_T_54661}; // @[Modules.scala 32:22:@8.4]
  assign _T_56479 = $signed(buffer_0_70) + $signed(buffer_0_71); // @[Modules.scala 50:57:@2416.4]
  assign _T_56480 = _T_56479[10:0]; // @[Modules.scala 50:57:@2417.4]
  assign buffer_0_427 = $signed(_T_56480); // @[Modules.scala 50:57:@2418.4]
  assign buffer_0_72 = {{6{_T_54664[4]}},_T_54664}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_73 = {{6{_T_54667[4]}},_T_54667}; // @[Modules.scala 32:22:@8.4]
  assign _T_56482 = $signed(buffer_0_72) + $signed(buffer_0_73); // @[Modules.scala 50:57:@2420.4]
  assign _T_56483 = _T_56482[10:0]; // @[Modules.scala 50:57:@2421.4]
  assign buffer_0_428 = $signed(_T_56483); // @[Modules.scala 50:57:@2422.4]
  assign buffer_0_74 = {{6{_T_54670[4]}},_T_54670}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_75 = {{6{_T_54677[4]}},_T_54677}; // @[Modules.scala 32:22:@8.4]
  assign _T_56485 = $signed(buffer_0_74) + $signed(buffer_0_75); // @[Modules.scala 50:57:@2424.4]
  assign _T_56486 = _T_56485[10:0]; // @[Modules.scala 50:57:@2425.4]
  assign buffer_0_429 = $signed(_T_56486); // @[Modules.scala 50:57:@2426.4]
  assign buffer_0_76 = {{6{_T_54684[4]}},_T_54684}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_77 = {{6{_T_54691[4]}},_T_54691}; // @[Modules.scala 32:22:@8.4]
  assign _T_56488 = $signed(buffer_0_76) + $signed(buffer_0_77); // @[Modules.scala 50:57:@2428.4]
  assign _T_56489 = _T_56488[10:0]; // @[Modules.scala 50:57:@2429.4]
  assign buffer_0_430 = $signed(_T_56489); // @[Modules.scala 50:57:@2430.4]
  assign buffer_0_78 = {{6{_T_54698[4]}},_T_54698}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_79 = {{6{_T_54705[4]}},_T_54705}; // @[Modules.scala 32:22:@8.4]
  assign _T_56491 = $signed(buffer_0_78) + $signed(buffer_0_79); // @[Modules.scala 50:57:@2432.4]
  assign _T_56492 = _T_56491[10:0]; // @[Modules.scala 50:57:@2433.4]
  assign buffer_0_431 = $signed(_T_56492); // @[Modules.scala 50:57:@2434.4]
  assign buffer_0_80 = {{6{_T_54712[4]}},_T_54712}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_81 = {{6{_T_54715[4]}},_T_54715}; // @[Modules.scala 32:22:@8.4]
  assign _T_56494 = $signed(buffer_0_80) + $signed(buffer_0_81); // @[Modules.scala 50:57:@2436.4]
  assign _T_56495 = _T_56494[10:0]; // @[Modules.scala 50:57:@2437.4]
  assign buffer_0_432 = $signed(_T_56495); // @[Modules.scala 50:57:@2438.4]
  assign buffer_0_82 = {{6{_T_54718[4]}},_T_54718}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_83 = {{6{_T_54725[4]}},_T_54725}; // @[Modules.scala 32:22:@8.4]
  assign _T_56497 = $signed(buffer_0_82) + $signed(buffer_0_83); // @[Modules.scala 50:57:@2440.4]
  assign _T_56498 = _T_56497[10:0]; // @[Modules.scala 50:57:@2441.4]
  assign buffer_0_433 = $signed(_T_56498); // @[Modules.scala 50:57:@2442.4]
  assign buffer_0_84 = {{6{_T_54732[4]}},_T_54732}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_85 = {{6{_T_54739[4]}},_T_54739}; // @[Modules.scala 32:22:@8.4]
  assign _T_56500 = $signed(buffer_0_84) + $signed(buffer_0_85); // @[Modules.scala 50:57:@2444.4]
  assign _T_56501 = _T_56500[10:0]; // @[Modules.scala 50:57:@2445.4]
  assign buffer_0_434 = $signed(_T_56501); // @[Modules.scala 50:57:@2446.4]
  assign buffer_0_86 = {{6{_T_54742[4]}},_T_54742}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_87 = {{6{_T_54749[4]}},_T_54749}; // @[Modules.scala 32:22:@8.4]
  assign _T_56503 = $signed(buffer_0_86) + $signed(buffer_0_87); // @[Modules.scala 50:57:@2448.4]
  assign _T_56504 = _T_56503[10:0]; // @[Modules.scala 50:57:@2449.4]
  assign buffer_0_435 = $signed(_T_56504); // @[Modules.scala 50:57:@2450.4]
  assign buffer_0_88 = {{6{_T_54756[4]}},_T_54756}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_89 = {{6{_T_54763[4]}},_T_54763}; // @[Modules.scala 32:22:@8.4]
  assign _T_56506 = $signed(buffer_0_88) + $signed(buffer_0_89); // @[Modules.scala 50:57:@2452.4]
  assign _T_56507 = _T_56506[10:0]; // @[Modules.scala 50:57:@2453.4]
  assign buffer_0_436 = $signed(_T_56507); // @[Modules.scala 50:57:@2454.4]
  assign buffer_0_90 = {{6{_T_54770[4]}},_T_54770}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_91 = {{6{_T_54777[4]}},_T_54777}; // @[Modules.scala 32:22:@8.4]
  assign _T_56509 = $signed(buffer_0_90) + $signed(buffer_0_91); // @[Modules.scala 50:57:@2456.4]
  assign _T_56510 = _T_56509[10:0]; // @[Modules.scala 50:57:@2457.4]
  assign buffer_0_437 = $signed(_T_56510); // @[Modules.scala 50:57:@2458.4]
  assign buffer_0_92 = {{6{_T_54784[4]}},_T_54784}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_93 = {{6{_T_54787[4]}},_T_54787}; // @[Modules.scala 32:22:@8.4]
  assign _T_56512 = $signed(buffer_0_92) + $signed(buffer_0_93); // @[Modules.scala 50:57:@2460.4]
  assign _T_56513 = _T_56512[10:0]; // @[Modules.scala 50:57:@2461.4]
  assign buffer_0_438 = $signed(_T_56513); // @[Modules.scala 50:57:@2462.4]
  assign buffer_0_94 = {{6{_T_54794[4]}},_T_54794}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_95 = {{6{_T_54797[4]}},_T_54797}; // @[Modules.scala 32:22:@8.4]
  assign _T_56515 = $signed(buffer_0_94) + $signed(buffer_0_95); // @[Modules.scala 50:57:@2464.4]
  assign _T_56516 = _T_56515[10:0]; // @[Modules.scala 50:57:@2465.4]
  assign buffer_0_439 = $signed(_T_56516); // @[Modules.scala 50:57:@2466.4]
  assign buffer_0_96 = {{6{_T_54804[4]}},_T_54804}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_97 = {{6{_T_54811[4]}},_T_54811}; // @[Modules.scala 32:22:@8.4]
  assign _T_56518 = $signed(buffer_0_96) + $signed(buffer_0_97); // @[Modules.scala 50:57:@2468.4]
  assign _T_56519 = _T_56518[10:0]; // @[Modules.scala 50:57:@2469.4]
  assign buffer_0_440 = $signed(_T_56519); // @[Modules.scala 50:57:@2470.4]
  assign buffer_0_98 = {{6{_T_54814[4]}},_T_54814}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_99 = {{6{_T_54817[4]}},_T_54817}; // @[Modules.scala 32:22:@8.4]
  assign _T_56521 = $signed(buffer_0_98) + $signed(buffer_0_99); // @[Modules.scala 50:57:@2472.4]
  assign _T_56522 = _T_56521[10:0]; // @[Modules.scala 50:57:@2473.4]
  assign buffer_0_441 = $signed(_T_56522); // @[Modules.scala 50:57:@2474.4]
  assign buffer_0_100 = {{6{_T_54824[4]}},_T_54824}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_101 = {{6{_T_54831[4]}},_T_54831}; // @[Modules.scala 32:22:@8.4]
  assign _T_56524 = $signed(buffer_0_100) + $signed(buffer_0_101); // @[Modules.scala 50:57:@2476.4]
  assign _T_56525 = _T_56524[10:0]; // @[Modules.scala 50:57:@2477.4]
  assign buffer_0_442 = $signed(_T_56525); // @[Modules.scala 50:57:@2478.4]
  assign buffer_0_102 = {{6{_T_54838[4]}},_T_54838}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_103 = {{6{_T_54845[4]}},_T_54845}; // @[Modules.scala 32:22:@8.4]
  assign _T_56527 = $signed(buffer_0_102) + $signed(buffer_0_103); // @[Modules.scala 50:57:@2480.4]
  assign _T_56528 = _T_56527[10:0]; // @[Modules.scala 50:57:@2481.4]
  assign buffer_0_443 = $signed(_T_56528); // @[Modules.scala 50:57:@2482.4]
  assign buffer_0_104 = {{6{_T_54852[4]}},_T_54852}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_105 = {{6{_T_54855[4]}},_T_54855}; // @[Modules.scala 32:22:@8.4]
  assign _T_56530 = $signed(buffer_0_104) + $signed(buffer_0_105); // @[Modules.scala 50:57:@2484.4]
  assign _T_56531 = _T_56530[10:0]; // @[Modules.scala 50:57:@2485.4]
  assign buffer_0_444 = $signed(_T_56531); // @[Modules.scala 50:57:@2486.4]
  assign buffer_0_106 = {{6{_T_54858[4]}},_T_54858}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_107 = {{6{_T_54865[4]}},_T_54865}; // @[Modules.scala 32:22:@8.4]
  assign _T_56533 = $signed(buffer_0_106) + $signed(buffer_0_107); // @[Modules.scala 50:57:@2488.4]
  assign _T_56534 = _T_56533[10:0]; // @[Modules.scala 50:57:@2489.4]
  assign buffer_0_445 = $signed(_T_56534); // @[Modules.scala 50:57:@2490.4]
  assign buffer_0_108 = {{6{_T_54872[4]}},_T_54872}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_109 = {{6{_T_54879[4]}},_T_54879}; // @[Modules.scala 32:22:@8.4]
  assign _T_56536 = $signed(buffer_0_108) + $signed(buffer_0_109); // @[Modules.scala 50:57:@2492.4]
  assign _T_56537 = _T_56536[10:0]; // @[Modules.scala 50:57:@2493.4]
  assign buffer_0_446 = $signed(_T_56537); // @[Modules.scala 50:57:@2494.4]
  assign buffer_0_110 = {{6{_T_54886[4]}},_T_54886}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_111 = {{6{_T_54893[4]}},_T_54893}; // @[Modules.scala 32:22:@8.4]
  assign _T_56539 = $signed(buffer_0_110) + $signed(buffer_0_111); // @[Modules.scala 50:57:@2496.4]
  assign _T_56540 = _T_56539[10:0]; // @[Modules.scala 50:57:@2497.4]
  assign buffer_0_447 = $signed(_T_56540); // @[Modules.scala 50:57:@2498.4]
  assign buffer_0_112 = {{6{_T_54900[4]}},_T_54900}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_113 = {{6{_T_54907[4]}},_T_54907}; // @[Modules.scala 32:22:@8.4]
  assign _T_56542 = $signed(buffer_0_112) + $signed(buffer_0_113); // @[Modules.scala 50:57:@2500.4]
  assign _T_56543 = _T_56542[10:0]; // @[Modules.scala 50:57:@2501.4]
  assign buffer_0_448 = $signed(_T_56543); // @[Modules.scala 50:57:@2502.4]
  assign buffer_0_114 = {{6{_T_54914[4]}},_T_54914}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_115 = {{6{_T_54921[4]}},_T_54921}; // @[Modules.scala 32:22:@8.4]
  assign _T_56545 = $signed(buffer_0_114) + $signed(buffer_0_115); // @[Modules.scala 50:57:@2504.4]
  assign _T_56546 = _T_56545[10:0]; // @[Modules.scala 50:57:@2505.4]
  assign buffer_0_449 = $signed(_T_56546); // @[Modules.scala 50:57:@2506.4]
  assign buffer_0_116 = {{6{_T_54928[4]}},_T_54928}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_117 = {{6{_T_54935[4]}},_T_54935}; // @[Modules.scala 32:22:@8.4]
  assign _T_56548 = $signed(buffer_0_116) + $signed(buffer_0_117); // @[Modules.scala 50:57:@2508.4]
  assign _T_56549 = _T_56548[10:0]; // @[Modules.scala 50:57:@2509.4]
  assign buffer_0_450 = $signed(_T_56549); // @[Modules.scala 50:57:@2510.4]
  assign buffer_0_118 = {{6{_T_54942[4]}},_T_54942}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_119 = {{6{_T_54949[4]}},_T_54949}; // @[Modules.scala 32:22:@8.4]
  assign _T_56551 = $signed(buffer_0_118) + $signed(buffer_0_119); // @[Modules.scala 50:57:@2512.4]
  assign _T_56552 = _T_56551[10:0]; // @[Modules.scala 50:57:@2513.4]
  assign buffer_0_451 = $signed(_T_56552); // @[Modules.scala 50:57:@2514.4]
  assign buffer_0_120 = {{6{_T_54956[4]}},_T_54956}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_121 = {{6{_T_54963[4]}},_T_54963}; // @[Modules.scala 32:22:@8.4]
  assign _T_56554 = $signed(buffer_0_120) + $signed(buffer_0_121); // @[Modules.scala 50:57:@2516.4]
  assign _T_56555 = _T_56554[10:0]; // @[Modules.scala 50:57:@2517.4]
  assign buffer_0_452 = $signed(_T_56555); // @[Modules.scala 50:57:@2518.4]
  assign buffer_0_122 = {{6{_T_54970[4]}},_T_54970}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_123 = {{6{_T_54977[4]}},_T_54977}; // @[Modules.scala 32:22:@8.4]
  assign _T_56557 = $signed(buffer_0_122) + $signed(buffer_0_123); // @[Modules.scala 50:57:@2520.4]
  assign _T_56558 = _T_56557[10:0]; // @[Modules.scala 50:57:@2521.4]
  assign buffer_0_453 = $signed(_T_56558); // @[Modules.scala 50:57:@2522.4]
  assign buffer_0_124 = {{6{_T_54984[4]}},_T_54984}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_125 = {{6{_T_54991[4]}},_T_54991}; // @[Modules.scala 32:22:@8.4]
  assign _T_56560 = $signed(buffer_0_124) + $signed(buffer_0_125); // @[Modules.scala 50:57:@2524.4]
  assign _T_56561 = _T_56560[10:0]; // @[Modules.scala 50:57:@2525.4]
  assign buffer_0_454 = $signed(_T_56561); // @[Modules.scala 50:57:@2526.4]
  assign buffer_0_126 = {{6{_T_54998[4]}},_T_54998}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_127 = {{6{_T_55005[4]}},_T_55005}; // @[Modules.scala 32:22:@8.4]
  assign _T_56563 = $signed(buffer_0_126) + $signed(buffer_0_127); // @[Modules.scala 50:57:@2528.4]
  assign _T_56564 = _T_56563[10:0]; // @[Modules.scala 50:57:@2529.4]
  assign buffer_0_455 = $signed(_T_56564); // @[Modules.scala 50:57:@2530.4]
  assign buffer_0_128 = {{6{_T_55012[4]}},_T_55012}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_129 = {{6{_T_55019[4]}},_T_55019}; // @[Modules.scala 32:22:@8.4]
  assign _T_56566 = $signed(buffer_0_128) + $signed(buffer_0_129); // @[Modules.scala 50:57:@2532.4]
  assign _T_56567 = _T_56566[10:0]; // @[Modules.scala 50:57:@2533.4]
  assign buffer_0_456 = $signed(_T_56567); // @[Modules.scala 50:57:@2534.4]
  assign buffer_0_130 = {{6{_T_55026[4]}},_T_55026}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_131 = {{6{_T_55029[4]}},_T_55029}; // @[Modules.scala 32:22:@8.4]
  assign _T_56569 = $signed(buffer_0_130) + $signed(buffer_0_131); // @[Modules.scala 50:57:@2536.4]
  assign _T_56570 = _T_56569[10:0]; // @[Modules.scala 50:57:@2537.4]
  assign buffer_0_457 = $signed(_T_56570); // @[Modules.scala 50:57:@2538.4]
  assign buffer_0_132 = {{6{_T_55036[4]}},_T_55036}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_133 = {{6{_T_55043[4]}},_T_55043}; // @[Modules.scala 32:22:@8.4]
  assign _T_56572 = $signed(buffer_0_132) + $signed(buffer_0_133); // @[Modules.scala 50:57:@2540.4]
  assign _T_56573 = _T_56572[10:0]; // @[Modules.scala 50:57:@2541.4]
  assign buffer_0_458 = $signed(_T_56573); // @[Modules.scala 50:57:@2542.4]
  assign buffer_0_134 = {{6{_T_55050[4]}},_T_55050}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_135 = {{6{_T_55057[4]}},_T_55057}; // @[Modules.scala 32:22:@8.4]
  assign _T_56575 = $signed(buffer_0_134) + $signed(buffer_0_135); // @[Modules.scala 50:57:@2544.4]
  assign _T_56576 = _T_56575[10:0]; // @[Modules.scala 50:57:@2545.4]
  assign buffer_0_459 = $signed(_T_56576); // @[Modules.scala 50:57:@2546.4]
  assign buffer_0_136 = {{6{_T_55064[4]}},_T_55064}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_137 = {{6{_T_55071[4]}},_T_55071}; // @[Modules.scala 32:22:@8.4]
  assign _T_56578 = $signed(buffer_0_136) + $signed(buffer_0_137); // @[Modules.scala 50:57:@2548.4]
  assign _T_56579 = _T_56578[10:0]; // @[Modules.scala 50:57:@2549.4]
  assign buffer_0_460 = $signed(_T_56579); // @[Modules.scala 50:57:@2550.4]
  assign buffer_0_138 = {{6{_T_55078[4]}},_T_55078}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_139 = {{6{_T_55085[4]}},_T_55085}; // @[Modules.scala 32:22:@8.4]
  assign _T_56581 = $signed(buffer_0_138) + $signed(buffer_0_139); // @[Modules.scala 50:57:@2552.4]
  assign _T_56582 = _T_56581[10:0]; // @[Modules.scala 50:57:@2553.4]
  assign buffer_0_461 = $signed(_T_56582); // @[Modules.scala 50:57:@2554.4]
  assign buffer_0_140 = {{6{_T_55092[4]}},_T_55092}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_141 = {{6{_T_55099[4]}},_T_55099}; // @[Modules.scala 32:22:@8.4]
  assign _T_56584 = $signed(buffer_0_140) + $signed(buffer_0_141); // @[Modules.scala 50:57:@2556.4]
  assign _T_56585 = _T_56584[10:0]; // @[Modules.scala 50:57:@2557.4]
  assign buffer_0_462 = $signed(_T_56585); // @[Modules.scala 50:57:@2558.4]
  assign buffer_0_142 = {{6{_T_55106[4]}},_T_55106}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_143 = {{6{_T_55113[4]}},_T_55113}; // @[Modules.scala 32:22:@8.4]
  assign _T_56587 = $signed(buffer_0_142) + $signed(buffer_0_143); // @[Modules.scala 50:57:@2560.4]
  assign _T_56588 = _T_56587[10:0]; // @[Modules.scala 50:57:@2561.4]
  assign buffer_0_463 = $signed(_T_56588); // @[Modules.scala 50:57:@2562.4]
  assign buffer_0_144 = {{6{_T_55120[4]}},_T_55120}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_145 = {{6{_T_55127[4]}},_T_55127}; // @[Modules.scala 32:22:@8.4]
  assign _T_56590 = $signed(buffer_0_144) + $signed(buffer_0_145); // @[Modules.scala 50:57:@2564.4]
  assign _T_56591 = _T_56590[10:0]; // @[Modules.scala 50:57:@2565.4]
  assign buffer_0_464 = $signed(_T_56591); // @[Modules.scala 50:57:@2566.4]
  assign buffer_0_146 = {{6{_T_55134[4]}},_T_55134}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_147 = {{6{_T_55141[4]}},_T_55141}; // @[Modules.scala 32:22:@8.4]
  assign _T_56593 = $signed(buffer_0_146) + $signed(buffer_0_147); // @[Modules.scala 50:57:@2568.4]
  assign _T_56594 = _T_56593[10:0]; // @[Modules.scala 50:57:@2569.4]
  assign buffer_0_465 = $signed(_T_56594); // @[Modules.scala 50:57:@2570.4]
  assign buffer_0_148 = {{6{_T_55148[4]}},_T_55148}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_149 = {{6{_T_55155[4]}},_T_55155}; // @[Modules.scala 32:22:@8.4]
  assign _T_56596 = $signed(buffer_0_148) + $signed(buffer_0_149); // @[Modules.scala 50:57:@2572.4]
  assign _T_56597 = _T_56596[10:0]; // @[Modules.scala 50:57:@2573.4]
  assign buffer_0_466 = $signed(_T_56597); // @[Modules.scala 50:57:@2574.4]
  assign buffer_0_150 = {{6{_T_55162[4]}},_T_55162}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_151 = {{6{_T_55169[4]}},_T_55169}; // @[Modules.scala 32:22:@8.4]
  assign _T_56599 = $signed(buffer_0_150) + $signed(buffer_0_151); // @[Modules.scala 50:57:@2576.4]
  assign _T_56600 = _T_56599[10:0]; // @[Modules.scala 50:57:@2577.4]
  assign buffer_0_467 = $signed(_T_56600); // @[Modules.scala 50:57:@2578.4]
  assign buffer_0_152 = {{6{_T_55176[4]}},_T_55176}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_153 = {{6{_T_55183[4]}},_T_55183}; // @[Modules.scala 32:22:@8.4]
  assign _T_56602 = $signed(buffer_0_152) + $signed(buffer_0_153); // @[Modules.scala 50:57:@2580.4]
  assign _T_56603 = _T_56602[10:0]; // @[Modules.scala 50:57:@2581.4]
  assign buffer_0_468 = $signed(_T_56603); // @[Modules.scala 50:57:@2582.4]
  assign buffer_0_154 = {{6{_T_55190[4]}},_T_55190}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_155 = {{6{_T_55197[4]}},_T_55197}; // @[Modules.scala 32:22:@8.4]
  assign _T_56605 = $signed(buffer_0_154) + $signed(buffer_0_155); // @[Modules.scala 50:57:@2584.4]
  assign _T_56606 = _T_56605[10:0]; // @[Modules.scala 50:57:@2585.4]
  assign buffer_0_469 = $signed(_T_56606); // @[Modules.scala 50:57:@2586.4]
  assign buffer_0_156 = {{6{_T_55204[4]}},_T_55204}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_157 = {{6{_T_55211[4]}},_T_55211}; // @[Modules.scala 32:22:@8.4]
  assign _T_56608 = $signed(buffer_0_156) + $signed(buffer_0_157); // @[Modules.scala 50:57:@2588.4]
  assign _T_56609 = _T_56608[10:0]; // @[Modules.scala 50:57:@2589.4]
  assign buffer_0_470 = $signed(_T_56609); // @[Modules.scala 50:57:@2590.4]
  assign buffer_0_158 = {{6{_T_55214[4]}},_T_55214}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_159 = {{6{_T_55217[4]}},_T_55217}; // @[Modules.scala 32:22:@8.4]
  assign _T_56611 = $signed(buffer_0_158) + $signed(buffer_0_159); // @[Modules.scala 50:57:@2592.4]
  assign _T_56612 = _T_56611[10:0]; // @[Modules.scala 50:57:@2593.4]
  assign buffer_0_471 = $signed(_T_56612); // @[Modules.scala 50:57:@2594.4]
  assign buffer_0_160 = {{6{_T_55224[4]}},_T_55224}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_161 = {{6{_T_55231[4]}},_T_55231}; // @[Modules.scala 32:22:@8.4]
  assign _T_56614 = $signed(buffer_0_160) + $signed(buffer_0_161); // @[Modules.scala 50:57:@2596.4]
  assign _T_56615 = _T_56614[10:0]; // @[Modules.scala 50:57:@2597.4]
  assign buffer_0_472 = $signed(_T_56615); // @[Modules.scala 50:57:@2598.4]
  assign buffer_0_162 = {{6{_T_55238[4]}},_T_55238}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_163 = {{6{_T_55245[4]}},_T_55245}; // @[Modules.scala 32:22:@8.4]
  assign _T_56617 = $signed(buffer_0_162) + $signed(buffer_0_163); // @[Modules.scala 50:57:@2600.4]
  assign _T_56618 = _T_56617[10:0]; // @[Modules.scala 50:57:@2601.4]
  assign buffer_0_473 = $signed(_T_56618); // @[Modules.scala 50:57:@2602.4]
  assign buffer_0_164 = {{6{_T_55248[4]}},_T_55248}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_165 = {{6{_T_55255[4]}},_T_55255}; // @[Modules.scala 32:22:@8.4]
  assign _T_56620 = $signed(buffer_0_164) + $signed(buffer_0_165); // @[Modules.scala 50:57:@2604.4]
  assign _T_56621 = _T_56620[10:0]; // @[Modules.scala 50:57:@2605.4]
  assign buffer_0_474 = $signed(_T_56621); // @[Modules.scala 50:57:@2606.4]
  assign buffer_0_166 = {{6{_T_55262[4]}},_T_55262}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_167 = {{6{_T_55269[4]}},_T_55269}; // @[Modules.scala 32:22:@8.4]
  assign _T_56623 = $signed(buffer_0_166) + $signed(buffer_0_167); // @[Modules.scala 50:57:@2608.4]
  assign _T_56624 = _T_56623[10:0]; // @[Modules.scala 50:57:@2609.4]
  assign buffer_0_475 = $signed(_T_56624); // @[Modules.scala 50:57:@2610.4]
  assign buffer_0_168 = {{6{_T_55272[4]}},_T_55272}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_169 = {{6{_T_55279[4]}},_T_55279}; // @[Modules.scala 32:22:@8.4]
  assign _T_56626 = $signed(buffer_0_168) + $signed(buffer_0_169); // @[Modules.scala 50:57:@2612.4]
  assign _T_56627 = _T_56626[10:0]; // @[Modules.scala 50:57:@2613.4]
  assign buffer_0_476 = $signed(_T_56627); // @[Modules.scala 50:57:@2614.4]
  assign buffer_0_170 = {{6{_T_55286[4]}},_T_55286}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_171 = {{6{_T_55289[4]}},_T_55289}; // @[Modules.scala 32:22:@8.4]
  assign _T_56629 = $signed(buffer_0_170) + $signed(buffer_0_171); // @[Modules.scala 50:57:@2616.4]
  assign _T_56630 = _T_56629[10:0]; // @[Modules.scala 50:57:@2617.4]
  assign buffer_0_477 = $signed(_T_56630); // @[Modules.scala 50:57:@2618.4]
  assign buffer_0_172 = {{6{_T_55292[4]}},_T_55292}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_173 = {{6{_T_55295[4]}},_T_55295}; // @[Modules.scala 32:22:@8.4]
  assign _T_56632 = $signed(buffer_0_172) + $signed(buffer_0_173); // @[Modules.scala 50:57:@2620.4]
  assign _T_56633 = _T_56632[10:0]; // @[Modules.scala 50:57:@2621.4]
  assign buffer_0_478 = $signed(_T_56633); // @[Modules.scala 50:57:@2622.4]
  assign buffer_0_174 = {{6{_T_55298[4]}},_T_55298}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_175 = {{6{_T_55301[4]}},_T_55301}; // @[Modules.scala 32:22:@8.4]
  assign _T_56635 = $signed(buffer_0_174) + $signed(buffer_0_175); // @[Modules.scala 50:57:@2624.4]
  assign _T_56636 = _T_56635[10:0]; // @[Modules.scala 50:57:@2625.4]
  assign buffer_0_479 = $signed(_T_56636); // @[Modules.scala 50:57:@2626.4]
  assign buffer_0_176 = {{6{_T_55304[4]}},_T_55304}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_177 = {{6{_T_55307[4]}},_T_55307}; // @[Modules.scala 32:22:@8.4]
  assign _T_56638 = $signed(buffer_0_176) + $signed(buffer_0_177); // @[Modules.scala 50:57:@2628.4]
  assign _T_56639 = _T_56638[10:0]; // @[Modules.scala 50:57:@2629.4]
  assign buffer_0_480 = $signed(_T_56639); // @[Modules.scala 50:57:@2630.4]
  assign buffer_0_178 = {{6{_T_55310[4]}},_T_55310}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_179 = {{6{_T_55313[4]}},_T_55313}; // @[Modules.scala 32:22:@8.4]
  assign _T_56641 = $signed(buffer_0_178) + $signed(buffer_0_179); // @[Modules.scala 50:57:@2632.4]
  assign _T_56642 = _T_56641[10:0]; // @[Modules.scala 50:57:@2633.4]
  assign buffer_0_481 = $signed(_T_56642); // @[Modules.scala 50:57:@2634.4]
  assign buffer_0_180 = {{6{_T_55320[4]}},_T_55320}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_181 = {{6{_T_55327[4]}},_T_55327}; // @[Modules.scala 32:22:@8.4]
  assign _T_56644 = $signed(buffer_0_180) + $signed(buffer_0_181); // @[Modules.scala 50:57:@2636.4]
  assign _T_56645 = _T_56644[10:0]; // @[Modules.scala 50:57:@2637.4]
  assign buffer_0_482 = $signed(_T_56645); // @[Modules.scala 50:57:@2638.4]
  assign buffer_0_182 = {{6{_T_55334[4]}},_T_55334}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_183 = {{6{_T_55341[4]}},_T_55341}; // @[Modules.scala 32:22:@8.4]
  assign _T_56647 = $signed(buffer_0_182) + $signed(buffer_0_183); // @[Modules.scala 50:57:@2640.4]
  assign _T_56648 = _T_56647[10:0]; // @[Modules.scala 50:57:@2641.4]
  assign buffer_0_483 = $signed(_T_56648); // @[Modules.scala 50:57:@2642.4]
  assign buffer_0_184 = {{6{_T_55344[4]}},_T_55344}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_185 = {{6{_T_55347[4]}},_T_55347}; // @[Modules.scala 32:22:@8.4]
  assign _T_56650 = $signed(buffer_0_184) + $signed(buffer_0_185); // @[Modules.scala 50:57:@2644.4]
  assign _T_56651 = _T_56650[10:0]; // @[Modules.scala 50:57:@2645.4]
  assign buffer_0_484 = $signed(_T_56651); // @[Modules.scala 50:57:@2646.4]
  assign buffer_0_186 = {{6{_T_55350[4]}},_T_55350}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_187 = {{6{_T_55353[4]}},_T_55353}; // @[Modules.scala 32:22:@8.4]
  assign _T_56653 = $signed(buffer_0_186) + $signed(buffer_0_187); // @[Modules.scala 50:57:@2648.4]
  assign _T_56654 = _T_56653[10:0]; // @[Modules.scala 50:57:@2649.4]
  assign buffer_0_485 = $signed(_T_56654); // @[Modules.scala 50:57:@2650.4]
  assign buffer_0_188 = {{6{_T_55356[4]}},_T_55356}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_189 = {{6{_T_55359[4]}},_T_55359}; // @[Modules.scala 32:22:@8.4]
  assign _T_56656 = $signed(buffer_0_188) + $signed(buffer_0_189); // @[Modules.scala 50:57:@2652.4]
  assign _T_56657 = _T_56656[10:0]; // @[Modules.scala 50:57:@2653.4]
  assign buffer_0_486 = $signed(_T_56657); // @[Modules.scala 50:57:@2654.4]
  assign buffer_0_190 = {{6{_T_55362[4]}},_T_55362}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_191 = {{6{_T_55365[4]}},_T_55365}; // @[Modules.scala 32:22:@8.4]
  assign _T_56659 = $signed(buffer_0_190) + $signed(buffer_0_191); // @[Modules.scala 50:57:@2656.4]
  assign _T_56660 = _T_56659[10:0]; // @[Modules.scala 50:57:@2657.4]
  assign buffer_0_487 = $signed(_T_56660); // @[Modules.scala 50:57:@2658.4]
  assign buffer_0_192 = {{6{_T_55372[4]}},_T_55372}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_193 = {{6{_T_55375[4]}},_T_55375}; // @[Modules.scala 32:22:@8.4]
  assign _T_56662 = $signed(buffer_0_192) + $signed(buffer_0_193); // @[Modules.scala 50:57:@2660.4]
  assign _T_56663 = _T_56662[10:0]; // @[Modules.scala 50:57:@2661.4]
  assign buffer_0_488 = $signed(_T_56663); // @[Modules.scala 50:57:@2662.4]
  assign buffer_0_194 = {{6{_T_55378[4]}},_T_55378}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_195 = {{6{_T_55385[4]}},_T_55385}; // @[Modules.scala 32:22:@8.4]
  assign _T_56665 = $signed(buffer_0_194) + $signed(buffer_0_195); // @[Modules.scala 50:57:@2664.4]
  assign _T_56666 = _T_56665[10:0]; // @[Modules.scala 50:57:@2665.4]
  assign buffer_0_489 = $signed(_T_56666); // @[Modules.scala 50:57:@2666.4]
  assign buffer_0_196 = {{6{_T_55392[4]}},_T_55392}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_197 = {{6{_T_55399[4]}},_T_55399}; // @[Modules.scala 32:22:@8.4]
  assign _T_56668 = $signed(buffer_0_196) + $signed(buffer_0_197); // @[Modules.scala 50:57:@2668.4]
  assign _T_56669 = _T_56668[10:0]; // @[Modules.scala 50:57:@2669.4]
  assign buffer_0_490 = $signed(_T_56669); // @[Modules.scala 50:57:@2670.4]
  assign buffer_0_198 = {{6{_T_55402[4]}},_T_55402}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_199 = {{6{_T_55405[4]}},_T_55405}; // @[Modules.scala 32:22:@8.4]
  assign _T_56671 = $signed(buffer_0_198) + $signed(buffer_0_199); // @[Modules.scala 50:57:@2672.4]
  assign _T_56672 = _T_56671[10:0]; // @[Modules.scala 50:57:@2673.4]
  assign buffer_0_491 = $signed(_T_56672); // @[Modules.scala 50:57:@2674.4]
  assign buffer_0_200 = {{6{_T_55408[4]}},_T_55408}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_201 = {{6{_T_55411[4]}},_T_55411}; // @[Modules.scala 32:22:@8.4]
  assign _T_56674 = $signed(buffer_0_200) + $signed(buffer_0_201); // @[Modules.scala 50:57:@2676.4]
  assign _T_56675 = _T_56674[10:0]; // @[Modules.scala 50:57:@2677.4]
  assign buffer_0_492 = $signed(_T_56675); // @[Modules.scala 50:57:@2678.4]
  assign buffer_0_202 = {{6{_T_55414[4]}},_T_55414}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_203 = {{6{_T_55417[4]}},_T_55417}; // @[Modules.scala 32:22:@8.4]
  assign _T_56677 = $signed(buffer_0_202) + $signed(buffer_0_203); // @[Modules.scala 50:57:@2680.4]
  assign _T_56678 = _T_56677[10:0]; // @[Modules.scala 50:57:@2681.4]
  assign buffer_0_493 = $signed(_T_56678); // @[Modules.scala 50:57:@2682.4]
  assign buffer_0_204 = {{6{_T_55420[4]}},_T_55420}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_205 = {{6{_T_55423[4]}},_T_55423}; // @[Modules.scala 32:22:@8.4]
  assign _T_56680 = $signed(buffer_0_204) + $signed(buffer_0_205); // @[Modules.scala 50:57:@2684.4]
  assign _T_56681 = _T_56680[10:0]; // @[Modules.scala 50:57:@2685.4]
  assign buffer_0_494 = $signed(_T_56681); // @[Modules.scala 50:57:@2686.4]
  assign buffer_0_206 = {{6{_T_55426[4]}},_T_55426}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_207 = {{6{_T_55429[4]}},_T_55429}; // @[Modules.scala 32:22:@8.4]
  assign _T_56683 = $signed(buffer_0_206) + $signed(buffer_0_207); // @[Modules.scala 50:57:@2688.4]
  assign _T_56684 = _T_56683[10:0]; // @[Modules.scala 50:57:@2689.4]
  assign buffer_0_495 = $signed(_T_56684); // @[Modules.scala 50:57:@2690.4]
  assign buffer_0_208 = {{6{_T_55432[4]}},_T_55432}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_209 = {{6{_T_55439[4]}},_T_55439}; // @[Modules.scala 32:22:@8.4]
  assign _T_56686 = $signed(buffer_0_208) + $signed(buffer_0_209); // @[Modules.scala 50:57:@2692.4]
  assign _T_56687 = _T_56686[10:0]; // @[Modules.scala 50:57:@2693.4]
  assign buffer_0_496 = $signed(_T_56687); // @[Modules.scala 50:57:@2694.4]
  assign buffer_0_210 = {{6{_T_55446[4]}},_T_55446}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_211 = {{6{_T_55453[4]}},_T_55453}; // @[Modules.scala 32:22:@8.4]
  assign _T_56689 = $signed(buffer_0_210) + $signed(buffer_0_211); // @[Modules.scala 50:57:@2696.4]
  assign _T_56690 = _T_56689[10:0]; // @[Modules.scala 50:57:@2697.4]
  assign buffer_0_497 = $signed(_T_56690); // @[Modules.scala 50:57:@2698.4]
  assign buffer_0_212 = {{6{_T_55460[4]}},_T_55460}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_213 = {{6{_T_55463[4]}},_T_55463}; // @[Modules.scala 32:22:@8.4]
  assign _T_56692 = $signed(buffer_0_212) + $signed(buffer_0_213); // @[Modules.scala 50:57:@2700.4]
  assign _T_56693 = _T_56692[10:0]; // @[Modules.scala 50:57:@2701.4]
  assign buffer_0_498 = $signed(_T_56693); // @[Modules.scala 50:57:@2702.4]
  assign buffer_0_214 = {{6{_T_55466[4]}},_T_55466}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_215 = {{6{_T_55469[4]}},_T_55469}; // @[Modules.scala 32:22:@8.4]
  assign _T_56695 = $signed(buffer_0_214) + $signed(buffer_0_215); // @[Modules.scala 50:57:@2704.4]
  assign _T_56696 = _T_56695[10:0]; // @[Modules.scala 50:57:@2705.4]
  assign buffer_0_499 = $signed(_T_56696); // @[Modules.scala 50:57:@2706.4]
  assign buffer_0_216 = {{6{_T_55472[4]}},_T_55472}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_217 = {{6{_T_55475[4]}},_T_55475}; // @[Modules.scala 32:22:@8.4]
  assign _T_56698 = $signed(buffer_0_216) + $signed(buffer_0_217); // @[Modules.scala 50:57:@2708.4]
  assign _T_56699 = _T_56698[10:0]; // @[Modules.scala 50:57:@2709.4]
  assign buffer_0_500 = $signed(_T_56699); // @[Modules.scala 50:57:@2710.4]
  assign buffer_0_218 = {{6{_T_55478[4]}},_T_55478}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_219 = {{6{_T_55481[4]}},_T_55481}; // @[Modules.scala 32:22:@8.4]
  assign _T_56701 = $signed(buffer_0_218) + $signed(buffer_0_219); // @[Modules.scala 50:57:@2712.4]
  assign _T_56702 = _T_56701[10:0]; // @[Modules.scala 50:57:@2713.4]
  assign buffer_0_501 = $signed(_T_56702); // @[Modules.scala 50:57:@2714.4]
  assign buffer_0_220 = {{6{_T_55484[4]}},_T_55484}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_221 = {{6{_T_55491[4]}},_T_55491}; // @[Modules.scala 32:22:@8.4]
  assign _T_56704 = $signed(buffer_0_220) + $signed(buffer_0_221); // @[Modules.scala 50:57:@2716.4]
  assign _T_56705 = _T_56704[10:0]; // @[Modules.scala 50:57:@2717.4]
  assign buffer_0_502 = $signed(_T_56705); // @[Modules.scala 50:57:@2718.4]
  assign buffer_0_222 = {{6{_T_55498[4]}},_T_55498}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_223 = {{6{_T_55505[4]}},_T_55505}; // @[Modules.scala 32:22:@8.4]
  assign _T_56707 = $signed(buffer_0_222) + $signed(buffer_0_223); // @[Modules.scala 50:57:@2720.4]
  assign _T_56708 = _T_56707[10:0]; // @[Modules.scala 50:57:@2721.4]
  assign buffer_0_503 = $signed(_T_56708); // @[Modules.scala 50:57:@2722.4]
  assign buffer_0_224 = {{6{_T_55508[4]}},_T_55508}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_225 = {{6{_T_55515[4]}},_T_55515}; // @[Modules.scala 32:22:@8.4]
  assign _T_56710 = $signed(buffer_0_224) + $signed(buffer_0_225); // @[Modules.scala 50:57:@2724.4]
  assign _T_56711 = _T_56710[10:0]; // @[Modules.scala 50:57:@2725.4]
  assign buffer_0_504 = $signed(_T_56711); // @[Modules.scala 50:57:@2726.4]
  assign buffer_0_226 = {{6{_T_55522[4]}},_T_55522}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_227 = {{6{_T_55525[4]}},_T_55525}; // @[Modules.scala 32:22:@8.4]
  assign _T_56713 = $signed(buffer_0_226) + $signed(buffer_0_227); // @[Modules.scala 50:57:@2728.4]
  assign _T_56714 = _T_56713[10:0]; // @[Modules.scala 50:57:@2729.4]
  assign buffer_0_505 = $signed(_T_56714); // @[Modules.scala 50:57:@2730.4]
  assign buffer_0_228 = {{6{_T_55528[4]}},_T_55528}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_229 = {{6{_T_55531[4]}},_T_55531}; // @[Modules.scala 32:22:@8.4]
  assign _T_56716 = $signed(buffer_0_228) + $signed(buffer_0_229); // @[Modules.scala 50:57:@2732.4]
  assign _T_56717 = _T_56716[10:0]; // @[Modules.scala 50:57:@2733.4]
  assign buffer_0_506 = $signed(_T_56717); // @[Modules.scala 50:57:@2734.4]
  assign buffer_0_230 = {{6{_T_55534[4]}},_T_55534}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_231 = {{6{_T_55537[4]}},_T_55537}; // @[Modules.scala 32:22:@8.4]
  assign _T_56719 = $signed(buffer_0_230) + $signed(buffer_0_231); // @[Modules.scala 50:57:@2736.4]
  assign _T_56720 = _T_56719[10:0]; // @[Modules.scala 50:57:@2737.4]
  assign buffer_0_507 = $signed(_T_56720); // @[Modules.scala 50:57:@2738.4]
  assign buffer_0_232 = {{6{_T_55540[4]}},_T_55540}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_233 = {{6{_T_55543[4]}},_T_55543}; // @[Modules.scala 32:22:@8.4]
  assign _T_56722 = $signed(buffer_0_232) + $signed(buffer_0_233); // @[Modules.scala 50:57:@2740.4]
  assign _T_56723 = _T_56722[10:0]; // @[Modules.scala 50:57:@2741.4]
  assign buffer_0_508 = $signed(_T_56723); // @[Modules.scala 50:57:@2742.4]
  assign buffer_0_234 = {{6{_T_55546[4]}},_T_55546}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_235 = {{6{_T_55553[4]}},_T_55553}; // @[Modules.scala 32:22:@8.4]
  assign _T_56725 = $signed(buffer_0_234) + $signed(buffer_0_235); // @[Modules.scala 50:57:@2744.4]
  assign _T_56726 = _T_56725[10:0]; // @[Modules.scala 50:57:@2745.4]
  assign buffer_0_509 = $signed(_T_56726); // @[Modules.scala 50:57:@2746.4]
  assign buffer_0_236 = {{6{_T_55560[4]}},_T_55560}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_237 = {{6{_T_55567[4]}},_T_55567}; // @[Modules.scala 32:22:@8.4]
  assign _T_56728 = $signed(buffer_0_236) + $signed(buffer_0_237); // @[Modules.scala 50:57:@2748.4]
  assign _T_56729 = _T_56728[10:0]; // @[Modules.scala 50:57:@2749.4]
  assign buffer_0_510 = $signed(_T_56729); // @[Modules.scala 50:57:@2750.4]
  assign buffer_0_238 = {{6{_T_55574[4]}},_T_55574}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_239 = {{6{_T_55577[4]}},_T_55577}; // @[Modules.scala 32:22:@8.4]
  assign _T_56731 = $signed(buffer_0_238) + $signed(buffer_0_239); // @[Modules.scala 50:57:@2752.4]
  assign _T_56732 = _T_56731[10:0]; // @[Modules.scala 50:57:@2753.4]
  assign buffer_0_511 = $signed(_T_56732); // @[Modules.scala 50:57:@2754.4]
  assign buffer_0_240 = {{6{_T_55584[4]}},_T_55584}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_241 = {{6{_T_55587[4]}},_T_55587}; // @[Modules.scala 32:22:@8.4]
  assign _T_56734 = $signed(buffer_0_240) + $signed(buffer_0_241); // @[Modules.scala 50:57:@2756.4]
  assign _T_56735 = _T_56734[10:0]; // @[Modules.scala 50:57:@2757.4]
  assign buffer_0_512 = $signed(_T_56735); // @[Modules.scala 50:57:@2758.4]
  assign buffer_0_242 = {{6{_T_55590[4]}},_T_55590}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_243 = {{6{_T_55593[4]}},_T_55593}; // @[Modules.scala 32:22:@8.4]
  assign _T_56737 = $signed(buffer_0_242) + $signed(buffer_0_243); // @[Modules.scala 50:57:@2760.4]
  assign _T_56738 = _T_56737[10:0]; // @[Modules.scala 50:57:@2761.4]
  assign buffer_0_513 = $signed(_T_56738); // @[Modules.scala 50:57:@2762.4]
  assign buffer_0_244 = {{6{_T_55600[4]}},_T_55600}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_245 = {{6{_T_55603[4]}},_T_55603}; // @[Modules.scala 32:22:@8.4]
  assign _T_56740 = $signed(buffer_0_244) + $signed(buffer_0_245); // @[Modules.scala 50:57:@2764.4]
  assign _T_56741 = _T_56740[10:0]; // @[Modules.scala 50:57:@2765.4]
  assign buffer_0_514 = $signed(_T_56741); // @[Modules.scala 50:57:@2766.4]
  assign buffer_0_246 = {{6{_T_55606[4]}},_T_55606}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_247 = {{6{_T_55609[4]}},_T_55609}; // @[Modules.scala 32:22:@8.4]
  assign _T_56743 = $signed(buffer_0_246) + $signed(buffer_0_247); // @[Modules.scala 50:57:@2768.4]
  assign _T_56744 = _T_56743[10:0]; // @[Modules.scala 50:57:@2769.4]
  assign buffer_0_515 = $signed(_T_56744); // @[Modules.scala 50:57:@2770.4]
  assign buffer_0_248 = {{6{_T_55616[4]}},_T_55616}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_249 = {{6{_T_55619[4]}},_T_55619}; // @[Modules.scala 32:22:@8.4]
  assign _T_56746 = $signed(buffer_0_248) + $signed(buffer_0_249); // @[Modules.scala 50:57:@2772.4]
  assign _T_56747 = _T_56746[10:0]; // @[Modules.scala 50:57:@2773.4]
  assign buffer_0_516 = $signed(_T_56747); // @[Modules.scala 50:57:@2774.4]
  assign buffer_0_250 = {{6{_T_55626[4]}},_T_55626}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_251 = {{6{_T_55633[4]}},_T_55633}; // @[Modules.scala 32:22:@8.4]
  assign _T_56749 = $signed(buffer_0_250) + $signed(buffer_0_251); // @[Modules.scala 50:57:@2776.4]
  assign _T_56750 = _T_56749[10:0]; // @[Modules.scala 50:57:@2777.4]
  assign buffer_0_517 = $signed(_T_56750); // @[Modules.scala 50:57:@2778.4]
  assign buffer_0_252 = {{6{_T_55640[4]}},_T_55640}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_253 = {{6{_T_55647[4]}},_T_55647}; // @[Modules.scala 32:22:@8.4]
  assign _T_56752 = $signed(buffer_0_252) + $signed(buffer_0_253); // @[Modules.scala 50:57:@2780.4]
  assign _T_56753 = _T_56752[10:0]; // @[Modules.scala 50:57:@2781.4]
  assign buffer_0_518 = $signed(_T_56753); // @[Modules.scala 50:57:@2782.4]
  assign buffer_0_254 = {{6{_T_55654[4]}},_T_55654}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_255 = {{6{_T_55661[4]}},_T_55661}; // @[Modules.scala 32:22:@8.4]
  assign _T_56755 = $signed(buffer_0_254) + $signed(buffer_0_255); // @[Modules.scala 50:57:@2784.4]
  assign _T_56756 = _T_56755[10:0]; // @[Modules.scala 50:57:@2785.4]
  assign buffer_0_519 = $signed(_T_56756); // @[Modules.scala 50:57:@2786.4]
  assign buffer_0_256 = {{6{_T_55664[4]}},_T_55664}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_257 = {{6{_T_55667[4]}},_T_55667}; // @[Modules.scala 32:22:@8.4]
  assign _T_56758 = $signed(buffer_0_256) + $signed(buffer_0_257); // @[Modules.scala 50:57:@2788.4]
  assign _T_56759 = _T_56758[10:0]; // @[Modules.scala 50:57:@2789.4]
  assign buffer_0_520 = $signed(_T_56759); // @[Modules.scala 50:57:@2790.4]
  assign buffer_0_258 = {{6{_T_55670[4]}},_T_55670}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_259 = {{6{_T_55673[4]}},_T_55673}; // @[Modules.scala 32:22:@8.4]
  assign _T_56761 = $signed(buffer_0_258) + $signed(buffer_0_259); // @[Modules.scala 50:57:@2792.4]
  assign _T_56762 = _T_56761[10:0]; // @[Modules.scala 50:57:@2793.4]
  assign buffer_0_521 = $signed(_T_56762); // @[Modules.scala 50:57:@2794.4]
  assign buffer_0_260 = {{6{_T_55680[4]}},_T_55680}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_261 = {{6{_T_55687[4]}},_T_55687}; // @[Modules.scala 32:22:@8.4]
  assign _T_56764 = $signed(buffer_0_260) + $signed(buffer_0_261); // @[Modules.scala 50:57:@2796.4]
  assign _T_56765 = _T_56764[10:0]; // @[Modules.scala 50:57:@2797.4]
  assign buffer_0_522 = $signed(_T_56765); // @[Modules.scala 50:57:@2798.4]
  assign buffer_0_262 = {{6{_T_55694[4]}},_T_55694}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_263 = {{6{_T_55697[4]}},_T_55697}; // @[Modules.scala 32:22:@8.4]
  assign _T_56767 = $signed(buffer_0_262) + $signed(buffer_0_263); // @[Modules.scala 50:57:@2800.4]
  assign _T_56768 = _T_56767[10:0]; // @[Modules.scala 50:57:@2801.4]
  assign buffer_0_523 = $signed(_T_56768); // @[Modules.scala 50:57:@2802.4]
  assign buffer_0_264 = {{6{_T_55700[4]}},_T_55700}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_265 = {{6{_T_55707[4]}},_T_55707}; // @[Modules.scala 32:22:@8.4]
  assign _T_56770 = $signed(buffer_0_264) + $signed(buffer_0_265); // @[Modules.scala 50:57:@2804.4]
  assign _T_56771 = _T_56770[10:0]; // @[Modules.scala 50:57:@2805.4]
  assign buffer_0_524 = $signed(_T_56771); // @[Modules.scala 50:57:@2806.4]
  assign buffer_0_266 = {{6{_T_55710[4]}},_T_55710}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_267 = {{6{_T_55717[4]}},_T_55717}; // @[Modules.scala 32:22:@8.4]
  assign _T_56773 = $signed(buffer_0_266) + $signed(buffer_0_267); // @[Modules.scala 50:57:@2808.4]
  assign _T_56774 = _T_56773[10:0]; // @[Modules.scala 50:57:@2809.4]
  assign buffer_0_525 = $signed(_T_56774); // @[Modules.scala 50:57:@2810.4]
  assign buffer_0_268 = {{6{_T_55724[4]}},_T_55724}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_269 = {{6{_T_55731[4]}},_T_55731}; // @[Modules.scala 32:22:@8.4]
  assign _T_56776 = $signed(buffer_0_268) + $signed(buffer_0_269); // @[Modules.scala 50:57:@2812.4]
  assign _T_56777 = _T_56776[10:0]; // @[Modules.scala 50:57:@2813.4]
  assign buffer_0_526 = $signed(_T_56777); // @[Modules.scala 50:57:@2814.4]
  assign buffer_0_270 = {{6{_T_55738[4]}},_T_55738}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_271 = {{6{_T_55745[4]}},_T_55745}; // @[Modules.scala 32:22:@8.4]
  assign _T_56779 = $signed(buffer_0_270) + $signed(buffer_0_271); // @[Modules.scala 50:57:@2816.4]
  assign _T_56780 = _T_56779[10:0]; // @[Modules.scala 50:57:@2817.4]
  assign buffer_0_527 = $signed(_T_56780); // @[Modules.scala 50:57:@2818.4]
  assign buffer_0_272 = {{6{_T_55752[4]}},_T_55752}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_273 = {{6{_T_55759[4]}},_T_55759}; // @[Modules.scala 32:22:@8.4]
  assign _T_56782 = $signed(buffer_0_272) + $signed(buffer_0_273); // @[Modules.scala 50:57:@2820.4]
  assign _T_56783 = _T_56782[10:0]; // @[Modules.scala 50:57:@2821.4]
  assign buffer_0_528 = $signed(_T_56783); // @[Modules.scala 50:57:@2822.4]
  assign buffer_0_274 = {{6{_T_55766[4]}},_T_55766}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_275 = {{6{_T_55769[4]}},_T_55769}; // @[Modules.scala 32:22:@8.4]
  assign _T_56785 = $signed(buffer_0_274) + $signed(buffer_0_275); // @[Modules.scala 50:57:@2824.4]
  assign _T_56786 = _T_56785[10:0]; // @[Modules.scala 50:57:@2825.4]
  assign buffer_0_529 = $signed(_T_56786); // @[Modules.scala 50:57:@2826.4]
  assign buffer_0_276 = {{6{_T_55772[4]}},_T_55772}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_277 = {{6{_T_55779[4]}},_T_55779}; // @[Modules.scala 32:22:@8.4]
  assign _T_56788 = $signed(buffer_0_276) + $signed(buffer_0_277); // @[Modules.scala 50:57:@2828.4]
  assign _T_56789 = _T_56788[10:0]; // @[Modules.scala 50:57:@2829.4]
  assign buffer_0_530 = $signed(_T_56789); // @[Modules.scala 50:57:@2830.4]
  assign buffer_0_278 = {{6{_T_55782[4]}},_T_55782}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_279 = {{6{_T_55789[4]}},_T_55789}; // @[Modules.scala 32:22:@8.4]
  assign _T_56791 = $signed(buffer_0_278) + $signed(buffer_0_279); // @[Modules.scala 50:57:@2832.4]
  assign _T_56792 = _T_56791[10:0]; // @[Modules.scala 50:57:@2833.4]
  assign buffer_0_531 = $signed(_T_56792); // @[Modules.scala 50:57:@2834.4]
  assign buffer_0_280 = {{6{_T_55796[4]}},_T_55796}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_281 = {{6{_T_55803[4]}},_T_55803}; // @[Modules.scala 32:22:@8.4]
  assign _T_56794 = $signed(buffer_0_280) + $signed(buffer_0_281); // @[Modules.scala 50:57:@2836.4]
  assign _T_56795 = _T_56794[10:0]; // @[Modules.scala 50:57:@2837.4]
  assign buffer_0_532 = $signed(_T_56795); // @[Modules.scala 50:57:@2838.4]
  assign buffer_0_282 = {{6{_T_55810[4]}},_T_55810}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_283 = {{6{_T_55817[4]}},_T_55817}; // @[Modules.scala 32:22:@8.4]
  assign _T_56797 = $signed(buffer_0_282) + $signed(buffer_0_283); // @[Modules.scala 50:57:@2840.4]
  assign _T_56798 = _T_56797[10:0]; // @[Modules.scala 50:57:@2841.4]
  assign buffer_0_533 = $signed(_T_56798); // @[Modules.scala 50:57:@2842.4]
  assign buffer_0_284 = {{6{_T_55824[4]}},_T_55824}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_285 = {{6{_T_55831[4]}},_T_55831}; // @[Modules.scala 32:22:@8.4]
  assign _T_56800 = $signed(buffer_0_284) + $signed(buffer_0_285); // @[Modules.scala 50:57:@2844.4]
  assign _T_56801 = _T_56800[10:0]; // @[Modules.scala 50:57:@2845.4]
  assign buffer_0_534 = $signed(_T_56801); // @[Modules.scala 50:57:@2846.4]
  assign buffer_0_286 = {{6{_T_55838[4]}},_T_55838}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_287 = {{6{_T_55845[4]}},_T_55845}; // @[Modules.scala 32:22:@8.4]
  assign _T_56803 = $signed(buffer_0_286) + $signed(buffer_0_287); // @[Modules.scala 50:57:@2848.4]
  assign _T_56804 = _T_56803[10:0]; // @[Modules.scala 50:57:@2849.4]
  assign buffer_0_535 = $signed(_T_56804); // @[Modules.scala 50:57:@2850.4]
  assign buffer_0_288 = {{6{_T_55848[4]}},_T_55848}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_289 = {{6{_T_55851[4]}},_T_55851}; // @[Modules.scala 32:22:@8.4]
  assign _T_56806 = $signed(buffer_0_288) + $signed(buffer_0_289); // @[Modules.scala 50:57:@2852.4]
  assign _T_56807 = _T_56806[10:0]; // @[Modules.scala 50:57:@2853.4]
  assign buffer_0_536 = $signed(_T_56807); // @[Modules.scala 50:57:@2854.4]
  assign buffer_0_290 = {{6{_T_55854[4]}},_T_55854}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_291 = {{6{_T_55861[4]}},_T_55861}; // @[Modules.scala 32:22:@8.4]
  assign _T_56809 = $signed(buffer_0_290) + $signed(buffer_0_291); // @[Modules.scala 50:57:@2856.4]
  assign _T_56810 = _T_56809[10:0]; // @[Modules.scala 50:57:@2857.4]
  assign buffer_0_537 = $signed(_T_56810); // @[Modules.scala 50:57:@2858.4]
  assign buffer_0_292 = {{6{_T_55864[4]}},_T_55864}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_293 = {{6{_T_55871[4]}},_T_55871}; // @[Modules.scala 32:22:@8.4]
  assign _T_56812 = $signed(buffer_0_292) + $signed(buffer_0_293); // @[Modules.scala 50:57:@2860.4]
  assign _T_56813 = _T_56812[10:0]; // @[Modules.scala 50:57:@2861.4]
  assign buffer_0_538 = $signed(_T_56813); // @[Modules.scala 50:57:@2862.4]
  assign buffer_0_294 = {{6{_T_55878[4]}},_T_55878}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_295 = {{6{_T_55885[4]}},_T_55885}; // @[Modules.scala 32:22:@8.4]
  assign _T_56815 = $signed(buffer_0_294) + $signed(buffer_0_295); // @[Modules.scala 50:57:@2864.4]
  assign _T_56816 = _T_56815[10:0]; // @[Modules.scala 50:57:@2865.4]
  assign buffer_0_539 = $signed(_T_56816); // @[Modules.scala 50:57:@2866.4]
  assign buffer_0_296 = {{6{_T_55892[4]}},_T_55892}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_297 = {{6{_T_55899[4]}},_T_55899}; // @[Modules.scala 32:22:@8.4]
  assign _T_56818 = $signed(buffer_0_296) + $signed(buffer_0_297); // @[Modules.scala 50:57:@2868.4]
  assign _T_56819 = _T_56818[10:0]; // @[Modules.scala 50:57:@2869.4]
  assign buffer_0_540 = $signed(_T_56819); // @[Modules.scala 50:57:@2870.4]
  assign buffer_0_298 = {{6{_T_55906[4]}},_T_55906}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_299 = {{6{_T_55913[4]}},_T_55913}; // @[Modules.scala 32:22:@8.4]
  assign _T_56821 = $signed(buffer_0_298) + $signed(buffer_0_299); // @[Modules.scala 50:57:@2872.4]
  assign _T_56822 = _T_56821[10:0]; // @[Modules.scala 50:57:@2873.4]
  assign buffer_0_541 = $signed(_T_56822); // @[Modules.scala 50:57:@2874.4]
  assign buffer_0_300 = {{6{_T_55916[4]}},_T_55916}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_301 = {{6{_T_55919[4]}},_T_55919}; // @[Modules.scala 32:22:@8.4]
  assign _T_56824 = $signed(buffer_0_300) + $signed(buffer_0_301); // @[Modules.scala 50:57:@2876.4]
  assign _T_56825 = _T_56824[10:0]; // @[Modules.scala 50:57:@2877.4]
  assign buffer_0_542 = $signed(_T_56825); // @[Modules.scala 50:57:@2878.4]
  assign buffer_0_302 = {{6{_T_55922[4]}},_T_55922}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_303 = {{6{_T_55925[4]}},_T_55925}; // @[Modules.scala 32:22:@8.4]
  assign _T_56827 = $signed(buffer_0_302) + $signed(buffer_0_303); // @[Modules.scala 50:57:@2880.4]
  assign _T_56828 = _T_56827[10:0]; // @[Modules.scala 50:57:@2881.4]
  assign buffer_0_543 = $signed(_T_56828); // @[Modules.scala 50:57:@2882.4]
  assign buffer_0_304 = {{6{_T_55932[4]}},_T_55932}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_305 = {{6{_T_55939[4]}},_T_55939}; // @[Modules.scala 32:22:@8.4]
  assign _T_56830 = $signed(buffer_0_304) + $signed(buffer_0_305); // @[Modules.scala 50:57:@2884.4]
  assign _T_56831 = _T_56830[10:0]; // @[Modules.scala 50:57:@2885.4]
  assign buffer_0_544 = $signed(_T_56831); // @[Modules.scala 50:57:@2886.4]
  assign buffer_0_306 = {{6{_T_55942[4]}},_T_55942}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_307 = {{6{_T_55949[4]}},_T_55949}; // @[Modules.scala 32:22:@8.4]
  assign _T_56833 = $signed(buffer_0_306) + $signed(buffer_0_307); // @[Modules.scala 50:57:@2888.4]
  assign _T_56834 = _T_56833[10:0]; // @[Modules.scala 50:57:@2889.4]
  assign buffer_0_545 = $signed(_T_56834); // @[Modules.scala 50:57:@2890.4]
  assign buffer_0_308 = {{6{_T_55956[4]}},_T_55956}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_309 = {{6{_T_55959[4]}},_T_55959}; // @[Modules.scala 32:22:@8.4]
  assign _T_56836 = $signed(buffer_0_308) + $signed(buffer_0_309); // @[Modules.scala 50:57:@2892.4]
  assign _T_56837 = _T_56836[10:0]; // @[Modules.scala 50:57:@2893.4]
  assign buffer_0_546 = $signed(_T_56837); // @[Modules.scala 50:57:@2894.4]
  assign buffer_0_310 = {{6{_T_55966[4]}},_T_55966}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_311 = {{6{_T_55973[4]}},_T_55973}; // @[Modules.scala 32:22:@8.4]
  assign _T_56839 = $signed(buffer_0_310) + $signed(buffer_0_311); // @[Modules.scala 50:57:@2896.4]
  assign _T_56840 = _T_56839[10:0]; // @[Modules.scala 50:57:@2897.4]
  assign buffer_0_547 = $signed(_T_56840); // @[Modules.scala 50:57:@2898.4]
  assign buffer_0_312 = {{6{_T_55980[4]}},_T_55980}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_313 = {{6{_T_55987[4]}},_T_55987}; // @[Modules.scala 32:22:@8.4]
  assign _T_56842 = $signed(buffer_0_312) + $signed(buffer_0_313); // @[Modules.scala 50:57:@2900.4]
  assign _T_56843 = _T_56842[10:0]; // @[Modules.scala 50:57:@2901.4]
  assign buffer_0_548 = $signed(_T_56843); // @[Modules.scala 50:57:@2902.4]
  assign buffer_0_314 = {{6{_T_55994[4]}},_T_55994}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_315 = {{6{_T_56001[4]}},_T_56001}; // @[Modules.scala 32:22:@8.4]
  assign _T_56845 = $signed(buffer_0_314) + $signed(buffer_0_315); // @[Modules.scala 50:57:@2904.4]
  assign _T_56846 = _T_56845[10:0]; // @[Modules.scala 50:57:@2905.4]
  assign buffer_0_549 = $signed(_T_56846); // @[Modules.scala 50:57:@2906.4]
  assign buffer_0_316 = {{6{_T_56008[4]}},_T_56008}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_317 = {{6{_T_56015[4]}},_T_56015}; // @[Modules.scala 32:22:@8.4]
  assign _T_56848 = $signed(buffer_0_316) + $signed(buffer_0_317); // @[Modules.scala 50:57:@2908.4]
  assign _T_56849 = _T_56848[10:0]; // @[Modules.scala 50:57:@2909.4]
  assign buffer_0_550 = $signed(_T_56849); // @[Modules.scala 50:57:@2910.4]
  assign buffer_0_318 = {{6{_T_56022[4]}},_T_56022}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_319 = {{6{_T_56029[4]}},_T_56029}; // @[Modules.scala 32:22:@8.4]
  assign _T_56851 = $signed(buffer_0_318) + $signed(buffer_0_319); // @[Modules.scala 50:57:@2912.4]
  assign _T_56852 = _T_56851[10:0]; // @[Modules.scala 50:57:@2913.4]
  assign buffer_0_551 = $signed(_T_56852); // @[Modules.scala 50:57:@2914.4]
  assign buffer_0_320 = {{6{_T_56032[4]}},_T_56032}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_321 = {{6{_T_56039[4]}},_T_56039}; // @[Modules.scala 32:22:@8.4]
  assign _T_56854 = $signed(buffer_0_320) + $signed(buffer_0_321); // @[Modules.scala 50:57:@2916.4]
  assign _T_56855 = _T_56854[10:0]; // @[Modules.scala 50:57:@2917.4]
  assign buffer_0_552 = $signed(_T_56855); // @[Modules.scala 50:57:@2918.4]
  assign buffer_0_322 = {{6{_T_56046[4]}},_T_56046}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_323 = {{6{_T_56049[4]}},_T_56049}; // @[Modules.scala 32:22:@8.4]
  assign _T_56857 = $signed(buffer_0_322) + $signed(buffer_0_323); // @[Modules.scala 50:57:@2920.4]
  assign _T_56858 = _T_56857[10:0]; // @[Modules.scala 50:57:@2921.4]
  assign buffer_0_553 = $signed(_T_56858); // @[Modules.scala 50:57:@2922.4]
  assign buffer_0_324 = {{6{_T_56056[4]}},_T_56056}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_325 = {{6{_T_56063[4]}},_T_56063}; // @[Modules.scala 32:22:@8.4]
  assign _T_56860 = $signed(buffer_0_324) + $signed(buffer_0_325); // @[Modules.scala 50:57:@2924.4]
  assign _T_56861 = _T_56860[10:0]; // @[Modules.scala 50:57:@2925.4]
  assign buffer_0_554 = $signed(_T_56861); // @[Modules.scala 50:57:@2926.4]
  assign buffer_0_326 = {{6{_T_56070[4]}},_T_56070}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_327 = {{6{_T_56077[4]}},_T_56077}; // @[Modules.scala 32:22:@8.4]
  assign _T_56863 = $signed(buffer_0_326) + $signed(buffer_0_327); // @[Modules.scala 50:57:@2928.4]
  assign _T_56864 = _T_56863[10:0]; // @[Modules.scala 50:57:@2929.4]
  assign buffer_0_555 = $signed(_T_56864); // @[Modules.scala 50:57:@2930.4]
  assign buffer_0_328 = {{6{_T_56084[4]}},_T_56084}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_329 = {{6{_T_56091[4]}},_T_56091}; // @[Modules.scala 32:22:@8.4]
  assign _T_56866 = $signed(buffer_0_328) + $signed(buffer_0_329); // @[Modules.scala 50:57:@2932.4]
  assign _T_56867 = _T_56866[10:0]; // @[Modules.scala 50:57:@2933.4]
  assign buffer_0_556 = $signed(_T_56867); // @[Modules.scala 50:57:@2934.4]
  assign buffer_0_330 = {{6{_T_56098[4]}},_T_56098}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_331 = {{6{_T_56105[4]}},_T_56105}; // @[Modules.scala 32:22:@8.4]
  assign _T_56869 = $signed(buffer_0_330) + $signed(buffer_0_331); // @[Modules.scala 50:57:@2936.4]
  assign _T_56870 = _T_56869[10:0]; // @[Modules.scala 50:57:@2937.4]
  assign buffer_0_557 = $signed(_T_56870); // @[Modules.scala 50:57:@2938.4]
  assign buffer_0_332 = {{6{_T_56108[4]}},_T_56108}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_333 = {{6{_T_56111[4]}},_T_56111}; // @[Modules.scala 32:22:@8.4]
  assign _T_56872 = $signed(buffer_0_332) + $signed(buffer_0_333); // @[Modules.scala 50:57:@2940.4]
  assign _T_56873 = _T_56872[10:0]; // @[Modules.scala 50:57:@2941.4]
  assign buffer_0_558 = $signed(_T_56873); // @[Modules.scala 50:57:@2942.4]
  assign buffer_0_334 = {{6{_T_56114[4]}},_T_56114}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_335 = {{6{_T_56121[4]}},_T_56121}; // @[Modules.scala 32:22:@8.4]
  assign _T_56875 = $signed(buffer_0_334) + $signed(buffer_0_335); // @[Modules.scala 50:57:@2944.4]
  assign _T_56876 = _T_56875[10:0]; // @[Modules.scala 50:57:@2945.4]
  assign buffer_0_559 = $signed(_T_56876); // @[Modules.scala 50:57:@2946.4]
  assign buffer_0_336 = {{6{_T_56128[4]}},_T_56128}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_337 = {{6{_T_56131[4]}},_T_56131}; // @[Modules.scala 32:22:@8.4]
  assign _T_56878 = $signed(buffer_0_336) + $signed(buffer_0_337); // @[Modules.scala 50:57:@2948.4]
  assign _T_56879 = _T_56878[10:0]; // @[Modules.scala 50:57:@2949.4]
  assign buffer_0_560 = $signed(_T_56879); // @[Modules.scala 50:57:@2950.4]
  assign buffer_0_338 = {{6{_T_56134[4]}},_T_56134}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_339 = {{6{_T_56137[4]}},_T_56137}; // @[Modules.scala 32:22:@8.4]
  assign _T_56881 = $signed(buffer_0_338) + $signed(buffer_0_339); // @[Modules.scala 50:57:@2952.4]
  assign _T_56882 = _T_56881[10:0]; // @[Modules.scala 50:57:@2953.4]
  assign buffer_0_561 = $signed(_T_56882); // @[Modules.scala 50:57:@2954.4]
  assign buffer_0_340 = {{6{_T_56140[4]}},_T_56140}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_341 = {{6{_T_56143[4]}},_T_56143}; // @[Modules.scala 32:22:@8.4]
  assign _T_56884 = $signed(buffer_0_340) + $signed(buffer_0_341); // @[Modules.scala 50:57:@2956.4]
  assign _T_56885 = _T_56884[10:0]; // @[Modules.scala 50:57:@2957.4]
  assign buffer_0_562 = $signed(_T_56885); // @[Modules.scala 50:57:@2958.4]
  assign buffer_0_342 = {{6{_T_56150[4]}},_T_56150}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_343 = {{6{_T_56157[4]}},_T_56157}; // @[Modules.scala 32:22:@8.4]
  assign _T_56887 = $signed(buffer_0_342) + $signed(buffer_0_343); // @[Modules.scala 50:57:@2960.4]
  assign _T_56888 = _T_56887[10:0]; // @[Modules.scala 50:57:@2961.4]
  assign buffer_0_563 = $signed(_T_56888); // @[Modules.scala 50:57:@2962.4]
  assign buffer_0_344 = {{6{_T_56160[4]}},_T_56160}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_345 = {{6{_T_56163[4]}},_T_56163}; // @[Modules.scala 32:22:@8.4]
  assign _T_56890 = $signed(buffer_0_344) + $signed(buffer_0_345); // @[Modules.scala 50:57:@2964.4]
  assign _T_56891 = _T_56890[10:0]; // @[Modules.scala 50:57:@2965.4]
  assign buffer_0_564 = $signed(_T_56891); // @[Modules.scala 50:57:@2966.4]
  assign buffer_0_346 = {{6{_T_56166[4]}},_T_56166}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_347 = {{6{_T_56169[4]}},_T_56169}; // @[Modules.scala 32:22:@8.4]
  assign _T_56893 = $signed(buffer_0_346) + $signed(buffer_0_347); // @[Modules.scala 50:57:@2968.4]
  assign _T_56894 = _T_56893[10:0]; // @[Modules.scala 50:57:@2969.4]
  assign buffer_0_565 = $signed(_T_56894); // @[Modules.scala 50:57:@2970.4]
  assign buffer_0_348 = {{6{_T_56172[4]}},_T_56172}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_349 = {{6{_T_56179[4]}},_T_56179}; // @[Modules.scala 32:22:@8.4]
  assign _T_56896 = $signed(buffer_0_348) + $signed(buffer_0_349); // @[Modules.scala 50:57:@2972.4]
  assign _T_56897 = _T_56896[10:0]; // @[Modules.scala 50:57:@2973.4]
  assign buffer_0_566 = $signed(_T_56897); // @[Modules.scala 50:57:@2974.4]
  assign buffer_0_350 = {{6{_T_56186[4]}},_T_56186}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_351 = {{6{_T_56189[4]}},_T_56189}; // @[Modules.scala 32:22:@8.4]
  assign _T_56899 = $signed(buffer_0_350) + $signed(buffer_0_351); // @[Modules.scala 50:57:@2976.4]
  assign _T_56900 = _T_56899[10:0]; // @[Modules.scala 50:57:@2977.4]
  assign buffer_0_567 = $signed(_T_56900); // @[Modules.scala 50:57:@2978.4]
  assign buffer_0_352 = {{6{_T_56192[4]}},_T_56192}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_353 = {{6{_T_56195[4]}},_T_56195}; // @[Modules.scala 32:22:@8.4]
  assign _T_56902 = $signed(buffer_0_352) + $signed(buffer_0_353); // @[Modules.scala 50:57:@2980.4]
  assign _T_56903 = _T_56902[10:0]; // @[Modules.scala 50:57:@2981.4]
  assign buffer_0_568 = $signed(_T_56903); // @[Modules.scala 50:57:@2982.4]
  assign buffer_0_354 = {{6{_T_56198[4]}},_T_56198}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_355 = {{6{_T_56201[4]}},_T_56201}; // @[Modules.scala 32:22:@8.4]
  assign _T_56905 = $signed(buffer_0_354) + $signed(buffer_0_355); // @[Modules.scala 50:57:@2984.4]
  assign _T_56906 = _T_56905[10:0]; // @[Modules.scala 50:57:@2985.4]
  assign buffer_0_569 = $signed(_T_56906); // @[Modules.scala 50:57:@2986.4]
  assign buffer_0_356 = {{6{_T_56204[4]}},_T_56204}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_357 = {{6{_T_56207[4]}},_T_56207}; // @[Modules.scala 32:22:@8.4]
  assign _T_56908 = $signed(buffer_0_356) + $signed(buffer_0_357); // @[Modules.scala 50:57:@2988.4]
  assign _T_56909 = _T_56908[10:0]; // @[Modules.scala 50:57:@2989.4]
  assign buffer_0_570 = $signed(_T_56909); // @[Modules.scala 50:57:@2990.4]
  assign buffer_0_358 = {{6{_T_56210[4]}},_T_56210}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_359 = {{6{_T_56213[4]}},_T_56213}; // @[Modules.scala 32:22:@8.4]
  assign _T_56911 = $signed(buffer_0_358) + $signed(buffer_0_359); // @[Modules.scala 50:57:@2992.4]
  assign _T_56912 = _T_56911[10:0]; // @[Modules.scala 50:57:@2993.4]
  assign buffer_0_571 = $signed(_T_56912); // @[Modules.scala 50:57:@2994.4]
  assign buffer_0_360 = {{6{_T_56216[4]}},_T_56216}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_361 = {{6{_T_56219[4]}},_T_56219}; // @[Modules.scala 32:22:@8.4]
  assign _T_56914 = $signed(buffer_0_360) + $signed(buffer_0_361); // @[Modules.scala 50:57:@2996.4]
  assign _T_56915 = _T_56914[10:0]; // @[Modules.scala 50:57:@2997.4]
  assign buffer_0_572 = $signed(_T_56915); // @[Modules.scala 50:57:@2998.4]
  assign buffer_0_362 = {{6{_T_56222[4]}},_T_56222}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_363 = {{6{_T_56229[4]}},_T_56229}; // @[Modules.scala 32:22:@8.4]
  assign _T_56917 = $signed(buffer_0_362) + $signed(buffer_0_363); // @[Modules.scala 50:57:@3000.4]
  assign _T_56918 = _T_56917[10:0]; // @[Modules.scala 50:57:@3001.4]
  assign buffer_0_573 = $signed(_T_56918); // @[Modules.scala 50:57:@3002.4]
  assign buffer_0_364 = {{6{_T_56232[4]}},_T_56232}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_365 = {{6{_T_56239[4]}},_T_56239}; // @[Modules.scala 32:22:@8.4]
  assign _T_56920 = $signed(buffer_0_364) + $signed(buffer_0_365); // @[Modules.scala 50:57:@3004.4]
  assign _T_56921 = _T_56920[10:0]; // @[Modules.scala 50:57:@3005.4]
  assign buffer_0_574 = $signed(_T_56921); // @[Modules.scala 50:57:@3006.4]
  assign buffer_0_366 = {{6{_T_56242[4]}},_T_56242}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_367 = {{6{_T_56245[4]}},_T_56245}; // @[Modules.scala 32:22:@8.4]
  assign _T_56923 = $signed(buffer_0_366) + $signed(buffer_0_367); // @[Modules.scala 50:57:@3008.4]
  assign _T_56924 = _T_56923[10:0]; // @[Modules.scala 50:57:@3009.4]
  assign buffer_0_575 = $signed(_T_56924); // @[Modules.scala 50:57:@3010.4]
  assign buffer_0_368 = {{6{_T_56252[4]}},_T_56252}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_369 = {{6{_T_56259[4]}},_T_56259}; // @[Modules.scala 32:22:@8.4]
  assign _T_56926 = $signed(buffer_0_368) + $signed(buffer_0_369); // @[Modules.scala 50:57:@3012.4]
  assign _T_56927 = _T_56926[10:0]; // @[Modules.scala 50:57:@3013.4]
  assign buffer_0_576 = $signed(_T_56927); // @[Modules.scala 50:57:@3014.4]
  assign buffer_0_370 = {{6{_T_56262[4]}},_T_56262}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_371 = {{6{_T_56265[4]}},_T_56265}; // @[Modules.scala 32:22:@8.4]
  assign _T_56929 = $signed(buffer_0_370) + $signed(buffer_0_371); // @[Modules.scala 50:57:@3016.4]
  assign _T_56930 = _T_56929[10:0]; // @[Modules.scala 50:57:@3017.4]
  assign buffer_0_577 = $signed(_T_56930); // @[Modules.scala 50:57:@3018.4]
  assign buffer_0_372 = {{6{_T_56272[4]}},_T_56272}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_373 = {{6{_T_56279[4]}},_T_56279}; // @[Modules.scala 32:22:@8.4]
  assign _T_56932 = $signed(buffer_0_372) + $signed(buffer_0_373); // @[Modules.scala 50:57:@3020.4]
  assign _T_56933 = _T_56932[10:0]; // @[Modules.scala 50:57:@3021.4]
  assign buffer_0_578 = $signed(_T_56933); // @[Modules.scala 50:57:@3022.4]
  assign buffer_0_374 = {{6{_T_56282[4]}},_T_56282}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_375 = {{6{_T_56285[4]}},_T_56285}; // @[Modules.scala 32:22:@8.4]
  assign _T_56935 = $signed(buffer_0_374) + $signed(buffer_0_375); // @[Modules.scala 50:57:@3024.4]
  assign _T_56936 = _T_56935[10:0]; // @[Modules.scala 50:57:@3025.4]
  assign buffer_0_579 = $signed(_T_56936); // @[Modules.scala 50:57:@3026.4]
  assign buffer_0_376 = {{6{_T_56288[4]}},_T_56288}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_377 = {{6{_T_56291[4]}},_T_56291}; // @[Modules.scala 32:22:@8.4]
  assign _T_56938 = $signed(buffer_0_376) + $signed(buffer_0_377); // @[Modules.scala 50:57:@3028.4]
  assign _T_56939 = _T_56938[10:0]; // @[Modules.scala 50:57:@3029.4]
  assign buffer_0_580 = $signed(_T_56939); // @[Modules.scala 50:57:@3030.4]
  assign buffer_0_378 = {{6{_T_56298[4]}},_T_56298}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_379 = {{6{_T_56305[4]}},_T_56305}; // @[Modules.scala 32:22:@8.4]
  assign _T_56941 = $signed(buffer_0_378) + $signed(buffer_0_379); // @[Modules.scala 50:57:@3032.4]
  assign _T_56942 = _T_56941[10:0]; // @[Modules.scala 50:57:@3033.4]
  assign buffer_0_581 = $signed(_T_56942); // @[Modules.scala 50:57:@3034.4]
  assign buffer_0_380 = {{6{_T_56308[4]}},_T_56308}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_381 = {{6{_T_56315[4]}},_T_56315}; // @[Modules.scala 32:22:@8.4]
  assign _T_56944 = $signed(buffer_0_380) + $signed(buffer_0_381); // @[Modules.scala 50:57:@3036.4]
  assign _T_56945 = _T_56944[10:0]; // @[Modules.scala 50:57:@3037.4]
  assign buffer_0_582 = $signed(_T_56945); // @[Modules.scala 50:57:@3038.4]
  assign buffer_0_382 = {{6{_T_56322[4]}},_T_56322}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_383 = {{6{_T_56329[4]}},_T_56329}; // @[Modules.scala 32:22:@8.4]
  assign _T_56947 = $signed(buffer_0_382) + $signed(buffer_0_383); // @[Modules.scala 50:57:@3040.4]
  assign _T_56948 = _T_56947[10:0]; // @[Modules.scala 50:57:@3041.4]
  assign buffer_0_583 = $signed(_T_56948); // @[Modules.scala 50:57:@3042.4]
  assign buffer_0_384 = {{6{_T_56332[4]}},_T_56332}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_385 = {{6{_T_56339[4]}},_T_56339}; // @[Modules.scala 32:22:@8.4]
  assign _T_56950 = $signed(buffer_0_384) + $signed(buffer_0_385); // @[Modules.scala 50:57:@3044.4]
  assign _T_56951 = _T_56950[10:0]; // @[Modules.scala 50:57:@3045.4]
  assign buffer_0_584 = $signed(_T_56951); // @[Modules.scala 50:57:@3046.4]
  assign buffer_0_386 = {{6{_T_56346[4]}},_T_56346}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_387 = {{6{_T_56353[4]}},_T_56353}; // @[Modules.scala 32:22:@8.4]
  assign _T_56953 = $signed(buffer_0_386) + $signed(buffer_0_387); // @[Modules.scala 50:57:@3048.4]
  assign _T_56954 = _T_56953[10:0]; // @[Modules.scala 50:57:@3049.4]
  assign buffer_0_585 = $signed(_T_56954); // @[Modules.scala 50:57:@3050.4]
  assign buffer_0_388 = {{6{_T_56356[4]}},_T_56356}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_389 = {{6{_T_56363[4]}},_T_56363}; // @[Modules.scala 32:22:@8.4]
  assign _T_56956 = $signed(buffer_0_388) + $signed(buffer_0_389); // @[Modules.scala 50:57:@3052.4]
  assign _T_56957 = _T_56956[10:0]; // @[Modules.scala 50:57:@3053.4]
  assign buffer_0_586 = $signed(_T_56957); // @[Modules.scala 50:57:@3054.4]
  assign buffer_0_390 = {{6{_T_56370[4]}},_T_56370}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_391 = {{6{_T_56373[4]}},_T_56373}; // @[Modules.scala 32:22:@8.4]
  assign _T_56959 = $signed(buffer_0_390) + $signed(buffer_0_391); // @[Modules.scala 50:57:@3056.4]
  assign _T_56960 = _T_56959[10:0]; // @[Modules.scala 50:57:@3057.4]
  assign buffer_0_587 = $signed(_T_56960); // @[Modules.scala 50:57:@3058.4]
  assign _T_56962 = $signed(buffer_0_392) + $signed(buffer_0_393); // @[Modules.scala 53:83:@3060.4]
  assign _T_56963 = _T_56962[10:0]; // @[Modules.scala 53:83:@3061.4]
  assign buffer_0_588 = $signed(_T_56963); // @[Modules.scala 53:83:@3062.4]
  assign _T_56965 = $signed(buffer_0_394) + $signed(buffer_0_395); // @[Modules.scala 53:83:@3064.4]
  assign _T_56966 = _T_56965[10:0]; // @[Modules.scala 53:83:@3065.4]
  assign buffer_0_589 = $signed(_T_56966); // @[Modules.scala 53:83:@3066.4]
  assign _T_56968 = $signed(buffer_0_396) + $signed(buffer_0_397); // @[Modules.scala 53:83:@3068.4]
  assign _T_56969 = _T_56968[10:0]; // @[Modules.scala 53:83:@3069.4]
  assign buffer_0_590 = $signed(_T_56969); // @[Modules.scala 53:83:@3070.4]
  assign _T_56971 = $signed(buffer_0_398) + $signed(buffer_0_399); // @[Modules.scala 53:83:@3072.4]
  assign _T_56972 = _T_56971[10:0]; // @[Modules.scala 53:83:@3073.4]
  assign buffer_0_591 = $signed(_T_56972); // @[Modules.scala 53:83:@3074.4]
  assign _T_56974 = $signed(buffer_0_400) + $signed(buffer_0_401); // @[Modules.scala 53:83:@3076.4]
  assign _T_56975 = _T_56974[10:0]; // @[Modules.scala 53:83:@3077.4]
  assign buffer_0_592 = $signed(_T_56975); // @[Modules.scala 53:83:@3078.4]
  assign _T_56977 = $signed(buffer_0_402) + $signed(buffer_0_403); // @[Modules.scala 53:83:@3080.4]
  assign _T_56978 = _T_56977[10:0]; // @[Modules.scala 53:83:@3081.4]
  assign buffer_0_593 = $signed(_T_56978); // @[Modules.scala 53:83:@3082.4]
  assign _T_56980 = $signed(buffer_0_404) + $signed(buffer_0_405); // @[Modules.scala 53:83:@3084.4]
  assign _T_56981 = _T_56980[10:0]; // @[Modules.scala 53:83:@3085.4]
  assign buffer_0_594 = $signed(_T_56981); // @[Modules.scala 53:83:@3086.4]
  assign _T_56983 = $signed(buffer_0_406) + $signed(buffer_0_407); // @[Modules.scala 53:83:@3088.4]
  assign _T_56984 = _T_56983[10:0]; // @[Modules.scala 53:83:@3089.4]
  assign buffer_0_595 = $signed(_T_56984); // @[Modules.scala 53:83:@3090.4]
  assign _T_56986 = $signed(buffer_0_408) + $signed(buffer_0_409); // @[Modules.scala 53:83:@3092.4]
  assign _T_56987 = _T_56986[10:0]; // @[Modules.scala 53:83:@3093.4]
  assign buffer_0_596 = $signed(_T_56987); // @[Modules.scala 53:83:@3094.4]
  assign _T_56989 = $signed(buffer_0_410) + $signed(buffer_0_411); // @[Modules.scala 53:83:@3096.4]
  assign _T_56990 = _T_56989[10:0]; // @[Modules.scala 53:83:@3097.4]
  assign buffer_0_597 = $signed(_T_56990); // @[Modules.scala 53:83:@3098.4]
  assign _T_56992 = $signed(buffer_0_412) + $signed(buffer_0_413); // @[Modules.scala 53:83:@3100.4]
  assign _T_56993 = _T_56992[10:0]; // @[Modules.scala 53:83:@3101.4]
  assign buffer_0_598 = $signed(_T_56993); // @[Modules.scala 53:83:@3102.4]
  assign _T_56995 = $signed(buffer_0_414) + $signed(buffer_0_415); // @[Modules.scala 53:83:@3104.4]
  assign _T_56996 = _T_56995[10:0]; // @[Modules.scala 53:83:@3105.4]
  assign buffer_0_599 = $signed(_T_56996); // @[Modules.scala 53:83:@3106.4]
  assign _T_56998 = $signed(buffer_0_416) + $signed(buffer_0_417); // @[Modules.scala 53:83:@3108.4]
  assign _T_56999 = _T_56998[10:0]; // @[Modules.scala 53:83:@3109.4]
  assign buffer_0_600 = $signed(_T_56999); // @[Modules.scala 53:83:@3110.4]
  assign _T_57001 = $signed(buffer_0_418) + $signed(buffer_0_419); // @[Modules.scala 53:83:@3112.4]
  assign _T_57002 = _T_57001[10:0]; // @[Modules.scala 53:83:@3113.4]
  assign buffer_0_601 = $signed(_T_57002); // @[Modules.scala 53:83:@3114.4]
  assign _T_57004 = $signed(buffer_0_420) + $signed(buffer_0_421); // @[Modules.scala 53:83:@3116.4]
  assign _T_57005 = _T_57004[10:0]; // @[Modules.scala 53:83:@3117.4]
  assign buffer_0_602 = $signed(_T_57005); // @[Modules.scala 53:83:@3118.4]
  assign _T_57007 = $signed(buffer_0_422) + $signed(buffer_0_423); // @[Modules.scala 53:83:@3120.4]
  assign _T_57008 = _T_57007[10:0]; // @[Modules.scala 53:83:@3121.4]
  assign buffer_0_603 = $signed(_T_57008); // @[Modules.scala 53:83:@3122.4]
  assign _T_57010 = $signed(buffer_0_424) + $signed(buffer_0_425); // @[Modules.scala 53:83:@3124.4]
  assign _T_57011 = _T_57010[10:0]; // @[Modules.scala 53:83:@3125.4]
  assign buffer_0_604 = $signed(_T_57011); // @[Modules.scala 53:83:@3126.4]
  assign _T_57013 = $signed(buffer_0_426) + $signed(buffer_0_427); // @[Modules.scala 53:83:@3128.4]
  assign _T_57014 = _T_57013[10:0]; // @[Modules.scala 53:83:@3129.4]
  assign buffer_0_605 = $signed(_T_57014); // @[Modules.scala 53:83:@3130.4]
  assign _T_57016 = $signed(buffer_0_428) + $signed(buffer_0_429); // @[Modules.scala 53:83:@3132.4]
  assign _T_57017 = _T_57016[10:0]; // @[Modules.scala 53:83:@3133.4]
  assign buffer_0_606 = $signed(_T_57017); // @[Modules.scala 53:83:@3134.4]
  assign _T_57019 = $signed(buffer_0_430) + $signed(buffer_0_431); // @[Modules.scala 53:83:@3136.4]
  assign _T_57020 = _T_57019[10:0]; // @[Modules.scala 53:83:@3137.4]
  assign buffer_0_607 = $signed(_T_57020); // @[Modules.scala 53:83:@3138.4]
  assign _T_57022 = $signed(buffer_0_432) + $signed(buffer_0_433); // @[Modules.scala 53:83:@3140.4]
  assign _T_57023 = _T_57022[10:0]; // @[Modules.scala 53:83:@3141.4]
  assign buffer_0_608 = $signed(_T_57023); // @[Modules.scala 53:83:@3142.4]
  assign _T_57025 = $signed(buffer_0_434) + $signed(buffer_0_435); // @[Modules.scala 53:83:@3144.4]
  assign _T_57026 = _T_57025[10:0]; // @[Modules.scala 53:83:@3145.4]
  assign buffer_0_609 = $signed(_T_57026); // @[Modules.scala 53:83:@3146.4]
  assign _T_57028 = $signed(buffer_0_436) + $signed(buffer_0_437); // @[Modules.scala 53:83:@3148.4]
  assign _T_57029 = _T_57028[10:0]; // @[Modules.scala 53:83:@3149.4]
  assign buffer_0_610 = $signed(_T_57029); // @[Modules.scala 53:83:@3150.4]
  assign _T_57031 = $signed(buffer_0_438) + $signed(buffer_0_439); // @[Modules.scala 53:83:@3152.4]
  assign _T_57032 = _T_57031[10:0]; // @[Modules.scala 53:83:@3153.4]
  assign buffer_0_611 = $signed(_T_57032); // @[Modules.scala 53:83:@3154.4]
  assign _T_57034 = $signed(buffer_0_440) + $signed(buffer_0_441); // @[Modules.scala 53:83:@3156.4]
  assign _T_57035 = _T_57034[10:0]; // @[Modules.scala 53:83:@3157.4]
  assign buffer_0_612 = $signed(_T_57035); // @[Modules.scala 53:83:@3158.4]
  assign _T_57037 = $signed(buffer_0_442) + $signed(buffer_0_443); // @[Modules.scala 53:83:@3160.4]
  assign _T_57038 = _T_57037[10:0]; // @[Modules.scala 53:83:@3161.4]
  assign buffer_0_613 = $signed(_T_57038); // @[Modules.scala 53:83:@3162.4]
  assign _T_57040 = $signed(buffer_0_444) + $signed(buffer_0_445); // @[Modules.scala 53:83:@3164.4]
  assign _T_57041 = _T_57040[10:0]; // @[Modules.scala 53:83:@3165.4]
  assign buffer_0_614 = $signed(_T_57041); // @[Modules.scala 53:83:@3166.4]
  assign _T_57043 = $signed(buffer_0_446) + $signed(buffer_0_447); // @[Modules.scala 53:83:@3168.4]
  assign _T_57044 = _T_57043[10:0]; // @[Modules.scala 53:83:@3169.4]
  assign buffer_0_615 = $signed(_T_57044); // @[Modules.scala 53:83:@3170.4]
  assign _T_57046 = $signed(buffer_0_448) + $signed(buffer_0_449); // @[Modules.scala 53:83:@3172.4]
  assign _T_57047 = _T_57046[10:0]; // @[Modules.scala 53:83:@3173.4]
  assign buffer_0_616 = $signed(_T_57047); // @[Modules.scala 53:83:@3174.4]
  assign _T_57049 = $signed(buffer_0_450) + $signed(buffer_0_451); // @[Modules.scala 53:83:@3176.4]
  assign _T_57050 = _T_57049[10:0]; // @[Modules.scala 53:83:@3177.4]
  assign buffer_0_617 = $signed(_T_57050); // @[Modules.scala 53:83:@3178.4]
  assign _T_57052 = $signed(buffer_0_452) + $signed(buffer_0_453); // @[Modules.scala 53:83:@3180.4]
  assign _T_57053 = _T_57052[10:0]; // @[Modules.scala 53:83:@3181.4]
  assign buffer_0_618 = $signed(_T_57053); // @[Modules.scala 53:83:@3182.4]
  assign _T_57055 = $signed(buffer_0_454) + $signed(buffer_0_455); // @[Modules.scala 53:83:@3184.4]
  assign _T_57056 = _T_57055[10:0]; // @[Modules.scala 53:83:@3185.4]
  assign buffer_0_619 = $signed(_T_57056); // @[Modules.scala 53:83:@3186.4]
  assign _T_57058 = $signed(buffer_0_456) + $signed(buffer_0_457); // @[Modules.scala 53:83:@3188.4]
  assign _T_57059 = _T_57058[10:0]; // @[Modules.scala 53:83:@3189.4]
  assign buffer_0_620 = $signed(_T_57059); // @[Modules.scala 53:83:@3190.4]
  assign _T_57061 = $signed(buffer_0_458) + $signed(buffer_0_459); // @[Modules.scala 53:83:@3192.4]
  assign _T_57062 = _T_57061[10:0]; // @[Modules.scala 53:83:@3193.4]
  assign buffer_0_621 = $signed(_T_57062); // @[Modules.scala 53:83:@3194.4]
  assign _T_57064 = $signed(buffer_0_460) + $signed(buffer_0_461); // @[Modules.scala 53:83:@3196.4]
  assign _T_57065 = _T_57064[10:0]; // @[Modules.scala 53:83:@3197.4]
  assign buffer_0_622 = $signed(_T_57065); // @[Modules.scala 53:83:@3198.4]
  assign _T_57067 = $signed(buffer_0_462) + $signed(buffer_0_463); // @[Modules.scala 53:83:@3200.4]
  assign _T_57068 = _T_57067[10:0]; // @[Modules.scala 53:83:@3201.4]
  assign buffer_0_623 = $signed(_T_57068); // @[Modules.scala 53:83:@3202.4]
  assign _T_57070 = $signed(buffer_0_464) + $signed(buffer_0_465); // @[Modules.scala 53:83:@3204.4]
  assign _T_57071 = _T_57070[10:0]; // @[Modules.scala 53:83:@3205.4]
  assign buffer_0_624 = $signed(_T_57071); // @[Modules.scala 53:83:@3206.4]
  assign _T_57073 = $signed(buffer_0_466) + $signed(buffer_0_467); // @[Modules.scala 53:83:@3208.4]
  assign _T_57074 = _T_57073[10:0]; // @[Modules.scala 53:83:@3209.4]
  assign buffer_0_625 = $signed(_T_57074); // @[Modules.scala 53:83:@3210.4]
  assign _T_57076 = $signed(buffer_0_468) + $signed(buffer_0_469); // @[Modules.scala 53:83:@3212.4]
  assign _T_57077 = _T_57076[10:0]; // @[Modules.scala 53:83:@3213.4]
  assign buffer_0_626 = $signed(_T_57077); // @[Modules.scala 53:83:@3214.4]
  assign _T_57079 = $signed(buffer_0_470) + $signed(buffer_0_471); // @[Modules.scala 53:83:@3216.4]
  assign _T_57080 = _T_57079[10:0]; // @[Modules.scala 53:83:@3217.4]
  assign buffer_0_627 = $signed(_T_57080); // @[Modules.scala 53:83:@3218.4]
  assign _T_57082 = $signed(buffer_0_472) + $signed(buffer_0_473); // @[Modules.scala 53:83:@3220.4]
  assign _T_57083 = _T_57082[10:0]; // @[Modules.scala 53:83:@3221.4]
  assign buffer_0_628 = $signed(_T_57083); // @[Modules.scala 53:83:@3222.4]
  assign _T_57085 = $signed(buffer_0_474) + $signed(buffer_0_475); // @[Modules.scala 53:83:@3224.4]
  assign _T_57086 = _T_57085[10:0]; // @[Modules.scala 53:83:@3225.4]
  assign buffer_0_629 = $signed(_T_57086); // @[Modules.scala 53:83:@3226.4]
  assign _T_57088 = $signed(buffer_0_476) + $signed(buffer_0_477); // @[Modules.scala 53:83:@3228.4]
  assign _T_57089 = _T_57088[10:0]; // @[Modules.scala 53:83:@3229.4]
  assign buffer_0_630 = $signed(_T_57089); // @[Modules.scala 53:83:@3230.4]
  assign _T_57091 = $signed(buffer_0_478) + $signed(buffer_0_479); // @[Modules.scala 53:83:@3232.4]
  assign _T_57092 = _T_57091[10:0]; // @[Modules.scala 53:83:@3233.4]
  assign buffer_0_631 = $signed(_T_57092); // @[Modules.scala 53:83:@3234.4]
  assign _T_57094 = $signed(buffer_0_480) + $signed(buffer_0_481); // @[Modules.scala 53:83:@3236.4]
  assign _T_57095 = _T_57094[10:0]; // @[Modules.scala 53:83:@3237.4]
  assign buffer_0_632 = $signed(_T_57095); // @[Modules.scala 53:83:@3238.4]
  assign _T_57097 = $signed(buffer_0_482) + $signed(buffer_0_483); // @[Modules.scala 53:83:@3240.4]
  assign _T_57098 = _T_57097[10:0]; // @[Modules.scala 53:83:@3241.4]
  assign buffer_0_633 = $signed(_T_57098); // @[Modules.scala 53:83:@3242.4]
  assign _T_57100 = $signed(buffer_0_484) + $signed(buffer_0_485); // @[Modules.scala 53:83:@3244.4]
  assign _T_57101 = _T_57100[10:0]; // @[Modules.scala 53:83:@3245.4]
  assign buffer_0_634 = $signed(_T_57101); // @[Modules.scala 53:83:@3246.4]
  assign _T_57103 = $signed(buffer_0_486) + $signed(buffer_0_487); // @[Modules.scala 53:83:@3248.4]
  assign _T_57104 = _T_57103[10:0]; // @[Modules.scala 53:83:@3249.4]
  assign buffer_0_635 = $signed(_T_57104); // @[Modules.scala 53:83:@3250.4]
  assign _T_57106 = $signed(buffer_0_488) + $signed(buffer_0_489); // @[Modules.scala 53:83:@3252.4]
  assign _T_57107 = _T_57106[10:0]; // @[Modules.scala 53:83:@3253.4]
  assign buffer_0_636 = $signed(_T_57107); // @[Modules.scala 53:83:@3254.4]
  assign _T_57109 = $signed(buffer_0_490) + $signed(buffer_0_491); // @[Modules.scala 53:83:@3256.4]
  assign _T_57110 = _T_57109[10:0]; // @[Modules.scala 53:83:@3257.4]
  assign buffer_0_637 = $signed(_T_57110); // @[Modules.scala 53:83:@3258.4]
  assign _T_57112 = $signed(buffer_0_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@3260.4]
  assign _T_57113 = _T_57112[10:0]; // @[Modules.scala 53:83:@3261.4]
  assign buffer_0_638 = $signed(_T_57113); // @[Modules.scala 53:83:@3262.4]
  assign _T_57115 = $signed(buffer_0_494) + $signed(buffer_0_495); // @[Modules.scala 53:83:@3264.4]
  assign _T_57116 = _T_57115[10:0]; // @[Modules.scala 53:83:@3265.4]
  assign buffer_0_639 = $signed(_T_57116); // @[Modules.scala 53:83:@3266.4]
  assign _T_57118 = $signed(buffer_0_496) + $signed(buffer_0_497); // @[Modules.scala 53:83:@3268.4]
  assign _T_57119 = _T_57118[10:0]; // @[Modules.scala 53:83:@3269.4]
  assign buffer_0_640 = $signed(_T_57119); // @[Modules.scala 53:83:@3270.4]
  assign _T_57121 = $signed(buffer_0_498) + $signed(buffer_0_499); // @[Modules.scala 53:83:@3272.4]
  assign _T_57122 = _T_57121[10:0]; // @[Modules.scala 53:83:@3273.4]
  assign buffer_0_641 = $signed(_T_57122); // @[Modules.scala 53:83:@3274.4]
  assign _T_57124 = $signed(buffer_0_500) + $signed(buffer_0_501); // @[Modules.scala 53:83:@3276.4]
  assign _T_57125 = _T_57124[10:0]; // @[Modules.scala 53:83:@3277.4]
  assign buffer_0_642 = $signed(_T_57125); // @[Modules.scala 53:83:@3278.4]
  assign _T_57127 = $signed(buffer_0_502) + $signed(buffer_0_503); // @[Modules.scala 53:83:@3280.4]
  assign _T_57128 = _T_57127[10:0]; // @[Modules.scala 53:83:@3281.4]
  assign buffer_0_643 = $signed(_T_57128); // @[Modules.scala 53:83:@3282.4]
  assign _T_57130 = $signed(buffer_0_504) + $signed(buffer_0_505); // @[Modules.scala 53:83:@3284.4]
  assign _T_57131 = _T_57130[10:0]; // @[Modules.scala 53:83:@3285.4]
  assign buffer_0_644 = $signed(_T_57131); // @[Modules.scala 53:83:@3286.4]
  assign _T_57133 = $signed(buffer_0_506) + $signed(buffer_0_507); // @[Modules.scala 53:83:@3288.4]
  assign _T_57134 = _T_57133[10:0]; // @[Modules.scala 53:83:@3289.4]
  assign buffer_0_645 = $signed(_T_57134); // @[Modules.scala 53:83:@3290.4]
  assign _T_57136 = $signed(buffer_0_508) + $signed(buffer_0_509); // @[Modules.scala 53:83:@3292.4]
  assign _T_57137 = _T_57136[10:0]; // @[Modules.scala 53:83:@3293.4]
  assign buffer_0_646 = $signed(_T_57137); // @[Modules.scala 53:83:@3294.4]
  assign _T_57139 = $signed(buffer_0_510) + $signed(buffer_0_511); // @[Modules.scala 53:83:@3296.4]
  assign _T_57140 = _T_57139[10:0]; // @[Modules.scala 53:83:@3297.4]
  assign buffer_0_647 = $signed(_T_57140); // @[Modules.scala 53:83:@3298.4]
  assign _T_57142 = $signed(buffer_0_512) + $signed(buffer_0_513); // @[Modules.scala 53:83:@3300.4]
  assign _T_57143 = _T_57142[10:0]; // @[Modules.scala 53:83:@3301.4]
  assign buffer_0_648 = $signed(_T_57143); // @[Modules.scala 53:83:@3302.4]
  assign _T_57145 = $signed(buffer_0_514) + $signed(buffer_0_515); // @[Modules.scala 53:83:@3304.4]
  assign _T_57146 = _T_57145[10:0]; // @[Modules.scala 53:83:@3305.4]
  assign buffer_0_649 = $signed(_T_57146); // @[Modules.scala 53:83:@3306.4]
  assign _T_57148 = $signed(buffer_0_516) + $signed(buffer_0_517); // @[Modules.scala 53:83:@3308.4]
  assign _T_57149 = _T_57148[10:0]; // @[Modules.scala 53:83:@3309.4]
  assign buffer_0_650 = $signed(_T_57149); // @[Modules.scala 53:83:@3310.4]
  assign _T_57151 = $signed(buffer_0_518) + $signed(buffer_0_519); // @[Modules.scala 53:83:@3312.4]
  assign _T_57152 = _T_57151[10:0]; // @[Modules.scala 53:83:@3313.4]
  assign buffer_0_651 = $signed(_T_57152); // @[Modules.scala 53:83:@3314.4]
  assign _T_57154 = $signed(buffer_0_520) + $signed(buffer_0_521); // @[Modules.scala 53:83:@3316.4]
  assign _T_57155 = _T_57154[10:0]; // @[Modules.scala 53:83:@3317.4]
  assign buffer_0_652 = $signed(_T_57155); // @[Modules.scala 53:83:@3318.4]
  assign _T_57157 = $signed(buffer_0_522) + $signed(buffer_0_523); // @[Modules.scala 53:83:@3320.4]
  assign _T_57158 = _T_57157[10:0]; // @[Modules.scala 53:83:@3321.4]
  assign buffer_0_653 = $signed(_T_57158); // @[Modules.scala 53:83:@3322.4]
  assign _T_57160 = $signed(buffer_0_524) + $signed(buffer_0_525); // @[Modules.scala 53:83:@3324.4]
  assign _T_57161 = _T_57160[10:0]; // @[Modules.scala 53:83:@3325.4]
  assign buffer_0_654 = $signed(_T_57161); // @[Modules.scala 53:83:@3326.4]
  assign _T_57163 = $signed(buffer_0_526) + $signed(buffer_0_527); // @[Modules.scala 53:83:@3328.4]
  assign _T_57164 = _T_57163[10:0]; // @[Modules.scala 53:83:@3329.4]
  assign buffer_0_655 = $signed(_T_57164); // @[Modules.scala 53:83:@3330.4]
  assign _T_57166 = $signed(buffer_0_528) + $signed(buffer_0_529); // @[Modules.scala 53:83:@3332.4]
  assign _T_57167 = _T_57166[10:0]; // @[Modules.scala 53:83:@3333.4]
  assign buffer_0_656 = $signed(_T_57167); // @[Modules.scala 53:83:@3334.4]
  assign _T_57169 = $signed(buffer_0_530) + $signed(buffer_0_531); // @[Modules.scala 53:83:@3336.4]
  assign _T_57170 = _T_57169[10:0]; // @[Modules.scala 53:83:@3337.4]
  assign buffer_0_657 = $signed(_T_57170); // @[Modules.scala 53:83:@3338.4]
  assign _T_57172 = $signed(buffer_0_532) + $signed(buffer_0_533); // @[Modules.scala 53:83:@3340.4]
  assign _T_57173 = _T_57172[10:0]; // @[Modules.scala 53:83:@3341.4]
  assign buffer_0_658 = $signed(_T_57173); // @[Modules.scala 53:83:@3342.4]
  assign _T_57175 = $signed(buffer_0_534) + $signed(buffer_0_535); // @[Modules.scala 53:83:@3344.4]
  assign _T_57176 = _T_57175[10:0]; // @[Modules.scala 53:83:@3345.4]
  assign buffer_0_659 = $signed(_T_57176); // @[Modules.scala 53:83:@3346.4]
  assign _T_57178 = $signed(buffer_0_536) + $signed(buffer_0_537); // @[Modules.scala 53:83:@3348.4]
  assign _T_57179 = _T_57178[10:0]; // @[Modules.scala 53:83:@3349.4]
  assign buffer_0_660 = $signed(_T_57179); // @[Modules.scala 53:83:@3350.4]
  assign _T_57181 = $signed(buffer_0_538) + $signed(buffer_0_539); // @[Modules.scala 53:83:@3352.4]
  assign _T_57182 = _T_57181[10:0]; // @[Modules.scala 53:83:@3353.4]
  assign buffer_0_661 = $signed(_T_57182); // @[Modules.scala 53:83:@3354.4]
  assign _T_57184 = $signed(buffer_0_540) + $signed(buffer_0_541); // @[Modules.scala 53:83:@3356.4]
  assign _T_57185 = _T_57184[10:0]; // @[Modules.scala 53:83:@3357.4]
  assign buffer_0_662 = $signed(_T_57185); // @[Modules.scala 53:83:@3358.4]
  assign _T_57187 = $signed(buffer_0_542) + $signed(buffer_0_543); // @[Modules.scala 53:83:@3360.4]
  assign _T_57188 = _T_57187[10:0]; // @[Modules.scala 53:83:@3361.4]
  assign buffer_0_663 = $signed(_T_57188); // @[Modules.scala 53:83:@3362.4]
  assign _T_57190 = $signed(buffer_0_544) + $signed(buffer_0_545); // @[Modules.scala 53:83:@3364.4]
  assign _T_57191 = _T_57190[10:0]; // @[Modules.scala 53:83:@3365.4]
  assign buffer_0_664 = $signed(_T_57191); // @[Modules.scala 53:83:@3366.4]
  assign _T_57193 = $signed(buffer_0_546) + $signed(buffer_0_547); // @[Modules.scala 53:83:@3368.4]
  assign _T_57194 = _T_57193[10:0]; // @[Modules.scala 53:83:@3369.4]
  assign buffer_0_665 = $signed(_T_57194); // @[Modules.scala 53:83:@3370.4]
  assign _T_57196 = $signed(buffer_0_548) + $signed(buffer_0_549); // @[Modules.scala 53:83:@3372.4]
  assign _T_57197 = _T_57196[10:0]; // @[Modules.scala 53:83:@3373.4]
  assign buffer_0_666 = $signed(_T_57197); // @[Modules.scala 53:83:@3374.4]
  assign _T_57199 = $signed(buffer_0_550) + $signed(buffer_0_551); // @[Modules.scala 53:83:@3376.4]
  assign _T_57200 = _T_57199[10:0]; // @[Modules.scala 53:83:@3377.4]
  assign buffer_0_667 = $signed(_T_57200); // @[Modules.scala 53:83:@3378.4]
  assign _T_57202 = $signed(buffer_0_552) + $signed(buffer_0_553); // @[Modules.scala 53:83:@3380.4]
  assign _T_57203 = _T_57202[10:0]; // @[Modules.scala 53:83:@3381.4]
  assign buffer_0_668 = $signed(_T_57203); // @[Modules.scala 53:83:@3382.4]
  assign _T_57205 = $signed(buffer_0_554) + $signed(buffer_0_555); // @[Modules.scala 53:83:@3384.4]
  assign _T_57206 = _T_57205[10:0]; // @[Modules.scala 53:83:@3385.4]
  assign buffer_0_669 = $signed(_T_57206); // @[Modules.scala 53:83:@3386.4]
  assign _T_57208 = $signed(buffer_0_556) + $signed(buffer_0_557); // @[Modules.scala 53:83:@3388.4]
  assign _T_57209 = _T_57208[10:0]; // @[Modules.scala 53:83:@3389.4]
  assign buffer_0_670 = $signed(_T_57209); // @[Modules.scala 53:83:@3390.4]
  assign _T_57211 = $signed(buffer_0_558) + $signed(buffer_0_559); // @[Modules.scala 53:83:@3392.4]
  assign _T_57212 = _T_57211[10:0]; // @[Modules.scala 53:83:@3393.4]
  assign buffer_0_671 = $signed(_T_57212); // @[Modules.scala 53:83:@3394.4]
  assign _T_57214 = $signed(buffer_0_560) + $signed(buffer_0_561); // @[Modules.scala 53:83:@3396.4]
  assign _T_57215 = _T_57214[10:0]; // @[Modules.scala 53:83:@3397.4]
  assign buffer_0_672 = $signed(_T_57215); // @[Modules.scala 53:83:@3398.4]
  assign _T_57217 = $signed(buffer_0_562) + $signed(buffer_0_563); // @[Modules.scala 53:83:@3400.4]
  assign _T_57218 = _T_57217[10:0]; // @[Modules.scala 53:83:@3401.4]
  assign buffer_0_673 = $signed(_T_57218); // @[Modules.scala 53:83:@3402.4]
  assign _T_57220 = $signed(buffer_0_564) + $signed(buffer_0_565); // @[Modules.scala 53:83:@3404.4]
  assign _T_57221 = _T_57220[10:0]; // @[Modules.scala 53:83:@3405.4]
  assign buffer_0_674 = $signed(_T_57221); // @[Modules.scala 53:83:@3406.4]
  assign _T_57223 = $signed(buffer_0_566) + $signed(buffer_0_567); // @[Modules.scala 53:83:@3408.4]
  assign _T_57224 = _T_57223[10:0]; // @[Modules.scala 53:83:@3409.4]
  assign buffer_0_675 = $signed(_T_57224); // @[Modules.scala 53:83:@3410.4]
  assign _T_57226 = $signed(buffer_0_568) + $signed(buffer_0_569); // @[Modules.scala 53:83:@3412.4]
  assign _T_57227 = _T_57226[10:0]; // @[Modules.scala 53:83:@3413.4]
  assign buffer_0_676 = $signed(_T_57227); // @[Modules.scala 53:83:@3414.4]
  assign _T_57229 = $signed(buffer_0_570) + $signed(buffer_0_571); // @[Modules.scala 53:83:@3416.4]
  assign _T_57230 = _T_57229[10:0]; // @[Modules.scala 53:83:@3417.4]
  assign buffer_0_677 = $signed(_T_57230); // @[Modules.scala 53:83:@3418.4]
  assign _T_57232 = $signed(buffer_0_572) + $signed(buffer_0_573); // @[Modules.scala 53:83:@3420.4]
  assign _T_57233 = _T_57232[10:0]; // @[Modules.scala 53:83:@3421.4]
  assign buffer_0_678 = $signed(_T_57233); // @[Modules.scala 53:83:@3422.4]
  assign _T_57235 = $signed(buffer_0_574) + $signed(buffer_0_575); // @[Modules.scala 53:83:@3424.4]
  assign _T_57236 = _T_57235[10:0]; // @[Modules.scala 53:83:@3425.4]
  assign buffer_0_679 = $signed(_T_57236); // @[Modules.scala 53:83:@3426.4]
  assign _T_57238 = $signed(buffer_0_576) + $signed(buffer_0_577); // @[Modules.scala 53:83:@3428.4]
  assign _T_57239 = _T_57238[10:0]; // @[Modules.scala 53:83:@3429.4]
  assign buffer_0_680 = $signed(_T_57239); // @[Modules.scala 53:83:@3430.4]
  assign _T_57241 = $signed(buffer_0_578) + $signed(buffer_0_579); // @[Modules.scala 53:83:@3432.4]
  assign _T_57242 = _T_57241[10:0]; // @[Modules.scala 53:83:@3433.4]
  assign buffer_0_681 = $signed(_T_57242); // @[Modules.scala 53:83:@3434.4]
  assign _T_57244 = $signed(buffer_0_580) + $signed(buffer_0_581); // @[Modules.scala 53:83:@3436.4]
  assign _T_57245 = _T_57244[10:0]; // @[Modules.scala 53:83:@3437.4]
  assign buffer_0_682 = $signed(_T_57245); // @[Modules.scala 53:83:@3438.4]
  assign _T_57247 = $signed(buffer_0_582) + $signed(buffer_0_583); // @[Modules.scala 53:83:@3440.4]
  assign _T_57248 = _T_57247[10:0]; // @[Modules.scala 53:83:@3441.4]
  assign buffer_0_683 = $signed(_T_57248); // @[Modules.scala 53:83:@3442.4]
  assign _T_57250 = $signed(buffer_0_584) + $signed(buffer_0_585); // @[Modules.scala 53:83:@3444.4]
  assign _T_57251 = _T_57250[10:0]; // @[Modules.scala 53:83:@3445.4]
  assign buffer_0_684 = $signed(_T_57251); // @[Modules.scala 53:83:@3446.4]
  assign _T_57253 = $signed(buffer_0_586) + $signed(buffer_0_587); // @[Modules.scala 53:83:@3448.4]
  assign _T_57254 = _T_57253[10:0]; // @[Modules.scala 53:83:@3449.4]
  assign buffer_0_685 = $signed(_T_57254); // @[Modules.scala 53:83:@3450.4]
  assign _T_57256 = $signed(buffer_0_588) + $signed(buffer_0_589); // @[Modules.scala 56:109:@3452.4]
  assign _T_57257 = _T_57256[10:0]; // @[Modules.scala 56:109:@3453.4]
  assign buffer_0_686 = $signed(_T_57257); // @[Modules.scala 56:109:@3454.4]
  assign _T_57259 = $signed(buffer_0_590) + $signed(buffer_0_591); // @[Modules.scala 56:109:@3456.4]
  assign _T_57260 = _T_57259[10:0]; // @[Modules.scala 56:109:@3457.4]
  assign buffer_0_687 = $signed(_T_57260); // @[Modules.scala 56:109:@3458.4]
  assign _T_57262 = $signed(buffer_0_592) + $signed(buffer_0_593); // @[Modules.scala 56:109:@3460.4]
  assign _T_57263 = _T_57262[10:0]; // @[Modules.scala 56:109:@3461.4]
  assign buffer_0_688 = $signed(_T_57263); // @[Modules.scala 56:109:@3462.4]
  assign _T_57265 = $signed(buffer_0_594) + $signed(buffer_0_595); // @[Modules.scala 56:109:@3464.4]
  assign _T_57266 = _T_57265[10:0]; // @[Modules.scala 56:109:@3465.4]
  assign buffer_0_689 = $signed(_T_57266); // @[Modules.scala 56:109:@3466.4]
  assign _T_57268 = $signed(buffer_0_596) + $signed(buffer_0_597); // @[Modules.scala 56:109:@3468.4]
  assign _T_57269 = _T_57268[10:0]; // @[Modules.scala 56:109:@3469.4]
  assign buffer_0_690 = $signed(_T_57269); // @[Modules.scala 56:109:@3470.4]
  assign _T_57271 = $signed(buffer_0_598) + $signed(buffer_0_599); // @[Modules.scala 56:109:@3472.4]
  assign _T_57272 = _T_57271[10:0]; // @[Modules.scala 56:109:@3473.4]
  assign buffer_0_691 = $signed(_T_57272); // @[Modules.scala 56:109:@3474.4]
  assign _T_57274 = $signed(buffer_0_600) + $signed(buffer_0_601); // @[Modules.scala 56:109:@3476.4]
  assign _T_57275 = _T_57274[10:0]; // @[Modules.scala 56:109:@3477.4]
  assign buffer_0_692 = $signed(_T_57275); // @[Modules.scala 56:109:@3478.4]
  assign _T_57277 = $signed(buffer_0_602) + $signed(buffer_0_603); // @[Modules.scala 56:109:@3480.4]
  assign _T_57278 = _T_57277[10:0]; // @[Modules.scala 56:109:@3481.4]
  assign buffer_0_693 = $signed(_T_57278); // @[Modules.scala 56:109:@3482.4]
  assign _T_57280 = $signed(buffer_0_604) + $signed(buffer_0_605); // @[Modules.scala 56:109:@3484.4]
  assign _T_57281 = _T_57280[10:0]; // @[Modules.scala 56:109:@3485.4]
  assign buffer_0_694 = $signed(_T_57281); // @[Modules.scala 56:109:@3486.4]
  assign _T_57283 = $signed(buffer_0_606) + $signed(buffer_0_607); // @[Modules.scala 56:109:@3488.4]
  assign _T_57284 = _T_57283[10:0]; // @[Modules.scala 56:109:@3489.4]
  assign buffer_0_695 = $signed(_T_57284); // @[Modules.scala 56:109:@3490.4]
  assign _T_57286 = $signed(buffer_0_608) + $signed(buffer_0_609); // @[Modules.scala 56:109:@3492.4]
  assign _T_57287 = _T_57286[10:0]; // @[Modules.scala 56:109:@3493.4]
  assign buffer_0_696 = $signed(_T_57287); // @[Modules.scala 56:109:@3494.4]
  assign _T_57289 = $signed(buffer_0_610) + $signed(buffer_0_611); // @[Modules.scala 56:109:@3496.4]
  assign _T_57290 = _T_57289[10:0]; // @[Modules.scala 56:109:@3497.4]
  assign buffer_0_697 = $signed(_T_57290); // @[Modules.scala 56:109:@3498.4]
  assign _T_57292 = $signed(buffer_0_612) + $signed(buffer_0_613); // @[Modules.scala 56:109:@3500.4]
  assign _T_57293 = _T_57292[10:0]; // @[Modules.scala 56:109:@3501.4]
  assign buffer_0_698 = $signed(_T_57293); // @[Modules.scala 56:109:@3502.4]
  assign _T_57295 = $signed(buffer_0_614) + $signed(buffer_0_615); // @[Modules.scala 56:109:@3504.4]
  assign _T_57296 = _T_57295[10:0]; // @[Modules.scala 56:109:@3505.4]
  assign buffer_0_699 = $signed(_T_57296); // @[Modules.scala 56:109:@3506.4]
  assign _T_57298 = $signed(buffer_0_616) + $signed(buffer_0_617); // @[Modules.scala 56:109:@3508.4]
  assign _T_57299 = _T_57298[10:0]; // @[Modules.scala 56:109:@3509.4]
  assign buffer_0_700 = $signed(_T_57299); // @[Modules.scala 56:109:@3510.4]
  assign _T_57301 = $signed(buffer_0_618) + $signed(buffer_0_619); // @[Modules.scala 56:109:@3512.4]
  assign _T_57302 = _T_57301[10:0]; // @[Modules.scala 56:109:@3513.4]
  assign buffer_0_701 = $signed(_T_57302); // @[Modules.scala 56:109:@3514.4]
  assign _T_57304 = $signed(buffer_0_620) + $signed(buffer_0_621); // @[Modules.scala 56:109:@3516.4]
  assign _T_57305 = _T_57304[10:0]; // @[Modules.scala 56:109:@3517.4]
  assign buffer_0_702 = $signed(_T_57305); // @[Modules.scala 56:109:@3518.4]
  assign _T_57307 = $signed(buffer_0_622) + $signed(buffer_0_623); // @[Modules.scala 56:109:@3520.4]
  assign _T_57308 = _T_57307[10:0]; // @[Modules.scala 56:109:@3521.4]
  assign buffer_0_703 = $signed(_T_57308); // @[Modules.scala 56:109:@3522.4]
  assign _T_57310 = $signed(buffer_0_624) + $signed(buffer_0_625); // @[Modules.scala 56:109:@3524.4]
  assign _T_57311 = _T_57310[10:0]; // @[Modules.scala 56:109:@3525.4]
  assign buffer_0_704 = $signed(_T_57311); // @[Modules.scala 56:109:@3526.4]
  assign _T_57313 = $signed(buffer_0_626) + $signed(buffer_0_627); // @[Modules.scala 56:109:@3528.4]
  assign _T_57314 = _T_57313[10:0]; // @[Modules.scala 56:109:@3529.4]
  assign buffer_0_705 = $signed(_T_57314); // @[Modules.scala 56:109:@3530.4]
  assign _T_57316 = $signed(buffer_0_628) + $signed(buffer_0_629); // @[Modules.scala 56:109:@3532.4]
  assign _T_57317 = _T_57316[10:0]; // @[Modules.scala 56:109:@3533.4]
  assign buffer_0_706 = $signed(_T_57317); // @[Modules.scala 56:109:@3534.4]
  assign _T_57319 = $signed(buffer_0_630) + $signed(buffer_0_631); // @[Modules.scala 56:109:@3536.4]
  assign _T_57320 = _T_57319[10:0]; // @[Modules.scala 56:109:@3537.4]
  assign buffer_0_707 = $signed(_T_57320); // @[Modules.scala 56:109:@3538.4]
  assign _T_57322 = $signed(buffer_0_632) + $signed(buffer_0_633); // @[Modules.scala 56:109:@3540.4]
  assign _T_57323 = _T_57322[10:0]; // @[Modules.scala 56:109:@3541.4]
  assign buffer_0_708 = $signed(_T_57323); // @[Modules.scala 56:109:@3542.4]
  assign _T_57325 = $signed(buffer_0_634) + $signed(buffer_0_635); // @[Modules.scala 56:109:@3544.4]
  assign _T_57326 = _T_57325[10:0]; // @[Modules.scala 56:109:@3545.4]
  assign buffer_0_709 = $signed(_T_57326); // @[Modules.scala 56:109:@3546.4]
  assign _T_57328 = $signed(buffer_0_636) + $signed(buffer_0_637); // @[Modules.scala 56:109:@3548.4]
  assign _T_57329 = _T_57328[10:0]; // @[Modules.scala 56:109:@3549.4]
  assign buffer_0_710 = $signed(_T_57329); // @[Modules.scala 56:109:@3550.4]
  assign _T_57331 = $signed(buffer_0_638) + $signed(buffer_0_639); // @[Modules.scala 56:109:@3552.4]
  assign _T_57332 = _T_57331[10:0]; // @[Modules.scala 56:109:@3553.4]
  assign buffer_0_711 = $signed(_T_57332); // @[Modules.scala 56:109:@3554.4]
  assign _T_57334 = $signed(buffer_0_640) + $signed(buffer_0_641); // @[Modules.scala 56:109:@3556.4]
  assign _T_57335 = _T_57334[10:0]; // @[Modules.scala 56:109:@3557.4]
  assign buffer_0_712 = $signed(_T_57335); // @[Modules.scala 56:109:@3558.4]
  assign _T_57337 = $signed(buffer_0_642) + $signed(buffer_0_643); // @[Modules.scala 56:109:@3560.4]
  assign _T_57338 = _T_57337[10:0]; // @[Modules.scala 56:109:@3561.4]
  assign buffer_0_713 = $signed(_T_57338); // @[Modules.scala 56:109:@3562.4]
  assign _T_57340 = $signed(buffer_0_644) + $signed(buffer_0_645); // @[Modules.scala 56:109:@3564.4]
  assign _T_57341 = _T_57340[10:0]; // @[Modules.scala 56:109:@3565.4]
  assign buffer_0_714 = $signed(_T_57341); // @[Modules.scala 56:109:@3566.4]
  assign _T_57343 = $signed(buffer_0_646) + $signed(buffer_0_647); // @[Modules.scala 56:109:@3568.4]
  assign _T_57344 = _T_57343[10:0]; // @[Modules.scala 56:109:@3569.4]
  assign buffer_0_715 = $signed(_T_57344); // @[Modules.scala 56:109:@3570.4]
  assign _T_57346 = $signed(buffer_0_648) + $signed(buffer_0_649); // @[Modules.scala 56:109:@3572.4]
  assign _T_57347 = _T_57346[10:0]; // @[Modules.scala 56:109:@3573.4]
  assign buffer_0_716 = $signed(_T_57347); // @[Modules.scala 56:109:@3574.4]
  assign _T_57349 = $signed(buffer_0_650) + $signed(buffer_0_651); // @[Modules.scala 56:109:@3576.4]
  assign _T_57350 = _T_57349[10:0]; // @[Modules.scala 56:109:@3577.4]
  assign buffer_0_717 = $signed(_T_57350); // @[Modules.scala 56:109:@3578.4]
  assign _T_57352 = $signed(buffer_0_652) + $signed(buffer_0_653); // @[Modules.scala 56:109:@3580.4]
  assign _T_57353 = _T_57352[10:0]; // @[Modules.scala 56:109:@3581.4]
  assign buffer_0_718 = $signed(_T_57353); // @[Modules.scala 56:109:@3582.4]
  assign _T_57355 = $signed(buffer_0_654) + $signed(buffer_0_655); // @[Modules.scala 56:109:@3584.4]
  assign _T_57356 = _T_57355[10:0]; // @[Modules.scala 56:109:@3585.4]
  assign buffer_0_719 = $signed(_T_57356); // @[Modules.scala 56:109:@3586.4]
  assign _T_57358 = $signed(buffer_0_656) + $signed(buffer_0_657); // @[Modules.scala 56:109:@3588.4]
  assign _T_57359 = _T_57358[10:0]; // @[Modules.scala 56:109:@3589.4]
  assign buffer_0_720 = $signed(_T_57359); // @[Modules.scala 56:109:@3590.4]
  assign _T_57361 = $signed(buffer_0_658) + $signed(buffer_0_659); // @[Modules.scala 56:109:@3592.4]
  assign _T_57362 = _T_57361[10:0]; // @[Modules.scala 56:109:@3593.4]
  assign buffer_0_721 = $signed(_T_57362); // @[Modules.scala 56:109:@3594.4]
  assign _T_57364 = $signed(buffer_0_660) + $signed(buffer_0_661); // @[Modules.scala 56:109:@3596.4]
  assign _T_57365 = _T_57364[10:0]; // @[Modules.scala 56:109:@3597.4]
  assign buffer_0_722 = $signed(_T_57365); // @[Modules.scala 56:109:@3598.4]
  assign _T_57367 = $signed(buffer_0_662) + $signed(buffer_0_663); // @[Modules.scala 56:109:@3600.4]
  assign _T_57368 = _T_57367[10:0]; // @[Modules.scala 56:109:@3601.4]
  assign buffer_0_723 = $signed(_T_57368); // @[Modules.scala 56:109:@3602.4]
  assign _T_57370 = $signed(buffer_0_664) + $signed(buffer_0_665); // @[Modules.scala 56:109:@3604.4]
  assign _T_57371 = _T_57370[10:0]; // @[Modules.scala 56:109:@3605.4]
  assign buffer_0_724 = $signed(_T_57371); // @[Modules.scala 56:109:@3606.4]
  assign _T_57373 = $signed(buffer_0_666) + $signed(buffer_0_667); // @[Modules.scala 56:109:@3608.4]
  assign _T_57374 = _T_57373[10:0]; // @[Modules.scala 56:109:@3609.4]
  assign buffer_0_725 = $signed(_T_57374); // @[Modules.scala 56:109:@3610.4]
  assign _T_57376 = $signed(buffer_0_668) + $signed(buffer_0_669); // @[Modules.scala 56:109:@3612.4]
  assign _T_57377 = _T_57376[10:0]; // @[Modules.scala 56:109:@3613.4]
  assign buffer_0_726 = $signed(_T_57377); // @[Modules.scala 56:109:@3614.4]
  assign _T_57379 = $signed(buffer_0_670) + $signed(buffer_0_671); // @[Modules.scala 56:109:@3616.4]
  assign _T_57380 = _T_57379[10:0]; // @[Modules.scala 56:109:@3617.4]
  assign buffer_0_727 = $signed(_T_57380); // @[Modules.scala 56:109:@3618.4]
  assign _T_57382 = $signed(buffer_0_672) + $signed(buffer_0_673); // @[Modules.scala 56:109:@3620.4]
  assign _T_57383 = _T_57382[10:0]; // @[Modules.scala 56:109:@3621.4]
  assign buffer_0_728 = $signed(_T_57383); // @[Modules.scala 56:109:@3622.4]
  assign _T_57385 = $signed(buffer_0_674) + $signed(buffer_0_675); // @[Modules.scala 56:109:@3624.4]
  assign _T_57386 = _T_57385[10:0]; // @[Modules.scala 56:109:@3625.4]
  assign buffer_0_729 = $signed(_T_57386); // @[Modules.scala 56:109:@3626.4]
  assign _T_57388 = $signed(buffer_0_676) + $signed(buffer_0_677); // @[Modules.scala 56:109:@3628.4]
  assign _T_57389 = _T_57388[10:0]; // @[Modules.scala 56:109:@3629.4]
  assign buffer_0_730 = $signed(_T_57389); // @[Modules.scala 56:109:@3630.4]
  assign _T_57391 = $signed(buffer_0_678) + $signed(buffer_0_679); // @[Modules.scala 56:109:@3632.4]
  assign _T_57392 = _T_57391[10:0]; // @[Modules.scala 56:109:@3633.4]
  assign buffer_0_731 = $signed(_T_57392); // @[Modules.scala 56:109:@3634.4]
  assign _T_57394 = $signed(buffer_0_680) + $signed(buffer_0_681); // @[Modules.scala 56:109:@3636.4]
  assign _T_57395 = _T_57394[10:0]; // @[Modules.scala 56:109:@3637.4]
  assign buffer_0_732 = $signed(_T_57395); // @[Modules.scala 56:109:@3638.4]
  assign _T_57397 = $signed(buffer_0_682) + $signed(buffer_0_683); // @[Modules.scala 56:109:@3640.4]
  assign _T_57398 = _T_57397[10:0]; // @[Modules.scala 56:109:@3641.4]
  assign buffer_0_733 = $signed(_T_57398); // @[Modules.scala 56:109:@3642.4]
  assign _T_57400 = $signed(buffer_0_684) + $signed(buffer_0_685); // @[Modules.scala 56:109:@3644.4]
  assign _T_57401 = _T_57400[10:0]; // @[Modules.scala 56:109:@3645.4]
  assign buffer_0_734 = $signed(_T_57401); // @[Modules.scala 56:109:@3646.4]
  assign _T_57403 = $signed(buffer_0_686) + $signed(buffer_0_687); // @[Modules.scala 63:156:@3649.4]
  assign _T_57404 = _T_57403[10:0]; // @[Modules.scala 63:156:@3650.4]
  assign buffer_0_736 = $signed(_T_57404); // @[Modules.scala 63:156:@3651.4]
  assign _T_57406 = $signed(buffer_0_736) + $signed(buffer_0_688); // @[Modules.scala 63:156:@3653.4]
  assign _T_57407 = _T_57406[10:0]; // @[Modules.scala 63:156:@3654.4]
  assign buffer_0_737 = $signed(_T_57407); // @[Modules.scala 63:156:@3655.4]
  assign _T_57409 = $signed(buffer_0_737) + $signed(buffer_0_689); // @[Modules.scala 63:156:@3657.4]
  assign _T_57410 = _T_57409[10:0]; // @[Modules.scala 63:156:@3658.4]
  assign buffer_0_738 = $signed(_T_57410); // @[Modules.scala 63:156:@3659.4]
  assign _T_57412 = $signed(buffer_0_738) + $signed(buffer_0_690); // @[Modules.scala 63:156:@3661.4]
  assign _T_57413 = _T_57412[10:0]; // @[Modules.scala 63:156:@3662.4]
  assign buffer_0_739 = $signed(_T_57413); // @[Modules.scala 63:156:@3663.4]
  assign _T_57415 = $signed(buffer_0_739) + $signed(buffer_0_691); // @[Modules.scala 63:156:@3665.4]
  assign _T_57416 = _T_57415[10:0]; // @[Modules.scala 63:156:@3666.4]
  assign buffer_0_740 = $signed(_T_57416); // @[Modules.scala 63:156:@3667.4]
  assign _T_57418 = $signed(buffer_0_740) + $signed(buffer_0_692); // @[Modules.scala 63:156:@3669.4]
  assign _T_57419 = _T_57418[10:0]; // @[Modules.scala 63:156:@3670.4]
  assign buffer_0_741 = $signed(_T_57419); // @[Modules.scala 63:156:@3671.4]
  assign _T_57421 = $signed(buffer_0_741) + $signed(buffer_0_693); // @[Modules.scala 63:156:@3673.4]
  assign _T_57422 = _T_57421[10:0]; // @[Modules.scala 63:156:@3674.4]
  assign buffer_0_742 = $signed(_T_57422); // @[Modules.scala 63:156:@3675.4]
  assign _T_57424 = $signed(buffer_0_742) + $signed(buffer_0_694); // @[Modules.scala 63:156:@3677.4]
  assign _T_57425 = _T_57424[10:0]; // @[Modules.scala 63:156:@3678.4]
  assign buffer_0_743 = $signed(_T_57425); // @[Modules.scala 63:156:@3679.4]
  assign _T_57427 = $signed(buffer_0_743) + $signed(buffer_0_695); // @[Modules.scala 63:156:@3681.4]
  assign _T_57428 = _T_57427[10:0]; // @[Modules.scala 63:156:@3682.4]
  assign buffer_0_744 = $signed(_T_57428); // @[Modules.scala 63:156:@3683.4]
  assign _T_57430 = $signed(buffer_0_744) + $signed(buffer_0_696); // @[Modules.scala 63:156:@3685.4]
  assign _T_57431 = _T_57430[10:0]; // @[Modules.scala 63:156:@3686.4]
  assign buffer_0_745 = $signed(_T_57431); // @[Modules.scala 63:156:@3687.4]
  assign _T_57433 = $signed(buffer_0_745) + $signed(buffer_0_697); // @[Modules.scala 63:156:@3689.4]
  assign _T_57434 = _T_57433[10:0]; // @[Modules.scala 63:156:@3690.4]
  assign buffer_0_746 = $signed(_T_57434); // @[Modules.scala 63:156:@3691.4]
  assign _T_57436 = $signed(buffer_0_746) + $signed(buffer_0_698); // @[Modules.scala 63:156:@3693.4]
  assign _T_57437 = _T_57436[10:0]; // @[Modules.scala 63:156:@3694.4]
  assign buffer_0_747 = $signed(_T_57437); // @[Modules.scala 63:156:@3695.4]
  assign _T_57439 = $signed(buffer_0_747) + $signed(buffer_0_699); // @[Modules.scala 63:156:@3697.4]
  assign _T_57440 = _T_57439[10:0]; // @[Modules.scala 63:156:@3698.4]
  assign buffer_0_748 = $signed(_T_57440); // @[Modules.scala 63:156:@3699.4]
  assign _T_57442 = $signed(buffer_0_748) + $signed(buffer_0_700); // @[Modules.scala 63:156:@3701.4]
  assign _T_57443 = _T_57442[10:0]; // @[Modules.scala 63:156:@3702.4]
  assign buffer_0_749 = $signed(_T_57443); // @[Modules.scala 63:156:@3703.4]
  assign _T_57445 = $signed(buffer_0_749) + $signed(buffer_0_701); // @[Modules.scala 63:156:@3705.4]
  assign _T_57446 = _T_57445[10:0]; // @[Modules.scala 63:156:@3706.4]
  assign buffer_0_750 = $signed(_T_57446); // @[Modules.scala 63:156:@3707.4]
  assign _T_57448 = $signed(buffer_0_750) + $signed(buffer_0_702); // @[Modules.scala 63:156:@3709.4]
  assign _T_57449 = _T_57448[10:0]; // @[Modules.scala 63:156:@3710.4]
  assign buffer_0_751 = $signed(_T_57449); // @[Modules.scala 63:156:@3711.4]
  assign _T_57451 = $signed(buffer_0_751) + $signed(buffer_0_703); // @[Modules.scala 63:156:@3713.4]
  assign _T_57452 = _T_57451[10:0]; // @[Modules.scala 63:156:@3714.4]
  assign buffer_0_752 = $signed(_T_57452); // @[Modules.scala 63:156:@3715.4]
  assign _T_57454 = $signed(buffer_0_752) + $signed(buffer_0_704); // @[Modules.scala 63:156:@3717.4]
  assign _T_57455 = _T_57454[10:0]; // @[Modules.scala 63:156:@3718.4]
  assign buffer_0_753 = $signed(_T_57455); // @[Modules.scala 63:156:@3719.4]
  assign _T_57457 = $signed(buffer_0_753) + $signed(buffer_0_705); // @[Modules.scala 63:156:@3721.4]
  assign _T_57458 = _T_57457[10:0]; // @[Modules.scala 63:156:@3722.4]
  assign buffer_0_754 = $signed(_T_57458); // @[Modules.scala 63:156:@3723.4]
  assign _T_57460 = $signed(buffer_0_754) + $signed(buffer_0_706); // @[Modules.scala 63:156:@3725.4]
  assign _T_57461 = _T_57460[10:0]; // @[Modules.scala 63:156:@3726.4]
  assign buffer_0_755 = $signed(_T_57461); // @[Modules.scala 63:156:@3727.4]
  assign _T_57463 = $signed(buffer_0_755) + $signed(buffer_0_707); // @[Modules.scala 63:156:@3729.4]
  assign _T_57464 = _T_57463[10:0]; // @[Modules.scala 63:156:@3730.4]
  assign buffer_0_756 = $signed(_T_57464); // @[Modules.scala 63:156:@3731.4]
  assign _T_57466 = $signed(buffer_0_756) + $signed(buffer_0_708); // @[Modules.scala 63:156:@3733.4]
  assign _T_57467 = _T_57466[10:0]; // @[Modules.scala 63:156:@3734.4]
  assign buffer_0_757 = $signed(_T_57467); // @[Modules.scala 63:156:@3735.4]
  assign _T_57469 = $signed(buffer_0_757) + $signed(buffer_0_709); // @[Modules.scala 63:156:@3737.4]
  assign _T_57470 = _T_57469[10:0]; // @[Modules.scala 63:156:@3738.4]
  assign buffer_0_758 = $signed(_T_57470); // @[Modules.scala 63:156:@3739.4]
  assign _T_57472 = $signed(buffer_0_758) + $signed(buffer_0_710); // @[Modules.scala 63:156:@3741.4]
  assign _T_57473 = _T_57472[10:0]; // @[Modules.scala 63:156:@3742.4]
  assign buffer_0_759 = $signed(_T_57473); // @[Modules.scala 63:156:@3743.4]
  assign _T_57475 = $signed(buffer_0_759) + $signed(buffer_0_711); // @[Modules.scala 63:156:@3745.4]
  assign _T_57476 = _T_57475[10:0]; // @[Modules.scala 63:156:@3746.4]
  assign buffer_0_760 = $signed(_T_57476); // @[Modules.scala 63:156:@3747.4]
  assign _T_57478 = $signed(buffer_0_760) + $signed(buffer_0_712); // @[Modules.scala 63:156:@3749.4]
  assign _T_57479 = _T_57478[10:0]; // @[Modules.scala 63:156:@3750.4]
  assign buffer_0_761 = $signed(_T_57479); // @[Modules.scala 63:156:@3751.4]
  assign _T_57481 = $signed(buffer_0_761) + $signed(buffer_0_713); // @[Modules.scala 63:156:@3753.4]
  assign _T_57482 = _T_57481[10:0]; // @[Modules.scala 63:156:@3754.4]
  assign buffer_0_762 = $signed(_T_57482); // @[Modules.scala 63:156:@3755.4]
  assign _T_57484 = $signed(buffer_0_762) + $signed(buffer_0_714); // @[Modules.scala 63:156:@3757.4]
  assign _T_57485 = _T_57484[10:0]; // @[Modules.scala 63:156:@3758.4]
  assign buffer_0_763 = $signed(_T_57485); // @[Modules.scala 63:156:@3759.4]
  assign _T_57487 = $signed(buffer_0_763) + $signed(buffer_0_715); // @[Modules.scala 63:156:@3761.4]
  assign _T_57488 = _T_57487[10:0]; // @[Modules.scala 63:156:@3762.4]
  assign buffer_0_764 = $signed(_T_57488); // @[Modules.scala 63:156:@3763.4]
  assign _T_57490 = $signed(buffer_0_764) + $signed(buffer_0_716); // @[Modules.scala 63:156:@3765.4]
  assign _T_57491 = _T_57490[10:0]; // @[Modules.scala 63:156:@3766.4]
  assign buffer_0_765 = $signed(_T_57491); // @[Modules.scala 63:156:@3767.4]
  assign _T_57493 = $signed(buffer_0_765) + $signed(buffer_0_717); // @[Modules.scala 63:156:@3769.4]
  assign _T_57494 = _T_57493[10:0]; // @[Modules.scala 63:156:@3770.4]
  assign buffer_0_766 = $signed(_T_57494); // @[Modules.scala 63:156:@3771.4]
  assign _T_57496 = $signed(buffer_0_766) + $signed(buffer_0_718); // @[Modules.scala 63:156:@3773.4]
  assign _T_57497 = _T_57496[10:0]; // @[Modules.scala 63:156:@3774.4]
  assign buffer_0_767 = $signed(_T_57497); // @[Modules.scala 63:156:@3775.4]
  assign _T_57499 = $signed(buffer_0_767) + $signed(buffer_0_719); // @[Modules.scala 63:156:@3777.4]
  assign _T_57500 = _T_57499[10:0]; // @[Modules.scala 63:156:@3778.4]
  assign buffer_0_768 = $signed(_T_57500); // @[Modules.scala 63:156:@3779.4]
  assign _T_57502 = $signed(buffer_0_768) + $signed(buffer_0_720); // @[Modules.scala 63:156:@3781.4]
  assign _T_57503 = _T_57502[10:0]; // @[Modules.scala 63:156:@3782.4]
  assign buffer_0_769 = $signed(_T_57503); // @[Modules.scala 63:156:@3783.4]
  assign _T_57505 = $signed(buffer_0_769) + $signed(buffer_0_721); // @[Modules.scala 63:156:@3785.4]
  assign _T_57506 = _T_57505[10:0]; // @[Modules.scala 63:156:@3786.4]
  assign buffer_0_770 = $signed(_T_57506); // @[Modules.scala 63:156:@3787.4]
  assign _T_57508 = $signed(buffer_0_770) + $signed(buffer_0_722); // @[Modules.scala 63:156:@3789.4]
  assign _T_57509 = _T_57508[10:0]; // @[Modules.scala 63:156:@3790.4]
  assign buffer_0_771 = $signed(_T_57509); // @[Modules.scala 63:156:@3791.4]
  assign _T_57511 = $signed(buffer_0_771) + $signed(buffer_0_723); // @[Modules.scala 63:156:@3793.4]
  assign _T_57512 = _T_57511[10:0]; // @[Modules.scala 63:156:@3794.4]
  assign buffer_0_772 = $signed(_T_57512); // @[Modules.scala 63:156:@3795.4]
  assign _T_57514 = $signed(buffer_0_772) + $signed(buffer_0_724); // @[Modules.scala 63:156:@3797.4]
  assign _T_57515 = _T_57514[10:0]; // @[Modules.scala 63:156:@3798.4]
  assign buffer_0_773 = $signed(_T_57515); // @[Modules.scala 63:156:@3799.4]
  assign _T_57517 = $signed(buffer_0_773) + $signed(buffer_0_725); // @[Modules.scala 63:156:@3801.4]
  assign _T_57518 = _T_57517[10:0]; // @[Modules.scala 63:156:@3802.4]
  assign buffer_0_774 = $signed(_T_57518); // @[Modules.scala 63:156:@3803.4]
  assign _T_57520 = $signed(buffer_0_774) + $signed(buffer_0_726); // @[Modules.scala 63:156:@3805.4]
  assign _T_57521 = _T_57520[10:0]; // @[Modules.scala 63:156:@3806.4]
  assign buffer_0_775 = $signed(_T_57521); // @[Modules.scala 63:156:@3807.4]
  assign _T_57523 = $signed(buffer_0_775) + $signed(buffer_0_727); // @[Modules.scala 63:156:@3809.4]
  assign _T_57524 = _T_57523[10:0]; // @[Modules.scala 63:156:@3810.4]
  assign buffer_0_776 = $signed(_T_57524); // @[Modules.scala 63:156:@3811.4]
  assign _T_57526 = $signed(buffer_0_776) + $signed(buffer_0_728); // @[Modules.scala 63:156:@3813.4]
  assign _T_57527 = _T_57526[10:0]; // @[Modules.scala 63:156:@3814.4]
  assign buffer_0_777 = $signed(_T_57527); // @[Modules.scala 63:156:@3815.4]
  assign _T_57529 = $signed(buffer_0_777) + $signed(buffer_0_729); // @[Modules.scala 63:156:@3817.4]
  assign _T_57530 = _T_57529[10:0]; // @[Modules.scala 63:156:@3818.4]
  assign buffer_0_778 = $signed(_T_57530); // @[Modules.scala 63:156:@3819.4]
  assign _T_57532 = $signed(buffer_0_778) + $signed(buffer_0_730); // @[Modules.scala 63:156:@3821.4]
  assign _T_57533 = _T_57532[10:0]; // @[Modules.scala 63:156:@3822.4]
  assign buffer_0_779 = $signed(_T_57533); // @[Modules.scala 63:156:@3823.4]
  assign _T_57535 = $signed(buffer_0_779) + $signed(buffer_0_731); // @[Modules.scala 63:156:@3825.4]
  assign _T_57536 = _T_57535[10:0]; // @[Modules.scala 63:156:@3826.4]
  assign buffer_0_780 = $signed(_T_57536); // @[Modules.scala 63:156:@3827.4]
  assign _T_57538 = $signed(buffer_0_780) + $signed(buffer_0_732); // @[Modules.scala 63:156:@3829.4]
  assign _T_57539 = _T_57538[10:0]; // @[Modules.scala 63:156:@3830.4]
  assign buffer_0_781 = $signed(_T_57539); // @[Modules.scala 63:156:@3831.4]
  assign _T_57541 = $signed(buffer_0_781) + $signed(buffer_0_733); // @[Modules.scala 63:156:@3833.4]
  assign _T_57542 = _T_57541[10:0]; // @[Modules.scala 63:156:@3834.4]
  assign buffer_0_782 = $signed(_T_57542); // @[Modules.scala 63:156:@3835.4]
  assign _T_57544 = $signed(buffer_0_782) + $signed(buffer_0_734); // @[Modules.scala 63:156:@3837.4]
  assign _T_57545 = _T_57544[10:0]; // @[Modules.scala 63:156:@3838.4]
  assign buffer_0_783 = $signed(_T_57545); // @[Modules.scala 63:156:@3839.4]
  assign _T_57551 = $signed(_T_54269) - $signed(io_in_1); // @[Modules.scala 46:47:@3845.4]
  assign _T_57552 = _T_57551[4:0]; // @[Modules.scala 46:47:@3846.4]
  assign _T_57553 = $signed(_T_57552); // @[Modules.scala 46:47:@3847.4]
  assign _T_57561 = $signed(io_in_4) + $signed(io_in_5); // @[Modules.scala 37:46:@3856.4]
  assign _T_57562 = _T_57561[4:0]; // @[Modules.scala 37:46:@3857.4]
  assign _T_57563 = $signed(_T_57562); // @[Modules.scala 37:46:@3858.4]
  assign _T_57564 = $signed(io_in_6) + $signed(io_in_7); // @[Modules.scala 37:46:@3860.4]
  assign _T_57565 = _T_57564[4:0]; // @[Modules.scala 37:46:@3861.4]
  assign _T_57566 = $signed(_T_57565); // @[Modules.scala 37:46:@3862.4]
  assign _T_57567 = $signed(io_in_8) + $signed(io_in_9); // @[Modules.scala 37:46:@3864.4]
  assign _T_57568 = _T_57567[4:0]; // @[Modules.scala 37:46:@3865.4]
  assign _T_57569 = $signed(_T_57568); // @[Modules.scala 37:46:@3866.4]
  assign _T_57577 = $signed(io_in_12) + $signed(io_in_13); // @[Modules.scala 37:46:@3875.4]
  assign _T_57578 = _T_57577[4:0]; // @[Modules.scala 37:46:@3876.4]
  assign _T_57579 = $signed(_T_57578); // @[Modules.scala 37:46:@3877.4]
  assign _T_57580 = $signed(io_in_14) + $signed(io_in_15); // @[Modules.scala 37:46:@3879.4]
  assign _T_57581 = _T_57580[4:0]; // @[Modules.scala 37:46:@3880.4]
  assign _T_57582 = $signed(_T_57581); // @[Modules.scala 37:46:@3881.4]
  assign _T_57583 = $signed(io_in_16) - $signed(io_in_17); // @[Modules.scala 40:46:@3883.4]
  assign _T_57584 = _T_57583[4:0]; // @[Modules.scala 40:46:@3884.4]
  assign _T_57585 = $signed(_T_57584); // @[Modules.scala 40:46:@3885.4]
  assign _T_57586 = $signed(io_in_18) - $signed(io_in_19); // @[Modules.scala 40:46:@3887.4]
  assign _T_57587 = _T_57586[4:0]; // @[Modules.scala 40:46:@3888.4]
  assign _T_57588 = $signed(_T_57587); // @[Modules.scala 40:46:@3889.4]
  assign _T_57592 = $signed(io_in_22) - $signed(io_in_23); // @[Modules.scala 40:46:@3895.4]
  assign _T_57593 = _T_57592[4:0]; // @[Modules.scala 40:46:@3896.4]
  assign _T_57594 = $signed(_T_57593); // @[Modules.scala 40:46:@3897.4]
  assign _T_57595 = $signed(io_in_24) + $signed(io_in_25); // @[Modules.scala 37:46:@3899.4]
  assign _T_57596 = _T_57595[4:0]; // @[Modules.scala 37:46:@3900.4]
  assign _T_57597 = $signed(_T_57596); // @[Modules.scala 37:46:@3901.4]
  assign _T_57599 = $signed(5'sh0) - $signed(io_in_26); // @[Modules.scala 46:37:@3903.4]
  assign _T_57600 = _T_57599[4:0]; // @[Modules.scala 46:37:@3904.4]
  assign _T_57601 = $signed(_T_57600); // @[Modules.scala 46:37:@3905.4]
  assign _T_57602 = $signed(_T_57601) - $signed(io_in_27); // @[Modules.scala 46:47:@3906.4]
  assign _T_57603 = _T_57602[4:0]; // @[Modules.scala 46:47:@3907.4]
  assign _T_57604 = $signed(_T_57603); // @[Modules.scala 46:47:@3908.4]
  assign _T_57605 = $signed(io_in_28) - $signed(io_in_29); // @[Modules.scala 40:46:@3910.4]
  assign _T_57606 = _T_57605[4:0]; // @[Modules.scala 40:46:@3911.4]
  assign _T_57607 = $signed(_T_57606); // @[Modules.scala 40:46:@3912.4]
  assign _T_57608 = $signed(io_in_30) + $signed(io_in_31); // @[Modules.scala 37:46:@3914.4]
  assign _T_57609 = _T_57608[4:0]; // @[Modules.scala 37:46:@3915.4]
  assign _T_57610 = $signed(_T_57609); // @[Modules.scala 37:46:@3916.4]
  assign _T_57614 = $signed(io_in_34) + $signed(io_in_35); // @[Modules.scala 37:46:@3922.4]
  assign _T_57615 = _T_57614[4:0]; // @[Modules.scala 37:46:@3923.4]
  assign _T_57616 = $signed(_T_57615); // @[Modules.scala 37:46:@3924.4]
  assign _T_57617 = $signed(io_in_36) + $signed(io_in_37); // @[Modules.scala 37:46:@3926.4]
  assign _T_57618 = _T_57617[4:0]; // @[Modules.scala 37:46:@3927.4]
  assign _T_57619 = $signed(_T_57618); // @[Modules.scala 37:46:@3928.4]
  assign _T_57620 = $signed(io_in_38) + $signed(io_in_39); // @[Modules.scala 37:46:@3930.4]
  assign _T_57621 = _T_57620[4:0]; // @[Modules.scala 37:46:@3931.4]
  assign _T_57622 = $signed(_T_57621); // @[Modules.scala 37:46:@3932.4]
  assign _T_57623 = $signed(io_in_40) + $signed(io_in_41); // @[Modules.scala 37:46:@3934.4]
  assign _T_57624 = _T_57623[4:0]; // @[Modules.scala 37:46:@3935.4]
  assign _T_57625 = $signed(_T_57624); // @[Modules.scala 37:46:@3936.4]
  assign _T_57626 = $signed(io_in_42) + $signed(io_in_43); // @[Modules.scala 37:46:@3938.4]
  assign _T_57627 = _T_57626[4:0]; // @[Modules.scala 37:46:@3939.4]
  assign _T_57628 = $signed(_T_57627); // @[Modules.scala 37:46:@3940.4]
  assign _T_57633 = $signed(_T_54407) + $signed(io_in_45); // @[Modules.scala 43:47:@3945.4]
  assign _T_57634 = _T_57633[4:0]; // @[Modules.scala 43:47:@3946.4]
  assign _T_57635 = $signed(_T_57634); // @[Modules.scala 43:47:@3947.4]
  assign _T_57636 = $signed(io_in_46) + $signed(io_in_47); // @[Modules.scala 37:46:@3949.4]
  assign _T_57637 = _T_57636[4:0]; // @[Modules.scala 37:46:@3950.4]
  assign _T_57638 = $signed(_T_57637); // @[Modules.scala 37:46:@3951.4]
  assign _T_57639 = $signed(io_in_48) + $signed(io_in_49); // @[Modules.scala 37:46:@3953.4]
  assign _T_57640 = _T_57639[4:0]; // @[Modules.scala 37:46:@3954.4]
  assign _T_57641 = $signed(_T_57640); // @[Modules.scala 37:46:@3955.4]
  assign _T_57642 = $signed(io_in_50) + $signed(io_in_51); // @[Modules.scala 37:46:@3957.4]
  assign _T_57643 = _T_57642[4:0]; // @[Modules.scala 37:46:@3958.4]
  assign _T_57644 = $signed(_T_57643); // @[Modules.scala 37:46:@3959.4]
  assign _T_57645 = $signed(io_in_52) - $signed(io_in_53); // @[Modules.scala 40:46:@3961.4]
  assign _T_57646 = _T_57645[4:0]; // @[Modules.scala 40:46:@3962.4]
  assign _T_57647 = $signed(_T_57646); // @[Modules.scala 40:46:@3963.4]
  assign _T_57649 = $signed(5'sh0) - $signed(io_in_54); // @[Modules.scala 43:37:@3965.4]
  assign _T_57650 = _T_57649[4:0]; // @[Modules.scala 43:37:@3966.4]
  assign _T_57651 = $signed(_T_57650); // @[Modules.scala 43:37:@3967.4]
  assign _T_57652 = $signed(_T_57651) + $signed(io_in_55); // @[Modules.scala 43:47:@3968.4]
  assign _T_57653 = _T_57652[4:0]; // @[Modules.scala 43:47:@3969.4]
  assign _T_57654 = $signed(_T_57653); // @[Modules.scala 43:47:@3970.4]
  assign _T_57656 = $signed(5'sh0) - $signed(io_in_56); // @[Modules.scala 43:37:@3972.4]
  assign _T_57657 = _T_57656[4:0]; // @[Modules.scala 43:37:@3973.4]
  assign _T_57658 = $signed(_T_57657); // @[Modules.scala 43:37:@3974.4]
  assign _T_57659 = $signed(_T_57658) + $signed(io_in_57); // @[Modules.scala 43:47:@3975.4]
  assign _T_57660 = _T_57659[4:0]; // @[Modules.scala 43:47:@3976.4]
  assign _T_57661 = $signed(_T_57660); // @[Modules.scala 43:47:@3977.4]
  assign _T_57662 = $signed(io_in_58) + $signed(io_in_59); // @[Modules.scala 37:46:@3979.4]
  assign _T_57663 = _T_57662[4:0]; // @[Modules.scala 37:46:@3980.4]
  assign _T_57664 = $signed(_T_57663); // @[Modules.scala 37:46:@3981.4]
  assign _T_57665 = $signed(io_in_60) + $signed(io_in_61); // @[Modules.scala 37:46:@3983.4]
  assign _T_57666 = _T_57665[4:0]; // @[Modules.scala 37:46:@3984.4]
  assign _T_57667 = $signed(_T_57666); // @[Modules.scala 37:46:@3985.4]
  assign _T_57668 = $signed(io_in_62) + $signed(io_in_63); // @[Modules.scala 37:46:@3987.4]
  assign _T_57669 = _T_57668[4:0]; // @[Modules.scala 37:46:@3988.4]
  assign _T_57670 = $signed(_T_57669); // @[Modules.scala 37:46:@3989.4]
  assign _T_57671 = $signed(io_in_64) + $signed(io_in_65); // @[Modules.scala 37:46:@3991.4]
  assign _T_57672 = _T_57671[4:0]; // @[Modules.scala 37:46:@3992.4]
  assign _T_57673 = $signed(_T_57672); // @[Modules.scala 37:46:@3993.4]
  assign _T_57674 = $signed(io_in_66) + $signed(io_in_67); // @[Modules.scala 37:46:@3995.4]
  assign _T_57675 = _T_57674[4:0]; // @[Modules.scala 37:46:@3996.4]
  assign _T_57676 = $signed(_T_57675); // @[Modules.scala 37:46:@3997.4]
  assign _T_57677 = $signed(io_in_68) + $signed(io_in_69); // @[Modules.scala 37:46:@3999.4]
  assign _T_57678 = _T_57677[4:0]; // @[Modules.scala 37:46:@4000.4]
  assign _T_57679 = $signed(_T_57678); // @[Modules.scala 37:46:@4001.4]
  assign _T_57680 = $signed(io_in_70) + $signed(io_in_71); // @[Modules.scala 37:46:@4003.4]
  assign _T_57681 = _T_57680[4:0]; // @[Modules.scala 37:46:@4004.4]
  assign _T_57682 = $signed(_T_57681); // @[Modules.scala 37:46:@4005.4]
  assign _T_57683 = $signed(io_in_72) + $signed(io_in_73); // @[Modules.scala 37:46:@4007.4]
  assign _T_57684 = _T_57683[4:0]; // @[Modules.scala 37:46:@4008.4]
  assign _T_57685 = $signed(_T_57684); // @[Modules.scala 37:46:@4009.4]
  assign _T_57686 = $signed(io_in_74) + $signed(io_in_75); // @[Modules.scala 37:46:@4011.4]
  assign _T_57687 = _T_57686[4:0]; // @[Modules.scala 37:46:@4012.4]
  assign _T_57688 = $signed(_T_57687); // @[Modules.scala 37:46:@4013.4]
  assign _T_57689 = $signed(io_in_76) + $signed(io_in_77); // @[Modules.scala 37:46:@4015.4]
  assign _T_57690 = _T_57689[4:0]; // @[Modules.scala 37:46:@4016.4]
  assign _T_57691 = $signed(_T_57690); // @[Modules.scala 37:46:@4017.4]
  assign _T_57695 = $signed(io_in_80) + $signed(io_in_81); // @[Modules.scala 37:46:@4023.4]
  assign _T_57696 = _T_57695[4:0]; // @[Modules.scala 37:46:@4024.4]
  assign _T_57697 = $signed(_T_57696); // @[Modules.scala 37:46:@4025.4]
  assign _T_57699 = $signed(5'sh0) - $signed(io_in_82); // @[Modules.scala 46:37:@4027.4]
  assign _T_57700 = _T_57699[4:0]; // @[Modules.scala 46:37:@4028.4]
  assign _T_57701 = $signed(_T_57700); // @[Modules.scala 46:37:@4029.4]
  assign _T_57702 = $signed(_T_57701) - $signed(io_in_83); // @[Modules.scala 46:47:@4030.4]
  assign _T_57703 = _T_57702[4:0]; // @[Modules.scala 46:47:@4031.4]
  assign _T_57704 = $signed(_T_57703); // @[Modules.scala 46:47:@4032.4]
  assign _T_57706 = $signed(5'sh0) - $signed(io_in_84); // @[Modules.scala 43:37:@4034.4]
  assign _T_57707 = _T_57706[4:0]; // @[Modules.scala 43:37:@4035.4]
  assign _T_57708 = $signed(_T_57707); // @[Modules.scala 43:37:@4036.4]
  assign _T_57709 = $signed(_T_57708) + $signed(io_in_85); // @[Modules.scala 43:47:@4037.4]
  assign _T_57710 = _T_57709[4:0]; // @[Modules.scala 43:47:@4038.4]
  assign _T_57711 = $signed(_T_57710); // @[Modules.scala 43:47:@4039.4]
  assign _T_57716 = $signed(_T_54526) + $signed(io_in_87); // @[Modules.scala 43:47:@4044.4]
  assign _T_57717 = _T_57716[4:0]; // @[Modules.scala 43:47:@4045.4]
  assign _T_57718 = $signed(_T_57717); // @[Modules.scala 43:47:@4046.4]
  assign _T_57725 = $signed(io_in_92) + $signed(io_in_93); // @[Modules.scala 37:46:@4056.4]
  assign _T_57726 = _T_57725[4:0]; // @[Modules.scala 37:46:@4057.4]
  assign _T_57727 = $signed(_T_57726); // @[Modules.scala 37:46:@4058.4]
  assign _T_57731 = $signed(io_in_96) + $signed(io_in_97); // @[Modules.scala 37:46:@4064.4]
  assign _T_57732 = _T_57731[4:0]; // @[Modules.scala 37:46:@4065.4]
  assign _T_57733 = $signed(_T_57732); // @[Modules.scala 37:46:@4066.4]
  assign _T_57749 = $signed(io_in_108) + $signed(io_in_109); // @[Modules.scala 37:46:@4088.4]
  assign _T_57750 = _T_57749[4:0]; // @[Modules.scala 37:46:@4089.4]
  assign _T_57751 = $signed(_T_57750); // @[Modules.scala 37:46:@4090.4]
  assign _T_57759 = $signed(_T_54577) - $signed(io_in_113); // @[Modules.scala 46:47:@4099.4]
  assign _T_57760 = _T_57759[4:0]; // @[Modules.scala 46:47:@4100.4]
  assign _T_57761 = $signed(_T_57760); // @[Modules.scala 46:47:@4101.4]
  assign _T_57766 = $signed(_T_54584) + $signed(io_in_115); // @[Modules.scala 43:47:@4106.4]
  assign _T_57767 = _T_57766[4:0]; // @[Modules.scala 43:47:@4107.4]
  assign _T_57768 = $signed(_T_57767); // @[Modules.scala 43:47:@4108.4]
  assign _T_57773 = $signed(5'sh0) - $signed(io_in_118); // @[Modules.scala 46:37:@4114.4]
  assign _T_57774 = _T_57773[4:0]; // @[Modules.scala 46:37:@4115.4]
  assign _T_57775 = $signed(_T_57774); // @[Modules.scala 46:37:@4116.4]
  assign _T_57776 = $signed(_T_57775) - $signed(io_in_119); // @[Modules.scala 46:47:@4117.4]
  assign _T_57777 = _T_57776[4:0]; // @[Modules.scala 46:47:@4118.4]
  assign _T_57778 = $signed(_T_57777); // @[Modules.scala 46:47:@4119.4]
  assign _T_57804 = $signed(_T_54618) + $signed(io_in_127); // @[Modules.scala 43:47:@4145.4]
  assign _T_57805 = _T_57804[4:0]; // @[Modules.scala 43:47:@4146.4]
  assign _T_57806 = $signed(_T_57805); // @[Modules.scala 43:47:@4147.4]
  assign _T_57807 = $signed(io_in_128) + $signed(io_in_129); // @[Modules.scala 37:46:@4149.4]
  assign _T_57808 = _T_57807[4:0]; // @[Modules.scala 37:46:@4150.4]
  assign _T_57809 = $signed(_T_57808); // @[Modules.scala 37:46:@4151.4]
  assign _T_57810 = $signed(io_in_130) + $signed(io_in_131); // @[Modules.scala 37:46:@4153.4]
  assign _T_57811 = _T_57810[4:0]; // @[Modules.scala 37:46:@4154.4]
  assign _T_57812 = $signed(_T_57811); // @[Modules.scala 37:46:@4155.4]
  assign _T_57814 = $signed(5'sh0) - $signed(io_in_132); // @[Modules.scala 43:37:@4157.4]
  assign _T_57815 = _T_57814[4:0]; // @[Modules.scala 43:37:@4158.4]
  assign _T_57816 = $signed(_T_57815); // @[Modules.scala 43:37:@4159.4]
  assign _T_57817 = $signed(_T_57816) + $signed(io_in_133); // @[Modules.scala 43:47:@4160.4]
  assign _T_57818 = _T_57817[4:0]; // @[Modules.scala 43:47:@4161.4]
  assign _T_57819 = $signed(_T_57818); // @[Modules.scala 43:47:@4162.4]
  assign _T_57823 = $signed(io_in_136) + $signed(io_in_137); // @[Modules.scala 37:46:@4168.4]
  assign _T_57824 = _T_57823[4:0]; // @[Modules.scala 37:46:@4169.4]
  assign _T_57825 = $signed(_T_57824); // @[Modules.scala 37:46:@4170.4]
  assign _T_57830 = $signed(_T_54648) + $signed(io_in_139); // @[Modules.scala 43:47:@4175.4]
  assign _T_57831 = _T_57830[4:0]; // @[Modules.scala 43:47:@4176.4]
  assign _T_57832 = $signed(_T_57831); // @[Modules.scala 43:47:@4177.4]
  assign _T_57833 = $signed(io_in_140) - $signed(io_in_141); // @[Modules.scala 40:46:@4179.4]
  assign _T_57834 = _T_57833[4:0]; // @[Modules.scala 40:46:@4180.4]
  assign _T_57835 = $signed(_T_57834); // @[Modules.scala 40:46:@4181.4]
  assign _T_57840 = $signed(_T_54658) + $signed(io_in_143); // @[Modules.scala 43:47:@4186.4]
  assign _T_57841 = _T_57840[4:0]; // @[Modules.scala 43:47:@4187.4]
  assign _T_57842 = $signed(_T_57841); // @[Modules.scala 43:47:@4188.4]
  assign _T_57844 = $signed(5'sh0) - $signed(io_in_144); // @[Modules.scala 46:37:@4190.4]
  assign _T_57845 = _T_57844[4:0]; // @[Modules.scala 46:37:@4191.4]
  assign _T_57846 = $signed(_T_57845); // @[Modules.scala 46:37:@4192.4]
  assign _T_57847 = $signed(_T_57846) - $signed(io_in_145); // @[Modules.scala 46:47:@4193.4]
  assign _T_57848 = _T_57847[4:0]; // @[Modules.scala 46:47:@4194.4]
  assign _T_57849 = $signed(_T_57848); // @[Modules.scala 46:47:@4195.4]
  assign _T_57851 = $signed(5'sh0) - $signed(io_in_146); // @[Modules.scala 46:37:@4197.4]
  assign _T_57852 = _T_57851[4:0]; // @[Modules.scala 46:37:@4198.4]
  assign _T_57853 = $signed(_T_57852); // @[Modules.scala 46:37:@4199.4]
  assign _T_57854 = $signed(_T_57853) - $signed(io_in_147); // @[Modules.scala 46:47:@4200.4]
  assign _T_57855 = _T_57854[4:0]; // @[Modules.scala 46:47:@4201.4]
  assign _T_57856 = $signed(_T_57855); // @[Modules.scala 46:47:@4202.4]
  assign _T_57857 = $signed(io_in_148) - $signed(io_in_149); // @[Modules.scala 40:46:@4204.4]
  assign _T_57858 = _T_57857[4:0]; // @[Modules.scala 40:46:@4205.4]
  assign _T_57859 = $signed(_T_57858); // @[Modules.scala 40:46:@4206.4]
  assign _T_57860 = $signed(io_in_150) - $signed(io_in_151); // @[Modules.scala 40:46:@4208.4]
  assign _T_57861 = _T_57860[4:0]; // @[Modules.scala 40:46:@4209.4]
  assign _T_57862 = $signed(_T_57861); // @[Modules.scala 40:46:@4210.4]
  assign _T_57877 = $signed(io_in_156) - $signed(io_in_157); // @[Modules.scala 40:46:@4226.4]
  assign _T_57878 = _T_57877[4:0]; // @[Modules.scala 40:46:@4227.4]
  assign _T_57879 = $signed(_T_57878); // @[Modules.scala 40:46:@4228.4]
  assign _T_57895 = $signed(5'sh0) - $signed(io_in_162); // @[Modules.scala 43:37:@4244.4]
  assign _T_57896 = _T_57895[4:0]; // @[Modules.scala 43:37:@4245.4]
  assign _T_57897 = $signed(_T_57896); // @[Modules.scala 43:37:@4246.4]
  assign _T_57898 = $signed(_T_57897) + $signed(io_in_163); // @[Modules.scala 43:47:@4247.4]
  assign _T_57899 = _T_57898[4:0]; // @[Modules.scala 43:47:@4248.4]
  assign _T_57900 = $signed(_T_57899); // @[Modules.scala 43:47:@4249.4]
  assign _T_57902 = $signed(5'sh0) - $signed(io_in_164); // @[Modules.scala 46:37:@4251.4]
  assign _T_57903 = _T_57902[4:0]; // @[Modules.scala 46:37:@4252.4]
  assign _T_57904 = $signed(_T_57903); // @[Modules.scala 46:37:@4253.4]
  assign _T_57905 = $signed(_T_57904) - $signed(io_in_165); // @[Modules.scala 46:47:@4254.4]
  assign _T_57906 = _T_57905[4:0]; // @[Modules.scala 46:47:@4255.4]
  assign _T_57907 = $signed(_T_57906); // @[Modules.scala 46:47:@4256.4]
  assign _T_57908 = $signed(io_in_166) + $signed(io_in_167); // @[Modules.scala 37:46:@4258.4]
  assign _T_57909 = _T_57908[4:0]; // @[Modules.scala 37:46:@4259.4]
  assign _T_57910 = $signed(_T_57909); // @[Modules.scala 37:46:@4260.4]
  assign _T_57915 = $signed(_T_54729) + $signed(io_in_169); // @[Modules.scala 43:47:@4265.4]
  assign _T_57916 = _T_57915[4:0]; // @[Modules.scala 43:47:@4266.4]
  assign _T_57917 = $signed(_T_57916); // @[Modules.scala 43:47:@4267.4]
  assign _T_57918 = $signed(io_in_170) + $signed(io_in_171); // @[Modules.scala 37:46:@4269.4]
  assign _T_57919 = _T_57918[4:0]; // @[Modules.scala 37:46:@4270.4]
  assign _T_57920 = $signed(_T_57919); // @[Modules.scala 37:46:@4271.4]
  assign _T_57924 = $signed(io_in_174) + $signed(io_in_175); // @[Modules.scala 37:46:@4277.4]
  assign _T_57925 = _T_57924[4:0]; // @[Modules.scala 37:46:@4278.4]
  assign _T_57926 = $signed(_T_57925); // @[Modules.scala 37:46:@4279.4]
  assign _T_57927 = $signed(io_in_176) + $signed(io_in_177); // @[Modules.scala 37:46:@4281.4]
  assign _T_57928 = _T_57927[4:0]; // @[Modules.scala 37:46:@4282.4]
  assign _T_57929 = $signed(_T_57928); // @[Modules.scala 37:46:@4283.4]
  assign _T_57930 = $signed(io_in_178) - $signed(io_in_179); // @[Modules.scala 40:46:@4285.4]
  assign _T_57931 = _T_57930[4:0]; // @[Modules.scala 40:46:@4286.4]
  assign _T_57932 = $signed(_T_57931); // @[Modules.scala 40:46:@4287.4]
  assign _T_57940 = $signed(io_in_182) - $signed(io_in_183); // @[Modules.scala 40:46:@4296.4]
  assign _T_57941 = _T_57940[4:0]; // @[Modules.scala 40:46:@4297.4]
  assign _T_57942 = $signed(_T_57941); // @[Modules.scala 40:46:@4298.4]
  assign _T_57953 = $signed(io_in_188) - $signed(io_in_189); // @[Modules.scala 40:46:@4311.4]
  assign _T_57954 = _T_57953[4:0]; // @[Modules.scala 40:46:@4312.4]
  assign _T_57955 = $signed(_T_57954); // @[Modules.scala 40:46:@4313.4]
  assign _T_57957 = $signed(5'sh0) - $signed(io_in_190); // @[Modules.scala 43:37:@4315.4]
  assign _T_57958 = _T_57957[4:0]; // @[Modules.scala 43:37:@4316.4]
  assign _T_57959 = $signed(_T_57958); // @[Modules.scala 43:37:@4317.4]
  assign _T_57960 = $signed(_T_57959) + $signed(io_in_191); // @[Modules.scala 43:47:@4318.4]
  assign _T_57961 = _T_57960[4:0]; // @[Modules.scala 43:47:@4319.4]
  assign _T_57962 = $signed(_T_57961); // @[Modules.scala 43:47:@4320.4]
  assign _T_57967 = $signed(_T_54801) + $signed(io_in_193); // @[Modules.scala 43:47:@4325.4]
  assign _T_57968 = _T_57967[4:0]; // @[Modules.scala 43:47:@4326.4]
  assign _T_57969 = $signed(_T_57968); // @[Modules.scala 43:47:@4327.4]
  assign _T_57974 = $signed(_T_54808) + $signed(io_in_195); // @[Modules.scala 43:47:@4332.4]
  assign _T_57975 = _T_57974[4:0]; // @[Modules.scala 43:47:@4333.4]
  assign _T_57976 = $signed(_T_57975); // @[Modules.scala 43:47:@4334.4]
  assign _T_57977 = $signed(io_in_196) + $signed(io_in_197); // @[Modules.scala 37:46:@4336.4]
  assign _T_57978 = _T_57977[4:0]; // @[Modules.scala 37:46:@4337.4]
  assign _T_57979 = $signed(_T_57978); // @[Modules.scala 37:46:@4338.4]
  assign _T_57981 = $signed(5'sh0) - $signed(io_in_198); // @[Modules.scala 43:37:@4340.4]
  assign _T_57982 = _T_57981[4:0]; // @[Modules.scala 43:37:@4341.4]
  assign _T_57983 = $signed(_T_57982); // @[Modules.scala 43:37:@4342.4]
  assign _T_57984 = $signed(_T_57983) + $signed(io_in_199); // @[Modules.scala 43:47:@4343.4]
  assign _T_57985 = _T_57984[4:0]; // @[Modules.scala 43:47:@4344.4]
  assign _T_57986 = $signed(_T_57985); // @[Modules.scala 43:47:@4345.4]
  assign _T_57991 = $signed(_T_54821) + $signed(io_in_201); // @[Modules.scala 43:47:@4350.4]
  assign _T_57992 = _T_57991[4:0]; // @[Modules.scala 43:47:@4351.4]
  assign _T_57993 = $signed(_T_57992); // @[Modules.scala 43:47:@4352.4]
  assign _T_57994 = $signed(io_in_202) + $signed(io_in_203); // @[Modules.scala 37:46:@4354.4]
  assign _T_57995 = _T_57994[4:0]; // @[Modules.scala 37:46:@4355.4]
  assign _T_57996 = $signed(_T_57995); // @[Modules.scala 37:46:@4356.4]
  assign _T_58001 = $signed(_T_54835) + $signed(io_in_205); // @[Modules.scala 43:47:@4361.4]
  assign _T_58002 = _T_58001[4:0]; // @[Modules.scala 43:47:@4362.4]
  assign _T_58003 = $signed(_T_58002); // @[Modules.scala 43:47:@4363.4]
  assign _T_58004 = $signed(io_in_206) - $signed(io_in_207); // @[Modules.scala 40:46:@4365.4]
  assign _T_58005 = _T_58004[4:0]; // @[Modules.scala 40:46:@4366.4]
  assign _T_58006 = $signed(_T_58005); // @[Modules.scala 40:46:@4367.4]
  assign _T_58007 = $signed(io_in_208) - $signed(io_in_209); // @[Modules.scala 40:46:@4369.4]
  assign _T_58008 = _T_58007[4:0]; // @[Modules.scala 40:46:@4370.4]
  assign _T_58009 = $signed(_T_58008); // @[Modules.scala 40:46:@4371.4]
  assign _T_58014 = $signed(5'sh0) - $signed(io_in_212); // @[Modules.scala 43:37:@4377.4]
  assign _T_58015 = _T_58014[4:0]; // @[Modules.scala 43:37:@4378.4]
  assign _T_58016 = $signed(_T_58015); // @[Modules.scala 43:37:@4379.4]
  assign _T_58017 = $signed(_T_58016) + $signed(io_in_213); // @[Modules.scala 43:47:@4380.4]
  assign _T_58018 = _T_58017[4:0]; // @[Modules.scala 43:47:@4381.4]
  assign _T_58019 = $signed(_T_58018); // @[Modules.scala 43:47:@4382.4]
  assign _T_58024 = $signed(_T_54862) + $signed(io_in_215); // @[Modules.scala 43:47:@4387.4]
  assign _T_58025 = _T_58024[4:0]; // @[Modules.scala 43:47:@4388.4]
  assign _T_58026 = $signed(_T_58025); // @[Modules.scala 43:47:@4389.4]
  assign _T_58031 = $signed(_T_54869) + $signed(io_in_217); // @[Modules.scala 43:47:@4394.4]
  assign _T_58032 = _T_58031[4:0]; // @[Modules.scala 43:47:@4395.4]
  assign _T_58033 = $signed(_T_58032); // @[Modules.scala 43:47:@4396.4]
  assign _T_58038 = $signed(_T_54876) + $signed(io_in_219); // @[Modules.scala 43:47:@4401.4]
  assign _T_58039 = _T_58038[4:0]; // @[Modules.scala 43:47:@4402.4]
  assign _T_58040 = $signed(_T_58039); // @[Modules.scala 43:47:@4403.4]
  assign _T_58041 = $signed(io_in_220) + $signed(io_in_221); // @[Modules.scala 37:46:@4405.4]
  assign _T_58042 = _T_58041[4:0]; // @[Modules.scala 37:46:@4406.4]
  assign _T_58043 = $signed(_T_58042); // @[Modules.scala 37:46:@4407.4]
  assign _T_58048 = $signed(_T_54890) + $signed(io_in_223); // @[Modules.scala 43:47:@4412.4]
  assign _T_58049 = _T_58048[4:0]; // @[Modules.scala 43:47:@4413.4]
  assign _T_58050 = $signed(_T_58049); // @[Modules.scala 43:47:@4414.4]
  assign _T_58051 = $signed(io_in_224) + $signed(io_in_225); // @[Modules.scala 37:46:@4416.4]
  assign _T_58052 = _T_58051[4:0]; // @[Modules.scala 37:46:@4417.4]
  assign _T_58053 = $signed(_T_58052); // @[Modules.scala 37:46:@4418.4]
  assign _T_58093 = $signed(_T_54939) - $signed(io_in_237); // @[Modules.scala 46:47:@4458.4]
  assign _T_58094 = _T_58093[4:0]; // @[Modules.scala 46:47:@4459.4]
  assign _T_58095 = $signed(_T_58094); // @[Modules.scala 46:47:@4460.4]
  assign _T_58103 = $signed(io_in_240) + $signed(io_in_241); // @[Modules.scala 37:46:@4469.4]
  assign _T_58104 = _T_58103[4:0]; // @[Modules.scala 37:46:@4470.4]
  assign _T_58105 = $signed(_T_58104); // @[Modules.scala 37:46:@4471.4]
  assign _T_58124 = $signed(_T_54974) + $signed(io_in_247); // @[Modules.scala 43:47:@4490.4]
  assign _T_58125 = _T_58124[4:0]; // @[Modules.scala 43:47:@4491.4]
  assign _T_58126 = $signed(_T_58125); // @[Modules.scala 43:47:@4492.4]
  assign _T_58127 = $signed(io_in_248) + $signed(io_in_249); // @[Modules.scala 37:46:@4494.4]
  assign _T_58128 = _T_58127[4:0]; // @[Modules.scala 37:46:@4495.4]
  assign _T_58129 = $signed(_T_58128); // @[Modules.scala 37:46:@4496.4]
  assign _T_58130 = $signed(io_in_250) + $signed(io_in_251); // @[Modules.scala 37:46:@4498.4]
  assign _T_58131 = _T_58130[4:0]; // @[Modules.scala 37:46:@4499.4]
  assign _T_58132 = $signed(_T_58131); // @[Modules.scala 37:46:@4500.4]
  assign _T_58137 = $signed(_T_54995) + $signed(io_in_253); // @[Modules.scala 43:47:@4505.4]
  assign _T_58138 = _T_58137[4:0]; // @[Modules.scala 43:47:@4506.4]
  assign _T_58139 = $signed(_T_58138); // @[Modules.scala 43:47:@4507.4]
  assign _T_58161 = $signed(io_in_260) - $signed(io_in_261); // @[Modules.scala 40:46:@4530.4]
  assign _T_58162 = _T_58161[4:0]; // @[Modules.scala 40:46:@4531.4]
  assign _T_58163 = $signed(_T_58162); // @[Modules.scala 40:46:@4532.4]
  assign _T_58165 = $signed(5'sh0) - $signed(io_in_262); // @[Modules.scala 46:37:@4534.4]
  assign _T_58166 = _T_58165[4:0]; // @[Modules.scala 46:37:@4535.4]
  assign _T_58167 = $signed(_T_58166); // @[Modules.scala 46:37:@4536.4]
  assign _T_58168 = $signed(_T_58167) - $signed(io_in_263); // @[Modules.scala 46:47:@4537.4]
  assign _T_58169 = _T_58168[4:0]; // @[Modules.scala 46:47:@4538.4]
  assign _T_58170 = $signed(_T_58169); // @[Modules.scala 46:47:@4539.4]
  assign _T_58178 = $signed(io_in_266) + $signed(io_in_267); // @[Modules.scala 37:46:@4548.4]
  assign _T_58179 = _T_58178[4:0]; // @[Modules.scala 37:46:@4549.4]
  assign _T_58180 = $signed(_T_58179); // @[Modules.scala 37:46:@4550.4]
  assign _T_58206 = $signed(_T_55068) + $signed(io_in_275); // @[Modules.scala 43:47:@4576.4]
  assign _T_58207 = _T_58206[4:0]; // @[Modules.scala 43:47:@4577.4]
  assign _T_58208 = $signed(_T_58207); // @[Modules.scala 43:47:@4578.4]
  assign _T_58209 = $signed(io_in_276) + $signed(io_in_277); // @[Modules.scala 37:46:@4580.4]
  assign _T_58210 = _T_58209[4:0]; // @[Modules.scala 37:46:@4581.4]
  assign _T_58211 = $signed(_T_58210); // @[Modules.scala 37:46:@4582.4]
  assign _T_58212 = $signed(io_in_278) + $signed(io_in_279); // @[Modules.scala 37:46:@4584.4]
  assign _T_58213 = _T_58212[4:0]; // @[Modules.scala 37:46:@4585.4]
  assign _T_58214 = $signed(_T_58213); // @[Modules.scala 37:46:@4586.4]
  assign _T_58219 = $signed(_T_55089) + $signed(io_in_281); // @[Modules.scala 43:47:@4591.4]
  assign _T_58220 = _T_58219[4:0]; // @[Modules.scala 43:47:@4592.4]
  assign _T_58221 = $signed(_T_58220); // @[Modules.scala 43:47:@4593.4]
  assign _T_58226 = $signed(_T_55096) + $signed(io_in_283); // @[Modules.scala 43:47:@4598.4]
  assign _T_58227 = _T_58226[4:0]; // @[Modules.scala 43:47:@4599.4]
  assign _T_58228 = $signed(_T_58227); // @[Modules.scala 43:47:@4600.4]
  assign _T_58257 = $signed(io_in_292) + $signed(io_in_293); // @[Modules.scala 37:46:@4630.4]
  assign _T_58258 = _T_58257[4:0]; // @[Modules.scala 37:46:@4631.4]
  assign _T_58259 = $signed(_T_58258); // @[Modules.scala 37:46:@4632.4]
  assign _T_58260 = $signed(io_in_294) - $signed(io_in_295); // @[Modules.scala 40:46:@4634.4]
  assign _T_58261 = _T_58260[4:0]; // @[Modules.scala 40:46:@4635.4]
  assign _T_58262 = $signed(_T_58261); // @[Modules.scala 40:46:@4636.4]
  assign _T_58288 = $signed(_T_55166) + $signed(io_in_303); // @[Modules.scala 43:47:@4662.4]
  assign _T_58289 = _T_58288[4:0]; // @[Modules.scala 43:47:@4663.4]
  assign _T_58290 = $signed(_T_58289); // @[Modules.scala 43:47:@4664.4]
  assign _T_58291 = $signed(io_in_304) + $signed(io_in_305); // @[Modules.scala 37:46:@4666.4]
  assign _T_58292 = _T_58291[4:0]; // @[Modules.scala 37:46:@4667.4]
  assign _T_58293 = $signed(_T_58292); // @[Modules.scala 37:46:@4668.4]
  assign _T_58294 = $signed(io_in_306) + $signed(io_in_307); // @[Modules.scala 37:46:@4670.4]
  assign _T_58295 = _T_58294[4:0]; // @[Modules.scala 37:46:@4671.4]
  assign _T_58296 = $signed(_T_58295); // @[Modules.scala 37:46:@4672.4]
  assign _T_58318 = $signed(io_in_314) - $signed(io_in_315); // @[Modules.scala 40:46:@4695.4]
  assign _T_58319 = _T_58318[4:0]; // @[Modules.scala 40:46:@4696.4]
  assign _T_58320 = $signed(_T_58319); // @[Modules.scala 40:46:@4697.4]
  assign _T_58322 = $signed(5'sh0) - $signed(io_in_316); // @[Modules.scala 46:37:@4699.4]
  assign _T_58323 = _T_58322[4:0]; // @[Modules.scala 46:37:@4700.4]
  assign _T_58324 = $signed(_T_58323); // @[Modules.scala 46:37:@4701.4]
  assign _T_58325 = $signed(_T_58324) - $signed(io_in_317); // @[Modules.scala 46:47:@4702.4]
  assign _T_58326 = _T_58325[4:0]; // @[Modules.scala 46:47:@4703.4]
  assign _T_58327 = $signed(_T_58326); // @[Modules.scala 46:47:@4704.4]
  assign _T_58331 = $signed(io_in_320) + $signed(io_in_321); // @[Modules.scala 37:46:@4710.4]
  assign _T_58332 = _T_58331[4:0]; // @[Modules.scala 37:46:@4711.4]
  assign _T_58333 = $signed(_T_58332); // @[Modules.scala 37:46:@4712.4]
  assign _T_58334 = $signed(io_in_322) - $signed(io_in_323); // @[Modules.scala 40:46:@4714.4]
  assign _T_58335 = _T_58334[4:0]; // @[Modules.scala 40:46:@4715.4]
  assign _T_58336 = $signed(_T_58335); // @[Modules.scala 40:46:@4716.4]
  assign _T_58341 = $signed(_T_55235) - $signed(io_in_325); // @[Modules.scala 46:47:@4721.4]
  assign _T_58342 = _T_58341[4:0]; // @[Modules.scala 46:47:@4722.4]
  assign _T_58343 = $signed(_T_58342); // @[Modules.scala 46:47:@4723.4]
  assign _T_58352 = $signed(5'sh0) - $signed(io_in_328); // @[Modules.scala 46:37:@4732.4]
  assign _T_58353 = _T_58352[4:0]; // @[Modules.scala 46:37:@4733.4]
  assign _T_58354 = $signed(_T_58353); // @[Modules.scala 46:37:@4734.4]
  assign _T_58355 = $signed(_T_58354) - $signed(io_in_329); // @[Modules.scala 46:47:@4735.4]
  assign _T_58356 = _T_58355[4:0]; // @[Modules.scala 46:47:@4736.4]
  assign _T_58357 = $signed(_T_58356); // @[Modules.scala 46:47:@4737.4]
  assign _T_58362 = $signed(_T_55252) + $signed(io_in_331); // @[Modules.scala 43:47:@4742.4]
  assign _T_58363 = _T_58362[4:0]; // @[Modules.scala 43:47:@4743.4]
  assign _T_58364 = $signed(_T_58363); // @[Modules.scala 43:47:@4744.4]
  assign _T_58365 = $signed(io_in_332) + $signed(io_in_333); // @[Modules.scala 37:46:@4746.4]
  assign _T_58366 = _T_58365[4:0]; // @[Modules.scala 37:46:@4747.4]
  assign _T_58367 = $signed(_T_58366); // @[Modules.scala 37:46:@4748.4]
  assign _T_58368 = $signed(io_in_334) + $signed(io_in_335); // @[Modules.scala 37:46:@4750.4]
  assign _T_58369 = _T_58368[4:0]; // @[Modules.scala 37:46:@4751.4]
  assign _T_58370 = $signed(_T_58369); // @[Modules.scala 37:46:@4752.4]
  assign _T_58401 = $signed(5'sh0) - $signed(io_in_350); // @[Modules.scala 46:37:@4788.4]
  assign _T_58402 = _T_58401[4:0]; // @[Modules.scala 46:37:@4789.4]
  assign _T_58403 = $signed(_T_58402); // @[Modules.scala 46:37:@4790.4]
  assign _T_58404 = $signed(_T_58403) - $signed(io_in_351); // @[Modules.scala 46:47:@4791.4]
  assign _T_58405 = _T_58404[4:0]; // @[Modules.scala 46:47:@4792.4]
  assign _T_58406 = $signed(_T_58405); // @[Modules.scala 46:47:@4793.4]
  assign _T_58408 = $signed(5'sh0) - $signed(io_in_352); // @[Modules.scala 46:37:@4795.4]
  assign _T_58409 = _T_58408[4:0]; // @[Modules.scala 46:37:@4796.4]
  assign _T_58410 = $signed(_T_58409); // @[Modules.scala 46:37:@4797.4]
  assign _T_58411 = $signed(_T_58410) - $signed(io_in_353); // @[Modules.scala 46:47:@4798.4]
  assign _T_58412 = _T_58411[4:0]; // @[Modules.scala 46:47:@4799.4]
  assign _T_58413 = $signed(_T_58412); // @[Modules.scala 46:47:@4800.4]
  assign _T_58415 = $signed(5'sh0) - $signed(io_in_354); // @[Modules.scala 46:37:@4802.4]
  assign _T_58416 = _T_58415[4:0]; // @[Modules.scala 46:37:@4803.4]
  assign _T_58417 = $signed(_T_58416); // @[Modules.scala 46:37:@4804.4]
  assign _T_58418 = $signed(_T_58417) - $signed(io_in_355); // @[Modules.scala 46:47:@4805.4]
  assign _T_58419 = _T_58418[4:0]; // @[Modules.scala 46:47:@4806.4]
  assign _T_58420 = $signed(_T_58419); // @[Modules.scala 46:47:@4807.4]
  assign _T_58422 = $signed(5'sh0) - $signed(io_in_356); // @[Modules.scala 46:37:@4809.4]
  assign _T_58423 = _T_58422[4:0]; // @[Modules.scala 46:37:@4810.4]
  assign _T_58424 = $signed(_T_58423); // @[Modules.scala 46:37:@4811.4]
  assign _T_58425 = $signed(_T_58424) - $signed(io_in_357); // @[Modules.scala 46:47:@4812.4]
  assign _T_58426 = _T_58425[4:0]; // @[Modules.scala 46:47:@4813.4]
  assign _T_58427 = $signed(_T_58426); // @[Modules.scala 46:47:@4814.4]
  assign _T_58429 = $signed(5'sh0) - $signed(io_in_358); // @[Modules.scala 43:37:@4816.4]
  assign _T_58430 = _T_58429[4:0]; // @[Modules.scala 43:37:@4817.4]
  assign _T_58431 = $signed(_T_58430); // @[Modules.scala 43:37:@4818.4]
  assign _T_58432 = $signed(_T_58431) + $signed(io_in_359); // @[Modules.scala 43:47:@4819.4]
  assign _T_58433 = _T_58432[4:0]; // @[Modules.scala 43:47:@4820.4]
  assign _T_58434 = $signed(_T_58433); // @[Modules.scala 43:47:@4821.4]
  assign _T_58435 = $signed(io_in_360) + $signed(io_in_361); // @[Modules.scala 37:46:@4823.4]
  assign _T_58436 = _T_58435[4:0]; // @[Modules.scala 37:46:@4824.4]
  assign _T_58437 = $signed(_T_58436); // @[Modules.scala 37:46:@4825.4]
  assign _T_58442 = $signed(_T_55324) - $signed(io_in_363); // @[Modules.scala 46:47:@4830.4]
  assign _T_58443 = _T_58442[4:0]; // @[Modules.scala 46:47:@4831.4]
  assign _T_58444 = $signed(_T_58443); // @[Modules.scala 46:47:@4832.4]
  assign _T_58460 = $signed(5'sh0) - $signed(io_in_368); // @[Modules.scala 43:37:@4848.4]
  assign _T_58461 = _T_58460[4:0]; // @[Modules.scala 43:37:@4849.4]
  assign _T_58462 = $signed(_T_58461); // @[Modules.scala 43:37:@4850.4]
  assign _T_58463 = $signed(_T_58462) + $signed(io_in_369); // @[Modules.scala 43:47:@4851.4]
  assign _T_58464 = _T_58463[4:0]; // @[Modules.scala 43:47:@4852.4]
  assign _T_58465 = $signed(_T_58464); // @[Modules.scala 43:47:@4853.4]
  assign _T_58479 = $signed(5'sh0) - $signed(io_in_378); // @[Modules.scala 46:37:@4871.4]
  assign _T_58480 = _T_58479[4:0]; // @[Modules.scala 46:37:@4872.4]
  assign _T_58481 = $signed(_T_58480); // @[Modules.scala 46:37:@4873.4]
  assign _T_58482 = $signed(_T_58481) - $signed(io_in_379); // @[Modules.scala 46:47:@4874.4]
  assign _T_58483 = _T_58482[4:0]; // @[Modules.scala 46:47:@4875.4]
  assign _T_58484 = $signed(_T_58483); // @[Modules.scala 46:47:@4876.4]
  assign _T_58486 = $signed(5'sh0) - $signed(io_in_380); // @[Modules.scala 46:37:@4878.4]
  assign _T_58487 = _T_58486[4:0]; // @[Modules.scala 46:37:@4879.4]
  assign _T_58488 = $signed(_T_58487); // @[Modules.scala 46:37:@4880.4]
  assign _T_58489 = $signed(_T_58488) - $signed(io_in_381); // @[Modules.scala 46:47:@4881.4]
  assign _T_58490 = _T_58489[4:0]; // @[Modules.scala 46:47:@4882.4]
  assign _T_58491 = $signed(_T_58490); // @[Modules.scala 46:47:@4883.4]
  assign _T_58493 = $signed(5'sh0) - $signed(io_in_382); // @[Modules.scala 46:37:@4885.4]
  assign _T_58494 = _T_58493[4:0]; // @[Modules.scala 46:37:@4886.4]
  assign _T_58495 = $signed(_T_58494); // @[Modules.scala 46:37:@4887.4]
  assign _T_58496 = $signed(_T_58495) - $signed(io_in_383); // @[Modules.scala 46:47:@4888.4]
  assign _T_58497 = _T_58496[4:0]; // @[Modules.scala 46:47:@4889.4]
  assign _T_58498 = $signed(_T_58497); // @[Modules.scala 46:47:@4890.4]
  assign _T_58516 = $signed(_T_55382) - $signed(io_in_391); // @[Modules.scala 46:47:@4910.4]
  assign _T_58517 = _T_58516[4:0]; // @[Modules.scala 46:47:@4911.4]
  assign _T_58518 = $signed(_T_58517); // @[Modules.scala 46:47:@4912.4]
  assign _T_58519 = $signed(io_in_392) + $signed(io_in_393); // @[Modules.scala 37:46:@4914.4]
  assign _T_58520 = _T_58519[4:0]; // @[Modules.scala 37:46:@4915.4]
  assign _T_58521 = $signed(_T_58520); // @[Modules.scala 37:46:@4916.4]
  assign _T_58530 = $signed(5'sh0) - $signed(io_in_396); // @[Modules.scala 43:37:@4925.4]
  assign _T_58531 = _T_58530[4:0]; // @[Modules.scala 43:37:@4926.4]
  assign _T_58532 = $signed(_T_58531); // @[Modules.scala 43:37:@4927.4]
  assign _T_58533 = $signed(_T_58532) + $signed(io_in_397); // @[Modules.scala 43:47:@4928.4]
  assign _T_58534 = _T_58533[4:0]; // @[Modules.scala 43:47:@4929.4]
  assign _T_58535 = $signed(_T_58534); // @[Modules.scala 43:47:@4930.4]
  assign _T_58545 = $signed(io_in_404) - $signed(io_in_405); // @[Modules.scala 40:46:@4944.4]
  assign _T_58546 = _T_58545[4:0]; // @[Modules.scala 40:46:@4945.4]
  assign _T_58547 = $signed(_T_58546); // @[Modules.scala 40:46:@4946.4]
  assign _T_58549 = $signed(5'sh0) - $signed(io_in_406); // @[Modules.scala 46:37:@4948.4]
  assign _T_58550 = _T_58549[4:0]; // @[Modules.scala 46:37:@4949.4]
  assign _T_58551 = $signed(_T_58550); // @[Modules.scala 46:37:@4950.4]
  assign _T_58552 = $signed(_T_58551) - $signed(io_in_407); // @[Modules.scala 46:47:@4951.4]
  assign _T_58553 = _T_58552[4:0]; // @[Modules.scala 46:47:@4952.4]
  assign _T_58554 = $signed(_T_58553); // @[Modules.scala 46:47:@4953.4]
  assign _T_58555 = $signed(io_in_408) - $signed(io_in_409); // @[Modules.scala 40:46:@4955.4]
  assign _T_58556 = _T_58555[4:0]; // @[Modules.scala 40:46:@4956.4]
  assign _T_58557 = $signed(_T_58556); // @[Modules.scala 40:46:@4957.4]
  assign _T_58559 = $signed(5'sh0) - $signed(io_in_410); // @[Modules.scala 46:37:@4959.4]
  assign _T_58560 = _T_58559[4:0]; // @[Modules.scala 46:37:@4960.4]
  assign _T_58561 = $signed(_T_58560); // @[Modules.scala 46:37:@4961.4]
  assign _T_58562 = $signed(_T_58561) - $signed(io_in_411); // @[Modules.scala 46:47:@4962.4]
  assign _T_58563 = _T_58562[4:0]; // @[Modules.scala 46:47:@4963.4]
  assign _T_58564 = $signed(_T_58563); // @[Modules.scala 46:47:@4964.4]
  assign _T_58578 = $signed(_T_55436) - $signed(io_in_419); // @[Modules.scala 46:47:@4981.4]
  assign _T_58579 = _T_58578[4:0]; // @[Modules.scala 46:47:@4982.4]
  assign _T_58580 = $signed(_T_58579); // @[Modules.scala 46:47:@4983.4]
  assign _T_58588 = $signed(io_in_422) - $signed(io_in_423); // @[Modules.scala 40:46:@4992.4]
  assign _T_58589 = _T_58588[4:0]; // @[Modules.scala 40:46:@4993.4]
  assign _T_58590 = $signed(_T_58589); // @[Modules.scala 40:46:@4994.4]
  assign _T_58599 = $signed(5'sh0) - $signed(io_in_426); // @[Modules.scala 46:37:@5003.4]
  assign _T_58600 = _T_58599[4:0]; // @[Modules.scala 46:37:@5004.4]
  assign _T_58601 = $signed(_T_58600); // @[Modules.scala 46:37:@5005.4]
  assign _T_58602 = $signed(_T_58601) - $signed(io_in_427); // @[Modules.scala 46:47:@5006.4]
  assign _T_58603 = _T_58602[4:0]; // @[Modules.scala 46:47:@5007.4]
  assign _T_58604 = $signed(_T_58603); // @[Modules.scala 46:47:@5008.4]
  assign _T_58612 = $signed(5'sh0) - $signed(io_in_432); // @[Modules.scala 46:37:@5018.4]
  assign _T_58613 = _T_58612[4:0]; // @[Modules.scala 46:37:@5019.4]
  assign _T_58614 = $signed(_T_58613); // @[Modules.scala 46:37:@5020.4]
  assign _T_58615 = $signed(_T_58614) - $signed(io_in_433); // @[Modules.scala 46:47:@5021.4]
  assign _T_58616 = _T_58615[4:0]; // @[Modules.scala 46:47:@5022.4]
  assign _T_58617 = $signed(_T_58616); // @[Modules.scala 46:47:@5023.4]
  assign _T_58619 = $signed(5'sh0) - $signed(io_in_434); // @[Modules.scala 46:37:@5025.4]
  assign _T_58620 = _T_58619[4:0]; // @[Modules.scala 46:37:@5026.4]
  assign _T_58621 = $signed(_T_58620); // @[Modules.scala 46:37:@5027.4]
  assign _T_58622 = $signed(_T_58621) - $signed(io_in_435); // @[Modules.scala 46:47:@5028.4]
  assign _T_58623 = _T_58622[4:0]; // @[Modules.scala 46:47:@5029.4]
  assign _T_58624 = $signed(_T_58623); // @[Modules.scala 46:47:@5030.4]
  assign _T_58626 = $signed(5'sh0) - $signed(io_in_436); // @[Modules.scala 46:37:@5032.4]
  assign _T_58627 = _T_58626[4:0]; // @[Modules.scala 46:37:@5033.4]
  assign _T_58628 = $signed(_T_58627); // @[Modules.scala 46:37:@5034.4]
  assign _T_58629 = $signed(_T_58628) - $signed(io_in_437); // @[Modules.scala 46:47:@5035.4]
  assign _T_58630 = _T_58629[4:0]; // @[Modules.scala 46:47:@5036.4]
  assign _T_58631 = $signed(_T_58630); // @[Modules.scala 46:47:@5037.4]
  assign _T_58633 = $signed(5'sh0) - $signed(io_in_438); // @[Modules.scala 43:37:@5039.4]
  assign _T_58634 = _T_58633[4:0]; // @[Modules.scala 43:37:@5040.4]
  assign _T_58635 = $signed(_T_58634); // @[Modules.scala 43:37:@5041.4]
  assign _T_58636 = $signed(_T_58635) + $signed(io_in_439); // @[Modules.scala 43:47:@5042.4]
  assign _T_58637 = _T_58636[4:0]; // @[Modules.scala 43:47:@5043.4]
  assign _T_58638 = $signed(_T_58637); // @[Modules.scala 43:47:@5044.4]
  assign _T_58639 = $signed(io_in_440) + $signed(io_in_441); // @[Modules.scala 37:46:@5046.4]
  assign _T_58640 = _T_58639[4:0]; // @[Modules.scala 37:46:@5047.4]
  assign _T_58641 = $signed(_T_58640); // @[Modules.scala 37:46:@5048.4]
  assign _T_58642 = $signed(io_in_442) + $signed(io_in_443); // @[Modules.scala 37:46:@5050.4]
  assign _T_58643 = _T_58642[4:0]; // @[Modules.scala 37:46:@5051.4]
  assign _T_58644 = $signed(_T_58643); // @[Modules.scala 37:46:@5052.4]
  assign _T_58645 = $signed(io_in_444) - $signed(io_in_445); // @[Modules.scala 40:46:@5054.4]
  assign _T_58646 = _T_58645[4:0]; // @[Modules.scala 40:46:@5055.4]
  assign _T_58647 = $signed(_T_58646); // @[Modules.scala 40:46:@5056.4]
  assign _T_58656 = $signed(5'sh0) - $signed(io_in_448); // @[Modules.scala 43:37:@5065.4]
  assign _T_58657 = _T_58656[4:0]; // @[Modules.scala 43:37:@5066.4]
  assign _T_58658 = $signed(_T_58657); // @[Modules.scala 43:37:@5067.4]
  assign _T_58659 = $signed(_T_58658) + $signed(io_in_449); // @[Modules.scala 43:47:@5068.4]
  assign _T_58660 = _T_58659[4:0]; // @[Modules.scala 43:47:@5069.4]
  assign _T_58661 = $signed(_T_58660); // @[Modules.scala 43:47:@5070.4]
  assign _T_58662 = $signed(io_in_450) + $signed(io_in_451); // @[Modules.scala 37:46:@5072.4]
  assign _T_58663 = _T_58662[4:0]; // @[Modules.scala 37:46:@5073.4]
  assign _T_58664 = $signed(_T_58663); // @[Modules.scala 37:46:@5074.4]
  assign _T_58669 = $signed(_T_55519) - $signed(io_in_453); // @[Modules.scala 46:47:@5079.4]
  assign _T_58670 = _T_58669[4:0]; // @[Modules.scala 46:47:@5080.4]
  assign _T_58671 = $signed(_T_58670); // @[Modules.scala 46:47:@5081.4]
  assign _T_58673 = $signed(5'sh0) - $signed(io_in_454); // @[Modules.scala 46:37:@5083.4]
  assign _T_58674 = _T_58673[4:0]; // @[Modules.scala 46:37:@5084.4]
  assign _T_58675 = $signed(_T_58674); // @[Modules.scala 46:37:@5085.4]
  assign _T_58676 = $signed(_T_58675) - $signed(io_in_455); // @[Modules.scala 46:47:@5086.4]
  assign _T_58677 = _T_58676[4:0]; // @[Modules.scala 46:47:@5087.4]
  assign _T_58678 = $signed(_T_58677); // @[Modules.scala 46:47:@5088.4]
  assign _T_58680 = $signed(5'sh0) - $signed(io_in_456); // @[Modules.scala 43:37:@5090.4]
  assign _T_58681 = _T_58680[4:0]; // @[Modules.scala 43:37:@5091.4]
  assign _T_58682 = $signed(_T_58681); // @[Modules.scala 43:37:@5092.4]
  assign _T_58683 = $signed(_T_58682) + $signed(io_in_457); // @[Modules.scala 43:47:@5093.4]
  assign _T_58684 = _T_58683[4:0]; // @[Modules.scala 43:47:@5094.4]
  assign _T_58685 = $signed(_T_58684); // @[Modules.scala 43:47:@5095.4]
  assign _T_58686 = $signed(io_in_458) - $signed(io_in_459); // @[Modules.scala 40:46:@5097.4]
  assign _T_58687 = _T_58686[4:0]; // @[Modules.scala 40:46:@5098.4]
  assign _T_58688 = $signed(_T_58687); // @[Modules.scala 40:46:@5099.4]
  assign _T_58690 = $signed(5'sh0) - $signed(io_in_460); // @[Modules.scala 46:37:@5101.4]
  assign _T_58691 = _T_58690[4:0]; // @[Modules.scala 46:37:@5102.4]
  assign _T_58692 = $signed(_T_58691); // @[Modules.scala 46:37:@5103.4]
  assign _T_58693 = $signed(_T_58692) - $signed(io_in_461); // @[Modules.scala 46:47:@5104.4]
  assign _T_58694 = _T_58693[4:0]; // @[Modules.scala 46:47:@5105.4]
  assign _T_58695 = $signed(_T_58694); // @[Modules.scala 46:47:@5106.4]
  assign _T_58697 = $signed(5'sh0) - $signed(io_in_462); // @[Modules.scala 46:37:@5108.4]
  assign _T_58698 = _T_58697[4:0]; // @[Modules.scala 46:37:@5109.4]
  assign _T_58699 = $signed(_T_58698); // @[Modules.scala 46:37:@5110.4]
  assign _T_58700 = $signed(_T_58699) - $signed(io_in_463); // @[Modules.scala 46:47:@5111.4]
  assign _T_58701 = _T_58700[4:0]; // @[Modules.scala 46:47:@5112.4]
  assign _T_58702 = $signed(_T_58701); // @[Modules.scala 46:47:@5113.4]
  assign _T_58704 = $signed(5'sh0) - $signed(io_in_464); // @[Modules.scala 46:37:@5115.4]
  assign _T_58705 = _T_58704[4:0]; // @[Modules.scala 46:37:@5116.4]
  assign _T_58706 = $signed(_T_58705); // @[Modules.scala 46:37:@5117.4]
  assign _T_58707 = $signed(_T_58706) - $signed(io_in_465); // @[Modules.scala 46:47:@5118.4]
  assign _T_58708 = _T_58707[4:0]; // @[Modules.scala 46:47:@5119.4]
  assign _T_58709 = $signed(_T_58708); // @[Modules.scala 46:47:@5120.4]
  assign _T_58711 = $signed(5'sh0) - $signed(io_in_466); // @[Modules.scala 43:37:@5122.4]
  assign _T_58712 = _T_58711[4:0]; // @[Modules.scala 43:37:@5123.4]
  assign _T_58713 = $signed(_T_58712); // @[Modules.scala 43:37:@5124.4]
  assign _T_58714 = $signed(_T_58713) + $signed(io_in_467); // @[Modules.scala 43:47:@5125.4]
  assign _T_58715 = _T_58714[4:0]; // @[Modules.scala 43:47:@5126.4]
  assign _T_58716 = $signed(_T_58715); // @[Modules.scala 43:47:@5127.4]
  assign _T_58717 = $signed(io_in_468) + $signed(io_in_469); // @[Modules.scala 37:46:@5129.4]
  assign _T_58718 = _T_58717[4:0]; // @[Modules.scala 37:46:@5130.4]
  assign _T_58719 = $signed(_T_58718); // @[Modules.scala 37:46:@5131.4]
  assign _T_58720 = $signed(io_in_470) + $signed(io_in_471); // @[Modules.scala 37:46:@5133.4]
  assign _T_58721 = _T_58720[4:0]; // @[Modules.scala 37:46:@5134.4]
  assign _T_58722 = $signed(_T_58721); // @[Modules.scala 37:46:@5135.4]
  assign _T_58723 = $signed(io_in_472) - $signed(io_in_473); // @[Modules.scala 40:46:@5137.4]
  assign _T_58724 = _T_58723[4:0]; // @[Modules.scala 40:46:@5138.4]
  assign _T_58725 = $signed(_T_58724); // @[Modules.scala 40:46:@5139.4]
  assign _T_58737 = $signed(_T_55571) + $signed(io_in_477); // @[Modules.scala 43:47:@5151.4]
  assign _T_58738 = _T_58737[4:0]; // @[Modules.scala 43:47:@5152.4]
  assign _T_58739 = $signed(_T_58738); // @[Modules.scala 43:47:@5153.4]
  assign _T_58740 = $signed(io_in_478) + $signed(io_in_479); // @[Modules.scala 37:46:@5155.4]
  assign _T_58741 = _T_58740[4:0]; // @[Modules.scala 37:46:@5156.4]
  assign _T_58742 = $signed(_T_58741); // @[Modules.scala 37:46:@5157.4]
  assign _T_58754 = $signed(5'sh0) - $signed(io_in_484); // @[Modules.scala 46:37:@5170.4]
  assign _T_58755 = _T_58754[4:0]; // @[Modules.scala 46:37:@5171.4]
  assign _T_58756 = $signed(_T_58755); // @[Modules.scala 46:37:@5172.4]
  assign _T_58757 = $signed(_T_58756) - $signed(io_in_485); // @[Modules.scala 46:47:@5173.4]
  assign _T_58758 = _T_58757[4:0]; // @[Modules.scala 46:47:@5174.4]
  assign _T_58759 = $signed(_T_58758); // @[Modules.scala 46:47:@5175.4]
  assign _T_58761 = $signed(5'sh0) - $signed(io_in_486); // @[Modules.scala 46:37:@5177.4]
  assign _T_58762 = _T_58761[4:0]; // @[Modules.scala 46:37:@5178.4]
  assign _T_58763 = $signed(_T_58762); // @[Modules.scala 46:37:@5179.4]
  assign _T_58764 = $signed(_T_58763) - $signed(io_in_487); // @[Modules.scala 46:47:@5180.4]
  assign _T_58765 = _T_58764[4:0]; // @[Modules.scala 46:47:@5181.4]
  assign _T_58766 = $signed(_T_58765); // @[Modules.scala 46:47:@5182.4]
  assign _T_58771 = $signed(_T_55597) - $signed(io_in_489); // @[Modules.scala 46:47:@5187.4]
  assign _T_58772 = _T_58771[4:0]; // @[Modules.scala 46:47:@5188.4]
  assign _T_58773 = $signed(_T_58772); // @[Modules.scala 46:47:@5189.4]
  assign _T_58775 = $signed(5'sh0) - $signed(io_in_490); // @[Modules.scala 46:37:@5191.4]
  assign _T_58776 = _T_58775[4:0]; // @[Modules.scala 46:37:@5192.4]
  assign _T_58777 = $signed(_T_58776); // @[Modules.scala 46:37:@5193.4]
  assign _T_58778 = $signed(_T_58777) - $signed(io_in_491); // @[Modules.scala 46:47:@5194.4]
  assign _T_58779 = _T_58778[4:0]; // @[Modules.scala 46:47:@5195.4]
  assign _T_58780 = $signed(_T_58779); // @[Modules.scala 46:47:@5196.4]
  assign _T_58782 = $signed(5'sh0) - $signed(io_in_492); // @[Modules.scala 46:37:@5198.4]
  assign _T_58783 = _T_58782[4:0]; // @[Modules.scala 46:37:@5199.4]
  assign _T_58784 = $signed(_T_58783); // @[Modules.scala 46:37:@5200.4]
  assign _T_58785 = $signed(_T_58784) - $signed(io_in_493); // @[Modules.scala 46:47:@5201.4]
  assign _T_58786 = _T_58785[4:0]; // @[Modules.scala 46:47:@5202.4]
  assign _T_58787 = $signed(_T_58786); // @[Modules.scala 46:47:@5203.4]
  assign _T_58788 = $signed(io_in_494) + $signed(io_in_495); // @[Modules.scala 37:46:@5205.4]
  assign _T_58789 = _T_58788[4:0]; // @[Modules.scala 37:46:@5206.4]
  assign _T_58790 = $signed(_T_58789); // @[Modules.scala 37:46:@5207.4]
  assign _T_58791 = $signed(io_in_496) + $signed(io_in_497); // @[Modules.scala 37:46:@5209.4]
  assign _T_58792 = _T_58791[4:0]; // @[Modules.scala 37:46:@5210.4]
  assign _T_58793 = $signed(_T_58792); // @[Modules.scala 37:46:@5211.4]
  assign _T_58815 = $signed(_T_55637) + $signed(io_in_505); // @[Modules.scala 43:47:@5234.4]
  assign _T_58816 = _T_58815[4:0]; // @[Modules.scala 43:47:@5235.4]
  assign _T_58817 = $signed(_T_58816); // @[Modules.scala 43:47:@5236.4]
  assign _T_58818 = $signed(io_in_506) + $signed(io_in_507); // @[Modules.scala 37:46:@5238.4]
  assign _T_58819 = _T_58818[4:0]; // @[Modules.scala 37:46:@5239.4]
  assign _T_58820 = $signed(_T_58819); // @[Modules.scala 37:46:@5240.4]
  assign _T_58821 = $signed(io_in_508) - $signed(io_in_509); // @[Modules.scala 40:46:@5242.4]
  assign _T_58822 = _T_58821[4:0]; // @[Modules.scala 40:46:@5243.4]
  assign _T_58823 = $signed(_T_58822); // @[Modules.scala 40:46:@5244.4]
  assign _T_58824 = $signed(io_in_510) + $signed(io_in_511); // @[Modules.scala 37:46:@5246.4]
  assign _T_58825 = _T_58824[4:0]; // @[Modules.scala 37:46:@5247.4]
  assign _T_58826 = $signed(_T_58825); // @[Modules.scala 37:46:@5248.4]
  assign _T_58828 = $signed(5'sh0) - $signed(io_in_512); // @[Modules.scala 46:37:@5250.4]
  assign _T_58829 = _T_58828[4:0]; // @[Modules.scala 46:37:@5251.4]
  assign _T_58830 = $signed(_T_58829); // @[Modules.scala 46:37:@5252.4]
  assign _T_58831 = $signed(_T_58830) - $signed(io_in_513); // @[Modules.scala 46:47:@5253.4]
  assign _T_58832 = _T_58831[4:0]; // @[Modules.scala 46:47:@5254.4]
  assign _T_58833 = $signed(_T_58832); // @[Modules.scala 46:47:@5255.4]
  assign _T_58838 = $signed(5'sh0) - $signed(io_in_516); // @[Modules.scala 46:37:@5261.4]
  assign _T_58839 = _T_58838[4:0]; // @[Modules.scala 46:37:@5262.4]
  assign _T_58840 = $signed(_T_58839); // @[Modules.scala 46:37:@5263.4]
  assign _T_58841 = $signed(_T_58840) - $signed(io_in_517); // @[Modules.scala 46:47:@5264.4]
  assign _T_58842 = _T_58841[4:0]; // @[Modules.scala 46:47:@5265.4]
  assign _T_58843 = $signed(_T_58842); // @[Modules.scala 46:47:@5266.4]
  assign _T_58845 = $signed(5'sh0) - $signed(io_in_518); // @[Modules.scala 46:37:@5268.4]
  assign _T_58846 = _T_58845[4:0]; // @[Modules.scala 46:37:@5269.4]
  assign _T_58847 = $signed(_T_58846); // @[Modules.scala 46:37:@5270.4]
  assign _T_58848 = $signed(_T_58847) - $signed(io_in_519); // @[Modules.scala 46:47:@5271.4]
  assign _T_58849 = _T_58848[4:0]; // @[Modules.scala 46:47:@5272.4]
  assign _T_58850 = $signed(_T_58849); // @[Modules.scala 46:47:@5273.4]
  assign _T_58851 = $signed(io_in_520) + $signed(io_in_521); // @[Modules.scala 37:46:@5275.4]
  assign _T_58852 = _T_58851[4:0]; // @[Modules.scala 37:46:@5276.4]
  assign _T_58853 = $signed(_T_58852); // @[Modules.scala 37:46:@5277.4]
  assign _T_58854 = $signed(io_in_522) + $signed(io_in_523); // @[Modules.scala 37:46:@5279.4]
  assign _T_58855 = _T_58854[4:0]; // @[Modules.scala 37:46:@5280.4]
  assign _T_58856 = $signed(_T_58855); // @[Modules.scala 37:46:@5281.4]
  assign _T_58857 = $signed(io_in_524) + $signed(io_in_525); // @[Modules.scala 37:46:@5283.4]
  assign _T_58858 = _T_58857[4:0]; // @[Modules.scala 37:46:@5284.4]
  assign _T_58859 = $signed(_T_58858); // @[Modules.scala 37:46:@5285.4]
  assign _T_58860 = $signed(io_in_526) - $signed(io_in_527); // @[Modules.scala 40:46:@5287.4]
  assign _T_58861 = _T_58860[4:0]; // @[Modules.scala 40:46:@5288.4]
  assign _T_58862 = $signed(_T_58861); // @[Modules.scala 40:46:@5289.4]
  assign _T_58864 = $signed(5'sh0) - $signed(io_in_528); // @[Modules.scala 46:37:@5291.4]
  assign _T_58865 = _T_58864[4:0]; // @[Modules.scala 46:37:@5292.4]
  assign _T_58866 = $signed(_T_58865); // @[Modules.scala 46:37:@5293.4]
  assign _T_58867 = $signed(_T_58866) - $signed(io_in_529); // @[Modules.scala 46:47:@5294.4]
  assign _T_58868 = _T_58867[4:0]; // @[Modules.scala 46:47:@5295.4]
  assign _T_58869 = $signed(_T_58868); // @[Modules.scala 46:47:@5296.4]
  assign _T_58877 = $signed(io_in_532) + $signed(io_in_533); // @[Modules.scala 37:46:@5305.4]
  assign _T_58878 = _T_58877[4:0]; // @[Modules.scala 37:46:@5306.4]
  assign _T_58879 = $signed(_T_58878); // @[Modules.scala 37:46:@5307.4]
  assign _T_58880 = $signed(io_in_534) + $signed(io_in_535); // @[Modules.scala 37:46:@5309.4]
  assign _T_58881 = _T_58880[4:0]; // @[Modules.scala 37:46:@5310.4]
  assign _T_58882 = $signed(_T_58881); // @[Modules.scala 37:46:@5311.4]
  assign _T_58883 = $signed(io_in_536) + $signed(io_in_537); // @[Modules.scala 37:46:@5313.4]
  assign _T_58884 = _T_58883[4:0]; // @[Modules.scala 37:46:@5314.4]
  assign _T_58885 = $signed(_T_58884); // @[Modules.scala 37:46:@5315.4]
  assign _T_58886 = $signed(io_in_538) + $signed(io_in_539); // @[Modules.scala 37:46:@5317.4]
  assign _T_58887 = _T_58886[4:0]; // @[Modules.scala 37:46:@5318.4]
  assign _T_58888 = $signed(_T_58887); // @[Modules.scala 37:46:@5319.4]
  assign _T_58889 = $signed(io_in_540) + $signed(io_in_541); // @[Modules.scala 37:46:@5321.4]
  assign _T_58890 = _T_58889[4:0]; // @[Modules.scala 37:46:@5322.4]
  assign _T_58891 = $signed(_T_58890); // @[Modules.scala 37:46:@5323.4]
  assign _T_58892 = $signed(io_in_542) + $signed(io_in_543); // @[Modules.scala 37:46:@5325.4]
  assign _T_58893 = _T_58892[4:0]; // @[Modules.scala 37:46:@5326.4]
  assign _T_58894 = $signed(_T_58893); // @[Modules.scala 37:46:@5327.4]
  assign _T_58895 = $signed(io_in_544) + $signed(io_in_545); // @[Modules.scala 37:46:@5329.4]
  assign _T_58896 = _T_58895[4:0]; // @[Modules.scala 37:46:@5330.4]
  assign _T_58897 = $signed(_T_58896); // @[Modules.scala 37:46:@5331.4]
  assign _T_58902 = $signed(_T_55756) + $signed(io_in_547); // @[Modules.scala 43:47:@5336.4]
  assign _T_58903 = _T_58902[4:0]; // @[Modules.scala 43:47:@5337.4]
  assign _T_58904 = $signed(_T_58903); // @[Modules.scala 43:47:@5338.4]
  assign _T_58905 = $signed(io_in_548) + $signed(io_in_549); // @[Modules.scala 37:46:@5340.4]
  assign _T_58906 = _T_58905[4:0]; // @[Modules.scala 37:46:@5341.4]
  assign _T_58907 = $signed(_T_58906); // @[Modules.scala 37:46:@5342.4]
  assign _T_58908 = $signed(io_in_550) + $signed(io_in_551); // @[Modules.scala 37:46:@5344.4]
  assign _T_58909 = _T_58908[4:0]; // @[Modules.scala 37:46:@5345.4]
  assign _T_58910 = $signed(_T_58909); // @[Modules.scala 37:46:@5346.4]
  assign _T_58914 = $signed(io_in_554) - $signed(io_in_555); // @[Modules.scala 40:46:@5352.4]
  assign _T_58915 = _T_58914[4:0]; // @[Modules.scala 40:46:@5353.4]
  assign _T_58916 = $signed(_T_58915); // @[Modules.scala 40:46:@5354.4]
  assign _T_58918 = $signed(5'sh0) - $signed(io_in_556); // @[Modules.scala 46:37:@5356.4]
  assign _T_58919 = _T_58918[4:0]; // @[Modules.scala 46:37:@5357.4]
  assign _T_58920 = $signed(_T_58919); // @[Modules.scala 46:37:@5358.4]
  assign _T_58921 = $signed(_T_58920) - $signed(io_in_557); // @[Modules.scala 46:47:@5359.4]
  assign _T_58922 = _T_58921[4:0]; // @[Modules.scala 46:47:@5360.4]
  assign _T_58923 = $signed(_T_58922); // @[Modules.scala 46:47:@5361.4]
  assign _T_58928 = $signed(_T_55786) - $signed(io_in_559); // @[Modules.scala 46:47:@5366.4]
  assign _T_58929 = _T_58928[4:0]; // @[Modules.scala 46:47:@5367.4]
  assign _T_58930 = $signed(_T_58929); // @[Modules.scala 46:47:@5368.4]
  assign _T_58935 = $signed(_T_55793) + $signed(io_in_561); // @[Modules.scala 43:47:@5373.4]
  assign _T_58936 = _T_58935[4:0]; // @[Modules.scala 43:47:@5374.4]
  assign _T_58937 = $signed(_T_58936); // @[Modules.scala 43:47:@5375.4]
  assign _T_58938 = $signed(io_in_562) + $signed(io_in_563); // @[Modules.scala 37:46:@5377.4]
  assign _T_58939 = _T_58938[4:0]; // @[Modules.scala 37:46:@5378.4]
  assign _T_58940 = $signed(_T_58939); // @[Modules.scala 37:46:@5379.4]
  assign _T_58941 = $signed(io_in_564) + $signed(io_in_565); // @[Modules.scala 37:46:@5381.4]
  assign _T_58942 = _T_58941[4:0]; // @[Modules.scala 37:46:@5382.4]
  assign _T_58943 = $signed(_T_58942); // @[Modules.scala 37:46:@5383.4]
  assign _T_58944 = $signed(io_in_566) - $signed(io_in_567); // @[Modules.scala 40:46:@5385.4]
  assign _T_58945 = _T_58944[4:0]; // @[Modules.scala 40:46:@5386.4]
  assign _T_58946 = $signed(_T_58945); // @[Modules.scala 40:46:@5387.4]
  assign _T_58947 = $signed(io_in_568) + $signed(io_in_569); // @[Modules.scala 37:46:@5389.4]
  assign _T_58948 = _T_58947[4:0]; // @[Modules.scala 37:46:@5390.4]
  assign _T_58949 = $signed(_T_58948); // @[Modules.scala 37:46:@5391.4]
  assign _T_58950 = $signed(io_in_570) + $signed(io_in_571); // @[Modules.scala 37:46:@5393.4]
  assign _T_58951 = _T_58950[4:0]; // @[Modules.scala 37:46:@5394.4]
  assign _T_58952 = $signed(_T_58951); // @[Modules.scala 37:46:@5395.4]
  assign _T_58953 = $signed(io_in_572) + $signed(io_in_573); // @[Modules.scala 37:46:@5397.4]
  assign _T_58954 = _T_58953[4:0]; // @[Modules.scala 37:46:@5398.4]
  assign _T_58955 = $signed(_T_58954); // @[Modules.scala 37:46:@5399.4]
  assign _T_58956 = $signed(io_in_574) + $signed(io_in_575); // @[Modules.scala 37:46:@5401.4]
  assign _T_58957 = _T_58956[4:0]; // @[Modules.scala 37:46:@5402.4]
  assign _T_58958 = $signed(_T_58957); // @[Modules.scala 37:46:@5403.4]
  assign _T_58959 = $signed(io_in_576) - $signed(io_in_577); // @[Modules.scala 40:46:@5405.4]
  assign _T_58960 = _T_58959[4:0]; // @[Modules.scala 40:46:@5406.4]
  assign _T_58961 = $signed(_T_58960); // @[Modules.scala 40:46:@5407.4]
  assign _T_58962 = $signed(io_in_578) + $signed(io_in_579); // @[Modules.scala 37:46:@5409.4]
  assign _T_58963 = _T_58962[4:0]; // @[Modules.scala 37:46:@5410.4]
  assign _T_58964 = $signed(_T_58963); // @[Modules.scala 37:46:@5411.4]
  assign _T_58968 = $signed(io_in_582) - $signed(io_in_583); // @[Modules.scala 40:46:@5417.4]
  assign _T_58969 = _T_58968[4:0]; // @[Modules.scala 40:46:@5418.4]
  assign _T_58970 = $signed(_T_58969); // @[Modules.scala 40:46:@5419.4]
  assign _T_58972 = $signed(5'sh0) - $signed(io_in_584); // @[Modules.scala 46:37:@5421.4]
  assign _T_58973 = _T_58972[4:0]; // @[Modules.scala 46:37:@5422.4]
  assign _T_58974 = $signed(_T_58973); // @[Modules.scala 46:37:@5423.4]
  assign _T_58975 = $signed(_T_58974) - $signed(io_in_585); // @[Modules.scala 46:47:@5424.4]
  assign _T_58976 = _T_58975[4:0]; // @[Modules.scala 46:47:@5425.4]
  assign _T_58977 = $signed(_T_58976); // @[Modules.scala 46:47:@5426.4]
  assign _T_58989 = $signed(_T_55875) - $signed(io_in_589); // @[Modules.scala 46:47:@5438.4]
  assign _T_58990 = _T_58989[4:0]; // @[Modules.scala 46:47:@5439.4]
  assign _T_58991 = $signed(_T_58990); // @[Modules.scala 46:47:@5440.4]
  assign _T_58992 = $signed(io_in_590) + $signed(io_in_591); // @[Modules.scala 37:46:@5442.4]
  assign _T_58993 = _T_58992[4:0]; // @[Modules.scala 37:46:@5443.4]
  assign _T_58994 = $signed(_T_58993); // @[Modules.scala 37:46:@5444.4]
  assign _T_58995 = $signed(io_in_592) + $signed(io_in_593); // @[Modules.scala 37:46:@5446.4]
  assign _T_58996 = _T_58995[4:0]; // @[Modules.scala 37:46:@5447.4]
  assign _T_58997 = $signed(_T_58996); // @[Modules.scala 37:46:@5448.4]
  assign _T_58998 = $signed(io_in_594) - $signed(io_in_595); // @[Modules.scala 40:46:@5450.4]
  assign _T_58999 = _T_58998[4:0]; // @[Modules.scala 40:46:@5451.4]
  assign _T_59000 = $signed(_T_58999); // @[Modules.scala 40:46:@5452.4]
  assign _T_59001 = $signed(io_in_596) - $signed(io_in_597); // @[Modules.scala 40:46:@5454.4]
  assign _T_59002 = _T_59001[4:0]; // @[Modules.scala 40:46:@5455.4]
  assign _T_59003 = $signed(_T_59002); // @[Modules.scala 40:46:@5456.4]
  assign _T_59004 = $signed(io_in_598) + $signed(io_in_599); // @[Modules.scala 37:46:@5458.4]
  assign _T_59005 = _T_59004[4:0]; // @[Modules.scala 37:46:@5459.4]
  assign _T_59006 = $signed(_T_59005); // @[Modules.scala 37:46:@5460.4]
  assign _T_59010 = $signed(io_in_602) + $signed(io_in_603); // @[Modules.scala 37:46:@5466.4]
  assign _T_59011 = _T_59010[4:0]; // @[Modules.scala 37:46:@5467.4]
  assign _T_59012 = $signed(_T_59011); // @[Modules.scala 37:46:@5468.4]
  assign _T_59034 = $signed(5'sh0) - $signed(io_in_612); // @[Modules.scala 46:37:@5492.4]
  assign _T_59035 = _T_59034[4:0]; // @[Modules.scala 46:37:@5493.4]
  assign _T_59036 = $signed(_T_59035); // @[Modules.scala 46:37:@5494.4]
  assign _T_59037 = $signed(_T_59036) - $signed(io_in_613); // @[Modules.scala 46:47:@5495.4]
  assign _T_59038 = _T_59037[4:0]; // @[Modules.scala 46:47:@5496.4]
  assign _T_59039 = $signed(_T_59038); // @[Modules.scala 46:47:@5497.4]
  assign _T_59051 = $signed(_T_55953) - $signed(io_in_617); // @[Modules.scala 46:47:@5509.4]
  assign _T_59052 = _T_59051[4:0]; // @[Modules.scala 46:47:@5510.4]
  assign _T_59053 = $signed(_T_59052); // @[Modules.scala 46:47:@5511.4]
  assign _T_59057 = $signed(io_in_620) - $signed(io_in_621); // @[Modules.scala 40:46:@5517.4]
  assign _T_59058 = _T_59057[4:0]; // @[Modules.scala 40:46:@5518.4]
  assign _T_59059 = $signed(_T_59058); // @[Modules.scala 40:46:@5519.4]
  assign _T_59067 = $signed(io_in_624) + $signed(io_in_625); // @[Modules.scala 37:46:@5528.4]
  assign _T_59068 = _T_59067[4:0]; // @[Modules.scala 37:46:@5529.4]
  assign _T_59069 = $signed(_T_59068); // @[Modules.scala 37:46:@5530.4]
  assign _T_59070 = $signed(io_in_626) + $signed(io_in_627); // @[Modules.scala 37:46:@5532.4]
  assign _T_59071 = _T_59070[4:0]; // @[Modules.scala 37:46:@5533.4]
  assign _T_59072 = $signed(_T_59071); // @[Modules.scala 37:46:@5534.4]
  assign _T_59073 = $signed(io_in_628) + $signed(io_in_629); // @[Modules.scala 37:46:@5536.4]
  assign _T_59074 = _T_59073[4:0]; // @[Modules.scala 37:46:@5537.4]
  assign _T_59075 = $signed(_T_59074); // @[Modules.scala 37:46:@5538.4]
  assign _T_59076 = $signed(io_in_630) + $signed(io_in_631); // @[Modules.scala 37:46:@5540.4]
  assign _T_59077 = _T_59076[4:0]; // @[Modules.scala 37:46:@5541.4]
  assign _T_59078 = $signed(_T_59077); // @[Modules.scala 37:46:@5542.4]
  assign _T_59079 = $signed(io_in_632) + $signed(io_in_633); // @[Modules.scala 37:46:@5544.4]
  assign _T_59080 = _T_59079[4:0]; // @[Modules.scala 37:46:@5545.4]
  assign _T_59081 = $signed(_T_59080); // @[Modules.scala 37:46:@5546.4]
  assign _T_59082 = $signed(io_in_634) - $signed(io_in_635); // @[Modules.scala 40:46:@5548.4]
  assign _T_59083 = _T_59082[4:0]; // @[Modules.scala 40:46:@5549.4]
  assign _T_59084 = $signed(_T_59083); // @[Modules.scala 40:46:@5550.4]
  assign _T_59085 = $signed(io_in_636) + $signed(io_in_637); // @[Modules.scala 37:46:@5552.4]
  assign _T_59086 = _T_59085[4:0]; // @[Modules.scala 37:46:@5553.4]
  assign _T_59087 = $signed(_T_59086); // @[Modules.scala 37:46:@5554.4]
  assign _T_59088 = $signed(io_in_638) - $signed(io_in_639); // @[Modules.scala 40:46:@5556.4]
  assign _T_59089 = _T_59088[4:0]; // @[Modules.scala 40:46:@5557.4]
  assign _T_59090 = $signed(_T_59089); // @[Modules.scala 40:46:@5558.4]
  assign _T_59092 = $signed(5'sh0) - $signed(io_in_640); // @[Modules.scala 46:37:@5560.4]
  assign _T_59093 = _T_59092[4:0]; // @[Modules.scala 46:37:@5561.4]
  assign _T_59094 = $signed(_T_59093); // @[Modules.scala 46:37:@5562.4]
  assign _T_59095 = $signed(_T_59094) - $signed(io_in_641); // @[Modules.scala 46:47:@5563.4]
  assign _T_59096 = _T_59095[4:0]; // @[Modules.scala 46:47:@5564.4]
  assign _T_59097 = $signed(_T_59096); // @[Modules.scala 46:47:@5565.4]
  assign _T_59098 = $signed(io_in_642) + $signed(io_in_643); // @[Modules.scala 37:46:@5567.4]
  assign _T_59099 = _T_59098[4:0]; // @[Modules.scala 37:46:@5568.4]
  assign _T_59100 = $signed(_T_59099); // @[Modules.scala 37:46:@5569.4]
  assign _T_59105 = $signed(_T_56043) - $signed(io_in_645); // @[Modules.scala 46:47:@5574.4]
  assign _T_59106 = _T_59105[4:0]; // @[Modules.scala 46:47:@5575.4]
  assign _T_59107 = $signed(_T_59106); // @[Modules.scala 46:47:@5576.4]
  assign _T_59111 = $signed(io_in_648) + $signed(io_in_649); // @[Modules.scala 37:46:@5582.4]
  assign _T_59112 = _T_59111[4:0]; // @[Modules.scala 37:46:@5583.4]
  assign _T_59113 = $signed(_T_59112); // @[Modules.scala 37:46:@5584.4]
  assign _T_59114 = $signed(io_in_650) + $signed(io_in_651); // @[Modules.scala 37:46:@5586.4]
  assign _T_59115 = _T_59114[4:0]; // @[Modules.scala 37:46:@5587.4]
  assign _T_59116 = $signed(_T_59115); // @[Modules.scala 37:46:@5588.4]
  assign _T_59117 = $signed(io_in_652) + $signed(io_in_653); // @[Modules.scala 37:46:@5590.4]
  assign _T_59118 = _T_59117[4:0]; // @[Modules.scala 37:46:@5591.4]
  assign _T_59119 = $signed(_T_59118); // @[Modules.scala 37:46:@5592.4]
  assign _T_59120 = $signed(io_in_654) + $signed(io_in_655); // @[Modules.scala 37:46:@5594.4]
  assign _T_59121 = _T_59120[4:0]; // @[Modules.scala 37:46:@5595.4]
  assign _T_59122 = $signed(_T_59121); // @[Modules.scala 37:46:@5596.4]
  assign _T_59123 = $signed(io_in_656) + $signed(io_in_657); // @[Modules.scala 37:46:@5598.4]
  assign _T_59124 = _T_59123[4:0]; // @[Modules.scala 37:46:@5599.4]
  assign _T_59125 = $signed(_T_59124); // @[Modules.scala 37:46:@5600.4]
  assign _T_59126 = $signed(io_in_658) + $signed(io_in_659); // @[Modules.scala 37:46:@5602.4]
  assign _T_59127 = _T_59126[4:0]; // @[Modules.scala 37:46:@5603.4]
  assign _T_59128 = $signed(_T_59127); // @[Modules.scala 37:46:@5604.4]
  assign _T_59136 = $signed(io_in_662) + $signed(io_in_663); // @[Modules.scala 37:46:@5613.4]
  assign _T_59137 = _T_59136[4:0]; // @[Modules.scala 37:46:@5614.4]
  assign _T_59138 = $signed(_T_59137); // @[Modules.scala 37:46:@5615.4]
  assign _T_59140 = $signed(5'sh0) - $signed(io_in_664); // @[Modules.scala 46:37:@5617.4]
  assign _T_59141 = _T_59140[4:0]; // @[Modules.scala 46:37:@5618.4]
  assign _T_59142 = $signed(_T_59141); // @[Modules.scala 46:37:@5619.4]
  assign _T_59143 = $signed(_T_59142) - $signed(io_in_665); // @[Modules.scala 46:47:@5620.4]
  assign _T_59144 = _T_59143[4:0]; // @[Modules.scala 46:47:@5621.4]
  assign _T_59145 = $signed(_T_59144); // @[Modules.scala 46:47:@5622.4]
  assign _T_59147 = $signed(5'sh0) - $signed(io_in_666); // @[Modules.scala 46:37:@5624.4]
  assign _T_59148 = _T_59147[4:0]; // @[Modules.scala 46:37:@5625.4]
  assign _T_59149 = $signed(_T_59148); // @[Modules.scala 46:37:@5626.4]
  assign _T_59150 = $signed(_T_59149) - $signed(io_in_667); // @[Modules.scala 46:47:@5627.4]
  assign _T_59151 = _T_59150[4:0]; // @[Modules.scala 46:47:@5628.4]
  assign _T_59152 = $signed(_T_59151); // @[Modules.scala 46:47:@5629.4]
  assign _T_59154 = $signed(5'sh0) - $signed(io_in_668); // @[Modules.scala 46:37:@5631.4]
  assign _T_59155 = _T_59154[4:0]; // @[Modules.scala 46:37:@5632.4]
  assign _T_59156 = $signed(_T_59155); // @[Modules.scala 46:37:@5633.4]
  assign _T_59157 = $signed(_T_59156) - $signed(io_in_669); // @[Modules.scala 46:47:@5634.4]
  assign _T_59158 = _T_59157[4:0]; // @[Modules.scala 46:47:@5635.4]
  assign _T_59159 = $signed(_T_59158); // @[Modules.scala 46:47:@5636.4]
  assign _T_59171 = $signed(_T_56125) - $signed(io_in_673); // @[Modules.scala 46:47:@5648.4]
  assign _T_59172 = _T_59171[4:0]; // @[Modules.scala 46:47:@5649.4]
  assign _T_59173 = $signed(_T_59172); // @[Modules.scala 46:47:@5650.4]
  assign _T_59174 = $signed(io_in_674) + $signed(io_in_675); // @[Modules.scala 37:46:@5652.4]
  assign _T_59175 = _T_59174[4:0]; // @[Modules.scala 37:46:@5653.4]
  assign _T_59176 = $signed(_T_59175); // @[Modules.scala 37:46:@5654.4]
  assign _T_59184 = $signed(5'sh0) - $signed(io_in_680); // @[Modules.scala 43:37:@5664.4]
  assign _T_59185 = _T_59184[4:0]; // @[Modules.scala 43:37:@5665.4]
  assign _T_59186 = $signed(_T_59185); // @[Modules.scala 43:37:@5666.4]
  assign _T_59187 = $signed(_T_59186) + $signed(io_in_681); // @[Modules.scala 43:47:@5667.4]
  assign _T_59188 = _T_59187[4:0]; // @[Modules.scala 43:47:@5668.4]
  assign _T_59189 = $signed(_T_59188); // @[Modules.scala 43:47:@5669.4]
  assign _T_59190 = $signed(io_in_682) + $signed(io_in_683); // @[Modules.scala 37:46:@5671.4]
  assign _T_59191 = _T_59190[4:0]; // @[Modules.scala 37:46:@5672.4]
  assign _T_59192 = $signed(_T_59191); // @[Modules.scala 37:46:@5673.4]
  assign _T_59193 = $signed(io_in_684) + $signed(io_in_685); // @[Modules.scala 37:46:@5675.4]
  assign _T_59194 = _T_59193[4:0]; // @[Modules.scala 37:46:@5676.4]
  assign _T_59195 = $signed(_T_59194); // @[Modules.scala 37:46:@5677.4]
  assign _T_59196 = $signed(io_in_686) - $signed(io_in_687); // @[Modules.scala 40:46:@5679.4]
  assign _T_59197 = _T_59196[4:0]; // @[Modules.scala 40:46:@5680.4]
  assign _T_59198 = $signed(_T_59197); // @[Modules.scala 40:46:@5681.4]
  assign _T_59199 = $signed(io_in_688) - $signed(io_in_689); // @[Modules.scala 40:46:@5683.4]
  assign _T_59200 = _T_59199[4:0]; // @[Modules.scala 40:46:@5684.4]
  assign _T_59201 = $signed(_T_59200); // @[Modules.scala 40:46:@5685.4]
  assign _T_59202 = $signed(io_in_690) - $signed(io_in_691); // @[Modules.scala 40:46:@5687.4]
  assign _T_59203 = _T_59202[4:0]; // @[Modules.scala 40:46:@5688.4]
  assign _T_59204 = $signed(_T_59203); // @[Modules.scala 40:46:@5689.4]
  assign _T_59206 = $signed(5'sh0) - $signed(io_in_692); // @[Modules.scala 46:37:@5691.4]
  assign _T_59207 = _T_59206[4:0]; // @[Modules.scala 46:37:@5692.4]
  assign _T_59208 = $signed(_T_59207); // @[Modules.scala 46:37:@5693.4]
  assign _T_59209 = $signed(_T_59208) - $signed(io_in_693); // @[Modules.scala 46:47:@5694.4]
  assign _T_59210 = _T_59209[4:0]; // @[Modules.scala 46:47:@5695.4]
  assign _T_59211 = $signed(_T_59210); // @[Modules.scala 46:47:@5696.4]
  assign _T_59213 = $signed(5'sh0) - $signed(io_in_694); // @[Modules.scala 43:37:@5698.4]
  assign _T_59214 = _T_59213[4:0]; // @[Modules.scala 43:37:@5699.4]
  assign _T_59215 = $signed(_T_59214); // @[Modules.scala 43:37:@5700.4]
  assign _T_59216 = $signed(_T_59215) + $signed(io_in_695); // @[Modules.scala 43:47:@5701.4]
  assign _T_59217 = _T_59216[4:0]; // @[Modules.scala 43:47:@5702.4]
  assign _T_59218 = $signed(_T_59217); // @[Modules.scala 43:47:@5703.4]
  assign _T_59219 = $signed(io_in_696) - $signed(io_in_697); // @[Modules.scala 40:46:@5705.4]
  assign _T_59220 = _T_59219[4:0]; // @[Modules.scala 40:46:@5706.4]
  assign _T_59221 = $signed(_T_59220); // @[Modules.scala 40:46:@5707.4]
  assign _T_59226 = $signed(_T_56176) - $signed(io_in_699); // @[Modules.scala 46:47:@5712.4]
  assign _T_59227 = _T_59226[4:0]; // @[Modules.scala 46:47:@5713.4]
  assign _T_59228 = $signed(_T_59227); // @[Modules.scala 46:47:@5714.4]
  assign _T_59229 = $signed(io_in_700) + $signed(io_in_701); // @[Modules.scala 37:46:@5716.4]
  assign _T_59230 = _T_59229[4:0]; // @[Modules.scala 37:46:@5717.4]
  assign _T_59231 = $signed(_T_59230); // @[Modules.scala 37:46:@5718.4]
  assign _T_59232 = $signed(io_in_702) + $signed(io_in_703); // @[Modules.scala 37:46:@5720.4]
  assign _T_59233 = _T_59232[4:0]; // @[Modules.scala 37:46:@5721.4]
  assign _T_59234 = $signed(_T_59233); // @[Modules.scala 37:46:@5722.4]
  assign _T_59242 = $signed(5'sh0) - $signed(io_in_708); // @[Modules.scala 46:37:@5732.4]
  assign _T_59243 = _T_59242[4:0]; // @[Modules.scala 46:37:@5733.4]
  assign _T_59244 = $signed(_T_59243); // @[Modules.scala 46:37:@5734.4]
  assign _T_59245 = $signed(_T_59244) - $signed(io_in_709); // @[Modules.scala 46:47:@5735.4]
  assign _T_59246 = _T_59245[4:0]; // @[Modules.scala 46:47:@5736.4]
  assign _T_59247 = $signed(_T_59246); // @[Modules.scala 46:47:@5737.4]
  assign _T_59249 = $signed(5'sh0) - $signed(io_in_710); // @[Modules.scala 43:37:@5739.4]
  assign _T_59250 = _T_59249[4:0]; // @[Modules.scala 43:37:@5740.4]
  assign _T_59251 = $signed(_T_59250); // @[Modules.scala 43:37:@5741.4]
  assign _T_59252 = $signed(_T_59251) + $signed(io_in_711); // @[Modules.scala 43:47:@5742.4]
  assign _T_59253 = _T_59252[4:0]; // @[Modules.scala 43:47:@5743.4]
  assign _T_59254 = $signed(_T_59253); // @[Modules.scala 43:47:@5744.4]
  assign _T_59256 = $signed(5'sh0) - $signed(io_in_712); // @[Modules.scala 46:37:@5746.4]
  assign _T_59257 = _T_59256[4:0]; // @[Modules.scala 46:37:@5747.4]
  assign _T_59258 = $signed(_T_59257); // @[Modules.scala 46:37:@5748.4]
  assign _T_59259 = $signed(_T_59258) - $signed(io_in_713); // @[Modules.scala 46:47:@5749.4]
  assign _T_59260 = _T_59259[4:0]; // @[Modules.scala 46:47:@5750.4]
  assign _T_59261 = $signed(_T_59260); // @[Modules.scala 46:47:@5751.4]
  assign _T_59263 = $signed(5'sh0) - $signed(io_in_714); // @[Modules.scala 43:37:@5753.4]
  assign _T_59264 = _T_59263[4:0]; // @[Modules.scala 43:37:@5754.4]
  assign _T_59265 = $signed(_T_59264); // @[Modules.scala 43:37:@5755.4]
  assign _T_59266 = $signed(_T_59265) + $signed(io_in_715); // @[Modules.scala 43:47:@5756.4]
  assign _T_59267 = _T_59266[4:0]; // @[Modules.scala 43:47:@5757.4]
  assign _T_59268 = $signed(_T_59267); // @[Modules.scala 43:47:@5758.4]
  assign _T_59269 = $signed(io_in_716) - $signed(io_in_717); // @[Modules.scala 40:46:@5760.4]
  assign _T_59270 = _T_59269[4:0]; // @[Modules.scala 40:46:@5761.4]
  assign _T_59271 = $signed(_T_59270); // @[Modules.scala 40:46:@5762.4]
  assign _T_59273 = $signed(5'sh0) - $signed(io_in_718); // @[Modules.scala 46:37:@5764.4]
  assign _T_59274 = _T_59273[4:0]; // @[Modules.scala 46:37:@5765.4]
  assign _T_59275 = $signed(_T_59274); // @[Modules.scala 46:37:@5766.4]
  assign _T_59276 = $signed(_T_59275) - $signed(io_in_719); // @[Modules.scala 46:47:@5767.4]
  assign _T_59277 = _T_59276[4:0]; // @[Modules.scala 46:47:@5768.4]
  assign _T_59278 = $signed(_T_59277); // @[Modules.scala 46:47:@5769.4]
  assign _T_59280 = $signed(5'sh0) - $signed(io_in_720); // @[Modules.scala 46:37:@5771.4]
  assign _T_59281 = _T_59280[4:0]; // @[Modules.scala 46:37:@5772.4]
  assign _T_59282 = $signed(_T_59281); // @[Modules.scala 46:37:@5773.4]
  assign _T_59283 = $signed(_T_59282) - $signed(io_in_721); // @[Modules.scala 46:47:@5774.4]
  assign _T_59284 = _T_59283[4:0]; // @[Modules.scala 46:47:@5775.4]
  assign _T_59285 = $signed(_T_59284); // @[Modules.scala 46:47:@5776.4]
  assign _T_59289 = $signed(io_in_724) + $signed(io_in_725); // @[Modules.scala 37:46:@5782.4]
  assign _T_59290 = _T_59289[4:0]; // @[Modules.scala 37:46:@5783.4]
  assign _T_59291 = $signed(_T_59290); // @[Modules.scala 37:46:@5784.4]
  assign _T_59292 = $signed(io_in_726) - $signed(io_in_727); // @[Modules.scala 40:46:@5786.4]
  assign _T_59293 = _T_59292[4:0]; // @[Modules.scala 40:46:@5787.4]
  assign _T_59294 = $signed(_T_59293); // @[Modules.scala 40:46:@5788.4]
  assign _T_59296 = $signed(5'sh0) - $signed(io_in_728); // @[Modules.scala 46:37:@5790.4]
  assign _T_59297 = _T_59296[4:0]; // @[Modules.scala 46:37:@5791.4]
  assign _T_59298 = $signed(_T_59297); // @[Modules.scala 46:37:@5792.4]
  assign _T_59299 = $signed(_T_59298) - $signed(io_in_729); // @[Modules.scala 46:47:@5793.4]
  assign _T_59300 = _T_59299[4:0]; // @[Modules.scala 46:47:@5794.4]
  assign _T_59301 = $signed(_T_59300); // @[Modules.scala 46:47:@5795.4]
  assign _T_59306 = $signed(_T_56236) - $signed(io_in_731); // @[Modules.scala 46:47:@5800.4]
  assign _T_59307 = _T_59306[4:0]; // @[Modules.scala 46:47:@5801.4]
  assign _T_59308 = $signed(_T_59307); // @[Modules.scala 46:47:@5802.4]
  assign _T_59310 = $signed(5'sh0) - $signed(io_in_732); // @[Modules.scala 46:37:@5804.4]
  assign _T_59311 = _T_59310[4:0]; // @[Modules.scala 46:37:@5805.4]
  assign _T_59312 = $signed(_T_59311); // @[Modules.scala 46:37:@5806.4]
  assign _T_59313 = $signed(_T_59312) - $signed(io_in_733); // @[Modules.scala 46:47:@5807.4]
  assign _T_59314 = _T_59313[4:0]; // @[Modules.scala 46:47:@5808.4]
  assign _T_59315 = $signed(_T_59314); // @[Modules.scala 46:47:@5809.4]
  assign _T_59317 = $signed(5'sh0) - $signed(io_in_734); // @[Modules.scala 46:37:@5811.4]
  assign _T_59318 = _T_59317[4:0]; // @[Modules.scala 46:37:@5812.4]
  assign _T_59319 = $signed(_T_59318); // @[Modules.scala 46:37:@5813.4]
  assign _T_59320 = $signed(_T_59319) - $signed(io_in_735); // @[Modules.scala 46:47:@5814.4]
  assign _T_59321 = _T_59320[4:0]; // @[Modules.scala 46:47:@5815.4]
  assign _T_59322 = $signed(_T_59321); // @[Modules.scala 46:47:@5816.4]
  assign _T_59338 = $signed(5'sh0) - $signed(io_in_740); // @[Modules.scala 46:37:@5832.4]
  assign _T_59339 = _T_59338[4:0]; // @[Modules.scala 46:37:@5833.4]
  assign _T_59340 = $signed(_T_59339); // @[Modules.scala 46:37:@5834.4]
  assign _T_59341 = $signed(_T_59340) - $signed(io_in_741); // @[Modules.scala 46:47:@5835.4]
  assign _T_59342 = _T_59341[4:0]; // @[Modules.scala 46:47:@5836.4]
  assign _T_59343 = $signed(_T_59342); // @[Modules.scala 46:47:@5837.4]
  assign _T_59345 = $signed(5'sh0) - $signed(io_in_742); // @[Modules.scala 46:37:@5839.4]
  assign _T_59346 = _T_59345[4:0]; // @[Modules.scala 46:37:@5840.4]
  assign _T_59347 = $signed(_T_59346); // @[Modules.scala 46:37:@5841.4]
  assign _T_59348 = $signed(_T_59347) - $signed(io_in_743); // @[Modules.scala 46:47:@5842.4]
  assign _T_59349 = _T_59348[4:0]; // @[Modules.scala 46:47:@5843.4]
  assign _T_59350 = $signed(_T_59349); // @[Modules.scala 46:47:@5844.4]
  assign _T_59377 = $signed(io_in_756) - $signed(io_in_757); // @[Modules.scala 40:46:@5876.4]
  assign _T_59378 = _T_59377[4:0]; // @[Modules.scala 40:46:@5877.4]
  assign _T_59379 = $signed(_T_59378); // @[Modules.scala 40:46:@5878.4]
  assign _T_59380 = $signed(io_in_758) + $signed(io_in_759); // @[Modules.scala 37:46:@5880.4]
  assign _T_59381 = _T_59380[4:0]; // @[Modules.scala 37:46:@5881.4]
  assign _T_59382 = $signed(_T_59381); // @[Modules.scala 37:46:@5882.4]
  assign _T_59383 = $signed(io_in_760) + $signed(io_in_761); // @[Modules.scala 37:46:@5884.4]
  assign _T_59384 = _T_59383[4:0]; // @[Modules.scala 37:46:@5885.4]
  assign _T_59385 = $signed(_T_59384); // @[Modules.scala 37:46:@5886.4]
  assign _T_59386 = $signed(io_in_762) + $signed(io_in_763); // @[Modules.scala 37:46:@5888.4]
  assign _T_59387 = _T_59386[4:0]; // @[Modules.scala 37:46:@5889.4]
  assign _T_59388 = $signed(_T_59387); // @[Modules.scala 37:46:@5890.4]
  assign _T_59396 = $signed(io_in_766) + $signed(io_in_767); // @[Modules.scala 37:46:@5899.4]
  assign _T_59397 = _T_59396[4:0]; // @[Modules.scala 37:46:@5900.4]
  assign _T_59398 = $signed(_T_59397); // @[Modules.scala 37:46:@5901.4]
  assign _T_59400 = $signed(5'sh0) - $signed(io_in_768); // @[Modules.scala 46:37:@5903.4]
  assign _T_59401 = _T_59400[4:0]; // @[Modules.scala 46:37:@5904.4]
  assign _T_59402 = $signed(_T_59401); // @[Modules.scala 46:37:@5905.4]
  assign _T_59403 = $signed(_T_59402) - $signed(io_in_769); // @[Modules.scala 46:47:@5906.4]
  assign _T_59404 = _T_59403[4:0]; // @[Modules.scala 46:47:@5907.4]
  assign _T_59405 = $signed(_T_59404); // @[Modules.scala 46:47:@5908.4]
  assign _T_59410 = $signed(_T_56336) - $signed(io_in_771); // @[Modules.scala 46:47:@5913.4]
  assign _T_59411 = _T_59410[4:0]; // @[Modules.scala 46:47:@5914.4]
  assign _T_59412 = $signed(_T_59411); // @[Modules.scala 46:47:@5915.4]
  assign _T_59428 = $signed(5'sh0) - $signed(io_in_776); // @[Modules.scala 46:37:@5931.4]
  assign _T_59429 = _T_59428[4:0]; // @[Modules.scala 46:37:@5932.4]
  assign _T_59430 = $signed(_T_59429); // @[Modules.scala 46:37:@5933.4]
  assign _T_59431 = $signed(_T_59430) - $signed(io_in_777); // @[Modules.scala 46:47:@5934.4]
  assign _T_59432 = _T_59431[4:0]; // @[Modules.scala 46:47:@5935.4]
  assign _T_59433 = $signed(_T_59432); // @[Modules.scala 46:47:@5936.4]
  assign _T_59441 = $signed(io_in_780) - $signed(io_in_781); // @[Modules.scala 40:46:@5945.4]
  assign _T_59442 = _T_59441[4:0]; // @[Modules.scala 40:46:@5946.4]
  assign _T_59443 = $signed(_T_59442); // @[Modules.scala 40:46:@5947.4]
  assign _T_59445 = $signed(5'sh0) - $signed(io_in_782); // @[Modules.scala 46:37:@5949.4]
  assign _T_59446 = _T_59445[4:0]; // @[Modules.scala 46:37:@5950.4]
  assign _T_59447 = $signed(_T_59446); // @[Modules.scala 46:37:@5951.4]
  assign _T_59448 = $signed(_T_59447) - $signed(io_in_783); // @[Modules.scala 46:47:@5952.4]
  assign _T_59449 = _T_59448[4:0]; // @[Modules.scala 46:47:@5953.4]
  assign _T_59450 = $signed(_T_59449); // @[Modules.scala 46:47:@5954.4]
  assign buffer_1_0 = {{6{_T_57553[4]}},_T_57553}; // @[Modules.scala 32:22:@8.4]
  assign _T_59451 = $signed(buffer_1_0) + $signed(buffer_0_1); // @[Modules.scala 50:57:@5956.4]
  assign _T_59452 = _T_59451[10:0]; // @[Modules.scala 50:57:@5957.4]
  assign buffer_1_392 = $signed(_T_59452); // @[Modules.scala 50:57:@5958.4]
  assign buffer_1_2 = {{6{_T_57563[4]}},_T_57563}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_3 = {{6{_T_57566[4]}},_T_57566}; // @[Modules.scala 32:22:@8.4]
  assign _T_59454 = $signed(buffer_1_2) + $signed(buffer_1_3); // @[Modules.scala 50:57:@5960.4]
  assign _T_59455 = _T_59454[10:0]; // @[Modules.scala 50:57:@5961.4]
  assign buffer_1_393 = $signed(_T_59455); // @[Modules.scala 50:57:@5962.4]
  assign buffer_1_4 = {{6{_T_57569[4]}},_T_57569}; // @[Modules.scala 32:22:@8.4]
  assign _T_59457 = $signed(buffer_1_4) + $signed(buffer_0_5); // @[Modules.scala 50:57:@5964.4]
  assign _T_59458 = _T_59457[10:0]; // @[Modules.scala 50:57:@5965.4]
  assign buffer_1_394 = $signed(_T_59458); // @[Modules.scala 50:57:@5966.4]
  assign buffer_1_6 = {{6{_T_57579[4]}},_T_57579}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_7 = {{6{_T_57582[4]}},_T_57582}; // @[Modules.scala 32:22:@8.4]
  assign _T_59460 = $signed(buffer_1_6) + $signed(buffer_1_7); // @[Modules.scala 50:57:@5968.4]
  assign _T_59461 = _T_59460[10:0]; // @[Modules.scala 50:57:@5969.4]
  assign buffer_1_395 = $signed(_T_59461); // @[Modules.scala 50:57:@5970.4]
  assign buffer_1_8 = {{6{_T_57585[4]}},_T_57585}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_9 = {{6{_T_57588[4]}},_T_57588}; // @[Modules.scala 32:22:@8.4]
  assign _T_59463 = $signed(buffer_1_8) + $signed(buffer_1_9); // @[Modules.scala 50:57:@5972.4]
  assign _T_59464 = _T_59463[10:0]; // @[Modules.scala 50:57:@5973.4]
  assign buffer_1_396 = $signed(_T_59464); // @[Modules.scala 50:57:@5974.4]
  assign buffer_1_11 = {{6{_T_57594[4]}},_T_57594}; // @[Modules.scala 32:22:@8.4]
  assign _T_59466 = $signed(buffer_0_10) + $signed(buffer_1_11); // @[Modules.scala 50:57:@5976.4]
  assign _T_59467 = _T_59466[10:0]; // @[Modules.scala 50:57:@5977.4]
  assign buffer_1_397 = $signed(_T_59467); // @[Modules.scala 50:57:@5978.4]
  assign buffer_1_12 = {{6{_T_57597[4]}},_T_57597}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_13 = {{6{_T_57604[4]}},_T_57604}; // @[Modules.scala 32:22:@8.4]
  assign _T_59469 = $signed(buffer_1_12) + $signed(buffer_1_13); // @[Modules.scala 50:57:@5980.4]
  assign _T_59470 = _T_59469[10:0]; // @[Modules.scala 50:57:@5981.4]
  assign buffer_1_398 = $signed(_T_59470); // @[Modules.scala 50:57:@5982.4]
  assign buffer_1_14 = {{6{_T_57607[4]}},_T_57607}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_15 = {{6{_T_57610[4]}},_T_57610}; // @[Modules.scala 32:22:@8.4]
  assign _T_59472 = $signed(buffer_1_14) + $signed(buffer_1_15); // @[Modules.scala 50:57:@5984.4]
  assign _T_59473 = _T_59472[10:0]; // @[Modules.scala 50:57:@5985.4]
  assign buffer_1_399 = $signed(_T_59473); // @[Modules.scala 50:57:@5986.4]
  assign buffer_1_17 = {{6{_T_57616[4]}},_T_57616}; // @[Modules.scala 32:22:@8.4]
  assign _T_59475 = $signed(buffer_0_16) + $signed(buffer_1_17); // @[Modules.scala 50:57:@5988.4]
  assign _T_59476 = _T_59475[10:0]; // @[Modules.scala 50:57:@5989.4]
  assign buffer_1_400 = $signed(_T_59476); // @[Modules.scala 50:57:@5990.4]
  assign buffer_1_18 = {{6{_T_57619[4]}},_T_57619}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_19 = {{6{_T_57622[4]}},_T_57622}; // @[Modules.scala 32:22:@8.4]
  assign _T_59478 = $signed(buffer_1_18) + $signed(buffer_1_19); // @[Modules.scala 50:57:@5992.4]
  assign _T_59479 = _T_59478[10:0]; // @[Modules.scala 50:57:@5993.4]
  assign buffer_1_401 = $signed(_T_59479); // @[Modules.scala 50:57:@5994.4]
  assign buffer_1_20 = {{6{_T_57625[4]}},_T_57625}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_21 = {{6{_T_57628[4]}},_T_57628}; // @[Modules.scala 32:22:@8.4]
  assign _T_59481 = $signed(buffer_1_20) + $signed(buffer_1_21); // @[Modules.scala 50:57:@5996.4]
  assign _T_59482 = _T_59481[10:0]; // @[Modules.scala 50:57:@5997.4]
  assign buffer_1_402 = $signed(_T_59482); // @[Modules.scala 50:57:@5998.4]
  assign buffer_1_22 = {{6{_T_57635[4]}},_T_57635}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_23 = {{6{_T_57638[4]}},_T_57638}; // @[Modules.scala 32:22:@8.4]
  assign _T_59484 = $signed(buffer_1_22) + $signed(buffer_1_23); // @[Modules.scala 50:57:@6000.4]
  assign _T_59485 = _T_59484[10:0]; // @[Modules.scala 50:57:@6001.4]
  assign buffer_1_403 = $signed(_T_59485); // @[Modules.scala 50:57:@6002.4]
  assign buffer_1_24 = {{6{_T_57641[4]}},_T_57641}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_25 = {{6{_T_57644[4]}},_T_57644}; // @[Modules.scala 32:22:@8.4]
  assign _T_59487 = $signed(buffer_1_24) + $signed(buffer_1_25); // @[Modules.scala 50:57:@6004.4]
  assign _T_59488 = _T_59487[10:0]; // @[Modules.scala 50:57:@6005.4]
  assign buffer_1_404 = $signed(_T_59488); // @[Modules.scala 50:57:@6006.4]
  assign buffer_1_26 = {{6{_T_57647[4]}},_T_57647}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_27 = {{6{_T_57654[4]}},_T_57654}; // @[Modules.scala 32:22:@8.4]
  assign _T_59490 = $signed(buffer_1_26) + $signed(buffer_1_27); // @[Modules.scala 50:57:@6008.4]
  assign _T_59491 = _T_59490[10:0]; // @[Modules.scala 50:57:@6009.4]
  assign buffer_1_405 = $signed(_T_59491); // @[Modules.scala 50:57:@6010.4]
  assign buffer_1_28 = {{6{_T_57661[4]}},_T_57661}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_29 = {{6{_T_57664[4]}},_T_57664}; // @[Modules.scala 32:22:@8.4]
  assign _T_59493 = $signed(buffer_1_28) + $signed(buffer_1_29); // @[Modules.scala 50:57:@6012.4]
  assign _T_59494 = _T_59493[10:0]; // @[Modules.scala 50:57:@6013.4]
  assign buffer_1_406 = $signed(_T_59494); // @[Modules.scala 50:57:@6014.4]
  assign buffer_1_30 = {{6{_T_57667[4]}},_T_57667}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_31 = {{6{_T_57670[4]}},_T_57670}; // @[Modules.scala 32:22:@8.4]
  assign _T_59496 = $signed(buffer_1_30) + $signed(buffer_1_31); // @[Modules.scala 50:57:@6016.4]
  assign _T_59497 = _T_59496[10:0]; // @[Modules.scala 50:57:@6017.4]
  assign buffer_1_407 = $signed(_T_59497); // @[Modules.scala 50:57:@6018.4]
  assign buffer_1_32 = {{6{_T_57673[4]}},_T_57673}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_33 = {{6{_T_57676[4]}},_T_57676}; // @[Modules.scala 32:22:@8.4]
  assign _T_59499 = $signed(buffer_1_32) + $signed(buffer_1_33); // @[Modules.scala 50:57:@6020.4]
  assign _T_59500 = _T_59499[10:0]; // @[Modules.scala 50:57:@6021.4]
  assign buffer_1_408 = $signed(_T_59500); // @[Modules.scala 50:57:@6022.4]
  assign buffer_1_34 = {{6{_T_57679[4]}},_T_57679}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_35 = {{6{_T_57682[4]}},_T_57682}; // @[Modules.scala 32:22:@8.4]
  assign _T_59502 = $signed(buffer_1_34) + $signed(buffer_1_35); // @[Modules.scala 50:57:@6024.4]
  assign _T_59503 = _T_59502[10:0]; // @[Modules.scala 50:57:@6025.4]
  assign buffer_1_409 = $signed(_T_59503); // @[Modules.scala 50:57:@6026.4]
  assign buffer_1_36 = {{6{_T_57685[4]}},_T_57685}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_37 = {{6{_T_57688[4]}},_T_57688}; // @[Modules.scala 32:22:@8.4]
  assign _T_59505 = $signed(buffer_1_36) + $signed(buffer_1_37); // @[Modules.scala 50:57:@6028.4]
  assign _T_59506 = _T_59505[10:0]; // @[Modules.scala 50:57:@6029.4]
  assign buffer_1_410 = $signed(_T_59506); // @[Modules.scala 50:57:@6030.4]
  assign buffer_1_38 = {{6{_T_57691[4]}},_T_57691}; // @[Modules.scala 32:22:@8.4]
  assign _T_59508 = $signed(buffer_1_38) + $signed(buffer_0_39); // @[Modules.scala 50:57:@6032.4]
  assign _T_59509 = _T_59508[10:0]; // @[Modules.scala 50:57:@6033.4]
  assign buffer_1_411 = $signed(_T_59509); // @[Modules.scala 50:57:@6034.4]
  assign buffer_1_40 = {{6{_T_57697[4]}},_T_57697}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_41 = {{6{_T_57704[4]}},_T_57704}; // @[Modules.scala 32:22:@8.4]
  assign _T_59511 = $signed(buffer_1_40) + $signed(buffer_1_41); // @[Modules.scala 50:57:@6036.4]
  assign _T_59512 = _T_59511[10:0]; // @[Modules.scala 50:57:@6037.4]
  assign buffer_1_412 = $signed(_T_59512); // @[Modules.scala 50:57:@6038.4]
  assign buffer_1_42 = {{6{_T_57711[4]}},_T_57711}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_43 = {{6{_T_57718[4]}},_T_57718}; // @[Modules.scala 32:22:@8.4]
  assign _T_59514 = $signed(buffer_1_42) + $signed(buffer_1_43); // @[Modules.scala 50:57:@6040.4]
  assign _T_59515 = _T_59514[10:0]; // @[Modules.scala 50:57:@6041.4]
  assign buffer_1_413 = $signed(_T_59515); // @[Modules.scala 50:57:@6042.4]
  assign buffer_1_46 = {{6{_T_57727[4]}},_T_57727}; // @[Modules.scala 32:22:@8.4]
  assign _T_59520 = $signed(buffer_1_46) + $signed(buffer_0_47); // @[Modules.scala 50:57:@6048.4]
  assign _T_59521 = _T_59520[10:0]; // @[Modules.scala 50:57:@6049.4]
  assign buffer_1_415 = $signed(_T_59521); // @[Modules.scala 50:57:@6050.4]
  assign buffer_1_48 = {{6{_T_57733[4]}},_T_57733}; // @[Modules.scala 32:22:@8.4]
  assign _T_59523 = $signed(buffer_1_48) + $signed(buffer_0_49); // @[Modules.scala 50:57:@6052.4]
  assign _T_59524 = _T_59523[10:0]; // @[Modules.scala 50:57:@6053.4]
  assign buffer_1_416 = $signed(_T_59524); // @[Modules.scala 50:57:@6054.4]
  assign buffer_1_54 = {{6{_T_57751[4]}},_T_57751}; // @[Modules.scala 32:22:@8.4]
  assign _T_59532 = $signed(buffer_1_54) + $signed(buffer_0_55); // @[Modules.scala 50:57:@6064.4]
  assign _T_59533 = _T_59532[10:0]; // @[Modules.scala 50:57:@6065.4]
  assign buffer_1_419 = $signed(_T_59533); // @[Modules.scala 50:57:@6066.4]
  assign buffer_1_56 = {{6{_T_57761[4]}},_T_57761}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_57 = {{6{_T_57768[4]}},_T_57768}; // @[Modules.scala 32:22:@8.4]
  assign _T_59535 = $signed(buffer_1_56) + $signed(buffer_1_57); // @[Modules.scala 50:57:@6068.4]
  assign _T_59536 = _T_59535[10:0]; // @[Modules.scala 50:57:@6069.4]
  assign buffer_1_420 = $signed(_T_59536); // @[Modules.scala 50:57:@6070.4]
  assign buffer_1_59 = {{6{_T_57778[4]}},_T_57778}; // @[Modules.scala 32:22:@8.4]
  assign _T_59538 = $signed(buffer_0_58) + $signed(buffer_1_59); // @[Modules.scala 50:57:@6072.4]
  assign _T_59539 = _T_59538[10:0]; // @[Modules.scala 50:57:@6073.4]
  assign buffer_1_421 = $signed(_T_59539); // @[Modules.scala 50:57:@6074.4]
  assign buffer_1_63 = {{6{_T_57806[4]}},_T_57806}; // @[Modules.scala 32:22:@8.4]
  assign _T_59544 = $signed(buffer_0_62) + $signed(buffer_1_63); // @[Modules.scala 50:57:@6080.4]
  assign _T_59545 = _T_59544[10:0]; // @[Modules.scala 50:57:@6081.4]
  assign buffer_1_423 = $signed(_T_59545); // @[Modules.scala 50:57:@6082.4]
  assign buffer_1_64 = {{6{_T_57809[4]}},_T_57809}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_65 = {{6{_T_57812[4]}},_T_57812}; // @[Modules.scala 32:22:@8.4]
  assign _T_59547 = $signed(buffer_1_64) + $signed(buffer_1_65); // @[Modules.scala 50:57:@6084.4]
  assign _T_59548 = _T_59547[10:0]; // @[Modules.scala 50:57:@6085.4]
  assign buffer_1_424 = $signed(_T_59548); // @[Modules.scala 50:57:@6086.4]
  assign buffer_1_66 = {{6{_T_57819[4]}},_T_57819}; // @[Modules.scala 32:22:@8.4]
  assign _T_59550 = $signed(buffer_1_66) + $signed(buffer_0_67); // @[Modules.scala 50:57:@6088.4]
  assign _T_59551 = _T_59550[10:0]; // @[Modules.scala 50:57:@6089.4]
  assign buffer_1_425 = $signed(_T_59551); // @[Modules.scala 50:57:@6090.4]
  assign buffer_1_68 = {{6{_T_57825[4]}},_T_57825}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_69 = {{6{_T_57832[4]}},_T_57832}; // @[Modules.scala 32:22:@8.4]
  assign _T_59553 = $signed(buffer_1_68) + $signed(buffer_1_69); // @[Modules.scala 50:57:@6092.4]
  assign _T_59554 = _T_59553[10:0]; // @[Modules.scala 50:57:@6093.4]
  assign buffer_1_426 = $signed(_T_59554); // @[Modules.scala 50:57:@6094.4]
  assign buffer_1_70 = {{6{_T_57835[4]}},_T_57835}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_71 = {{6{_T_57842[4]}},_T_57842}; // @[Modules.scala 32:22:@8.4]
  assign _T_59556 = $signed(buffer_1_70) + $signed(buffer_1_71); // @[Modules.scala 50:57:@6096.4]
  assign _T_59557 = _T_59556[10:0]; // @[Modules.scala 50:57:@6097.4]
  assign buffer_1_427 = $signed(_T_59557); // @[Modules.scala 50:57:@6098.4]
  assign buffer_1_72 = {{6{_T_57849[4]}},_T_57849}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_73 = {{6{_T_57856[4]}},_T_57856}; // @[Modules.scala 32:22:@8.4]
  assign _T_59559 = $signed(buffer_1_72) + $signed(buffer_1_73); // @[Modules.scala 50:57:@6100.4]
  assign _T_59560 = _T_59559[10:0]; // @[Modules.scala 50:57:@6101.4]
  assign buffer_1_428 = $signed(_T_59560); // @[Modules.scala 50:57:@6102.4]
  assign buffer_1_74 = {{6{_T_57859[4]}},_T_57859}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_75 = {{6{_T_57862[4]}},_T_57862}; // @[Modules.scala 32:22:@8.4]
  assign _T_59562 = $signed(buffer_1_74) + $signed(buffer_1_75); // @[Modules.scala 50:57:@6104.4]
  assign _T_59563 = _T_59562[10:0]; // @[Modules.scala 50:57:@6105.4]
  assign buffer_1_429 = $signed(_T_59563); // @[Modules.scala 50:57:@6106.4]
  assign buffer_1_78 = {{6{_T_57879[4]}},_T_57879}; // @[Modules.scala 32:22:@8.4]
  assign _T_59568 = $signed(buffer_1_78) + $signed(buffer_0_79); // @[Modules.scala 50:57:@6112.4]
  assign _T_59569 = _T_59568[10:0]; // @[Modules.scala 50:57:@6113.4]
  assign buffer_1_431 = $signed(_T_59569); // @[Modules.scala 50:57:@6114.4]
  assign buffer_1_81 = {{6{_T_57900[4]}},_T_57900}; // @[Modules.scala 32:22:@8.4]
  assign _T_59571 = $signed(buffer_0_80) + $signed(buffer_1_81); // @[Modules.scala 50:57:@6116.4]
  assign _T_59572 = _T_59571[10:0]; // @[Modules.scala 50:57:@6117.4]
  assign buffer_1_432 = $signed(_T_59572); // @[Modules.scala 50:57:@6118.4]
  assign buffer_1_82 = {{6{_T_57907[4]}},_T_57907}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_83 = {{6{_T_57910[4]}},_T_57910}; // @[Modules.scala 32:22:@8.4]
  assign _T_59574 = $signed(buffer_1_82) + $signed(buffer_1_83); // @[Modules.scala 50:57:@6120.4]
  assign _T_59575 = _T_59574[10:0]; // @[Modules.scala 50:57:@6121.4]
  assign buffer_1_433 = $signed(_T_59575); // @[Modules.scala 50:57:@6122.4]
  assign buffer_1_84 = {{6{_T_57917[4]}},_T_57917}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_85 = {{6{_T_57920[4]}},_T_57920}; // @[Modules.scala 32:22:@8.4]
  assign _T_59577 = $signed(buffer_1_84) + $signed(buffer_1_85); // @[Modules.scala 50:57:@6124.4]
  assign _T_59578 = _T_59577[10:0]; // @[Modules.scala 50:57:@6125.4]
  assign buffer_1_434 = $signed(_T_59578); // @[Modules.scala 50:57:@6126.4]
  assign buffer_1_87 = {{6{_T_57926[4]}},_T_57926}; // @[Modules.scala 32:22:@8.4]
  assign _T_59580 = $signed(buffer_0_86) + $signed(buffer_1_87); // @[Modules.scala 50:57:@6128.4]
  assign _T_59581 = _T_59580[10:0]; // @[Modules.scala 50:57:@6129.4]
  assign buffer_1_435 = $signed(_T_59581); // @[Modules.scala 50:57:@6130.4]
  assign buffer_1_88 = {{6{_T_57929[4]}},_T_57929}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_89 = {{6{_T_57932[4]}},_T_57932}; // @[Modules.scala 32:22:@8.4]
  assign _T_59583 = $signed(buffer_1_88) + $signed(buffer_1_89); // @[Modules.scala 50:57:@6132.4]
  assign _T_59584 = _T_59583[10:0]; // @[Modules.scala 50:57:@6133.4]
  assign buffer_1_436 = $signed(_T_59584); // @[Modules.scala 50:57:@6134.4]
  assign buffer_1_91 = {{6{_T_57942[4]}},_T_57942}; // @[Modules.scala 32:22:@8.4]
  assign _T_59586 = $signed(buffer_0_90) + $signed(buffer_1_91); // @[Modules.scala 50:57:@6136.4]
  assign _T_59587 = _T_59586[10:0]; // @[Modules.scala 50:57:@6137.4]
  assign buffer_1_437 = $signed(_T_59587); // @[Modules.scala 50:57:@6138.4]
  assign buffer_1_94 = {{6{_T_57955[4]}},_T_57955}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_95 = {{6{_T_57962[4]}},_T_57962}; // @[Modules.scala 32:22:@8.4]
  assign _T_59592 = $signed(buffer_1_94) + $signed(buffer_1_95); // @[Modules.scala 50:57:@6144.4]
  assign _T_59593 = _T_59592[10:0]; // @[Modules.scala 50:57:@6145.4]
  assign buffer_1_439 = $signed(_T_59593); // @[Modules.scala 50:57:@6146.4]
  assign buffer_1_96 = {{6{_T_57969[4]}},_T_57969}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_97 = {{6{_T_57976[4]}},_T_57976}; // @[Modules.scala 32:22:@8.4]
  assign _T_59595 = $signed(buffer_1_96) + $signed(buffer_1_97); // @[Modules.scala 50:57:@6148.4]
  assign _T_59596 = _T_59595[10:0]; // @[Modules.scala 50:57:@6149.4]
  assign buffer_1_440 = $signed(_T_59596); // @[Modules.scala 50:57:@6150.4]
  assign buffer_1_98 = {{6{_T_57979[4]}},_T_57979}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_99 = {{6{_T_57986[4]}},_T_57986}; // @[Modules.scala 32:22:@8.4]
  assign _T_59598 = $signed(buffer_1_98) + $signed(buffer_1_99); // @[Modules.scala 50:57:@6152.4]
  assign _T_59599 = _T_59598[10:0]; // @[Modules.scala 50:57:@6153.4]
  assign buffer_1_441 = $signed(_T_59599); // @[Modules.scala 50:57:@6154.4]
  assign buffer_1_100 = {{6{_T_57993[4]}},_T_57993}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_101 = {{6{_T_57996[4]}},_T_57996}; // @[Modules.scala 32:22:@8.4]
  assign _T_59601 = $signed(buffer_1_100) + $signed(buffer_1_101); // @[Modules.scala 50:57:@6156.4]
  assign _T_59602 = _T_59601[10:0]; // @[Modules.scala 50:57:@6157.4]
  assign buffer_1_442 = $signed(_T_59602); // @[Modules.scala 50:57:@6158.4]
  assign buffer_1_102 = {{6{_T_58003[4]}},_T_58003}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_103 = {{6{_T_58006[4]}},_T_58006}; // @[Modules.scala 32:22:@8.4]
  assign _T_59604 = $signed(buffer_1_102) + $signed(buffer_1_103); // @[Modules.scala 50:57:@6160.4]
  assign _T_59605 = _T_59604[10:0]; // @[Modules.scala 50:57:@6161.4]
  assign buffer_1_443 = $signed(_T_59605); // @[Modules.scala 50:57:@6162.4]
  assign buffer_1_104 = {{6{_T_58009[4]}},_T_58009}; // @[Modules.scala 32:22:@8.4]
  assign _T_59607 = $signed(buffer_1_104) + $signed(buffer_0_105); // @[Modules.scala 50:57:@6164.4]
  assign _T_59608 = _T_59607[10:0]; // @[Modules.scala 50:57:@6165.4]
  assign buffer_1_444 = $signed(_T_59608); // @[Modules.scala 50:57:@6166.4]
  assign buffer_1_106 = {{6{_T_58019[4]}},_T_58019}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_107 = {{6{_T_58026[4]}},_T_58026}; // @[Modules.scala 32:22:@8.4]
  assign _T_59610 = $signed(buffer_1_106) + $signed(buffer_1_107); // @[Modules.scala 50:57:@6168.4]
  assign _T_59611 = _T_59610[10:0]; // @[Modules.scala 50:57:@6169.4]
  assign buffer_1_445 = $signed(_T_59611); // @[Modules.scala 50:57:@6170.4]
  assign buffer_1_108 = {{6{_T_58033[4]}},_T_58033}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_109 = {{6{_T_58040[4]}},_T_58040}; // @[Modules.scala 32:22:@8.4]
  assign _T_59613 = $signed(buffer_1_108) + $signed(buffer_1_109); // @[Modules.scala 50:57:@6172.4]
  assign _T_59614 = _T_59613[10:0]; // @[Modules.scala 50:57:@6173.4]
  assign buffer_1_446 = $signed(_T_59614); // @[Modules.scala 50:57:@6174.4]
  assign buffer_1_110 = {{6{_T_58043[4]}},_T_58043}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_111 = {{6{_T_58050[4]}},_T_58050}; // @[Modules.scala 32:22:@8.4]
  assign _T_59616 = $signed(buffer_1_110) + $signed(buffer_1_111); // @[Modules.scala 50:57:@6176.4]
  assign _T_59617 = _T_59616[10:0]; // @[Modules.scala 50:57:@6177.4]
  assign buffer_1_447 = $signed(_T_59617); // @[Modules.scala 50:57:@6178.4]
  assign buffer_1_112 = {{6{_T_58053[4]}},_T_58053}; // @[Modules.scala 32:22:@8.4]
  assign _T_59619 = $signed(buffer_1_112) + $signed(buffer_0_113); // @[Modules.scala 50:57:@6180.4]
  assign _T_59620 = _T_59619[10:0]; // @[Modules.scala 50:57:@6181.4]
  assign buffer_1_448 = $signed(_T_59620); // @[Modules.scala 50:57:@6182.4]
  assign buffer_1_118 = {{6{_T_58095[4]}},_T_58095}; // @[Modules.scala 32:22:@8.4]
  assign _T_59628 = $signed(buffer_1_118) + $signed(buffer_0_119); // @[Modules.scala 50:57:@6192.4]
  assign _T_59629 = _T_59628[10:0]; // @[Modules.scala 50:57:@6193.4]
  assign buffer_1_451 = $signed(_T_59629); // @[Modules.scala 50:57:@6194.4]
  assign buffer_1_120 = {{6{_T_58105[4]}},_T_58105}; // @[Modules.scala 32:22:@8.4]
  assign _T_59631 = $signed(buffer_1_120) + $signed(buffer_0_121); // @[Modules.scala 50:57:@6196.4]
  assign _T_59632 = _T_59631[10:0]; // @[Modules.scala 50:57:@6197.4]
  assign buffer_1_452 = $signed(_T_59632); // @[Modules.scala 50:57:@6198.4]
  assign buffer_1_123 = {{6{_T_58126[4]}},_T_58126}; // @[Modules.scala 32:22:@8.4]
  assign _T_59634 = $signed(buffer_0_122) + $signed(buffer_1_123); // @[Modules.scala 50:57:@6200.4]
  assign _T_59635 = _T_59634[10:0]; // @[Modules.scala 50:57:@6201.4]
  assign buffer_1_453 = $signed(_T_59635); // @[Modules.scala 50:57:@6202.4]
  assign buffer_1_124 = {{6{_T_58129[4]}},_T_58129}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_125 = {{6{_T_58132[4]}},_T_58132}; // @[Modules.scala 32:22:@8.4]
  assign _T_59637 = $signed(buffer_1_124) + $signed(buffer_1_125); // @[Modules.scala 50:57:@6204.4]
  assign _T_59638 = _T_59637[10:0]; // @[Modules.scala 50:57:@6205.4]
  assign buffer_1_454 = $signed(_T_59638); // @[Modules.scala 50:57:@6206.4]
  assign buffer_1_126 = {{6{_T_58139[4]}},_T_58139}; // @[Modules.scala 32:22:@8.4]
  assign _T_59640 = $signed(buffer_1_126) + $signed(buffer_0_127); // @[Modules.scala 50:57:@6208.4]
  assign _T_59641 = _T_59640[10:0]; // @[Modules.scala 50:57:@6209.4]
  assign buffer_1_455 = $signed(_T_59641); // @[Modules.scala 50:57:@6210.4]
  assign buffer_1_130 = {{6{_T_58163[4]}},_T_58163}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_131 = {{6{_T_58170[4]}},_T_58170}; // @[Modules.scala 32:22:@8.4]
  assign _T_59646 = $signed(buffer_1_130) + $signed(buffer_1_131); // @[Modules.scala 50:57:@6216.4]
  assign _T_59647 = _T_59646[10:0]; // @[Modules.scala 50:57:@6217.4]
  assign buffer_1_457 = $signed(_T_59647); // @[Modules.scala 50:57:@6218.4]
  assign buffer_1_133 = {{6{_T_58180[4]}},_T_58180}; // @[Modules.scala 32:22:@8.4]
  assign _T_59649 = $signed(buffer_0_132) + $signed(buffer_1_133); // @[Modules.scala 50:57:@6220.4]
  assign _T_59650 = _T_59649[10:0]; // @[Modules.scala 50:57:@6221.4]
  assign buffer_1_458 = $signed(_T_59650); // @[Modules.scala 50:57:@6222.4]
  assign buffer_1_137 = {{6{_T_58208[4]}},_T_58208}; // @[Modules.scala 32:22:@8.4]
  assign _T_59655 = $signed(buffer_0_136) + $signed(buffer_1_137); // @[Modules.scala 50:57:@6228.4]
  assign _T_59656 = _T_59655[10:0]; // @[Modules.scala 50:57:@6229.4]
  assign buffer_1_460 = $signed(_T_59656); // @[Modules.scala 50:57:@6230.4]
  assign buffer_1_138 = {{6{_T_58211[4]}},_T_58211}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_139 = {{6{_T_58214[4]}},_T_58214}; // @[Modules.scala 32:22:@8.4]
  assign _T_59658 = $signed(buffer_1_138) + $signed(buffer_1_139); // @[Modules.scala 50:57:@6232.4]
  assign _T_59659 = _T_59658[10:0]; // @[Modules.scala 50:57:@6233.4]
  assign buffer_1_461 = $signed(_T_59659); // @[Modules.scala 50:57:@6234.4]
  assign buffer_1_140 = {{6{_T_58221[4]}},_T_58221}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_141 = {{6{_T_58228[4]}},_T_58228}; // @[Modules.scala 32:22:@8.4]
  assign _T_59661 = $signed(buffer_1_140) + $signed(buffer_1_141); // @[Modules.scala 50:57:@6236.4]
  assign _T_59662 = _T_59661[10:0]; // @[Modules.scala 50:57:@6237.4]
  assign buffer_1_462 = $signed(_T_59662); // @[Modules.scala 50:57:@6238.4]
  assign buffer_1_146 = {{6{_T_58259[4]}},_T_58259}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_147 = {{6{_T_58262[4]}},_T_58262}; // @[Modules.scala 32:22:@8.4]
  assign _T_59670 = $signed(buffer_1_146) + $signed(buffer_1_147); // @[Modules.scala 50:57:@6248.4]
  assign _T_59671 = _T_59670[10:0]; // @[Modules.scala 50:57:@6249.4]
  assign buffer_1_465 = $signed(_T_59671); // @[Modules.scala 50:57:@6250.4]
  assign buffer_1_151 = {{6{_T_58290[4]}},_T_58290}; // @[Modules.scala 32:22:@8.4]
  assign _T_59676 = $signed(buffer_0_150) + $signed(buffer_1_151); // @[Modules.scala 50:57:@6256.4]
  assign _T_59677 = _T_59676[10:0]; // @[Modules.scala 50:57:@6257.4]
  assign buffer_1_467 = $signed(_T_59677); // @[Modules.scala 50:57:@6258.4]
  assign buffer_1_152 = {{6{_T_58293[4]}},_T_58293}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_153 = {{6{_T_58296[4]}},_T_58296}; // @[Modules.scala 32:22:@8.4]
  assign _T_59679 = $signed(buffer_1_152) + $signed(buffer_1_153); // @[Modules.scala 50:57:@6260.4]
  assign _T_59680 = _T_59679[10:0]; // @[Modules.scala 50:57:@6261.4]
  assign buffer_1_468 = $signed(_T_59680); // @[Modules.scala 50:57:@6262.4]
  assign buffer_1_157 = {{6{_T_58320[4]}},_T_58320}; // @[Modules.scala 32:22:@8.4]
  assign _T_59685 = $signed(buffer_0_156) + $signed(buffer_1_157); // @[Modules.scala 50:57:@6268.4]
  assign _T_59686 = _T_59685[10:0]; // @[Modules.scala 50:57:@6269.4]
  assign buffer_1_470 = $signed(_T_59686); // @[Modules.scala 50:57:@6270.4]
  assign buffer_1_158 = {{6{_T_58327[4]}},_T_58327}; // @[Modules.scala 32:22:@8.4]
  assign _T_59688 = $signed(buffer_1_158) + $signed(buffer_0_159); // @[Modules.scala 50:57:@6272.4]
  assign _T_59689 = _T_59688[10:0]; // @[Modules.scala 50:57:@6273.4]
  assign buffer_1_471 = $signed(_T_59689); // @[Modules.scala 50:57:@6274.4]
  assign buffer_1_160 = {{6{_T_58333[4]}},_T_58333}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_161 = {{6{_T_58336[4]}},_T_58336}; // @[Modules.scala 32:22:@8.4]
  assign _T_59691 = $signed(buffer_1_160) + $signed(buffer_1_161); // @[Modules.scala 50:57:@6276.4]
  assign _T_59692 = _T_59691[10:0]; // @[Modules.scala 50:57:@6277.4]
  assign buffer_1_472 = $signed(_T_59692); // @[Modules.scala 50:57:@6278.4]
  assign buffer_1_162 = {{6{_T_58343[4]}},_T_58343}; // @[Modules.scala 32:22:@8.4]
  assign _T_59694 = $signed(buffer_1_162) + $signed(buffer_0_163); // @[Modules.scala 50:57:@6280.4]
  assign _T_59695 = _T_59694[10:0]; // @[Modules.scala 50:57:@6281.4]
  assign buffer_1_473 = $signed(_T_59695); // @[Modules.scala 50:57:@6282.4]
  assign buffer_1_164 = {{6{_T_58357[4]}},_T_58357}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_165 = {{6{_T_58364[4]}},_T_58364}; // @[Modules.scala 32:22:@8.4]
  assign _T_59697 = $signed(buffer_1_164) + $signed(buffer_1_165); // @[Modules.scala 50:57:@6284.4]
  assign _T_59698 = _T_59697[10:0]; // @[Modules.scala 50:57:@6285.4]
  assign buffer_1_474 = $signed(_T_59698); // @[Modules.scala 50:57:@6286.4]
  assign buffer_1_166 = {{6{_T_58367[4]}},_T_58367}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_167 = {{6{_T_58370[4]}},_T_58370}; // @[Modules.scala 32:22:@8.4]
  assign _T_59700 = $signed(buffer_1_166) + $signed(buffer_1_167); // @[Modules.scala 50:57:@6288.4]
  assign _T_59701 = _T_59700[10:0]; // @[Modules.scala 50:57:@6289.4]
  assign buffer_1_475 = $signed(_T_59701); // @[Modules.scala 50:57:@6290.4]
  assign buffer_1_175 = {{6{_T_58406[4]}},_T_58406}; // @[Modules.scala 32:22:@8.4]
  assign _T_59712 = $signed(buffer_0_174) + $signed(buffer_1_175); // @[Modules.scala 50:57:@6304.4]
  assign _T_59713 = _T_59712[10:0]; // @[Modules.scala 50:57:@6305.4]
  assign buffer_1_479 = $signed(_T_59713); // @[Modules.scala 50:57:@6306.4]
  assign buffer_1_176 = {{6{_T_58413[4]}},_T_58413}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_177 = {{6{_T_58420[4]}},_T_58420}; // @[Modules.scala 32:22:@8.4]
  assign _T_59715 = $signed(buffer_1_176) + $signed(buffer_1_177); // @[Modules.scala 50:57:@6308.4]
  assign _T_59716 = _T_59715[10:0]; // @[Modules.scala 50:57:@6309.4]
  assign buffer_1_480 = $signed(_T_59716); // @[Modules.scala 50:57:@6310.4]
  assign buffer_1_178 = {{6{_T_58427[4]}},_T_58427}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_179 = {{6{_T_58434[4]}},_T_58434}; // @[Modules.scala 32:22:@8.4]
  assign _T_59718 = $signed(buffer_1_178) + $signed(buffer_1_179); // @[Modules.scala 50:57:@6312.4]
  assign _T_59719 = _T_59718[10:0]; // @[Modules.scala 50:57:@6313.4]
  assign buffer_1_481 = $signed(_T_59719); // @[Modules.scala 50:57:@6314.4]
  assign buffer_1_180 = {{6{_T_58437[4]}},_T_58437}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_181 = {{6{_T_58444[4]}},_T_58444}; // @[Modules.scala 32:22:@8.4]
  assign _T_59721 = $signed(buffer_1_180) + $signed(buffer_1_181); // @[Modules.scala 50:57:@6316.4]
  assign _T_59722 = _T_59721[10:0]; // @[Modules.scala 50:57:@6317.4]
  assign buffer_1_482 = $signed(_T_59722); // @[Modules.scala 50:57:@6318.4]
  assign buffer_1_184 = {{6{_T_58465[4]}},_T_58465}; // @[Modules.scala 32:22:@8.4]
  assign _T_59727 = $signed(buffer_1_184) + $signed(buffer_0_185); // @[Modules.scala 50:57:@6324.4]
  assign _T_59728 = _T_59727[10:0]; // @[Modules.scala 50:57:@6325.4]
  assign buffer_1_484 = $signed(_T_59728); // @[Modules.scala 50:57:@6326.4]
  assign buffer_1_189 = {{6{_T_58484[4]}},_T_58484}; // @[Modules.scala 32:22:@8.4]
  assign _T_59733 = $signed(buffer_0_188) + $signed(buffer_1_189); // @[Modules.scala 50:57:@6332.4]
  assign _T_59734 = _T_59733[10:0]; // @[Modules.scala 50:57:@6333.4]
  assign buffer_1_486 = $signed(_T_59734); // @[Modules.scala 50:57:@6334.4]
  assign buffer_1_190 = {{6{_T_58491[4]}},_T_58491}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_191 = {{6{_T_58498[4]}},_T_58498}; // @[Modules.scala 32:22:@8.4]
  assign _T_59736 = $signed(buffer_1_190) + $signed(buffer_1_191); // @[Modules.scala 50:57:@6336.4]
  assign _T_59737 = _T_59736[10:0]; // @[Modules.scala 50:57:@6337.4]
  assign buffer_1_487 = $signed(_T_59737); // @[Modules.scala 50:57:@6338.4]
  assign buffer_1_195 = {{6{_T_58518[4]}},_T_58518}; // @[Modules.scala 32:22:@8.4]
  assign _T_59742 = $signed(buffer_0_194) + $signed(buffer_1_195); // @[Modules.scala 50:57:@6344.4]
  assign _T_59743 = _T_59742[10:0]; // @[Modules.scala 50:57:@6345.4]
  assign buffer_1_489 = $signed(_T_59743); // @[Modules.scala 50:57:@6346.4]
  assign buffer_1_196 = {{6{_T_58521[4]}},_T_58521}; // @[Modules.scala 32:22:@8.4]
  assign _T_59745 = $signed(buffer_1_196) + $signed(buffer_0_197); // @[Modules.scala 50:57:@6348.4]
  assign _T_59746 = _T_59745[10:0]; // @[Modules.scala 50:57:@6349.4]
  assign buffer_1_490 = $signed(_T_59746); // @[Modules.scala 50:57:@6350.4]
  assign buffer_1_198 = {{6{_T_58535[4]}},_T_58535}; // @[Modules.scala 32:22:@8.4]
  assign _T_59748 = $signed(buffer_1_198) + $signed(buffer_0_199); // @[Modules.scala 50:57:@6352.4]
  assign _T_59749 = _T_59748[10:0]; // @[Modules.scala 50:57:@6353.4]
  assign buffer_1_491 = $signed(_T_59749); // @[Modules.scala 50:57:@6354.4]
  assign buffer_1_202 = {{6{_T_58547[4]}},_T_58547}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_203 = {{6{_T_58554[4]}},_T_58554}; // @[Modules.scala 32:22:@8.4]
  assign _T_59754 = $signed(buffer_1_202) + $signed(buffer_1_203); // @[Modules.scala 50:57:@6360.4]
  assign _T_59755 = _T_59754[10:0]; // @[Modules.scala 50:57:@6361.4]
  assign buffer_1_493 = $signed(_T_59755); // @[Modules.scala 50:57:@6362.4]
  assign buffer_1_204 = {{6{_T_58557[4]}},_T_58557}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_205 = {{6{_T_58564[4]}},_T_58564}; // @[Modules.scala 32:22:@8.4]
  assign _T_59757 = $signed(buffer_1_204) + $signed(buffer_1_205); // @[Modules.scala 50:57:@6364.4]
  assign _T_59758 = _T_59757[10:0]; // @[Modules.scala 50:57:@6365.4]
  assign buffer_1_494 = $signed(_T_59758); // @[Modules.scala 50:57:@6366.4]
  assign buffer_1_209 = {{6{_T_58580[4]}},_T_58580}; // @[Modules.scala 32:22:@8.4]
  assign _T_59763 = $signed(buffer_0_208) + $signed(buffer_1_209); // @[Modules.scala 50:57:@6372.4]
  assign _T_59764 = _T_59763[10:0]; // @[Modules.scala 50:57:@6373.4]
  assign buffer_1_496 = $signed(_T_59764); // @[Modules.scala 50:57:@6374.4]
  assign buffer_1_211 = {{6{_T_58590[4]}},_T_58590}; // @[Modules.scala 32:22:@8.4]
  assign _T_59766 = $signed(buffer_0_210) + $signed(buffer_1_211); // @[Modules.scala 50:57:@6376.4]
  assign _T_59767 = _T_59766[10:0]; // @[Modules.scala 50:57:@6377.4]
  assign buffer_1_497 = $signed(_T_59767); // @[Modules.scala 50:57:@6378.4]
  assign buffer_1_213 = {{6{_T_58604[4]}},_T_58604}; // @[Modules.scala 32:22:@8.4]
  assign _T_59769 = $signed(buffer_0_212) + $signed(buffer_1_213); // @[Modules.scala 50:57:@6380.4]
  assign _T_59770 = _T_59769[10:0]; // @[Modules.scala 50:57:@6381.4]
  assign buffer_1_498 = $signed(_T_59770); // @[Modules.scala 50:57:@6382.4]
  assign buffer_1_216 = {{6{_T_58617[4]}},_T_58617}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_217 = {{6{_T_58624[4]}},_T_58624}; // @[Modules.scala 32:22:@8.4]
  assign _T_59775 = $signed(buffer_1_216) + $signed(buffer_1_217); // @[Modules.scala 50:57:@6388.4]
  assign _T_59776 = _T_59775[10:0]; // @[Modules.scala 50:57:@6389.4]
  assign buffer_1_500 = $signed(_T_59776); // @[Modules.scala 50:57:@6390.4]
  assign buffer_1_218 = {{6{_T_58631[4]}},_T_58631}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_219 = {{6{_T_58638[4]}},_T_58638}; // @[Modules.scala 32:22:@8.4]
  assign _T_59778 = $signed(buffer_1_218) + $signed(buffer_1_219); // @[Modules.scala 50:57:@6392.4]
  assign _T_59779 = _T_59778[10:0]; // @[Modules.scala 50:57:@6393.4]
  assign buffer_1_501 = $signed(_T_59779); // @[Modules.scala 50:57:@6394.4]
  assign buffer_1_220 = {{6{_T_58641[4]}},_T_58641}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_221 = {{6{_T_58644[4]}},_T_58644}; // @[Modules.scala 32:22:@8.4]
  assign _T_59781 = $signed(buffer_1_220) + $signed(buffer_1_221); // @[Modules.scala 50:57:@6396.4]
  assign _T_59782 = _T_59781[10:0]; // @[Modules.scala 50:57:@6397.4]
  assign buffer_1_502 = $signed(_T_59782); // @[Modules.scala 50:57:@6398.4]
  assign buffer_1_222 = {{6{_T_58647[4]}},_T_58647}; // @[Modules.scala 32:22:@8.4]
  assign _T_59784 = $signed(buffer_1_222) + $signed(buffer_0_223); // @[Modules.scala 50:57:@6400.4]
  assign _T_59785 = _T_59784[10:0]; // @[Modules.scala 50:57:@6401.4]
  assign buffer_1_503 = $signed(_T_59785); // @[Modules.scala 50:57:@6402.4]
  assign buffer_1_224 = {{6{_T_58661[4]}},_T_58661}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_225 = {{6{_T_58664[4]}},_T_58664}; // @[Modules.scala 32:22:@8.4]
  assign _T_59787 = $signed(buffer_1_224) + $signed(buffer_1_225); // @[Modules.scala 50:57:@6404.4]
  assign _T_59788 = _T_59787[10:0]; // @[Modules.scala 50:57:@6405.4]
  assign buffer_1_504 = $signed(_T_59788); // @[Modules.scala 50:57:@6406.4]
  assign buffer_1_226 = {{6{_T_58671[4]}},_T_58671}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_227 = {{6{_T_58678[4]}},_T_58678}; // @[Modules.scala 32:22:@8.4]
  assign _T_59790 = $signed(buffer_1_226) + $signed(buffer_1_227); // @[Modules.scala 50:57:@6408.4]
  assign _T_59791 = _T_59790[10:0]; // @[Modules.scala 50:57:@6409.4]
  assign buffer_1_505 = $signed(_T_59791); // @[Modules.scala 50:57:@6410.4]
  assign buffer_1_228 = {{6{_T_58685[4]}},_T_58685}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_229 = {{6{_T_58688[4]}},_T_58688}; // @[Modules.scala 32:22:@8.4]
  assign _T_59793 = $signed(buffer_1_228) + $signed(buffer_1_229); // @[Modules.scala 50:57:@6412.4]
  assign _T_59794 = _T_59793[10:0]; // @[Modules.scala 50:57:@6413.4]
  assign buffer_1_506 = $signed(_T_59794); // @[Modules.scala 50:57:@6414.4]
  assign buffer_1_230 = {{6{_T_58695[4]}},_T_58695}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_231 = {{6{_T_58702[4]}},_T_58702}; // @[Modules.scala 32:22:@8.4]
  assign _T_59796 = $signed(buffer_1_230) + $signed(buffer_1_231); // @[Modules.scala 50:57:@6416.4]
  assign _T_59797 = _T_59796[10:0]; // @[Modules.scala 50:57:@6417.4]
  assign buffer_1_507 = $signed(_T_59797); // @[Modules.scala 50:57:@6418.4]
  assign buffer_1_232 = {{6{_T_58709[4]}},_T_58709}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_233 = {{6{_T_58716[4]}},_T_58716}; // @[Modules.scala 32:22:@8.4]
  assign _T_59799 = $signed(buffer_1_232) + $signed(buffer_1_233); // @[Modules.scala 50:57:@6420.4]
  assign _T_59800 = _T_59799[10:0]; // @[Modules.scala 50:57:@6421.4]
  assign buffer_1_508 = $signed(_T_59800); // @[Modules.scala 50:57:@6422.4]
  assign buffer_1_234 = {{6{_T_58719[4]}},_T_58719}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_235 = {{6{_T_58722[4]}},_T_58722}; // @[Modules.scala 32:22:@8.4]
  assign _T_59802 = $signed(buffer_1_234) + $signed(buffer_1_235); // @[Modules.scala 50:57:@6424.4]
  assign _T_59803 = _T_59802[10:0]; // @[Modules.scala 50:57:@6425.4]
  assign buffer_1_509 = $signed(_T_59803); // @[Modules.scala 50:57:@6426.4]
  assign buffer_1_236 = {{6{_T_58725[4]}},_T_58725}; // @[Modules.scala 32:22:@8.4]
  assign _T_59805 = $signed(buffer_1_236) + $signed(buffer_0_237); // @[Modules.scala 50:57:@6428.4]
  assign _T_59806 = _T_59805[10:0]; // @[Modules.scala 50:57:@6429.4]
  assign buffer_1_510 = $signed(_T_59806); // @[Modules.scala 50:57:@6430.4]
  assign buffer_1_238 = {{6{_T_58739[4]}},_T_58739}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_239 = {{6{_T_58742[4]}},_T_58742}; // @[Modules.scala 32:22:@8.4]
  assign _T_59808 = $signed(buffer_1_238) + $signed(buffer_1_239); // @[Modules.scala 50:57:@6432.4]
  assign _T_59809 = _T_59808[10:0]; // @[Modules.scala 50:57:@6433.4]
  assign buffer_1_511 = $signed(_T_59809); // @[Modules.scala 50:57:@6434.4]
  assign buffer_1_242 = {{6{_T_58759[4]}},_T_58759}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_243 = {{6{_T_58766[4]}},_T_58766}; // @[Modules.scala 32:22:@8.4]
  assign _T_59814 = $signed(buffer_1_242) + $signed(buffer_1_243); // @[Modules.scala 50:57:@6440.4]
  assign _T_59815 = _T_59814[10:0]; // @[Modules.scala 50:57:@6441.4]
  assign buffer_1_513 = $signed(_T_59815); // @[Modules.scala 50:57:@6442.4]
  assign buffer_1_244 = {{6{_T_58773[4]}},_T_58773}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_245 = {{6{_T_58780[4]}},_T_58780}; // @[Modules.scala 32:22:@8.4]
  assign _T_59817 = $signed(buffer_1_244) + $signed(buffer_1_245); // @[Modules.scala 50:57:@6444.4]
  assign _T_59818 = _T_59817[10:0]; // @[Modules.scala 50:57:@6445.4]
  assign buffer_1_514 = $signed(_T_59818); // @[Modules.scala 50:57:@6446.4]
  assign buffer_1_246 = {{6{_T_58787[4]}},_T_58787}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_247 = {{6{_T_58790[4]}},_T_58790}; // @[Modules.scala 32:22:@8.4]
  assign _T_59820 = $signed(buffer_1_246) + $signed(buffer_1_247); // @[Modules.scala 50:57:@6448.4]
  assign _T_59821 = _T_59820[10:0]; // @[Modules.scala 50:57:@6449.4]
  assign buffer_1_515 = $signed(_T_59821); // @[Modules.scala 50:57:@6450.4]
  assign buffer_1_248 = {{6{_T_58793[4]}},_T_58793}; // @[Modules.scala 32:22:@8.4]
  assign _T_59823 = $signed(buffer_1_248) + $signed(buffer_0_249); // @[Modules.scala 50:57:@6452.4]
  assign _T_59824 = _T_59823[10:0]; // @[Modules.scala 50:57:@6453.4]
  assign buffer_1_516 = $signed(_T_59824); // @[Modules.scala 50:57:@6454.4]
  assign buffer_1_252 = {{6{_T_58817[4]}},_T_58817}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_253 = {{6{_T_58820[4]}},_T_58820}; // @[Modules.scala 32:22:@8.4]
  assign _T_59829 = $signed(buffer_1_252) + $signed(buffer_1_253); // @[Modules.scala 50:57:@6460.4]
  assign _T_59830 = _T_59829[10:0]; // @[Modules.scala 50:57:@6461.4]
  assign buffer_1_518 = $signed(_T_59830); // @[Modules.scala 50:57:@6462.4]
  assign buffer_1_254 = {{6{_T_58823[4]}},_T_58823}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_255 = {{6{_T_58826[4]}},_T_58826}; // @[Modules.scala 32:22:@8.4]
  assign _T_59832 = $signed(buffer_1_254) + $signed(buffer_1_255); // @[Modules.scala 50:57:@6464.4]
  assign _T_59833 = _T_59832[10:0]; // @[Modules.scala 50:57:@6465.4]
  assign buffer_1_519 = $signed(_T_59833); // @[Modules.scala 50:57:@6466.4]
  assign buffer_1_256 = {{6{_T_58833[4]}},_T_58833}; // @[Modules.scala 32:22:@8.4]
  assign _T_59835 = $signed(buffer_1_256) + $signed(buffer_0_257); // @[Modules.scala 50:57:@6468.4]
  assign _T_59836 = _T_59835[10:0]; // @[Modules.scala 50:57:@6469.4]
  assign buffer_1_520 = $signed(_T_59836); // @[Modules.scala 50:57:@6470.4]
  assign buffer_1_258 = {{6{_T_58843[4]}},_T_58843}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_259 = {{6{_T_58850[4]}},_T_58850}; // @[Modules.scala 32:22:@8.4]
  assign _T_59838 = $signed(buffer_1_258) + $signed(buffer_1_259); // @[Modules.scala 50:57:@6472.4]
  assign _T_59839 = _T_59838[10:0]; // @[Modules.scala 50:57:@6473.4]
  assign buffer_1_521 = $signed(_T_59839); // @[Modules.scala 50:57:@6474.4]
  assign buffer_1_260 = {{6{_T_58853[4]}},_T_58853}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_261 = {{6{_T_58856[4]}},_T_58856}; // @[Modules.scala 32:22:@8.4]
  assign _T_59841 = $signed(buffer_1_260) + $signed(buffer_1_261); // @[Modules.scala 50:57:@6476.4]
  assign _T_59842 = _T_59841[10:0]; // @[Modules.scala 50:57:@6477.4]
  assign buffer_1_522 = $signed(_T_59842); // @[Modules.scala 50:57:@6478.4]
  assign buffer_1_262 = {{6{_T_58859[4]}},_T_58859}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_263 = {{6{_T_58862[4]}},_T_58862}; // @[Modules.scala 32:22:@8.4]
  assign _T_59844 = $signed(buffer_1_262) + $signed(buffer_1_263); // @[Modules.scala 50:57:@6480.4]
  assign _T_59845 = _T_59844[10:0]; // @[Modules.scala 50:57:@6481.4]
  assign buffer_1_523 = $signed(_T_59845); // @[Modules.scala 50:57:@6482.4]
  assign buffer_1_264 = {{6{_T_58869[4]}},_T_58869}; // @[Modules.scala 32:22:@8.4]
  assign _T_59847 = $signed(buffer_1_264) + $signed(buffer_0_265); // @[Modules.scala 50:57:@6484.4]
  assign _T_59848 = _T_59847[10:0]; // @[Modules.scala 50:57:@6485.4]
  assign buffer_1_524 = $signed(_T_59848); // @[Modules.scala 50:57:@6486.4]
  assign buffer_1_266 = {{6{_T_58879[4]}},_T_58879}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_267 = {{6{_T_58882[4]}},_T_58882}; // @[Modules.scala 32:22:@8.4]
  assign _T_59850 = $signed(buffer_1_266) + $signed(buffer_1_267); // @[Modules.scala 50:57:@6488.4]
  assign _T_59851 = _T_59850[10:0]; // @[Modules.scala 50:57:@6489.4]
  assign buffer_1_525 = $signed(_T_59851); // @[Modules.scala 50:57:@6490.4]
  assign buffer_1_268 = {{6{_T_58885[4]}},_T_58885}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_269 = {{6{_T_58888[4]}},_T_58888}; // @[Modules.scala 32:22:@8.4]
  assign _T_59853 = $signed(buffer_1_268) + $signed(buffer_1_269); // @[Modules.scala 50:57:@6492.4]
  assign _T_59854 = _T_59853[10:0]; // @[Modules.scala 50:57:@6493.4]
  assign buffer_1_526 = $signed(_T_59854); // @[Modules.scala 50:57:@6494.4]
  assign buffer_1_270 = {{6{_T_58891[4]}},_T_58891}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_271 = {{6{_T_58894[4]}},_T_58894}; // @[Modules.scala 32:22:@8.4]
  assign _T_59856 = $signed(buffer_1_270) + $signed(buffer_1_271); // @[Modules.scala 50:57:@6496.4]
  assign _T_59857 = _T_59856[10:0]; // @[Modules.scala 50:57:@6497.4]
  assign buffer_1_527 = $signed(_T_59857); // @[Modules.scala 50:57:@6498.4]
  assign buffer_1_272 = {{6{_T_58897[4]}},_T_58897}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_273 = {{6{_T_58904[4]}},_T_58904}; // @[Modules.scala 32:22:@8.4]
  assign _T_59859 = $signed(buffer_1_272) + $signed(buffer_1_273); // @[Modules.scala 50:57:@6500.4]
  assign _T_59860 = _T_59859[10:0]; // @[Modules.scala 50:57:@6501.4]
  assign buffer_1_528 = $signed(_T_59860); // @[Modules.scala 50:57:@6502.4]
  assign buffer_1_274 = {{6{_T_58907[4]}},_T_58907}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_275 = {{6{_T_58910[4]}},_T_58910}; // @[Modules.scala 32:22:@8.4]
  assign _T_59862 = $signed(buffer_1_274) + $signed(buffer_1_275); // @[Modules.scala 50:57:@6504.4]
  assign _T_59863 = _T_59862[10:0]; // @[Modules.scala 50:57:@6505.4]
  assign buffer_1_529 = $signed(_T_59863); // @[Modules.scala 50:57:@6506.4]
  assign buffer_1_277 = {{6{_T_58916[4]}},_T_58916}; // @[Modules.scala 32:22:@8.4]
  assign _T_59865 = $signed(buffer_0_276) + $signed(buffer_1_277); // @[Modules.scala 50:57:@6508.4]
  assign _T_59866 = _T_59865[10:0]; // @[Modules.scala 50:57:@6509.4]
  assign buffer_1_530 = $signed(_T_59866); // @[Modules.scala 50:57:@6510.4]
  assign buffer_1_278 = {{6{_T_58923[4]}},_T_58923}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_279 = {{6{_T_58930[4]}},_T_58930}; // @[Modules.scala 32:22:@8.4]
  assign _T_59868 = $signed(buffer_1_278) + $signed(buffer_1_279); // @[Modules.scala 50:57:@6512.4]
  assign _T_59869 = _T_59868[10:0]; // @[Modules.scala 50:57:@6513.4]
  assign buffer_1_531 = $signed(_T_59869); // @[Modules.scala 50:57:@6514.4]
  assign buffer_1_280 = {{6{_T_58937[4]}},_T_58937}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_281 = {{6{_T_58940[4]}},_T_58940}; // @[Modules.scala 32:22:@8.4]
  assign _T_59871 = $signed(buffer_1_280) + $signed(buffer_1_281); // @[Modules.scala 50:57:@6516.4]
  assign _T_59872 = _T_59871[10:0]; // @[Modules.scala 50:57:@6517.4]
  assign buffer_1_532 = $signed(_T_59872); // @[Modules.scala 50:57:@6518.4]
  assign buffer_1_282 = {{6{_T_58943[4]}},_T_58943}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_283 = {{6{_T_58946[4]}},_T_58946}; // @[Modules.scala 32:22:@8.4]
  assign _T_59874 = $signed(buffer_1_282) + $signed(buffer_1_283); // @[Modules.scala 50:57:@6520.4]
  assign _T_59875 = _T_59874[10:0]; // @[Modules.scala 50:57:@6521.4]
  assign buffer_1_533 = $signed(_T_59875); // @[Modules.scala 50:57:@6522.4]
  assign buffer_1_284 = {{6{_T_58949[4]}},_T_58949}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_285 = {{6{_T_58952[4]}},_T_58952}; // @[Modules.scala 32:22:@8.4]
  assign _T_59877 = $signed(buffer_1_284) + $signed(buffer_1_285); // @[Modules.scala 50:57:@6524.4]
  assign _T_59878 = _T_59877[10:0]; // @[Modules.scala 50:57:@6525.4]
  assign buffer_1_534 = $signed(_T_59878); // @[Modules.scala 50:57:@6526.4]
  assign buffer_1_286 = {{6{_T_58955[4]}},_T_58955}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_287 = {{6{_T_58958[4]}},_T_58958}; // @[Modules.scala 32:22:@8.4]
  assign _T_59880 = $signed(buffer_1_286) + $signed(buffer_1_287); // @[Modules.scala 50:57:@6528.4]
  assign _T_59881 = _T_59880[10:0]; // @[Modules.scala 50:57:@6529.4]
  assign buffer_1_535 = $signed(_T_59881); // @[Modules.scala 50:57:@6530.4]
  assign buffer_1_288 = {{6{_T_58961[4]}},_T_58961}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_289 = {{6{_T_58964[4]}},_T_58964}; // @[Modules.scala 32:22:@8.4]
  assign _T_59883 = $signed(buffer_1_288) + $signed(buffer_1_289); // @[Modules.scala 50:57:@6532.4]
  assign _T_59884 = _T_59883[10:0]; // @[Modules.scala 50:57:@6533.4]
  assign buffer_1_536 = $signed(_T_59884); // @[Modules.scala 50:57:@6534.4]
  assign buffer_1_291 = {{6{_T_58970[4]}},_T_58970}; // @[Modules.scala 32:22:@8.4]
  assign _T_59886 = $signed(buffer_0_290) + $signed(buffer_1_291); // @[Modules.scala 50:57:@6536.4]
  assign _T_59887 = _T_59886[10:0]; // @[Modules.scala 50:57:@6537.4]
  assign buffer_1_537 = $signed(_T_59887); // @[Modules.scala 50:57:@6538.4]
  assign buffer_1_292 = {{6{_T_58977[4]}},_T_58977}; // @[Modules.scala 32:22:@8.4]
  assign _T_59889 = $signed(buffer_1_292) + $signed(buffer_0_293); // @[Modules.scala 50:57:@6540.4]
  assign _T_59890 = _T_59889[10:0]; // @[Modules.scala 50:57:@6541.4]
  assign buffer_1_538 = $signed(_T_59890); // @[Modules.scala 50:57:@6542.4]
  assign buffer_1_294 = {{6{_T_58991[4]}},_T_58991}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_295 = {{6{_T_58994[4]}},_T_58994}; // @[Modules.scala 32:22:@8.4]
  assign _T_59892 = $signed(buffer_1_294) + $signed(buffer_1_295); // @[Modules.scala 50:57:@6544.4]
  assign _T_59893 = _T_59892[10:0]; // @[Modules.scala 50:57:@6545.4]
  assign buffer_1_539 = $signed(_T_59893); // @[Modules.scala 50:57:@6546.4]
  assign buffer_1_296 = {{6{_T_58997[4]}},_T_58997}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_297 = {{6{_T_59000[4]}},_T_59000}; // @[Modules.scala 32:22:@8.4]
  assign _T_59895 = $signed(buffer_1_296) + $signed(buffer_1_297); // @[Modules.scala 50:57:@6548.4]
  assign _T_59896 = _T_59895[10:0]; // @[Modules.scala 50:57:@6549.4]
  assign buffer_1_540 = $signed(_T_59896); // @[Modules.scala 50:57:@6550.4]
  assign buffer_1_298 = {{6{_T_59003[4]}},_T_59003}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_299 = {{6{_T_59006[4]}},_T_59006}; // @[Modules.scala 32:22:@8.4]
  assign _T_59898 = $signed(buffer_1_298) + $signed(buffer_1_299); // @[Modules.scala 50:57:@6552.4]
  assign _T_59899 = _T_59898[10:0]; // @[Modules.scala 50:57:@6553.4]
  assign buffer_1_541 = $signed(_T_59899); // @[Modules.scala 50:57:@6554.4]
  assign buffer_1_301 = {{6{_T_59012[4]}},_T_59012}; // @[Modules.scala 32:22:@8.4]
  assign _T_59901 = $signed(buffer_0_300) + $signed(buffer_1_301); // @[Modules.scala 50:57:@6556.4]
  assign _T_59902 = _T_59901[10:0]; // @[Modules.scala 50:57:@6557.4]
  assign buffer_1_542 = $signed(_T_59902); // @[Modules.scala 50:57:@6558.4]
  assign buffer_1_306 = {{6{_T_59039[4]}},_T_59039}; // @[Modules.scala 32:22:@8.4]
  assign _T_59910 = $signed(buffer_1_306) + $signed(buffer_0_307); // @[Modules.scala 50:57:@6568.4]
  assign _T_59911 = _T_59910[10:0]; // @[Modules.scala 50:57:@6569.4]
  assign buffer_1_545 = $signed(_T_59911); // @[Modules.scala 50:57:@6570.4]
  assign buffer_1_308 = {{6{_T_59053[4]}},_T_59053}; // @[Modules.scala 32:22:@8.4]
  assign _T_59913 = $signed(buffer_1_308) + $signed(buffer_0_309); // @[Modules.scala 50:57:@6572.4]
  assign _T_59914 = _T_59913[10:0]; // @[Modules.scala 50:57:@6573.4]
  assign buffer_1_546 = $signed(_T_59914); // @[Modules.scala 50:57:@6574.4]
  assign buffer_1_310 = {{6{_T_59059[4]}},_T_59059}; // @[Modules.scala 32:22:@8.4]
  assign _T_59916 = $signed(buffer_1_310) + $signed(buffer_0_311); // @[Modules.scala 50:57:@6576.4]
  assign _T_59917 = _T_59916[10:0]; // @[Modules.scala 50:57:@6577.4]
  assign buffer_1_547 = $signed(_T_59917); // @[Modules.scala 50:57:@6578.4]
  assign buffer_1_312 = {{6{_T_59069[4]}},_T_59069}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_313 = {{6{_T_59072[4]}},_T_59072}; // @[Modules.scala 32:22:@8.4]
  assign _T_59919 = $signed(buffer_1_312) + $signed(buffer_1_313); // @[Modules.scala 50:57:@6580.4]
  assign _T_59920 = _T_59919[10:0]; // @[Modules.scala 50:57:@6581.4]
  assign buffer_1_548 = $signed(_T_59920); // @[Modules.scala 50:57:@6582.4]
  assign buffer_1_314 = {{6{_T_59075[4]}},_T_59075}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_315 = {{6{_T_59078[4]}},_T_59078}; // @[Modules.scala 32:22:@8.4]
  assign _T_59922 = $signed(buffer_1_314) + $signed(buffer_1_315); // @[Modules.scala 50:57:@6584.4]
  assign _T_59923 = _T_59922[10:0]; // @[Modules.scala 50:57:@6585.4]
  assign buffer_1_549 = $signed(_T_59923); // @[Modules.scala 50:57:@6586.4]
  assign buffer_1_316 = {{6{_T_59081[4]}},_T_59081}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_317 = {{6{_T_59084[4]}},_T_59084}; // @[Modules.scala 32:22:@8.4]
  assign _T_59925 = $signed(buffer_1_316) + $signed(buffer_1_317); // @[Modules.scala 50:57:@6588.4]
  assign _T_59926 = _T_59925[10:0]; // @[Modules.scala 50:57:@6589.4]
  assign buffer_1_550 = $signed(_T_59926); // @[Modules.scala 50:57:@6590.4]
  assign buffer_1_318 = {{6{_T_59087[4]}},_T_59087}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_319 = {{6{_T_59090[4]}},_T_59090}; // @[Modules.scala 32:22:@8.4]
  assign _T_59928 = $signed(buffer_1_318) + $signed(buffer_1_319); // @[Modules.scala 50:57:@6592.4]
  assign _T_59929 = _T_59928[10:0]; // @[Modules.scala 50:57:@6593.4]
  assign buffer_1_551 = $signed(_T_59929); // @[Modules.scala 50:57:@6594.4]
  assign buffer_1_320 = {{6{_T_59097[4]}},_T_59097}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_321 = {{6{_T_59100[4]}},_T_59100}; // @[Modules.scala 32:22:@8.4]
  assign _T_59931 = $signed(buffer_1_320) + $signed(buffer_1_321); // @[Modules.scala 50:57:@6596.4]
  assign _T_59932 = _T_59931[10:0]; // @[Modules.scala 50:57:@6597.4]
  assign buffer_1_552 = $signed(_T_59932); // @[Modules.scala 50:57:@6598.4]
  assign buffer_1_322 = {{6{_T_59107[4]}},_T_59107}; // @[Modules.scala 32:22:@8.4]
  assign _T_59934 = $signed(buffer_1_322) + $signed(buffer_0_323); // @[Modules.scala 50:57:@6600.4]
  assign _T_59935 = _T_59934[10:0]; // @[Modules.scala 50:57:@6601.4]
  assign buffer_1_553 = $signed(_T_59935); // @[Modules.scala 50:57:@6602.4]
  assign buffer_1_324 = {{6{_T_59113[4]}},_T_59113}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_325 = {{6{_T_59116[4]}},_T_59116}; // @[Modules.scala 32:22:@8.4]
  assign _T_59937 = $signed(buffer_1_324) + $signed(buffer_1_325); // @[Modules.scala 50:57:@6604.4]
  assign _T_59938 = _T_59937[10:0]; // @[Modules.scala 50:57:@6605.4]
  assign buffer_1_554 = $signed(_T_59938); // @[Modules.scala 50:57:@6606.4]
  assign buffer_1_326 = {{6{_T_59119[4]}},_T_59119}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_327 = {{6{_T_59122[4]}},_T_59122}; // @[Modules.scala 32:22:@8.4]
  assign _T_59940 = $signed(buffer_1_326) + $signed(buffer_1_327); // @[Modules.scala 50:57:@6608.4]
  assign _T_59941 = _T_59940[10:0]; // @[Modules.scala 50:57:@6609.4]
  assign buffer_1_555 = $signed(_T_59941); // @[Modules.scala 50:57:@6610.4]
  assign buffer_1_328 = {{6{_T_59125[4]}},_T_59125}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_329 = {{6{_T_59128[4]}},_T_59128}; // @[Modules.scala 32:22:@8.4]
  assign _T_59943 = $signed(buffer_1_328) + $signed(buffer_1_329); // @[Modules.scala 50:57:@6612.4]
  assign _T_59944 = _T_59943[10:0]; // @[Modules.scala 50:57:@6613.4]
  assign buffer_1_556 = $signed(_T_59944); // @[Modules.scala 50:57:@6614.4]
  assign buffer_1_331 = {{6{_T_59138[4]}},_T_59138}; // @[Modules.scala 32:22:@8.4]
  assign _T_59946 = $signed(buffer_0_330) + $signed(buffer_1_331); // @[Modules.scala 50:57:@6616.4]
  assign _T_59947 = _T_59946[10:0]; // @[Modules.scala 50:57:@6617.4]
  assign buffer_1_557 = $signed(_T_59947); // @[Modules.scala 50:57:@6618.4]
  assign buffer_1_332 = {{6{_T_59145[4]}},_T_59145}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_333 = {{6{_T_59152[4]}},_T_59152}; // @[Modules.scala 32:22:@8.4]
  assign _T_59949 = $signed(buffer_1_332) + $signed(buffer_1_333); // @[Modules.scala 50:57:@6620.4]
  assign _T_59950 = _T_59949[10:0]; // @[Modules.scala 50:57:@6621.4]
  assign buffer_1_558 = $signed(_T_59950); // @[Modules.scala 50:57:@6622.4]
  assign buffer_1_334 = {{6{_T_59159[4]}},_T_59159}; // @[Modules.scala 32:22:@8.4]
  assign _T_59952 = $signed(buffer_1_334) + $signed(buffer_0_335); // @[Modules.scala 50:57:@6624.4]
  assign _T_59953 = _T_59952[10:0]; // @[Modules.scala 50:57:@6625.4]
  assign buffer_1_559 = $signed(_T_59953); // @[Modules.scala 50:57:@6626.4]
  assign buffer_1_336 = {{6{_T_59173[4]}},_T_59173}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_337 = {{6{_T_59176[4]}},_T_59176}; // @[Modules.scala 32:22:@8.4]
  assign _T_59955 = $signed(buffer_1_336) + $signed(buffer_1_337); // @[Modules.scala 50:57:@6628.4]
  assign _T_59956 = _T_59955[10:0]; // @[Modules.scala 50:57:@6629.4]
  assign buffer_1_560 = $signed(_T_59956); // @[Modules.scala 50:57:@6630.4]
  assign buffer_1_340 = {{6{_T_59189[4]}},_T_59189}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_341 = {{6{_T_59192[4]}},_T_59192}; // @[Modules.scala 32:22:@8.4]
  assign _T_59961 = $signed(buffer_1_340) + $signed(buffer_1_341); // @[Modules.scala 50:57:@6636.4]
  assign _T_59962 = _T_59961[10:0]; // @[Modules.scala 50:57:@6637.4]
  assign buffer_1_562 = $signed(_T_59962); // @[Modules.scala 50:57:@6638.4]
  assign buffer_1_342 = {{6{_T_59195[4]}},_T_59195}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_343 = {{6{_T_59198[4]}},_T_59198}; // @[Modules.scala 32:22:@8.4]
  assign _T_59964 = $signed(buffer_1_342) + $signed(buffer_1_343); // @[Modules.scala 50:57:@6640.4]
  assign _T_59965 = _T_59964[10:0]; // @[Modules.scala 50:57:@6641.4]
  assign buffer_1_563 = $signed(_T_59965); // @[Modules.scala 50:57:@6642.4]
  assign buffer_1_344 = {{6{_T_59201[4]}},_T_59201}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_345 = {{6{_T_59204[4]}},_T_59204}; // @[Modules.scala 32:22:@8.4]
  assign _T_59967 = $signed(buffer_1_344) + $signed(buffer_1_345); // @[Modules.scala 50:57:@6644.4]
  assign _T_59968 = _T_59967[10:0]; // @[Modules.scala 50:57:@6645.4]
  assign buffer_1_564 = $signed(_T_59968); // @[Modules.scala 50:57:@6646.4]
  assign buffer_1_346 = {{6{_T_59211[4]}},_T_59211}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_347 = {{6{_T_59218[4]}},_T_59218}; // @[Modules.scala 32:22:@8.4]
  assign _T_59970 = $signed(buffer_1_346) + $signed(buffer_1_347); // @[Modules.scala 50:57:@6648.4]
  assign _T_59971 = _T_59970[10:0]; // @[Modules.scala 50:57:@6649.4]
  assign buffer_1_565 = $signed(_T_59971); // @[Modules.scala 50:57:@6650.4]
  assign buffer_1_348 = {{6{_T_59221[4]}},_T_59221}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_349 = {{6{_T_59228[4]}},_T_59228}; // @[Modules.scala 32:22:@8.4]
  assign _T_59973 = $signed(buffer_1_348) + $signed(buffer_1_349); // @[Modules.scala 50:57:@6652.4]
  assign _T_59974 = _T_59973[10:0]; // @[Modules.scala 50:57:@6653.4]
  assign buffer_1_566 = $signed(_T_59974); // @[Modules.scala 50:57:@6654.4]
  assign buffer_1_350 = {{6{_T_59231[4]}},_T_59231}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_351 = {{6{_T_59234[4]}},_T_59234}; // @[Modules.scala 32:22:@8.4]
  assign _T_59976 = $signed(buffer_1_350) + $signed(buffer_1_351); // @[Modules.scala 50:57:@6656.4]
  assign _T_59977 = _T_59976[10:0]; // @[Modules.scala 50:57:@6657.4]
  assign buffer_1_567 = $signed(_T_59977); // @[Modules.scala 50:57:@6658.4]
  assign buffer_1_354 = {{6{_T_59247[4]}},_T_59247}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_355 = {{6{_T_59254[4]}},_T_59254}; // @[Modules.scala 32:22:@8.4]
  assign _T_59982 = $signed(buffer_1_354) + $signed(buffer_1_355); // @[Modules.scala 50:57:@6664.4]
  assign _T_59983 = _T_59982[10:0]; // @[Modules.scala 50:57:@6665.4]
  assign buffer_1_569 = $signed(_T_59983); // @[Modules.scala 50:57:@6666.4]
  assign buffer_1_356 = {{6{_T_59261[4]}},_T_59261}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_357 = {{6{_T_59268[4]}},_T_59268}; // @[Modules.scala 32:22:@8.4]
  assign _T_59985 = $signed(buffer_1_356) + $signed(buffer_1_357); // @[Modules.scala 50:57:@6668.4]
  assign _T_59986 = _T_59985[10:0]; // @[Modules.scala 50:57:@6669.4]
  assign buffer_1_570 = $signed(_T_59986); // @[Modules.scala 50:57:@6670.4]
  assign buffer_1_358 = {{6{_T_59271[4]}},_T_59271}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_359 = {{6{_T_59278[4]}},_T_59278}; // @[Modules.scala 32:22:@8.4]
  assign _T_59988 = $signed(buffer_1_358) + $signed(buffer_1_359); // @[Modules.scala 50:57:@6672.4]
  assign _T_59989 = _T_59988[10:0]; // @[Modules.scala 50:57:@6673.4]
  assign buffer_1_571 = $signed(_T_59989); // @[Modules.scala 50:57:@6674.4]
  assign buffer_1_360 = {{6{_T_59285[4]}},_T_59285}; // @[Modules.scala 32:22:@8.4]
  assign _T_59991 = $signed(buffer_1_360) + $signed(buffer_0_361); // @[Modules.scala 50:57:@6676.4]
  assign _T_59992 = _T_59991[10:0]; // @[Modules.scala 50:57:@6677.4]
  assign buffer_1_572 = $signed(_T_59992); // @[Modules.scala 50:57:@6678.4]
  assign buffer_1_362 = {{6{_T_59291[4]}},_T_59291}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_363 = {{6{_T_59294[4]}},_T_59294}; // @[Modules.scala 32:22:@8.4]
  assign _T_59994 = $signed(buffer_1_362) + $signed(buffer_1_363); // @[Modules.scala 50:57:@6680.4]
  assign _T_59995 = _T_59994[10:0]; // @[Modules.scala 50:57:@6681.4]
  assign buffer_1_573 = $signed(_T_59995); // @[Modules.scala 50:57:@6682.4]
  assign buffer_1_364 = {{6{_T_59301[4]}},_T_59301}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_365 = {{6{_T_59308[4]}},_T_59308}; // @[Modules.scala 32:22:@8.4]
  assign _T_59997 = $signed(buffer_1_364) + $signed(buffer_1_365); // @[Modules.scala 50:57:@6684.4]
  assign _T_59998 = _T_59997[10:0]; // @[Modules.scala 50:57:@6685.4]
  assign buffer_1_574 = $signed(_T_59998); // @[Modules.scala 50:57:@6686.4]
  assign buffer_1_366 = {{6{_T_59315[4]}},_T_59315}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_367 = {{6{_T_59322[4]}},_T_59322}; // @[Modules.scala 32:22:@8.4]
  assign _T_60000 = $signed(buffer_1_366) + $signed(buffer_1_367); // @[Modules.scala 50:57:@6688.4]
  assign _T_60001 = _T_60000[10:0]; // @[Modules.scala 50:57:@6689.4]
  assign buffer_1_575 = $signed(_T_60001); // @[Modules.scala 50:57:@6690.4]
  assign buffer_1_370 = {{6{_T_59343[4]}},_T_59343}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_371 = {{6{_T_59350[4]}},_T_59350}; // @[Modules.scala 32:22:@8.4]
  assign _T_60006 = $signed(buffer_1_370) + $signed(buffer_1_371); // @[Modules.scala 50:57:@6696.4]
  assign _T_60007 = _T_60006[10:0]; // @[Modules.scala 50:57:@6697.4]
  assign buffer_1_577 = $signed(_T_60007); // @[Modules.scala 50:57:@6698.4]
  assign buffer_1_378 = {{6{_T_59379[4]}},_T_59379}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_379 = {{6{_T_59382[4]}},_T_59382}; // @[Modules.scala 32:22:@8.4]
  assign _T_60018 = $signed(buffer_1_378) + $signed(buffer_1_379); // @[Modules.scala 50:57:@6712.4]
  assign _T_60019 = _T_60018[10:0]; // @[Modules.scala 50:57:@6713.4]
  assign buffer_1_581 = $signed(_T_60019); // @[Modules.scala 50:57:@6714.4]
  assign buffer_1_380 = {{6{_T_59385[4]}},_T_59385}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_381 = {{6{_T_59388[4]}},_T_59388}; // @[Modules.scala 32:22:@8.4]
  assign _T_60021 = $signed(buffer_1_380) + $signed(buffer_1_381); // @[Modules.scala 50:57:@6716.4]
  assign _T_60022 = _T_60021[10:0]; // @[Modules.scala 50:57:@6717.4]
  assign buffer_1_582 = $signed(_T_60022); // @[Modules.scala 50:57:@6718.4]
  assign buffer_1_383 = {{6{_T_59398[4]}},_T_59398}; // @[Modules.scala 32:22:@8.4]
  assign _T_60024 = $signed(buffer_0_382) + $signed(buffer_1_383); // @[Modules.scala 50:57:@6720.4]
  assign _T_60025 = _T_60024[10:0]; // @[Modules.scala 50:57:@6721.4]
  assign buffer_1_583 = $signed(_T_60025); // @[Modules.scala 50:57:@6722.4]
  assign buffer_1_384 = {{6{_T_59405[4]}},_T_59405}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_385 = {{6{_T_59412[4]}},_T_59412}; // @[Modules.scala 32:22:@8.4]
  assign _T_60027 = $signed(buffer_1_384) + $signed(buffer_1_385); // @[Modules.scala 50:57:@6724.4]
  assign _T_60028 = _T_60027[10:0]; // @[Modules.scala 50:57:@6725.4]
  assign buffer_1_584 = $signed(_T_60028); // @[Modules.scala 50:57:@6726.4]
  assign buffer_1_388 = {{6{_T_59433[4]}},_T_59433}; // @[Modules.scala 32:22:@8.4]
  assign _T_60033 = $signed(buffer_1_388) + $signed(buffer_0_389); // @[Modules.scala 50:57:@6732.4]
  assign _T_60034 = _T_60033[10:0]; // @[Modules.scala 50:57:@6733.4]
  assign buffer_1_586 = $signed(_T_60034); // @[Modules.scala 50:57:@6734.4]
  assign buffer_1_390 = {{6{_T_59443[4]}},_T_59443}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_391 = {{6{_T_59450[4]}},_T_59450}; // @[Modules.scala 32:22:@8.4]
  assign _T_60036 = $signed(buffer_1_390) + $signed(buffer_1_391); // @[Modules.scala 50:57:@6736.4]
  assign _T_60037 = _T_60036[10:0]; // @[Modules.scala 50:57:@6737.4]
  assign buffer_1_587 = $signed(_T_60037); // @[Modules.scala 50:57:@6738.4]
  assign _T_60039 = $signed(buffer_1_392) + $signed(buffer_1_393); // @[Modules.scala 53:83:@6740.4]
  assign _T_60040 = _T_60039[10:0]; // @[Modules.scala 53:83:@6741.4]
  assign buffer_1_588 = $signed(_T_60040); // @[Modules.scala 53:83:@6742.4]
  assign _T_60042 = $signed(buffer_1_394) + $signed(buffer_1_395); // @[Modules.scala 53:83:@6744.4]
  assign _T_60043 = _T_60042[10:0]; // @[Modules.scala 53:83:@6745.4]
  assign buffer_1_589 = $signed(_T_60043); // @[Modules.scala 53:83:@6746.4]
  assign _T_60045 = $signed(buffer_1_396) + $signed(buffer_1_397); // @[Modules.scala 53:83:@6748.4]
  assign _T_60046 = _T_60045[10:0]; // @[Modules.scala 53:83:@6749.4]
  assign buffer_1_590 = $signed(_T_60046); // @[Modules.scala 53:83:@6750.4]
  assign _T_60048 = $signed(buffer_1_398) + $signed(buffer_1_399); // @[Modules.scala 53:83:@6752.4]
  assign _T_60049 = _T_60048[10:0]; // @[Modules.scala 53:83:@6753.4]
  assign buffer_1_591 = $signed(_T_60049); // @[Modules.scala 53:83:@6754.4]
  assign _T_60051 = $signed(buffer_1_400) + $signed(buffer_1_401); // @[Modules.scala 53:83:@6756.4]
  assign _T_60052 = _T_60051[10:0]; // @[Modules.scala 53:83:@6757.4]
  assign buffer_1_592 = $signed(_T_60052); // @[Modules.scala 53:83:@6758.4]
  assign _T_60054 = $signed(buffer_1_402) + $signed(buffer_1_403); // @[Modules.scala 53:83:@6760.4]
  assign _T_60055 = _T_60054[10:0]; // @[Modules.scala 53:83:@6761.4]
  assign buffer_1_593 = $signed(_T_60055); // @[Modules.scala 53:83:@6762.4]
  assign _T_60057 = $signed(buffer_1_404) + $signed(buffer_1_405); // @[Modules.scala 53:83:@6764.4]
  assign _T_60058 = _T_60057[10:0]; // @[Modules.scala 53:83:@6765.4]
  assign buffer_1_594 = $signed(_T_60058); // @[Modules.scala 53:83:@6766.4]
  assign _T_60060 = $signed(buffer_1_406) + $signed(buffer_1_407); // @[Modules.scala 53:83:@6768.4]
  assign _T_60061 = _T_60060[10:0]; // @[Modules.scala 53:83:@6769.4]
  assign buffer_1_595 = $signed(_T_60061); // @[Modules.scala 53:83:@6770.4]
  assign _T_60063 = $signed(buffer_1_408) + $signed(buffer_1_409); // @[Modules.scala 53:83:@6772.4]
  assign _T_60064 = _T_60063[10:0]; // @[Modules.scala 53:83:@6773.4]
  assign buffer_1_596 = $signed(_T_60064); // @[Modules.scala 53:83:@6774.4]
  assign _T_60066 = $signed(buffer_1_410) + $signed(buffer_1_411); // @[Modules.scala 53:83:@6776.4]
  assign _T_60067 = _T_60066[10:0]; // @[Modules.scala 53:83:@6777.4]
  assign buffer_1_597 = $signed(_T_60067); // @[Modules.scala 53:83:@6778.4]
  assign _T_60069 = $signed(buffer_1_412) + $signed(buffer_1_413); // @[Modules.scala 53:83:@6780.4]
  assign _T_60070 = _T_60069[10:0]; // @[Modules.scala 53:83:@6781.4]
  assign buffer_1_598 = $signed(_T_60070); // @[Modules.scala 53:83:@6782.4]
  assign _T_60072 = $signed(buffer_0_414) + $signed(buffer_1_415); // @[Modules.scala 53:83:@6784.4]
  assign _T_60073 = _T_60072[10:0]; // @[Modules.scala 53:83:@6785.4]
  assign buffer_1_599 = $signed(_T_60073); // @[Modules.scala 53:83:@6786.4]
  assign _T_60075 = $signed(buffer_1_416) + $signed(buffer_0_417); // @[Modules.scala 53:83:@6788.4]
  assign _T_60076 = _T_60075[10:0]; // @[Modules.scala 53:83:@6789.4]
  assign buffer_1_600 = $signed(_T_60076); // @[Modules.scala 53:83:@6790.4]
  assign _T_60078 = $signed(buffer_0_418) + $signed(buffer_1_419); // @[Modules.scala 53:83:@6792.4]
  assign _T_60079 = _T_60078[10:0]; // @[Modules.scala 53:83:@6793.4]
  assign buffer_1_601 = $signed(_T_60079); // @[Modules.scala 53:83:@6794.4]
  assign _T_60081 = $signed(buffer_1_420) + $signed(buffer_1_421); // @[Modules.scala 53:83:@6796.4]
  assign _T_60082 = _T_60081[10:0]; // @[Modules.scala 53:83:@6797.4]
  assign buffer_1_602 = $signed(_T_60082); // @[Modules.scala 53:83:@6798.4]
  assign _T_60084 = $signed(buffer_0_422) + $signed(buffer_1_423); // @[Modules.scala 53:83:@6800.4]
  assign _T_60085 = _T_60084[10:0]; // @[Modules.scala 53:83:@6801.4]
  assign buffer_1_603 = $signed(_T_60085); // @[Modules.scala 53:83:@6802.4]
  assign _T_60087 = $signed(buffer_1_424) + $signed(buffer_1_425); // @[Modules.scala 53:83:@6804.4]
  assign _T_60088 = _T_60087[10:0]; // @[Modules.scala 53:83:@6805.4]
  assign buffer_1_604 = $signed(_T_60088); // @[Modules.scala 53:83:@6806.4]
  assign _T_60090 = $signed(buffer_1_426) + $signed(buffer_1_427); // @[Modules.scala 53:83:@6808.4]
  assign _T_60091 = _T_60090[10:0]; // @[Modules.scala 53:83:@6809.4]
  assign buffer_1_605 = $signed(_T_60091); // @[Modules.scala 53:83:@6810.4]
  assign _T_60093 = $signed(buffer_1_428) + $signed(buffer_1_429); // @[Modules.scala 53:83:@6812.4]
  assign _T_60094 = _T_60093[10:0]; // @[Modules.scala 53:83:@6813.4]
  assign buffer_1_606 = $signed(_T_60094); // @[Modules.scala 53:83:@6814.4]
  assign _T_60096 = $signed(buffer_0_430) + $signed(buffer_1_431); // @[Modules.scala 53:83:@6816.4]
  assign _T_60097 = _T_60096[10:0]; // @[Modules.scala 53:83:@6817.4]
  assign buffer_1_607 = $signed(_T_60097); // @[Modules.scala 53:83:@6818.4]
  assign _T_60099 = $signed(buffer_1_432) + $signed(buffer_1_433); // @[Modules.scala 53:83:@6820.4]
  assign _T_60100 = _T_60099[10:0]; // @[Modules.scala 53:83:@6821.4]
  assign buffer_1_608 = $signed(_T_60100); // @[Modules.scala 53:83:@6822.4]
  assign _T_60102 = $signed(buffer_1_434) + $signed(buffer_1_435); // @[Modules.scala 53:83:@6824.4]
  assign _T_60103 = _T_60102[10:0]; // @[Modules.scala 53:83:@6825.4]
  assign buffer_1_609 = $signed(_T_60103); // @[Modules.scala 53:83:@6826.4]
  assign _T_60105 = $signed(buffer_1_436) + $signed(buffer_1_437); // @[Modules.scala 53:83:@6828.4]
  assign _T_60106 = _T_60105[10:0]; // @[Modules.scala 53:83:@6829.4]
  assign buffer_1_610 = $signed(_T_60106); // @[Modules.scala 53:83:@6830.4]
  assign _T_60108 = $signed(buffer_0_438) + $signed(buffer_1_439); // @[Modules.scala 53:83:@6832.4]
  assign _T_60109 = _T_60108[10:0]; // @[Modules.scala 53:83:@6833.4]
  assign buffer_1_611 = $signed(_T_60109); // @[Modules.scala 53:83:@6834.4]
  assign _T_60111 = $signed(buffer_1_440) + $signed(buffer_1_441); // @[Modules.scala 53:83:@6836.4]
  assign _T_60112 = _T_60111[10:0]; // @[Modules.scala 53:83:@6837.4]
  assign buffer_1_612 = $signed(_T_60112); // @[Modules.scala 53:83:@6838.4]
  assign _T_60114 = $signed(buffer_1_442) + $signed(buffer_1_443); // @[Modules.scala 53:83:@6840.4]
  assign _T_60115 = _T_60114[10:0]; // @[Modules.scala 53:83:@6841.4]
  assign buffer_1_613 = $signed(_T_60115); // @[Modules.scala 53:83:@6842.4]
  assign _T_60117 = $signed(buffer_1_444) + $signed(buffer_1_445); // @[Modules.scala 53:83:@6844.4]
  assign _T_60118 = _T_60117[10:0]; // @[Modules.scala 53:83:@6845.4]
  assign buffer_1_614 = $signed(_T_60118); // @[Modules.scala 53:83:@6846.4]
  assign _T_60120 = $signed(buffer_1_446) + $signed(buffer_1_447); // @[Modules.scala 53:83:@6848.4]
  assign _T_60121 = _T_60120[10:0]; // @[Modules.scala 53:83:@6849.4]
  assign buffer_1_615 = $signed(_T_60121); // @[Modules.scala 53:83:@6850.4]
  assign _T_60123 = $signed(buffer_1_448) + $signed(buffer_0_449); // @[Modules.scala 53:83:@6852.4]
  assign _T_60124 = _T_60123[10:0]; // @[Modules.scala 53:83:@6853.4]
  assign buffer_1_616 = $signed(_T_60124); // @[Modules.scala 53:83:@6854.4]
  assign _T_60126 = $signed(buffer_0_450) + $signed(buffer_1_451); // @[Modules.scala 53:83:@6856.4]
  assign _T_60127 = _T_60126[10:0]; // @[Modules.scala 53:83:@6857.4]
  assign buffer_1_617 = $signed(_T_60127); // @[Modules.scala 53:83:@6858.4]
  assign _T_60129 = $signed(buffer_1_452) + $signed(buffer_1_453); // @[Modules.scala 53:83:@6860.4]
  assign _T_60130 = _T_60129[10:0]; // @[Modules.scala 53:83:@6861.4]
  assign buffer_1_618 = $signed(_T_60130); // @[Modules.scala 53:83:@6862.4]
  assign _T_60132 = $signed(buffer_1_454) + $signed(buffer_1_455); // @[Modules.scala 53:83:@6864.4]
  assign _T_60133 = _T_60132[10:0]; // @[Modules.scala 53:83:@6865.4]
  assign buffer_1_619 = $signed(_T_60133); // @[Modules.scala 53:83:@6866.4]
  assign _T_60135 = $signed(buffer_0_456) + $signed(buffer_1_457); // @[Modules.scala 53:83:@6868.4]
  assign _T_60136 = _T_60135[10:0]; // @[Modules.scala 53:83:@6869.4]
  assign buffer_1_620 = $signed(_T_60136); // @[Modules.scala 53:83:@6870.4]
  assign _T_60138 = $signed(buffer_1_458) + $signed(buffer_0_459); // @[Modules.scala 53:83:@6872.4]
  assign _T_60139 = _T_60138[10:0]; // @[Modules.scala 53:83:@6873.4]
  assign buffer_1_621 = $signed(_T_60139); // @[Modules.scala 53:83:@6874.4]
  assign _T_60141 = $signed(buffer_1_460) + $signed(buffer_1_461); // @[Modules.scala 53:83:@6876.4]
  assign _T_60142 = _T_60141[10:0]; // @[Modules.scala 53:83:@6877.4]
  assign buffer_1_622 = $signed(_T_60142); // @[Modules.scala 53:83:@6878.4]
  assign _T_60144 = $signed(buffer_1_462) + $signed(buffer_0_463); // @[Modules.scala 53:83:@6880.4]
  assign _T_60145 = _T_60144[10:0]; // @[Modules.scala 53:83:@6881.4]
  assign buffer_1_623 = $signed(_T_60145); // @[Modules.scala 53:83:@6882.4]
  assign _T_60147 = $signed(buffer_0_464) + $signed(buffer_1_465); // @[Modules.scala 53:83:@6884.4]
  assign _T_60148 = _T_60147[10:0]; // @[Modules.scala 53:83:@6885.4]
  assign buffer_1_624 = $signed(_T_60148); // @[Modules.scala 53:83:@6886.4]
  assign _T_60150 = $signed(buffer_0_466) + $signed(buffer_1_467); // @[Modules.scala 53:83:@6888.4]
  assign _T_60151 = _T_60150[10:0]; // @[Modules.scala 53:83:@6889.4]
  assign buffer_1_625 = $signed(_T_60151); // @[Modules.scala 53:83:@6890.4]
  assign _T_60153 = $signed(buffer_1_468) + $signed(buffer_0_469); // @[Modules.scala 53:83:@6892.4]
  assign _T_60154 = _T_60153[10:0]; // @[Modules.scala 53:83:@6893.4]
  assign buffer_1_626 = $signed(_T_60154); // @[Modules.scala 53:83:@6894.4]
  assign _T_60156 = $signed(buffer_1_470) + $signed(buffer_1_471); // @[Modules.scala 53:83:@6896.4]
  assign _T_60157 = _T_60156[10:0]; // @[Modules.scala 53:83:@6897.4]
  assign buffer_1_627 = $signed(_T_60157); // @[Modules.scala 53:83:@6898.4]
  assign _T_60159 = $signed(buffer_1_472) + $signed(buffer_1_473); // @[Modules.scala 53:83:@6900.4]
  assign _T_60160 = _T_60159[10:0]; // @[Modules.scala 53:83:@6901.4]
  assign buffer_1_628 = $signed(_T_60160); // @[Modules.scala 53:83:@6902.4]
  assign _T_60162 = $signed(buffer_1_474) + $signed(buffer_1_475); // @[Modules.scala 53:83:@6904.4]
  assign _T_60163 = _T_60162[10:0]; // @[Modules.scala 53:83:@6905.4]
  assign buffer_1_629 = $signed(_T_60163); // @[Modules.scala 53:83:@6906.4]
  assign _T_60168 = $signed(buffer_0_478) + $signed(buffer_1_479); // @[Modules.scala 53:83:@6912.4]
  assign _T_60169 = _T_60168[10:0]; // @[Modules.scala 53:83:@6913.4]
  assign buffer_1_631 = $signed(_T_60169); // @[Modules.scala 53:83:@6914.4]
  assign _T_60171 = $signed(buffer_1_480) + $signed(buffer_1_481); // @[Modules.scala 53:83:@6916.4]
  assign _T_60172 = _T_60171[10:0]; // @[Modules.scala 53:83:@6917.4]
  assign buffer_1_632 = $signed(_T_60172); // @[Modules.scala 53:83:@6918.4]
  assign _T_60174 = $signed(buffer_1_482) + $signed(buffer_0_483); // @[Modules.scala 53:83:@6920.4]
  assign _T_60175 = _T_60174[10:0]; // @[Modules.scala 53:83:@6921.4]
  assign buffer_1_633 = $signed(_T_60175); // @[Modules.scala 53:83:@6922.4]
  assign _T_60177 = $signed(buffer_1_484) + $signed(buffer_0_485); // @[Modules.scala 53:83:@6924.4]
  assign _T_60178 = _T_60177[10:0]; // @[Modules.scala 53:83:@6925.4]
  assign buffer_1_634 = $signed(_T_60178); // @[Modules.scala 53:83:@6926.4]
  assign _T_60180 = $signed(buffer_1_486) + $signed(buffer_1_487); // @[Modules.scala 53:83:@6928.4]
  assign _T_60181 = _T_60180[10:0]; // @[Modules.scala 53:83:@6929.4]
  assign buffer_1_635 = $signed(_T_60181); // @[Modules.scala 53:83:@6930.4]
  assign _T_60183 = $signed(buffer_0_488) + $signed(buffer_1_489); // @[Modules.scala 53:83:@6932.4]
  assign _T_60184 = _T_60183[10:0]; // @[Modules.scala 53:83:@6933.4]
  assign buffer_1_636 = $signed(_T_60184); // @[Modules.scala 53:83:@6934.4]
  assign _T_60186 = $signed(buffer_1_490) + $signed(buffer_1_491); // @[Modules.scala 53:83:@6936.4]
  assign _T_60187 = _T_60186[10:0]; // @[Modules.scala 53:83:@6937.4]
  assign buffer_1_637 = $signed(_T_60187); // @[Modules.scala 53:83:@6938.4]
  assign _T_60189 = $signed(buffer_0_492) + $signed(buffer_1_493); // @[Modules.scala 53:83:@6940.4]
  assign _T_60190 = _T_60189[10:0]; // @[Modules.scala 53:83:@6941.4]
  assign buffer_1_638 = $signed(_T_60190); // @[Modules.scala 53:83:@6942.4]
  assign _T_60192 = $signed(buffer_1_494) + $signed(buffer_0_495); // @[Modules.scala 53:83:@6944.4]
  assign _T_60193 = _T_60192[10:0]; // @[Modules.scala 53:83:@6945.4]
  assign buffer_1_639 = $signed(_T_60193); // @[Modules.scala 53:83:@6946.4]
  assign _T_60195 = $signed(buffer_1_496) + $signed(buffer_1_497); // @[Modules.scala 53:83:@6948.4]
  assign _T_60196 = _T_60195[10:0]; // @[Modules.scala 53:83:@6949.4]
  assign buffer_1_640 = $signed(_T_60196); // @[Modules.scala 53:83:@6950.4]
  assign _T_60198 = $signed(buffer_1_498) + $signed(buffer_0_499); // @[Modules.scala 53:83:@6952.4]
  assign _T_60199 = _T_60198[10:0]; // @[Modules.scala 53:83:@6953.4]
  assign buffer_1_641 = $signed(_T_60199); // @[Modules.scala 53:83:@6954.4]
  assign _T_60201 = $signed(buffer_1_500) + $signed(buffer_1_501); // @[Modules.scala 53:83:@6956.4]
  assign _T_60202 = _T_60201[10:0]; // @[Modules.scala 53:83:@6957.4]
  assign buffer_1_642 = $signed(_T_60202); // @[Modules.scala 53:83:@6958.4]
  assign _T_60204 = $signed(buffer_1_502) + $signed(buffer_1_503); // @[Modules.scala 53:83:@6960.4]
  assign _T_60205 = _T_60204[10:0]; // @[Modules.scala 53:83:@6961.4]
  assign buffer_1_643 = $signed(_T_60205); // @[Modules.scala 53:83:@6962.4]
  assign _T_60207 = $signed(buffer_1_504) + $signed(buffer_1_505); // @[Modules.scala 53:83:@6964.4]
  assign _T_60208 = _T_60207[10:0]; // @[Modules.scala 53:83:@6965.4]
  assign buffer_1_644 = $signed(_T_60208); // @[Modules.scala 53:83:@6966.4]
  assign _T_60210 = $signed(buffer_1_506) + $signed(buffer_1_507); // @[Modules.scala 53:83:@6968.4]
  assign _T_60211 = _T_60210[10:0]; // @[Modules.scala 53:83:@6969.4]
  assign buffer_1_645 = $signed(_T_60211); // @[Modules.scala 53:83:@6970.4]
  assign _T_60213 = $signed(buffer_1_508) + $signed(buffer_1_509); // @[Modules.scala 53:83:@6972.4]
  assign _T_60214 = _T_60213[10:0]; // @[Modules.scala 53:83:@6973.4]
  assign buffer_1_646 = $signed(_T_60214); // @[Modules.scala 53:83:@6974.4]
  assign _T_60216 = $signed(buffer_1_510) + $signed(buffer_1_511); // @[Modules.scala 53:83:@6976.4]
  assign _T_60217 = _T_60216[10:0]; // @[Modules.scala 53:83:@6977.4]
  assign buffer_1_647 = $signed(_T_60217); // @[Modules.scala 53:83:@6978.4]
  assign _T_60219 = $signed(buffer_0_512) + $signed(buffer_1_513); // @[Modules.scala 53:83:@6980.4]
  assign _T_60220 = _T_60219[10:0]; // @[Modules.scala 53:83:@6981.4]
  assign buffer_1_648 = $signed(_T_60220); // @[Modules.scala 53:83:@6982.4]
  assign _T_60222 = $signed(buffer_1_514) + $signed(buffer_1_515); // @[Modules.scala 53:83:@6984.4]
  assign _T_60223 = _T_60222[10:0]; // @[Modules.scala 53:83:@6985.4]
  assign buffer_1_649 = $signed(_T_60223); // @[Modules.scala 53:83:@6986.4]
  assign _T_60225 = $signed(buffer_1_516) + $signed(buffer_0_517); // @[Modules.scala 53:83:@6988.4]
  assign _T_60226 = _T_60225[10:0]; // @[Modules.scala 53:83:@6989.4]
  assign buffer_1_650 = $signed(_T_60226); // @[Modules.scala 53:83:@6990.4]
  assign _T_60228 = $signed(buffer_1_518) + $signed(buffer_1_519); // @[Modules.scala 53:83:@6992.4]
  assign _T_60229 = _T_60228[10:0]; // @[Modules.scala 53:83:@6993.4]
  assign buffer_1_651 = $signed(_T_60229); // @[Modules.scala 53:83:@6994.4]
  assign _T_60231 = $signed(buffer_1_520) + $signed(buffer_1_521); // @[Modules.scala 53:83:@6996.4]
  assign _T_60232 = _T_60231[10:0]; // @[Modules.scala 53:83:@6997.4]
  assign buffer_1_652 = $signed(_T_60232); // @[Modules.scala 53:83:@6998.4]
  assign _T_60234 = $signed(buffer_1_522) + $signed(buffer_1_523); // @[Modules.scala 53:83:@7000.4]
  assign _T_60235 = _T_60234[10:0]; // @[Modules.scala 53:83:@7001.4]
  assign buffer_1_653 = $signed(_T_60235); // @[Modules.scala 53:83:@7002.4]
  assign _T_60237 = $signed(buffer_1_524) + $signed(buffer_1_525); // @[Modules.scala 53:83:@7004.4]
  assign _T_60238 = _T_60237[10:0]; // @[Modules.scala 53:83:@7005.4]
  assign buffer_1_654 = $signed(_T_60238); // @[Modules.scala 53:83:@7006.4]
  assign _T_60240 = $signed(buffer_1_526) + $signed(buffer_1_527); // @[Modules.scala 53:83:@7008.4]
  assign _T_60241 = _T_60240[10:0]; // @[Modules.scala 53:83:@7009.4]
  assign buffer_1_655 = $signed(_T_60241); // @[Modules.scala 53:83:@7010.4]
  assign _T_60243 = $signed(buffer_1_528) + $signed(buffer_1_529); // @[Modules.scala 53:83:@7012.4]
  assign _T_60244 = _T_60243[10:0]; // @[Modules.scala 53:83:@7013.4]
  assign buffer_1_656 = $signed(_T_60244); // @[Modules.scala 53:83:@7014.4]
  assign _T_60246 = $signed(buffer_1_530) + $signed(buffer_1_531); // @[Modules.scala 53:83:@7016.4]
  assign _T_60247 = _T_60246[10:0]; // @[Modules.scala 53:83:@7017.4]
  assign buffer_1_657 = $signed(_T_60247); // @[Modules.scala 53:83:@7018.4]
  assign _T_60249 = $signed(buffer_1_532) + $signed(buffer_1_533); // @[Modules.scala 53:83:@7020.4]
  assign _T_60250 = _T_60249[10:0]; // @[Modules.scala 53:83:@7021.4]
  assign buffer_1_658 = $signed(_T_60250); // @[Modules.scala 53:83:@7022.4]
  assign _T_60252 = $signed(buffer_1_534) + $signed(buffer_1_535); // @[Modules.scala 53:83:@7024.4]
  assign _T_60253 = _T_60252[10:0]; // @[Modules.scala 53:83:@7025.4]
  assign buffer_1_659 = $signed(_T_60253); // @[Modules.scala 53:83:@7026.4]
  assign _T_60255 = $signed(buffer_1_536) + $signed(buffer_1_537); // @[Modules.scala 53:83:@7028.4]
  assign _T_60256 = _T_60255[10:0]; // @[Modules.scala 53:83:@7029.4]
  assign buffer_1_660 = $signed(_T_60256); // @[Modules.scala 53:83:@7030.4]
  assign _T_60258 = $signed(buffer_1_538) + $signed(buffer_1_539); // @[Modules.scala 53:83:@7032.4]
  assign _T_60259 = _T_60258[10:0]; // @[Modules.scala 53:83:@7033.4]
  assign buffer_1_661 = $signed(_T_60259); // @[Modules.scala 53:83:@7034.4]
  assign _T_60261 = $signed(buffer_1_540) + $signed(buffer_1_541); // @[Modules.scala 53:83:@7036.4]
  assign _T_60262 = _T_60261[10:0]; // @[Modules.scala 53:83:@7037.4]
  assign buffer_1_662 = $signed(_T_60262); // @[Modules.scala 53:83:@7038.4]
  assign _T_60264 = $signed(buffer_1_542) + $signed(buffer_0_543); // @[Modules.scala 53:83:@7040.4]
  assign _T_60265 = _T_60264[10:0]; // @[Modules.scala 53:83:@7041.4]
  assign buffer_1_663 = $signed(_T_60265); // @[Modules.scala 53:83:@7042.4]
  assign _T_60267 = $signed(buffer_0_544) + $signed(buffer_1_545); // @[Modules.scala 53:83:@7044.4]
  assign _T_60268 = _T_60267[10:0]; // @[Modules.scala 53:83:@7045.4]
  assign buffer_1_664 = $signed(_T_60268); // @[Modules.scala 53:83:@7046.4]
  assign _T_60270 = $signed(buffer_1_546) + $signed(buffer_1_547); // @[Modules.scala 53:83:@7048.4]
  assign _T_60271 = _T_60270[10:0]; // @[Modules.scala 53:83:@7049.4]
  assign buffer_1_665 = $signed(_T_60271); // @[Modules.scala 53:83:@7050.4]
  assign _T_60273 = $signed(buffer_1_548) + $signed(buffer_1_549); // @[Modules.scala 53:83:@7052.4]
  assign _T_60274 = _T_60273[10:0]; // @[Modules.scala 53:83:@7053.4]
  assign buffer_1_666 = $signed(_T_60274); // @[Modules.scala 53:83:@7054.4]
  assign _T_60276 = $signed(buffer_1_550) + $signed(buffer_1_551); // @[Modules.scala 53:83:@7056.4]
  assign _T_60277 = _T_60276[10:0]; // @[Modules.scala 53:83:@7057.4]
  assign buffer_1_667 = $signed(_T_60277); // @[Modules.scala 53:83:@7058.4]
  assign _T_60279 = $signed(buffer_1_552) + $signed(buffer_1_553); // @[Modules.scala 53:83:@7060.4]
  assign _T_60280 = _T_60279[10:0]; // @[Modules.scala 53:83:@7061.4]
  assign buffer_1_668 = $signed(_T_60280); // @[Modules.scala 53:83:@7062.4]
  assign _T_60282 = $signed(buffer_1_554) + $signed(buffer_1_555); // @[Modules.scala 53:83:@7064.4]
  assign _T_60283 = _T_60282[10:0]; // @[Modules.scala 53:83:@7065.4]
  assign buffer_1_669 = $signed(_T_60283); // @[Modules.scala 53:83:@7066.4]
  assign _T_60285 = $signed(buffer_1_556) + $signed(buffer_1_557); // @[Modules.scala 53:83:@7068.4]
  assign _T_60286 = _T_60285[10:0]; // @[Modules.scala 53:83:@7069.4]
  assign buffer_1_670 = $signed(_T_60286); // @[Modules.scala 53:83:@7070.4]
  assign _T_60288 = $signed(buffer_1_558) + $signed(buffer_1_559); // @[Modules.scala 53:83:@7072.4]
  assign _T_60289 = _T_60288[10:0]; // @[Modules.scala 53:83:@7073.4]
  assign buffer_1_671 = $signed(_T_60289); // @[Modules.scala 53:83:@7074.4]
  assign _T_60291 = $signed(buffer_1_560) + $signed(buffer_0_561); // @[Modules.scala 53:83:@7076.4]
  assign _T_60292 = _T_60291[10:0]; // @[Modules.scala 53:83:@7077.4]
  assign buffer_1_672 = $signed(_T_60292); // @[Modules.scala 53:83:@7078.4]
  assign _T_60294 = $signed(buffer_1_562) + $signed(buffer_1_563); // @[Modules.scala 53:83:@7080.4]
  assign _T_60295 = _T_60294[10:0]; // @[Modules.scala 53:83:@7081.4]
  assign buffer_1_673 = $signed(_T_60295); // @[Modules.scala 53:83:@7082.4]
  assign _T_60297 = $signed(buffer_1_564) + $signed(buffer_1_565); // @[Modules.scala 53:83:@7084.4]
  assign _T_60298 = _T_60297[10:0]; // @[Modules.scala 53:83:@7085.4]
  assign buffer_1_674 = $signed(_T_60298); // @[Modules.scala 53:83:@7086.4]
  assign _T_60300 = $signed(buffer_1_566) + $signed(buffer_1_567); // @[Modules.scala 53:83:@7088.4]
  assign _T_60301 = _T_60300[10:0]; // @[Modules.scala 53:83:@7089.4]
  assign buffer_1_675 = $signed(_T_60301); // @[Modules.scala 53:83:@7090.4]
  assign _T_60303 = $signed(buffer_0_568) + $signed(buffer_1_569); // @[Modules.scala 53:83:@7092.4]
  assign _T_60304 = _T_60303[10:0]; // @[Modules.scala 53:83:@7093.4]
  assign buffer_1_676 = $signed(_T_60304); // @[Modules.scala 53:83:@7094.4]
  assign _T_60306 = $signed(buffer_1_570) + $signed(buffer_1_571); // @[Modules.scala 53:83:@7096.4]
  assign _T_60307 = _T_60306[10:0]; // @[Modules.scala 53:83:@7097.4]
  assign buffer_1_677 = $signed(_T_60307); // @[Modules.scala 53:83:@7098.4]
  assign _T_60309 = $signed(buffer_1_572) + $signed(buffer_1_573); // @[Modules.scala 53:83:@7100.4]
  assign _T_60310 = _T_60309[10:0]; // @[Modules.scala 53:83:@7101.4]
  assign buffer_1_678 = $signed(_T_60310); // @[Modules.scala 53:83:@7102.4]
  assign _T_60312 = $signed(buffer_1_574) + $signed(buffer_1_575); // @[Modules.scala 53:83:@7104.4]
  assign _T_60313 = _T_60312[10:0]; // @[Modules.scala 53:83:@7105.4]
  assign buffer_1_679 = $signed(_T_60313); // @[Modules.scala 53:83:@7106.4]
  assign _T_60315 = $signed(buffer_0_576) + $signed(buffer_1_577); // @[Modules.scala 53:83:@7108.4]
  assign _T_60316 = _T_60315[10:0]; // @[Modules.scala 53:83:@7109.4]
  assign buffer_1_680 = $signed(_T_60316); // @[Modules.scala 53:83:@7110.4]
  assign _T_60321 = $signed(buffer_0_580) + $signed(buffer_1_581); // @[Modules.scala 53:83:@7116.4]
  assign _T_60322 = _T_60321[10:0]; // @[Modules.scala 53:83:@7117.4]
  assign buffer_1_682 = $signed(_T_60322); // @[Modules.scala 53:83:@7118.4]
  assign _T_60324 = $signed(buffer_1_582) + $signed(buffer_1_583); // @[Modules.scala 53:83:@7120.4]
  assign _T_60325 = _T_60324[10:0]; // @[Modules.scala 53:83:@7121.4]
  assign buffer_1_683 = $signed(_T_60325); // @[Modules.scala 53:83:@7122.4]
  assign _T_60327 = $signed(buffer_1_584) + $signed(buffer_0_585); // @[Modules.scala 53:83:@7124.4]
  assign _T_60328 = _T_60327[10:0]; // @[Modules.scala 53:83:@7125.4]
  assign buffer_1_684 = $signed(_T_60328); // @[Modules.scala 53:83:@7126.4]
  assign _T_60330 = $signed(buffer_1_586) + $signed(buffer_1_587); // @[Modules.scala 53:83:@7128.4]
  assign _T_60331 = _T_60330[10:0]; // @[Modules.scala 53:83:@7129.4]
  assign buffer_1_685 = $signed(_T_60331); // @[Modules.scala 53:83:@7130.4]
  assign _T_60333 = $signed(buffer_1_588) + $signed(buffer_1_589); // @[Modules.scala 56:109:@7132.4]
  assign _T_60334 = _T_60333[10:0]; // @[Modules.scala 56:109:@7133.4]
  assign buffer_1_686 = $signed(_T_60334); // @[Modules.scala 56:109:@7134.4]
  assign _T_60336 = $signed(buffer_1_590) + $signed(buffer_1_591); // @[Modules.scala 56:109:@7136.4]
  assign _T_60337 = _T_60336[10:0]; // @[Modules.scala 56:109:@7137.4]
  assign buffer_1_687 = $signed(_T_60337); // @[Modules.scala 56:109:@7138.4]
  assign _T_60339 = $signed(buffer_1_592) + $signed(buffer_1_593); // @[Modules.scala 56:109:@7140.4]
  assign _T_60340 = _T_60339[10:0]; // @[Modules.scala 56:109:@7141.4]
  assign buffer_1_688 = $signed(_T_60340); // @[Modules.scala 56:109:@7142.4]
  assign _T_60342 = $signed(buffer_1_594) + $signed(buffer_1_595); // @[Modules.scala 56:109:@7144.4]
  assign _T_60343 = _T_60342[10:0]; // @[Modules.scala 56:109:@7145.4]
  assign buffer_1_689 = $signed(_T_60343); // @[Modules.scala 56:109:@7146.4]
  assign _T_60345 = $signed(buffer_1_596) + $signed(buffer_1_597); // @[Modules.scala 56:109:@7148.4]
  assign _T_60346 = _T_60345[10:0]; // @[Modules.scala 56:109:@7149.4]
  assign buffer_1_690 = $signed(_T_60346); // @[Modules.scala 56:109:@7150.4]
  assign _T_60348 = $signed(buffer_1_598) + $signed(buffer_1_599); // @[Modules.scala 56:109:@7152.4]
  assign _T_60349 = _T_60348[10:0]; // @[Modules.scala 56:109:@7153.4]
  assign buffer_1_691 = $signed(_T_60349); // @[Modules.scala 56:109:@7154.4]
  assign _T_60351 = $signed(buffer_1_600) + $signed(buffer_1_601); // @[Modules.scala 56:109:@7156.4]
  assign _T_60352 = _T_60351[10:0]; // @[Modules.scala 56:109:@7157.4]
  assign buffer_1_692 = $signed(_T_60352); // @[Modules.scala 56:109:@7158.4]
  assign _T_60354 = $signed(buffer_1_602) + $signed(buffer_1_603); // @[Modules.scala 56:109:@7160.4]
  assign _T_60355 = _T_60354[10:0]; // @[Modules.scala 56:109:@7161.4]
  assign buffer_1_693 = $signed(_T_60355); // @[Modules.scala 56:109:@7162.4]
  assign _T_60357 = $signed(buffer_1_604) + $signed(buffer_1_605); // @[Modules.scala 56:109:@7164.4]
  assign _T_60358 = _T_60357[10:0]; // @[Modules.scala 56:109:@7165.4]
  assign buffer_1_694 = $signed(_T_60358); // @[Modules.scala 56:109:@7166.4]
  assign _T_60360 = $signed(buffer_1_606) + $signed(buffer_1_607); // @[Modules.scala 56:109:@7168.4]
  assign _T_60361 = _T_60360[10:0]; // @[Modules.scala 56:109:@7169.4]
  assign buffer_1_695 = $signed(_T_60361); // @[Modules.scala 56:109:@7170.4]
  assign _T_60363 = $signed(buffer_1_608) + $signed(buffer_1_609); // @[Modules.scala 56:109:@7172.4]
  assign _T_60364 = _T_60363[10:0]; // @[Modules.scala 56:109:@7173.4]
  assign buffer_1_696 = $signed(_T_60364); // @[Modules.scala 56:109:@7174.4]
  assign _T_60366 = $signed(buffer_1_610) + $signed(buffer_1_611); // @[Modules.scala 56:109:@7176.4]
  assign _T_60367 = _T_60366[10:0]; // @[Modules.scala 56:109:@7177.4]
  assign buffer_1_697 = $signed(_T_60367); // @[Modules.scala 56:109:@7178.4]
  assign _T_60369 = $signed(buffer_1_612) + $signed(buffer_1_613); // @[Modules.scala 56:109:@7180.4]
  assign _T_60370 = _T_60369[10:0]; // @[Modules.scala 56:109:@7181.4]
  assign buffer_1_698 = $signed(_T_60370); // @[Modules.scala 56:109:@7182.4]
  assign _T_60372 = $signed(buffer_1_614) + $signed(buffer_1_615); // @[Modules.scala 56:109:@7184.4]
  assign _T_60373 = _T_60372[10:0]; // @[Modules.scala 56:109:@7185.4]
  assign buffer_1_699 = $signed(_T_60373); // @[Modules.scala 56:109:@7186.4]
  assign _T_60375 = $signed(buffer_1_616) + $signed(buffer_1_617); // @[Modules.scala 56:109:@7188.4]
  assign _T_60376 = _T_60375[10:0]; // @[Modules.scala 56:109:@7189.4]
  assign buffer_1_700 = $signed(_T_60376); // @[Modules.scala 56:109:@7190.4]
  assign _T_60378 = $signed(buffer_1_618) + $signed(buffer_1_619); // @[Modules.scala 56:109:@7192.4]
  assign _T_60379 = _T_60378[10:0]; // @[Modules.scala 56:109:@7193.4]
  assign buffer_1_701 = $signed(_T_60379); // @[Modules.scala 56:109:@7194.4]
  assign _T_60381 = $signed(buffer_1_620) + $signed(buffer_1_621); // @[Modules.scala 56:109:@7196.4]
  assign _T_60382 = _T_60381[10:0]; // @[Modules.scala 56:109:@7197.4]
  assign buffer_1_702 = $signed(_T_60382); // @[Modules.scala 56:109:@7198.4]
  assign _T_60384 = $signed(buffer_1_622) + $signed(buffer_1_623); // @[Modules.scala 56:109:@7200.4]
  assign _T_60385 = _T_60384[10:0]; // @[Modules.scala 56:109:@7201.4]
  assign buffer_1_703 = $signed(_T_60385); // @[Modules.scala 56:109:@7202.4]
  assign _T_60387 = $signed(buffer_1_624) + $signed(buffer_1_625); // @[Modules.scala 56:109:@7204.4]
  assign _T_60388 = _T_60387[10:0]; // @[Modules.scala 56:109:@7205.4]
  assign buffer_1_704 = $signed(_T_60388); // @[Modules.scala 56:109:@7206.4]
  assign _T_60390 = $signed(buffer_1_626) + $signed(buffer_1_627); // @[Modules.scala 56:109:@7208.4]
  assign _T_60391 = _T_60390[10:0]; // @[Modules.scala 56:109:@7209.4]
  assign buffer_1_705 = $signed(_T_60391); // @[Modules.scala 56:109:@7210.4]
  assign _T_60393 = $signed(buffer_1_628) + $signed(buffer_1_629); // @[Modules.scala 56:109:@7212.4]
  assign _T_60394 = _T_60393[10:0]; // @[Modules.scala 56:109:@7213.4]
  assign buffer_1_706 = $signed(_T_60394); // @[Modules.scala 56:109:@7214.4]
  assign _T_60396 = $signed(buffer_0_630) + $signed(buffer_1_631); // @[Modules.scala 56:109:@7216.4]
  assign _T_60397 = _T_60396[10:0]; // @[Modules.scala 56:109:@7217.4]
  assign buffer_1_707 = $signed(_T_60397); // @[Modules.scala 56:109:@7218.4]
  assign _T_60399 = $signed(buffer_1_632) + $signed(buffer_1_633); // @[Modules.scala 56:109:@7220.4]
  assign _T_60400 = _T_60399[10:0]; // @[Modules.scala 56:109:@7221.4]
  assign buffer_1_708 = $signed(_T_60400); // @[Modules.scala 56:109:@7222.4]
  assign _T_60402 = $signed(buffer_1_634) + $signed(buffer_1_635); // @[Modules.scala 56:109:@7224.4]
  assign _T_60403 = _T_60402[10:0]; // @[Modules.scala 56:109:@7225.4]
  assign buffer_1_709 = $signed(_T_60403); // @[Modules.scala 56:109:@7226.4]
  assign _T_60405 = $signed(buffer_1_636) + $signed(buffer_1_637); // @[Modules.scala 56:109:@7228.4]
  assign _T_60406 = _T_60405[10:0]; // @[Modules.scala 56:109:@7229.4]
  assign buffer_1_710 = $signed(_T_60406); // @[Modules.scala 56:109:@7230.4]
  assign _T_60408 = $signed(buffer_1_638) + $signed(buffer_1_639); // @[Modules.scala 56:109:@7232.4]
  assign _T_60409 = _T_60408[10:0]; // @[Modules.scala 56:109:@7233.4]
  assign buffer_1_711 = $signed(_T_60409); // @[Modules.scala 56:109:@7234.4]
  assign _T_60411 = $signed(buffer_1_640) + $signed(buffer_1_641); // @[Modules.scala 56:109:@7236.4]
  assign _T_60412 = _T_60411[10:0]; // @[Modules.scala 56:109:@7237.4]
  assign buffer_1_712 = $signed(_T_60412); // @[Modules.scala 56:109:@7238.4]
  assign _T_60414 = $signed(buffer_1_642) + $signed(buffer_1_643); // @[Modules.scala 56:109:@7240.4]
  assign _T_60415 = _T_60414[10:0]; // @[Modules.scala 56:109:@7241.4]
  assign buffer_1_713 = $signed(_T_60415); // @[Modules.scala 56:109:@7242.4]
  assign _T_60417 = $signed(buffer_1_644) + $signed(buffer_1_645); // @[Modules.scala 56:109:@7244.4]
  assign _T_60418 = _T_60417[10:0]; // @[Modules.scala 56:109:@7245.4]
  assign buffer_1_714 = $signed(_T_60418); // @[Modules.scala 56:109:@7246.4]
  assign _T_60420 = $signed(buffer_1_646) + $signed(buffer_1_647); // @[Modules.scala 56:109:@7248.4]
  assign _T_60421 = _T_60420[10:0]; // @[Modules.scala 56:109:@7249.4]
  assign buffer_1_715 = $signed(_T_60421); // @[Modules.scala 56:109:@7250.4]
  assign _T_60423 = $signed(buffer_1_648) + $signed(buffer_1_649); // @[Modules.scala 56:109:@7252.4]
  assign _T_60424 = _T_60423[10:0]; // @[Modules.scala 56:109:@7253.4]
  assign buffer_1_716 = $signed(_T_60424); // @[Modules.scala 56:109:@7254.4]
  assign _T_60426 = $signed(buffer_1_650) + $signed(buffer_1_651); // @[Modules.scala 56:109:@7256.4]
  assign _T_60427 = _T_60426[10:0]; // @[Modules.scala 56:109:@7257.4]
  assign buffer_1_717 = $signed(_T_60427); // @[Modules.scala 56:109:@7258.4]
  assign _T_60429 = $signed(buffer_1_652) + $signed(buffer_1_653); // @[Modules.scala 56:109:@7260.4]
  assign _T_60430 = _T_60429[10:0]; // @[Modules.scala 56:109:@7261.4]
  assign buffer_1_718 = $signed(_T_60430); // @[Modules.scala 56:109:@7262.4]
  assign _T_60432 = $signed(buffer_1_654) + $signed(buffer_1_655); // @[Modules.scala 56:109:@7264.4]
  assign _T_60433 = _T_60432[10:0]; // @[Modules.scala 56:109:@7265.4]
  assign buffer_1_719 = $signed(_T_60433); // @[Modules.scala 56:109:@7266.4]
  assign _T_60435 = $signed(buffer_1_656) + $signed(buffer_1_657); // @[Modules.scala 56:109:@7268.4]
  assign _T_60436 = _T_60435[10:0]; // @[Modules.scala 56:109:@7269.4]
  assign buffer_1_720 = $signed(_T_60436); // @[Modules.scala 56:109:@7270.4]
  assign _T_60438 = $signed(buffer_1_658) + $signed(buffer_1_659); // @[Modules.scala 56:109:@7272.4]
  assign _T_60439 = _T_60438[10:0]; // @[Modules.scala 56:109:@7273.4]
  assign buffer_1_721 = $signed(_T_60439); // @[Modules.scala 56:109:@7274.4]
  assign _T_60441 = $signed(buffer_1_660) + $signed(buffer_1_661); // @[Modules.scala 56:109:@7276.4]
  assign _T_60442 = _T_60441[10:0]; // @[Modules.scala 56:109:@7277.4]
  assign buffer_1_722 = $signed(_T_60442); // @[Modules.scala 56:109:@7278.4]
  assign _T_60444 = $signed(buffer_1_662) + $signed(buffer_1_663); // @[Modules.scala 56:109:@7280.4]
  assign _T_60445 = _T_60444[10:0]; // @[Modules.scala 56:109:@7281.4]
  assign buffer_1_723 = $signed(_T_60445); // @[Modules.scala 56:109:@7282.4]
  assign _T_60447 = $signed(buffer_1_664) + $signed(buffer_1_665); // @[Modules.scala 56:109:@7284.4]
  assign _T_60448 = _T_60447[10:0]; // @[Modules.scala 56:109:@7285.4]
  assign buffer_1_724 = $signed(_T_60448); // @[Modules.scala 56:109:@7286.4]
  assign _T_60450 = $signed(buffer_1_666) + $signed(buffer_1_667); // @[Modules.scala 56:109:@7288.4]
  assign _T_60451 = _T_60450[10:0]; // @[Modules.scala 56:109:@7289.4]
  assign buffer_1_725 = $signed(_T_60451); // @[Modules.scala 56:109:@7290.4]
  assign _T_60453 = $signed(buffer_1_668) + $signed(buffer_1_669); // @[Modules.scala 56:109:@7292.4]
  assign _T_60454 = _T_60453[10:0]; // @[Modules.scala 56:109:@7293.4]
  assign buffer_1_726 = $signed(_T_60454); // @[Modules.scala 56:109:@7294.4]
  assign _T_60456 = $signed(buffer_1_670) + $signed(buffer_1_671); // @[Modules.scala 56:109:@7296.4]
  assign _T_60457 = _T_60456[10:0]; // @[Modules.scala 56:109:@7297.4]
  assign buffer_1_727 = $signed(_T_60457); // @[Modules.scala 56:109:@7298.4]
  assign _T_60459 = $signed(buffer_1_672) + $signed(buffer_1_673); // @[Modules.scala 56:109:@7300.4]
  assign _T_60460 = _T_60459[10:0]; // @[Modules.scala 56:109:@7301.4]
  assign buffer_1_728 = $signed(_T_60460); // @[Modules.scala 56:109:@7302.4]
  assign _T_60462 = $signed(buffer_1_674) + $signed(buffer_1_675); // @[Modules.scala 56:109:@7304.4]
  assign _T_60463 = _T_60462[10:0]; // @[Modules.scala 56:109:@7305.4]
  assign buffer_1_729 = $signed(_T_60463); // @[Modules.scala 56:109:@7306.4]
  assign _T_60465 = $signed(buffer_1_676) + $signed(buffer_1_677); // @[Modules.scala 56:109:@7308.4]
  assign _T_60466 = _T_60465[10:0]; // @[Modules.scala 56:109:@7309.4]
  assign buffer_1_730 = $signed(_T_60466); // @[Modules.scala 56:109:@7310.4]
  assign _T_60468 = $signed(buffer_1_678) + $signed(buffer_1_679); // @[Modules.scala 56:109:@7312.4]
  assign _T_60469 = _T_60468[10:0]; // @[Modules.scala 56:109:@7313.4]
  assign buffer_1_731 = $signed(_T_60469); // @[Modules.scala 56:109:@7314.4]
  assign _T_60471 = $signed(buffer_1_680) + $signed(buffer_0_681); // @[Modules.scala 56:109:@7316.4]
  assign _T_60472 = _T_60471[10:0]; // @[Modules.scala 56:109:@7317.4]
  assign buffer_1_732 = $signed(_T_60472); // @[Modules.scala 56:109:@7318.4]
  assign _T_60474 = $signed(buffer_1_682) + $signed(buffer_1_683); // @[Modules.scala 56:109:@7320.4]
  assign _T_60475 = _T_60474[10:0]; // @[Modules.scala 56:109:@7321.4]
  assign buffer_1_733 = $signed(_T_60475); // @[Modules.scala 56:109:@7322.4]
  assign _T_60477 = $signed(buffer_1_684) + $signed(buffer_1_685); // @[Modules.scala 56:109:@7324.4]
  assign _T_60478 = _T_60477[10:0]; // @[Modules.scala 56:109:@7325.4]
  assign buffer_1_734 = $signed(_T_60478); // @[Modules.scala 56:109:@7326.4]
  assign _T_60480 = $signed(buffer_1_686) + $signed(buffer_1_687); // @[Modules.scala 63:156:@7329.4]
  assign _T_60481 = _T_60480[10:0]; // @[Modules.scala 63:156:@7330.4]
  assign buffer_1_736 = $signed(_T_60481); // @[Modules.scala 63:156:@7331.4]
  assign _T_60483 = $signed(buffer_1_736) + $signed(buffer_1_688); // @[Modules.scala 63:156:@7333.4]
  assign _T_60484 = _T_60483[10:0]; // @[Modules.scala 63:156:@7334.4]
  assign buffer_1_737 = $signed(_T_60484); // @[Modules.scala 63:156:@7335.4]
  assign _T_60486 = $signed(buffer_1_737) + $signed(buffer_1_689); // @[Modules.scala 63:156:@7337.4]
  assign _T_60487 = _T_60486[10:0]; // @[Modules.scala 63:156:@7338.4]
  assign buffer_1_738 = $signed(_T_60487); // @[Modules.scala 63:156:@7339.4]
  assign _T_60489 = $signed(buffer_1_738) + $signed(buffer_1_690); // @[Modules.scala 63:156:@7341.4]
  assign _T_60490 = _T_60489[10:0]; // @[Modules.scala 63:156:@7342.4]
  assign buffer_1_739 = $signed(_T_60490); // @[Modules.scala 63:156:@7343.4]
  assign _T_60492 = $signed(buffer_1_739) + $signed(buffer_1_691); // @[Modules.scala 63:156:@7345.4]
  assign _T_60493 = _T_60492[10:0]; // @[Modules.scala 63:156:@7346.4]
  assign buffer_1_740 = $signed(_T_60493); // @[Modules.scala 63:156:@7347.4]
  assign _T_60495 = $signed(buffer_1_740) + $signed(buffer_1_692); // @[Modules.scala 63:156:@7349.4]
  assign _T_60496 = _T_60495[10:0]; // @[Modules.scala 63:156:@7350.4]
  assign buffer_1_741 = $signed(_T_60496); // @[Modules.scala 63:156:@7351.4]
  assign _T_60498 = $signed(buffer_1_741) + $signed(buffer_1_693); // @[Modules.scala 63:156:@7353.4]
  assign _T_60499 = _T_60498[10:0]; // @[Modules.scala 63:156:@7354.4]
  assign buffer_1_742 = $signed(_T_60499); // @[Modules.scala 63:156:@7355.4]
  assign _T_60501 = $signed(buffer_1_742) + $signed(buffer_1_694); // @[Modules.scala 63:156:@7357.4]
  assign _T_60502 = _T_60501[10:0]; // @[Modules.scala 63:156:@7358.4]
  assign buffer_1_743 = $signed(_T_60502); // @[Modules.scala 63:156:@7359.4]
  assign _T_60504 = $signed(buffer_1_743) + $signed(buffer_1_695); // @[Modules.scala 63:156:@7361.4]
  assign _T_60505 = _T_60504[10:0]; // @[Modules.scala 63:156:@7362.4]
  assign buffer_1_744 = $signed(_T_60505); // @[Modules.scala 63:156:@7363.4]
  assign _T_60507 = $signed(buffer_1_744) + $signed(buffer_1_696); // @[Modules.scala 63:156:@7365.4]
  assign _T_60508 = _T_60507[10:0]; // @[Modules.scala 63:156:@7366.4]
  assign buffer_1_745 = $signed(_T_60508); // @[Modules.scala 63:156:@7367.4]
  assign _T_60510 = $signed(buffer_1_745) + $signed(buffer_1_697); // @[Modules.scala 63:156:@7369.4]
  assign _T_60511 = _T_60510[10:0]; // @[Modules.scala 63:156:@7370.4]
  assign buffer_1_746 = $signed(_T_60511); // @[Modules.scala 63:156:@7371.4]
  assign _T_60513 = $signed(buffer_1_746) + $signed(buffer_1_698); // @[Modules.scala 63:156:@7373.4]
  assign _T_60514 = _T_60513[10:0]; // @[Modules.scala 63:156:@7374.4]
  assign buffer_1_747 = $signed(_T_60514); // @[Modules.scala 63:156:@7375.4]
  assign _T_60516 = $signed(buffer_1_747) + $signed(buffer_1_699); // @[Modules.scala 63:156:@7377.4]
  assign _T_60517 = _T_60516[10:0]; // @[Modules.scala 63:156:@7378.4]
  assign buffer_1_748 = $signed(_T_60517); // @[Modules.scala 63:156:@7379.4]
  assign _T_60519 = $signed(buffer_1_748) + $signed(buffer_1_700); // @[Modules.scala 63:156:@7381.4]
  assign _T_60520 = _T_60519[10:0]; // @[Modules.scala 63:156:@7382.4]
  assign buffer_1_749 = $signed(_T_60520); // @[Modules.scala 63:156:@7383.4]
  assign _T_60522 = $signed(buffer_1_749) + $signed(buffer_1_701); // @[Modules.scala 63:156:@7385.4]
  assign _T_60523 = _T_60522[10:0]; // @[Modules.scala 63:156:@7386.4]
  assign buffer_1_750 = $signed(_T_60523); // @[Modules.scala 63:156:@7387.4]
  assign _T_60525 = $signed(buffer_1_750) + $signed(buffer_1_702); // @[Modules.scala 63:156:@7389.4]
  assign _T_60526 = _T_60525[10:0]; // @[Modules.scala 63:156:@7390.4]
  assign buffer_1_751 = $signed(_T_60526); // @[Modules.scala 63:156:@7391.4]
  assign _T_60528 = $signed(buffer_1_751) + $signed(buffer_1_703); // @[Modules.scala 63:156:@7393.4]
  assign _T_60529 = _T_60528[10:0]; // @[Modules.scala 63:156:@7394.4]
  assign buffer_1_752 = $signed(_T_60529); // @[Modules.scala 63:156:@7395.4]
  assign _T_60531 = $signed(buffer_1_752) + $signed(buffer_1_704); // @[Modules.scala 63:156:@7397.4]
  assign _T_60532 = _T_60531[10:0]; // @[Modules.scala 63:156:@7398.4]
  assign buffer_1_753 = $signed(_T_60532); // @[Modules.scala 63:156:@7399.4]
  assign _T_60534 = $signed(buffer_1_753) + $signed(buffer_1_705); // @[Modules.scala 63:156:@7401.4]
  assign _T_60535 = _T_60534[10:0]; // @[Modules.scala 63:156:@7402.4]
  assign buffer_1_754 = $signed(_T_60535); // @[Modules.scala 63:156:@7403.4]
  assign _T_60537 = $signed(buffer_1_754) + $signed(buffer_1_706); // @[Modules.scala 63:156:@7405.4]
  assign _T_60538 = _T_60537[10:0]; // @[Modules.scala 63:156:@7406.4]
  assign buffer_1_755 = $signed(_T_60538); // @[Modules.scala 63:156:@7407.4]
  assign _T_60540 = $signed(buffer_1_755) + $signed(buffer_1_707); // @[Modules.scala 63:156:@7409.4]
  assign _T_60541 = _T_60540[10:0]; // @[Modules.scala 63:156:@7410.4]
  assign buffer_1_756 = $signed(_T_60541); // @[Modules.scala 63:156:@7411.4]
  assign _T_60543 = $signed(buffer_1_756) + $signed(buffer_1_708); // @[Modules.scala 63:156:@7413.4]
  assign _T_60544 = _T_60543[10:0]; // @[Modules.scala 63:156:@7414.4]
  assign buffer_1_757 = $signed(_T_60544); // @[Modules.scala 63:156:@7415.4]
  assign _T_60546 = $signed(buffer_1_757) + $signed(buffer_1_709); // @[Modules.scala 63:156:@7417.4]
  assign _T_60547 = _T_60546[10:0]; // @[Modules.scala 63:156:@7418.4]
  assign buffer_1_758 = $signed(_T_60547); // @[Modules.scala 63:156:@7419.4]
  assign _T_60549 = $signed(buffer_1_758) + $signed(buffer_1_710); // @[Modules.scala 63:156:@7421.4]
  assign _T_60550 = _T_60549[10:0]; // @[Modules.scala 63:156:@7422.4]
  assign buffer_1_759 = $signed(_T_60550); // @[Modules.scala 63:156:@7423.4]
  assign _T_60552 = $signed(buffer_1_759) + $signed(buffer_1_711); // @[Modules.scala 63:156:@7425.4]
  assign _T_60553 = _T_60552[10:0]; // @[Modules.scala 63:156:@7426.4]
  assign buffer_1_760 = $signed(_T_60553); // @[Modules.scala 63:156:@7427.4]
  assign _T_60555 = $signed(buffer_1_760) + $signed(buffer_1_712); // @[Modules.scala 63:156:@7429.4]
  assign _T_60556 = _T_60555[10:0]; // @[Modules.scala 63:156:@7430.4]
  assign buffer_1_761 = $signed(_T_60556); // @[Modules.scala 63:156:@7431.4]
  assign _T_60558 = $signed(buffer_1_761) + $signed(buffer_1_713); // @[Modules.scala 63:156:@7433.4]
  assign _T_60559 = _T_60558[10:0]; // @[Modules.scala 63:156:@7434.4]
  assign buffer_1_762 = $signed(_T_60559); // @[Modules.scala 63:156:@7435.4]
  assign _T_60561 = $signed(buffer_1_762) + $signed(buffer_1_714); // @[Modules.scala 63:156:@7437.4]
  assign _T_60562 = _T_60561[10:0]; // @[Modules.scala 63:156:@7438.4]
  assign buffer_1_763 = $signed(_T_60562); // @[Modules.scala 63:156:@7439.4]
  assign _T_60564 = $signed(buffer_1_763) + $signed(buffer_1_715); // @[Modules.scala 63:156:@7441.4]
  assign _T_60565 = _T_60564[10:0]; // @[Modules.scala 63:156:@7442.4]
  assign buffer_1_764 = $signed(_T_60565); // @[Modules.scala 63:156:@7443.4]
  assign _T_60567 = $signed(buffer_1_764) + $signed(buffer_1_716); // @[Modules.scala 63:156:@7445.4]
  assign _T_60568 = _T_60567[10:0]; // @[Modules.scala 63:156:@7446.4]
  assign buffer_1_765 = $signed(_T_60568); // @[Modules.scala 63:156:@7447.4]
  assign _T_60570 = $signed(buffer_1_765) + $signed(buffer_1_717); // @[Modules.scala 63:156:@7449.4]
  assign _T_60571 = _T_60570[10:0]; // @[Modules.scala 63:156:@7450.4]
  assign buffer_1_766 = $signed(_T_60571); // @[Modules.scala 63:156:@7451.4]
  assign _T_60573 = $signed(buffer_1_766) + $signed(buffer_1_718); // @[Modules.scala 63:156:@7453.4]
  assign _T_60574 = _T_60573[10:0]; // @[Modules.scala 63:156:@7454.4]
  assign buffer_1_767 = $signed(_T_60574); // @[Modules.scala 63:156:@7455.4]
  assign _T_60576 = $signed(buffer_1_767) + $signed(buffer_1_719); // @[Modules.scala 63:156:@7457.4]
  assign _T_60577 = _T_60576[10:0]; // @[Modules.scala 63:156:@7458.4]
  assign buffer_1_768 = $signed(_T_60577); // @[Modules.scala 63:156:@7459.4]
  assign _T_60579 = $signed(buffer_1_768) + $signed(buffer_1_720); // @[Modules.scala 63:156:@7461.4]
  assign _T_60580 = _T_60579[10:0]; // @[Modules.scala 63:156:@7462.4]
  assign buffer_1_769 = $signed(_T_60580); // @[Modules.scala 63:156:@7463.4]
  assign _T_60582 = $signed(buffer_1_769) + $signed(buffer_1_721); // @[Modules.scala 63:156:@7465.4]
  assign _T_60583 = _T_60582[10:0]; // @[Modules.scala 63:156:@7466.4]
  assign buffer_1_770 = $signed(_T_60583); // @[Modules.scala 63:156:@7467.4]
  assign _T_60585 = $signed(buffer_1_770) + $signed(buffer_1_722); // @[Modules.scala 63:156:@7469.4]
  assign _T_60586 = _T_60585[10:0]; // @[Modules.scala 63:156:@7470.4]
  assign buffer_1_771 = $signed(_T_60586); // @[Modules.scala 63:156:@7471.4]
  assign _T_60588 = $signed(buffer_1_771) + $signed(buffer_1_723); // @[Modules.scala 63:156:@7473.4]
  assign _T_60589 = _T_60588[10:0]; // @[Modules.scala 63:156:@7474.4]
  assign buffer_1_772 = $signed(_T_60589); // @[Modules.scala 63:156:@7475.4]
  assign _T_60591 = $signed(buffer_1_772) + $signed(buffer_1_724); // @[Modules.scala 63:156:@7477.4]
  assign _T_60592 = _T_60591[10:0]; // @[Modules.scala 63:156:@7478.4]
  assign buffer_1_773 = $signed(_T_60592); // @[Modules.scala 63:156:@7479.4]
  assign _T_60594 = $signed(buffer_1_773) + $signed(buffer_1_725); // @[Modules.scala 63:156:@7481.4]
  assign _T_60595 = _T_60594[10:0]; // @[Modules.scala 63:156:@7482.4]
  assign buffer_1_774 = $signed(_T_60595); // @[Modules.scala 63:156:@7483.4]
  assign _T_60597 = $signed(buffer_1_774) + $signed(buffer_1_726); // @[Modules.scala 63:156:@7485.4]
  assign _T_60598 = _T_60597[10:0]; // @[Modules.scala 63:156:@7486.4]
  assign buffer_1_775 = $signed(_T_60598); // @[Modules.scala 63:156:@7487.4]
  assign _T_60600 = $signed(buffer_1_775) + $signed(buffer_1_727); // @[Modules.scala 63:156:@7489.4]
  assign _T_60601 = _T_60600[10:0]; // @[Modules.scala 63:156:@7490.4]
  assign buffer_1_776 = $signed(_T_60601); // @[Modules.scala 63:156:@7491.4]
  assign _T_60603 = $signed(buffer_1_776) + $signed(buffer_1_728); // @[Modules.scala 63:156:@7493.4]
  assign _T_60604 = _T_60603[10:0]; // @[Modules.scala 63:156:@7494.4]
  assign buffer_1_777 = $signed(_T_60604); // @[Modules.scala 63:156:@7495.4]
  assign _T_60606 = $signed(buffer_1_777) + $signed(buffer_1_729); // @[Modules.scala 63:156:@7497.4]
  assign _T_60607 = _T_60606[10:0]; // @[Modules.scala 63:156:@7498.4]
  assign buffer_1_778 = $signed(_T_60607); // @[Modules.scala 63:156:@7499.4]
  assign _T_60609 = $signed(buffer_1_778) + $signed(buffer_1_730); // @[Modules.scala 63:156:@7501.4]
  assign _T_60610 = _T_60609[10:0]; // @[Modules.scala 63:156:@7502.4]
  assign buffer_1_779 = $signed(_T_60610); // @[Modules.scala 63:156:@7503.4]
  assign _T_60612 = $signed(buffer_1_779) + $signed(buffer_1_731); // @[Modules.scala 63:156:@7505.4]
  assign _T_60613 = _T_60612[10:0]; // @[Modules.scala 63:156:@7506.4]
  assign buffer_1_780 = $signed(_T_60613); // @[Modules.scala 63:156:@7507.4]
  assign _T_60615 = $signed(buffer_1_780) + $signed(buffer_1_732); // @[Modules.scala 63:156:@7509.4]
  assign _T_60616 = _T_60615[10:0]; // @[Modules.scala 63:156:@7510.4]
  assign buffer_1_781 = $signed(_T_60616); // @[Modules.scala 63:156:@7511.4]
  assign _T_60618 = $signed(buffer_1_781) + $signed(buffer_1_733); // @[Modules.scala 63:156:@7513.4]
  assign _T_60619 = _T_60618[10:0]; // @[Modules.scala 63:156:@7514.4]
  assign buffer_1_782 = $signed(_T_60619); // @[Modules.scala 63:156:@7515.4]
  assign _T_60621 = $signed(buffer_1_782) + $signed(buffer_1_734); // @[Modules.scala 63:156:@7517.4]
  assign _T_60622 = _T_60621[10:0]; // @[Modules.scala 63:156:@7518.4]
  assign buffer_1_783 = $signed(_T_60622); // @[Modules.scala 63:156:@7519.4]
  assign _T_60638 = $signed(io_in_4) - $signed(io_in_5); // @[Modules.scala 40:46:@7536.4]
  assign _T_60639 = _T_60638[4:0]; // @[Modules.scala 40:46:@7537.4]
  assign _T_60640 = $signed(_T_60639); // @[Modules.scala 40:46:@7538.4]
  assign _T_60645 = $signed(_T_54290) - $signed(io_in_7); // @[Modules.scala 46:47:@7543.4]
  assign _T_60646 = _T_60645[4:0]; // @[Modules.scala 46:47:@7544.4]
  assign _T_60647 = $signed(_T_60646); // @[Modules.scala 46:47:@7545.4]
  assign _T_60648 = $signed(io_in_8) - $signed(io_in_9); // @[Modules.scala 40:46:@7547.4]
  assign _T_60649 = _T_60648[4:0]; // @[Modules.scala 40:46:@7548.4]
  assign _T_60650 = $signed(_T_60649); // @[Modules.scala 40:46:@7549.4]
  assign _T_60651 = $signed(io_in_10) + $signed(io_in_11); // @[Modules.scala 37:46:@7551.4]
  assign _T_60652 = _T_60651[4:0]; // @[Modules.scala 37:46:@7552.4]
  assign _T_60653 = $signed(_T_60652); // @[Modules.scala 37:46:@7553.4]
  assign _T_60675 = $signed(_T_54328) + $signed(io_in_19); // @[Modules.scala 43:47:@7576.4]
  assign _T_60676 = _T_60675[4:0]; // @[Modules.scala 43:47:@7577.4]
  assign _T_60677 = $signed(_T_60676); // @[Modules.scala 43:47:@7578.4]
  assign _T_60678 = $signed(io_in_20) - $signed(io_in_21); // @[Modules.scala 40:46:@7580.4]
  assign _T_60679 = _T_60678[4:0]; // @[Modules.scala 40:46:@7581.4]
  assign _T_60680 = $signed(_T_60679); // @[Modules.scala 40:46:@7582.4]
  assign _T_60681 = $signed(io_in_22) + $signed(io_in_23); // @[Modules.scala 37:46:@7584.4]
  assign _T_60682 = _T_60681[4:0]; // @[Modules.scala 37:46:@7585.4]
  assign _T_60683 = $signed(_T_60682); // @[Modules.scala 37:46:@7586.4]
  assign _T_60688 = $signed(_T_54345) - $signed(io_in_25); // @[Modules.scala 46:47:@7591.4]
  assign _T_60689 = _T_60688[4:0]; // @[Modules.scala 46:47:@7592.4]
  assign _T_60690 = $signed(_T_60689); // @[Modules.scala 46:47:@7593.4]
  assign _T_60701 = $signed(io_in_30) - $signed(io_in_31); // @[Modules.scala 40:46:@7606.4]
  assign _T_60702 = _T_60701[4:0]; // @[Modules.scala 40:46:@7607.4]
  assign _T_60703 = $signed(_T_60702); // @[Modules.scala 40:46:@7608.4]
  assign _T_60705 = $signed(5'sh0) - $signed(io_in_32); // @[Modules.scala 46:37:@7610.4]
  assign _T_60706 = _T_60705[4:0]; // @[Modules.scala 46:37:@7611.4]
  assign _T_60707 = $signed(_T_60706); // @[Modules.scala 46:37:@7612.4]
  assign _T_60708 = $signed(_T_60707) - $signed(io_in_33); // @[Modules.scala 46:47:@7613.4]
  assign _T_60709 = _T_60708[4:0]; // @[Modules.scala 46:47:@7614.4]
  assign _T_60710 = $signed(_T_60709); // @[Modules.scala 46:47:@7615.4]
  assign _T_60720 = $signed(io_in_40) - $signed(io_in_41); // @[Modules.scala 40:46:@7629.4]
  assign _T_60721 = _T_60720[4:0]; // @[Modules.scala 40:46:@7630.4]
  assign _T_60722 = $signed(_T_60721); // @[Modules.scala 40:46:@7631.4]
  assign _T_60743 = $signed(5'sh0) - $signed(io_in_52); // @[Modules.scala 46:37:@7656.4]
  assign _T_60744 = _T_60743[4:0]; // @[Modules.scala 46:37:@7657.4]
  assign _T_60745 = $signed(_T_60744); // @[Modules.scala 46:37:@7658.4]
  assign _T_60746 = $signed(_T_60745) - $signed(io_in_53); // @[Modules.scala 46:47:@7659.4]
  assign _T_60747 = _T_60746[4:0]; // @[Modules.scala 46:47:@7660.4]
  assign _T_60748 = $signed(_T_60747); // @[Modules.scala 46:47:@7661.4]
  assign _T_60756 = $signed(io_in_56) + $signed(io_in_57); // @[Modules.scala 37:46:@7670.4]
  assign _T_60757 = _T_60756[4:0]; // @[Modules.scala 37:46:@7671.4]
  assign _T_60758 = $signed(_T_60757); // @[Modules.scala 37:46:@7672.4]
  assign _T_60763 = $signed(_T_54444) + $signed(io_in_59); // @[Modules.scala 43:47:@7677.4]
  assign _T_60764 = _T_60763[4:0]; // @[Modules.scala 43:47:@7678.4]
  assign _T_60765 = $signed(_T_60764); // @[Modules.scala 43:47:@7679.4]
  assign _T_60777 = $signed(_T_54458) + $signed(io_in_63); // @[Modules.scala 43:47:@7691.4]
  assign _T_60778 = _T_60777[4:0]; // @[Modules.scala 43:47:@7692.4]
  assign _T_60779 = $signed(_T_60778); // @[Modules.scala 43:47:@7693.4]
  assign _T_60793 = $signed(_T_54486) + $signed(io_in_71); // @[Modules.scala 43:47:@7710.4]
  assign _T_60794 = _T_60793[4:0]; // @[Modules.scala 43:47:@7711.4]
  assign _T_60795 = $signed(_T_60794); // @[Modules.scala 43:47:@7712.4]
  assign _T_60805 = $signed(io_in_78) - $signed(io_in_79); // @[Modules.scala 40:46:@7726.4]
  assign _T_60806 = _T_60805[4:0]; // @[Modules.scala 40:46:@7727.4]
  assign _T_60807 = $signed(_T_60806); // @[Modules.scala 40:46:@7728.4]
  assign _T_60815 = $signed(io_in_82) + $signed(io_in_83); // @[Modules.scala 37:46:@7737.4]
  assign _T_60816 = _T_60815[4:0]; // @[Modules.scala 37:46:@7738.4]
  assign _T_60817 = $signed(_T_60816); // @[Modules.scala 37:46:@7739.4]
  assign _T_60822 = $signed(_T_57708) - $signed(io_in_85); // @[Modules.scala 46:47:@7744.4]
  assign _T_60823 = _T_60822[4:0]; // @[Modules.scala 46:47:@7745.4]
  assign _T_60824 = $signed(_T_60823); // @[Modules.scala 46:47:@7746.4]
  assign _T_60832 = $signed(io_in_88) - $signed(io_in_89); // @[Modules.scala 40:46:@7755.4]
  assign _T_60833 = _T_60832[4:0]; // @[Modules.scala 40:46:@7756.4]
  assign _T_60834 = $signed(_T_60833); // @[Modules.scala 40:46:@7757.4]
  assign _T_60842 = $signed(5'sh0) - $signed(io_in_94); // @[Modules.scala 46:37:@7767.4]
  assign _T_60843 = _T_60842[4:0]; // @[Modules.scala 46:37:@7768.4]
  assign _T_60844 = $signed(_T_60843); // @[Modules.scala 46:37:@7769.4]
  assign _T_60845 = $signed(_T_60844) - $signed(io_in_95); // @[Modules.scala 46:47:@7770.4]
  assign _T_60846 = _T_60845[4:0]; // @[Modules.scala 46:47:@7771.4]
  assign _T_60847 = $signed(_T_60846); // @[Modules.scala 46:47:@7772.4]
  assign _T_60852 = $signed(_T_54549) - $signed(io_in_97); // @[Modules.scala 46:47:@7777.4]
  assign _T_60853 = _T_60852[4:0]; // @[Modules.scala 46:47:@7778.4]
  assign _T_60854 = $signed(_T_60853); // @[Modules.scala 46:47:@7779.4]
  assign _T_60856 = $signed(5'sh0) - $signed(io_in_98); // @[Modules.scala 46:37:@7781.4]
  assign _T_60857 = _T_60856[4:0]; // @[Modules.scala 46:37:@7782.4]
  assign _T_60858 = $signed(_T_60857); // @[Modules.scala 46:37:@7783.4]
  assign _T_60859 = $signed(_T_60858) - $signed(io_in_99); // @[Modules.scala 46:47:@7784.4]
  assign _T_60860 = _T_60859[4:0]; // @[Modules.scala 46:47:@7785.4]
  assign _T_60861 = $signed(_T_60860); // @[Modules.scala 46:47:@7786.4]
  assign _T_60862 = $signed(io_in_100) - $signed(io_in_101); // @[Modules.scala 40:46:@7788.4]
  assign _T_60863 = _T_60862[4:0]; // @[Modules.scala 40:46:@7789.4]
  assign _T_60864 = $signed(_T_60863); // @[Modules.scala 40:46:@7790.4]
  assign _T_60875 = $signed(5'sh0) - $signed(io_in_108); // @[Modules.scala 46:37:@7804.4]
  assign _T_60876 = _T_60875[4:0]; // @[Modules.scala 46:37:@7805.4]
  assign _T_60877 = $signed(_T_60876); // @[Modules.scala 46:37:@7806.4]
  assign _T_60878 = $signed(_T_60877) - $signed(io_in_109); // @[Modules.scala 46:47:@7807.4]
  assign _T_60879 = _T_60878[4:0]; // @[Modules.scala 46:47:@7808.4]
  assign _T_60880 = $signed(_T_60879); // @[Modules.scala 46:47:@7809.4]
  assign _T_60882 = $signed(5'sh0) - $signed(io_in_110); // @[Modules.scala 46:37:@7811.4]
  assign _T_60883 = _T_60882[4:0]; // @[Modules.scala 46:37:@7812.4]
  assign _T_60884 = $signed(_T_60883); // @[Modules.scala 46:37:@7813.4]
  assign _T_60885 = $signed(_T_60884) - $signed(io_in_111); // @[Modules.scala 46:47:@7814.4]
  assign _T_60886 = _T_60885[4:0]; // @[Modules.scala 46:47:@7815.4]
  assign _T_60887 = $signed(_T_60886); // @[Modules.scala 46:47:@7816.4]
  assign _T_60903 = $signed(5'sh0) - $signed(io_in_116); // @[Modules.scala 46:37:@7832.4]
  assign _T_60904 = _T_60903[4:0]; // @[Modules.scala 46:37:@7833.4]
  assign _T_60905 = $signed(_T_60904); // @[Modules.scala 46:37:@7834.4]
  assign _T_60906 = $signed(_T_60905) - $signed(io_in_117); // @[Modules.scala 46:47:@7835.4]
  assign _T_60907 = _T_60906[4:0]; // @[Modules.scala 46:47:@7836.4]
  assign _T_60908 = $signed(_T_60907); // @[Modules.scala 46:47:@7837.4]
  assign _T_60955 = $signed(_T_54632) - $signed(io_in_131); // @[Modules.scala 46:47:@7884.4]
  assign _T_60956 = _T_60955[4:0]; // @[Modules.scala 46:47:@7885.4]
  assign _T_60957 = $signed(_T_60956); // @[Modules.scala 46:47:@7886.4]
  assign _T_60979 = $signed(5'sh0) - $signed(io_in_140); // @[Modules.scala 43:37:@7910.4]
  assign _T_60980 = _T_60979[4:0]; // @[Modules.scala 43:37:@7911.4]
  assign _T_60981 = $signed(_T_60980); // @[Modules.scala 43:37:@7912.4]
  assign _T_60982 = $signed(_T_60981) + $signed(io_in_141); // @[Modules.scala 43:47:@7913.4]
  assign _T_60983 = _T_60982[4:0]; // @[Modules.scala 43:47:@7914.4]
  assign _T_60984 = $signed(_T_60983); // @[Modules.scala 43:47:@7915.4]
  assign _T_60985 = $signed(io_in_142) - $signed(io_in_143); // @[Modules.scala 40:46:@7917.4]
  assign _T_60986 = _T_60985[4:0]; // @[Modules.scala 40:46:@7918.4]
  assign _T_60987 = $signed(_T_60986); // @[Modules.scala 40:46:@7919.4]
  assign _T_61003 = $signed(5'sh0) - $signed(io_in_148); // @[Modules.scala 46:37:@7935.4]
  assign _T_61004 = _T_61003[4:0]; // @[Modules.scala 46:37:@7936.4]
  assign _T_61005 = $signed(_T_61004); // @[Modules.scala 46:37:@7937.4]
  assign _T_61006 = $signed(_T_61005) - $signed(io_in_149); // @[Modules.scala 46:47:@7938.4]
  assign _T_61007 = _T_61006[4:0]; // @[Modules.scala 46:47:@7939.4]
  assign _T_61008 = $signed(_T_61007); // @[Modules.scala 46:47:@7940.4]
  assign _T_61041 = $signed(_T_54702) + $signed(io_in_159); // @[Modules.scala 43:47:@7973.4]
  assign _T_61042 = _T_61041[4:0]; // @[Modules.scala 43:47:@7974.4]
  assign _T_61043 = $signed(_T_61042); // @[Modules.scala 43:47:@7975.4]
  assign _T_61044 = $signed(io_in_160) + $signed(io_in_161); // @[Modules.scala 37:46:@7977.4]
  assign _T_61045 = _T_61044[4:0]; // @[Modules.scala 37:46:@7978.4]
  assign _T_61046 = $signed(_T_61045); // @[Modules.scala 37:46:@7979.4]
  assign _T_61050 = $signed(io_in_164) + $signed(io_in_165); // @[Modules.scala 37:46:@7985.4]
  assign _T_61051 = _T_61050[4:0]; // @[Modules.scala 37:46:@7986.4]
  assign _T_61052 = $signed(_T_61051); // @[Modules.scala 37:46:@7987.4]
  assign _T_61056 = $signed(io_in_168) - $signed(io_in_169); // @[Modules.scala 40:46:@7993.4]
  assign _T_61057 = _T_61056[4:0]; // @[Modules.scala 40:46:@7994.4]
  assign _T_61058 = $signed(_T_61057); // @[Modules.scala 40:46:@7995.4]
  assign _T_61067 = $signed(5'sh0) - $signed(io_in_172); // @[Modules.scala 46:37:@8004.4]
  assign _T_61068 = _T_61067[4:0]; // @[Modules.scala 46:37:@8005.4]
  assign _T_61069 = $signed(_T_61068); // @[Modules.scala 46:37:@8006.4]
  assign _T_61070 = $signed(_T_61069) - $signed(io_in_173); // @[Modules.scala 46:47:@8007.4]
  assign _T_61071 = _T_61070[4:0]; // @[Modules.scala 46:47:@8008.4]
  assign _T_61072 = $signed(_T_61071); // @[Modules.scala 46:47:@8009.4]
  assign _T_61116 = $signed(5'sh0) - $signed(io_in_186); // @[Modules.scala 46:37:@8053.4]
  assign _T_61117 = _T_61116[4:0]; // @[Modules.scala 46:37:@8054.4]
  assign _T_61118 = $signed(_T_61117); // @[Modules.scala 46:37:@8055.4]
  assign _T_61119 = $signed(_T_61118) - $signed(io_in_187); // @[Modules.scala 46:47:@8056.4]
  assign _T_61120 = _T_61119[4:0]; // @[Modules.scala 46:47:@8057.4]
  assign _T_61121 = $signed(_T_61120); // @[Modules.scala 46:47:@8058.4]
  assign _T_61129 = $signed(io_in_190) + $signed(io_in_191); // @[Modules.scala 37:46:@8067.4]
  assign _T_61130 = _T_61129[4:0]; // @[Modules.scala 37:46:@8068.4]
  assign _T_61131 = $signed(_T_61130); // @[Modules.scala 37:46:@8069.4]
  assign _T_61132 = $signed(io_in_192) + $signed(io_in_193); // @[Modules.scala 37:46:@8071.4]
  assign _T_61133 = _T_61132[4:0]; // @[Modules.scala 37:46:@8072.4]
  assign _T_61134 = $signed(_T_61133); // @[Modules.scala 37:46:@8073.4]
  assign _T_61135 = $signed(io_in_194) + $signed(io_in_195); // @[Modules.scala 37:46:@8075.4]
  assign _T_61136 = _T_61135[4:0]; // @[Modules.scala 37:46:@8076.4]
  assign _T_61137 = $signed(_T_61136); // @[Modules.scala 37:46:@8077.4]
  assign _T_61145 = $signed(_T_57983) - $signed(io_in_199); // @[Modules.scala 46:47:@8086.4]
  assign _T_61146 = _T_61145[4:0]; // @[Modules.scala 46:47:@8087.4]
  assign _T_61147 = $signed(_T_61146); // @[Modules.scala 46:47:@8088.4]
  assign _T_61173 = $signed(_T_54842) - $signed(io_in_207); // @[Modules.scala 46:47:@8114.4]
  assign _T_61174 = _T_61173[4:0]; // @[Modules.scala 46:47:@8115.4]
  assign _T_61175 = $signed(_T_61174); // @[Modules.scala 46:47:@8116.4]
  assign _T_61180 = $signed(_T_54849) - $signed(io_in_209); // @[Modules.scala 46:47:@8121.4]
  assign _T_61181 = _T_61180[4:0]; // @[Modules.scala 46:47:@8122.4]
  assign _T_61182 = $signed(_T_61181); // @[Modules.scala 46:47:@8123.4]
  assign _T_61189 = $signed(io_in_214) + $signed(io_in_215); // @[Modules.scala 37:46:@8133.4]
  assign _T_61190 = _T_61189[4:0]; // @[Modules.scala 37:46:@8134.4]
  assign _T_61191 = $signed(_T_61190); // @[Modules.scala 37:46:@8135.4]
  assign _T_61199 = $signed(io_in_218) + $signed(io_in_219); // @[Modules.scala 37:46:@8144.4]
  assign _T_61200 = _T_61199[4:0]; // @[Modules.scala 37:46:@8145.4]
  assign _T_61201 = $signed(_T_61200); // @[Modules.scala 37:46:@8146.4]
  assign _T_61205 = $signed(io_in_222) + $signed(io_in_223); // @[Modules.scala 37:46:@8152.4]
  assign _T_61206 = _T_61205[4:0]; // @[Modules.scala 37:46:@8153.4]
  assign _T_61207 = $signed(_T_61206); // @[Modules.scala 37:46:@8154.4]
  assign _T_61247 = $signed(_T_54932) + $signed(io_in_235); // @[Modules.scala 43:47:@8194.4]
  assign _T_61248 = _T_61247[4:0]; // @[Modules.scala 43:47:@8195.4]
  assign _T_61249 = $signed(_T_61248); // @[Modules.scala 43:47:@8196.4]
  assign _T_61330 = $signed(_T_55023) + $signed(io_in_261); // @[Modules.scala 43:47:@8279.4]
  assign _T_61331 = _T_61330[4:0]; // @[Modules.scala 43:47:@8280.4]
  assign _T_61332 = $signed(_T_61331); // @[Modules.scala 43:47:@8281.4]
  assign _T_61337 = $signed(_T_58167) + $signed(io_in_263); // @[Modules.scala 43:47:@8286.4]
  assign _T_61338 = _T_61337[4:0]; // @[Modules.scala 43:47:@8287.4]
  assign _T_61339 = $signed(_T_61338); // @[Modules.scala 43:47:@8288.4]
  assign _T_61413 = $signed(_T_55110) + $signed(io_in_287); // @[Modules.scala 43:47:@8364.4]
  assign _T_61414 = _T_61413[4:0]; // @[Modules.scala 43:47:@8365.4]
  assign _T_61415 = $signed(_T_61414); // @[Modules.scala 43:47:@8366.4]
  assign _T_61416 = $signed(io_in_288) + $signed(io_in_289); // @[Modules.scala 37:46:@8368.4]
  assign _T_61417 = _T_61416[4:0]; // @[Modules.scala 37:46:@8369.4]
  assign _T_61418 = $signed(_T_61417); // @[Modules.scala 37:46:@8370.4]
  assign _T_61419 = $signed(io_in_290) + $signed(io_in_291); // @[Modules.scala 37:46:@8372.4]
  assign _T_61420 = _T_61419[4:0]; // @[Modules.scala 37:46:@8373.4]
  assign _T_61421 = $signed(_T_61420); // @[Modules.scala 37:46:@8374.4]
  assign _T_61468 = $signed(_T_55173) + $signed(io_in_305); // @[Modules.scala 43:47:@8421.4]
  assign _T_61469 = _T_61468[4:0]; // @[Modules.scala 43:47:@8422.4]
  assign _T_61470 = $signed(_T_61469); // @[Modules.scala 43:47:@8423.4]
  assign _T_61495 = $signed(io_in_314) + $signed(io_in_315); // @[Modules.scala 37:46:@8450.4]
  assign _T_61496 = _T_61495[4:0]; // @[Modules.scala 37:46:@8451.4]
  assign _T_61497 = $signed(_T_61496); // @[Modules.scala 37:46:@8452.4]
  assign _T_61504 = $signed(io_in_320) - $signed(io_in_321); // @[Modules.scala 40:46:@8462.4]
  assign _T_61505 = _T_61504[4:0]; // @[Modules.scala 40:46:@8463.4]
  assign _T_61506 = $signed(_T_61505); // @[Modules.scala 40:46:@8464.4]
  assign _T_61542 = $signed(_T_55259) + $signed(io_in_333); // @[Modules.scala 43:47:@8501.4]
  assign _T_61543 = _T_61542[4:0]; // @[Modules.scala 43:47:@8502.4]
  assign _T_61544 = $signed(_T_61543); // @[Modules.scala 43:47:@8503.4]
  assign _T_61587 = $signed(io_in_354) - $signed(io_in_355); // @[Modules.scala 40:46:@8554.4]
  assign _T_61588 = _T_61587[4:0]; // @[Modules.scala 40:46:@8555.4]
  assign _T_61589 = $signed(_T_61588); // @[Modules.scala 40:46:@8556.4]
  assign _T_61601 = $signed(_T_58431) - $signed(io_in_359); // @[Modules.scala 46:47:@8568.4]
  assign _T_61602 = _T_61601[4:0]; // @[Modules.scala 46:47:@8569.4]
  assign _T_61603 = $signed(_T_61602); // @[Modules.scala 46:47:@8570.4]
  assign _T_61608 = $signed(_T_55317) + $signed(io_in_361); // @[Modules.scala 43:47:@8575.4]
  assign _T_61609 = _T_61608[4:0]; // @[Modules.scala 43:47:@8576.4]
  assign _T_61610 = $signed(_T_61609); // @[Modules.scala 43:47:@8577.4]
  assign _T_61611 = $signed(io_in_362) - $signed(io_in_363); // @[Modules.scala 40:46:@8579.4]
  assign _T_61612 = _T_61611[4:0]; // @[Modules.scala 40:46:@8580.4]
  assign _T_61613 = $signed(_T_61612); // @[Modules.scala 40:46:@8581.4]
  assign _T_61656 = $signed(io_in_384) + $signed(io_in_385); // @[Modules.scala 37:46:@8632.4]
  assign _T_61657 = _T_61656[4:0]; // @[Modules.scala 37:46:@8633.4]
  assign _T_61658 = $signed(_T_61657); // @[Modules.scala 37:46:@8634.4]
  assign _T_61660 = $signed(5'sh0) - $signed(io_in_386); // @[Modules.scala 46:37:@8636.4]
  assign _T_61661 = _T_61660[4:0]; // @[Modules.scala 46:37:@8637.4]
  assign _T_61662 = $signed(_T_61661); // @[Modules.scala 46:37:@8638.4]
  assign _T_61663 = $signed(_T_61662) - $signed(io_in_387); // @[Modules.scala 46:47:@8639.4]
  assign _T_61664 = _T_61663[4:0]; // @[Modules.scala 46:47:@8640.4]
  assign _T_61665 = $signed(_T_61664); // @[Modules.scala 46:47:@8641.4]
  assign _T_61667 = $signed(5'sh0) - $signed(io_in_388); // @[Modules.scala 46:37:@8643.4]
  assign _T_61668 = _T_61667[4:0]; // @[Modules.scala 46:37:@8644.4]
  assign _T_61669 = $signed(_T_61668); // @[Modules.scala 46:37:@8645.4]
  assign _T_61670 = $signed(_T_61669) - $signed(io_in_389); // @[Modules.scala 46:47:@8646.4]
  assign _T_61671 = _T_61670[4:0]; // @[Modules.scala 46:47:@8647.4]
  assign _T_61672 = $signed(_T_61671); // @[Modules.scala 46:47:@8648.4]
  assign _T_61715 = $signed(_T_58561) + $signed(io_in_411); // @[Modules.scala 43:47:@8699.4]
  assign _T_61716 = _T_61715[4:0]; // @[Modules.scala 43:47:@8700.4]
  assign _T_61717 = $signed(_T_61716); // @[Modules.scala 43:47:@8701.4]
  assign _T_61725 = $signed(5'sh0) - $signed(io_in_416); // @[Modules.scala 46:37:@8711.4]
  assign _T_61726 = _T_61725[4:0]; // @[Modules.scala 46:37:@8712.4]
  assign _T_61727 = $signed(_T_61726); // @[Modules.scala 46:37:@8713.4]
  assign _T_61728 = $signed(_T_61727) - $signed(io_in_417); // @[Modules.scala 46:47:@8714.4]
  assign _T_61729 = _T_61728[4:0]; // @[Modules.scala 46:47:@8715.4]
  assign _T_61730 = $signed(_T_61729); // @[Modules.scala 46:47:@8716.4]
  assign _T_61745 = $signed(io_in_422) + $signed(io_in_423); // @[Modules.scala 37:46:@8732.4]
  assign _T_61746 = _T_61745[4:0]; // @[Modules.scala 37:46:@8733.4]
  assign _T_61747 = $signed(_T_61746); // @[Modules.scala 37:46:@8734.4]
  assign _T_61752 = $signed(_T_55457) - $signed(io_in_425); // @[Modules.scala 46:47:@8739.4]
  assign _T_61753 = _T_61752[4:0]; // @[Modules.scala 46:47:@8740.4]
  assign _T_61754 = $signed(_T_61753); // @[Modules.scala 46:47:@8741.4]
  assign _T_61762 = $signed(5'sh0) - $signed(io_in_430); // @[Modules.scala 46:37:@8751.4]
  assign _T_61763 = _T_61762[4:0]; // @[Modules.scala 46:37:@8752.4]
  assign _T_61764 = $signed(_T_61763); // @[Modules.scala 46:37:@8753.4]
  assign _T_61765 = $signed(_T_61764) - $signed(io_in_431); // @[Modules.scala 46:47:@8754.4]
  assign _T_61766 = _T_61765[4:0]; // @[Modules.scala 46:47:@8755.4]
  assign _T_61767 = $signed(_T_61766); // @[Modules.scala 46:47:@8756.4]
  assign _T_61785 = $signed(_T_58635) - $signed(io_in_439); // @[Modules.scala 46:47:@8776.4]
  assign _T_61786 = _T_61785[4:0]; // @[Modules.scala 46:47:@8777.4]
  assign _T_61787 = $signed(_T_61786); // @[Modules.scala 46:47:@8778.4]
  assign _T_61789 = $signed(5'sh0) - $signed(io_in_440); // @[Modules.scala 46:37:@8780.4]
  assign _T_61790 = _T_61789[4:0]; // @[Modules.scala 46:37:@8781.4]
  assign _T_61791 = $signed(_T_61790); // @[Modules.scala 46:37:@8782.4]
  assign _T_61792 = $signed(_T_61791) - $signed(io_in_441); // @[Modules.scala 46:47:@8783.4]
  assign _T_61793 = _T_61792[4:0]; // @[Modules.scala 46:47:@8784.4]
  assign _T_61794 = $signed(_T_61793); // @[Modules.scala 46:47:@8785.4]
  assign _T_61837 = $signed(_T_58675) + $signed(io_in_455); // @[Modules.scala 43:47:@8829.4]
  assign _T_61838 = _T_61837[4:0]; // @[Modules.scala 43:47:@8830.4]
  assign _T_61839 = $signed(_T_61838); // @[Modules.scala 43:47:@8831.4]
  assign _T_61840 = $signed(io_in_456) - $signed(io_in_457); // @[Modules.scala 40:46:@8833.4]
  assign _T_61841 = _T_61840[4:0]; // @[Modules.scala 40:46:@8834.4]
  assign _T_61842 = $signed(_T_61841); // @[Modules.scala 40:46:@8835.4]
  assign _T_61844 = $signed(5'sh0) - $signed(io_in_458); // @[Modules.scala 46:37:@8837.4]
  assign _T_61845 = _T_61844[4:0]; // @[Modules.scala 46:37:@8838.4]
  assign _T_61846 = $signed(_T_61845); // @[Modules.scala 46:37:@8839.4]
  assign _T_61847 = $signed(_T_61846) - $signed(io_in_459); // @[Modules.scala 46:47:@8840.4]
  assign _T_61848 = _T_61847[4:0]; // @[Modules.scala 46:47:@8841.4]
  assign _T_61849 = $signed(_T_61848); // @[Modules.scala 46:47:@8842.4]
  assign _T_61850 = $signed(io_in_460) + $signed(io_in_461); // @[Modules.scala 37:46:@8844.4]
  assign _T_61851 = _T_61850[4:0]; // @[Modules.scala 37:46:@8845.4]
  assign _T_61852 = $signed(_T_61851); // @[Modules.scala 37:46:@8846.4]
  assign _T_61860 = $signed(_T_58706) + $signed(io_in_465); // @[Modules.scala 43:47:@8855.4]
  assign _T_61861 = _T_61860[4:0]; // @[Modules.scala 43:47:@8856.4]
  assign _T_61862 = $signed(_T_61861); // @[Modules.scala 43:47:@8857.4]
  assign _T_61867 = $signed(5'sh0) - $signed(io_in_468); // @[Modules.scala 46:37:@8863.4]
  assign _T_61868 = _T_61867[4:0]; // @[Modules.scala 46:37:@8864.4]
  assign _T_61869 = $signed(_T_61868); // @[Modules.scala 46:37:@8865.4]
  assign _T_61870 = $signed(_T_61869) - $signed(io_in_469); // @[Modules.scala 46:47:@8866.4]
  assign _T_61871 = _T_61870[4:0]; // @[Modules.scala 46:47:@8867.4]
  assign _T_61872 = $signed(_T_61871); // @[Modules.scala 46:47:@8868.4]
  assign _T_61890 = $signed(io_in_476) + $signed(io_in_477); // @[Modules.scala 37:46:@8888.4]
  assign _T_61891 = _T_61890[4:0]; // @[Modules.scala 37:46:@8889.4]
  assign _T_61892 = $signed(_T_61891); // @[Modules.scala 37:46:@8890.4]
  assign _T_61904 = $signed(5'sh0) - $signed(io_in_482); // @[Modules.scala 46:37:@8903.4]
  assign _T_61905 = _T_61904[4:0]; // @[Modules.scala 46:37:@8904.4]
  assign _T_61906 = $signed(_T_61905); // @[Modules.scala 46:37:@8905.4]
  assign _T_61907 = $signed(_T_61906) - $signed(io_in_483); // @[Modules.scala 46:47:@8906.4]
  assign _T_61908 = _T_61907[4:0]; // @[Modules.scala 46:47:@8907.4]
  assign _T_61909 = $signed(_T_61908); // @[Modules.scala 46:47:@8908.4]
  assign _T_61914 = $signed(_T_58756) + $signed(io_in_485); // @[Modules.scala 43:47:@8913.4]
  assign _T_61915 = _T_61914[4:0]; // @[Modules.scala 43:47:@8914.4]
  assign _T_61916 = $signed(_T_61915); // @[Modules.scala 43:47:@8915.4]
  assign _T_61920 = $signed(io_in_488) + $signed(io_in_489); // @[Modules.scala 37:46:@8921.4]
  assign _T_61921 = _T_61920[4:0]; // @[Modules.scala 37:46:@8922.4]
  assign _T_61922 = $signed(_T_61921); // @[Modules.scala 37:46:@8923.4]
  assign _T_61940 = $signed(5'sh0) - $signed(io_in_498); // @[Modules.scala 46:37:@8944.4]
  assign _T_61941 = _T_61940[4:0]; // @[Modules.scala 46:37:@8945.4]
  assign _T_61942 = $signed(_T_61941); // @[Modules.scala 46:37:@8946.4]
  assign _T_61943 = $signed(_T_61942) - $signed(io_in_499); // @[Modules.scala 46:47:@8947.4]
  assign _T_61944 = _T_61943[4:0]; // @[Modules.scala 46:47:@8948.4]
  assign _T_61945 = $signed(_T_61944); // @[Modules.scala 46:47:@8949.4]
  assign _T_61971 = $signed(_T_55644) - $signed(io_in_507); // @[Modules.scala 46:47:@8975.4]
  assign _T_61972 = _T_61971[4:0]; // @[Modules.scala 46:47:@8976.4]
  assign _T_61973 = $signed(_T_61972); // @[Modules.scala 46:47:@8977.4]
  assign _T_61998 = $signed(io_in_516) + $signed(io_in_517); // @[Modules.scala 37:46:@9004.4]
  assign _T_61999 = _T_61998[4:0]; // @[Modules.scala 37:46:@9005.4]
  assign _T_62000 = $signed(_T_61999); // @[Modules.scala 37:46:@9006.4]
  assign _T_62001 = $signed(io_in_518) - $signed(io_in_519); // @[Modules.scala 40:46:@9008.4]
  assign _T_62002 = _T_62001[4:0]; // @[Modules.scala 40:46:@9009.4]
  assign _T_62003 = $signed(_T_62002); // @[Modules.scala 40:46:@9010.4]
  assign _T_62008 = $signed(_T_55677) - $signed(io_in_521); // @[Modules.scala 46:47:@9015.4]
  assign _T_62009 = _T_62008[4:0]; // @[Modules.scala 46:47:@9016.4]
  assign _T_62010 = $signed(_T_62009); // @[Modules.scala 46:47:@9017.4]
  assign _T_62022 = $signed(_T_55691) - $signed(io_in_525); // @[Modules.scala 46:47:@9029.4]
  assign _T_62023 = _T_62022[4:0]; // @[Modules.scala 46:47:@9030.4]
  assign _T_62024 = $signed(_T_62023); // @[Modules.scala 46:47:@9031.4]
  assign _T_62026 = $signed(5'sh0) - $signed(io_in_526); // @[Modules.scala 46:37:@9033.4]
  assign _T_62027 = _T_62026[4:0]; // @[Modules.scala 46:37:@9034.4]
  assign _T_62028 = $signed(_T_62027); // @[Modules.scala 46:37:@9035.4]
  assign _T_62029 = $signed(_T_62028) - $signed(io_in_527); // @[Modules.scala 46:47:@9036.4]
  assign _T_62030 = _T_62029[4:0]; // @[Modules.scala 46:47:@9037.4]
  assign _T_62031 = $signed(_T_62030); // @[Modules.scala 46:47:@9038.4]
  assign _T_62047 = $signed(5'sh0) - $signed(io_in_532); // @[Modules.scala 46:37:@9054.4]
  assign _T_62048 = _T_62047[4:0]; // @[Modules.scala 46:37:@9055.4]
  assign _T_62049 = $signed(_T_62048); // @[Modules.scala 46:37:@9056.4]
  assign _T_62050 = $signed(_T_62049) - $signed(io_in_533); // @[Modules.scala 46:47:@9057.4]
  assign _T_62051 = _T_62050[4:0]; // @[Modules.scala 46:47:@9058.4]
  assign _T_62052 = $signed(_T_62051); // @[Modules.scala 46:47:@9059.4]
  assign _T_62057 = $signed(_T_55714) - $signed(io_in_535); // @[Modules.scala 46:47:@9064.4]
  assign _T_62058 = _T_62057[4:0]; // @[Modules.scala 46:47:@9065.4]
  assign _T_62059 = $signed(_T_62058); // @[Modules.scala 46:47:@9066.4]
  assign _T_62092 = $signed(_T_55749) + $signed(io_in_545); // @[Modules.scala 43:47:@9099.4]
  assign _T_62093 = _T_62092[4:0]; // @[Modules.scala 43:47:@9100.4]
  assign _T_62094 = $signed(_T_62093); // @[Modules.scala 43:47:@9101.4]
  assign _T_62106 = $signed(_T_55763) + $signed(io_in_549); // @[Modules.scala 43:47:@9113.4]
  assign _T_62107 = _T_62106[4:0]; // @[Modules.scala 43:47:@9114.4]
  assign _T_62108 = $signed(_T_62107); // @[Modules.scala 43:47:@9115.4]
  assign _T_62110 = $signed(5'sh0) - $signed(io_in_550); // @[Modules.scala 43:37:@9117.4]
  assign _T_62111 = _T_62110[4:0]; // @[Modules.scala 43:37:@9118.4]
  assign _T_62112 = $signed(_T_62111); // @[Modules.scala 43:37:@9119.4]
  assign _T_62113 = $signed(_T_62112) + $signed(io_in_551); // @[Modules.scala 43:47:@9120.4]
  assign _T_62114 = _T_62113[4:0]; // @[Modules.scala 43:47:@9121.4]
  assign _T_62115 = $signed(_T_62114); // @[Modules.scala 43:47:@9122.4]
  assign _T_62116 = $signed(io_in_552) + $signed(io_in_553); // @[Modules.scala 37:46:@9124.4]
  assign _T_62117 = _T_62116[4:0]; // @[Modules.scala 37:46:@9125.4]
  assign _T_62118 = $signed(_T_62117); // @[Modules.scala 37:46:@9126.4]
  assign _T_62140 = $signed(io_in_560) - $signed(io_in_561); // @[Modules.scala 40:46:@9149.4]
  assign _T_62141 = _T_62140[4:0]; // @[Modules.scala 40:46:@9150.4]
  assign _T_62142 = $signed(_T_62141); // @[Modules.scala 40:46:@9151.4]
  assign _T_62182 = $signed(_T_55835) - $signed(io_in_573); // @[Modules.scala 46:47:@9191.4]
  assign _T_62183 = _T_62182[4:0]; // @[Modules.scala 46:47:@9192.4]
  assign _T_62184 = $signed(_T_62183); // @[Modules.scala 46:47:@9193.4]
  assign _T_62195 = $signed(5'sh0) - $signed(io_in_580); // @[Modules.scala 46:37:@9207.4]
  assign _T_62196 = _T_62195[4:0]; // @[Modules.scala 46:37:@9208.4]
  assign _T_62197 = $signed(_T_62196); // @[Modules.scala 46:37:@9209.4]
  assign _T_62198 = $signed(_T_62197) - $signed(io_in_581); // @[Modules.scala 46:47:@9210.4]
  assign _T_62199 = _T_62198[4:0]; // @[Modules.scala 46:47:@9211.4]
  assign _T_62200 = $signed(_T_62199); // @[Modules.scala 46:47:@9212.4]
  assign _T_62222 = $signed(io_in_588) - $signed(io_in_589); // @[Modules.scala 40:46:@9235.4]
  assign _T_62223 = _T_62222[4:0]; // @[Modules.scala 40:46:@9236.4]
  assign _T_62224 = $signed(_T_62223); // @[Modules.scala 40:46:@9237.4]
  assign _T_62225 = $signed(io_in_590) - $signed(io_in_591); // @[Modules.scala 40:46:@9239.4]
  assign _T_62226 = _T_62225[4:0]; // @[Modules.scala 40:46:@9240.4]
  assign _T_62227 = $signed(_T_62226); // @[Modules.scala 40:46:@9241.4]
  assign _T_62239 = $signed(_T_55896) + $signed(io_in_595); // @[Modules.scala 43:47:@9253.4]
  assign _T_62240 = _T_62239[4:0]; // @[Modules.scala 43:47:@9254.4]
  assign _T_62241 = $signed(_T_62240); // @[Modules.scala 43:47:@9255.4]
  assign _T_62242 = $signed(io_in_596) + $signed(io_in_597); // @[Modules.scala 37:46:@9257.4]
  assign _T_62243 = _T_62242[4:0]; // @[Modules.scala 37:46:@9258.4]
  assign _T_62244 = $signed(_T_62243); // @[Modules.scala 37:46:@9259.4]
  assign _T_62245 = $signed(io_in_598) - $signed(io_in_599); // @[Modules.scala 40:46:@9261.4]
  assign _T_62246 = _T_62245[4:0]; // @[Modules.scala 40:46:@9262.4]
  assign _T_62247 = $signed(_T_62246); // @[Modules.scala 40:46:@9263.4]
  assign _T_62249 = $signed(5'sh0) - $signed(io_in_600); // @[Modules.scala 43:37:@9265.4]
  assign _T_62250 = _T_62249[4:0]; // @[Modules.scala 43:37:@9266.4]
  assign _T_62251 = $signed(_T_62250); // @[Modules.scala 43:37:@9267.4]
  assign _T_62252 = $signed(_T_62251) + $signed(io_in_601); // @[Modules.scala 43:47:@9268.4]
  assign _T_62253 = _T_62252[4:0]; // @[Modules.scala 43:47:@9269.4]
  assign _T_62254 = $signed(_T_62253); // @[Modules.scala 43:47:@9270.4]
  assign _T_62259 = $signed(5'sh0) - $signed(io_in_604); // @[Modules.scala 43:37:@9276.4]
  assign _T_62260 = _T_62259[4:0]; // @[Modules.scala 43:37:@9277.4]
  assign _T_62261 = $signed(_T_62260); // @[Modules.scala 43:37:@9278.4]
  assign _T_62262 = $signed(_T_62261) + $signed(io_in_605); // @[Modules.scala 43:47:@9279.4]
  assign _T_62263 = _T_62262[4:0]; // @[Modules.scala 43:47:@9280.4]
  assign _T_62264 = $signed(_T_62263); // @[Modules.scala 43:47:@9281.4]
  assign _T_62266 = $signed(5'sh0) - $signed(io_in_606); // @[Modules.scala 46:37:@9283.4]
  assign _T_62267 = _T_62266[4:0]; // @[Modules.scala 46:37:@9284.4]
  assign _T_62268 = $signed(_T_62267); // @[Modules.scala 46:37:@9285.4]
  assign _T_62269 = $signed(_T_62268) - $signed(io_in_607); // @[Modules.scala 46:47:@9286.4]
  assign _T_62270 = _T_62269[4:0]; // @[Modules.scala 46:47:@9287.4]
  assign _T_62271 = $signed(_T_62270); // @[Modules.scala 46:47:@9288.4]
  assign _T_62272 = $signed(io_in_608) + $signed(io_in_609); // @[Modules.scala 37:46:@9290.4]
  assign _T_62273 = _T_62272[4:0]; // @[Modules.scala 37:46:@9291.4]
  assign _T_62274 = $signed(_T_62273); // @[Modules.scala 37:46:@9292.4]
  assign _T_62275 = $signed(io_in_610) - $signed(io_in_611); // @[Modules.scala 40:46:@9294.4]
  assign _T_62276 = _T_62275[4:0]; // @[Modules.scala 40:46:@9295.4]
  assign _T_62277 = $signed(_T_62276); // @[Modules.scala 40:46:@9296.4]
  assign _T_62292 = $signed(io_in_616) + $signed(io_in_617); // @[Modules.scala 37:46:@9312.4]
  assign _T_62293 = _T_62292[4:0]; // @[Modules.scala 37:46:@9313.4]
  assign _T_62294 = $signed(_T_62293); // @[Modules.scala 37:46:@9314.4]
  assign _T_62296 = $signed(5'sh0) - $signed(io_in_618); // @[Modules.scala 46:37:@9316.4]
  assign _T_62297 = _T_62296[4:0]; // @[Modules.scala 46:37:@9317.4]
  assign _T_62298 = $signed(_T_62297); // @[Modules.scala 46:37:@9318.4]
  assign _T_62299 = $signed(_T_62298) - $signed(io_in_619); // @[Modules.scala 46:47:@9319.4]
  assign _T_62300 = _T_62299[4:0]; // @[Modules.scala 46:47:@9320.4]
  assign _T_62301 = $signed(_T_62300); // @[Modules.scala 46:47:@9321.4]
  assign _T_62316 = $signed(io_in_624) - $signed(io_in_625); // @[Modules.scala 40:46:@9337.4]
  assign _T_62317 = _T_62316[4:0]; // @[Modules.scala 40:46:@9338.4]
  assign _T_62318 = $signed(_T_62317); // @[Modules.scala 40:46:@9339.4]
  assign _T_62343 = $signed(io_in_634) + $signed(io_in_635); // @[Modules.scala 37:46:@9366.4]
  assign _T_62344 = _T_62343[4:0]; // @[Modules.scala 37:46:@9367.4]
  assign _T_62345 = $signed(_T_62344); // @[Modules.scala 37:46:@9368.4]
  assign _T_62362 = $signed(io_in_644) - $signed(io_in_645); // @[Modules.scala 40:46:@9389.4]
  assign _T_62363 = _T_62362[4:0]; // @[Modules.scala 40:46:@9390.4]
  assign _T_62364 = $signed(_T_62363); // @[Modules.scala 40:46:@9391.4]
  assign _T_62365 = $signed(io_in_646) - $signed(io_in_647); // @[Modules.scala 40:46:@9393.4]
  assign _T_62366 = _T_62365[4:0]; // @[Modules.scala 40:46:@9394.4]
  assign _T_62367 = $signed(_T_62366); // @[Modules.scala 40:46:@9395.4]
  assign _T_62372 = $signed(_T_56053) + $signed(io_in_649); // @[Modules.scala 43:47:@9400.4]
  assign _T_62373 = _T_62372[4:0]; // @[Modules.scala 43:47:@9401.4]
  assign _T_62374 = $signed(_T_62373); // @[Modules.scala 43:47:@9402.4]
  assign _T_62375 = $signed(io_in_650) - $signed(io_in_651); // @[Modules.scala 40:46:@9404.4]
  assign _T_62376 = _T_62375[4:0]; // @[Modules.scala 40:46:@9405.4]
  assign _T_62377 = $signed(_T_62376); // @[Modules.scala 40:46:@9406.4]
  assign _T_62388 = $signed(io_in_656) - $signed(io_in_657); // @[Modules.scala 40:46:@9419.4]
  assign _T_62389 = _T_62388[4:0]; // @[Modules.scala 40:46:@9420.4]
  assign _T_62390 = $signed(_T_62389); // @[Modules.scala 40:46:@9421.4]
  assign _T_62394 = $signed(io_in_660) + $signed(io_in_661); // @[Modules.scala 37:46:@9427.4]
  assign _T_62395 = _T_62394[4:0]; // @[Modules.scala 37:46:@9428.4]
  assign _T_62396 = $signed(_T_62395); // @[Modules.scala 37:46:@9429.4]
  assign _T_62413 = $signed(io_in_670) + $signed(io_in_671); // @[Modules.scala 37:46:@9450.4]
  assign _T_62414 = _T_62413[4:0]; // @[Modules.scala 37:46:@9451.4]
  assign _T_62415 = $signed(_T_62414); // @[Modules.scala 37:46:@9452.4]
  assign _T_62427 = $signed(5'sh0) - $signed(io_in_676); // @[Modules.scala 46:37:@9465.4]
  assign _T_62428 = _T_62427[4:0]; // @[Modules.scala 46:37:@9466.4]
  assign _T_62429 = $signed(_T_62428); // @[Modules.scala 46:37:@9467.4]
  assign _T_62430 = $signed(_T_62429) - $signed(io_in_677); // @[Modules.scala 46:47:@9468.4]
  assign _T_62431 = _T_62430[4:0]; // @[Modules.scala 46:47:@9469.4]
  assign _T_62432 = $signed(_T_62431); // @[Modules.scala 46:47:@9470.4]
  assign _T_62434 = $signed(5'sh0) - $signed(io_in_678); // @[Modules.scala 46:37:@9472.4]
  assign _T_62435 = _T_62434[4:0]; // @[Modules.scala 46:37:@9473.4]
  assign _T_62436 = $signed(_T_62435); // @[Modules.scala 46:37:@9474.4]
  assign _T_62437 = $signed(_T_62436) - $signed(io_in_679); // @[Modules.scala 46:47:@9475.4]
  assign _T_62438 = _T_62437[4:0]; // @[Modules.scala 46:47:@9476.4]
  assign _T_62439 = $signed(_T_62438); // @[Modules.scala 46:47:@9477.4]
  assign _T_62444 = $signed(_T_59186) - $signed(io_in_681); // @[Modules.scala 46:47:@9482.4]
  assign _T_62445 = _T_62444[4:0]; // @[Modules.scala 46:47:@9483.4]
  assign _T_62446 = $signed(_T_62445); // @[Modules.scala 46:47:@9484.4]
  assign _T_62448 = $signed(5'sh0) - $signed(io_in_682); // @[Modules.scala 46:37:@9486.4]
  assign _T_62449 = _T_62448[4:0]; // @[Modules.scala 46:37:@9487.4]
  assign _T_62450 = $signed(_T_62449); // @[Modules.scala 46:37:@9488.4]
  assign _T_62451 = $signed(_T_62450) - $signed(io_in_683); // @[Modules.scala 46:47:@9489.4]
  assign _T_62452 = _T_62451[4:0]; // @[Modules.scala 46:47:@9490.4]
  assign _T_62453 = $signed(_T_62452); // @[Modules.scala 46:47:@9491.4]
  assign _T_62454 = $signed(io_in_684) - $signed(io_in_685); // @[Modules.scala 40:46:@9493.4]
  assign _T_62455 = _T_62454[4:0]; // @[Modules.scala 40:46:@9494.4]
  assign _T_62456 = $signed(_T_62455); // @[Modules.scala 40:46:@9495.4]
  assign _T_62465 = $signed(5'sh0) - $signed(io_in_688); // @[Modules.scala 43:37:@9504.4]
  assign _T_62466 = _T_62465[4:0]; // @[Modules.scala 43:37:@9505.4]
  assign _T_62467 = $signed(_T_62466); // @[Modules.scala 43:37:@9506.4]
  assign _T_62468 = $signed(_T_62467) + $signed(io_in_689); // @[Modules.scala 43:47:@9507.4]
  assign _T_62469 = _T_62468[4:0]; // @[Modules.scala 43:47:@9508.4]
  assign _T_62470 = $signed(_T_62469); // @[Modules.scala 43:47:@9509.4]
  assign _T_62481 = $signed(5'sh0) - $signed(io_in_696); // @[Modules.scala 46:37:@9523.4]
  assign _T_62482 = _T_62481[4:0]; // @[Modules.scala 46:37:@9524.4]
  assign _T_62483 = $signed(_T_62482); // @[Modules.scala 46:37:@9525.4]
  assign _T_62484 = $signed(_T_62483) - $signed(io_in_697); // @[Modules.scala 46:47:@9526.4]
  assign _T_62485 = _T_62484[4:0]; // @[Modules.scala 46:47:@9527.4]
  assign _T_62486 = $signed(_T_62485); // @[Modules.scala 46:47:@9528.4]
  assign _T_62498 = $signed(_T_56183) - $signed(io_in_701); // @[Modules.scala 46:47:@9540.4]
  assign _T_62499 = _T_62498[4:0]; // @[Modules.scala 46:47:@9541.4]
  assign _T_62500 = $signed(_T_62499); // @[Modules.scala 46:47:@9542.4]
  assign _T_62505 = $signed(5'sh0) - $signed(io_in_704); // @[Modules.scala 46:37:@9548.4]
  assign _T_62506 = _T_62505[4:0]; // @[Modules.scala 46:37:@9549.4]
  assign _T_62507 = $signed(_T_62506); // @[Modules.scala 46:37:@9550.4]
  assign _T_62508 = $signed(_T_62507) - $signed(io_in_705); // @[Modules.scala 46:47:@9551.4]
  assign _T_62509 = _T_62508[4:0]; // @[Modules.scala 46:47:@9552.4]
  assign _T_62510 = $signed(_T_62509); // @[Modules.scala 46:47:@9553.4]
  assign _T_62512 = $signed(5'sh0) - $signed(io_in_706); // @[Modules.scala 46:37:@9555.4]
  assign _T_62513 = _T_62512[4:0]; // @[Modules.scala 46:37:@9556.4]
  assign _T_62514 = $signed(_T_62513); // @[Modules.scala 46:37:@9557.4]
  assign _T_62515 = $signed(_T_62514) - $signed(io_in_707); // @[Modules.scala 46:47:@9558.4]
  assign _T_62516 = _T_62515[4:0]; // @[Modules.scala 46:47:@9559.4]
  assign _T_62517 = $signed(_T_62516); // @[Modules.scala 46:47:@9560.4]
  assign _T_62529 = $signed(_T_59251) - $signed(io_in_711); // @[Modules.scala 46:47:@9572.4]
  assign _T_62530 = _T_62529[4:0]; // @[Modules.scala 46:47:@9573.4]
  assign _T_62531 = $signed(_T_62530); // @[Modules.scala 46:47:@9574.4]
  assign _T_62543 = $signed(_T_59265) - $signed(io_in_715); // @[Modules.scala 46:47:@9586.4]
  assign _T_62544 = _T_62543[4:0]; // @[Modules.scala 46:47:@9587.4]
  assign _T_62545 = $signed(_T_62544); // @[Modules.scala 46:47:@9588.4]
  assign _T_62547 = $signed(5'sh0) - $signed(io_in_716); // @[Modules.scala 46:37:@9590.4]
  assign _T_62548 = _T_62547[4:0]; // @[Modules.scala 46:37:@9591.4]
  assign _T_62549 = $signed(_T_62548); // @[Modules.scala 46:37:@9592.4]
  assign _T_62550 = $signed(_T_62549) - $signed(io_in_717); // @[Modules.scala 46:47:@9593.4]
  assign _T_62551 = _T_62550[4:0]; // @[Modules.scala 46:47:@9594.4]
  assign _T_62552 = $signed(_T_62551); // @[Modules.scala 46:47:@9595.4]
  assign _T_62576 = $signed(io_in_728) + $signed(io_in_729); // @[Modules.scala 37:46:@9623.4]
  assign _T_62577 = _T_62576[4:0]; // @[Modules.scala 37:46:@9624.4]
  assign _T_62578 = $signed(_T_62577); // @[Modules.scala 37:46:@9625.4]
  assign _T_62579 = $signed(io_in_730) + $signed(io_in_731); // @[Modules.scala 37:46:@9627.4]
  assign _T_62580 = _T_62579[4:0]; // @[Modules.scala 37:46:@9628.4]
  assign _T_62581 = $signed(_T_62580); // @[Modules.scala 37:46:@9629.4]
  assign _T_62582 = $signed(io_in_732) - $signed(io_in_733); // @[Modules.scala 40:46:@9631.4]
  assign _T_62583 = _T_62582[4:0]; // @[Modules.scala 40:46:@9632.4]
  assign _T_62584 = $signed(_T_62583); // @[Modules.scala 40:46:@9633.4]
  assign _T_62634 = $signed(io_in_748) - $signed(io_in_749); // @[Modules.scala 40:46:@9684.4]
  assign _T_62635 = _T_62634[4:0]; // @[Modules.scala 40:46:@9685.4]
  assign _T_62636 = $signed(_T_62635); // @[Modules.scala 40:46:@9686.4]
  assign _T_62638 = $signed(5'sh0) - $signed(io_in_750); // @[Modules.scala 43:37:@9688.4]
  assign _T_62639 = _T_62638[4:0]; // @[Modules.scala 43:37:@9689.4]
  assign _T_62640 = $signed(_T_62639); // @[Modules.scala 43:37:@9690.4]
  assign _T_62641 = $signed(_T_62640) + $signed(io_in_751); // @[Modules.scala 43:47:@9691.4]
  assign _T_62642 = _T_62641[4:0]; // @[Modules.scala 43:47:@9692.4]
  assign _T_62643 = $signed(_T_62642); // @[Modules.scala 43:47:@9693.4]
  assign _T_62647 = $signed(io_in_754) - $signed(io_in_755); // @[Modules.scala 40:46:@9699.4]
  assign _T_62648 = _T_62647[4:0]; // @[Modules.scala 40:46:@9700.4]
  assign _T_62649 = $signed(_T_62648); // @[Modules.scala 40:46:@9701.4]
  assign _T_62654 = $signed(_T_56295) - $signed(io_in_757); // @[Modules.scala 46:47:@9706.4]
  assign _T_62655 = _T_62654[4:0]; // @[Modules.scala 46:47:@9707.4]
  assign _T_62656 = $signed(_T_62655); // @[Modules.scala 46:47:@9708.4]
  assign _T_62733 = $signed(_T_59447) + $signed(io_in_783); // @[Modules.scala 43:47:@9788.4]
  assign _T_62734 = _T_62733[4:0]; // @[Modules.scala 43:47:@9789.4]
  assign _T_62735 = $signed(_T_62734); // @[Modules.scala 43:47:@9790.4]
  assign buffer_2_2 = {{6{_T_60640[4]}},_T_60640}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_3 = {{6{_T_60647[4]}},_T_60647}; // @[Modules.scala 32:22:@8.4]
  assign _T_62739 = $signed(buffer_2_2) + $signed(buffer_2_3); // @[Modules.scala 50:57:@9796.4]
  assign _T_62740 = _T_62739[10:0]; // @[Modules.scala 50:57:@9797.4]
  assign buffer_2_393 = $signed(_T_62740); // @[Modules.scala 50:57:@9798.4]
  assign buffer_2_4 = {{6{_T_60650[4]}},_T_60650}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_5 = {{6{_T_60653[4]}},_T_60653}; // @[Modules.scala 32:22:@8.4]
  assign _T_62742 = $signed(buffer_2_4) + $signed(buffer_2_5); // @[Modules.scala 50:57:@9800.4]
  assign _T_62743 = _T_62742[10:0]; // @[Modules.scala 50:57:@9801.4]
  assign buffer_2_394 = $signed(_T_62743); // @[Modules.scala 50:57:@9802.4]
  assign buffer_2_9 = {{6{_T_60677[4]}},_T_60677}; // @[Modules.scala 32:22:@8.4]
  assign _T_62748 = $signed(buffer_1_8) + $signed(buffer_2_9); // @[Modules.scala 50:57:@9808.4]
  assign _T_62749 = _T_62748[10:0]; // @[Modules.scala 50:57:@9809.4]
  assign buffer_2_396 = $signed(_T_62749); // @[Modules.scala 50:57:@9810.4]
  assign buffer_2_10 = {{6{_T_60680[4]}},_T_60680}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_11 = {{6{_T_60683[4]}},_T_60683}; // @[Modules.scala 32:22:@8.4]
  assign _T_62751 = $signed(buffer_2_10) + $signed(buffer_2_11); // @[Modules.scala 50:57:@9812.4]
  assign _T_62752 = _T_62751[10:0]; // @[Modules.scala 50:57:@9813.4]
  assign buffer_2_397 = $signed(_T_62752); // @[Modules.scala 50:57:@9814.4]
  assign buffer_2_12 = {{6{_T_60690[4]}},_T_60690}; // @[Modules.scala 32:22:@8.4]
  assign _T_62754 = $signed(buffer_2_12) + $signed(buffer_0_13); // @[Modules.scala 50:57:@9816.4]
  assign _T_62755 = _T_62754[10:0]; // @[Modules.scala 50:57:@9817.4]
  assign buffer_2_398 = $signed(_T_62755); // @[Modules.scala 50:57:@9818.4]
  assign buffer_2_15 = {{6{_T_60703[4]}},_T_60703}; // @[Modules.scala 32:22:@8.4]
  assign _T_62757 = $signed(buffer_0_14) + $signed(buffer_2_15); // @[Modules.scala 50:57:@9820.4]
  assign _T_62758 = _T_62757[10:0]; // @[Modules.scala 50:57:@9821.4]
  assign buffer_2_399 = $signed(_T_62758); // @[Modules.scala 50:57:@9822.4]
  assign buffer_2_16 = {{6{_T_60710[4]}},_T_60710}; // @[Modules.scala 32:22:@8.4]
  assign _T_62760 = $signed(buffer_2_16) + $signed(buffer_1_17); // @[Modules.scala 50:57:@9824.4]
  assign _T_62761 = _T_62760[10:0]; // @[Modules.scala 50:57:@9825.4]
  assign buffer_2_400 = $signed(_T_62761); // @[Modules.scala 50:57:@9826.4]
  assign buffer_2_20 = {{6{_T_60722[4]}},_T_60722}; // @[Modules.scala 32:22:@8.4]
  assign _T_62766 = $signed(buffer_2_20) + $signed(buffer_1_21); // @[Modules.scala 50:57:@9832.4]
  assign _T_62767 = _T_62766[10:0]; // @[Modules.scala 50:57:@9833.4]
  assign buffer_2_402 = $signed(_T_62767); // @[Modules.scala 50:57:@9834.4]
  assign _T_62769 = $signed(buffer_0_22) + $signed(buffer_1_23); // @[Modules.scala 50:57:@9836.4]
  assign _T_62770 = _T_62769[10:0]; // @[Modules.scala 50:57:@9837.4]
  assign buffer_2_403 = $signed(_T_62770); // @[Modules.scala 50:57:@9838.4]
  assign buffer_2_26 = {{6{_T_60748[4]}},_T_60748}; // @[Modules.scala 32:22:@8.4]
  assign _T_62775 = $signed(buffer_2_26) + $signed(buffer_1_27); // @[Modules.scala 50:57:@9844.4]
  assign _T_62776 = _T_62775[10:0]; // @[Modules.scala 50:57:@9845.4]
  assign buffer_2_405 = $signed(_T_62776); // @[Modules.scala 50:57:@9846.4]
  assign buffer_2_28 = {{6{_T_60758[4]}},_T_60758}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_29 = {{6{_T_60765[4]}},_T_60765}; // @[Modules.scala 32:22:@8.4]
  assign _T_62778 = $signed(buffer_2_28) + $signed(buffer_2_29); // @[Modules.scala 50:57:@9848.4]
  assign _T_62779 = _T_62778[10:0]; // @[Modules.scala 50:57:@9849.4]
  assign buffer_2_406 = $signed(_T_62779); // @[Modules.scala 50:57:@9850.4]
  assign buffer_2_31 = {{6{_T_60779[4]}},_T_60779}; // @[Modules.scala 32:22:@8.4]
  assign _T_62781 = $signed(buffer_0_30) + $signed(buffer_2_31); // @[Modules.scala 50:57:@9852.4]
  assign _T_62782 = _T_62781[10:0]; // @[Modules.scala 50:57:@9853.4]
  assign buffer_2_407 = $signed(_T_62782); // @[Modules.scala 50:57:@9854.4]
  assign buffer_2_35 = {{6{_T_60795[4]}},_T_60795}; // @[Modules.scala 32:22:@8.4]
  assign _T_62787 = $signed(buffer_1_34) + $signed(buffer_2_35); // @[Modules.scala 50:57:@9860.4]
  assign _T_62788 = _T_62787[10:0]; // @[Modules.scala 50:57:@9861.4]
  assign buffer_2_409 = $signed(_T_62788); // @[Modules.scala 50:57:@9862.4]
  assign buffer_2_39 = {{6{_T_60807[4]}},_T_60807}; // @[Modules.scala 32:22:@8.4]
  assign _T_62793 = $signed(buffer_1_38) + $signed(buffer_2_39); // @[Modules.scala 50:57:@9868.4]
  assign _T_62794 = _T_62793[10:0]; // @[Modules.scala 50:57:@9869.4]
  assign buffer_2_411 = $signed(_T_62794); // @[Modules.scala 50:57:@9870.4]
  assign buffer_2_41 = {{6{_T_60817[4]}},_T_60817}; // @[Modules.scala 32:22:@8.4]
  assign _T_62796 = $signed(buffer_0_40) + $signed(buffer_2_41); // @[Modules.scala 50:57:@9872.4]
  assign _T_62797 = _T_62796[10:0]; // @[Modules.scala 50:57:@9873.4]
  assign buffer_2_412 = $signed(_T_62797); // @[Modules.scala 50:57:@9874.4]
  assign buffer_2_42 = {{6{_T_60824[4]}},_T_60824}; // @[Modules.scala 32:22:@8.4]
  assign _T_62799 = $signed(buffer_2_42) + $signed(buffer_1_43); // @[Modules.scala 50:57:@9876.4]
  assign _T_62800 = _T_62799[10:0]; // @[Modules.scala 50:57:@9877.4]
  assign buffer_2_413 = $signed(_T_62800); // @[Modules.scala 50:57:@9878.4]
  assign buffer_2_44 = {{6{_T_60834[4]}},_T_60834}; // @[Modules.scala 32:22:@8.4]
  assign _T_62802 = $signed(buffer_2_44) + $signed(buffer_0_45); // @[Modules.scala 50:57:@9880.4]
  assign _T_62803 = _T_62802[10:0]; // @[Modules.scala 50:57:@9881.4]
  assign buffer_2_414 = $signed(_T_62803); // @[Modules.scala 50:57:@9882.4]
  assign buffer_2_47 = {{6{_T_60847[4]}},_T_60847}; // @[Modules.scala 32:22:@8.4]
  assign _T_62805 = $signed(buffer_1_46) + $signed(buffer_2_47); // @[Modules.scala 50:57:@9884.4]
  assign _T_62806 = _T_62805[10:0]; // @[Modules.scala 50:57:@9885.4]
  assign buffer_2_415 = $signed(_T_62806); // @[Modules.scala 50:57:@9886.4]
  assign buffer_2_48 = {{6{_T_60854[4]}},_T_60854}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_49 = {{6{_T_60861[4]}},_T_60861}; // @[Modules.scala 32:22:@8.4]
  assign _T_62808 = $signed(buffer_2_48) + $signed(buffer_2_49); // @[Modules.scala 50:57:@9888.4]
  assign _T_62809 = _T_62808[10:0]; // @[Modules.scala 50:57:@9889.4]
  assign buffer_2_416 = $signed(_T_62809); // @[Modules.scala 50:57:@9890.4]
  assign buffer_2_50 = {{6{_T_60864[4]}},_T_60864}; // @[Modules.scala 32:22:@8.4]
  assign _T_62811 = $signed(buffer_2_50) + $signed(buffer_0_51); // @[Modules.scala 50:57:@9892.4]
  assign _T_62812 = _T_62811[10:0]; // @[Modules.scala 50:57:@9893.4]
  assign buffer_2_417 = $signed(_T_62812); // @[Modules.scala 50:57:@9894.4]
  assign buffer_2_54 = {{6{_T_60880[4]}},_T_60880}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_55 = {{6{_T_60887[4]}},_T_60887}; // @[Modules.scala 32:22:@8.4]
  assign _T_62817 = $signed(buffer_2_54) + $signed(buffer_2_55); // @[Modules.scala 50:57:@9900.4]
  assign _T_62818 = _T_62817[10:0]; // @[Modules.scala 50:57:@9901.4]
  assign buffer_2_419 = $signed(_T_62818); // @[Modules.scala 50:57:@9902.4]
  assign buffer_2_58 = {{6{_T_60908[4]}},_T_60908}; // @[Modules.scala 32:22:@8.4]
  assign _T_62823 = $signed(buffer_2_58) + $signed(buffer_1_59); // @[Modules.scala 50:57:@9908.4]
  assign _T_62824 = _T_62823[10:0]; // @[Modules.scala 50:57:@9909.4]
  assign buffer_2_421 = $signed(_T_62824); // @[Modules.scala 50:57:@9910.4]
  assign buffer_2_65 = {{6{_T_60957[4]}},_T_60957}; // @[Modules.scala 32:22:@8.4]
  assign _T_62832 = $signed(buffer_0_64) + $signed(buffer_2_65); // @[Modules.scala 50:57:@9920.4]
  assign _T_62833 = _T_62832[10:0]; // @[Modules.scala 50:57:@9921.4]
  assign buffer_2_424 = $signed(_T_62833); // @[Modules.scala 50:57:@9922.4]
  assign buffer_2_70 = {{6{_T_60984[4]}},_T_60984}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_71 = {{6{_T_60987[4]}},_T_60987}; // @[Modules.scala 32:22:@8.4]
  assign _T_62841 = $signed(buffer_2_70) + $signed(buffer_2_71); // @[Modules.scala 50:57:@9932.4]
  assign _T_62842 = _T_62841[10:0]; // @[Modules.scala 50:57:@9933.4]
  assign buffer_2_427 = $signed(_T_62842); // @[Modules.scala 50:57:@9934.4]
  assign buffer_2_74 = {{6{_T_61008[4]}},_T_61008}; // @[Modules.scala 32:22:@8.4]
  assign _T_62847 = $signed(buffer_2_74) + $signed(buffer_0_75); // @[Modules.scala 50:57:@9940.4]
  assign _T_62848 = _T_62847[10:0]; // @[Modules.scala 50:57:@9941.4]
  assign buffer_2_429 = $signed(_T_62848); // @[Modules.scala 50:57:@9942.4]
  assign buffer_2_79 = {{6{_T_61043[4]}},_T_61043}; // @[Modules.scala 32:22:@8.4]
  assign _T_62853 = $signed(buffer_0_78) + $signed(buffer_2_79); // @[Modules.scala 50:57:@9948.4]
  assign _T_62854 = _T_62853[10:0]; // @[Modules.scala 50:57:@9949.4]
  assign buffer_2_431 = $signed(_T_62854); // @[Modules.scala 50:57:@9950.4]
  assign buffer_2_80 = {{6{_T_61046[4]}},_T_61046}; // @[Modules.scala 32:22:@8.4]
  assign _T_62856 = $signed(buffer_2_80) + $signed(buffer_0_81); // @[Modules.scala 50:57:@9952.4]
  assign _T_62857 = _T_62856[10:0]; // @[Modules.scala 50:57:@9953.4]
  assign buffer_2_432 = $signed(_T_62857); // @[Modules.scala 50:57:@9954.4]
  assign buffer_2_82 = {{6{_T_61052[4]}},_T_61052}; // @[Modules.scala 32:22:@8.4]
  assign _T_62859 = $signed(buffer_2_82) + $signed(buffer_1_83); // @[Modules.scala 50:57:@9956.4]
  assign _T_62860 = _T_62859[10:0]; // @[Modules.scala 50:57:@9957.4]
  assign buffer_2_433 = $signed(_T_62860); // @[Modules.scala 50:57:@9958.4]
  assign buffer_2_84 = {{6{_T_61058[4]}},_T_61058}; // @[Modules.scala 32:22:@8.4]
  assign _T_62862 = $signed(buffer_2_84) + $signed(buffer_0_85); // @[Modules.scala 50:57:@9960.4]
  assign _T_62863 = _T_62862[10:0]; // @[Modules.scala 50:57:@9961.4]
  assign buffer_2_434 = $signed(_T_62863); // @[Modules.scala 50:57:@9962.4]
  assign buffer_2_86 = {{6{_T_61072[4]}},_T_61072}; // @[Modules.scala 32:22:@8.4]
  assign _T_62865 = $signed(buffer_2_86) + $signed(buffer_0_87); // @[Modules.scala 50:57:@9964.4]
  assign _T_62866 = _T_62865[10:0]; // @[Modules.scala 50:57:@9965.4]
  assign buffer_2_435 = $signed(_T_62866); // @[Modules.scala 50:57:@9966.4]
  assign buffer_2_93 = {{6{_T_61121[4]}},_T_61121}; // @[Modules.scala 32:22:@8.4]
  assign _T_62874 = $signed(buffer_0_92) + $signed(buffer_2_93); // @[Modules.scala 50:57:@9976.4]
  assign _T_62875 = _T_62874[10:0]; // @[Modules.scala 50:57:@9977.4]
  assign buffer_2_438 = $signed(_T_62875); // @[Modules.scala 50:57:@9978.4]
  assign buffer_2_95 = {{6{_T_61131[4]}},_T_61131}; // @[Modules.scala 32:22:@8.4]
  assign _T_62877 = $signed(buffer_0_94) + $signed(buffer_2_95); // @[Modules.scala 50:57:@9980.4]
  assign _T_62878 = _T_62877[10:0]; // @[Modules.scala 50:57:@9981.4]
  assign buffer_2_439 = $signed(_T_62878); // @[Modules.scala 50:57:@9982.4]
  assign buffer_2_96 = {{6{_T_61134[4]}},_T_61134}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_97 = {{6{_T_61137[4]}},_T_61137}; // @[Modules.scala 32:22:@8.4]
  assign _T_62880 = $signed(buffer_2_96) + $signed(buffer_2_97); // @[Modules.scala 50:57:@9984.4]
  assign _T_62881 = _T_62880[10:0]; // @[Modules.scala 50:57:@9985.4]
  assign buffer_2_440 = $signed(_T_62881); // @[Modules.scala 50:57:@9986.4]
  assign buffer_2_99 = {{6{_T_61147[4]}},_T_61147}; // @[Modules.scala 32:22:@8.4]
  assign _T_62883 = $signed(buffer_0_98) + $signed(buffer_2_99); // @[Modules.scala 50:57:@9988.4]
  assign _T_62884 = _T_62883[10:0]; // @[Modules.scala 50:57:@9989.4]
  assign buffer_2_441 = $signed(_T_62884); // @[Modules.scala 50:57:@9990.4]
  assign buffer_2_103 = {{6{_T_61175[4]}},_T_61175}; // @[Modules.scala 32:22:@8.4]
  assign _T_62889 = $signed(buffer_0_102) + $signed(buffer_2_103); // @[Modules.scala 50:57:@9996.4]
  assign _T_62890 = _T_62889[10:0]; // @[Modules.scala 50:57:@9997.4]
  assign buffer_2_443 = $signed(_T_62890); // @[Modules.scala 50:57:@9998.4]
  assign buffer_2_104 = {{6{_T_61182[4]}},_T_61182}; // @[Modules.scala 32:22:@8.4]
  assign _T_62892 = $signed(buffer_2_104) + $signed(buffer_0_105); // @[Modules.scala 50:57:@10000.4]
  assign _T_62893 = _T_62892[10:0]; // @[Modules.scala 50:57:@10001.4]
  assign buffer_2_444 = $signed(_T_62893); // @[Modules.scala 50:57:@10002.4]
  assign buffer_2_107 = {{6{_T_61191[4]}},_T_61191}; // @[Modules.scala 32:22:@8.4]
  assign _T_62895 = $signed(buffer_0_106) + $signed(buffer_2_107); // @[Modules.scala 50:57:@10004.4]
  assign _T_62896 = _T_62895[10:0]; // @[Modules.scala 50:57:@10005.4]
  assign buffer_2_445 = $signed(_T_62896); // @[Modules.scala 50:57:@10006.4]
  assign buffer_2_109 = {{6{_T_61201[4]}},_T_61201}; // @[Modules.scala 32:22:@8.4]
  assign _T_62898 = $signed(buffer_1_108) + $signed(buffer_2_109); // @[Modules.scala 50:57:@10008.4]
  assign _T_62899 = _T_62898[10:0]; // @[Modules.scala 50:57:@10009.4]
  assign buffer_2_446 = $signed(_T_62899); // @[Modules.scala 50:57:@10010.4]
  assign buffer_2_111 = {{6{_T_61207[4]}},_T_61207}; // @[Modules.scala 32:22:@8.4]
  assign _T_62901 = $signed(buffer_1_110) + $signed(buffer_2_111); // @[Modules.scala 50:57:@10012.4]
  assign _T_62902 = _T_62901[10:0]; // @[Modules.scala 50:57:@10013.4]
  assign buffer_2_447 = $signed(_T_62902); // @[Modules.scala 50:57:@10014.4]
  assign buffer_2_117 = {{6{_T_61249[4]}},_T_61249}; // @[Modules.scala 32:22:@8.4]
  assign _T_62910 = $signed(buffer_0_116) + $signed(buffer_2_117); // @[Modules.scala 50:57:@10024.4]
  assign _T_62911 = _T_62910[10:0]; // @[Modules.scala 50:57:@10025.4]
  assign buffer_2_450 = $signed(_T_62911); // @[Modules.scala 50:57:@10026.4]
  assign buffer_2_130 = {{6{_T_61332[4]}},_T_61332}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_131 = {{6{_T_61339[4]}},_T_61339}; // @[Modules.scala 32:22:@8.4]
  assign _T_62931 = $signed(buffer_2_130) + $signed(buffer_2_131); // @[Modules.scala 50:57:@10052.4]
  assign _T_62932 = _T_62931[10:0]; // @[Modules.scala 50:57:@10053.4]
  assign buffer_2_457 = $signed(_T_62932); // @[Modules.scala 50:57:@10054.4]
  assign buffer_2_143 = {{6{_T_61415[4]}},_T_61415}; // @[Modules.scala 32:22:@8.4]
  assign _T_62949 = $signed(buffer_0_142) + $signed(buffer_2_143); // @[Modules.scala 50:57:@10076.4]
  assign _T_62950 = _T_62949[10:0]; // @[Modules.scala 50:57:@10077.4]
  assign buffer_2_463 = $signed(_T_62950); // @[Modules.scala 50:57:@10078.4]
  assign buffer_2_144 = {{6{_T_61418[4]}},_T_61418}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_145 = {{6{_T_61421[4]}},_T_61421}; // @[Modules.scala 32:22:@8.4]
  assign _T_62952 = $signed(buffer_2_144) + $signed(buffer_2_145); // @[Modules.scala 50:57:@10080.4]
  assign _T_62953 = _T_62952[10:0]; // @[Modules.scala 50:57:@10081.4]
  assign buffer_2_464 = $signed(_T_62953); // @[Modules.scala 50:57:@10082.4]
  assign buffer_2_152 = {{6{_T_61470[4]}},_T_61470}; // @[Modules.scala 32:22:@8.4]
  assign _T_62964 = $signed(buffer_2_152) + $signed(buffer_1_153); // @[Modules.scala 50:57:@10096.4]
  assign _T_62965 = _T_62964[10:0]; // @[Modules.scala 50:57:@10097.4]
  assign buffer_2_468 = $signed(_T_62965); // @[Modules.scala 50:57:@10098.4]
  assign buffer_2_157 = {{6{_T_61497[4]}},_T_61497}; // @[Modules.scala 32:22:@8.4]
  assign _T_62970 = $signed(buffer_0_156) + $signed(buffer_2_157); // @[Modules.scala 50:57:@10104.4]
  assign _T_62971 = _T_62970[10:0]; // @[Modules.scala 50:57:@10105.4]
  assign buffer_2_470 = $signed(_T_62971); // @[Modules.scala 50:57:@10106.4]
  assign buffer_2_160 = {{6{_T_61506[4]}},_T_61506}; // @[Modules.scala 32:22:@8.4]
  assign _T_62976 = $signed(buffer_2_160) + $signed(buffer_1_161); // @[Modules.scala 50:57:@10112.4]
  assign _T_62977 = _T_62976[10:0]; // @[Modules.scala 50:57:@10113.4]
  assign buffer_2_472 = $signed(_T_62977); // @[Modules.scala 50:57:@10114.4]
  assign _T_62982 = $signed(buffer_1_164) + $signed(buffer_0_165); // @[Modules.scala 50:57:@10120.4]
  assign _T_62983 = _T_62982[10:0]; // @[Modules.scala 50:57:@10121.4]
  assign buffer_2_474 = $signed(_T_62983); // @[Modules.scala 50:57:@10122.4]
  assign buffer_2_166 = {{6{_T_61544[4]}},_T_61544}; // @[Modules.scala 32:22:@8.4]
  assign _T_62985 = $signed(buffer_2_166) + $signed(buffer_1_167); // @[Modules.scala 50:57:@10124.4]
  assign _T_62986 = _T_62985[10:0]; // @[Modules.scala 50:57:@10125.4]
  assign buffer_2_475 = $signed(_T_62986); // @[Modules.scala 50:57:@10126.4]
  assign buffer_2_177 = {{6{_T_61589[4]}},_T_61589}; // @[Modules.scala 32:22:@8.4]
  assign _T_63000 = $signed(buffer_1_176) + $signed(buffer_2_177); // @[Modules.scala 50:57:@10144.4]
  assign _T_63001 = _T_63000[10:0]; // @[Modules.scala 50:57:@10145.4]
  assign buffer_2_480 = $signed(_T_63001); // @[Modules.scala 50:57:@10146.4]
  assign buffer_2_179 = {{6{_T_61603[4]}},_T_61603}; // @[Modules.scala 32:22:@8.4]
  assign _T_63003 = $signed(buffer_1_178) + $signed(buffer_2_179); // @[Modules.scala 50:57:@10148.4]
  assign _T_63004 = _T_63003[10:0]; // @[Modules.scala 50:57:@10149.4]
  assign buffer_2_481 = $signed(_T_63004); // @[Modules.scala 50:57:@10150.4]
  assign buffer_2_180 = {{6{_T_61610[4]}},_T_61610}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_181 = {{6{_T_61613[4]}},_T_61613}; // @[Modules.scala 32:22:@8.4]
  assign _T_63006 = $signed(buffer_2_180) + $signed(buffer_2_181); // @[Modules.scala 50:57:@10152.4]
  assign _T_63007 = _T_63006[10:0]; // @[Modules.scala 50:57:@10153.4]
  assign buffer_2_482 = $signed(_T_63007); // @[Modules.scala 50:57:@10154.4]
  assign buffer_2_192 = {{6{_T_61658[4]}},_T_61658}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_193 = {{6{_T_61665[4]}},_T_61665}; // @[Modules.scala 32:22:@8.4]
  assign _T_63024 = $signed(buffer_2_192) + $signed(buffer_2_193); // @[Modules.scala 50:57:@10176.4]
  assign _T_63025 = _T_63024[10:0]; // @[Modules.scala 50:57:@10177.4]
  assign buffer_2_488 = $signed(_T_63025); // @[Modules.scala 50:57:@10178.4]
  assign buffer_2_194 = {{6{_T_61672[4]}},_T_61672}; // @[Modules.scala 32:22:@8.4]
  assign _T_63027 = $signed(buffer_2_194) + $signed(buffer_1_195); // @[Modules.scala 50:57:@10180.4]
  assign _T_63028 = _T_63027[10:0]; // @[Modules.scala 50:57:@10181.4]
  assign buffer_2_489 = $signed(_T_63028); // @[Modules.scala 50:57:@10182.4]
  assign buffer_2_205 = {{6{_T_61717[4]}},_T_61717}; // @[Modules.scala 32:22:@8.4]
  assign _T_63042 = $signed(buffer_0_204) + $signed(buffer_2_205); // @[Modules.scala 50:57:@10200.4]
  assign _T_63043 = _T_63042[10:0]; // @[Modules.scala 50:57:@10201.4]
  assign buffer_2_494 = $signed(_T_63043); // @[Modules.scala 50:57:@10202.4]
  assign buffer_2_208 = {{6{_T_61730[4]}},_T_61730}; // @[Modules.scala 32:22:@8.4]
  assign _T_63048 = $signed(buffer_2_208) + $signed(buffer_1_209); // @[Modules.scala 50:57:@10208.4]
  assign _T_63049 = _T_63048[10:0]; // @[Modules.scala 50:57:@10209.4]
  assign buffer_2_496 = $signed(_T_63049); // @[Modules.scala 50:57:@10210.4]
  assign buffer_2_211 = {{6{_T_61747[4]}},_T_61747}; // @[Modules.scala 32:22:@8.4]
  assign _T_63051 = $signed(buffer_0_210) + $signed(buffer_2_211); // @[Modules.scala 50:57:@10212.4]
  assign _T_63052 = _T_63051[10:0]; // @[Modules.scala 50:57:@10213.4]
  assign buffer_2_497 = $signed(_T_63052); // @[Modules.scala 50:57:@10214.4]
  assign buffer_2_212 = {{6{_T_61754[4]}},_T_61754}; // @[Modules.scala 32:22:@8.4]
  assign _T_63054 = $signed(buffer_2_212) + $signed(buffer_0_213); // @[Modules.scala 50:57:@10216.4]
  assign _T_63055 = _T_63054[10:0]; // @[Modules.scala 50:57:@10217.4]
  assign buffer_2_498 = $signed(_T_63055); // @[Modules.scala 50:57:@10218.4]
  assign buffer_2_215 = {{6{_T_61767[4]}},_T_61767}; // @[Modules.scala 32:22:@8.4]
  assign _T_63057 = $signed(buffer_0_214) + $signed(buffer_2_215); // @[Modules.scala 50:57:@10220.4]
  assign _T_63058 = _T_63057[10:0]; // @[Modules.scala 50:57:@10221.4]
  assign buffer_2_499 = $signed(_T_63058); // @[Modules.scala 50:57:@10222.4]
  assign buffer_2_219 = {{6{_T_61787[4]}},_T_61787}; // @[Modules.scala 32:22:@8.4]
  assign _T_63063 = $signed(buffer_1_218) + $signed(buffer_2_219); // @[Modules.scala 50:57:@10228.4]
  assign _T_63064 = _T_63063[10:0]; // @[Modules.scala 50:57:@10229.4]
  assign buffer_2_501 = $signed(_T_63064); // @[Modules.scala 50:57:@10230.4]
  assign buffer_2_220 = {{6{_T_61794[4]}},_T_61794}; // @[Modules.scala 32:22:@8.4]
  assign _T_63066 = $signed(buffer_2_220) + $signed(buffer_1_221); // @[Modules.scala 50:57:@10232.4]
  assign _T_63067 = _T_63066[10:0]; // @[Modules.scala 50:57:@10233.4]
  assign buffer_2_502 = $signed(_T_63067); // @[Modules.scala 50:57:@10234.4]
  assign _T_63072 = $signed(buffer_1_224) + $signed(buffer_0_225); // @[Modules.scala 50:57:@10240.4]
  assign _T_63073 = _T_63072[10:0]; // @[Modules.scala 50:57:@10241.4]
  assign buffer_2_504 = $signed(_T_63073); // @[Modules.scala 50:57:@10242.4]
  assign buffer_2_227 = {{6{_T_61839[4]}},_T_61839}; // @[Modules.scala 32:22:@8.4]
  assign _T_63075 = $signed(buffer_1_226) + $signed(buffer_2_227); // @[Modules.scala 50:57:@10244.4]
  assign _T_63076 = _T_63075[10:0]; // @[Modules.scala 50:57:@10245.4]
  assign buffer_2_505 = $signed(_T_63076); // @[Modules.scala 50:57:@10246.4]
  assign buffer_2_228 = {{6{_T_61842[4]}},_T_61842}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_229 = {{6{_T_61849[4]}},_T_61849}; // @[Modules.scala 32:22:@8.4]
  assign _T_63078 = $signed(buffer_2_228) + $signed(buffer_2_229); // @[Modules.scala 50:57:@10248.4]
  assign _T_63079 = _T_63078[10:0]; // @[Modules.scala 50:57:@10249.4]
  assign buffer_2_506 = $signed(_T_63079); // @[Modules.scala 50:57:@10250.4]
  assign buffer_2_230 = {{6{_T_61852[4]}},_T_61852}; // @[Modules.scala 32:22:@8.4]
  assign _T_63081 = $signed(buffer_2_230) + $signed(buffer_0_231); // @[Modules.scala 50:57:@10252.4]
  assign _T_63082 = _T_63081[10:0]; // @[Modules.scala 50:57:@10253.4]
  assign buffer_2_507 = $signed(_T_63082); // @[Modules.scala 50:57:@10254.4]
  assign buffer_2_232 = {{6{_T_61862[4]}},_T_61862}; // @[Modules.scala 32:22:@8.4]
  assign _T_63084 = $signed(buffer_2_232) + $signed(buffer_0_233); // @[Modules.scala 50:57:@10256.4]
  assign _T_63085 = _T_63084[10:0]; // @[Modules.scala 50:57:@10257.4]
  assign buffer_2_508 = $signed(_T_63085); // @[Modules.scala 50:57:@10258.4]
  assign buffer_2_234 = {{6{_T_61872[4]}},_T_61872}; // @[Modules.scala 32:22:@8.4]
  assign _T_63087 = $signed(buffer_2_234) + $signed(buffer_1_235); // @[Modules.scala 50:57:@10260.4]
  assign _T_63088 = _T_63087[10:0]; // @[Modules.scala 50:57:@10261.4]
  assign buffer_2_509 = $signed(_T_63088); // @[Modules.scala 50:57:@10262.4]
  assign buffer_2_238 = {{6{_T_61892[4]}},_T_61892}; // @[Modules.scala 32:22:@8.4]
  assign _T_63093 = $signed(buffer_2_238) + $signed(buffer_0_239); // @[Modules.scala 50:57:@10268.4]
  assign _T_63094 = _T_63093[10:0]; // @[Modules.scala 50:57:@10269.4]
  assign buffer_2_511 = $signed(_T_63094); // @[Modules.scala 50:57:@10270.4]
  assign buffer_2_241 = {{6{_T_61909[4]}},_T_61909}; // @[Modules.scala 32:22:@8.4]
  assign _T_63096 = $signed(buffer_0_240) + $signed(buffer_2_241); // @[Modules.scala 50:57:@10272.4]
  assign _T_63097 = _T_63096[10:0]; // @[Modules.scala 50:57:@10273.4]
  assign buffer_2_512 = $signed(_T_63097); // @[Modules.scala 50:57:@10274.4]
  assign buffer_2_242 = {{6{_T_61916[4]}},_T_61916}; // @[Modules.scala 32:22:@8.4]
  assign _T_63099 = $signed(buffer_2_242) + $signed(buffer_0_243); // @[Modules.scala 50:57:@10276.4]
  assign _T_63100 = _T_63099[10:0]; // @[Modules.scala 50:57:@10277.4]
  assign buffer_2_513 = $signed(_T_63100); // @[Modules.scala 50:57:@10278.4]
  assign buffer_2_244 = {{6{_T_61922[4]}},_T_61922}; // @[Modules.scala 32:22:@8.4]
  assign _T_63102 = $signed(buffer_2_244) + $signed(buffer_0_245); // @[Modules.scala 50:57:@10280.4]
  assign _T_63103 = _T_63102[10:0]; // @[Modules.scala 50:57:@10281.4]
  assign buffer_2_514 = $signed(_T_63103); // @[Modules.scala 50:57:@10282.4]
  assign buffer_2_249 = {{6{_T_61945[4]}},_T_61945}; // @[Modules.scala 32:22:@8.4]
  assign _T_63108 = $signed(buffer_1_248) + $signed(buffer_2_249); // @[Modules.scala 50:57:@10288.4]
  assign _T_63109 = _T_63108[10:0]; // @[Modules.scala 50:57:@10289.4]
  assign buffer_2_516 = $signed(_T_63109); // @[Modules.scala 50:57:@10290.4]
  assign buffer_2_253 = {{6{_T_61973[4]}},_T_61973}; // @[Modules.scala 32:22:@8.4]
  assign _T_63114 = $signed(buffer_0_252) + $signed(buffer_2_253); // @[Modules.scala 50:57:@10296.4]
  assign _T_63115 = _T_63114[10:0]; // @[Modules.scala 50:57:@10297.4]
  assign buffer_2_518 = $signed(_T_63115); // @[Modules.scala 50:57:@10298.4]
  assign buffer_2_258 = {{6{_T_62000[4]}},_T_62000}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_259 = {{6{_T_62003[4]}},_T_62003}; // @[Modules.scala 32:22:@8.4]
  assign _T_63123 = $signed(buffer_2_258) + $signed(buffer_2_259); // @[Modules.scala 50:57:@10308.4]
  assign _T_63124 = _T_63123[10:0]; // @[Modules.scala 50:57:@10309.4]
  assign buffer_2_521 = $signed(_T_63124); // @[Modules.scala 50:57:@10310.4]
  assign buffer_2_260 = {{6{_T_62010[4]}},_T_62010}; // @[Modules.scala 32:22:@8.4]
  assign _T_63126 = $signed(buffer_2_260) + $signed(buffer_0_261); // @[Modules.scala 50:57:@10312.4]
  assign _T_63127 = _T_63126[10:0]; // @[Modules.scala 50:57:@10313.4]
  assign buffer_2_522 = $signed(_T_63127); // @[Modules.scala 50:57:@10314.4]
  assign buffer_2_262 = {{6{_T_62024[4]}},_T_62024}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_263 = {{6{_T_62031[4]}},_T_62031}; // @[Modules.scala 32:22:@8.4]
  assign _T_63129 = $signed(buffer_2_262) + $signed(buffer_2_263); // @[Modules.scala 50:57:@10316.4]
  assign _T_63130 = _T_63129[10:0]; // @[Modules.scala 50:57:@10317.4]
  assign buffer_2_523 = $signed(_T_63130); // @[Modules.scala 50:57:@10318.4]
  assign buffer_2_266 = {{6{_T_62052[4]}},_T_62052}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_267 = {{6{_T_62059[4]}},_T_62059}; // @[Modules.scala 32:22:@8.4]
  assign _T_63135 = $signed(buffer_2_266) + $signed(buffer_2_267); // @[Modules.scala 50:57:@10324.4]
  assign _T_63136 = _T_63135[10:0]; // @[Modules.scala 50:57:@10325.4]
  assign buffer_2_525 = $signed(_T_63136); // @[Modules.scala 50:57:@10326.4]
  assign buffer_2_272 = {{6{_T_62094[4]}},_T_62094}; // @[Modules.scala 32:22:@8.4]
  assign _T_63144 = $signed(buffer_2_272) + $signed(buffer_1_273); // @[Modules.scala 50:57:@10336.4]
  assign _T_63145 = _T_63144[10:0]; // @[Modules.scala 50:57:@10337.4]
  assign buffer_2_528 = $signed(_T_63145); // @[Modules.scala 50:57:@10338.4]
  assign buffer_2_274 = {{6{_T_62108[4]}},_T_62108}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_275 = {{6{_T_62115[4]}},_T_62115}; // @[Modules.scala 32:22:@8.4]
  assign _T_63147 = $signed(buffer_2_274) + $signed(buffer_2_275); // @[Modules.scala 50:57:@10340.4]
  assign _T_63148 = _T_63147[10:0]; // @[Modules.scala 50:57:@10341.4]
  assign buffer_2_529 = $signed(_T_63148); // @[Modules.scala 50:57:@10342.4]
  assign buffer_2_276 = {{6{_T_62118[4]}},_T_62118}; // @[Modules.scala 32:22:@8.4]
  assign _T_63150 = $signed(buffer_2_276) + $signed(buffer_0_277); // @[Modules.scala 50:57:@10344.4]
  assign _T_63151 = _T_63150[10:0]; // @[Modules.scala 50:57:@10345.4]
  assign buffer_2_530 = $signed(_T_63151); // @[Modules.scala 50:57:@10346.4]
  assign _T_63153 = $signed(buffer_1_278) + $signed(buffer_0_279); // @[Modules.scala 50:57:@10348.4]
  assign _T_63154 = _T_63153[10:0]; // @[Modules.scala 50:57:@10349.4]
  assign buffer_2_531 = $signed(_T_63154); // @[Modules.scala 50:57:@10350.4]
  assign buffer_2_280 = {{6{_T_62142[4]}},_T_62142}; // @[Modules.scala 32:22:@8.4]
  assign _T_63156 = $signed(buffer_2_280) + $signed(buffer_0_281); // @[Modules.scala 50:57:@10352.4]
  assign _T_63157 = _T_63156[10:0]; // @[Modules.scala 50:57:@10353.4]
  assign buffer_2_532 = $signed(_T_63157); // @[Modules.scala 50:57:@10354.4]
  assign buffer_2_286 = {{6{_T_62184[4]}},_T_62184}; // @[Modules.scala 32:22:@8.4]
  assign _T_63165 = $signed(buffer_2_286) + $signed(buffer_1_287); // @[Modules.scala 50:57:@10364.4]
  assign _T_63166 = _T_63165[10:0]; // @[Modules.scala 50:57:@10365.4]
  assign buffer_2_535 = $signed(_T_63166); // @[Modules.scala 50:57:@10366.4]
  assign _T_63168 = $signed(buffer_0_288) + $signed(buffer_1_289); // @[Modules.scala 50:57:@10368.4]
  assign _T_63169 = _T_63168[10:0]; // @[Modules.scala 50:57:@10369.4]
  assign buffer_2_536 = $signed(_T_63169); // @[Modules.scala 50:57:@10370.4]
  assign buffer_2_290 = {{6{_T_62200[4]}},_T_62200}; // @[Modules.scala 32:22:@8.4]
  assign _T_63171 = $signed(buffer_2_290) + $signed(buffer_0_291); // @[Modules.scala 50:57:@10372.4]
  assign _T_63172 = _T_63171[10:0]; // @[Modules.scala 50:57:@10373.4]
  assign buffer_2_537 = $signed(_T_63172); // @[Modules.scala 50:57:@10374.4]
  assign buffer_2_294 = {{6{_T_62224[4]}},_T_62224}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_295 = {{6{_T_62227[4]}},_T_62227}; // @[Modules.scala 32:22:@8.4]
  assign _T_63177 = $signed(buffer_2_294) + $signed(buffer_2_295); // @[Modules.scala 50:57:@10380.4]
  assign _T_63178 = _T_63177[10:0]; // @[Modules.scala 50:57:@10381.4]
  assign buffer_2_539 = $signed(_T_63178); // @[Modules.scala 50:57:@10382.4]
  assign buffer_2_297 = {{6{_T_62241[4]}},_T_62241}; // @[Modules.scala 32:22:@8.4]
  assign _T_63180 = $signed(buffer_0_296) + $signed(buffer_2_297); // @[Modules.scala 50:57:@10384.4]
  assign _T_63181 = _T_63180[10:0]; // @[Modules.scala 50:57:@10385.4]
  assign buffer_2_540 = $signed(_T_63181); // @[Modules.scala 50:57:@10386.4]
  assign buffer_2_298 = {{6{_T_62244[4]}},_T_62244}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_299 = {{6{_T_62247[4]}},_T_62247}; // @[Modules.scala 32:22:@8.4]
  assign _T_63183 = $signed(buffer_2_298) + $signed(buffer_2_299); // @[Modules.scala 50:57:@10388.4]
  assign _T_63184 = _T_63183[10:0]; // @[Modules.scala 50:57:@10389.4]
  assign buffer_2_541 = $signed(_T_63184); // @[Modules.scala 50:57:@10390.4]
  assign buffer_2_300 = {{6{_T_62254[4]}},_T_62254}; // @[Modules.scala 32:22:@8.4]
  assign _T_63186 = $signed(buffer_2_300) + $signed(buffer_1_301); // @[Modules.scala 50:57:@10392.4]
  assign _T_63187 = _T_63186[10:0]; // @[Modules.scala 50:57:@10393.4]
  assign buffer_2_542 = $signed(_T_63187); // @[Modules.scala 50:57:@10394.4]
  assign buffer_2_302 = {{6{_T_62264[4]}},_T_62264}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_303 = {{6{_T_62271[4]}},_T_62271}; // @[Modules.scala 32:22:@8.4]
  assign _T_63189 = $signed(buffer_2_302) + $signed(buffer_2_303); // @[Modules.scala 50:57:@10396.4]
  assign _T_63190 = _T_63189[10:0]; // @[Modules.scala 50:57:@10397.4]
  assign buffer_2_543 = $signed(_T_63190); // @[Modules.scala 50:57:@10398.4]
  assign buffer_2_304 = {{6{_T_62274[4]}},_T_62274}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_305 = {{6{_T_62277[4]}},_T_62277}; // @[Modules.scala 32:22:@8.4]
  assign _T_63192 = $signed(buffer_2_304) + $signed(buffer_2_305); // @[Modules.scala 50:57:@10400.4]
  assign _T_63193 = _T_63192[10:0]; // @[Modules.scala 50:57:@10401.4]
  assign buffer_2_544 = $signed(_T_63193); // @[Modules.scala 50:57:@10402.4]
  assign buffer_2_308 = {{6{_T_62294[4]}},_T_62294}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_309 = {{6{_T_62301[4]}},_T_62301}; // @[Modules.scala 32:22:@8.4]
  assign _T_63198 = $signed(buffer_2_308) + $signed(buffer_2_309); // @[Modules.scala 50:57:@10408.4]
  assign _T_63199 = _T_63198[10:0]; // @[Modules.scala 50:57:@10409.4]
  assign buffer_2_546 = $signed(_T_63199); // @[Modules.scala 50:57:@10410.4]
  assign buffer_2_312 = {{6{_T_62318[4]}},_T_62318}; // @[Modules.scala 32:22:@8.4]
  assign _T_63204 = $signed(buffer_2_312) + $signed(buffer_0_313); // @[Modules.scala 50:57:@10416.4]
  assign _T_63205 = _T_63204[10:0]; // @[Modules.scala 50:57:@10417.4]
  assign buffer_2_548 = $signed(_T_63205); // @[Modules.scala 50:57:@10418.4]
  assign buffer_2_317 = {{6{_T_62345[4]}},_T_62345}; // @[Modules.scala 32:22:@8.4]
  assign _T_63210 = $signed(buffer_1_316) + $signed(buffer_2_317); // @[Modules.scala 50:57:@10424.4]
  assign _T_63211 = _T_63210[10:0]; // @[Modules.scala 50:57:@10425.4]
  assign buffer_2_550 = $signed(_T_63211); // @[Modules.scala 50:57:@10426.4]
  assign buffer_2_322 = {{6{_T_62364[4]}},_T_62364}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_323 = {{6{_T_62367[4]}},_T_62367}; // @[Modules.scala 32:22:@8.4]
  assign _T_63219 = $signed(buffer_2_322) + $signed(buffer_2_323); // @[Modules.scala 50:57:@10436.4]
  assign _T_63220 = _T_63219[10:0]; // @[Modules.scala 50:57:@10437.4]
  assign buffer_2_553 = $signed(_T_63220); // @[Modules.scala 50:57:@10438.4]
  assign buffer_2_324 = {{6{_T_62374[4]}},_T_62374}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_325 = {{6{_T_62377[4]}},_T_62377}; // @[Modules.scala 32:22:@8.4]
  assign _T_63222 = $signed(buffer_2_324) + $signed(buffer_2_325); // @[Modules.scala 50:57:@10440.4]
  assign _T_63223 = _T_63222[10:0]; // @[Modules.scala 50:57:@10441.4]
  assign buffer_2_554 = $signed(_T_63223); // @[Modules.scala 50:57:@10442.4]
  assign _T_63225 = $signed(buffer_1_326) + $signed(buffer_0_327); // @[Modules.scala 50:57:@10444.4]
  assign _T_63226 = _T_63225[10:0]; // @[Modules.scala 50:57:@10445.4]
  assign buffer_2_555 = $signed(_T_63226); // @[Modules.scala 50:57:@10446.4]
  assign buffer_2_328 = {{6{_T_62390[4]}},_T_62390}; // @[Modules.scala 32:22:@8.4]
  assign _T_63228 = $signed(buffer_2_328) + $signed(buffer_1_329); // @[Modules.scala 50:57:@10448.4]
  assign _T_63229 = _T_63228[10:0]; // @[Modules.scala 50:57:@10449.4]
  assign buffer_2_556 = $signed(_T_63229); // @[Modules.scala 50:57:@10450.4]
  assign buffer_2_330 = {{6{_T_62396[4]}},_T_62396}; // @[Modules.scala 32:22:@8.4]
  assign _T_63231 = $signed(buffer_2_330) + $signed(buffer_1_331); // @[Modules.scala 50:57:@10452.4]
  assign _T_63232 = _T_63231[10:0]; // @[Modules.scala 50:57:@10453.4]
  assign buffer_2_557 = $signed(_T_63232); // @[Modules.scala 50:57:@10454.4]
  assign buffer_2_335 = {{6{_T_62415[4]}},_T_62415}; // @[Modules.scala 32:22:@8.4]
  assign _T_63237 = $signed(buffer_1_334) + $signed(buffer_2_335); // @[Modules.scala 50:57:@10460.4]
  assign _T_63238 = _T_63237[10:0]; // @[Modules.scala 50:57:@10461.4]
  assign buffer_2_559 = $signed(_T_63238); // @[Modules.scala 50:57:@10462.4]
  assign _T_63240 = $signed(buffer_1_336) + $signed(buffer_0_337); // @[Modules.scala 50:57:@10464.4]
  assign _T_63241 = _T_63240[10:0]; // @[Modules.scala 50:57:@10465.4]
  assign buffer_2_560 = $signed(_T_63241); // @[Modules.scala 50:57:@10466.4]
  assign buffer_2_338 = {{6{_T_62432[4]}},_T_62432}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_339 = {{6{_T_62439[4]}},_T_62439}; // @[Modules.scala 32:22:@8.4]
  assign _T_63243 = $signed(buffer_2_338) + $signed(buffer_2_339); // @[Modules.scala 50:57:@10468.4]
  assign _T_63244 = _T_63243[10:0]; // @[Modules.scala 50:57:@10469.4]
  assign buffer_2_561 = $signed(_T_63244); // @[Modules.scala 50:57:@10470.4]
  assign buffer_2_340 = {{6{_T_62446[4]}},_T_62446}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_341 = {{6{_T_62453[4]}},_T_62453}; // @[Modules.scala 32:22:@8.4]
  assign _T_63246 = $signed(buffer_2_340) + $signed(buffer_2_341); // @[Modules.scala 50:57:@10472.4]
  assign _T_63247 = _T_63246[10:0]; // @[Modules.scala 50:57:@10473.4]
  assign buffer_2_562 = $signed(_T_63247); // @[Modules.scala 50:57:@10474.4]
  assign buffer_2_342 = {{6{_T_62456[4]}},_T_62456}; // @[Modules.scala 32:22:@8.4]
  assign _T_63249 = $signed(buffer_2_342) + $signed(buffer_0_343); // @[Modules.scala 50:57:@10476.4]
  assign _T_63250 = _T_63249[10:0]; // @[Modules.scala 50:57:@10477.4]
  assign buffer_2_563 = $signed(_T_63250); // @[Modules.scala 50:57:@10478.4]
  assign buffer_2_344 = {{6{_T_62470[4]}},_T_62470}; // @[Modules.scala 32:22:@8.4]
  assign _T_63252 = $signed(buffer_2_344) + $signed(buffer_0_345); // @[Modules.scala 50:57:@10480.4]
  assign _T_63253 = _T_63252[10:0]; // @[Modules.scala 50:57:@10481.4]
  assign buffer_2_564 = $signed(_T_63253); // @[Modules.scala 50:57:@10482.4]
  assign buffer_2_348 = {{6{_T_62486[4]}},_T_62486}; // @[Modules.scala 32:22:@8.4]
  assign _T_63258 = $signed(buffer_2_348) + $signed(buffer_0_349); // @[Modules.scala 50:57:@10488.4]
  assign _T_63259 = _T_63258[10:0]; // @[Modules.scala 50:57:@10489.4]
  assign buffer_2_566 = $signed(_T_63259); // @[Modules.scala 50:57:@10490.4]
  assign buffer_2_350 = {{6{_T_62500[4]}},_T_62500}; // @[Modules.scala 32:22:@8.4]
  assign _T_63261 = $signed(buffer_2_350) + $signed(buffer_0_351); // @[Modules.scala 50:57:@10492.4]
  assign _T_63262 = _T_63261[10:0]; // @[Modules.scala 50:57:@10493.4]
  assign buffer_2_567 = $signed(_T_63262); // @[Modules.scala 50:57:@10494.4]
  assign buffer_2_352 = {{6{_T_62510[4]}},_T_62510}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_353 = {{6{_T_62517[4]}},_T_62517}; // @[Modules.scala 32:22:@8.4]
  assign _T_63264 = $signed(buffer_2_352) + $signed(buffer_2_353); // @[Modules.scala 50:57:@10496.4]
  assign _T_63265 = _T_63264[10:0]; // @[Modules.scala 50:57:@10497.4]
  assign buffer_2_568 = $signed(_T_63265); // @[Modules.scala 50:57:@10498.4]
  assign buffer_2_355 = {{6{_T_62531[4]}},_T_62531}; // @[Modules.scala 32:22:@8.4]
  assign _T_63267 = $signed(buffer_1_354) + $signed(buffer_2_355); // @[Modules.scala 50:57:@10500.4]
  assign _T_63268 = _T_63267[10:0]; // @[Modules.scala 50:57:@10501.4]
  assign buffer_2_569 = $signed(_T_63268); // @[Modules.scala 50:57:@10502.4]
  assign buffer_2_357 = {{6{_T_62545[4]}},_T_62545}; // @[Modules.scala 32:22:@8.4]
  assign _T_63270 = $signed(buffer_1_356) + $signed(buffer_2_357); // @[Modules.scala 50:57:@10504.4]
  assign _T_63271 = _T_63270[10:0]; // @[Modules.scala 50:57:@10505.4]
  assign buffer_2_570 = $signed(_T_63271); // @[Modules.scala 50:57:@10506.4]
  assign buffer_2_358 = {{6{_T_62552[4]}},_T_62552}; // @[Modules.scala 32:22:@8.4]
  assign _T_63273 = $signed(buffer_2_358) + $signed(buffer_1_359); // @[Modules.scala 50:57:@10508.4]
  assign _T_63274 = _T_63273[10:0]; // @[Modules.scala 50:57:@10509.4]
  assign buffer_2_571 = $signed(_T_63274); // @[Modules.scala 50:57:@10510.4]
  assign buffer_2_364 = {{6{_T_62578[4]}},_T_62578}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_365 = {{6{_T_62581[4]}},_T_62581}; // @[Modules.scala 32:22:@8.4]
  assign _T_63282 = $signed(buffer_2_364) + $signed(buffer_2_365); // @[Modules.scala 50:57:@10520.4]
  assign _T_63283 = _T_63282[10:0]; // @[Modules.scala 50:57:@10521.4]
  assign buffer_2_574 = $signed(_T_63283); // @[Modules.scala 50:57:@10522.4]
  assign buffer_2_366 = {{6{_T_62584[4]}},_T_62584}; // @[Modules.scala 32:22:@8.4]
  assign _T_63285 = $signed(buffer_2_366) + $signed(buffer_1_367); // @[Modules.scala 50:57:@10524.4]
  assign _T_63286 = _T_63285[10:0]; // @[Modules.scala 50:57:@10525.4]
  assign buffer_2_575 = $signed(_T_63286); // @[Modules.scala 50:57:@10526.4]
  assign buffer_2_374 = {{6{_T_62636[4]}},_T_62636}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_375 = {{6{_T_62643[4]}},_T_62643}; // @[Modules.scala 32:22:@8.4]
  assign _T_63297 = $signed(buffer_2_374) + $signed(buffer_2_375); // @[Modules.scala 50:57:@10540.4]
  assign _T_63298 = _T_63297[10:0]; // @[Modules.scala 50:57:@10541.4]
  assign buffer_2_579 = $signed(_T_63298); // @[Modules.scala 50:57:@10542.4]
  assign buffer_2_377 = {{6{_T_62649[4]}},_T_62649}; // @[Modules.scala 32:22:@8.4]
  assign _T_63300 = $signed(buffer_0_376) + $signed(buffer_2_377); // @[Modules.scala 50:57:@10544.4]
  assign _T_63301 = _T_63300[10:0]; // @[Modules.scala 50:57:@10545.4]
  assign buffer_2_580 = $signed(_T_63301); // @[Modules.scala 50:57:@10546.4]
  assign buffer_2_378 = {{6{_T_62656[4]}},_T_62656}; // @[Modules.scala 32:22:@8.4]
  assign _T_63303 = $signed(buffer_2_378) + $signed(buffer_1_379); // @[Modules.scala 50:57:@10548.4]
  assign _T_63304 = _T_63303[10:0]; // @[Modules.scala 50:57:@10549.4]
  assign buffer_2_581 = $signed(_T_63304); // @[Modules.scala 50:57:@10550.4]
  assign buffer_2_391 = {{6{_T_62735[4]}},_T_62735}; // @[Modules.scala 32:22:@8.4]
  assign _T_63321 = $signed(buffer_1_390) + $signed(buffer_2_391); // @[Modules.scala 50:57:@10572.4]
  assign _T_63322 = _T_63321[10:0]; // @[Modules.scala 50:57:@10573.4]
  assign buffer_2_587 = $signed(_T_63322); // @[Modules.scala 50:57:@10574.4]
  assign _T_63324 = $signed(buffer_0_392) + $signed(buffer_2_393); // @[Modules.scala 53:83:@10576.4]
  assign _T_63325 = _T_63324[10:0]; // @[Modules.scala 53:83:@10577.4]
  assign buffer_2_588 = $signed(_T_63325); // @[Modules.scala 53:83:@10578.4]
  assign _T_63327 = $signed(buffer_2_394) + $signed(buffer_0_395); // @[Modules.scala 53:83:@10580.4]
  assign _T_63328 = _T_63327[10:0]; // @[Modules.scala 53:83:@10581.4]
  assign buffer_2_589 = $signed(_T_63328); // @[Modules.scala 53:83:@10582.4]
  assign _T_63330 = $signed(buffer_2_396) + $signed(buffer_2_397); // @[Modules.scala 53:83:@10584.4]
  assign _T_63331 = _T_63330[10:0]; // @[Modules.scala 53:83:@10585.4]
  assign buffer_2_590 = $signed(_T_63331); // @[Modules.scala 53:83:@10586.4]
  assign _T_63333 = $signed(buffer_2_398) + $signed(buffer_2_399); // @[Modules.scala 53:83:@10588.4]
  assign _T_63334 = _T_63333[10:0]; // @[Modules.scala 53:83:@10589.4]
  assign buffer_2_591 = $signed(_T_63334); // @[Modules.scala 53:83:@10590.4]
  assign _T_63336 = $signed(buffer_2_400) + $signed(buffer_1_401); // @[Modules.scala 53:83:@10592.4]
  assign _T_63337 = _T_63336[10:0]; // @[Modules.scala 53:83:@10593.4]
  assign buffer_2_592 = $signed(_T_63337); // @[Modules.scala 53:83:@10594.4]
  assign _T_63339 = $signed(buffer_2_402) + $signed(buffer_2_403); // @[Modules.scala 53:83:@10596.4]
  assign _T_63340 = _T_63339[10:0]; // @[Modules.scala 53:83:@10597.4]
  assign buffer_2_593 = $signed(_T_63340); // @[Modules.scala 53:83:@10598.4]
  assign _T_63342 = $signed(buffer_1_404) + $signed(buffer_2_405); // @[Modules.scala 53:83:@10600.4]
  assign _T_63343 = _T_63342[10:0]; // @[Modules.scala 53:83:@10601.4]
  assign buffer_2_594 = $signed(_T_63343); // @[Modules.scala 53:83:@10602.4]
  assign _T_63345 = $signed(buffer_2_406) + $signed(buffer_2_407); // @[Modules.scala 53:83:@10604.4]
  assign _T_63346 = _T_63345[10:0]; // @[Modules.scala 53:83:@10605.4]
  assign buffer_2_595 = $signed(_T_63346); // @[Modules.scala 53:83:@10606.4]
  assign _T_63348 = $signed(buffer_1_408) + $signed(buffer_2_409); // @[Modules.scala 53:83:@10608.4]
  assign _T_63349 = _T_63348[10:0]; // @[Modules.scala 53:83:@10609.4]
  assign buffer_2_596 = $signed(_T_63349); // @[Modules.scala 53:83:@10610.4]
  assign _T_63351 = $signed(buffer_1_410) + $signed(buffer_2_411); // @[Modules.scala 53:83:@10612.4]
  assign _T_63352 = _T_63351[10:0]; // @[Modules.scala 53:83:@10613.4]
  assign buffer_2_597 = $signed(_T_63352); // @[Modules.scala 53:83:@10614.4]
  assign _T_63354 = $signed(buffer_2_412) + $signed(buffer_2_413); // @[Modules.scala 53:83:@10616.4]
  assign _T_63355 = _T_63354[10:0]; // @[Modules.scala 53:83:@10617.4]
  assign buffer_2_598 = $signed(_T_63355); // @[Modules.scala 53:83:@10618.4]
  assign _T_63357 = $signed(buffer_2_414) + $signed(buffer_2_415); // @[Modules.scala 53:83:@10620.4]
  assign _T_63358 = _T_63357[10:0]; // @[Modules.scala 53:83:@10621.4]
  assign buffer_2_599 = $signed(_T_63358); // @[Modules.scala 53:83:@10622.4]
  assign _T_63360 = $signed(buffer_2_416) + $signed(buffer_2_417); // @[Modules.scala 53:83:@10624.4]
  assign _T_63361 = _T_63360[10:0]; // @[Modules.scala 53:83:@10625.4]
  assign buffer_2_600 = $signed(_T_63361); // @[Modules.scala 53:83:@10626.4]
  assign _T_63363 = $signed(buffer_0_418) + $signed(buffer_2_419); // @[Modules.scala 53:83:@10628.4]
  assign _T_63364 = _T_63363[10:0]; // @[Modules.scala 53:83:@10629.4]
  assign buffer_2_601 = $signed(_T_63364); // @[Modules.scala 53:83:@10630.4]
  assign _T_63366 = $signed(buffer_0_420) + $signed(buffer_2_421); // @[Modules.scala 53:83:@10632.4]
  assign _T_63367 = _T_63366[10:0]; // @[Modules.scala 53:83:@10633.4]
  assign buffer_2_602 = $signed(_T_63367); // @[Modules.scala 53:83:@10634.4]
  assign _T_63372 = $signed(buffer_2_424) + $signed(buffer_1_425); // @[Modules.scala 53:83:@10640.4]
  assign _T_63373 = _T_63372[10:0]; // @[Modules.scala 53:83:@10641.4]
  assign buffer_2_604 = $signed(_T_63373); // @[Modules.scala 53:83:@10642.4]
  assign _T_63375 = $signed(buffer_0_426) + $signed(buffer_2_427); // @[Modules.scala 53:83:@10644.4]
  assign _T_63376 = _T_63375[10:0]; // @[Modules.scala 53:83:@10645.4]
  assign buffer_2_605 = $signed(_T_63376); // @[Modules.scala 53:83:@10646.4]
  assign _T_63378 = $signed(buffer_1_428) + $signed(buffer_2_429); // @[Modules.scala 53:83:@10648.4]
  assign _T_63379 = _T_63378[10:0]; // @[Modules.scala 53:83:@10649.4]
  assign buffer_2_606 = $signed(_T_63379); // @[Modules.scala 53:83:@10650.4]
  assign _T_63381 = $signed(buffer_0_430) + $signed(buffer_2_431); // @[Modules.scala 53:83:@10652.4]
  assign _T_63382 = _T_63381[10:0]; // @[Modules.scala 53:83:@10653.4]
  assign buffer_2_607 = $signed(_T_63382); // @[Modules.scala 53:83:@10654.4]
  assign _T_63384 = $signed(buffer_2_432) + $signed(buffer_2_433); // @[Modules.scala 53:83:@10656.4]
  assign _T_63385 = _T_63384[10:0]; // @[Modules.scala 53:83:@10657.4]
  assign buffer_2_608 = $signed(_T_63385); // @[Modules.scala 53:83:@10658.4]
  assign _T_63387 = $signed(buffer_2_434) + $signed(buffer_2_435); // @[Modules.scala 53:83:@10660.4]
  assign _T_63388 = _T_63387[10:0]; // @[Modules.scala 53:83:@10661.4]
  assign buffer_2_609 = $signed(_T_63388); // @[Modules.scala 53:83:@10662.4]
  assign _T_63393 = $signed(buffer_2_438) + $signed(buffer_2_439); // @[Modules.scala 53:83:@10668.4]
  assign _T_63394 = _T_63393[10:0]; // @[Modules.scala 53:83:@10669.4]
  assign buffer_2_611 = $signed(_T_63394); // @[Modules.scala 53:83:@10670.4]
  assign _T_63396 = $signed(buffer_2_440) + $signed(buffer_2_441); // @[Modules.scala 53:83:@10672.4]
  assign _T_63397 = _T_63396[10:0]; // @[Modules.scala 53:83:@10673.4]
  assign buffer_2_612 = $signed(_T_63397); // @[Modules.scala 53:83:@10674.4]
  assign _T_63399 = $signed(buffer_0_442) + $signed(buffer_2_443); // @[Modules.scala 53:83:@10676.4]
  assign _T_63400 = _T_63399[10:0]; // @[Modules.scala 53:83:@10677.4]
  assign buffer_2_613 = $signed(_T_63400); // @[Modules.scala 53:83:@10678.4]
  assign _T_63402 = $signed(buffer_2_444) + $signed(buffer_2_445); // @[Modules.scala 53:83:@10680.4]
  assign _T_63403 = _T_63402[10:0]; // @[Modules.scala 53:83:@10681.4]
  assign buffer_2_614 = $signed(_T_63403); // @[Modules.scala 53:83:@10682.4]
  assign _T_63405 = $signed(buffer_2_446) + $signed(buffer_2_447); // @[Modules.scala 53:83:@10684.4]
  assign _T_63406 = _T_63405[10:0]; // @[Modules.scala 53:83:@10685.4]
  assign buffer_2_615 = $signed(_T_63406); // @[Modules.scala 53:83:@10686.4]
  assign _T_63411 = $signed(buffer_2_450) + $signed(buffer_1_451); // @[Modules.scala 53:83:@10692.4]
  assign _T_63412 = _T_63411[10:0]; // @[Modules.scala 53:83:@10693.4]
  assign buffer_2_617 = $signed(_T_63412); // @[Modules.scala 53:83:@10694.4]
  assign _T_63414 = $signed(buffer_0_452) + $signed(buffer_1_453); // @[Modules.scala 53:83:@10696.4]
  assign _T_63415 = _T_63414[10:0]; // @[Modules.scala 53:83:@10697.4]
  assign buffer_2_618 = $signed(_T_63415); // @[Modules.scala 53:83:@10698.4]
  assign _T_63417 = $signed(buffer_1_454) + $signed(buffer_0_455); // @[Modules.scala 53:83:@10700.4]
  assign _T_63418 = _T_63417[10:0]; // @[Modules.scala 53:83:@10701.4]
  assign buffer_2_619 = $signed(_T_63418); // @[Modules.scala 53:83:@10702.4]
  assign _T_63420 = $signed(buffer_0_456) + $signed(buffer_2_457); // @[Modules.scala 53:83:@10704.4]
  assign _T_63421 = _T_63420[10:0]; // @[Modules.scala 53:83:@10705.4]
  assign buffer_2_620 = $signed(_T_63421); // @[Modules.scala 53:83:@10706.4]
  assign _T_63426 = $signed(buffer_0_460) + $signed(buffer_1_461); // @[Modules.scala 53:83:@10712.4]
  assign _T_63427 = _T_63426[10:0]; // @[Modules.scala 53:83:@10713.4]
  assign buffer_2_622 = $signed(_T_63427); // @[Modules.scala 53:83:@10714.4]
  assign _T_63429 = $signed(buffer_0_462) + $signed(buffer_2_463); // @[Modules.scala 53:83:@10716.4]
  assign _T_63430 = _T_63429[10:0]; // @[Modules.scala 53:83:@10717.4]
  assign buffer_2_623 = $signed(_T_63430); // @[Modules.scala 53:83:@10718.4]
  assign _T_63432 = $signed(buffer_2_464) + $signed(buffer_0_465); // @[Modules.scala 53:83:@10720.4]
  assign _T_63433 = _T_63432[10:0]; // @[Modules.scala 53:83:@10721.4]
  assign buffer_2_624 = $signed(_T_63433); // @[Modules.scala 53:83:@10722.4]
  assign _T_63438 = $signed(buffer_2_468) + $signed(buffer_0_469); // @[Modules.scala 53:83:@10728.4]
  assign _T_63439 = _T_63438[10:0]; // @[Modules.scala 53:83:@10729.4]
  assign buffer_2_626 = $signed(_T_63439); // @[Modules.scala 53:83:@10730.4]
  assign _T_63441 = $signed(buffer_2_470) + $signed(buffer_0_471); // @[Modules.scala 53:83:@10732.4]
  assign _T_63442 = _T_63441[10:0]; // @[Modules.scala 53:83:@10733.4]
  assign buffer_2_627 = $signed(_T_63442); // @[Modules.scala 53:83:@10734.4]
  assign _T_63444 = $signed(buffer_2_472) + $signed(buffer_1_473); // @[Modules.scala 53:83:@10736.4]
  assign _T_63445 = _T_63444[10:0]; // @[Modules.scala 53:83:@10737.4]
  assign buffer_2_628 = $signed(_T_63445); // @[Modules.scala 53:83:@10738.4]
  assign _T_63447 = $signed(buffer_2_474) + $signed(buffer_2_475); // @[Modules.scala 53:83:@10740.4]
  assign _T_63448 = _T_63447[10:0]; // @[Modules.scala 53:83:@10741.4]
  assign buffer_2_629 = $signed(_T_63448); // @[Modules.scala 53:83:@10742.4]
  assign _T_63456 = $signed(buffer_2_480) + $signed(buffer_2_481); // @[Modules.scala 53:83:@10752.4]
  assign _T_63457 = _T_63456[10:0]; // @[Modules.scala 53:83:@10753.4]
  assign buffer_2_632 = $signed(_T_63457); // @[Modules.scala 53:83:@10754.4]
  assign _T_63459 = $signed(buffer_2_482) + $signed(buffer_0_483); // @[Modules.scala 53:83:@10756.4]
  assign _T_63460 = _T_63459[10:0]; // @[Modules.scala 53:83:@10757.4]
  assign buffer_2_633 = $signed(_T_63460); // @[Modules.scala 53:83:@10758.4]
  assign _T_63468 = $signed(buffer_2_488) + $signed(buffer_2_489); // @[Modules.scala 53:83:@10768.4]
  assign _T_63469 = _T_63468[10:0]; // @[Modules.scala 53:83:@10769.4]
  assign buffer_2_636 = $signed(_T_63469); // @[Modules.scala 53:83:@10770.4]
  assign _T_63471 = $signed(buffer_1_490) + $signed(buffer_0_491); // @[Modules.scala 53:83:@10772.4]
  assign _T_63472 = _T_63471[10:0]; // @[Modules.scala 53:83:@10773.4]
  assign buffer_2_637 = $signed(_T_63472); // @[Modules.scala 53:83:@10774.4]
  assign _T_63477 = $signed(buffer_2_494) + $signed(buffer_0_495); // @[Modules.scala 53:83:@10780.4]
  assign _T_63478 = _T_63477[10:0]; // @[Modules.scala 53:83:@10781.4]
  assign buffer_2_639 = $signed(_T_63478); // @[Modules.scala 53:83:@10782.4]
  assign _T_63480 = $signed(buffer_2_496) + $signed(buffer_2_497); // @[Modules.scala 53:83:@10784.4]
  assign _T_63481 = _T_63480[10:0]; // @[Modules.scala 53:83:@10785.4]
  assign buffer_2_640 = $signed(_T_63481); // @[Modules.scala 53:83:@10786.4]
  assign _T_63483 = $signed(buffer_2_498) + $signed(buffer_2_499); // @[Modules.scala 53:83:@10788.4]
  assign _T_63484 = _T_63483[10:0]; // @[Modules.scala 53:83:@10789.4]
  assign buffer_2_641 = $signed(_T_63484); // @[Modules.scala 53:83:@10790.4]
  assign _T_63486 = $signed(buffer_0_500) + $signed(buffer_2_501); // @[Modules.scala 53:83:@10792.4]
  assign _T_63487 = _T_63486[10:0]; // @[Modules.scala 53:83:@10793.4]
  assign buffer_2_642 = $signed(_T_63487); // @[Modules.scala 53:83:@10794.4]
  assign _T_63489 = $signed(buffer_2_502) + $signed(buffer_0_503); // @[Modules.scala 53:83:@10796.4]
  assign _T_63490 = _T_63489[10:0]; // @[Modules.scala 53:83:@10797.4]
  assign buffer_2_643 = $signed(_T_63490); // @[Modules.scala 53:83:@10798.4]
  assign _T_63492 = $signed(buffer_2_504) + $signed(buffer_2_505); // @[Modules.scala 53:83:@10800.4]
  assign _T_63493 = _T_63492[10:0]; // @[Modules.scala 53:83:@10801.4]
  assign buffer_2_644 = $signed(_T_63493); // @[Modules.scala 53:83:@10802.4]
  assign _T_63495 = $signed(buffer_2_506) + $signed(buffer_2_507); // @[Modules.scala 53:83:@10804.4]
  assign _T_63496 = _T_63495[10:0]; // @[Modules.scala 53:83:@10805.4]
  assign buffer_2_645 = $signed(_T_63496); // @[Modules.scala 53:83:@10806.4]
  assign _T_63498 = $signed(buffer_2_508) + $signed(buffer_2_509); // @[Modules.scala 53:83:@10808.4]
  assign _T_63499 = _T_63498[10:0]; // @[Modules.scala 53:83:@10809.4]
  assign buffer_2_646 = $signed(_T_63499); // @[Modules.scala 53:83:@10810.4]
  assign _T_63501 = $signed(buffer_0_510) + $signed(buffer_2_511); // @[Modules.scala 53:83:@10812.4]
  assign _T_63502 = _T_63501[10:0]; // @[Modules.scala 53:83:@10813.4]
  assign buffer_2_647 = $signed(_T_63502); // @[Modules.scala 53:83:@10814.4]
  assign _T_63504 = $signed(buffer_2_512) + $signed(buffer_2_513); // @[Modules.scala 53:83:@10816.4]
  assign _T_63505 = _T_63504[10:0]; // @[Modules.scala 53:83:@10817.4]
  assign buffer_2_648 = $signed(_T_63505); // @[Modules.scala 53:83:@10818.4]
  assign _T_63507 = $signed(buffer_2_514) + $signed(buffer_1_515); // @[Modules.scala 53:83:@10820.4]
  assign _T_63508 = _T_63507[10:0]; // @[Modules.scala 53:83:@10821.4]
  assign buffer_2_649 = $signed(_T_63508); // @[Modules.scala 53:83:@10822.4]
  assign _T_63510 = $signed(buffer_2_516) + $signed(buffer_0_517); // @[Modules.scala 53:83:@10824.4]
  assign _T_63511 = _T_63510[10:0]; // @[Modules.scala 53:83:@10825.4]
  assign buffer_2_650 = $signed(_T_63511); // @[Modules.scala 53:83:@10826.4]
  assign _T_63513 = $signed(buffer_2_518) + $signed(buffer_0_519); // @[Modules.scala 53:83:@10828.4]
  assign _T_63514 = _T_63513[10:0]; // @[Modules.scala 53:83:@10829.4]
  assign buffer_2_651 = $signed(_T_63514); // @[Modules.scala 53:83:@10830.4]
  assign _T_63516 = $signed(buffer_1_520) + $signed(buffer_2_521); // @[Modules.scala 53:83:@10832.4]
  assign _T_63517 = _T_63516[10:0]; // @[Modules.scala 53:83:@10833.4]
  assign buffer_2_652 = $signed(_T_63517); // @[Modules.scala 53:83:@10834.4]
  assign _T_63519 = $signed(buffer_2_522) + $signed(buffer_2_523); // @[Modules.scala 53:83:@10836.4]
  assign _T_63520 = _T_63519[10:0]; // @[Modules.scala 53:83:@10837.4]
  assign buffer_2_653 = $signed(_T_63520); // @[Modules.scala 53:83:@10838.4]
  assign _T_63522 = $signed(buffer_1_524) + $signed(buffer_2_525); // @[Modules.scala 53:83:@10840.4]
  assign _T_63523 = _T_63522[10:0]; // @[Modules.scala 53:83:@10841.4]
  assign buffer_2_654 = $signed(_T_63523); // @[Modules.scala 53:83:@10842.4]
  assign _T_63528 = $signed(buffer_2_528) + $signed(buffer_2_529); // @[Modules.scala 53:83:@10848.4]
  assign _T_63529 = _T_63528[10:0]; // @[Modules.scala 53:83:@10849.4]
  assign buffer_2_656 = $signed(_T_63529); // @[Modules.scala 53:83:@10850.4]
  assign _T_63531 = $signed(buffer_2_530) + $signed(buffer_2_531); // @[Modules.scala 53:83:@10852.4]
  assign _T_63532 = _T_63531[10:0]; // @[Modules.scala 53:83:@10853.4]
  assign buffer_2_657 = $signed(_T_63532); // @[Modules.scala 53:83:@10854.4]
  assign _T_63534 = $signed(buffer_2_532) + $signed(buffer_0_533); // @[Modules.scala 53:83:@10856.4]
  assign _T_63535 = _T_63534[10:0]; // @[Modules.scala 53:83:@10857.4]
  assign buffer_2_658 = $signed(_T_63535); // @[Modules.scala 53:83:@10858.4]
  assign _T_63537 = $signed(buffer_0_534) + $signed(buffer_2_535); // @[Modules.scala 53:83:@10860.4]
  assign _T_63538 = _T_63537[10:0]; // @[Modules.scala 53:83:@10861.4]
  assign buffer_2_659 = $signed(_T_63538); // @[Modules.scala 53:83:@10862.4]
  assign _T_63540 = $signed(buffer_2_536) + $signed(buffer_2_537); // @[Modules.scala 53:83:@10864.4]
  assign _T_63541 = _T_63540[10:0]; // @[Modules.scala 53:83:@10865.4]
  assign buffer_2_660 = $signed(_T_63541); // @[Modules.scala 53:83:@10866.4]
  assign _T_63543 = $signed(buffer_1_538) + $signed(buffer_2_539); // @[Modules.scala 53:83:@10868.4]
  assign _T_63544 = _T_63543[10:0]; // @[Modules.scala 53:83:@10869.4]
  assign buffer_2_661 = $signed(_T_63544); // @[Modules.scala 53:83:@10870.4]
  assign _T_63546 = $signed(buffer_2_540) + $signed(buffer_2_541); // @[Modules.scala 53:83:@10872.4]
  assign _T_63547 = _T_63546[10:0]; // @[Modules.scala 53:83:@10873.4]
  assign buffer_2_662 = $signed(_T_63547); // @[Modules.scala 53:83:@10874.4]
  assign _T_63549 = $signed(buffer_2_542) + $signed(buffer_2_543); // @[Modules.scala 53:83:@10876.4]
  assign _T_63550 = _T_63549[10:0]; // @[Modules.scala 53:83:@10877.4]
  assign buffer_2_663 = $signed(_T_63550); // @[Modules.scala 53:83:@10878.4]
  assign _T_63552 = $signed(buffer_2_544) + $signed(buffer_1_545); // @[Modules.scala 53:83:@10880.4]
  assign _T_63553 = _T_63552[10:0]; // @[Modules.scala 53:83:@10881.4]
  assign buffer_2_664 = $signed(_T_63553); // @[Modules.scala 53:83:@10882.4]
  assign _T_63555 = $signed(buffer_2_546) + $signed(buffer_0_547); // @[Modules.scala 53:83:@10884.4]
  assign _T_63556 = _T_63555[10:0]; // @[Modules.scala 53:83:@10885.4]
  assign buffer_2_665 = $signed(_T_63556); // @[Modules.scala 53:83:@10886.4]
  assign _T_63558 = $signed(buffer_2_548) + $signed(buffer_0_549); // @[Modules.scala 53:83:@10888.4]
  assign _T_63559 = _T_63558[10:0]; // @[Modules.scala 53:83:@10889.4]
  assign buffer_2_666 = $signed(_T_63559); // @[Modules.scala 53:83:@10890.4]
  assign _T_63561 = $signed(buffer_2_550) + $signed(buffer_1_551); // @[Modules.scala 53:83:@10892.4]
  assign _T_63562 = _T_63561[10:0]; // @[Modules.scala 53:83:@10893.4]
  assign buffer_2_667 = $signed(_T_63562); // @[Modules.scala 53:83:@10894.4]
  assign _T_63564 = $signed(buffer_1_552) + $signed(buffer_2_553); // @[Modules.scala 53:83:@10896.4]
  assign _T_63565 = _T_63564[10:0]; // @[Modules.scala 53:83:@10897.4]
  assign buffer_2_668 = $signed(_T_63565); // @[Modules.scala 53:83:@10898.4]
  assign _T_63567 = $signed(buffer_2_554) + $signed(buffer_2_555); // @[Modules.scala 53:83:@10900.4]
  assign _T_63568 = _T_63567[10:0]; // @[Modules.scala 53:83:@10901.4]
  assign buffer_2_669 = $signed(_T_63568); // @[Modules.scala 53:83:@10902.4]
  assign _T_63570 = $signed(buffer_2_556) + $signed(buffer_2_557); // @[Modules.scala 53:83:@10904.4]
  assign _T_63571 = _T_63570[10:0]; // @[Modules.scala 53:83:@10905.4]
  assign buffer_2_670 = $signed(_T_63571); // @[Modules.scala 53:83:@10906.4]
  assign _T_63573 = $signed(buffer_0_558) + $signed(buffer_2_559); // @[Modules.scala 53:83:@10908.4]
  assign _T_63574 = _T_63573[10:0]; // @[Modules.scala 53:83:@10909.4]
  assign buffer_2_671 = $signed(_T_63574); // @[Modules.scala 53:83:@10910.4]
  assign _T_63576 = $signed(buffer_2_560) + $signed(buffer_2_561); // @[Modules.scala 53:83:@10912.4]
  assign _T_63577 = _T_63576[10:0]; // @[Modules.scala 53:83:@10913.4]
  assign buffer_2_672 = $signed(_T_63577); // @[Modules.scala 53:83:@10914.4]
  assign _T_63579 = $signed(buffer_2_562) + $signed(buffer_2_563); // @[Modules.scala 53:83:@10916.4]
  assign _T_63580 = _T_63579[10:0]; // @[Modules.scala 53:83:@10917.4]
  assign buffer_2_673 = $signed(_T_63580); // @[Modules.scala 53:83:@10918.4]
  assign _T_63582 = $signed(buffer_2_564) + $signed(buffer_0_565); // @[Modules.scala 53:83:@10920.4]
  assign _T_63583 = _T_63582[10:0]; // @[Modules.scala 53:83:@10921.4]
  assign buffer_2_674 = $signed(_T_63583); // @[Modules.scala 53:83:@10922.4]
  assign _T_63585 = $signed(buffer_2_566) + $signed(buffer_2_567); // @[Modules.scala 53:83:@10924.4]
  assign _T_63586 = _T_63585[10:0]; // @[Modules.scala 53:83:@10925.4]
  assign buffer_2_675 = $signed(_T_63586); // @[Modules.scala 53:83:@10926.4]
  assign _T_63588 = $signed(buffer_2_568) + $signed(buffer_2_569); // @[Modules.scala 53:83:@10928.4]
  assign _T_63589 = _T_63588[10:0]; // @[Modules.scala 53:83:@10929.4]
  assign buffer_2_676 = $signed(_T_63589); // @[Modules.scala 53:83:@10930.4]
  assign _T_63591 = $signed(buffer_2_570) + $signed(buffer_2_571); // @[Modules.scala 53:83:@10932.4]
  assign _T_63592 = _T_63591[10:0]; // @[Modules.scala 53:83:@10933.4]
  assign buffer_2_677 = $signed(_T_63592); // @[Modules.scala 53:83:@10934.4]
  assign _T_63597 = $signed(buffer_2_574) + $signed(buffer_2_575); // @[Modules.scala 53:83:@10940.4]
  assign _T_63598 = _T_63597[10:0]; // @[Modules.scala 53:83:@10941.4]
  assign buffer_2_679 = $signed(_T_63598); // @[Modules.scala 53:83:@10942.4]
  assign _T_63603 = $signed(buffer_0_578) + $signed(buffer_2_579); // @[Modules.scala 53:83:@10948.4]
  assign _T_63604 = _T_63603[10:0]; // @[Modules.scala 53:83:@10949.4]
  assign buffer_2_681 = $signed(_T_63604); // @[Modules.scala 53:83:@10950.4]
  assign _T_63606 = $signed(buffer_2_580) + $signed(buffer_2_581); // @[Modules.scala 53:83:@10952.4]
  assign _T_63607 = _T_63606[10:0]; // @[Modules.scala 53:83:@10953.4]
  assign buffer_2_682 = $signed(_T_63607); // @[Modules.scala 53:83:@10954.4]
  assign _T_63615 = $signed(buffer_1_586) + $signed(buffer_2_587); // @[Modules.scala 53:83:@10964.4]
  assign _T_63616 = _T_63615[10:0]; // @[Modules.scala 53:83:@10965.4]
  assign buffer_2_685 = $signed(_T_63616); // @[Modules.scala 53:83:@10966.4]
  assign _T_63618 = $signed(buffer_2_588) + $signed(buffer_2_589); // @[Modules.scala 56:109:@10968.4]
  assign _T_63619 = _T_63618[10:0]; // @[Modules.scala 56:109:@10969.4]
  assign buffer_2_686 = $signed(_T_63619); // @[Modules.scala 56:109:@10970.4]
  assign _T_63621 = $signed(buffer_2_590) + $signed(buffer_2_591); // @[Modules.scala 56:109:@10972.4]
  assign _T_63622 = _T_63621[10:0]; // @[Modules.scala 56:109:@10973.4]
  assign buffer_2_687 = $signed(_T_63622); // @[Modules.scala 56:109:@10974.4]
  assign _T_63624 = $signed(buffer_2_592) + $signed(buffer_2_593); // @[Modules.scala 56:109:@10976.4]
  assign _T_63625 = _T_63624[10:0]; // @[Modules.scala 56:109:@10977.4]
  assign buffer_2_688 = $signed(_T_63625); // @[Modules.scala 56:109:@10978.4]
  assign _T_63627 = $signed(buffer_2_594) + $signed(buffer_2_595); // @[Modules.scala 56:109:@10980.4]
  assign _T_63628 = _T_63627[10:0]; // @[Modules.scala 56:109:@10981.4]
  assign buffer_2_689 = $signed(_T_63628); // @[Modules.scala 56:109:@10982.4]
  assign _T_63630 = $signed(buffer_2_596) + $signed(buffer_2_597); // @[Modules.scala 56:109:@10984.4]
  assign _T_63631 = _T_63630[10:0]; // @[Modules.scala 56:109:@10985.4]
  assign buffer_2_690 = $signed(_T_63631); // @[Modules.scala 56:109:@10986.4]
  assign _T_63633 = $signed(buffer_2_598) + $signed(buffer_2_599); // @[Modules.scala 56:109:@10988.4]
  assign _T_63634 = _T_63633[10:0]; // @[Modules.scala 56:109:@10989.4]
  assign buffer_2_691 = $signed(_T_63634); // @[Modules.scala 56:109:@10990.4]
  assign _T_63636 = $signed(buffer_2_600) + $signed(buffer_2_601); // @[Modules.scala 56:109:@10992.4]
  assign _T_63637 = _T_63636[10:0]; // @[Modules.scala 56:109:@10993.4]
  assign buffer_2_692 = $signed(_T_63637); // @[Modules.scala 56:109:@10994.4]
  assign _T_63639 = $signed(buffer_2_602) + $signed(buffer_0_603); // @[Modules.scala 56:109:@10996.4]
  assign _T_63640 = _T_63639[10:0]; // @[Modules.scala 56:109:@10997.4]
  assign buffer_2_693 = $signed(_T_63640); // @[Modules.scala 56:109:@10998.4]
  assign _T_63642 = $signed(buffer_2_604) + $signed(buffer_2_605); // @[Modules.scala 56:109:@11000.4]
  assign _T_63643 = _T_63642[10:0]; // @[Modules.scala 56:109:@11001.4]
  assign buffer_2_694 = $signed(_T_63643); // @[Modules.scala 56:109:@11002.4]
  assign _T_63645 = $signed(buffer_2_606) + $signed(buffer_2_607); // @[Modules.scala 56:109:@11004.4]
  assign _T_63646 = _T_63645[10:0]; // @[Modules.scala 56:109:@11005.4]
  assign buffer_2_695 = $signed(_T_63646); // @[Modules.scala 56:109:@11006.4]
  assign _T_63648 = $signed(buffer_2_608) + $signed(buffer_2_609); // @[Modules.scala 56:109:@11008.4]
  assign _T_63649 = _T_63648[10:0]; // @[Modules.scala 56:109:@11009.4]
  assign buffer_2_696 = $signed(_T_63649); // @[Modules.scala 56:109:@11010.4]
  assign _T_63651 = $signed(buffer_0_610) + $signed(buffer_2_611); // @[Modules.scala 56:109:@11012.4]
  assign _T_63652 = _T_63651[10:0]; // @[Modules.scala 56:109:@11013.4]
  assign buffer_2_697 = $signed(_T_63652); // @[Modules.scala 56:109:@11014.4]
  assign _T_63654 = $signed(buffer_2_612) + $signed(buffer_2_613); // @[Modules.scala 56:109:@11016.4]
  assign _T_63655 = _T_63654[10:0]; // @[Modules.scala 56:109:@11017.4]
  assign buffer_2_698 = $signed(_T_63655); // @[Modules.scala 56:109:@11018.4]
  assign _T_63657 = $signed(buffer_2_614) + $signed(buffer_2_615); // @[Modules.scala 56:109:@11020.4]
  assign _T_63658 = _T_63657[10:0]; // @[Modules.scala 56:109:@11021.4]
  assign buffer_2_699 = $signed(_T_63658); // @[Modules.scala 56:109:@11022.4]
  assign _T_63660 = $signed(buffer_0_616) + $signed(buffer_2_617); // @[Modules.scala 56:109:@11024.4]
  assign _T_63661 = _T_63660[10:0]; // @[Modules.scala 56:109:@11025.4]
  assign buffer_2_700 = $signed(_T_63661); // @[Modules.scala 56:109:@11026.4]
  assign _T_63663 = $signed(buffer_2_618) + $signed(buffer_2_619); // @[Modules.scala 56:109:@11028.4]
  assign _T_63664 = _T_63663[10:0]; // @[Modules.scala 56:109:@11029.4]
  assign buffer_2_701 = $signed(_T_63664); // @[Modules.scala 56:109:@11030.4]
  assign _T_63666 = $signed(buffer_2_620) + $signed(buffer_0_621); // @[Modules.scala 56:109:@11032.4]
  assign _T_63667 = _T_63666[10:0]; // @[Modules.scala 56:109:@11033.4]
  assign buffer_2_702 = $signed(_T_63667); // @[Modules.scala 56:109:@11034.4]
  assign _T_63669 = $signed(buffer_2_622) + $signed(buffer_2_623); // @[Modules.scala 56:109:@11036.4]
  assign _T_63670 = _T_63669[10:0]; // @[Modules.scala 56:109:@11037.4]
  assign buffer_2_703 = $signed(_T_63670); // @[Modules.scala 56:109:@11038.4]
  assign _T_63672 = $signed(buffer_2_624) + $signed(buffer_0_625); // @[Modules.scala 56:109:@11040.4]
  assign _T_63673 = _T_63672[10:0]; // @[Modules.scala 56:109:@11041.4]
  assign buffer_2_704 = $signed(_T_63673); // @[Modules.scala 56:109:@11042.4]
  assign _T_63675 = $signed(buffer_2_626) + $signed(buffer_2_627); // @[Modules.scala 56:109:@11044.4]
  assign _T_63676 = _T_63675[10:0]; // @[Modules.scala 56:109:@11045.4]
  assign buffer_2_705 = $signed(_T_63676); // @[Modules.scala 56:109:@11046.4]
  assign _T_63678 = $signed(buffer_2_628) + $signed(buffer_2_629); // @[Modules.scala 56:109:@11048.4]
  assign _T_63679 = _T_63678[10:0]; // @[Modules.scala 56:109:@11049.4]
  assign buffer_2_706 = $signed(_T_63679); // @[Modules.scala 56:109:@11050.4]
  assign _T_63684 = $signed(buffer_2_632) + $signed(buffer_2_633); // @[Modules.scala 56:109:@11056.4]
  assign _T_63685 = _T_63684[10:0]; // @[Modules.scala 56:109:@11057.4]
  assign buffer_2_708 = $signed(_T_63685); // @[Modules.scala 56:109:@11058.4]
  assign _T_63687 = $signed(buffer_1_634) + $signed(buffer_0_635); // @[Modules.scala 56:109:@11060.4]
  assign _T_63688 = _T_63687[10:0]; // @[Modules.scala 56:109:@11061.4]
  assign buffer_2_709 = $signed(_T_63688); // @[Modules.scala 56:109:@11062.4]
  assign _T_63690 = $signed(buffer_2_636) + $signed(buffer_2_637); // @[Modules.scala 56:109:@11064.4]
  assign _T_63691 = _T_63690[10:0]; // @[Modules.scala 56:109:@11065.4]
  assign buffer_2_710 = $signed(_T_63691); // @[Modules.scala 56:109:@11066.4]
  assign _T_63693 = $signed(buffer_0_638) + $signed(buffer_2_639); // @[Modules.scala 56:109:@11068.4]
  assign _T_63694 = _T_63693[10:0]; // @[Modules.scala 56:109:@11069.4]
  assign buffer_2_711 = $signed(_T_63694); // @[Modules.scala 56:109:@11070.4]
  assign _T_63696 = $signed(buffer_2_640) + $signed(buffer_2_641); // @[Modules.scala 56:109:@11072.4]
  assign _T_63697 = _T_63696[10:0]; // @[Modules.scala 56:109:@11073.4]
  assign buffer_2_712 = $signed(_T_63697); // @[Modules.scala 56:109:@11074.4]
  assign _T_63699 = $signed(buffer_2_642) + $signed(buffer_2_643); // @[Modules.scala 56:109:@11076.4]
  assign _T_63700 = _T_63699[10:0]; // @[Modules.scala 56:109:@11077.4]
  assign buffer_2_713 = $signed(_T_63700); // @[Modules.scala 56:109:@11078.4]
  assign _T_63702 = $signed(buffer_2_644) + $signed(buffer_2_645); // @[Modules.scala 56:109:@11080.4]
  assign _T_63703 = _T_63702[10:0]; // @[Modules.scala 56:109:@11081.4]
  assign buffer_2_714 = $signed(_T_63703); // @[Modules.scala 56:109:@11082.4]
  assign _T_63705 = $signed(buffer_2_646) + $signed(buffer_2_647); // @[Modules.scala 56:109:@11084.4]
  assign _T_63706 = _T_63705[10:0]; // @[Modules.scala 56:109:@11085.4]
  assign buffer_2_715 = $signed(_T_63706); // @[Modules.scala 56:109:@11086.4]
  assign _T_63708 = $signed(buffer_2_648) + $signed(buffer_2_649); // @[Modules.scala 56:109:@11088.4]
  assign _T_63709 = _T_63708[10:0]; // @[Modules.scala 56:109:@11089.4]
  assign buffer_2_716 = $signed(_T_63709); // @[Modules.scala 56:109:@11090.4]
  assign _T_63711 = $signed(buffer_2_650) + $signed(buffer_2_651); // @[Modules.scala 56:109:@11092.4]
  assign _T_63712 = _T_63711[10:0]; // @[Modules.scala 56:109:@11093.4]
  assign buffer_2_717 = $signed(_T_63712); // @[Modules.scala 56:109:@11094.4]
  assign _T_63714 = $signed(buffer_2_652) + $signed(buffer_2_653); // @[Modules.scala 56:109:@11096.4]
  assign _T_63715 = _T_63714[10:0]; // @[Modules.scala 56:109:@11097.4]
  assign buffer_2_718 = $signed(_T_63715); // @[Modules.scala 56:109:@11098.4]
  assign _T_63717 = $signed(buffer_2_654) + $signed(buffer_0_655); // @[Modules.scala 56:109:@11100.4]
  assign _T_63718 = _T_63717[10:0]; // @[Modules.scala 56:109:@11101.4]
  assign buffer_2_719 = $signed(_T_63718); // @[Modules.scala 56:109:@11102.4]
  assign _T_63720 = $signed(buffer_2_656) + $signed(buffer_2_657); // @[Modules.scala 56:109:@11104.4]
  assign _T_63721 = _T_63720[10:0]; // @[Modules.scala 56:109:@11105.4]
  assign buffer_2_720 = $signed(_T_63721); // @[Modules.scala 56:109:@11106.4]
  assign _T_63723 = $signed(buffer_2_658) + $signed(buffer_2_659); // @[Modules.scala 56:109:@11108.4]
  assign _T_63724 = _T_63723[10:0]; // @[Modules.scala 56:109:@11109.4]
  assign buffer_2_721 = $signed(_T_63724); // @[Modules.scala 56:109:@11110.4]
  assign _T_63726 = $signed(buffer_2_660) + $signed(buffer_2_661); // @[Modules.scala 56:109:@11112.4]
  assign _T_63727 = _T_63726[10:0]; // @[Modules.scala 56:109:@11113.4]
  assign buffer_2_722 = $signed(_T_63727); // @[Modules.scala 56:109:@11114.4]
  assign _T_63729 = $signed(buffer_2_662) + $signed(buffer_2_663); // @[Modules.scala 56:109:@11116.4]
  assign _T_63730 = _T_63729[10:0]; // @[Modules.scala 56:109:@11117.4]
  assign buffer_2_723 = $signed(_T_63730); // @[Modules.scala 56:109:@11118.4]
  assign _T_63732 = $signed(buffer_2_664) + $signed(buffer_2_665); // @[Modules.scala 56:109:@11120.4]
  assign _T_63733 = _T_63732[10:0]; // @[Modules.scala 56:109:@11121.4]
  assign buffer_2_724 = $signed(_T_63733); // @[Modules.scala 56:109:@11122.4]
  assign _T_63735 = $signed(buffer_2_666) + $signed(buffer_2_667); // @[Modules.scala 56:109:@11124.4]
  assign _T_63736 = _T_63735[10:0]; // @[Modules.scala 56:109:@11125.4]
  assign buffer_2_725 = $signed(_T_63736); // @[Modules.scala 56:109:@11126.4]
  assign _T_63738 = $signed(buffer_2_668) + $signed(buffer_2_669); // @[Modules.scala 56:109:@11128.4]
  assign _T_63739 = _T_63738[10:0]; // @[Modules.scala 56:109:@11129.4]
  assign buffer_2_726 = $signed(_T_63739); // @[Modules.scala 56:109:@11130.4]
  assign _T_63741 = $signed(buffer_2_670) + $signed(buffer_2_671); // @[Modules.scala 56:109:@11132.4]
  assign _T_63742 = _T_63741[10:0]; // @[Modules.scala 56:109:@11133.4]
  assign buffer_2_727 = $signed(_T_63742); // @[Modules.scala 56:109:@11134.4]
  assign _T_63744 = $signed(buffer_2_672) + $signed(buffer_2_673); // @[Modules.scala 56:109:@11136.4]
  assign _T_63745 = _T_63744[10:0]; // @[Modules.scala 56:109:@11137.4]
  assign buffer_2_728 = $signed(_T_63745); // @[Modules.scala 56:109:@11138.4]
  assign _T_63747 = $signed(buffer_2_674) + $signed(buffer_2_675); // @[Modules.scala 56:109:@11140.4]
  assign _T_63748 = _T_63747[10:0]; // @[Modules.scala 56:109:@11141.4]
  assign buffer_2_729 = $signed(_T_63748); // @[Modules.scala 56:109:@11142.4]
  assign _T_63750 = $signed(buffer_2_676) + $signed(buffer_2_677); // @[Modules.scala 56:109:@11144.4]
  assign _T_63751 = _T_63750[10:0]; // @[Modules.scala 56:109:@11145.4]
  assign buffer_2_730 = $signed(_T_63751); // @[Modules.scala 56:109:@11146.4]
  assign _T_63753 = $signed(buffer_0_678) + $signed(buffer_2_679); // @[Modules.scala 56:109:@11148.4]
  assign _T_63754 = _T_63753[10:0]; // @[Modules.scala 56:109:@11149.4]
  assign buffer_2_731 = $signed(_T_63754); // @[Modules.scala 56:109:@11150.4]
  assign _T_63756 = $signed(buffer_1_680) + $signed(buffer_2_681); // @[Modules.scala 56:109:@11152.4]
  assign _T_63757 = _T_63756[10:0]; // @[Modules.scala 56:109:@11153.4]
  assign buffer_2_732 = $signed(_T_63757); // @[Modules.scala 56:109:@11154.4]
  assign _T_63759 = $signed(buffer_2_682) + $signed(buffer_0_683); // @[Modules.scala 56:109:@11156.4]
  assign _T_63760 = _T_63759[10:0]; // @[Modules.scala 56:109:@11157.4]
  assign buffer_2_733 = $signed(_T_63760); // @[Modules.scala 56:109:@11158.4]
  assign _T_63762 = $signed(buffer_1_684) + $signed(buffer_2_685); // @[Modules.scala 56:109:@11160.4]
  assign _T_63763 = _T_63762[10:0]; // @[Modules.scala 56:109:@11161.4]
  assign buffer_2_734 = $signed(_T_63763); // @[Modules.scala 56:109:@11162.4]
  assign _T_63765 = $signed(buffer_2_686) + $signed(buffer_2_687); // @[Modules.scala 63:156:@11165.4]
  assign _T_63766 = _T_63765[10:0]; // @[Modules.scala 63:156:@11166.4]
  assign buffer_2_736 = $signed(_T_63766); // @[Modules.scala 63:156:@11167.4]
  assign _T_63768 = $signed(buffer_2_736) + $signed(buffer_2_688); // @[Modules.scala 63:156:@11169.4]
  assign _T_63769 = _T_63768[10:0]; // @[Modules.scala 63:156:@11170.4]
  assign buffer_2_737 = $signed(_T_63769); // @[Modules.scala 63:156:@11171.4]
  assign _T_63771 = $signed(buffer_2_737) + $signed(buffer_2_689); // @[Modules.scala 63:156:@11173.4]
  assign _T_63772 = _T_63771[10:0]; // @[Modules.scala 63:156:@11174.4]
  assign buffer_2_738 = $signed(_T_63772); // @[Modules.scala 63:156:@11175.4]
  assign _T_63774 = $signed(buffer_2_738) + $signed(buffer_2_690); // @[Modules.scala 63:156:@11177.4]
  assign _T_63775 = _T_63774[10:0]; // @[Modules.scala 63:156:@11178.4]
  assign buffer_2_739 = $signed(_T_63775); // @[Modules.scala 63:156:@11179.4]
  assign _T_63777 = $signed(buffer_2_739) + $signed(buffer_2_691); // @[Modules.scala 63:156:@11181.4]
  assign _T_63778 = _T_63777[10:0]; // @[Modules.scala 63:156:@11182.4]
  assign buffer_2_740 = $signed(_T_63778); // @[Modules.scala 63:156:@11183.4]
  assign _T_63780 = $signed(buffer_2_740) + $signed(buffer_2_692); // @[Modules.scala 63:156:@11185.4]
  assign _T_63781 = _T_63780[10:0]; // @[Modules.scala 63:156:@11186.4]
  assign buffer_2_741 = $signed(_T_63781); // @[Modules.scala 63:156:@11187.4]
  assign _T_63783 = $signed(buffer_2_741) + $signed(buffer_2_693); // @[Modules.scala 63:156:@11189.4]
  assign _T_63784 = _T_63783[10:0]; // @[Modules.scala 63:156:@11190.4]
  assign buffer_2_742 = $signed(_T_63784); // @[Modules.scala 63:156:@11191.4]
  assign _T_63786 = $signed(buffer_2_742) + $signed(buffer_2_694); // @[Modules.scala 63:156:@11193.4]
  assign _T_63787 = _T_63786[10:0]; // @[Modules.scala 63:156:@11194.4]
  assign buffer_2_743 = $signed(_T_63787); // @[Modules.scala 63:156:@11195.4]
  assign _T_63789 = $signed(buffer_2_743) + $signed(buffer_2_695); // @[Modules.scala 63:156:@11197.4]
  assign _T_63790 = _T_63789[10:0]; // @[Modules.scala 63:156:@11198.4]
  assign buffer_2_744 = $signed(_T_63790); // @[Modules.scala 63:156:@11199.4]
  assign _T_63792 = $signed(buffer_2_744) + $signed(buffer_2_696); // @[Modules.scala 63:156:@11201.4]
  assign _T_63793 = _T_63792[10:0]; // @[Modules.scala 63:156:@11202.4]
  assign buffer_2_745 = $signed(_T_63793); // @[Modules.scala 63:156:@11203.4]
  assign _T_63795 = $signed(buffer_2_745) + $signed(buffer_2_697); // @[Modules.scala 63:156:@11205.4]
  assign _T_63796 = _T_63795[10:0]; // @[Modules.scala 63:156:@11206.4]
  assign buffer_2_746 = $signed(_T_63796); // @[Modules.scala 63:156:@11207.4]
  assign _T_63798 = $signed(buffer_2_746) + $signed(buffer_2_698); // @[Modules.scala 63:156:@11209.4]
  assign _T_63799 = _T_63798[10:0]; // @[Modules.scala 63:156:@11210.4]
  assign buffer_2_747 = $signed(_T_63799); // @[Modules.scala 63:156:@11211.4]
  assign _T_63801 = $signed(buffer_2_747) + $signed(buffer_2_699); // @[Modules.scala 63:156:@11213.4]
  assign _T_63802 = _T_63801[10:0]; // @[Modules.scala 63:156:@11214.4]
  assign buffer_2_748 = $signed(_T_63802); // @[Modules.scala 63:156:@11215.4]
  assign _T_63804 = $signed(buffer_2_748) + $signed(buffer_2_700); // @[Modules.scala 63:156:@11217.4]
  assign _T_63805 = _T_63804[10:0]; // @[Modules.scala 63:156:@11218.4]
  assign buffer_2_749 = $signed(_T_63805); // @[Modules.scala 63:156:@11219.4]
  assign _T_63807 = $signed(buffer_2_749) + $signed(buffer_2_701); // @[Modules.scala 63:156:@11221.4]
  assign _T_63808 = _T_63807[10:0]; // @[Modules.scala 63:156:@11222.4]
  assign buffer_2_750 = $signed(_T_63808); // @[Modules.scala 63:156:@11223.4]
  assign _T_63810 = $signed(buffer_2_750) + $signed(buffer_2_702); // @[Modules.scala 63:156:@11225.4]
  assign _T_63811 = _T_63810[10:0]; // @[Modules.scala 63:156:@11226.4]
  assign buffer_2_751 = $signed(_T_63811); // @[Modules.scala 63:156:@11227.4]
  assign _T_63813 = $signed(buffer_2_751) + $signed(buffer_2_703); // @[Modules.scala 63:156:@11229.4]
  assign _T_63814 = _T_63813[10:0]; // @[Modules.scala 63:156:@11230.4]
  assign buffer_2_752 = $signed(_T_63814); // @[Modules.scala 63:156:@11231.4]
  assign _T_63816 = $signed(buffer_2_752) + $signed(buffer_2_704); // @[Modules.scala 63:156:@11233.4]
  assign _T_63817 = _T_63816[10:0]; // @[Modules.scala 63:156:@11234.4]
  assign buffer_2_753 = $signed(_T_63817); // @[Modules.scala 63:156:@11235.4]
  assign _T_63819 = $signed(buffer_2_753) + $signed(buffer_2_705); // @[Modules.scala 63:156:@11237.4]
  assign _T_63820 = _T_63819[10:0]; // @[Modules.scala 63:156:@11238.4]
  assign buffer_2_754 = $signed(_T_63820); // @[Modules.scala 63:156:@11239.4]
  assign _T_63822 = $signed(buffer_2_754) + $signed(buffer_2_706); // @[Modules.scala 63:156:@11241.4]
  assign _T_63823 = _T_63822[10:0]; // @[Modules.scala 63:156:@11242.4]
  assign buffer_2_755 = $signed(_T_63823); // @[Modules.scala 63:156:@11243.4]
  assign _T_63825 = $signed(buffer_2_755) + $signed(buffer_0_707); // @[Modules.scala 63:156:@11245.4]
  assign _T_63826 = _T_63825[10:0]; // @[Modules.scala 63:156:@11246.4]
  assign buffer_2_756 = $signed(_T_63826); // @[Modules.scala 63:156:@11247.4]
  assign _T_63828 = $signed(buffer_2_756) + $signed(buffer_2_708); // @[Modules.scala 63:156:@11249.4]
  assign _T_63829 = _T_63828[10:0]; // @[Modules.scala 63:156:@11250.4]
  assign buffer_2_757 = $signed(_T_63829); // @[Modules.scala 63:156:@11251.4]
  assign _T_63831 = $signed(buffer_2_757) + $signed(buffer_2_709); // @[Modules.scala 63:156:@11253.4]
  assign _T_63832 = _T_63831[10:0]; // @[Modules.scala 63:156:@11254.4]
  assign buffer_2_758 = $signed(_T_63832); // @[Modules.scala 63:156:@11255.4]
  assign _T_63834 = $signed(buffer_2_758) + $signed(buffer_2_710); // @[Modules.scala 63:156:@11257.4]
  assign _T_63835 = _T_63834[10:0]; // @[Modules.scala 63:156:@11258.4]
  assign buffer_2_759 = $signed(_T_63835); // @[Modules.scala 63:156:@11259.4]
  assign _T_63837 = $signed(buffer_2_759) + $signed(buffer_2_711); // @[Modules.scala 63:156:@11261.4]
  assign _T_63838 = _T_63837[10:0]; // @[Modules.scala 63:156:@11262.4]
  assign buffer_2_760 = $signed(_T_63838); // @[Modules.scala 63:156:@11263.4]
  assign _T_63840 = $signed(buffer_2_760) + $signed(buffer_2_712); // @[Modules.scala 63:156:@11265.4]
  assign _T_63841 = _T_63840[10:0]; // @[Modules.scala 63:156:@11266.4]
  assign buffer_2_761 = $signed(_T_63841); // @[Modules.scala 63:156:@11267.4]
  assign _T_63843 = $signed(buffer_2_761) + $signed(buffer_2_713); // @[Modules.scala 63:156:@11269.4]
  assign _T_63844 = _T_63843[10:0]; // @[Modules.scala 63:156:@11270.4]
  assign buffer_2_762 = $signed(_T_63844); // @[Modules.scala 63:156:@11271.4]
  assign _T_63846 = $signed(buffer_2_762) + $signed(buffer_2_714); // @[Modules.scala 63:156:@11273.4]
  assign _T_63847 = _T_63846[10:0]; // @[Modules.scala 63:156:@11274.4]
  assign buffer_2_763 = $signed(_T_63847); // @[Modules.scala 63:156:@11275.4]
  assign _T_63849 = $signed(buffer_2_763) + $signed(buffer_2_715); // @[Modules.scala 63:156:@11277.4]
  assign _T_63850 = _T_63849[10:0]; // @[Modules.scala 63:156:@11278.4]
  assign buffer_2_764 = $signed(_T_63850); // @[Modules.scala 63:156:@11279.4]
  assign _T_63852 = $signed(buffer_2_764) + $signed(buffer_2_716); // @[Modules.scala 63:156:@11281.4]
  assign _T_63853 = _T_63852[10:0]; // @[Modules.scala 63:156:@11282.4]
  assign buffer_2_765 = $signed(_T_63853); // @[Modules.scala 63:156:@11283.4]
  assign _T_63855 = $signed(buffer_2_765) + $signed(buffer_2_717); // @[Modules.scala 63:156:@11285.4]
  assign _T_63856 = _T_63855[10:0]; // @[Modules.scala 63:156:@11286.4]
  assign buffer_2_766 = $signed(_T_63856); // @[Modules.scala 63:156:@11287.4]
  assign _T_63858 = $signed(buffer_2_766) + $signed(buffer_2_718); // @[Modules.scala 63:156:@11289.4]
  assign _T_63859 = _T_63858[10:0]; // @[Modules.scala 63:156:@11290.4]
  assign buffer_2_767 = $signed(_T_63859); // @[Modules.scala 63:156:@11291.4]
  assign _T_63861 = $signed(buffer_2_767) + $signed(buffer_2_719); // @[Modules.scala 63:156:@11293.4]
  assign _T_63862 = _T_63861[10:0]; // @[Modules.scala 63:156:@11294.4]
  assign buffer_2_768 = $signed(_T_63862); // @[Modules.scala 63:156:@11295.4]
  assign _T_63864 = $signed(buffer_2_768) + $signed(buffer_2_720); // @[Modules.scala 63:156:@11297.4]
  assign _T_63865 = _T_63864[10:0]; // @[Modules.scala 63:156:@11298.4]
  assign buffer_2_769 = $signed(_T_63865); // @[Modules.scala 63:156:@11299.4]
  assign _T_63867 = $signed(buffer_2_769) + $signed(buffer_2_721); // @[Modules.scala 63:156:@11301.4]
  assign _T_63868 = _T_63867[10:0]; // @[Modules.scala 63:156:@11302.4]
  assign buffer_2_770 = $signed(_T_63868); // @[Modules.scala 63:156:@11303.4]
  assign _T_63870 = $signed(buffer_2_770) + $signed(buffer_2_722); // @[Modules.scala 63:156:@11305.4]
  assign _T_63871 = _T_63870[10:0]; // @[Modules.scala 63:156:@11306.4]
  assign buffer_2_771 = $signed(_T_63871); // @[Modules.scala 63:156:@11307.4]
  assign _T_63873 = $signed(buffer_2_771) + $signed(buffer_2_723); // @[Modules.scala 63:156:@11309.4]
  assign _T_63874 = _T_63873[10:0]; // @[Modules.scala 63:156:@11310.4]
  assign buffer_2_772 = $signed(_T_63874); // @[Modules.scala 63:156:@11311.4]
  assign _T_63876 = $signed(buffer_2_772) + $signed(buffer_2_724); // @[Modules.scala 63:156:@11313.4]
  assign _T_63877 = _T_63876[10:0]; // @[Modules.scala 63:156:@11314.4]
  assign buffer_2_773 = $signed(_T_63877); // @[Modules.scala 63:156:@11315.4]
  assign _T_63879 = $signed(buffer_2_773) + $signed(buffer_2_725); // @[Modules.scala 63:156:@11317.4]
  assign _T_63880 = _T_63879[10:0]; // @[Modules.scala 63:156:@11318.4]
  assign buffer_2_774 = $signed(_T_63880); // @[Modules.scala 63:156:@11319.4]
  assign _T_63882 = $signed(buffer_2_774) + $signed(buffer_2_726); // @[Modules.scala 63:156:@11321.4]
  assign _T_63883 = _T_63882[10:0]; // @[Modules.scala 63:156:@11322.4]
  assign buffer_2_775 = $signed(_T_63883); // @[Modules.scala 63:156:@11323.4]
  assign _T_63885 = $signed(buffer_2_775) + $signed(buffer_2_727); // @[Modules.scala 63:156:@11325.4]
  assign _T_63886 = _T_63885[10:0]; // @[Modules.scala 63:156:@11326.4]
  assign buffer_2_776 = $signed(_T_63886); // @[Modules.scala 63:156:@11327.4]
  assign _T_63888 = $signed(buffer_2_776) + $signed(buffer_2_728); // @[Modules.scala 63:156:@11329.4]
  assign _T_63889 = _T_63888[10:0]; // @[Modules.scala 63:156:@11330.4]
  assign buffer_2_777 = $signed(_T_63889); // @[Modules.scala 63:156:@11331.4]
  assign _T_63891 = $signed(buffer_2_777) + $signed(buffer_2_729); // @[Modules.scala 63:156:@11333.4]
  assign _T_63892 = _T_63891[10:0]; // @[Modules.scala 63:156:@11334.4]
  assign buffer_2_778 = $signed(_T_63892); // @[Modules.scala 63:156:@11335.4]
  assign _T_63894 = $signed(buffer_2_778) + $signed(buffer_2_730); // @[Modules.scala 63:156:@11337.4]
  assign _T_63895 = _T_63894[10:0]; // @[Modules.scala 63:156:@11338.4]
  assign buffer_2_779 = $signed(_T_63895); // @[Modules.scala 63:156:@11339.4]
  assign _T_63897 = $signed(buffer_2_779) + $signed(buffer_2_731); // @[Modules.scala 63:156:@11341.4]
  assign _T_63898 = _T_63897[10:0]; // @[Modules.scala 63:156:@11342.4]
  assign buffer_2_780 = $signed(_T_63898); // @[Modules.scala 63:156:@11343.4]
  assign _T_63900 = $signed(buffer_2_780) + $signed(buffer_2_732); // @[Modules.scala 63:156:@11345.4]
  assign _T_63901 = _T_63900[10:0]; // @[Modules.scala 63:156:@11346.4]
  assign buffer_2_781 = $signed(_T_63901); // @[Modules.scala 63:156:@11347.4]
  assign _T_63903 = $signed(buffer_2_781) + $signed(buffer_2_733); // @[Modules.scala 63:156:@11349.4]
  assign _T_63904 = _T_63903[10:0]; // @[Modules.scala 63:156:@11350.4]
  assign buffer_2_782 = $signed(_T_63904); // @[Modules.scala 63:156:@11351.4]
  assign _T_63906 = $signed(buffer_2_782) + $signed(buffer_2_734); // @[Modules.scala 63:156:@11353.4]
  assign _T_63907 = _T_63906[10:0]; // @[Modules.scala 63:156:@11354.4]
  assign buffer_2_783 = $signed(_T_63907); // @[Modules.scala 63:156:@11355.4]
  assign _T_63909 = $signed(io_in_0) - $signed(io_in_1); // @[Modules.scala 40:46:@11358.4]
  assign _T_63910 = _T_63909[4:0]; // @[Modules.scala 40:46:@11359.4]
  assign _T_63911 = $signed(_T_63910); // @[Modules.scala 40:46:@11360.4]
  assign _T_63912 = $signed(io_in_2) - $signed(io_in_3); // @[Modules.scala 40:46:@11362.4]
  assign _T_63913 = _T_63912[4:0]; // @[Modules.scala 40:46:@11363.4]
  assign _T_63914 = $signed(_T_63913); // @[Modules.scala 40:46:@11364.4]
  assign _T_63925 = $signed(_T_54297) - $signed(io_in_9); // @[Modules.scala 46:47:@11377.4]
  assign _T_63926 = _T_63925[4:0]; // @[Modules.scala 46:47:@11378.4]
  assign _T_63927 = $signed(_T_63926); // @[Modules.scala 46:47:@11379.4]
  assign _T_63928 = $signed(io_in_10) - $signed(io_in_11); // @[Modules.scala 40:46:@11381.4]
  assign _T_63929 = _T_63928[4:0]; // @[Modules.scala 40:46:@11382.4]
  assign _T_63930 = $signed(_T_63929); // @[Modules.scala 40:46:@11383.4]
  assign _T_63957 = $signed(io_in_24) - $signed(io_in_25); // @[Modules.scala 40:46:@11415.4]
  assign _T_63958 = _T_63957[4:0]; // @[Modules.scala 40:46:@11416.4]
  assign _T_63959 = $signed(_T_63958); // @[Modules.scala 40:46:@11417.4]
  assign _T_63960 = $signed(io_in_26) + $signed(io_in_27); // @[Modules.scala 37:46:@11419.4]
  assign _T_63961 = _T_63960[4:0]; // @[Modules.scala 37:46:@11420.4]
  assign _T_63962 = $signed(_T_63961); // @[Modules.scala 37:46:@11421.4]
  assign _T_63963 = $signed(io_in_28) + $signed(io_in_29); // @[Modules.scala 37:46:@11423.4]
  assign _T_63964 = _T_63963[4:0]; // @[Modules.scala 37:46:@11424.4]
  assign _T_63965 = $signed(_T_63964); // @[Modules.scala 37:46:@11425.4]
  assign _T_63970 = $signed(_T_54362) - $signed(io_in_31); // @[Modules.scala 46:47:@11430.4]
  assign _T_63971 = _T_63970[4:0]; // @[Modules.scala 46:47:@11431.4]
  assign _T_63972 = $signed(_T_63971); // @[Modules.scala 46:47:@11432.4]
  assign _T_63973 = $signed(io_in_32) - $signed(io_in_33); // @[Modules.scala 40:46:@11434.4]
  assign _T_63974 = _T_63973[4:0]; // @[Modules.scala 40:46:@11435.4]
  assign _T_63975 = $signed(_T_63974); // @[Modules.scala 40:46:@11436.4]
  assign _T_64031 = $signed(_T_60745) + $signed(io_in_53); // @[Modules.scala 43:47:@11495.4]
  assign _T_64032 = _T_64031[4:0]; // @[Modules.scala 43:47:@11496.4]
  assign _T_64033 = $signed(_T_64032); // @[Modules.scala 43:47:@11497.4]
  assign _T_64038 = $signed(_T_57651) - $signed(io_in_55); // @[Modules.scala 46:47:@11502.4]
  assign _T_64039 = _T_64038[4:0]; // @[Modules.scala 46:47:@11503.4]
  assign _T_64040 = $signed(_T_64039); // @[Modules.scala 46:47:@11504.4]
  assign _T_64045 = $signed(_T_57658) - $signed(io_in_57); // @[Modules.scala 46:47:@11509.4]
  assign _T_64046 = _T_64045[4:0]; // @[Modules.scala 46:47:@11510.4]
  assign _T_64047 = $signed(_T_64046); // @[Modules.scala 46:47:@11511.4]
  assign _T_64048 = $signed(io_in_58) - $signed(io_in_59); // @[Modules.scala 40:46:@11513.4]
  assign _T_64049 = _T_64048[4:0]; // @[Modules.scala 40:46:@11514.4]
  assign _T_64050 = $signed(_T_64049); // @[Modules.scala 40:46:@11515.4]
  assign _T_64055 = $signed(_T_54451) + $signed(io_in_61); // @[Modules.scala 43:47:@11520.4]
  assign _T_64056 = _T_64055[4:0]; // @[Modules.scala 43:47:@11521.4]
  assign _T_64057 = $signed(_T_64056); // @[Modules.scala 43:47:@11522.4]
  assign _T_64069 = $signed(_T_54465) - $signed(io_in_65); // @[Modules.scala 46:47:@11534.4]
  assign _T_64070 = _T_64069[4:0]; // @[Modules.scala 46:47:@11535.4]
  assign _T_64071 = $signed(_T_64070); // @[Modules.scala 46:47:@11536.4]
  assign _T_64104 = $signed(_T_54500) - $signed(io_in_75); // @[Modules.scala 46:47:@11569.4]
  assign _T_64105 = _T_64104[4:0]; // @[Modules.scala 46:47:@11570.4]
  assign _T_64106 = $signed(_T_64105); // @[Modules.scala 46:47:@11571.4]
  assign _T_64108 = $signed(5'sh0) - $signed(io_in_76); // @[Modules.scala 46:37:@11573.4]
  assign _T_64109 = _T_64108[4:0]; // @[Modules.scala 46:37:@11574.4]
  assign _T_64110 = $signed(_T_64109); // @[Modules.scala 46:37:@11575.4]
  assign _T_64111 = $signed(_T_64110) - $signed(io_in_77); // @[Modules.scala 46:47:@11576.4]
  assign _T_64112 = _T_64111[4:0]; // @[Modules.scala 46:47:@11577.4]
  assign _T_64113 = $signed(_T_64112); // @[Modules.scala 46:47:@11578.4]
  assign _T_64115 = $signed(5'sh0) - $signed(io_in_78); // @[Modules.scala 46:37:@11580.4]
  assign _T_64116 = _T_64115[4:0]; // @[Modules.scala 46:37:@11581.4]
  assign _T_64117 = $signed(_T_64116); // @[Modules.scala 46:37:@11582.4]
  assign _T_64118 = $signed(_T_64117) - $signed(io_in_79); // @[Modules.scala 46:47:@11583.4]
  assign _T_64119 = _T_64118[4:0]; // @[Modules.scala 46:47:@11584.4]
  assign _T_64120 = $signed(_T_64119); // @[Modules.scala 46:47:@11585.4]
  assign _T_64130 = $signed(io_in_86) - $signed(io_in_87); // @[Modules.scala 40:46:@11599.4]
  assign _T_64131 = _T_64130[4:0]; // @[Modules.scala 40:46:@11600.4]
  assign _T_64132 = $signed(_T_64131); // @[Modules.scala 40:46:@11601.4]
  assign _T_64134 = $signed(5'sh0) - $signed(io_in_88); // @[Modules.scala 46:37:@11603.4]
  assign _T_64135 = _T_64134[4:0]; // @[Modules.scala 46:37:@11604.4]
  assign _T_64136 = $signed(_T_64135); // @[Modules.scala 46:37:@11605.4]
  assign _T_64137 = $signed(_T_64136) - $signed(io_in_89); // @[Modules.scala 46:47:@11606.4]
  assign _T_64138 = _T_64137[4:0]; // @[Modules.scala 46:47:@11607.4]
  assign _T_64139 = $signed(_T_64138); // @[Modules.scala 46:47:@11608.4]
  assign _T_64141 = $signed(5'sh0) - $signed(io_in_90); // @[Modules.scala 46:37:@11610.4]
  assign _T_64142 = _T_64141[4:0]; // @[Modules.scala 46:37:@11611.4]
  assign _T_64143 = $signed(_T_64142); // @[Modules.scala 46:37:@11612.4]
  assign _T_64144 = $signed(_T_64143) - $signed(io_in_91); // @[Modules.scala 46:47:@11613.4]
  assign _T_64145 = _T_64144[4:0]; // @[Modules.scala 46:47:@11614.4]
  assign _T_64146 = $signed(_T_64145); // @[Modules.scala 46:47:@11615.4]
  assign _T_64151 = $signed(_T_54539) - $signed(io_in_93); // @[Modules.scala 46:47:@11620.4]
  assign _T_64152 = _T_64151[4:0]; // @[Modules.scala 46:47:@11621.4]
  assign _T_64153 = $signed(_T_64152); // @[Modules.scala 46:47:@11622.4]
  assign _T_64160 = $signed(io_in_98) - $signed(io_in_99); // @[Modules.scala 40:46:@11632.4]
  assign _T_64161 = _T_64160[4:0]; // @[Modules.scala 40:46:@11633.4]
  assign _T_64162 = $signed(_T_64161); // @[Modules.scala 40:46:@11634.4]
  assign _T_64167 = $signed(5'sh0) - $signed(io_in_102); // @[Modules.scala 46:37:@11640.4]
  assign _T_64168 = _T_64167[4:0]; // @[Modules.scala 46:37:@11641.4]
  assign _T_64169 = $signed(_T_64168); // @[Modules.scala 46:37:@11642.4]
  assign _T_64170 = $signed(_T_64169) - $signed(io_in_103); // @[Modules.scala 46:47:@11643.4]
  assign _T_64171 = _T_64170[4:0]; // @[Modules.scala 46:47:@11644.4]
  assign _T_64172 = $signed(_T_64171); // @[Modules.scala 46:47:@11645.4]
  assign _T_64174 = $signed(5'sh0) - $signed(io_in_104); // @[Modules.scala 46:37:@11647.4]
  assign _T_64175 = _T_64174[4:0]; // @[Modules.scala 46:37:@11648.4]
  assign _T_64176 = $signed(_T_64175); // @[Modules.scala 46:37:@11649.4]
  assign _T_64177 = $signed(_T_64176) - $signed(io_in_105); // @[Modules.scala 46:47:@11650.4]
  assign _T_64178 = _T_64177[4:0]; // @[Modules.scala 46:47:@11651.4]
  assign _T_64179 = $signed(_T_64178); // @[Modules.scala 46:47:@11652.4]
  assign _T_64181 = $signed(5'sh0) - $signed(io_in_106); // @[Modules.scala 46:37:@11654.4]
  assign _T_64182 = _T_64181[4:0]; // @[Modules.scala 46:37:@11655.4]
  assign _T_64183 = $signed(_T_64182); // @[Modules.scala 46:37:@11656.4]
  assign _T_64184 = $signed(_T_64183) - $signed(io_in_107); // @[Modules.scala 46:47:@11657.4]
  assign _T_64185 = _T_64184[4:0]; // @[Modules.scala 46:47:@11658.4]
  assign _T_64186 = $signed(_T_64185); // @[Modules.scala 46:47:@11659.4]
  assign _T_64191 = $signed(_T_60877) + $signed(io_in_109); // @[Modules.scala 43:47:@11664.4]
  assign _T_64192 = _T_64191[4:0]; // @[Modules.scala 43:47:@11665.4]
  assign _T_64193 = $signed(_T_64192); // @[Modules.scala 43:47:@11666.4]
  assign _T_64194 = $signed(io_in_110) - $signed(io_in_111); // @[Modules.scala 40:46:@11668.4]
  assign _T_64195 = _T_64194[4:0]; // @[Modules.scala 40:46:@11669.4]
  assign _T_64196 = $signed(_T_64195); // @[Modules.scala 40:46:@11670.4]
  assign _T_64197 = $signed(io_in_112) - $signed(io_in_113); // @[Modules.scala 40:46:@11672.4]
  assign _T_64198 = _T_64197[4:0]; // @[Modules.scala 40:46:@11673.4]
  assign _T_64199 = $signed(_T_64198); // @[Modules.scala 40:46:@11674.4]
  assign _T_64200 = $signed(io_in_114) + $signed(io_in_115); // @[Modules.scala 37:46:@11676.4]
  assign _T_64201 = _T_64200[4:0]; // @[Modules.scala 37:46:@11677.4]
  assign _T_64202 = $signed(_T_64201); // @[Modules.scala 37:46:@11678.4]
  assign _T_64213 = $signed(io_in_120) + $signed(io_in_121); // @[Modules.scala 37:46:@11691.4]
  assign _T_64214 = _T_64213[4:0]; // @[Modules.scala 37:46:@11692.4]
  assign _T_64215 = $signed(_T_64214); // @[Modules.scala 37:46:@11693.4]
  assign _T_64216 = $signed(io_in_122) + $signed(io_in_123); // @[Modules.scala 37:46:@11695.4]
  assign _T_64217 = _T_64216[4:0]; // @[Modules.scala 37:46:@11696.4]
  assign _T_64218 = $signed(_T_64217); // @[Modules.scala 37:46:@11697.4]
  assign _T_64219 = $signed(io_in_124) + $signed(io_in_125); // @[Modules.scala 37:46:@11699.4]
  assign _T_64220 = _T_64219[4:0]; // @[Modules.scala 37:46:@11700.4]
  assign _T_64221 = $signed(_T_64220); // @[Modules.scala 37:46:@11701.4]
  assign _T_64222 = $signed(io_in_126) + $signed(io_in_127); // @[Modules.scala 37:46:@11703.4]
  assign _T_64223 = _T_64222[4:0]; // @[Modules.scala 37:46:@11704.4]
  assign _T_64224 = $signed(_T_64223); // @[Modules.scala 37:46:@11705.4]
  assign _T_64235 = $signed(_T_57816) - $signed(io_in_133); // @[Modules.scala 46:47:@11718.4]
  assign _T_64236 = _T_64235[4:0]; // @[Modules.scala 46:47:@11719.4]
  assign _T_64237 = $signed(_T_64236); // @[Modules.scala 46:47:@11720.4]
  assign _T_64238 = $signed(io_in_134) - $signed(io_in_135); // @[Modules.scala 40:46:@11722.4]
  assign _T_64239 = _T_64238[4:0]; // @[Modules.scala 40:46:@11723.4]
  assign _T_64240 = $signed(_T_64239); // @[Modules.scala 40:46:@11724.4]
  assign _T_64244 = $signed(io_in_138) - $signed(io_in_139); // @[Modules.scala 40:46:@11730.4]
  assign _T_64245 = _T_64244[4:0]; // @[Modules.scala 40:46:@11731.4]
  assign _T_64246 = $signed(_T_64245); // @[Modules.scala 40:46:@11732.4]
  assign _T_64261 = $signed(_T_57846) + $signed(io_in_145); // @[Modules.scala 43:47:@11748.4]
  assign _T_64262 = _T_64261[4:0]; // @[Modules.scala 43:47:@11749.4]
  assign _T_64263 = $signed(_T_64262); // @[Modules.scala 43:47:@11750.4]
  assign _T_64270 = $signed(io_in_150) + $signed(io_in_151); // @[Modules.scala 37:46:@11760.4]
  assign _T_64271 = _T_64270[4:0]; // @[Modules.scala 37:46:@11761.4]
  assign _T_64272 = $signed(_T_64271); // @[Modules.scala 37:46:@11762.4]
  assign _T_64277 = $signed(_T_54681) + $signed(io_in_153); // @[Modules.scala 43:47:@11767.4]
  assign _T_64278 = _T_64277[4:0]; // @[Modules.scala 43:47:@11768.4]
  assign _T_64279 = $signed(_T_64278); // @[Modules.scala 43:47:@11769.4]
  assign _T_64280 = $signed(io_in_154) + $signed(io_in_155); // @[Modules.scala 37:46:@11771.4]
  assign _T_64281 = _T_64280[4:0]; // @[Modules.scala 37:46:@11772.4]
  assign _T_64282 = $signed(_T_64281); // @[Modules.scala 37:46:@11773.4]
  assign _T_64286 = $signed(io_in_158) + $signed(io_in_159); // @[Modules.scala 37:46:@11779.4]
  assign _T_64287 = _T_64286[4:0]; // @[Modules.scala 37:46:@11780.4]
  assign _T_64288 = $signed(_T_64287); // @[Modules.scala 37:46:@11781.4]
  assign _T_64311 = $signed(io_in_172) + $signed(io_in_173); // @[Modules.scala 37:46:@11810.4]
  assign _T_64312 = _T_64311[4:0]; // @[Modules.scala 37:46:@11811.4]
  assign _T_64313 = $signed(_T_64312); // @[Modules.scala 37:46:@11812.4]
  assign _T_64320 = $signed(io_in_178) + $signed(io_in_179); // @[Modules.scala 37:46:@11822.4]
  assign _T_64321 = _T_64320[4:0]; // @[Modules.scala 37:46:@11823.4]
  assign _T_64322 = $signed(_T_64321); // @[Modules.scala 37:46:@11824.4]
  assign _T_64323 = $signed(io_in_180) + $signed(io_in_181); // @[Modules.scala 37:46:@11826.4]
  assign _T_64324 = _T_64323[4:0]; // @[Modules.scala 37:46:@11827.4]
  assign _T_64325 = $signed(_T_64324); // @[Modules.scala 37:46:@11828.4]
  assign _T_64333 = $signed(io_in_184) - $signed(io_in_185); // @[Modules.scala 40:46:@11837.4]
  assign _T_64334 = _T_64333[4:0]; // @[Modules.scala 40:46:@11838.4]
  assign _T_64335 = $signed(_T_64334); // @[Modules.scala 40:46:@11839.4]
  assign _T_64336 = $signed(io_in_186) - $signed(io_in_187); // @[Modules.scala 40:46:@11841.4]
  assign _T_64337 = _T_64336[4:0]; // @[Modules.scala 40:46:@11842.4]
  assign _T_64338 = $signed(_T_64337); // @[Modules.scala 40:46:@11843.4]
  assign _T_64352 = $signed(5'sh0) - $signed(io_in_196); // @[Modules.scala 43:37:@11861.4]
  assign _T_64353 = _T_64352[4:0]; // @[Modules.scala 43:37:@11862.4]
  assign _T_64354 = $signed(_T_64353); // @[Modules.scala 43:37:@11863.4]
  assign _T_64355 = $signed(_T_64354) + $signed(io_in_197); // @[Modules.scala 43:47:@11864.4]
  assign _T_64356 = _T_64355[4:0]; // @[Modules.scala 43:47:@11865.4]
  assign _T_64357 = $signed(_T_64356); // @[Modules.scala 43:47:@11866.4]
  assign _T_64358 = $signed(io_in_198) + $signed(io_in_199); // @[Modules.scala 37:46:@11868.4]
  assign _T_64359 = _T_64358[4:0]; // @[Modules.scala 37:46:@11869.4]
  assign _T_64360 = $signed(_T_64359); // @[Modules.scala 37:46:@11870.4]
  assign _T_64361 = $signed(io_in_200) + $signed(io_in_201); // @[Modules.scala 37:46:@11872.4]
  assign _T_64362 = _T_64361[4:0]; // @[Modules.scala 37:46:@11873.4]
  assign _T_64363 = $signed(_T_64362); // @[Modules.scala 37:46:@11874.4]
  assign _T_64374 = $signed(io_in_206) + $signed(io_in_207); // @[Modules.scala 37:46:@11887.4]
  assign _T_64375 = _T_64374[4:0]; // @[Modules.scala 37:46:@11888.4]
  assign _T_64376 = $signed(_T_64375); // @[Modules.scala 37:46:@11889.4]
  assign _T_64377 = $signed(io_in_208) + $signed(io_in_209); // @[Modules.scala 37:46:@11891.4]
  assign _T_64378 = _T_64377[4:0]; // @[Modules.scala 37:46:@11892.4]
  assign _T_64379 = $signed(_T_64378); // @[Modules.scala 37:46:@11893.4]
  assign _T_64380 = $signed(io_in_210) - $signed(io_in_211); // @[Modules.scala 40:46:@11895.4]
  assign _T_64381 = _T_64380[4:0]; // @[Modules.scala 40:46:@11896.4]
  assign _T_64382 = $signed(_T_64381); // @[Modules.scala 40:46:@11897.4]
  assign _T_64383 = $signed(io_in_212) + $signed(io_in_213); // @[Modules.scala 37:46:@11899.4]
  assign _T_64384 = _T_64383[4:0]; // @[Modules.scala 37:46:@11900.4]
  assign _T_64385 = $signed(_T_64384); // @[Modules.scala 37:46:@11901.4]
  assign _T_64396 = $signed(io_in_218) - $signed(io_in_219); // @[Modules.scala 40:46:@11914.4]
  assign _T_64397 = _T_64396[4:0]; // @[Modules.scala 40:46:@11915.4]
  assign _T_64398 = $signed(_T_64397); // @[Modules.scala 40:46:@11916.4]
  assign _T_64408 = $signed(io_in_226) + $signed(io_in_227); // @[Modules.scala 37:46:@11930.4]
  assign _T_64409 = _T_64408[4:0]; // @[Modules.scala 37:46:@11931.4]
  assign _T_64410 = $signed(_T_64409); // @[Modules.scala 37:46:@11932.4]
  assign _T_64411 = $signed(io_in_228) + $signed(io_in_229); // @[Modules.scala 37:46:@11934.4]
  assign _T_64412 = _T_64411[4:0]; // @[Modules.scala 37:46:@11935.4]
  assign _T_64413 = $signed(_T_64412); // @[Modules.scala 37:46:@11936.4]
  assign _T_64418 = $signed(_T_54918) + $signed(io_in_231); // @[Modules.scala 43:47:@11941.4]
  assign _T_64419 = _T_64418[4:0]; // @[Modules.scala 43:47:@11942.4]
  assign _T_64420 = $signed(_T_64419); // @[Modules.scala 43:47:@11943.4]
  assign _T_64421 = $signed(io_in_232) - $signed(io_in_233); // @[Modules.scala 40:46:@11945.4]
  assign _T_64422 = _T_64421[4:0]; // @[Modules.scala 40:46:@11946.4]
  assign _T_64423 = $signed(_T_64422); // @[Modules.scala 40:46:@11947.4]
  assign _T_64424 = $signed(io_in_234) + $signed(io_in_235); // @[Modules.scala 37:46:@11949.4]
  assign _T_64425 = _T_64424[4:0]; // @[Modules.scala 37:46:@11950.4]
  assign _T_64426 = $signed(_T_64425); // @[Modules.scala 37:46:@11951.4]
  assign _T_64427 = $signed(io_in_236) + $signed(io_in_237); // @[Modules.scala 37:46:@11953.4]
  assign _T_64428 = _T_64427[4:0]; // @[Modules.scala 37:46:@11954.4]
  assign _T_64429 = $signed(_T_64428); // @[Modules.scala 37:46:@11955.4]
  assign _T_64430 = $signed(io_in_238) + $signed(io_in_239); // @[Modules.scala 37:46:@11957.4]
  assign _T_64431 = _T_64430[4:0]; // @[Modules.scala 37:46:@11958.4]
  assign _T_64432 = $signed(_T_64431); // @[Modules.scala 37:46:@11959.4]
  assign _T_64436 = $signed(io_in_242) + $signed(io_in_243); // @[Modules.scala 37:46:@11965.4]
  assign _T_64437 = _T_64436[4:0]; // @[Modules.scala 37:46:@11966.4]
  assign _T_64438 = $signed(_T_64437); // @[Modules.scala 37:46:@11967.4]
  assign _T_64439 = $signed(io_in_244) - $signed(io_in_245); // @[Modules.scala 40:46:@11969.4]
  assign _T_64440 = _T_64439[4:0]; // @[Modules.scala 40:46:@11970.4]
  assign _T_64441 = $signed(_T_64440); // @[Modules.scala 40:46:@11971.4]
  assign _T_64442 = $signed(io_in_246) + $signed(io_in_247); // @[Modules.scala 37:46:@11973.4]
  assign _T_64443 = _T_64442[4:0]; // @[Modules.scala 37:46:@11974.4]
  assign _T_64444 = $signed(_T_64443); // @[Modules.scala 37:46:@11975.4]
  assign _T_64451 = $signed(io_in_252) + $signed(io_in_253); // @[Modules.scala 37:46:@11985.4]
  assign _T_64452 = _T_64451[4:0]; // @[Modules.scala 37:46:@11986.4]
  assign _T_64453 = $signed(_T_64452); // @[Modules.scala 37:46:@11987.4]
  assign _T_64454 = $signed(io_in_254) + $signed(io_in_255); // @[Modules.scala 37:46:@11989.4]
  assign _T_64455 = _T_64454[4:0]; // @[Modules.scala 37:46:@11990.4]
  assign _T_64456 = $signed(_T_64455); // @[Modules.scala 37:46:@11991.4]
  assign _T_64457 = $signed(io_in_256) + $signed(io_in_257); // @[Modules.scala 37:46:@11993.4]
  assign _T_64458 = _T_64457[4:0]; // @[Modules.scala 37:46:@11994.4]
  assign _T_64459 = $signed(_T_64458); // @[Modules.scala 37:46:@11995.4]
  assign _T_64481 = $signed(io_in_264) + $signed(io_in_265); // @[Modules.scala 37:46:@12018.4]
  assign _T_64482 = _T_64481[4:0]; // @[Modules.scala 37:46:@12019.4]
  assign _T_64483 = $signed(_T_64482); // @[Modules.scala 37:46:@12020.4]
  assign _T_64487 = $signed(io_in_268) + $signed(io_in_269); // @[Modules.scala 37:46:@12026.4]
  assign _T_64488 = _T_64487[4:0]; // @[Modules.scala 37:46:@12027.4]
  assign _T_64489 = $signed(_T_64488); // @[Modules.scala 37:46:@12028.4]
  assign _T_64490 = $signed(io_in_270) + $signed(io_in_271); // @[Modules.scala 37:46:@12030.4]
  assign _T_64491 = _T_64490[4:0]; // @[Modules.scala 37:46:@12031.4]
  assign _T_64492 = $signed(_T_64491); // @[Modules.scala 37:46:@12032.4]
  assign _T_64493 = $signed(io_in_272) + $signed(io_in_273); // @[Modules.scala 37:46:@12034.4]
  assign _T_64494 = _T_64493[4:0]; // @[Modules.scala 37:46:@12035.4]
  assign _T_64495 = $signed(_T_64494); // @[Modules.scala 37:46:@12036.4]
  assign _T_64496 = $signed(io_in_274) + $signed(io_in_275); // @[Modules.scala 37:46:@12038.4]
  assign _T_64497 = _T_64496[4:0]; // @[Modules.scala 37:46:@12039.4]
  assign _T_64498 = $signed(_T_64497); // @[Modules.scala 37:46:@12040.4]
  assign _T_64505 = $signed(io_in_280) + $signed(io_in_281); // @[Modules.scala 37:46:@12050.4]
  assign _T_64506 = _T_64505[4:0]; // @[Modules.scala 37:46:@12051.4]
  assign _T_64507 = $signed(_T_64506); // @[Modules.scala 37:46:@12052.4]
  assign _T_64508 = $signed(io_in_282) + $signed(io_in_283); // @[Modules.scala 37:46:@12054.4]
  assign _T_64509 = _T_64508[4:0]; // @[Modules.scala 37:46:@12055.4]
  assign _T_64510 = $signed(_T_64509); // @[Modules.scala 37:46:@12056.4]
  assign _T_64511 = $signed(io_in_284) - $signed(io_in_285); // @[Modules.scala 40:46:@12058.4]
  assign _T_64512 = _T_64511[4:0]; // @[Modules.scala 40:46:@12059.4]
  assign _T_64513 = $signed(_T_64512); // @[Modules.scala 40:46:@12060.4]
  assign _T_64525 = $signed(_T_55117) - $signed(io_in_289); // @[Modules.scala 46:47:@12072.4]
  assign _T_64526 = _T_64525[4:0]; // @[Modules.scala 46:47:@12073.4]
  assign _T_64527 = $signed(_T_64526); // @[Modules.scala 46:47:@12074.4]
  assign _T_64546 = $signed(_T_55138) + $signed(io_in_295); // @[Modules.scala 43:47:@12093.4]
  assign _T_64547 = _T_64546[4:0]; // @[Modules.scala 43:47:@12094.4]
  assign _T_64548 = $signed(_T_64547); // @[Modules.scala 43:47:@12095.4]
  assign _T_64549 = $signed(io_in_296) + $signed(io_in_297); // @[Modules.scala 37:46:@12097.4]
  assign _T_64550 = _T_64549[4:0]; // @[Modules.scala 37:46:@12098.4]
  assign _T_64551 = $signed(_T_64550); // @[Modules.scala 37:46:@12099.4]
  assign _T_64552 = $signed(io_in_298) - $signed(io_in_299); // @[Modules.scala 40:46:@12101.4]
  assign _T_64553 = _T_64552[4:0]; // @[Modules.scala 40:46:@12102.4]
  assign _T_64554 = $signed(_T_64553); // @[Modules.scala 40:46:@12103.4]
  assign _T_64555 = $signed(io_in_300) - $signed(io_in_301); // @[Modules.scala 40:46:@12105.4]
  assign _T_64556 = _T_64555[4:0]; // @[Modules.scala 40:46:@12106.4]
  assign _T_64557 = $signed(_T_64556); // @[Modules.scala 40:46:@12107.4]
  assign _T_64575 = $signed(_T_55187) + $signed(io_in_309); // @[Modules.scala 43:47:@12127.4]
  assign _T_64576 = _T_64575[4:0]; // @[Modules.scala 43:47:@12128.4]
  assign _T_64577 = $signed(_T_64576); // @[Modules.scala 43:47:@12129.4]
  assign _T_64578 = $signed(io_in_310) + $signed(io_in_311); // @[Modules.scala 37:46:@12131.4]
  assign _T_64579 = _T_64578[4:0]; // @[Modules.scala 37:46:@12132.4]
  assign _T_64580 = $signed(_T_64579); // @[Modules.scala 37:46:@12133.4]
  assign _T_64592 = $signed(_T_55208) - $signed(io_in_315); // @[Modules.scala 46:47:@12145.4]
  assign _T_64593 = _T_64592[4:0]; // @[Modules.scala 46:47:@12146.4]
  assign _T_64594 = $signed(_T_64593); // @[Modules.scala 46:47:@12147.4]
  assign _T_64603 = $signed(5'sh0) - $signed(io_in_318); // @[Modules.scala 46:37:@12156.4]
  assign _T_64604 = _T_64603[4:0]; // @[Modules.scala 46:37:@12157.4]
  assign _T_64605 = $signed(_T_64604); // @[Modules.scala 46:37:@12158.4]
  assign _T_64606 = $signed(_T_64605) - $signed(io_in_319); // @[Modules.scala 46:47:@12159.4]
  assign _T_64607 = _T_64606[4:0]; // @[Modules.scala 46:47:@12160.4]
  assign _T_64608 = $signed(_T_64607); // @[Modules.scala 46:47:@12161.4]
  assign _T_64658 = $signed(io_in_334) - $signed(io_in_335); // @[Modules.scala 40:46:@12212.4]
  assign _T_64659 = _T_64658[4:0]; // @[Modules.scala 40:46:@12213.4]
  assign _T_64660 = $signed(_T_64659); // @[Modules.scala 40:46:@12214.4]
  assign _T_64662 = $signed(5'sh0) - $signed(io_in_336); // @[Modules.scala 43:37:@12216.4]
  assign _T_64663 = _T_64662[4:0]; // @[Modules.scala 43:37:@12217.4]
  assign _T_64664 = $signed(_T_64663); // @[Modules.scala 43:37:@12218.4]
  assign _T_64665 = $signed(_T_64664) + $signed(io_in_337); // @[Modules.scala 43:47:@12219.4]
  assign _T_64666 = _T_64665[4:0]; // @[Modules.scala 43:47:@12220.4]
  assign _T_64667 = $signed(_T_64666); // @[Modules.scala 43:47:@12221.4]
  assign _T_64668 = $signed(io_in_338) - $signed(io_in_339); // @[Modules.scala 40:46:@12223.4]
  assign _T_64669 = _T_64668[4:0]; // @[Modules.scala 40:46:@12224.4]
  assign _T_64670 = $signed(_T_64669); // @[Modules.scala 40:46:@12225.4]
  assign _T_64675 = $signed(_T_55283) - $signed(io_in_341); // @[Modules.scala 46:47:@12230.4]
  assign _T_64676 = _T_64675[4:0]; // @[Modules.scala 46:47:@12231.4]
  assign _T_64677 = $signed(_T_64676); // @[Modules.scala 46:47:@12232.4]
  assign _T_64679 = $signed(5'sh0) - $signed(io_in_342); // @[Modules.scala 46:37:@12234.4]
  assign _T_64680 = _T_64679[4:0]; // @[Modules.scala 46:37:@12235.4]
  assign _T_64681 = $signed(_T_64680); // @[Modules.scala 46:37:@12236.4]
  assign _T_64682 = $signed(_T_64681) - $signed(io_in_343); // @[Modules.scala 46:47:@12237.4]
  assign _T_64683 = _T_64682[4:0]; // @[Modules.scala 46:47:@12238.4]
  assign _T_64684 = $signed(_T_64683); // @[Modules.scala 46:47:@12239.4]
  assign _T_64686 = $signed(5'sh0) - $signed(io_in_344); // @[Modules.scala 46:37:@12241.4]
  assign _T_64687 = _T_64686[4:0]; // @[Modules.scala 46:37:@12242.4]
  assign _T_64688 = $signed(_T_64687); // @[Modules.scala 46:37:@12243.4]
  assign _T_64689 = $signed(_T_64688) - $signed(io_in_345); // @[Modules.scala 46:47:@12244.4]
  assign _T_64690 = _T_64689[4:0]; // @[Modules.scala 46:47:@12245.4]
  assign _T_64691 = $signed(_T_64690); // @[Modules.scala 46:47:@12246.4]
  assign _T_64693 = $signed(5'sh0) - $signed(io_in_346); // @[Modules.scala 46:37:@12248.4]
  assign _T_64694 = _T_64693[4:0]; // @[Modules.scala 46:37:@12249.4]
  assign _T_64695 = $signed(_T_64694); // @[Modules.scala 46:37:@12250.4]
  assign _T_64696 = $signed(_T_64695) - $signed(io_in_347); // @[Modules.scala 46:47:@12251.4]
  assign _T_64697 = _T_64696[4:0]; // @[Modules.scala 46:47:@12252.4]
  assign _T_64698 = $signed(_T_64697); // @[Modules.scala 46:47:@12253.4]
  assign _T_64700 = $signed(5'sh0) - $signed(io_in_348); // @[Modules.scala 46:37:@12255.4]
  assign _T_64701 = _T_64700[4:0]; // @[Modules.scala 46:37:@12256.4]
  assign _T_64702 = $signed(_T_64701); // @[Modules.scala 46:37:@12257.4]
  assign _T_64703 = $signed(_T_64702) - $signed(io_in_349); // @[Modules.scala 46:47:@12258.4]
  assign _T_64704 = _T_64703[4:0]; // @[Modules.scala 46:47:@12259.4]
  assign _T_64705 = $signed(_T_64704); // @[Modules.scala 46:47:@12260.4]
  assign _T_64755 = $signed(_T_55331) + $signed(io_in_365); // @[Modules.scala 43:47:@12311.4]
  assign _T_64756 = _T_64755[4:0]; // @[Modules.scala 43:47:@12312.4]
  assign _T_64757 = $signed(_T_64756); // @[Modules.scala 43:47:@12313.4]
  assign _T_64758 = $signed(io_in_366) - $signed(io_in_367); // @[Modules.scala 40:46:@12315.4]
  assign _T_64759 = _T_64758[4:0]; // @[Modules.scala 40:46:@12316.4]
  assign _T_64760 = $signed(_T_64759); // @[Modules.scala 40:46:@12317.4]
  assign _T_64765 = $signed(_T_58462) - $signed(io_in_369); // @[Modules.scala 46:47:@12322.4]
  assign _T_64766 = _T_64765[4:0]; // @[Modules.scala 46:47:@12323.4]
  assign _T_64767 = $signed(_T_64766); // @[Modules.scala 46:47:@12324.4]
  assign _T_64769 = $signed(5'sh0) - $signed(io_in_370); // @[Modules.scala 46:37:@12326.4]
  assign _T_64770 = _T_64769[4:0]; // @[Modules.scala 46:37:@12327.4]
  assign _T_64771 = $signed(_T_64770); // @[Modules.scala 46:37:@12328.4]
  assign _T_64772 = $signed(_T_64771) - $signed(io_in_371); // @[Modules.scala 46:47:@12329.4]
  assign _T_64773 = _T_64772[4:0]; // @[Modules.scala 46:47:@12330.4]
  assign _T_64774 = $signed(_T_64773); // @[Modules.scala 46:47:@12331.4]
  assign _T_64776 = $signed(5'sh0) - $signed(io_in_372); // @[Modules.scala 46:37:@12333.4]
  assign _T_64777 = _T_64776[4:0]; // @[Modules.scala 46:37:@12334.4]
  assign _T_64778 = $signed(_T_64777); // @[Modules.scala 46:37:@12335.4]
  assign _T_64779 = $signed(_T_64778) - $signed(io_in_373); // @[Modules.scala 46:47:@12336.4]
  assign _T_64780 = _T_64779[4:0]; // @[Modules.scala 46:47:@12337.4]
  assign _T_64781 = $signed(_T_64780); // @[Modules.scala 46:47:@12338.4]
  assign _T_64783 = $signed(5'sh0) - $signed(io_in_374); // @[Modules.scala 43:37:@12340.4]
  assign _T_64784 = _T_64783[4:0]; // @[Modules.scala 43:37:@12341.4]
  assign _T_64785 = $signed(_T_64784); // @[Modules.scala 43:37:@12342.4]
  assign _T_64786 = $signed(_T_64785) + $signed(io_in_375); // @[Modules.scala 43:47:@12343.4]
  assign _T_64787 = _T_64786[4:0]; // @[Modules.scala 43:47:@12344.4]
  assign _T_64788 = $signed(_T_64787); // @[Modules.scala 43:47:@12345.4]
  assign _T_64790 = $signed(5'sh0) - $signed(io_in_376); // @[Modules.scala 46:37:@12347.4]
  assign _T_64791 = _T_64790[4:0]; // @[Modules.scala 46:37:@12348.4]
  assign _T_64792 = $signed(_T_64791); // @[Modules.scala 46:37:@12349.4]
  assign _T_64793 = $signed(_T_64792) - $signed(io_in_377); // @[Modules.scala 46:47:@12350.4]
  assign _T_64794 = _T_64793[4:0]; // @[Modules.scala 46:47:@12351.4]
  assign _T_64795 = $signed(_T_64794); // @[Modules.scala 46:47:@12352.4]
  assign _T_64807 = $signed(_T_58488) + $signed(io_in_381); // @[Modules.scala 43:47:@12364.4]
  assign _T_64808 = _T_64807[4:0]; // @[Modules.scala 43:47:@12365.4]
  assign _T_64809 = $signed(_T_64808); // @[Modules.scala 43:47:@12366.4]
  assign _T_64821 = $signed(_T_55369) - $signed(io_in_385); // @[Modules.scala 46:47:@12378.4]
  assign _T_64822 = _T_64821[4:0]; // @[Modules.scala 46:47:@12379.4]
  assign _T_64823 = $signed(_T_64822); // @[Modules.scala 46:47:@12380.4]
  assign _T_64838 = $signed(io_in_390) + $signed(io_in_391); // @[Modules.scala 37:46:@12396.4]
  assign _T_64839 = _T_64838[4:0]; // @[Modules.scala 37:46:@12397.4]
  assign _T_64840 = $signed(_T_64839); // @[Modules.scala 37:46:@12398.4]
  assign _T_64844 = $signed(io_in_394) - $signed(io_in_395); // @[Modules.scala 40:46:@12404.4]
  assign _T_64845 = _T_64844[4:0]; // @[Modules.scala 40:46:@12405.4]
  assign _T_64846 = $signed(_T_64845); // @[Modules.scala 40:46:@12406.4]
  assign _T_64851 = $signed(_T_58532) - $signed(io_in_397); // @[Modules.scala 46:47:@12411.4]
  assign _T_64852 = _T_64851[4:0]; // @[Modules.scala 46:47:@12412.4]
  assign _T_64853 = $signed(_T_64852); // @[Modules.scala 46:47:@12413.4]
  assign _T_64855 = $signed(5'sh0) - $signed(io_in_398); // @[Modules.scala 46:37:@12415.4]
  assign _T_64856 = _T_64855[4:0]; // @[Modules.scala 46:37:@12416.4]
  assign _T_64857 = $signed(_T_64856); // @[Modules.scala 46:37:@12417.4]
  assign _T_64858 = $signed(_T_64857) - $signed(io_in_399); // @[Modules.scala 46:47:@12418.4]
  assign _T_64859 = _T_64858[4:0]; // @[Modules.scala 46:47:@12419.4]
  assign _T_64860 = $signed(_T_64859); // @[Modules.scala 46:47:@12420.4]
  assign _T_64862 = $signed(5'sh0) - $signed(io_in_400); // @[Modules.scala 43:37:@12422.4]
  assign _T_64863 = _T_64862[4:0]; // @[Modules.scala 43:37:@12423.4]
  assign _T_64864 = $signed(_T_64863); // @[Modules.scala 43:37:@12424.4]
  assign _T_64865 = $signed(_T_64864) + $signed(io_in_401); // @[Modules.scala 43:47:@12425.4]
  assign _T_64866 = _T_64865[4:0]; // @[Modules.scala 43:47:@12426.4]
  assign _T_64867 = $signed(_T_64866); // @[Modules.scala 43:47:@12427.4]
  assign _T_64868 = $signed(io_in_402) - $signed(io_in_403); // @[Modules.scala 40:46:@12429.4]
  assign _T_64869 = _T_64868[4:0]; // @[Modules.scala 40:46:@12430.4]
  assign _T_64870 = $signed(_T_64869); // @[Modules.scala 40:46:@12431.4]
  assign _T_64872 = $signed(5'sh0) - $signed(io_in_404); // @[Modules.scala 46:37:@12433.4]
  assign _T_64873 = _T_64872[4:0]; // @[Modules.scala 46:37:@12434.4]
  assign _T_64874 = $signed(_T_64873); // @[Modules.scala 46:37:@12435.4]
  assign _T_64875 = $signed(_T_64874) - $signed(io_in_405); // @[Modules.scala 46:47:@12436.4]
  assign _T_64876 = _T_64875[4:0]; // @[Modules.scala 46:47:@12437.4]
  assign _T_64877 = $signed(_T_64876); // @[Modules.scala 46:47:@12438.4]
  assign _T_64886 = $signed(5'sh0) - $signed(io_in_408); // @[Modules.scala 46:37:@12447.4]
  assign _T_64887 = _T_64886[4:0]; // @[Modules.scala 46:37:@12448.4]
  assign _T_64888 = $signed(_T_64887); // @[Modules.scala 46:37:@12449.4]
  assign _T_64889 = $signed(_T_64888) - $signed(io_in_409); // @[Modules.scala 46:47:@12450.4]
  assign _T_64890 = _T_64889[4:0]; // @[Modules.scala 46:47:@12451.4]
  assign _T_64891 = $signed(_T_64890); // @[Modules.scala 46:47:@12452.4]
  assign _T_64892 = $signed(io_in_410) - $signed(io_in_411); // @[Modules.scala 40:46:@12454.4]
  assign _T_64893 = _T_64892[4:0]; // @[Modules.scala 40:46:@12455.4]
  assign _T_64894 = $signed(_T_64893); // @[Modules.scala 40:46:@12456.4]
  assign _T_64896 = $signed(5'sh0) - $signed(io_in_412); // @[Modules.scala 46:37:@12458.4]
  assign _T_64897 = _T_64896[4:0]; // @[Modules.scala 46:37:@12459.4]
  assign _T_64898 = $signed(_T_64897); // @[Modules.scala 46:37:@12460.4]
  assign _T_64899 = $signed(_T_64898) - $signed(io_in_413); // @[Modules.scala 46:47:@12461.4]
  assign _T_64900 = _T_64899[4:0]; // @[Modules.scala 46:47:@12462.4]
  assign _T_64901 = $signed(_T_64900); // @[Modules.scala 46:47:@12463.4]
  assign _T_64903 = $signed(5'sh0) - $signed(io_in_414); // @[Modules.scala 46:37:@12465.4]
  assign _T_64904 = _T_64903[4:0]; // @[Modules.scala 46:37:@12466.4]
  assign _T_64905 = $signed(_T_64904); // @[Modules.scala 46:37:@12467.4]
  assign _T_64906 = $signed(_T_64905) - $signed(io_in_415); // @[Modules.scala 46:47:@12468.4]
  assign _T_64907 = _T_64906[4:0]; // @[Modules.scala 46:47:@12469.4]
  assign _T_64908 = $signed(_T_64907); // @[Modules.scala 46:47:@12470.4]
  assign _T_64913 = $signed(_T_61727) + $signed(io_in_417); // @[Modules.scala 43:47:@12475.4]
  assign _T_64914 = _T_64913[4:0]; // @[Modules.scala 43:47:@12476.4]
  assign _T_64915 = $signed(_T_64914); // @[Modules.scala 43:47:@12477.4]
  assign _T_64916 = $signed(io_in_418) + $signed(io_in_419); // @[Modules.scala 37:46:@12479.4]
  assign _T_64917 = _T_64916[4:0]; // @[Modules.scala 37:46:@12480.4]
  assign _T_64918 = $signed(_T_64917); // @[Modules.scala 37:46:@12481.4]
  assign _T_64919 = $signed(io_in_420) - $signed(io_in_421); // @[Modules.scala 40:46:@12483.4]
  assign _T_64920 = _T_64919[4:0]; // @[Modules.scala 40:46:@12484.4]
  assign _T_64921 = $signed(_T_64920); // @[Modules.scala 40:46:@12485.4]
  assign _T_64925 = $signed(io_in_424) + $signed(io_in_425); // @[Modules.scala 37:46:@12491.4]
  assign _T_64926 = _T_64925[4:0]; // @[Modules.scala 37:46:@12492.4]
  assign _T_64927 = $signed(_T_64926); // @[Modules.scala 37:46:@12493.4]
  assign _T_64932 = $signed(_T_58601) + $signed(io_in_427); // @[Modules.scala 43:47:@12498.4]
  assign _T_64933 = _T_64932[4:0]; // @[Modules.scala 43:47:@12499.4]
  assign _T_64934 = $signed(_T_64933); // @[Modules.scala 43:47:@12500.4]
  assign _T_64977 = $signed(_T_61791) + $signed(io_in_441); // @[Modules.scala 43:47:@12544.4]
  assign _T_64978 = _T_64977[4:0]; // @[Modules.scala 43:47:@12545.4]
  assign _T_64979 = $signed(_T_64978); // @[Modules.scala 43:47:@12546.4]
  assign _T_64984 = $signed(_T_55488) - $signed(io_in_443); // @[Modules.scala 46:47:@12551.4]
  assign _T_64985 = _T_64984[4:0]; // @[Modules.scala 46:47:@12552.4]
  assign _T_64986 = $signed(_T_64985); // @[Modules.scala 46:47:@12553.4]
  assign _T_64987 = $signed(io_in_444) + $signed(io_in_445); // @[Modules.scala 37:46:@12555.4]
  assign _T_64988 = _T_64987[4:0]; // @[Modules.scala 37:46:@12556.4]
  assign _T_64989 = $signed(_T_64988); // @[Modules.scala 37:46:@12557.4]
  assign _T_64990 = $signed(io_in_446) + $signed(io_in_447); // @[Modules.scala 37:46:@12559.4]
  assign _T_64991 = _T_64990[4:0]; // @[Modules.scala 37:46:@12560.4]
  assign _T_64992 = $signed(_T_64991); // @[Modules.scala 37:46:@12561.4]
  assign _T_64993 = $signed(io_in_448) - $signed(io_in_449); // @[Modules.scala 40:46:@12563.4]
  assign _T_64994 = _T_64993[4:0]; // @[Modules.scala 40:46:@12564.4]
  assign _T_64995 = $signed(_T_64994); // @[Modules.scala 40:46:@12565.4]
  assign _T_64999 = $signed(io_in_452) + $signed(io_in_453); // @[Modules.scala 37:46:@12571.4]
  assign _T_65000 = _T_64999[4:0]; // @[Modules.scala 37:46:@12572.4]
  assign _T_65001 = $signed(_T_65000); // @[Modules.scala 37:46:@12573.4]
  assign _T_65009 = $signed(_T_58682) - $signed(io_in_457); // @[Modules.scala 46:47:@12582.4]
  assign _T_65010 = _T_65009[4:0]; // @[Modules.scala 46:47:@12583.4]
  assign _T_65011 = $signed(_T_65010); // @[Modules.scala 46:47:@12584.4]
  assign _T_65049 = $signed(io_in_472) + $signed(io_in_473); // @[Modules.scala 37:46:@12626.4]
  assign _T_65050 = _T_65049[4:0]; // @[Modules.scala 37:46:@12627.4]
  assign _T_65051 = $signed(_T_65050); // @[Modules.scala 37:46:@12628.4]
  assign _T_65052 = $signed(io_in_474) + $signed(io_in_475); // @[Modules.scala 37:46:@12630.4]
  assign _T_65053 = _T_65052[4:0]; // @[Modules.scala 37:46:@12631.4]
  assign _T_65054 = $signed(_T_65053); // @[Modules.scala 37:46:@12632.4]
  assign _T_65065 = $signed(io_in_480) + $signed(io_in_481); // @[Modules.scala 37:46:@12645.4]
  assign _T_65066 = _T_65065[4:0]; // @[Modules.scala 37:46:@12646.4]
  assign _T_65067 = $signed(_T_65066); // @[Modules.scala 37:46:@12647.4]
  assign _T_65068 = $signed(io_in_482) - $signed(io_in_483); // @[Modules.scala 40:46:@12649.4]
  assign _T_65069 = _T_65068[4:0]; // @[Modules.scala 40:46:@12650.4]
  assign _T_65070 = $signed(_T_65069); // @[Modules.scala 40:46:@12651.4]
  assign _T_65103 = $signed(_T_58784) + $signed(io_in_493); // @[Modules.scala 43:47:@12684.4]
  assign _T_65104 = _T_65103[4:0]; // @[Modules.scala 43:47:@12685.4]
  assign _T_65105 = $signed(_T_65104); // @[Modules.scala 43:47:@12686.4]
  assign _T_65115 = $signed(io_in_500) + $signed(io_in_501); // @[Modules.scala 37:46:@12700.4]
  assign _T_65116 = _T_65115[4:0]; // @[Modules.scala 37:46:@12701.4]
  assign _T_65117 = $signed(_T_65116); // @[Modules.scala 37:46:@12702.4]
  assign _T_65118 = $signed(io_in_502) + $signed(io_in_503); // @[Modules.scala 37:46:@12704.4]
  assign _T_65119 = _T_65118[4:0]; // @[Modules.scala 37:46:@12705.4]
  assign _T_65120 = $signed(_T_65119); // @[Modules.scala 37:46:@12706.4]
  assign _T_65121 = $signed(io_in_504) - $signed(io_in_505); // @[Modules.scala 40:46:@12708.4]
  assign _T_65122 = _T_65121[4:0]; // @[Modules.scala 40:46:@12709.4]
  assign _T_65123 = $signed(_T_65122); // @[Modules.scala 40:46:@12710.4]
  assign _T_65127 = $signed(io_in_508) + $signed(io_in_509); // @[Modules.scala 37:46:@12716.4]
  assign _T_65128 = _T_65127[4:0]; // @[Modules.scala 37:46:@12717.4]
  assign _T_65129 = $signed(_T_65128); // @[Modules.scala 37:46:@12718.4]
  assign _T_65141 = $signed(5'sh0) - $signed(io_in_514); // @[Modules.scala 46:37:@12731.4]
  assign _T_65142 = _T_65141[4:0]; // @[Modules.scala 46:37:@12732.4]
  assign _T_65143 = $signed(_T_65142); // @[Modules.scala 46:37:@12733.4]
  assign _T_65144 = $signed(_T_65143) - $signed(io_in_515); // @[Modules.scala 46:47:@12734.4]
  assign _T_65145 = _T_65144[4:0]; // @[Modules.scala 46:47:@12735.4]
  assign _T_65146 = $signed(_T_65145); // @[Modules.scala 46:47:@12736.4]
  assign _T_65180 = $signed(io_in_530) + $signed(io_in_531); // @[Modules.scala 37:46:@12775.4]
  assign _T_65181 = _T_65180[4:0]; // @[Modules.scala 37:46:@12776.4]
  assign _T_65182 = $signed(_T_65181); // @[Modules.scala 37:46:@12777.4]
  assign _T_65195 = $signed(io_in_540) - $signed(io_in_541); // @[Modules.scala 40:46:@12795.4]
  assign _T_65196 = _T_65195[4:0]; // @[Modules.scala 40:46:@12796.4]
  assign _T_65197 = $signed(_T_65196); // @[Modules.scala 40:46:@12797.4]
  assign _T_65202 = $signed(_T_55742) - $signed(io_in_543); // @[Modules.scala 46:47:@12802.4]
  assign _T_65203 = _T_65202[4:0]; // @[Modules.scala 46:47:@12803.4]
  assign _T_65204 = $signed(_T_65203); // @[Modules.scala 46:47:@12804.4]
  assign _T_65212 = $signed(io_in_546) - $signed(io_in_547); // @[Modules.scala 40:46:@12813.4]
  assign _T_65213 = _T_65212[4:0]; // @[Modules.scala 40:46:@12814.4]
  assign _T_65214 = $signed(_T_65213); // @[Modules.scala 40:46:@12815.4]
  assign _T_65226 = $signed(_T_62112) - $signed(io_in_551); // @[Modules.scala 46:47:@12827.4]
  assign _T_65227 = _T_65226[4:0]; // @[Modules.scala 46:47:@12828.4]
  assign _T_65228 = $signed(_T_65227); // @[Modules.scala 46:47:@12829.4]
  assign _T_65232 = $signed(io_in_554) + $signed(io_in_555); // @[Modules.scala 37:46:@12835.4]
  assign _T_65233 = _T_65232[4:0]; // @[Modules.scala 37:46:@12836.4]
  assign _T_65234 = $signed(_T_65233); // @[Modules.scala 37:46:@12837.4]
  assign _T_65235 = $signed(io_in_556) + $signed(io_in_557); // @[Modules.scala 37:46:@12839.4]
  assign _T_65236 = _T_65235[4:0]; // @[Modules.scala 37:46:@12840.4]
  assign _T_65237 = $signed(_T_65236); // @[Modules.scala 37:46:@12841.4]
  assign _T_65238 = $signed(io_in_558) - $signed(io_in_559); // @[Modules.scala 40:46:@12843.4]
  assign _T_65239 = _T_65238[4:0]; // @[Modules.scala 40:46:@12844.4]
  assign _T_65240 = $signed(_T_65239); // @[Modules.scala 40:46:@12845.4]
  assign _T_65250 = $signed(io_in_566) + $signed(io_in_567); // @[Modules.scala 37:46:@12859.4]
  assign _T_65251 = _T_65250[4:0]; // @[Modules.scala 37:46:@12860.4]
  assign _T_65252 = $signed(_T_65251); // @[Modules.scala 37:46:@12861.4]
  assign _T_65259 = $signed(io_in_572) - $signed(io_in_573); // @[Modules.scala 40:46:@12871.4]
  assign _T_65260 = _T_65259[4:0]; // @[Modules.scala 40:46:@12872.4]
  assign _T_65261 = $signed(_T_65260); // @[Modules.scala 40:46:@12873.4]
  assign _T_65278 = $signed(io_in_582) + $signed(io_in_583); // @[Modules.scala 37:46:@12894.4]
  assign _T_65279 = _T_65278[4:0]; // @[Modules.scala 37:46:@12895.4]
  assign _T_65280 = $signed(_T_65279); // @[Modules.scala 37:46:@12896.4]
  assign _T_65284 = $signed(io_in_586) + $signed(io_in_587); // @[Modules.scala 37:46:@12902.4]
  assign _T_65285 = _T_65284[4:0]; // @[Modules.scala 37:46:@12903.4]
  assign _T_65286 = $signed(_T_65285); // @[Modules.scala 37:46:@12904.4]
  assign _T_65300 = $signed(io_in_594) + $signed(io_in_595); // @[Modules.scala 37:46:@12921.4]
  assign _T_65301 = _T_65300[4:0]; // @[Modules.scala 37:46:@12922.4]
  assign _T_65302 = $signed(_T_65301); // @[Modules.scala 37:46:@12923.4]
  assign _T_65321 = $signed(5'sh0) - $signed(io_in_602); // @[Modules.scala 46:37:@12943.4]
  assign _T_65322 = _T_65321[4:0]; // @[Modules.scala 46:37:@12944.4]
  assign _T_65323 = $signed(_T_65322); // @[Modules.scala 46:37:@12945.4]
  assign _T_65324 = $signed(_T_65323) - $signed(io_in_603); // @[Modules.scala 46:47:@12946.4]
  assign _T_65325 = _T_65324[4:0]; // @[Modules.scala 46:47:@12947.4]
  assign _T_65326 = $signed(_T_65325); // @[Modules.scala 46:47:@12948.4]
  assign _T_65341 = $signed(_T_55929) + $signed(io_in_609); // @[Modules.scala 43:47:@12964.4]
  assign _T_65342 = _T_65341[4:0]; // @[Modules.scala 43:47:@12965.4]
  assign _T_65343 = $signed(_T_65342); // @[Modules.scala 43:47:@12966.4]
  assign _T_65344 = $signed(io_in_610) + $signed(io_in_611); // @[Modules.scala 37:46:@12968.4]
  assign _T_65345 = _T_65344[4:0]; // @[Modules.scala 37:46:@12969.4]
  assign _T_65346 = $signed(_T_65345); // @[Modules.scala 37:46:@12970.4]
  assign _T_65350 = $signed(io_in_614) - $signed(io_in_615); // @[Modules.scala 40:46:@12976.4]
  assign _T_65351 = _T_65350[4:0]; // @[Modules.scala 40:46:@12977.4]
  assign _T_65352 = $signed(_T_65351); // @[Modules.scala 40:46:@12978.4]
  assign _T_65363 = $signed(io_in_620) + $signed(io_in_621); // @[Modules.scala 37:46:@12991.4]
  assign _T_65364 = _T_65363[4:0]; // @[Modules.scala 37:46:@12992.4]
  assign _T_65365 = $signed(_T_65364); // @[Modules.scala 37:46:@12993.4]
  assign _T_65380 = $signed(_T_55984) + $signed(io_in_627); // @[Modules.scala 43:47:@13009.4]
  assign _T_65381 = _T_65380[4:0]; // @[Modules.scala 43:47:@13010.4]
  assign _T_65382 = $signed(_T_65381); // @[Modules.scala 43:47:@13011.4]
  assign _T_65386 = $signed(io_in_630) - $signed(io_in_631); // @[Modules.scala 40:46:@13017.4]
  assign _T_65387 = _T_65386[4:0]; // @[Modules.scala 40:46:@13018.4]
  assign _T_65388 = $signed(_T_65387); // @[Modules.scala 40:46:@13019.4]
  assign _T_65389 = $signed(io_in_632) - $signed(io_in_633); // @[Modules.scala 40:46:@13021.4]
  assign _T_65390 = _T_65389[4:0]; // @[Modules.scala 40:46:@13022.4]
  assign _T_65391 = $signed(_T_65390); // @[Modules.scala 40:46:@13023.4]
  assign _T_65396 = $signed(_T_56012) + $signed(io_in_635); // @[Modules.scala 43:47:@13028.4]
  assign _T_65397 = _T_65396[4:0]; // @[Modules.scala 43:47:@13029.4]
  assign _T_65398 = $signed(_T_65397); // @[Modules.scala 43:47:@13030.4]
  assign _T_65402 = $signed(io_in_638) + $signed(io_in_639); // @[Modules.scala 37:46:@13036.4]
  assign _T_65403 = _T_65402[4:0]; // @[Modules.scala 37:46:@13037.4]
  assign _T_65404 = $signed(_T_65403); // @[Modules.scala 37:46:@13038.4]
  assign _T_65408 = $signed(io_in_642) - $signed(io_in_643); // @[Modules.scala 40:46:@13044.4]
  assign _T_65409 = _T_65408[4:0]; // @[Modules.scala 40:46:@13045.4]
  assign _T_65410 = $signed(_T_65409); // @[Modules.scala 40:46:@13046.4]
  assign _T_65424 = $signed(_T_56060) + $signed(io_in_651); // @[Modules.scala 43:47:@13063.4]
  assign _T_65425 = _T_65424[4:0]; // @[Modules.scala 43:47:@13064.4]
  assign _T_65426 = $signed(_T_65425); // @[Modules.scala 43:47:@13065.4]
  assign _T_65431 = $signed(_T_56067) + $signed(io_in_653); // @[Modules.scala 43:47:@13070.4]
  assign _T_65432 = _T_65431[4:0]; // @[Modules.scala 43:47:@13071.4]
  assign _T_65433 = $signed(_T_65432); // @[Modules.scala 43:47:@13072.4]
  assign _T_65458 = $signed(_T_56102) - $signed(io_in_663); // @[Modules.scala 46:47:@13099.4]
  assign _T_65459 = _T_65458[4:0]; // @[Modules.scala 46:47:@13100.4]
  assign _T_65460 = $signed(_T_65459); // @[Modules.scala 46:47:@13101.4]
  assign _T_65468 = $signed(io_in_666) - $signed(io_in_667); // @[Modules.scala 40:46:@13110.4]
  assign _T_65469 = _T_65468[4:0]; // @[Modules.scala 40:46:@13111.4]
  assign _T_65470 = $signed(_T_65469); // @[Modules.scala 40:46:@13112.4]
  assign _T_65474 = $signed(io_in_670) - $signed(io_in_671); // @[Modules.scala 40:46:@13118.4]
  assign _T_65475 = _T_65474[4:0]; // @[Modules.scala 40:46:@13119.4]
  assign _T_65476 = $signed(_T_65475); // @[Modules.scala 40:46:@13120.4]
  assign _T_65477 = $signed(io_in_672) - $signed(io_in_673); // @[Modules.scala 40:46:@13122.4]
  assign _T_65478 = _T_65477[4:0]; // @[Modules.scala 40:46:@13123.4]
  assign _T_65479 = $signed(_T_65478); // @[Modules.scala 40:46:@13124.4]
  assign _T_65481 = $signed(5'sh0) - $signed(io_in_674); // @[Modules.scala 43:37:@13126.4]
  assign _T_65482 = _T_65481[4:0]; // @[Modules.scala 43:37:@13127.4]
  assign _T_65483 = $signed(_T_65482); // @[Modules.scala 43:37:@13128.4]
  assign _T_65484 = $signed(_T_65483) + $signed(io_in_675); // @[Modules.scala 43:47:@13129.4]
  assign _T_65485 = _T_65484[4:0]; // @[Modules.scala 43:47:@13130.4]
  assign _T_65486 = $signed(_T_65485); // @[Modules.scala 43:47:@13131.4]
  assign _T_65503 = $signed(_T_56147) + $signed(io_in_685); // @[Modules.scala 43:47:@13152.4]
  assign _T_65504 = _T_65503[4:0]; // @[Modules.scala 43:47:@13153.4]
  assign _T_65505 = $signed(_T_65504); // @[Modules.scala 43:47:@13154.4]
  assign _T_65506 = $signed(io_in_686) + $signed(io_in_687); // @[Modules.scala 37:46:@13156.4]
  assign _T_65507 = _T_65506[4:0]; // @[Modules.scala 37:46:@13157.4]
  assign _T_65508 = $signed(_T_65507); // @[Modules.scala 37:46:@13158.4]
  assign _T_65513 = $signed(_T_62467) - $signed(io_in_689); // @[Modules.scala 46:47:@13163.4]
  assign _T_65514 = _T_65513[4:0]; // @[Modules.scala 46:47:@13164.4]
  assign _T_65515 = $signed(_T_65514); // @[Modules.scala 46:47:@13165.4]
  assign _T_65517 = $signed(5'sh0) - $signed(io_in_690); // @[Modules.scala 46:37:@13167.4]
  assign _T_65518 = _T_65517[4:0]; // @[Modules.scala 46:37:@13168.4]
  assign _T_65519 = $signed(_T_65518); // @[Modules.scala 46:37:@13169.4]
  assign _T_65520 = $signed(_T_65519) - $signed(io_in_691); // @[Modules.scala 46:47:@13170.4]
  assign _T_65521 = _T_65520[4:0]; // @[Modules.scala 46:47:@13171.4]
  assign _T_65522 = $signed(_T_65521); // @[Modules.scala 46:47:@13172.4]
  assign _T_65534 = $signed(_T_59215) - $signed(io_in_695); // @[Modules.scala 46:47:@13184.4]
  assign _T_65535 = _T_65534[4:0]; // @[Modules.scala 46:47:@13185.4]
  assign _T_65536 = $signed(_T_65535); // @[Modules.scala 46:47:@13186.4]
  assign _T_65544 = $signed(io_in_698) + $signed(io_in_699); // @[Modules.scala 37:46:@13195.4]
  assign _T_65545 = _T_65544[4:0]; // @[Modules.scala 37:46:@13196.4]
  assign _T_65546 = $signed(_T_65545); // @[Modules.scala 37:46:@13197.4]
  assign _T_65555 = $signed(5'sh0) - $signed(io_in_702); // @[Modules.scala 43:37:@13206.4]
  assign _T_65556 = _T_65555[4:0]; // @[Modules.scala 43:37:@13207.4]
  assign _T_65557 = $signed(_T_65556); // @[Modules.scala 43:37:@13208.4]
  assign _T_65558 = $signed(_T_65557) + $signed(io_in_703); // @[Modules.scala 43:47:@13209.4]
  assign _T_65559 = _T_65558[4:0]; // @[Modules.scala 43:47:@13210.4]
  assign _T_65560 = $signed(_T_65559); // @[Modules.scala 43:47:@13211.4]
  assign _T_65570 = $signed(io_in_710) + $signed(io_in_711); // @[Modules.scala 37:46:@13225.4]
  assign _T_65571 = _T_65570[4:0]; // @[Modules.scala 37:46:@13226.4]
  assign _T_65572 = $signed(_T_65571); // @[Modules.scala 37:46:@13227.4]
  assign _T_65597 = $signed(5'sh0) - $signed(io_in_722); // @[Modules.scala 46:37:@13255.4]
  assign _T_65598 = _T_65597[4:0]; // @[Modules.scala 46:37:@13256.4]
  assign _T_65599 = $signed(_T_65598); // @[Modules.scala 46:37:@13257.4]
  assign _T_65600 = $signed(_T_65599) - $signed(io_in_723); // @[Modules.scala 46:47:@13258.4]
  assign _T_65601 = _T_65600[4:0]; // @[Modules.scala 46:47:@13259.4]
  assign _T_65602 = $signed(_T_65601); // @[Modules.scala 46:47:@13260.4]
  assign _T_65612 = $signed(io_in_730) - $signed(io_in_731); // @[Modules.scala 40:46:@13274.4]
  assign _T_65613 = _T_65612[4:0]; // @[Modules.scala 40:46:@13275.4]
  assign _T_65614 = $signed(_T_65613); // @[Modules.scala 40:46:@13276.4]
  assign _T_65621 = $signed(io_in_736) + $signed(io_in_737); // @[Modules.scala 37:46:@13286.4]
  assign _T_65622 = _T_65621[4:0]; // @[Modules.scala 37:46:@13287.4]
  assign _T_65623 = $signed(_T_65622); // @[Modules.scala 37:46:@13288.4]
  assign _T_65624 = $signed(io_in_738) + $signed(io_in_739); // @[Modules.scala 37:46:@13290.4]
  assign _T_65625 = _T_65624[4:0]; // @[Modules.scala 37:46:@13291.4]
  assign _T_65626 = $signed(_T_65625); // @[Modules.scala 37:46:@13292.4]
  assign _T_65627 = $signed(io_in_740) + $signed(io_in_741); // @[Modules.scala 37:46:@13294.4]
  assign _T_65628 = _T_65627[4:0]; // @[Modules.scala 37:46:@13295.4]
  assign _T_65629 = $signed(_T_65628); // @[Modules.scala 37:46:@13296.4]
  assign _T_65634 = $signed(_T_59347) + $signed(io_in_743); // @[Modules.scala 43:47:@13301.4]
  assign _T_65635 = _T_65634[4:0]; // @[Modules.scala 43:47:@13302.4]
  assign _T_65636 = $signed(_T_65635); // @[Modules.scala 43:47:@13303.4]
  assign _T_65637 = $signed(io_in_744) + $signed(io_in_745); // @[Modules.scala 37:46:@13305.4]
  assign _T_65638 = _T_65637[4:0]; // @[Modules.scala 37:46:@13306.4]
  assign _T_65639 = $signed(_T_65638); // @[Modules.scala 37:46:@13307.4]
  assign _T_65640 = $signed(io_in_746) + $signed(io_in_747); // @[Modules.scala 37:46:@13309.4]
  assign _T_65641 = _T_65640[4:0]; // @[Modules.scala 37:46:@13310.4]
  assign _T_65642 = $signed(_T_65641); // @[Modules.scala 37:46:@13311.4]
  assign _T_65644 = $signed(5'sh0) - $signed(io_in_748); // @[Modules.scala 46:37:@13313.4]
  assign _T_65645 = _T_65644[4:0]; // @[Modules.scala 46:37:@13314.4]
  assign _T_65646 = $signed(_T_65645); // @[Modules.scala 46:37:@13315.4]
  assign _T_65647 = $signed(_T_65646) - $signed(io_in_749); // @[Modules.scala 46:47:@13316.4]
  assign _T_65648 = _T_65647[4:0]; // @[Modules.scala 46:47:@13317.4]
  assign _T_65649 = $signed(_T_65648); // @[Modules.scala 46:47:@13318.4]
  assign _T_65653 = $signed(io_in_752) - $signed(io_in_753); // @[Modules.scala 40:46:@13324.4]
  assign _T_65654 = _T_65653[4:0]; // @[Modules.scala 40:46:@13325.4]
  assign _T_65655 = $signed(_T_65654); // @[Modules.scala 40:46:@13326.4]
  assign _T_65657 = $signed(5'sh0) - $signed(io_in_754); // @[Modules.scala 43:37:@13328.4]
  assign _T_65658 = _T_65657[4:0]; // @[Modules.scala 43:37:@13329.4]
  assign _T_65659 = $signed(_T_65658); // @[Modules.scala 43:37:@13330.4]
  assign _T_65660 = $signed(_T_65659) + $signed(io_in_755); // @[Modules.scala 43:47:@13331.4]
  assign _T_65661 = _T_65660[4:0]; // @[Modules.scala 43:47:@13332.4]
  assign _T_65662 = $signed(_T_65661); // @[Modules.scala 43:47:@13333.4]
  assign _T_65663 = $signed(io_in_756) + $signed(io_in_757); // @[Modules.scala 37:46:@13335.4]
  assign _T_65664 = _T_65663[4:0]; // @[Modules.scala 37:46:@13336.4]
  assign _T_65665 = $signed(_T_65664); // @[Modules.scala 37:46:@13337.4]
  assign _T_65679 = $signed(io_in_764) + $signed(io_in_765); // @[Modules.scala 37:46:@13354.4]
  assign _T_65680 = _T_65679[4:0]; // @[Modules.scala 37:46:@13355.4]
  assign _T_65681 = $signed(_T_65680); // @[Modules.scala 37:46:@13356.4]
  assign _T_65685 = $signed(io_in_768) + $signed(io_in_769); // @[Modules.scala 37:46:@13362.4]
  assign _T_65686 = _T_65685[4:0]; // @[Modules.scala 37:46:@13363.4]
  assign _T_65687 = $signed(_T_65686); // @[Modules.scala 37:46:@13364.4]
  assign _T_65688 = $signed(io_in_770) + $signed(io_in_771); // @[Modules.scala 37:46:@13366.4]
  assign _T_65689 = _T_65688[4:0]; // @[Modules.scala 37:46:@13367.4]
  assign _T_65690 = $signed(_T_65689); // @[Modules.scala 37:46:@13368.4]
  assign _T_65691 = $signed(io_in_772) + $signed(io_in_773); // @[Modules.scala 37:46:@13370.4]
  assign _T_65692 = _T_65691[4:0]; // @[Modules.scala 37:46:@13371.4]
  assign _T_65693 = $signed(_T_65692); // @[Modules.scala 37:46:@13372.4]
  assign _T_65694 = $signed(io_in_774) + $signed(io_in_775); // @[Modules.scala 37:46:@13374.4]
  assign _T_65695 = _T_65694[4:0]; // @[Modules.scala 37:46:@13375.4]
  assign _T_65696 = $signed(_T_65695); // @[Modules.scala 37:46:@13376.4]
  assign _T_65708 = $signed(_T_56360) + $signed(io_in_779); // @[Modules.scala 43:47:@13388.4]
  assign _T_65709 = _T_65708[4:0]; // @[Modules.scala 43:47:@13389.4]
  assign _T_65710 = $signed(_T_65709); // @[Modules.scala 43:47:@13390.4]
  assign buffer_3_0 = {{6{_T_63911[4]}},_T_63911}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_1 = {{6{_T_63914[4]}},_T_63914}; // @[Modules.scala 32:22:@8.4]
  assign _T_65717 = $signed(buffer_3_0) + $signed(buffer_3_1); // @[Modules.scala 50:57:@13400.4]
  assign _T_65718 = _T_65717[10:0]; // @[Modules.scala 50:57:@13401.4]
  assign buffer_3_392 = $signed(_T_65718); // @[Modules.scala 50:57:@13402.4]
  assign buffer_3_4 = {{6{_T_63927[4]}},_T_63927}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_5 = {{6{_T_63930[4]}},_T_63930}; // @[Modules.scala 32:22:@8.4]
  assign _T_65723 = $signed(buffer_3_4) + $signed(buffer_3_5); // @[Modules.scala 50:57:@13408.4]
  assign _T_65724 = _T_65723[10:0]; // @[Modules.scala 50:57:@13409.4]
  assign buffer_3_394 = $signed(_T_65724); // @[Modules.scala 50:57:@13410.4]
  assign _T_65729 = $signed(buffer_1_8) + $signed(buffer_0_9); // @[Modules.scala 50:57:@13416.4]
  assign _T_65730 = _T_65729[10:0]; // @[Modules.scala 50:57:@13417.4]
  assign buffer_3_396 = $signed(_T_65730); // @[Modules.scala 50:57:@13418.4]
  assign _T_65732 = $signed(buffer_2_10) + $signed(buffer_0_11); // @[Modules.scala 50:57:@13420.4]
  assign _T_65733 = _T_65732[10:0]; // @[Modules.scala 50:57:@13421.4]
  assign buffer_3_397 = $signed(_T_65733); // @[Modules.scala 50:57:@13422.4]
  assign buffer_3_12 = {{6{_T_63959[4]}},_T_63959}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_13 = {{6{_T_63962[4]}},_T_63962}; // @[Modules.scala 32:22:@8.4]
  assign _T_65735 = $signed(buffer_3_12) + $signed(buffer_3_13); // @[Modules.scala 50:57:@13424.4]
  assign _T_65736 = _T_65735[10:0]; // @[Modules.scala 50:57:@13425.4]
  assign buffer_3_398 = $signed(_T_65736); // @[Modules.scala 50:57:@13426.4]
  assign buffer_3_14 = {{6{_T_63965[4]}},_T_63965}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_15 = {{6{_T_63972[4]}},_T_63972}; // @[Modules.scala 32:22:@8.4]
  assign _T_65738 = $signed(buffer_3_14) + $signed(buffer_3_15); // @[Modules.scala 50:57:@13428.4]
  assign _T_65739 = _T_65738[10:0]; // @[Modules.scala 50:57:@13429.4]
  assign buffer_3_399 = $signed(_T_65739); // @[Modules.scala 50:57:@13430.4]
  assign buffer_3_16 = {{6{_T_63975[4]}},_T_63975}; // @[Modules.scala 32:22:@8.4]
  assign _T_65741 = $signed(buffer_3_16) + $signed(buffer_0_17); // @[Modules.scala 50:57:@13432.4]
  assign _T_65742 = _T_65741[10:0]; // @[Modules.scala 50:57:@13433.4]
  assign buffer_3_400 = $signed(_T_65742); // @[Modules.scala 50:57:@13434.4]
  assign _T_65750 = $signed(buffer_1_22) + $signed(buffer_0_23); // @[Modules.scala 50:57:@13444.4]
  assign _T_65751 = _T_65750[10:0]; // @[Modules.scala 50:57:@13445.4]
  assign buffer_3_403 = $signed(_T_65751); // @[Modules.scala 50:57:@13446.4]
  assign _T_65753 = $signed(buffer_0_24) + $signed(buffer_1_25); // @[Modules.scala 50:57:@13448.4]
  assign _T_65754 = _T_65753[10:0]; // @[Modules.scala 50:57:@13449.4]
  assign buffer_3_404 = $signed(_T_65754); // @[Modules.scala 50:57:@13450.4]
  assign buffer_3_26 = {{6{_T_64033[4]}},_T_64033}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_27 = {{6{_T_64040[4]}},_T_64040}; // @[Modules.scala 32:22:@8.4]
  assign _T_65756 = $signed(buffer_3_26) + $signed(buffer_3_27); // @[Modules.scala 50:57:@13452.4]
  assign _T_65757 = _T_65756[10:0]; // @[Modules.scala 50:57:@13453.4]
  assign buffer_3_405 = $signed(_T_65757); // @[Modules.scala 50:57:@13454.4]
  assign buffer_3_28 = {{6{_T_64047[4]}},_T_64047}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_29 = {{6{_T_64050[4]}},_T_64050}; // @[Modules.scala 32:22:@8.4]
  assign _T_65759 = $signed(buffer_3_28) + $signed(buffer_3_29); // @[Modules.scala 50:57:@13456.4]
  assign _T_65760 = _T_65759[10:0]; // @[Modules.scala 50:57:@13457.4]
  assign buffer_3_406 = $signed(_T_65760); // @[Modules.scala 50:57:@13458.4]
  assign buffer_3_30 = {{6{_T_64057[4]}},_T_64057}; // @[Modules.scala 32:22:@8.4]
  assign _T_65762 = $signed(buffer_3_30) + $signed(buffer_0_31); // @[Modules.scala 50:57:@13460.4]
  assign _T_65763 = _T_65762[10:0]; // @[Modules.scala 50:57:@13461.4]
  assign buffer_3_407 = $signed(_T_65763); // @[Modules.scala 50:57:@13462.4]
  assign buffer_3_32 = {{6{_T_64071[4]}},_T_64071}; // @[Modules.scala 32:22:@8.4]
  assign _T_65765 = $signed(buffer_3_32) + $signed(buffer_0_33); // @[Modules.scala 50:57:@13464.4]
  assign _T_65766 = _T_65765[10:0]; // @[Modules.scala 50:57:@13465.4]
  assign buffer_3_408 = $signed(_T_65766); // @[Modules.scala 50:57:@13466.4]
  assign buffer_3_37 = {{6{_T_64106[4]}},_T_64106}; // @[Modules.scala 32:22:@8.4]
  assign _T_65771 = $signed(buffer_0_36) + $signed(buffer_3_37); // @[Modules.scala 50:57:@13472.4]
  assign _T_65772 = _T_65771[10:0]; // @[Modules.scala 50:57:@13473.4]
  assign buffer_3_410 = $signed(_T_65772); // @[Modules.scala 50:57:@13474.4]
  assign buffer_3_38 = {{6{_T_64113[4]}},_T_64113}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_39 = {{6{_T_64120[4]}},_T_64120}; // @[Modules.scala 32:22:@8.4]
  assign _T_65774 = $signed(buffer_3_38) + $signed(buffer_3_39); // @[Modules.scala 50:57:@13476.4]
  assign _T_65775 = _T_65774[10:0]; // @[Modules.scala 50:57:@13477.4]
  assign buffer_3_411 = $signed(_T_65775); // @[Modules.scala 50:57:@13478.4]
  assign _T_65777 = $signed(buffer_1_40) + $signed(buffer_2_41); // @[Modules.scala 50:57:@13480.4]
  assign _T_65778 = _T_65777[10:0]; // @[Modules.scala 50:57:@13481.4]
  assign buffer_3_412 = $signed(_T_65778); // @[Modules.scala 50:57:@13482.4]
  assign buffer_3_43 = {{6{_T_64132[4]}},_T_64132}; // @[Modules.scala 32:22:@8.4]
  assign _T_65780 = $signed(buffer_0_42) + $signed(buffer_3_43); // @[Modules.scala 50:57:@13484.4]
  assign _T_65781 = _T_65780[10:0]; // @[Modules.scala 50:57:@13485.4]
  assign buffer_3_413 = $signed(_T_65781); // @[Modules.scala 50:57:@13486.4]
  assign buffer_3_44 = {{6{_T_64139[4]}},_T_64139}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_45 = {{6{_T_64146[4]}},_T_64146}; // @[Modules.scala 32:22:@8.4]
  assign _T_65783 = $signed(buffer_3_44) + $signed(buffer_3_45); // @[Modules.scala 50:57:@13488.4]
  assign _T_65784 = _T_65783[10:0]; // @[Modules.scala 50:57:@13489.4]
  assign buffer_3_414 = $signed(_T_65784); // @[Modules.scala 50:57:@13490.4]
  assign buffer_3_46 = {{6{_T_64153[4]}},_T_64153}; // @[Modules.scala 32:22:@8.4]
  assign _T_65786 = $signed(buffer_3_46) + $signed(buffer_0_47); // @[Modules.scala 50:57:@13492.4]
  assign _T_65787 = _T_65786[10:0]; // @[Modules.scala 50:57:@13493.4]
  assign buffer_3_415 = $signed(_T_65787); // @[Modules.scala 50:57:@13494.4]
  assign buffer_3_49 = {{6{_T_64162[4]}},_T_64162}; // @[Modules.scala 32:22:@8.4]
  assign _T_65789 = $signed(buffer_1_48) + $signed(buffer_3_49); // @[Modules.scala 50:57:@13496.4]
  assign _T_65790 = _T_65789[10:0]; // @[Modules.scala 50:57:@13497.4]
  assign buffer_3_416 = $signed(_T_65790); // @[Modules.scala 50:57:@13498.4]
  assign buffer_3_51 = {{6{_T_64172[4]}},_T_64172}; // @[Modules.scala 32:22:@8.4]
  assign _T_65792 = $signed(buffer_0_50) + $signed(buffer_3_51); // @[Modules.scala 50:57:@13500.4]
  assign _T_65793 = _T_65792[10:0]; // @[Modules.scala 50:57:@13501.4]
  assign buffer_3_417 = $signed(_T_65793); // @[Modules.scala 50:57:@13502.4]
  assign buffer_3_52 = {{6{_T_64179[4]}},_T_64179}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_53 = {{6{_T_64186[4]}},_T_64186}; // @[Modules.scala 32:22:@8.4]
  assign _T_65795 = $signed(buffer_3_52) + $signed(buffer_3_53); // @[Modules.scala 50:57:@13504.4]
  assign _T_65796 = _T_65795[10:0]; // @[Modules.scala 50:57:@13505.4]
  assign buffer_3_418 = $signed(_T_65796); // @[Modules.scala 50:57:@13506.4]
  assign buffer_3_54 = {{6{_T_64193[4]}},_T_64193}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_55 = {{6{_T_64196[4]}},_T_64196}; // @[Modules.scala 32:22:@8.4]
  assign _T_65798 = $signed(buffer_3_54) + $signed(buffer_3_55); // @[Modules.scala 50:57:@13508.4]
  assign _T_65799 = _T_65798[10:0]; // @[Modules.scala 50:57:@13509.4]
  assign buffer_3_419 = $signed(_T_65799); // @[Modules.scala 50:57:@13510.4]
  assign buffer_3_56 = {{6{_T_64199[4]}},_T_64199}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_57 = {{6{_T_64202[4]}},_T_64202}; // @[Modules.scala 32:22:@8.4]
  assign _T_65801 = $signed(buffer_3_56) + $signed(buffer_3_57); // @[Modules.scala 50:57:@13512.4]
  assign _T_65802 = _T_65801[10:0]; // @[Modules.scala 50:57:@13513.4]
  assign buffer_3_420 = $signed(_T_65802); // @[Modules.scala 50:57:@13514.4]
  assign _T_65804 = $signed(buffer_2_58) + $signed(buffer_0_59); // @[Modules.scala 50:57:@13516.4]
  assign _T_65805 = _T_65804[10:0]; // @[Modules.scala 50:57:@13517.4]
  assign buffer_3_421 = $signed(_T_65805); // @[Modules.scala 50:57:@13518.4]
  assign buffer_3_60 = {{6{_T_64215[4]}},_T_64215}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_61 = {{6{_T_64218[4]}},_T_64218}; // @[Modules.scala 32:22:@8.4]
  assign _T_65807 = $signed(buffer_3_60) + $signed(buffer_3_61); // @[Modules.scala 50:57:@13520.4]
  assign _T_65808 = _T_65807[10:0]; // @[Modules.scala 50:57:@13521.4]
  assign buffer_3_422 = $signed(_T_65808); // @[Modules.scala 50:57:@13522.4]
  assign buffer_3_62 = {{6{_T_64221[4]}},_T_64221}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_63 = {{6{_T_64224[4]}},_T_64224}; // @[Modules.scala 32:22:@8.4]
  assign _T_65810 = $signed(buffer_3_62) + $signed(buffer_3_63); // @[Modules.scala 50:57:@13524.4]
  assign _T_65811 = _T_65810[10:0]; // @[Modules.scala 50:57:@13525.4]
  assign buffer_3_423 = $signed(_T_65811); // @[Modules.scala 50:57:@13526.4]
  assign buffer_3_66 = {{6{_T_64237[4]}},_T_64237}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_67 = {{6{_T_64240[4]}},_T_64240}; // @[Modules.scala 32:22:@8.4]
  assign _T_65816 = $signed(buffer_3_66) + $signed(buffer_3_67); // @[Modules.scala 50:57:@13532.4]
  assign _T_65817 = _T_65816[10:0]; // @[Modules.scala 50:57:@13533.4]
  assign buffer_3_425 = $signed(_T_65817); // @[Modules.scala 50:57:@13534.4]
  assign buffer_3_69 = {{6{_T_64246[4]}},_T_64246}; // @[Modules.scala 32:22:@8.4]
  assign _T_65819 = $signed(buffer_1_68) + $signed(buffer_3_69); // @[Modules.scala 50:57:@13536.4]
  assign _T_65820 = _T_65819[10:0]; // @[Modules.scala 50:57:@13537.4]
  assign buffer_3_426 = $signed(_T_65820); // @[Modules.scala 50:57:@13538.4]
  assign _T_65822 = $signed(buffer_0_70) + $signed(buffer_1_71); // @[Modules.scala 50:57:@13540.4]
  assign _T_65823 = _T_65822[10:0]; // @[Modules.scala 50:57:@13541.4]
  assign buffer_3_427 = $signed(_T_65823); // @[Modules.scala 50:57:@13542.4]
  assign buffer_3_72 = {{6{_T_64263[4]}},_T_64263}; // @[Modules.scala 32:22:@8.4]
  assign _T_65825 = $signed(buffer_3_72) + $signed(buffer_0_73); // @[Modules.scala 50:57:@13544.4]
  assign _T_65826 = _T_65825[10:0]; // @[Modules.scala 50:57:@13545.4]
  assign buffer_3_428 = $signed(_T_65826); // @[Modules.scala 50:57:@13546.4]
  assign buffer_3_75 = {{6{_T_64272[4]}},_T_64272}; // @[Modules.scala 32:22:@8.4]
  assign _T_65828 = $signed(buffer_0_74) + $signed(buffer_3_75); // @[Modules.scala 50:57:@13548.4]
  assign _T_65829 = _T_65828[10:0]; // @[Modules.scala 50:57:@13549.4]
  assign buffer_3_429 = $signed(_T_65829); // @[Modules.scala 50:57:@13550.4]
  assign buffer_3_76 = {{6{_T_64279[4]}},_T_64279}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_77 = {{6{_T_64282[4]}},_T_64282}; // @[Modules.scala 32:22:@8.4]
  assign _T_65831 = $signed(buffer_3_76) + $signed(buffer_3_77); // @[Modules.scala 50:57:@13552.4]
  assign _T_65832 = _T_65831[10:0]; // @[Modules.scala 50:57:@13553.4]
  assign buffer_3_430 = $signed(_T_65832); // @[Modules.scala 50:57:@13554.4]
  assign buffer_3_79 = {{6{_T_64288[4]}},_T_64288}; // @[Modules.scala 32:22:@8.4]
  assign _T_65834 = $signed(buffer_1_78) + $signed(buffer_3_79); // @[Modules.scala 50:57:@13556.4]
  assign _T_65835 = _T_65834[10:0]; // @[Modules.scala 50:57:@13557.4]
  assign buffer_3_431 = $signed(_T_65835); // @[Modules.scala 50:57:@13558.4]
  assign buffer_3_86 = {{6{_T_64313[4]}},_T_64313}; // @[Modules.scala 32:22:@8.4]
  assign _T_65846 = $signed(buffer_3_86) + $signed(buffer_1_87); // @[Modules.scala 50:57:@13572.4]
  assign _T_65847 = _T_65846[10:0]; // @[Modules.scala 50:57:@13573.4]
  assign buffer_3_435 = $signed(_T_65847); // @[Modules.scala 50:57:@13574.4]
  assign buffer_3_89 = {{6{_T_64322[4]}},_T_64322}; // @[Modules.scala 32:22:@8.4]
  assign _T_65849 = $signed(buffer_1_88) + $signed(buffer_3_89); // @[Modules.scala 50:57:@13576.4]
  assign _T_65850 = _T_65849[10:0]; // @[Modules.scala 50:57:@13577.4]
  assign buffer_3_436 = $signed(_T_65850); // @[Modules.scala 50:57:@13578.4]
  assign buffer_3_90 = {{6{_T_64325[4]}},_T_64325}; // @[Modules.scala 32:22:@8.4]
  assign _T_65852 = $signed(buffer_3_90) + $signed(buffer_0_91); // @[Modules.scala 50:57:@13580.4]
  assign _T_65853 = _T_65852[10:0]; // @[Modules.scala 50:57:@13581.4]
  assign buffer_3_437 = $signed(_T_65853); // @[Modules.scala 50:57:@13582.4]
  assign buffer_3_92 = {{6{_T_64335[4]}},_T_64335}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_93 = {{6{_T_64338[4]}},_T_64338}; // @[Modules.scala 32:22:@8.4]
  assign _T_65855 = $signed(buffer_3_92) + $signed(buffer_3_93); // @[Modules.scala 50:57:@13584.4]
  assign _T_65856 = _T_65855[10:0]; // @[Modules.scala 50:57:@13585.4]
  assign buffer_3_438 = $signed(_T_65856); // @[Modules.scala 50:57:@13586.4]
  assign _T_65858 = $signed(buffer_1_94) + $signed(buffer_0_95); // @[Modules.scala 50:57:@13588.4]
  assign _T_65859 = _T_65858[10:0]; // @[Modules.scala 50:57:@13589.4]
  assign buffer_3_439 = $signed(_T_65859); // @[Modules.scala 50:57:@13590.4]
  assign buffer_3_98 = {{6{_T_64357[4]}},_T_64357}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_99 = {{6{_T_64360[4]}},_T_64360}; // @[Modules.scala 32:22:@8.4]
  assign _T_65864 = $signed(buffer_3_98) + $signed(buffer_3_99); // @[Modules.scala 50:57:@13596.4]
  assign _T_65865 = _T_65864[10:0]; // @[Modules.scala 50:57:@13597.4]
  assign buffer_3_441 = $signed(_T_65865); // @[Modules.scala 50:57:@13598.4]
  assign buffer_3_100 = {{6{_T_64363[4]}},_T_64363}; // @[Modules.scala 32:22:@8.4]
  assign _T_65867 = $signed(buffer_3_100) + $signed(buffer_1_101); // @[Modules.scala 50:57:@13600.4]
  assign _T_65868 = _T_65867[10:0]; // @[Modules.scala 50:57:@13601.4]
  assign buffer_3_442 = $signed(_T_65868); // @[Modules.scala 50:57:@13602.4]
  assign buffer_3_103 = {{6{_T_64376[4]}},_T_64376}; // @[Modules.scala 32:22:@8.4]
  assign _T_65870 = $signed(buffer_1_102) + $signed(buffer_3_103); // @[Modules.scala 50:57:@13604.4]
  assign _T_65871 = _T_65870[10:0]; // @[Modules.scala 50:57:@13605.4]
  assign buffer_3_443 = $signed(_T_65871); // @[Modules.scala 50:57:@13606.4]
  assign buffer_3_104 = {{6{_T_64379[4]}},_T_64379}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_105 = {{6{_T_64382[4]}},_T_64382}; // @[Modules.scala 32:22:@8.4]
  assign _T_65873 = $signed(buffer_3_104) + $signed(buffer_3_105); // @[Modules.scala 50:57:@13608.4]
  assign _T_65874 = _T_65873[10:0]; // @[Modules.scala 50:57:@13609.4]
  assign buffer_3_444 = $signed(_T_65874); // @[Modules.scala 50:57:@13610.4]
  assign buffer_3_106 = {{6{_T_64385[4]}},_T_64385}; // @[Modules.scala 32:22:@8.4]
  assign _T_65876 = $signed(buffer_3_106) + $signed(buffer_2_107); // @[Modules.scala 50:57:@13612.4]
  assign _T_65877 = _T_65876[10:0]; // @[Modules.scala 50:57:@13613.4]
  assign buffer_3_445 = $signed(_T_65877); // @[Modules.scala 50:57:@13614.4]
  assign buffer_3_109 = {{6{_T_64398[4]}},_T_64398}; // @[Modules.scala 32:22:@8.4]
  assign _T_65879 = $signed(buffer_1_108) + $signed(buffer_3_109); // @[Modules.scala 50:57:@13616.4]
  assign _T_65880 = _T_65879[10:0]; // @[Modules.scala 50:57:@13617.4]
  assign buffer_3_446 = $signed(_T_65880); // @[Modules.scala 50:57:@13618.4]
  assign buffer_3_113 = {{6{_T_64410[4]}},_T_64410}; // @[Modules.scala 32:22:@8.4]
  assign _T_65885 = $signed(buffer_1_112) + $signed(buffer_3_113); // @[Modules.scala 50:57:@13624.4]
  assign _T_65886 = _T_65885[10:0]; // @[Modules.scala 50:57:@13625.4]
  assign buffer_3_448 = $signed(_T_65886); // @[Modules.scala 50:57:@13626.4]
  assign buffer_3_114 = {{6{_T_64413[4]}},_T_64413}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_115 = {{6{_T_64420[4]}},_T_64420}; // @[Modules.scala 32:22:@8.4]
  assign _T_65888 = $signed(buffer_3_114) + $signed(buffer_3_115); // @[Modules.scala 50:57:@13628.4]
  assign _T_65889 = _T_65888[10:0]; // @[Modules.scala 50:57:@13629.4]
  assign buffer_3_449 = $signed(_T_65889); // @[Modules.scala 50:57:@13630.4]
  assign buffer_3_116 = {{6{_T_64423[4]}},_T_64423}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_117 = {{6{_T_64426[4]}},_T_64426}; // @[Modules.scala 32:22:@8.4]
  assign _T_65891 = $signed(buffer_3_116) + $signed(buffer_3_117); // @[Modules.scala 50:57:@13632.4]
  assign _T_65892 = _T_65891[10:0]; // @[Modules.scala 50:57:@13633.4]
  assign buffer_3_450 = $signed(_T_65892); // @[Modules.scala 50:57:@13634.4]
  assign buffer_3_118 = {{6{_T_64429[4]}},_T_64429}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_119 = {{6{_T_64432[4]}},_T_64432}; // @[Modules.scala 32:22:@8.4]
  assign _T_65894 = $signed(buffer_3_118) + $signed(buffer_3_119); // @[Modules.scala 50:57:@13636.4]
  assign _T_65895 = _T_65894[10:0]; // @[Modules.scala 50:57:@13637.4]
  assign buffer_3_451 = $signed(_T_65895); // @[Modules.scala 50:57:@13638.4]
  assign buffer_3_121 = {{6{_T_64438[4]}},_T_64438}; // @[Modules.scala 32:22:@8.4]
  assign _T_65897 = $signed(buffer_1_120) + $signed(buffer_3_121); // @[Modules.scala 50:57:@13640.4]
  assign _T_65898 = _T_65897[10:0]; // @[Modules.scala 50:57:@13641.4]
  assign buffer_3_452 = $signed(_T_65898); // @[Modules.scala 50:57:@13642.4]
  assign buffer_3_122 = {{6{_T_64441[4]}},_T_64441}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_123 = {{6{_T_64444[4]}},_T_64444}; // @[Modules.scala 32:22:@8.4]
  assign _T_65900 = $signed(buffer_3_122) + $signed(buffer_3_123); // @[Modules.scala 50:57:@13644.4]
  assign _T_65901 = _T_65900[10:0]; // @[Modules.scala 50:57:@13645.4]
  assign buffer_3_453 = $signed(_T_65901); // @[Modules.scala 50:57:@13646.4]
  assign buffer_3_126 = {{6{_T_64453[4]}},_T_64453}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_127 = {{6{_T_64456[4]}},_T_64456}; // @[Modules.scala 32:22:@8.4]
  assign _T_65906 = $signed(buffer_3_126) + $signed(buffer_3_127); // @[Modules.scala 50:57:@13652.4]
  assign _T_65907 = _T_65906[10:0]; // @[Modules.scala 50:57:@13653.4]
  assign buffer_3_455 = $signed(_T_65907); // @[Modules.scala 50:57:@13654.4]
  assign buffer_3_128 = {{6{_T_64459[4]}},_T_64459}; // @[Modules.scala 32:22:@8.4]
  assign _T_65909 = $signed(buffer_3_128) + $signed(buffer_0_129); // @[Modules.scala 50:57:@13656.4]
  assign _T_65910 = _T_65909[10:0]; // @[Modules.scala 50:57:@13657.4]
  assign buffer_3_456 = $signed(_T_65910); // @[Modules.scala 50:57:@13658.4]
  assign buffer_3_132 = {{6{_T_64483[4]}},_T_64483}; // @[Modules.scala 32:22:@8.4]
  assign _T_65915 = $signed(buffer_3_132) + $signed(buffer_1_133); // @[Modules.scala 50:57:@13664.4]
  assign _T_65916 = _T_65915[10:0]; // @[Modules.scala 50:57:@13665.4]
  assign buffer_3_458 = $signed(_T_65916); // @[Modules.scala 50:57:@13666.4]
  assign buffer_3_134 = {{6{_T_64489[4]}},_T_64489}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_135 = {{6{_T_64492[4]}},_T_64492}; // @[Modules.scala 32:22:@8.4]
  assign _T_65918 = $signed(buffer_3_134) + $signed(buffer_3_135); // @[Modules.scala 50:57:@13668.4]
  assign _T_65919 = _T_65918[10:0]; // @[Modules.scala 50:57:@13669.4]
  assign buffer_3_459 = $signed(_T_65919); // @[Modules.scala 50:57:@13670.4]
  assign buffer_3_136 = {{6{_T_64495[4]}},_T_64495}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_137 = {{6{_T_64498[4]}},_T_64498}; // @[Modules.scala 32:22:@8.4]
  assign _T_65921 = $signed(buffer_3_136) + $signed(buffer_3_137); // @[Modules.scala 50:57:@13672.4]
  assign _T_65922 = _T_65921[10:0]; // @[Modules.scala 50:57:@13673.4]
  assign buffer_3_460 = $signed(_T_65922); // @[Modules.scala 50:57:@13674.4]
  assign buffer_3_140 = {{6{_T_64507[4]}},_T_64507}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_141 = {{6{_T_64510[4]}},_T_64510}; // @[Modules.scala 32:22:@8.4]
  assign _T_65927 = $signed(buffer_3_140) + $signed(buffer_3_141); // @[Modules.scala 50:57:@13680.4]
  assign _T_65928 = _T_65927[10:0]; // @[Modules.scala 50:57:@13681.4]
  assign buffer_3_462 = $signed(_T_65928); // @[Modules.scala 50:57:@13682.4]
  assign buffer_3_142 = {{6{_T_64513[4]}},_T_64513}; // @[Modules.scala 32:22:@8.4]
  assign _T_65930 = $signed(buffer_3_142) + $signed(buffer_0_143); // @[Modules.scala 50:57:@13684.4]
  assign _T_65931 = _T_65930[10:0]; // @[Modules.scala 50:57:@13685.4]
  assign buffer_3_463 = $signed(_T_65931); // @[Modules.scala 50:57:@13686.4]
  assign buffer_3_144 = {{6{_T_64527[4]}},_T_64527}; // @[Modules.scala 32:22:@8.4]
  assign _T_65933 = $signed(buffer_3_144) + $signed(buffer_0_145); // @[Modules.scala 50:57:@13688.4]
  assign _T_65934 = _T_65933[10:0]; // @[Modules.scala 50:57:@13689.4]
  assign buffer_3_464 = $signed(_T_65934); // @[Modules.scala 50:57:@13690.4]
  assign buffer_3_147 = {{6{_T_64548[4]}},_T_64548}; // @[Modules.scala 32:22:@8.4]
  assign _T_65936 = $signed(buffer_0_146) + $signed(buffer_3_147); // @[Modules.scala 50:57:@13692.4]
  assign _T_65937 = _T_65936[10:0]; // @[Modules.scala 50:57:@13693.4]
  assign buffer_3_465 = $signed(_T_65937); // @[Modules.scala 50:57:@13694.4]
  assign buffer_3_148 = {{6{_T_64551[4]}},_T_64551}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_149 = {{6{_T_64554[4]}},_T_64554}; // @[Modules.scala 32:22:@8.4]
  assign _T_65939 = $signed(buffer_3_148) + $signed(buffer_3_149); // @[Modules.scala 50:57:@13696.4]
  assign _T_65940 = _T_65939[10:0]; // @[Modules.scala 50:57:@13697.4]
  assign buffer_3_466 = $signed(_T_65940); // @[Modules.scala 50:57:@13698.4]
  assign buffer_3_150 = {{6{_T_64557[4]}},_T_64557}; // @[Modules.scala 32:22:@8.4]
  assign _T_65942 = $signed(buffer_3_150) + $signed(buffer_0_151); // @[Modules.scala 50:57:@13700.4]
  assign _T_65943 = _T_65942[10:0]; // @[Modules.scala 50:57:@13701.4]
  assign buffer_3_467 = $signed(_T_65943); // @[Modules.scala 50:57:@13702.4]
  assign buffer_3_154 = {{6{_T_64577[4]}},_T_64577}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_155 = {{6{_T_64580[4]}},_T_64580}; // @[Modules.scala 32:22:@8.4]
  assign _T_65948 = $signed(buffer_3_154) + $signed(buffer_3_155); // @[Modules.scala 50:57:@13708.4]
  assign _T_65949 = _T_65948[10:0]; // @[Modules.scala 50:57:@13709.4]
  assign buffer_3_469 = $signed(_T_65949); // @[Modules.scala 50:57:@13710.4]
  assign buffer_3_157 = {{6{_T_64594[4]}},_T_64594}; // @[Modules.scala 32:22:@8.4]
  assign _T_65951 = $signed(buffer_0_156) + $signed(buffer_3_157); // @[Modules.scala 50:57:@13712.4]
  assign _T_65952 = _T_65951[10:0]; // @[Modules.scala 50:57:@13713.4]
  assign buffer_3_470 = $signed(_T_65952); // @[Modules.scala 50:57:@13714.4]
  assign buffer_3_159 = {{6{_T_64608[4]}},_T_64608}; // @[Modules.scala 32:22:@8.4]
  assign _T_65954 = $signed(buffer_1_158) + $signed(buffer_3_159); // @[Modules.scala 50:57:@13716.4]
  assign _T_65955 = _T_65954[10:0]; // @[Modules.scala 50:57:@13717.4]
  assign buffer_3_471 = $signed(_T_65955); // @[Modules.scala 50:57:@13718.4]
  assign buffer_3_167 = {{6{_T_64660[4]}},_T_64660}; // @[Modules.scala 32:22:@8.4]
  assign _T_65966 = $signed(buffer_0_166) + $signed(buffer_3_167); // @[Modules.scala 50:57:@13732.4]
  assign _T_65967 = _T_65966[10:0]; // @[Modules.scala 50:57:@13733.4]
  assign buffer_3_475 = $signed(_T_65967); // @[Modules.scala 50:57:@13734.4]
  assign buffer_3_168 = {{6{_T_64667[4]}},_T_64667}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_169 = {{6{_T_64670[4]}},_T_64670}; // @[Modules.scala 32:22:@8.4]
  assign _T_65969 = $signed(buffer_3_168) + $signed(buffer_3_169); // @[Modules.scala 50:57:@13736.4]
  assign _T_65970 = _T_65969[10:0]; // @[Modules.scala 50:57:@13737.4]
  assign buffer_3_476 = $signed(_T_65970); // @[Modules.scala 50:57:@13738.4]
  assign buffer_3_170 = {{6{_T_64677[4]}},_T_64677}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_171 = {{6{_T_64684[4]}},_T_64684}; // @[Modules.scala 32:22:@8.4]
  assign _T_65972 = $signed(buffer_3_170) + $signed(buffer_3_171); // @[Modules.scala 50:57:@13740.4]
  assign _T_65973 = _T_65972[10:0]; // @[Modules.scala 50:57:@13741.4]
  assign buffer_3_477 = $signed(_T_65973); // @[Modules.scala 50:57:@13742.4]
  assign buffer_3_172 = {{6{_T_64691[4]}},_T_64691}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_173 = {{6{_T_64698[4]}},_T_64698}; // @[Modules.scala 32:22:@8.4]
  assign _T_65975 = $signed(buffer_3_172) + $signed(buffer_3_173); // @[Modules.scala 50:57:@13744.4]
  assign _T_65976 = _T_65975[10:0]; // @[Modules.scala 50:57:@13745.4]
  assign buffer_3_478 = $signed(_T_65976); // @[Modules.scala 50:57:@13746.4]
  assign buffer_3_174 = {{6{_T_64705[4]}},_T_64705}; // @[Modules.scala 32:22:@8.4]
  assign _T_65978 = $signed(buffer_3_174) + $signed(buffer_1_175); // @[Modules.scala 50:57:@13748.4]
  assign _T_65979 = _T_65978[10:0]; // @[Modules.scala 50:57:@13749.4]
  assign buffer_3_479 = $signed(_T_65979); // @[Modules.scala 50:57:@13750.4]
  assign _T_65987 = $signed(buffer_0_180) + $signed(buffer_1_181); // @[Modules.scala 50:57:@13760.4]
  assign _T_65988 = _T_65987[10:0]; // @[Modules.scala 50:57:@13761.4]
  assign buffer_3_482 = $signed(_T_65988); // @[Modules.scala 50:57:@13762.4]
  assign buffer_3_182 = {{6{_T_64757[4]}},_T_64757}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_183 = {{6{_T_64760[4]}},_T_64760}; // @[Modules.scala 32:22:@8.4]
  assign _T_65990 = $signed(buffer_3_182) + $signed(buffer_3_183); // @[Modules.scala 50:57:@13764.4]
  assign _T_65991 = _T_65990[10:0]; // @[Modules.scala 50:57:@13765.4]
  assign buffer_3_483 = $signed(_T_65991); // @[Modules.scala 50:57:@13766.4]
  assign buffer_3_184 = {{6{_T_64767[4]}},_T_64767}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_185 = {{6{_T_64774[4]}},_T_64774}; // @[Modules.scala 32:22:@8.4]
  assign _T_65993 = $signed(buffer_3_184) + $signed(buffer_3_185); // @[Modules.scala 50:57:@13768.4]
  assign _T_65994 = _T_65993[10:0]; // @[Modules.scala 50:57:@13769.4]
  assign buffer_3_484 = $signed(_T_65994); // @[Modules.scala 50:57:@13770.4]
  assign buffer_3_186 = {{6{_T_64781[4]}},_T_64781}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_187 = {{6{_T_64788[4]}},_T_64788}; // @[Modules.scala 32:22:@8.4]
  assign _T_65996 = $signed(buffer_3_186) + $signed(buffer_3_187); // @[Modules.scala 50:57:@13772.4]
  assign _T_65997 = _T_65996[10:0]; // @[Modules.scala 50:57:@13773.4]
  assign buffer_3_485 = $signed(_T_65997); // @[Modules.scala 50:57:@13774.4]
  assign buffer_3_188 = {{6{_T_64795[4]}},_T_64795}; // @[Modules.scala 32:22:@8.4]
  assign _T_65999 = $signed(buffer_3_188) + $signed(buffer_1_189); // @[Modules.scala 50:57:@13776.4]
  assign _T_66000 = _T_65999[10:0]; // @[Modules.scala 50:57:@13777.4]
  assign buffer_3_486 = $signed(_T_66000); // @[Modules.scala 50:57:@13778.4]
  assign buffer_3_190 = {{6{_T_64809[4]}},_T_64809}; // @[Modules.scala 32:22:@8.4]
  assign _T_66002 = $signed(buffer_3_190) + $signed(buffer_1_191); // @[Modules.scala 50:57:@13780.4]
  assign _T_66003 = _T_66002[10:0]; // @[Modules.scala 50:57:@13781.4]
  assign buffer_3_487 = $signed(_T_66003); // @[Modules.scala 50:57:@13782.4]
  assign buffer_3_192 = {{6{_T_64823[4]}},_T_64823}; // @[Modules.scala 32:22:@8.4]
  assign _T_66005 = $signed(buffer_3_192) + $signed(buffer_2_193); // @[Modules.scala 50:57:@13784.4]
  assign _T_66006 = _T_66005[10:0]; // @[Modules.scala 50:57:@13785.4]
  assign buffer_3_488 = $signed(_T_66006); // @[Modules.scala 50:57:@13786.4]
  assign buffer_3_195 = {{6{_T_64840[4]}},_T_64840}; // @[Modules.scala 32:22:@8.4]
  assign _T_66008 = $signed(buffer_2_194) + $signed(buffer_3_195); // @[Modules.scala 50:57:@13788.4]
  assign _T_66009 = _T_66008[10:0]; // @[Modules.scala 50:57:@13789.4]
  assign buffer_3_489 = $signed(_T_66009); // @[Modules.scala 50:57:@13790.4]
  assign buffer_3_197 = {{6{_T_64846[4]}},_T_64846}; // @[Modules.scala 32:22:@8.4]
  assign _T_66011 = $signed(buffer_1_196) + $signed(buffer_3_197); // @[Modules.scala 50:57:@13792.4]
  assign _T_66012 = _T_66011[10:0]; // @[Modules.scala 50:57:@13793.4]
  assign buffer_3_490 = $signed(_T_66012); // @[Modules.scala 50:57:@13794.4]
  assign buffer_3_198 = {{6{_T_64853[4]}},_T_64853}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_199 = {{6{_T_64860[4]}},_T_64860}; // @[Modules.scala 32:22:@8.4]
  assign _T_66014 = $signed(buffer_3_198) + $signed(buffer_3_199); // @[Modules.scala 50:57:@13796.4]
  assign _T_66015 = _T_66014[10:0]; // @[Modules.scala 50:57:@13797.4]
  assign buffer_3_491 = $signed(_T_66015); // @[Modules.scala 50:57:@13798.4]
  assign buffer_3_200 = {{6{_T_64867[4]}},_T_64867}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_201 = {{6{_T_64870[4]}},_T_64870}; // @[Modules.scala 32:22:@8.4]
  assign _T_66017 = $signed(buffer_3_200) + $signed(buffer_3_201); // @[Modules.scala 50:57:@13800.4]
  assign _T_66018 = _T_66017[10:0]; // @[Modules.scala 50:57:@13801.4]
  assign buffer_3_492 = $signed(_T_66018); // @[Modules.scala 50:57:@13802.4]
  assign buffer_3_202 = {{6{_T_64877[4]}},_T_64877}; // @[Modules.scala 32:22:@8.4]
  assign _T_66020 = $signed(buffer_3_202) + $signed(buffer_1_203); // @[Modules.scala 50:57:@13804.4]
  assign _T_66021 = _T_66020[10:0]; // @[Modules.scala 50:57:@13805.4]
  assign buffer_3_493 = $signed(_T_66021); // @[Modules.scala 50:57:@13806.4]
  assign buffer_3_204 = {{6{_T_64891[4]}},_T_64891}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_205 = {{6{_T_64894[4]}},_T_64894}; // @[Modules.scala 32:22:@8.4]
  assign _T_66023 = $signed(buffer_3_204) + $signed(buffer_3_205); // @[Modules.scala 50:57:@13808.4]
  assign _T_66024 = _T_66023[10:0]; // @[Modules.scala 50:57:@13809.4]
  assign buffer_3_494 = $signed(_T_66024); // @[Modules.scala 50:57:@13810.4]
  assign buffer_3_206 = {{6{_T_64901[4]}},_T_64901}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_207 = {{6{_T_64908[4]}},_T_64908}; // @[Modules.scala 32:22:@8.4]
  assign _T_66026 = $signed(buffer_3_206) + $signed(buffer_3_207); // @[Modules.scala 50:57:@13812.4]
  assign _T_66027 = _T_66026[10:0]; // @[Modules.scala 50:57:@13813.4]
  assign buffer_3_495 = $signed(_T_66027); // @[Modules.scala 50:57:@13814.4]
  assign buffer_3_208 = {{6{_T_64915[4]}},_T_64915}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_209 = {{6{_T_64918[4]}},_T_64918}; // @[Modules.scala 32:22:@8.4]
  assign _T_66029 = $signed(buffer_3_208) + $signed(buffer_3_209); // @[Modules.scala 50:57:@13816.4]
  assign _T_66030 = _T_66029[10:0]; // @[Modules.scala 50:57:@13817.4]
  assign buffer_3_496 = $signed(_T_66030); // @[Modules.scala 50:57:@13818.4]
  assign buffer_3_210 = {{6{_T_64921[4]}},_T_64921}; // @[Modules.scala 32:22:@8.4]
  assign _T_66032 = $signed(buffer_3_210) + $signed(buffer_2_211); // @[Modules.scala 50:57:@13820.4]
  assign _T_66033 = _T_66032[10:0]; // @[Modules.scala 50:57:@13821.4]
  assign buffer_3_497 = $signed(_T_66033); // @[Modules.scala 50:57:@13822.4]
  assign buffer_3_212 = {{6{_T_64927[4]}},_T_64927}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_213 = {{6{_T_64934[4]}},_T_64934}; // @[Modules.scala 32:22:@8.4]
  assign _T_66035 = $signed(buffer_3_212) + $signed(buffer_3_213); // @[Modules.scala 50:57:@13824.4]
  assign _T_66036 = _T_66035[10:0]; // @[Modules.scala 50:57:@13825.4]
  assign buffer_3_498 = $signed(_T_66036); // @[Modules.scala 50:57:@13826.4]
  assign buffer_3_220 = {{6{_T_64979[4]}},_T_64979}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_221 = {{6{_T_64986[4]}},_T_64986}; // @[Modules.scala 32:22:@8.4]
  assign _T_66047 = $signed(buffer_3_220) + $signed(buffer_3_221); // @[Modules.scala 50:57:@13840.4]
  assign _T_66048 = _T_66047[10:0]; // @[Modules.scala 50:57:@13841.4]
  assign buffer_3_502 = $signed(_T_66048); // @[Modules.scala 50:57:@13842.4]
  assign buffer_3_222 = {{6{_T_64989[4]}},_T_64989}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_223 = {{6{_T_64992[4]}},_T_64992}; // @[Modules.scala 32:22:@8.4]
  assign _T_66050 = $signed(buffer_3_222) + $signed(buffer_3_223); // @[Modules.scala 50:57:@13844.4]
  assign _T_66051 = _T_66050[10:0]; // @[Modules.scala 50:57:@13845.4]
  assign buffer_3_503 = $signed(_T_66051); // @[Modules.scala 50:57:@13846.4]
  assign buffer_3_224 = {{6{_T_64995[4]}},_T_64995}; // @[Modules.scala 32:22:@8.4]
  assign _T_66053 = $signed(buffer_3_224) + $signed(buffer_1_225); // @[Modules.scala 50:57:@13848.4]
  assign _T_66054 = _T_66053[10:0]; // @[Modules.scala 50:57:@13849.4]
  assign buffer_3_504 = $signed(_T_66054); // @[Modules.scala 50:57:@13850.4]
  assign buffer_3_226 = {{6{_T_65001[4]}},_T_65001}; // @[Modules.scala 32:22:@8.4]
  assign _T_66056 = $signed(buffer_3_226) + $signed(buffer_0_227); // @[Modules.scala 50:57:@13852.4]
  assign _T_66057 = _T_66056[10:0]; // @[Modules.scala 50:57:@13853.4]
  assign buffer_3_505 = $signed(_T_66057); // @[Modules.scala 50:57:@13854.4]
  assign buffer_3_228 = {{6{_T_65011[4]}},_T_65011}; // @[Modules.scala 32:22:@8.4]
  assign _T_66059 = $signed(buffer_3_228) + $signed(buffer_2_229); // @[Modules.scala 50:57:@13856.4]
  assign _T_66060 = _T_66059[10:0]; // @[Modules.scala 50:57:@13857.4]
  assign buffer_3_506 = $signed(_T_66060); // @[Modules.scala 50:57:@13858.4]
  assign _T_66065 = $signed(buffer_1_232) + $signed(buffer_0_233); // @[Modules.scala 50:57:@13864.4]
  assign _T_66066 = _T_66065[10:0]; // @[Modules.scala 50:57:@13865.4]
  assign buffer_3_508 = $signed(_T_66066); // @[Modules.scala 50:57:@13866.4]
  assign buffer_3_236 = {{6{_T_65051[4]}},_T_65051}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_237 = {{6{_T_65054[4]}},_T_65054}; // @[Modules.scala 32:22:@8.4]
  assign _T_66071 = $signed(buffer_3_236) + $signed(buffer_3_237); // @[Modules.scala 50:57:@13872.4]
  assign _T_66072 = _T_66071[10:0]; // @[Modules.scala 50:57:@13873.4]
  assign buffer_3_510 = $signed(_T_66072); // @[Modules.scala 50:57:@13874.4]
  assign _T_66074 = $signed(buffer_0_238) + $signed(buffer_1_239); // @[Modules.scala 50:57:@13876.4]
  assign _T_66075 = _T_66074[10:0]; // @[Modules.scala 50:57:@13877.4]
  assign buffer_3_511 = $signed(_T_66075); // @[Modules.scala 50:57:@13878.4]
  assign buffer_3_240 = {{6{_T_65067[4]}},_T_65067}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_241 = {{6{_T_65070[4]}},_T_65070}; // @[Modules.scala 32:22:@8.4]
  assign _T_66077 = $signed(buffer_3_240) + $signed(buffer_3_241); // @[Modules.scala 50:57:@13880.4]
  assign _T_66078 = _T_66077[10:0]; // @[Modules.scala 50:57:@13881.4]
  assign buffer_3_512 = $signed(_T_66078); // @[Modules.scala 50:57:@13882.4]
  assign buffer_3_246 = {{6{_T_65105[4]}},_T_65105}; // @[Modules.scala 32:22:@8.4]
  assign _T_66086 = $signed(buffer_3_246) + $signed(buffer_1_247); // @[Modules.scala 50:57:@13892.4]
  assign _T_66087 = _T_66086[10:0]; // @[Modules.scala 50:57:@13893.4]
  assign buffer_3_515 = $signed(_T_66087); // @[Modules.scala 50:57:@13894.4]
  assign buffer_3_250 = {{6{_T_65117[4]}},_T_65117}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_251 = {{6{_T_65120[4]}},_T_65120}; // @[Modules.scala 32:22:@8.4]
  assign _T_66092 = $signed(buffer_3_250) + $signed(buffer_3_251); // @[Modules.scala 50:57:@13900.4]
  assign _T_66093 = _T_66092[10:0]; // @[Modules.scala 50:57:@13901.4]
  assign buffer_3_517 = $signed(_T_66093); // @[Modules.scala 50:57:@13902.4]
  assign buffer_3_252 = {{6{_T_65123[4]}},_T_65123}; // @[Modules.scala 32:22:@8.4]
  assign _T_66095 = $signed(buffer_3_252) + $signed(buffer_1_253); // @[Modules.scala 50:57:@13904.4]
  assign _T_66096 = _T_66095[10:0]; // @[Modules.scala 50:57:@13905.4]
  assign buffer_3_518 = $signed(_T_66096); // @[Modules.scala 50:57:@13906.4]
  assign buffer_3_254 = {{6{_T_65129[4]}},_T_65129}; // @[Modules.scala 32:22:@8.4]
  assign _T_66098 = $signed(buffer_3_254) + $signed(buffer_1_255); // @[Modules.scala 50:57:@13908.4]
  assign _T_66099 = _T_66098[10:0]; // @[Modules.scala 50:57:@13909.4]
  assign buffer_3_519 = $signed(_T_66099); // @[Modules.scala 50:57:@13910.4]
  assign buffer_3_257 = {{6{_T_65146[4]}},_T_65146}; // @[Modules.scala 32:22:@8.4]
  assign _T_66101 = $signed(buffer_1_256) + $signed(buffer_3_257); // @[Modules.scala 50:57:@13912.4]
  assign _T_66102 = _T_66101[10:0]; // @[Modules.scala 50:57:@13913.4]
  assign buffer_3_520 = $signed(_T_66102); // @[Modules.scala 50:57:@13914.4]
  assign buffer_3_265 = {{6{_T_65182[4]}},_T_65182}; // @[Modules.scala 32:22:@8.4]
  assign _T_66113 = $signed(buffer_0_264) + $signed(buffer_3_265); // @[Modules.scala 50:57:@13928.4]
  assign _T_66114 = _T_66113[10:0]; // @[Modules.scala 50:57:@13929.4]
  assign buffer_3_524 = $signed(_T_66114); // @[Modules.scala 50:57:@13930.4]
  assign buffer_3_270 = {{6{_T_65197[4]}},_T_65197}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_271 = {{6{_T_65204[4]}},_T_65204}; // @[Modules.scala 32:22:@8.4]
  assign _T_66122 = $signed(buffer_3_270) + $signed(buffer_3_271); // @[Modules.scala 50:57:@13940.4]
  assign _T_66123 = _T_66122[10:0]; // @[Modules.scala 50:57:@13941.4]
  assign buffer_3_527 = $signed(_T_66123); // @[Modules.scala 50:57:@13942.4]
  assign buffer_3_273 = {{6{_T_65214[4]}},_T_65214}; // @[Modules.scala 32:22:@8.4]
  assign _T_66125 = $signed(buffer_0_272) + $signed(buffer_3_273); // @[Modules.scala 50:57:@13944.4]
  assign _T_66126 = _T_66125[10:0]; // @[Modules.scala 50:57:@13945.4]
  assign buffer_3_528 = $signed(_T_66126); // @[Modules.scala 50:57:@13946.4]
  assign buffer_3_275 = {{6{_T_65228[4]}},_T_65228}; // @[Modules.scala 32:22:@8.4]
  assign _T_66128 = $signed(buffer_0_274) + $signed(buffer_3_275); // @[Modules.scala 50:57:@13948.4]
  assign _T_66129 = _T_66128[10:0]; // @[Modules.scala 50:57:@13949.4]
  assign buffer_3_529 = $signed(_T_66129); // @[Modules.scala 50:57:@13950.4]
  assign buffer_3_277 = {{6{_T_65234[4]}},_T_65234}; // @[Modules.scala 32:22:@8.4]
  assign _T_66131 = $signed(buffer_2_276) + $signed(buffer_3_277); // @[Modules.scala 50:57:@13952.4]
  assign _T_66132 = _T_66131[10:0]; // @[Modules.scala 50:57:@13953.4]
  assign buffer_3_530 = $signed(_T_66132); // @[Modules.scala 50:57:@13954.4]
  assign buffer_3_278 = {{6{_T_65237[4]}},_T_65237}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_279 = {{6{_T_65240[4]}},_T_65240}; // @[Modules.scala 32:22:@8.4]
  assign _T_66134 = $signed(buffer_3_278) + $signed(buffer_3_279); // @[Modules.scala 50:57:@13956.4]
  assign _T_66135 = _T_66134[10:0]; // @[Modules.scala 50:57:@13957.4]
  assign buffer_3_531 = $signed(_T_66135); // @[Modules.scala 50:57:@13958.4]
  assign _T_66137 = $signed(buffer_2_280) + $signed(buffer_1_281); // @[Modules.scala 50:57:@13960.4]
  assign _T_66138 = _T_66137[10:0]; // @[Modules.scala 50:57:@13961.4]
  assign buffer_3_532 = $signed(_T_66138); // @[Modules.scala 50:57:@13962.4]
  assign buffer_3_283 = {{6{_T_65252[4]}},_T_65252}; // @[Modules.scala 32:22:@8.4]
  assign _T_66140 = $signed(buffer_1_282) + $signed(buffer_3_283); // @[Modules.scala 50:57:@13964.4]
  assign _T_66141 = _T_66140[10:0]; // @[Modules.scala 50:57:@13965.4]
  assign buffer_3_533 = $signed(_T_66141); // @[Modules.scala 50:57:@13966.4]
  assign buffer_3_286 = {{6{_T_65261[4]}},_T_65261}; // @[Modules.scala 32:22:@8.4]
  assign _T_66146 = $signed(buffer_3_286) + $signed(buffer_0_287); // @[Modules.scala 50:57:@13972.4]
  assign _T_66147 = _T_66146[10:0]; // @[Modules.scala 50:57:@13973.4]
  assign buffer_3_535 = $signed(_T_66147); // @[Modules.scala 50:57:@13974.4]
  assign _T_66149 = $signed(buffer_1_288) + $signed(buffer_0_289); // @[Modules.scala 50:57:@13976.4]
  assign _T_66150 = _T_66149[10:0]; // @[Modules.scala 50:57:@13977.4]
  assign buffer_3_536 = $signed(_T_66150); // @[Modules.scala 50:57:@13978.4]
  assign buffer_3_291 = {{6{_T_65280[4]}},_T_65280}; // @[Modules.scala 32:22:@8.4]
  assign _T_66152 = $signed(buffer_0_290) + $signed(buffer_3_291); // @[Modules.scala 50:57:@13980.4]
  assign _T_66153 = _T_66152[10:0]; // @[Modules.scala 50:57:@13981.4]
  assign buffer_3_537 = $signed(_T_66153); // @[Modules.scala 50:57:@13982.4]
  assign buffer_3_293 = {{6{_T_65286[4]}},_T_65286}; // @[Modules.scala 32:22:@8.4]
  assign _T_66155 = $signed(buffer_0_292) + $signed(buffer_3_293); // @[Modules.scala 50:57:@13984.4]
  assign _T_66156 = _T_66155[10:0]; // @[Modules.scala 50:57:@13985.4]
  assign buffer_3_538 = $signed(_T_66156); // @[Modules.scala 50:57:@13986.4]
  assign buffer_3_297 = {{6{_T_65302[4]}},_T_65302}; // @[Modules.scala 32:22:@8.4]
  assign _T_66161 = $signed(buffer_1_296) + $signed(buffer_3_297); // @[Modules.scala 50:57:@13992.4]
  assign _T_66162 = _T_66161[10:0]; // @[Modules.scala 50:57:@13993.4]
  assign buffer_3_540 = $signed(_T_66162); // @[Modules.scala 50:57:@13994.4]
  assign _T_66164 = $signed(buffer_1_298) + $signed(buffer_0_299); // @[Modules.scala 50:57:@13996.4]
  assign _T_66165 = _T_66164[10:0]; // @[Modules.scala 50:57:@13997.4]
  assign buffer_3_541 = $signed(_T_66165); // @[Modules.scala 50:57:@13998.4]
  assign buffer_3_301 = {{6{_T_65326[4]}},_T_65326}; // @[Modules.scala 32:22:@8.4]
  assign _T_66167 = $signed(buffer_2_300) + $signed(buffer_3_301); // @[Modules.scala 50:57:@14000.4]
  assign _T_66168 = _T_66167[10:0]; // @[Modules.scala 50:57:@14001.4]
  assign buffer_3_542 = $signed(_T_66168); // @[Modules.scala 50:57:@14002.4]
  assign _T_66170 = $signed(buffer_2_302) + $signed(buffer_0_303); // @[Modules.scala 50:57:@14004.4]
  assign _T_66171 = _T_66170[10:0]; // @[Modules.scala 50:57:@14005.4]
  assign buffer_3_543 = $signed(_T_66171); // @[Modules.scala 50:57:@14006.4]
  assign buffer_3_304 = {{6{_T_65343[4]}},_T_65343}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_305 = {{6{_T_65346[4]}},_T_65346}; // @[Modules.scala 32:22:@8.4]
  assign _T_66173 = $signed(buffer_3_304) + $signed(buffer_3_305); // @[Modules.scala 50:57:@14008.4]
  assign _T_66174 = _T_66173[10:0]; // @[Modules.scala 50:57:@14009.4]
  assign buffer_3_544 = $signed(_T_66174); // @[Modules.scala 50:57:@14010.4]
  assign buffer_3_307 = {{6{_T_65352[4]}},_T_65352}; // @[Modules.scala 32:22:@8.4]
  assign _T_66176 = $signed(buffer_0_306) + $signed(buffer_3_307); // @[Modules.scala 50:57:@14012.4]
  assign _T_66177 = _T_66176[10:0]; // @[Modules.scala 50:57:@14013.4]
  assign buffer_3_545 = $signed(_T_66177); // @[Modules.scala 50:57:@14014.4]
  assign buffer_3_310 = {{6{_T_65365[4]}},_T_65365}; // @[Modules.scala 32:22:@8.4]
  assign _T_66182 = $signed(buffer_3_310) + $signed(buffer_0_311); // @[Modules.scala 50:57:@14020.4]
  assign _T_66183 = _T_66182[10:0]; // @[Modules.scala 50:57:@14021.4]
  assign buffer_3_547 = $signed(_T_66183); // @[Modules.scala 50:57:@14022.4]
  assign buffer_3_313 = {{6{_T_65382[4]}},_T_65382}; // @[Modules.scala 32:22:@8.4]
  assign _T_66185 = $signed(buffer_1_312) + $signed(buffer_3_313); // @[Modules.scala 50:57:@14024.4]
  assign _T_66186 = _T_66185[10:0]; // @[Modules.scala 50:57:@14025.4]
  assign buffer_3_548 = $signed(_T_66186); // @[Modules.scala 50:57:@14026.4]
  assign buffer_3_315 = {{6{_T_65388[4]}},_T_65388}; // @[Modules.scala 32:22:@8.4]
  assign _T_66188 = $signed(buffer_1_314) + $signed(buffer_3_315); // @[Modules.scala 50:57:@14028.4]
  assign _T_66189 = _T_66188[10:0]; // @[Modules.scala 50:57:@14029.4]
  assign buffer_3_549 = $signed(_T_66189); // @[Modules.scala 50:57:@14030.4]
  assign buffer_3_316 = {{6{_T_65391[4]}},_T_65391}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_317 = {{6{_T_65398[4]}},_T_65398}; // @[Modules.scala 32:22:@8.4]
  assign _T_66191 = $signed(buffer_3_316) + $signed(buffer_3_317); // @[Modules.scala 50:57:@14032.4]
  assign _T_66192 = _T_66191[10:0]; // @[Modules.scala 50:57:@14033.4]
  assign buffer_3_550 = $signed(_T_66192); // @[Modules.scala 50:57:@14034.4]
  assign buffer_3_319 = {{6{_T_65404[4]}},_T_65404}; // @[Modules.scala 32:22:@8.4]
  assign _T_66194 = $signed(buffer_1_318) + $signed(buffer_3_319); // @[Modules.scala 50:57:@14036.4]
  assign _T_66195 = _T_66194[10:0]; // @[Modules.scala 50:57:@14037.4]
  assign buffer_3_551 = $signed(_T_66195); // @[Modules.scala 50:57:@14038.4]
  assign buffer_3_321 = {{6{_T_65410[4]}},_T_65410}; // @[Modules.scala 32:22:@8.4]
  assign _T_66197 = $signed(buffer_0_320) + $signed(buffer_3_321); // @[Modules.scala 50:57:@14040.4]
  assign _T_66198 = _T_66197[10:0]; // @[Modules.scala 50:57:@14041.4]
  assign buffer_3_552 = $signed(_T_66198); // @[Modules.scala 50:57:@14042.4]
  assign _T_66200 = $signed(buffer_2_322) + $signed(buffer_0_323); // @[Modules.scala 50:57:@14044.4]
  assign _T_66201 = _T_66200[10:0]; // @[Modules.scala 50:57:@14045.4]
  assign buffer_3_553 = $signed(_T_66201); // @[Modules.scala 50:57:@14046.4]
  assign buffer_3_325 = {{6{_T_65426[4]}},_T_65426}; // @[Modules.scala 32:22:@8.4]
  assign _T_66203 = $signed(buffer_1_324) + $signed(buffer_3_325); // @[Modules.scala 50:57:@14048.4]
  assign _T_66204 = _T_66203[10:0]; // @[Modules.scala 50:57:@14049.4]
  assign buffer_3_554 = $signed(_T_66204); // @[Modules.scala 50:57:@14050.4]
  assign buffer_3_326 = {{6{_T_65433[4]}},_T_65433}; // @[Modules.scala 32:22:@8.4]
  assign _T_66206 = $signed(buffer_3_326) + $signed(buffer_1_327); // @[Modules.scala 50:57:@14052.4]
  assign _T_66207 = _T_66206[10:0]; // @[Modules.scala 50:57:@14053.4]
  assign buffer_3_555 = $signed(_T_66207); // @[Modules.scala 50:57:@14054.4]
  assign _T_66209 = $signed(buffer_2_328) + $signed(buffer_0_329); // @[Modules.scala 50:57:@14056.4]
  assign _T_66210 = _T_66209[10:0]; // @[Modules.scala 50:57:@14057.4]
  assign buffer_3_556 = $signed(_T_66210); // @[Modules.scala 50:57:@14058.4]
  assign buffer_3_331 = {{6{_T_65460[4]}},_T_65460}; // @[Modules.scala 32:22:@8.4]
  assign _T_66212 = $signed(buffer_0_330) + $signed(buffer_3_331); // @[Modules.scala 50:57:@14060.4]
  assign _T_66213 = _T_66212[10:0]; // @[Modules.scala 50:57:@14061.4]
  assign buffer_3_557 = $signed(_T_66213); // @[Modules.scala 50:57:@14062.4]
  assign buffer_3_333 = {{6{_T_65470[4]}},_T_65470}; // @[Modules.scala 32:22:@8.4]
  assign _T_66215 = $signed(buffer_1_332) + $signed(buffer_3_333); // @[Modules.scala 50:57:@14064.4]
  assign _T_66216 = _T_66215[10:0]; // @[Modules.scala 50:57:@14065.4]
  assign buffer_3_558 = $signed(_T_66216); // @[Modules.scala 50:57:@14066.4]
  assign buffer_3_335 = {{6{_T_65476[4]}},_T_65476}; // @[Modules.scala 32:22:@8.4]
  assign _T_66218 = $signed(buffer_0_334) + $signed(buffer_3_335); // @[Modules.scala 50:57:@14068.4]
  assign _T_66219 = _T_66218[10:0]; // @[Modules.scala 50:57:@14069.4]
  assign buffer_3_559 = $signed(_T_66219); // @[Modules.scala 50:57:@14070.4]
  assign buffer_3_336 = {{6{_T_65479[4]}},_T_65479}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_337 = {{6{_T_65486[4]}},_T_65486}; // @[Modules.scala 32:22:@8.4]
  assign _T_66221 = $signed(buffer_3_336) + $signed(buffer_3_337); // @[Modules.scala 50:57:@14072.4]
  assign _T_66222 = _T_66221[10:0]; // @[Modules.scala 50:57:@14073.4]
  assign buffer_3_560 = $signed(_T_66222); // @[Modules.scala 50:57:@14074.4]
  assign _T_66227 = $signed(buffer_0_340) + $signed(buffer_1_341); // @[Modules.scala 50:57:@14080.4]
  assign _T_66228 = _T_66227[10:0]; // @[Modules.scala 50:57:@14081.4]
  assign buffer_3_562 = $signed(_T_66228); // @[Modules.scala 50:57:@14082.4]
  assign buffer_3_342 = {{6{_T_65505[4]}},_T_65505}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_343 = {{6{_T_65508[4]}},_T_65508}; // @[Modules.scala 32:22:@8.4]
  assign _T_66230 = $signed(buffer_3_342) + $signed(buffer_3_343); // @[Modules.scala 50:57:@14084.4]
  assign _T_66231 = _T_66230[10:0]; // @[Modules.scala 50:57:@14085.4]
  assign buffer_3_563 = $signed(_T_66231); // @[Modules.scala 50:57:@14086.4]
  assign buffer_3_344 = {{6{_T_65515[4]}},_T_65515}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_345 = {{6{_T_65522[4]}},_T_65522}; // @[Modules.scala 32:22:@8.4]
  assign _T_66233 = $signed(buffer_3_344) + $signed(buffer_3_345); // @[Modules.scala 50:57:@14088.4]
  assign _T_66234 = _T_66233[10:0]; // @[Modules.scala 50:57:@14089.4]
  assign buffer_3_564 = $signed(_T_66234); // @[Modules.scala 50:57:@14090.4]
  assign buffer_3_347 = {{6{_T_65536[4]}},_T_65536}; // @[Modules.scala 32:22:@8.4]
  assign _T_66236 = $signed(buffer_1_346) + $signed(buffer_3_347); // @[Modules.scala 50:57:@14092.4]
  assign _T_66237 = _T_66236[10:0]; // @[Modules.scala 50:57:@14093.4]
  assign buffer_3_565 = $signed(_T_66237); // @[Modules.scala 50:57:@14094.4]
  assign buffer_3_349 = {{6{_T_65546[4]}},_T_65546}; // @[Modules.scala 32:22:@8.4]
  assign _T_66239 = $signed(buffer_2_348) + $signed(buffer_3_349); // @[Modules.scala 50:57:@14096.4]
  assign _T_66240 = _T_66239[10:0]; // @[Modules.scala 50:57:@14097.4]
  assign buffer_3_566 = $signed(_T_66240); // @[Modules.scala 50:57:@14098.4]
  assign buffer_3_351 = {{6{_T_65560[4]}},_T_65560}; // @[Modules.scala 32:22:@8.4]
  assign _T_66242 = $signed(buffer_0_350) + $signed(buffer_3_351); // @[Modules.scala 50:57:@14100.4]
  assign _T_66243 = _T_66242[10:0]; // @[Modules.scala 50:57:@14101.4]
  assign buffer_3_567 = $signed(_T_66243); // @[Modules.scala 50:57:@14102.4]
  assign buffer_3_355 = {{6{_T_65572[4]}},_T_65572}; // @[Modules.scala 32:22:@8.4]
  assign _T_66248 = $signed(buffer_0_354) + $signed(buffer_3_355); // @[Modules.scala 50:57:@14108.4]
  assign _T_66249 = _T_66248[10:0]; // @[Modules.scala 50:57:@14109.4]
  assign buffer_3_569 = $signed(_T_66249); // @[Modules.scala 50:57:@14110.4]
  assign buffer_3_361 = {{6{_T_65602[4]}},_T_65602}; // @[Modules.scala 32:22:@8.4]
  assign _T_66257 = $signed(buffer_1_360) + $signed(buffer_3_361); // @[Modules.scala 50:57:@14120.4]
  assign _T_66258 = _T_66257[10:0]; // @[Modules.scala 50:57:@14121.4]
  assign buffer_3_572 = $signed(_T_66258); // @[Modules.scala 50:57:@14122.4]
  assign _T_66260 = $signed(buffer_0_362) + $signed(buffer_1_363); // @[Modules.scala 50:57:@14124.4]
  assign _T_66261 = _T_66260[10:0]; // @[Modules.scala 50:57:@14125.4]
  assign buffer_3_573 = $signed(_T_66261); // @[Modules.scala 50:57:@14126.4]
  assign buffer_3_365 = {{6{_T_65614[4]}},_T_65614}; // @[Modules.scala 32:22:@8.4]
  assign _T_66263 = $signed(buffer_2_364) + $signed(buffer_3_365); // @[Modules.scala 50:57:@14128.4]
  assign _T_66264 = _T_66263[10:0]; // @[Modules.scala 50:57:@14129.4]
  assign buffer_3_574 = $signed(_T_66264); // @[Modules.scala 50:57:@14130.4]
  assign buffer_3_368 = {{6{_T_65623[4]}},_T_65623}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_369 = {{6{_T_65626[4]}},_T_65626}; // @[Modules.scala 32:22:@8.4]
  assign _T_66269 = $signed(buffer_3_368) + $signed(buffer_3_369); // @[Modules.scala 50:57:@14136.4]
  assign _T_66270 = _T_66269[10:0]; // @[Modules.scala 50:57:@14137.4]
  assign buffer_3_576 = $signed(_T_66270); // @[Modules.scala 50:57:@14138.4]
  assign buffer_3_370 = {{6{_T_65629[4]}},_T_65629}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_371 = {{6{_T_65636[4]}},_T_65636}; // @[Modules.scala 32:22:@8.4]
  assign _T_66272 = $signed(buffer_3_370) + $signed(buffer_3_371); // @[Modules.scala 50:57:@14140.4]
  assign _T_66273 = _T_66272[10:0]; // @[Modules.scala 50:57:@14141.4]
  assign buffer_3_577 = $signed(_T_66273); // @[Modules.scala 50:57:@14142.4]
  assign buffer_3_372 = {{6{_T_65639[4]}},_T_65639}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_373 = {{6{_T_65642[4]}},_T_65642}; // @[Modules.scala 32:22:@8.4]
  assign _T_66275 = $signed(buffer_3_372) + $signed(buffer_3_373); // @[Modules.scala 50:57:@14144.4]
  assign _T_66276 = _T_66275[10:0]; // @[Modules.scala 50:57:@14145.4]
  assign buffer_3_578 = $signed(_T_66276); // @[Modules.scala 50:57:@14146.4]
  assign buffer_3_374 = {{6{_T_65649[4]}},_T_65649}; // @[Modules.scala 32:22:@8.4]
  assign _T_66278 = $signed(buffer_3_374) + $signed(buffer_0_375); // @[Modules.scala 50:57:@14148.4]
  assign _T_66279 = _T_66278[10:0]; // @[Modules.scala 50:57:@14149.4]
  assign buffer_3_579 = $signed(_T_66279); // @[Modules.scala 50:57:@14150.4]
  assign buffer_3_376 = {{6{_T_65655[4]}},_T_65655}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_377 = {{6{_T_65662[4]}},_T_65662}; // @[Modules.scala 32:22:@8.4]
  assign _T_66281 = $signed(buffer_3_376) + $signed(buffer_3_377); // @[Modules.scala 50:57:@14152.4]
  assign _T_66282 = _T_66281[10:0]; // @[Modules.scala 50:57:@14153.4]
  assign buffer_3_580 = $signed(_T_66282); // @[Modules.scala 50:57:@14154.4]
  assign buffer_3_378 = {{6{_T_65665[4]}},_T_65665}; // @[Modules.scala 32:22:@8.4]
  assign _T_66284 = $signed(buffer_3_378) + $signed(buffer_0_379); // @[Modules.scala 50:57:@14156.4]
  assign _T_66285 = _T_66284[10:0]; // @[Modules.scala 50:57:@14157.4]
  assign buffer_3_581 = $signed(_T_66285); // @[Modules.scala 50:57:@14158.4]
  assign buffer_3_382 = {{6{_T_65681[4]}},_T_65681}; // @[Modules.scala 32:22:@8.4]
  assign _T_66290 = $signed(buffer_3_382) + $signed(buffer_1_383); // @[Modules.scala 50:57:@14164.4]
  assign _T_66291 = _T_66290[10:0]; // @[Modules.scala 50:57:@14165.4]
  assign buffer_3_583 = $signed(_T_66291); // @[Modules.scala 50:57:@14166.4]
  assign buffer_3_384 = {{6{_T_65687[4]}},_T_65687}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_385 = {{6{_T_65690[4]}},_T_65690}; // @[Modules.scala 32:22:@8.4]
  assign _T_66293 = $signed(buffer_3_384) + $signed(buffer_3_385); // @[Modules.scala 50:57:@14168.4]
  assign _T_66294 = _T_66293[10:0]; // @[Modules.scala 50:57:@14169.4]
  assign buffer_3_584 = $signed(_T_66294); // @[Modules.scala 50:57:@14170.4]
  assign buffer_3_386 = {{6{_T_65693[4]}},_T_65693}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_387 = {{6{_T_65696[4]}},_T_65696}; // @[Modules.scala 32:22:@8.4]
  assign _T_66296 = $signed(buffer_3_386) + $signed(buffer_3_387); // @[Modules.scala 50:57:@14172.4]
  assign _T_66297 = _T_66296[10:0]; // @[Modules.scala 50:57:@14173.4]
  assign buffer_3_585 = $signed(_T_66297); // @[Modules.scala 50:57:@14174.4]
  assign buffer_3_389 = {{6{_T_65710[4]}},_T_65710}; // @[Modules.scala 32:22:@8.4]
  assign _T_66299 = $signed(buffer_1_388) + $signed(buffer_3_389); // @[Modules.scala 50:57:@14176.4]
  assign _T_66300 = _T_66299[10:0]; // @[Modules.scala 50:57:@14177.4]
  assign buffer_3_586 = $signed(_T_66300); // @[Modules.scala 50:57:@14178.4]
  assign _T_66302 = $signed(buffer_1_390) + $signed(buffer_0_391); // @[Modules.scala 50:57:@14180.4]
  assign _T_66303 = _T_66302[10:0]; // @[Modules.scala 50:57:@14181.4]
  assign buffer_3_587 = $signed(_T_66303); // @[Modules.scala 50:57:@14182.4]
  assign _T_66305 = $signed(buffer_3_392) + $signed(buffer_1_393); // @[Modules.scala 53:83:@14184.4]
  assign _T_66306 = _T_66305[10:0]; // @[Modules.scala 53:83:@14185.4]
  assign buffer_3_588 = $signed(_T_66306); // @[Modules.scala 53:83:@14186.4]
  assign _T_66308 = $signed(buffer_3_394) + $signed(buffer_1_395); // @[Modules.scala 53:83:@14188.4]
  assign _T_66309 = _T_66308[10:0]; // @[Modules.scala 53:83:@14189.4]
  assign buffer_3_589 = $signed(_T_66309); // @[Modules.scala 53:83:@14190.4]
  assign _T_66311 = $signed(buffer_3_396) + $signed(buffer_3_397); // @[Modules.scala 53:83:@14192.4]
  assign _T_66312 = _T_66311[10:0]; // @[Modules.scala 53:83:@14193.4]
  assign buffer_3_590 = $signed(_T_66312); // @[Modules.scala 53:83:@14194.4]
  assign _T_66314 = $signed(buffer_3_398) + $signed(buffer_3_399); // @[Modules.scala 53:83:@14196.4]
  assign _T_66315 = _T_66314[10:0]; // @[Modules.scala 53:83:@14197.4]
  assign buffer_3_591 = $signed(_T_66315); // @[Modules.scala 53:83:@14198.4]
  assign _T_66317 = $signed(buffer_3_400) + $signed(buffer_1_401); // @[Modules.scala 53:83:@14200.4]
  assign _T_66318 = _T_66317[10:0]; // @[Modules.scala 53:83:@14201.4]
  assign buffer_3_592 = $signed(_T_66318); // @[Modules.scala 53:83:@14202.4]
  assign _T_66320 = $signed(buffer_0_402) + $signed(buffer_3_403); // @[Modules.scala 53:83:@14204.4]
  assign _T_66321 = _T_66320[10:0]; // @[Modules.scala 53:83:@14205.4]
  assign buffer_3_593 = $signed(_T_66321); // @[Modules.scala 53:83:@14206.4]
  assign _T_66323 = $signed(buffer_3_404) + $signed(buffer_3_405); // @[Modules.scala 53:83:@14208.4]
  assign _T_66324 = _T_66323[10:0]; // @[Modules.scala 53:83:@14209.4]
  assign buffer_3_594 = $signed(_T_66324); // @[Modules.scala 53:83:@14210.4]
  assign _T_66326 = $signed(buffer_3_406) + $signed(buffer_3_407); // @[Modules.scala 53:83:@14212.4]
  assign _T_66327 = _T_66326[10:0]; // @[Modules.scala 53:83:@14213.4]
  assign buffer_3_595 = $signed(_T_66327); // @[Modules.scala 53:83:@14214.4]
  assign _T_66329 = $signed(buffer_3_408) + $signed(buffer_0_409); // @[Modules.scala 53:83:@14216.4]
  assign _T_66330 = _T_66329[10:0]; // @[Modules.scala 53:83:@14217.4]
  assign buffer_3_596 = $signed(_T_66330); // @[Modules.scala 53:83:@14218.4]
  assign _T_66332 = $signed(buffer_3_410) + $signed(buffer_3_411); // @[Modules.scala 53:83:@14220.4]
  assign _T_66333 = _T_66332[10:0]; // @[Modules.scala 53:83:@14221.4]
  assign buffer_3_597 = $signed(_T_66333); // @[Modules.scala 53:83:@14222.4]
  assign _T_66335 = $signed(buffer_3_412) + $signed(buffer_3_413); // @[Modules.scala 53:83:@14224.4]
  assign _T_66336 = _T_66335[10:0]; // @[Modules.scala 53:83:@14225.4]
  assign buffer_3_598 = $signed(_T_66336); // @[Modules.scala 53:83:@14226.4]
  assign _T_66338 = $signed(buffer_3_414) + $signed(buffer_3_415); // @[Modules.scala 53:83:@14228.4]
  assign _T_66339 = _T_66338[10:0]; // @[Modules.scala 53:83:@14229.4]
  assign buffer_3_599 = $signed(_T_66339); // @[Modules.scala 53:83:@14230.4]
  assign _T_66341 = $signed(buffer_3_416) + $signed(buffer_3_417); // @[Modules.scala 53:83:@14232.4]
  assign _T_66342 = _T_66341[10:0]; // @[Modules.scala 53:83:@14233.4]
  assign buffer_3_600 = $signed(_T_66342); // @[Modules.scala 53:83:@14234.4]
  assign _T_66344 = $signed(buffer_3_418) + $signed(buffer_3_419); // @[Modules.scala 53:83:@14236.4]
  assign _T_66345 = _T_66344[10:0]; // @[Modules.scala 53:83:@14237.4]
  assign buffer_3_601 = $signed(_T_66345); // @[Modules.scala 53:83:@14238.4]
  assign _T_66347 = $signed(buffer_3_420) + $signed(buffer_3_421); // @[Modules.scala 53:83:@14240.4]
  assign _T_66348 = _T_66347[10:0]; // @[Modules.scala 53:83:@14241.4]
  assign buffer_3_602 = $signed(_T_66348); // @[Modules.scala 53:83:@14242.4]
  assign _T_66350 = $signed(buffer_3_422) + $signed(buffer_3_423); // @[Modules.scala 53:83:@14244.4]
  assign _T_66351 = _T_66350[10:0]; // @[Modules.scala 53:83:@14245.4]
  assign buffer_3_603 = $signed(_T_66351); // @[Modules.scala 53:83:@14246.4]
  assign _T_66353 = $signed(buffer_1_424) + $signed(buffer_3_425); // @[Modules.scala 53:83:@14248.4]
  assign _T_66354 = _T_66353[10:0]; // @[Modules.scala 53:83:@14249.4]
  assign buffer_3_604 = $signed(_T_66354); // @[Modules.scala 53:83:@14250.4]
  assign _T_66356 = $signed(buffer_3_426) + $signed(buffer_3_427); // @[Modules.scala 53:83:@14252.4]
  assign _T_66357 = _T_66356[10:0]; // @[Modules.scala 53:83:@14253.4]
  assign buffer_3_605 = $signed(_T_66357); // @[Modules.scala 53:83:@14254.4]
  assign _T_66359 = $signed(buffer_3_428) + $signed(buffer_3_429); // @[Modules.scala 53:83:@14256.4]
  assign _T_66360 = _T_66359[10:0]; // @[Modules.scala 53:83:@14257.4]
  assign buffer_3_606 = $signed(_T_66360); // @[Modules.scala 53:83:@14258.4]
  assign _T_66362 = $signed(buffer_3_430) + $signed(buffer_3_431); // @[Modules.scala 53:83:@14260.4]
  assign _T_66363 = _T_66362[10:0]; // @[Modules.scala 53:83:@14261.4]
  assign buffer_3_607 = $signed(_T_66363); // @[Modules.scala 53:83:@14262.4]
  assign _T_66368 = $signed(buffer_1_434) + $signed(buffer_3_435); // @[Modules.scala 53:83:@14268.4]
  assign _T_66369 = _T_66368[10:0]; // @[Modules.scala 53:83:@14269.4]
  assign buffer_3_609 = $signed(_T_66369); // @[Modules.scala 53:83:@14270.4]
  assign _T_66371 = $signed(buffer_3_436) + $signed(buffer_3_437); // @[Modules.scala 53:83:@14272.4]
  assign _T_66372 = _T_66371[10:0]; // @[Modules.scala 53:83:@14273.4]
  assign buffer_3_610 = $signed(_T_66372); // @[Modules.scala 53:83:@14274.4]
  assign _T_66374 = $signed(buffer_3_438) + $signed(buffer_3_439); // @[Modules.scala 53:83:@14276.4]
  assign _T_66375 = _T_66374[10:0]; // @[Modules.scala 53:83:@14277.4]
  assign buffer_3_611 = $signed(_T_66375); // @[Modules.scala 53:83:@14278.4]
  assign _T_66377 = $signed(buffer_2_440) + $signed(buffer_3_441); // @[Modules.scala 53:83:@14280.4]
  assign _T_66378 = _T_66377[10:0]; // @[Modules.scala 53:83:@14281.4]
  assign buffer_3_612 = $signed(_T_66378); // @[Modules.scala 53:83:@14282.4]
  assign _T_66380 = $signed(buffer_3_442) + $signed(buffer_3_443); // @[Modules.scala 53:83:@14284.4]
  assign _T_66381 = _T_66380[10:0]; // @[Modules.scala 53:83:@14285.4]
  assign buffer_3_613 = $signed(_T_66381); // @[Modules.scala 53:83:@14286.4]
  assign _T_66383 = $signed(buffer_3_444) + $signed(buffer_3_445); // @[Modules.scala 53:83:@14288.4]
  assign _T_66384 = _T_66383[10:0]; // @[Modules.scala 53:83:@14289.4]
  assign buffer_3_614 = $signed(_T_66384); // @[Modules.scala 53:83:@14290.4]
  assign _T_66386 = $signed(buffer_3_446) + $signed(buffer_2_447); // @[Modules.scala 53:83:@14292.4]
  assign _T_66387 = _T_66386[10:0]; // @[Modules.scala 53:83:@14293.4]
  assign buffer_3_615 = $signed(_T_66387); // @[Modules.scala 53:83:@14294.4]
  assign _T_66389 = $signed(buffer_3_448) + $signed(buffer_3_449); // @[Modules.scala 53:83:@14296.4]
  assign _T_66390 = _T_66389[10:0]; // @[Modules.scala 53:83:@14297.4]
  assign buffer_3_616 = $signed(_T_66390); // @[Modules.scala 53:83:@14298.4]
  assign _T_66392 = $signed(buffer_3_450) + $signed(buffer_3_451); // @[Modules.scala 53:83:@14300.4]
  assign _T_66393 = _T_66392[10:0]; // @[Modules.scala 53:83:@14301.4]
  assign buffer_3_617 = $signed(_T_66393); // @[Modules.scala 53:83:@14302.4]
  assign _T_66395 = $signed(buffer_3_452) + $signed(buffer_3_453); // @[Modules.scala 53:83:@14304.4]
  assign _T_66396 = _T_66395[10:0]; // @[Modules.scala 53:83:@14305.4]
  assign buffer_3_618 = $signed(_T_66396); // @[Modules.scala 53:83:@14306.4]
  assign _T_66398 = $signed(buffer_1_454) + $signed(buffer_3_455); // @[Modules.scala 53:83:@14308.4]
  assign _T_66399 = _T_66398[10:0]; // @[Modules.scala 53:83:@14309.4]
  assign buffer_3_619 = $signed(_T_66399); // @[Modules.scala 53:83:@14310.4]
  assign _T_66401 = $signed(buffer_3_456) + $signed(buffer_2_457); // @[Modules.scala 53:83:@14312.4]
  assign _T_66402 = _T_66401[10:0]; // @[Modules.scala 53:83:@14313.4]
  assign buffer_3_620 = $signed(_T_66402); // @[Modules.scala 53:83:@14314.4]
  assign _T_66404 = $signed(buffer_3_458) + $signed(buffer_3_459); // @[Modules.scala 53:83:@14316.4]
  assign _T_66405 = _T_66404[10:0]; // @[Modules.scala 53:83:@14317.4]
  assign buffer_3_621 = $signed(_T_66405); // @[Modules.scala 53:83:@14318.4]
  assign _T_66407 = $signed(buffer_3_460) + $signed(buffer_1_461); // @[Modules.scala 53:83:@14320.4]
  assign _T_66408 = _T_66407[10:0]; // @[Modules.scala 53:83:@14321.4]
  assign buffer_3_622 = $signed(_T_66408); // @[Modules.scala 53:83:@14322.4]
  assign _T_66410 = $signed(buffer_3_462) + $signed(buffer_3_463); // @[Modules.scala 53:83:@14324.4]
  assign _T_66411 = _T_66410[10:0]; // @[Modules.scala 53:83:@14325.4]
  assign buffer_3_623 = $signed(_T_66411); // @[Modules.scala 53:83:@14326.4]
  assign _T_66413 = $signed(buffer_3_464) + $signed(buffer_3_465); // @[Modules.scala 53:83:@14328.4]
  assign _T_66414 = _T_66413[10:0]; // @[Modules.scala 53:83:@14329.4]
  assign buffer_3_624 = $signed(_T_66414); // @[Modules.scala 53:83:@14330.4]
  assign _T_66416 = $signed(buffer_3_466) + $signed(buffer_3_467); // @[Modules.scala 53:83:@14332.4]
  assign _T_66417 = _T_66416[10:0]; // @[Modules.scala 53:83:@14333.4]
  assign buffer_3_625 = $signed(_T_66417); // @[Modules.scala 53:83:@14334.4]
  assign _T_66419 = $signed(buffer_1_468) + $signed(buffer_3_469); // @[Modules.scala 53:83:@14336.4]
  assign _T_66420 = _T_66419[10:0]; // @[Modules.scala 53:83:@14337.4]
  assign buffer_3_626 = $signed(_T_66420); // @[Modules.scala 53:83:@14338.4]
  assign _T_66422 = $signed(buffer_3_470) + $signed(buffer_3_471); // @[Modules.scala 53:83:@14340.4]
  assign _T_66423 = _T_66422[10:0]; // @[Modules.scala 53:83:@14341.4]
  assign buffer_3_627 = $signed(_T_66423); // @[Modules.scala 53:83:@14342.4]
  assign _T_66425 = $signed(buffer_0_472) + $signed(buffer_1_473); // @[Modules.scala 53:83:@14344.4]
  assign _T_66426 = _T_66425[10:0]; // @[Modules.scala 53:83:@14345.4]
  assign buffer_3_628 = $signed(_T_66426); // @[Modules.scala 53:83:@14346.4]
  assign _T_66428 = $signed(buffer_2_474) + $signed(buffer_3_475); // @[Modules.scala 53:83:@14348.4]
  assign _T_66429 = _T_66428[10:0]; // @[Modules.scala 53:83:@14349.4]
  assign buffer_3_629 = $signed(_T_66429); // @[Modules.scala 53:83:@14350.4]
  assign _T_66431 = $signed(buffer_3_476) + $signed(buffer_3_477); // @[Modules.scala 53:83:@14352.4]
  assign _T_66432 = _T_66431[10:0]; // @[Modules.scala 53:83:@14353.4]
  assign buffer_3_630 = $signed(_T_66432); // @[Modules.scala 53:83:@14354.4]
  assign _T_66434 = $signed(buffer_3_478) + $signed(buffer_3_479); // @[Modules.scala 53:83:@14356.4]
  assign _T_66435 = _T_66434[10:0]; // @[Modules.scala 53:83:@14357.4]
  assign buffer_3_631 = $signed(_T_66435); // @[Modules.scala 53:83:@14358.4]
  assign _T_66440 = $signed(buffer_3_482) + $signed(buffer_3_483); // @[Modules.scala 53:83:@14364.4]
  assign _T_66441 = _T_66440[10:0]; // @[Modules.scala 53:83:@14365.4]
  assign buffer_3_633 = $signed(_T_66441); // @[Modules.scala 53:83:@14366.4]
  assign _T_66443 = $signed(buffer_3_484) + $signed(buffer_3_485); // @[Modules.scala 53:83:@14368.4]
  assign _T_66444 = _T_66443[10:0]; // @[Modules.scala 53:83:@14369.4]
  assign buffer_3_634 = $signed(_T_66444); // @[Modules.scala 53:83:@14370.4]
  assign _T_66446 = $signed(buffer_3_486) + $signed(buffer_3_487); // @[Modules.scala 53:83:@14372.4]
  assign _T_66447 = _T_66446[10:0]; // @[Modules.scala 53:83:@14373.4]
  assign buffer_3_635 = $signed(_T_66447); // @[Modules.scala 53:83:@14374.4]
  assign _T_66449 = $signed(buffer_3_488) + $signed(buffer_3_489); // @[Modules.scala 53:83:@14376.4]
  assign _T_66450 = _T_66449[10:0]; // @[Modules.scala 53:83:@14377.4]
  assign buffer_3_636 = $signed(_T_66450); // @[Modules.scala 53:83:@14378.4]
  assign _T_66452 = $signed(buffer_3_490) + $signed(buffer_3_491); // @[Modules.scala 53:83:@14380.4]
  assign _T_66453 = _T_66452[10:0]; // @[Modules.scala 53:83:@14381.4]
  assign buffer_3_637 = $signed(_T_66453); // @[Modules.scala 53:83:@14382.4]
  assign _T_66455 = $signed(buffer_3_492) + $signed(buffer_3_493); // @[Modules.scala 53:83:@14384.4]
  assign _T_66456 = _T_66455[10:0]; // @[Modules.scala 53:83:@14385.4]
  assign buffer_3_638 = $signed(_T_66456); // @[Modules.scala 53:83:@14386.4]
  assign _T_66458 = $signed(buffer_3_494) + $signed(buffer_3_495); // @[Modules.scala 53:83:@14388.4]
  assign _T_66459 = _T_66458[10:0]; // @[Modules.scala 53:83:@14389.4]
  assign buffer_3_639 = $signed(_T_66459); // @[Modules.scala 53:83:@14390.4]
  assign _T_66461 = $signed(buffer_3_496) + $signed(buffer_3_497); // @[Modules.scala 53:83:@14392.4]
  assign _T_66462 = _T_66461[10:0]; // @[Modules.scala 53:83:@14393.4]
  assign buffer_3_640 = $signed(_T_66462); // @[Modules.scala 53:83:@14394.4]
  assign _T_66464 = $signed(buffer_3_498) + $signed(buffer_2_499); // @[Modules.scala 53:83:@14396.4]
  assign _T_66465 = _T_66464[10:0]; // @[Modules.scala 53:83:@14397.4]
  assign buffer_3_641 = $signed(_T_66465); // @[Modules.scala 53:83:@14398.4]
  assign _T_66467 = $signed(buffer_1_500) + $signed(buffer_2_501); // @[Modules.scala 53:83:@14400.4]
  assign _T_66468 = _T_66467[10:0]; // @[Modules.scala 53:83:@14401.4]
  assign buffer_3_642 = $signed(_T_66468); // @[Modules.scala 53:83:@14402.4]
  assign _T_66470 = $signed(buffer_3_502) + $signed(buffer_3_503); // @[Modules.scala 53:83:@14404.4]
  assign _T_66471 = _T_66470[10:0]; // @[Modules.scala 53:83:@14405.4]
  assign buffer_3_643 = $signed(_T_66471); // @[Modules.scala 53:83:@14406.4]
  assign _T_66473 = $signed(buffer_3_504) + $signed(buffer_3_505); // @[Modules.scala 53:83:@14408.4]
  assign _T_66474 = _T_66473[10:0]; // @[Modules.scala 53:83:@14409.4]
  assign buffer_3_644 = $signed(_T_66474); // @[Modules.scala 53:83:@14410.4]
  assign _T_66476 = $signed(buffer_3_506) + $signed(buffer_1_507); // @[Modules.scala 53:83:@14412.4]
  assign _T_66477 = _T_66476[10:0]; // @[Modules.scala 53:83:@14413.4]
  assign buffer_3_645 = $signed(_T_66477); // @[Modules.scala 53:83:@14414.4]
  assign _T_66479 = $signed(buffer_3_508) + $signed(buffer_1_509); // @[Modules.scala 53:83:@14416.4]
  assign _T_66480 = _T_66479[10:0]; // @[Modules.scala 53:83:@14417.4]
  assign buffer_3_646 = $signed(_T_66480); // @[Modules.scala 53:83:@14418.4]
  assign _T_66482 = $signed(buffer_3_510) + $signed(buffer_3_511); // @[Modules.scala 53:83:@14420.4]
  assign _T_66483 = _T_66482[10:0]; // @[Modules.scala 53:83:@14421.4]
  assign buffer_3_647 = $signed(_T_66483); // @[Modules.scala 53:83:@14422.4]
  assign _T_66485 = $signed(buffer_3_512) + $signed(buffer_1_513); // @[Modules.scala 53:83:@14424.4]
  assign _T_66486 = _T_66485[10:0]; // @[Modules.scala 53:83:@14425.4]
  assign buffer_3_648 = $signed(_T_66486); // @[Modules.scala 53:83:@14426.4]
  assign _T_66488 = $signed(buffer_1_514) + $signed(buffer_3_515); // @[Modules.scala 53:83:@14428.4]
  assign _T_66489 = _T_66488[10:0]; // @[Modules.scala 53:83:@14429.4]
  assign buffer_3_649 = $signed(_T_66489); // @[Modules.scala 53:83:@14430.4]
  assign _T_66491 = $signed(buffer_1_516) + $signed(buffer_3_517); // @[Modules.scala 53:83:@14432.4]
  assign _T_66492 = _T_66491[10:0]; // @[Modules.scala 53:83:@14433.4]
  assign buffer_3_650 = $signed(_T_66492); // @[Modules.scala 53:83:@14434.4]
  assign _T_66494 = $signed(buffer_3_518) + $signed(buffer_3_519); // @[Modules.scala 53:83:@14436.4]
  assign _T_66495 = _T_66494[10:0]; // @[Modules.scala 53:83:@14437.4]
  assign buffer_3_651 = $signed(_T_66495); // @[Modules.scala 53:83:@14438.4]
  assign _T_66497 = $signed(buffer_3_520) + $signed(buffer_1_521); // @[Modules.scala 53:83:@14440.4]
  assign _T_66498 = _T_66497[10:0]; // @[Modules.scala 53:83:@14441.4]
  assign buffer_3_652 = $signed(_T_66498); // @[Modules.scala 53:83:@14442.4]
  assign _T_66500 = $signed(buffer_1_522) + $signed(buffer_0_523); // @[Modules.scala 53:83:@14444.4]
  assign _T_66501 = _T_66500[10:0]; // @[Modules.scala 53:83:@14445.4]
  assign buffer_3_653 = $signed(_T_66501); // @[Modules.scala 53:83:@14446.4]
  assign _T_66503 = $signed(buffer_3_524) + $signed(buffer_1_525); // @[Modules.scala 53:83:@14448.4]
  assign _T_66504 = _T_66503[10:0]; // @[Modules.scala 53:83:@14449.4]
  assign buffer_3_654 = $signed(_T_66504); // @[Modules.scala 53:83:@14450.4]
  assign _T_66506 = $signed(buffer_1_526) + $signed(buffer_3_527); // @[Modules.scala 53:83:@14452.4]
  assign _T_66507 = _T_66506[10:0]; // @[Modules.scala 53:83:@14453.4]
  assign buffer_3_655 = $signed(_T_66507); // @[Modules.scala 53:83:@14454.4]
  assign _T_66509 = $signed(buffer_3_528) + $signed(buffer_3_529); // @[Modules.scala 53:83:@14456.4]
  assign _T_66510 = _T_66509[10:0]; // @[Modules.scala 53:83:@14457.4]
  assign buffer_3_656 = $signed(_T_66510); // @[Modules.scala 53:83:@14458.4]
  assign _T_66512 = $signed(buffer_3_530) + $signed(buffer_3_531); // @[Modules.scala 53:83:@14460.4]
  assign _T_66513 = _T_66512[10:0]; // @[Modules.scala 53:83:@14461.4]
  assign buffer_3_657 = $signed(_T_66513); // @[Modules.scala 53:83:@14462.4]
  assign _T_66515 = $signed(buffer_3_532) + $signed(buffer_3_533); // @[Modules.scala 53:83:@14464.4]
  assign _T_66516 = _T_66515[10:0]; // @[Modules.scala 53:83:@14465.4]
  assign buffer_3_658 = $signed(_T_66516); // @[Modules.scala 53:83:@14466.4]
  assign _T_66518 = $signed(buffer_1_534) + $signed(buffer_3_535); // @[Modules.scala 53:83:@14468.4]
  assign _T_66519 = _T_66518[10:0]; // @[Modules.scala 53:83:@14469.4]
  assign buffer_3_659 = $signed(_T_66519); // @[Modules.scala 53:83:@14470.4]
  assign _T_66521 = $signed(buffer_3_536) + $signed(buffer_3_537); // @[Modules.scala 53:83:@14472.4]
  assign _T_66522 = _T_66521[10:0]; // @[Modules.scala 53:83:@14473.4]
  assign buffer_3_660 = $signed(_T_66522); // @[Modules.scala 53:83:@14474.4]
  assign _T_66524 = $signed(buffer_3_538) + $signed(buffer_1_539); // @[Modules.scala 53:83:@14476.4]
  assign _T_66525 = _T_66524[10:0]; // @[Modules.scala 53:83:@14477.4]
  assign buffer_3_661 = $signed(_T_66525); // @[Modules.scala 53:83:@14478.4]
  assign _T_66527 = $signed(buffer_3_540) + $signed(buffer_3_541); // @[Modules.scala 53:83:@14480.4]
  assign _T_66528 = _T_66527[10:0]; // @[Modules.scala 53:83:@14481.4]
  assign buffer_3_662 = $signed(_T_66528); // @[Modules.scala 53:83:@14482.4]
  assign _T_66530 = $signed(buffer_3_542) + $signed(buffer_3_543); // @[Modules.scala 53:83:@14484.4]
  assign _T_66531 = _T_66530[10:0]; // @[Modules.scala 53:83:@14485.4]
  assign buffer_3_663 = $signed(_T_66531); // @[Modules.scala 53:83:@14486.4]
  assign _T_66533 = $signed(buffer_3_544) + $signed(buffer_3_545); // @[Modules.scala 53:83:@14488.4]
  assign _T_66534 = _T_66533[10:0]; // @[Modules.scala 53:83:@14489.4]
  assign buffer_3_664 = $signed(_T_66534); // @[Modules.scala 53:83:@14490.4]
  assign _T_66536 = $signed(buffer_1_546) + $signed(buffer_3_547); // @[Modules.scala 53:83:@14492.4]
  assign _T_66537 = _T_66536[10:0]; // @[Modules.scala 53:83:@14493.4]
  assign buffer_3_665 = $signed(_T_66537); // @[Modules.scala 53:83:@14494.4]
  assign _T_66539 = $signed(buffer_3_548) + $signed(buffer_3_549); // @[Modules.scala 53:83:@14496.4]
  assign _T_66540 = _T_66539[10:0]; // @[Modules.scala 53:83:@14497.4]
  assign buffer_3_666 = $signed(_T_66540); // @[Modules.scala 53:83:@14498.4]
  assign _T_66542 = $signed(buffer_3_550) + $signed(buffer_3_551); // @[Modules.scala 53:83:@14500.4]
  assign _T_66543 = _T_66542[10:0]; // @[Modules.scala 53:83:@14501.4]
  assign buffer_3_667 = $signed(_T_66543); // @[Modules.scala 53:83:@14502.4]
  assign _T_66545 = $signed(buffer_3_552) + $signed(buffer_3_553); // @[Modules.scala 53:83:@14504.4]
  assign _T_66546 = _T_66545[10:0]; // @[Modules.scala 53:83:@14505.4]
  assign buffer_3_668 = $signed(_T_66546); // @[Modules.scala 53:83:@14506.4]
  assign _T_66548 = $signed(buffer_3_554) + $signed(buffer_3_555); // @[Modules.scala 53:83:@14508.4]
  assign _T_66549 = _T_66548[10:0]; // @[Modules.scala 53:83:@14509.4]
  assign buffer_3_669 = $signed(_T_66549); // @[Modules.scala 53:83:@14510.4]
  assign _T_66551 = $signed(buffer_3_556) + $signed(buffer_3_557); // @[Modules.scala 53:83:@14512.4]
  assign _T_66552 = _T_66551[10:0]; // @[Modules.scala 53:83:@14513.4]
  assign buffer_3_670 = $signed(_T_66552); // @[Modules.scala 53:83:@14514.4]
  assign _T_66554 = $signed(buffer_3_558) + $signed(buffer_3_559); // @[Modules.scala 53:83:@14516.4]
  assign _T_66555 = _T_66554[10:0]; // @[Modules.scala 53:83:@14517.4]
  assign buffer_3_671 = $signed(_T_66555); // @[Modules.scala 53:83:@14518.4]
  assign _T_66557 = $signed(buffer_3_560) + $signed(buffer_0_561); // @[Modules.scala 53:83:@14520.4]
  assign _T_66558 = _T_66557[10:0]; // @[Modules.scala 53:83:@14521.4]
  assign buffer_3_672 = $signed(_T_66558); // @[Modules.scala 53:83:@14522.4]
  assign _T_66560 = $signed(buffer_3_562) + $signed(buffer_3_563); // @[Modules.scala 53:83:@14524.4]
  assign _T_66561 = _T_66560[10:0]; // @[Modules.scala 53:83:@14525.4]
  assign buffer_3_673 = $signed(_T_66561); // @[Modules.scala 53:83:@14526.4]
  assign _T_66563 = $signed(buffer_3_564) + $signed(buffer_3_565); // @[Modules.scala 53:83:@14528.4]
  assign _T_66564 = _T_66563[10:0]; // @[Modules.scala 53:83:@14529.4]
  assign buffer_3_674 = $signed(_T_66564); // @[Modules.scala 53:83:@14530.4]
  assign _T_66566 = $signed(buffer_3_566) + $signed(buffer_3_567); // @[Modules.scala 53:83:@14532.4]
  assign _T_66567 = _T_66566[10:0]; // @[Modules.scala 53:83:@14533.4]
  assign buffer_3_675 = $signed(_T_66567); // @[Modules.scala 53:83:@14534.4]
  assign _T_66569 = $signed(buffer_0_568) + $signed(buffer_3_569); // @[Modules.scala 53:83:@14536.4]
  assign _T_66570 = _T_66569[10:0]; // @[Modules.scala 53:83:@14537.4]
  assign buffer_3_676 = $signed(_T_66570); // @[Modules.scala 53:83:@14538.4]
  assign _T_66572 = $signed(buffer_0_570) + $signed(buffer_1_571); // @[Modules.scala 53:83:@14540.4]
  assign _T_66573 = _T_66572[10:0]; // @[Modules.scala 53:83:@14541.4]
  assign buffer_3_677 = $signed(_T_66573); // @[Modules.scala 53:83:@14542.4]
  assign _T_66575 = $signed(buffer_3_572) + $signed(buffer_3_573); // @[Modules.scala 53:83:@14544.4]
  assign _T_66576 = _T_66575[10:0]; // @[Modules.scala 53:83:@14545.4]
  assign buffer_3_678 = $signed(_T_66576); // @[Modules.scala 53:83:@14546.4]
  assign _T_66578 = $signed(buffer_3_574) + $signed(buffer_0_575); // @[Modules.scala 53:83:@14548.4]
  assign _T_66579 = _T_66578[10:0]; // @[Modules.scala 53:83:@14549.4]
  assign buffer_3_679 = $signed(_T_66579); // @[Modules.scala 53:83:@14550.4]
  assign _T_66581 = $signed(buffer_3_576) + $signed(buffer_3_577); // @[Modules.scala 53:83:@14552.4]
  assign _T_66582 = _T_66581[10:0]; // @[Modules.scala 53:83:@14553.4]
  assign buffer_3_680 = $signed(_T_66582); // @[Modules.scala 53:83:@14554.4]
  assign _T_66584 = $signed(buffer_3_578) + $signed(buffer_3_579); // @[Modules.scala 53:83:@14556.4]
  assign _T_66585 = _T_66584[10:0]; // @[Modules.scala 53:83:@14557.4]
  assign buffer_3_681 = $signed(_T_66585); // @[Modules.scala 53:83:@14558.4]
  assign _T_66587 = $signed(buffer_3_580) + $signed(buffer_3_581); // @[Modules.scala 53:83:@14560.4]
  assign _T_66588 = _T_66587[10:0]; // @[Modules.scala 53:83:@14561.4]
  assign buffer_3_682 = $signed(_T_66588); // @[Modules.scala 53:83:@14562.4]
  assign _T_66590 = $signed(buffer_1_582) + $signed(buffer_3_583); // @[Modules.scala 53:83:@14564.4]
  assign _T_66591 = _T_66590[10:0]; // @[Modules.scala 53:83:@14565.4]
  assign buffer_3_683 = $signed(_T_66591); // @[Modules.scala 53:83:@14566.4]
  assign _T_66593 = $signed(buffer_3_584) + $signed(buffer_3_585); // @[Modules.scala 53:83:@14568.4]
  assign _T_66594 = _T_66593[10:0]; // @[Modules.scala 53:83:@14569.4]
  assign buffer_3_684 = $signed(_T_66594); // @[Modules.scala 53:83:@14570.4]
  assign _T_66596 = $signed(buffer_3_586) + $signed(buffer_3_587); // @[Modules.scala 53:83:@14572.4]
  assign _T_66597 = _T_66596[10:0]; // @[Modules.scala 53:83:@14573.4]
  assign buffer_3_685 = $signed(_T_66597); // @[Modules.scala 53:83:@14574.4]
  assign _T_66599 = $signed(buffer_3_588) + $signed(buffer_3_589); // @[Modules.scala 56:109:@14576.4]
  assign _T_66600 = _T_66599[10:0]; // @[Modules.scala 56:109:@14577.4]
  assign buffer_3_686 = $signed(_T_66600); // @[Modules.scala 56:109:@14578.4]
  assign _T_66602 = $signed(buffer_3_590) + $signed(buffer_3_591); // @[Modules.scala 56:109:@14580.4]
  assign _T_66603 = _T_66602[10:0]; // @[Modules.scala 56:109:@14581.4]
  assign buffer_3_687 = $signed(_T_66603); // @[Modules.scala 56:109:@14582.4]
  assign _T_66605 = $signed(buffer_3_592) + $signed(buffer_3_593); // @[Modules.scala 56:109:@14584.4]
  assign _T_66606 = _T_66605[10:0]; // @[Modules.scala 56:109:@14585.4]
  assign buffer_3_688 = $signed(_T_66606); // @[Modules.scala 56:109:@14586.4]
  assign _T_66608 = $signed(buffer_3_594) + $signed(buffer_3_595); // @[Modules.scala 56:109:@14588.4]
  assign _T_66609 = _T_66608[10:0]; // @[Modules.scala 56:109:@14589.4]
  assign buffer_3_689 = $signed(_T_66609); // @[Modules.scala 56:109:@14590.4]
  assign _T_66611 = $signed(buffer_3_596) + $signed(buffer_3_597); // @[Modules.scala 56:109:@14592.4]
  assign _T_66612 = _T_66611[10:0]; // @[Modules.scala 56:109:@14593.4]
  assign buffer_3_690 = $signed(_T_66612); // @[Modules.scala 56:109:@14594.4]
  assign _T_66614 = $signed(buffer_3_598) + $signed(buffer_3_599); // @[Modules.scala 56:109:@14596.4]
  assign _T_66615 = _T_66614[10:0]; // @[Modules.scala 56:109:@14597.4]
  assign buffer_3_691 = $signed(_T_66615); // @[Modules.scala 56:109:@14598.4]
  assign _T_66617 = $signed(buffer_3_600) + $signed(buffer_3_601); // @[Modules.scala 56:109:@14600.4]
  assign _T_66618 = _T_66617[10:0]; // @[Modules.scala 56:109:@14601.4]
  assign buffer_3_692 = $signed(_T_66618); // @[Modules.scala 56:109:@14602.4]
  assign _T_66620 = $signed(buffer_3_602) + $signed(buffer_3_603); // @[Modules.scala 56:109:@14604.4]
  assign _T_66621 = _T_66620[10:0]; // @[Modules.scala 56:109:@14605.4]
  assign buffer_3_693 = $signed(_T_66621); // @[Modules.scala 56:109:@14606.4]
  assign _T_66623 = $signed(buffer_3_604) + $signed(buffer_3_605); // @[Modules.scala 56:109:@14608.4]
  assign _T_66624 = _T_66623[10:0]; // @[Modules.scala 56:109:@14609.4]
  assign buffer_3_694 = $signed(_T_66624); // @[Modules.scala 56:109:@14610.4]
  assign _T_66626 = $signed(buffer_3_606) + $signed(buffer_3_607); // @[Modules.scala 56:109:@14612.4]
  assign _T_66627 = _T_66626[10:0]; // @[Modules.scala 56:109:@14613.4]
  assign buffer_3_695 = $signed(_T_66627); // @[Modules.scala 56:109:@14614.4]
  assign _T_66629 = $signed(buffer_2_608) + $signed(buffer_3_609); // @[Modules.scala 56:109:@14616.4]
  assign _T_66630 = _T_66629[10:0]; // @[Modules.scala 56:109:@14617.4]
  assign buffer_3_696 = $signed(_T_66630); // @[Modules.scala 56:109:@14618.4]
  assign _T_66632 = $signed(buffer_3_610) + $signed(buffer_3_611); // @[Modules.scala 56:109:@14620.4]
  assign _T_66633 = _T_66632[10:0]; // @[Modules.scala 56:109:@14621.4]
  assign buffer_3_697 = $signed(_T_66633); // @[Modules.scala 56:109:@14622.4]
  assign _T_66635 = $signed(buffer_3_612) + $signed(buffer_3_613); // @[Modules.scala 56:109:@14624.4]
  assign _T_66636 = _T_66635[10:0]; // @[Modules.scala 56:109:@14625.4]
  assign buffer_3_698 = $signed(_T_66636); // @[Modules.scala 56:109:@14626.4]
  assign _T_66638 = $signed(buffer_3_614) + $signed(buffer_3_615); // @[Modules.scala 56:109:@14628.4]
  assign _T_66639 = _T_66638[10:0]; // @[Modules.scala 56:109:@14629.4]
  assign buffer_3_699 = $signed(_T_66639); // @[Modules.scala 56:109:@14630.4]
  assign _T_66641 = $signed(buffer_3_616) + $signed(buffer_3_617); // @[Modules.scala 56:109:@14632.4]
  assign _T_66642 = _T_66641[10:0]; // @[Modules.scala 56:109:@14633.4]
  assign buffer_3_700 = $signed(_T_66642); // @[Modules.scala 56:109:@14634.4]
  assign _T_66644 = $signed(buffer_3_618) + $signed(buffer_3_619); // @[Modules.scala 56:109:@14636.4]
  assign _T_66645 = _T_66644[10:0]; // @[Modules.scala 56:109:@14637.4]
  assign buffer_3_701 = $signed(_T_66645); // @[Modules.scala 56:109:@14638.4]
  assign _T_66647 = $signed(buffer_3_620) + $signed(buffer_3_621); // @[Modules.scala 56:109:@14640.4]
  assign _T_66648 = _T_66647[10:0]; // @[Modules.scala 56:109:@14641.4]
  assign buffer_3_702 = $signed(_T_66648); // @[Modules.scala 56:109:@14642.4]
  assign _T_66650 = $signed(buffer_3_622) + $signed(buffer_3_623); // @[Modules.scala 56:109:@14644.4]
  assign _T_66651 = _T_66650[10:0]; // @[Modules.scala 56:109:@14645.4]
  assign buffer_3_703 = $signed(_T_66651); // @[Modules.scala 56:109:@14646.4]
  assign _T_66653 = $signed(buffer_3_624) + $signed(buffer_3_625); // @[Modules.scala 56:109:@14648.4]
  assign _T_66654 = _T_66653[10:0]; // @[Modules.scala 56:109:@14649.4]
  assign buffer_3_704 = $signed(_T_66654); // @[Modules.scala 56:109:@14650.4]
  assign _T_66656 = $signed(buffer_3_626) + $signed(buffer_3_627); // @[Modules.scala 56:109:@14652.4]
  assign _T_66657 = _T_66656[10:0]; // @[Modules.scala 56:109:@14653.4]
  assign buffer_3_705 = $signed(_T_66657); // @[Modules.scala 56:109:@14654.4]
  assign _T_66659 = $signed(buffer_3_628) + $signed(buffer_3_629); // @[Modules.scala 56:109:@14656.4]
  assign _T_66660 = _T_66659[10:0]; // @[Modules.scala 56:109:@14657.4]
  assign buffer_3_706 = $signed(_T_66660); // @[Modules.scala 56:109:@14658.4]
  assign _T_66662 = $signed(buffer_3_630) + $signed(buffer_3_631); // @[Modules.scala 56:109:@14660.4]
  assign _T_66663 = _T_66662[10:0]; // @[Modules.scala 56:109:@14661.4]
  assign buffer_3_707 = $signed(_T_66663); // @[Modules.scala 56:109:@14662.4]
  assign _T_66665 = $signed(buffer_2_632) + $signed(buffer_3_633); // @[Modules.scala 56:109:@14664.4]
  assign _T_66666 = _T_66665[10:0]; // @[Modules.scala 56:109:@14665.4]
  assign buffer_3_708 = $signed(_T_66666); // @[Modules.scala 56:109:@14666.4]
  assign _T_66668 = $signed(buffer_3_634) + $signed(buffer_3_635); // @[Modules.scala 56:109:@14668.4]
  assign _T_66669 = _T_66668[10:0]; // @[Modules.scala 56:109:@14669.4]
  assign buffer_3_709 = $signed(_T_66669); // @[Modules.scala 56:109:@14670.4]
  assign _T_66671 = $signed(buffer_3_636) + $signed(buffer_3_637); // @[Modules.scala 56:109:@14672.4]
  assign _T_66672 = _T_66671[10:0]; // @[Modules.scala 56:109:@14673.4]
  assign buffer_3_710 = $signed(_T_66672); // @[Modules.scala 56:109:@14674.4]
  assign _T_66674 = $signed(buffer_3_638) + $signed(buffer_3_639); // @[Modules.scala 56:109:@14676.4]
  assign _T_66675 = _T_66674[10:0]; // @[Modules.scala 56:109:@14677.4]
  assign buffer_3_711 = $signed(_T_66675); // @[Modules.scala 56:109:@14678.4]
  assign _T_66677 = $signed(buffer_3_640) + $signed(buffer_3_641); // @[Modules.scala 56:109:@14680.4]
  assign _T_66678 = _T_66677[10:0]; // @[Modules.scala 56:109:@14681.4]
  assign buffer_3_712 = $signed(_T_66678); // @[Modules.scala 56:109:@14682.4]
  assign _T_66680 = $signed(buffer_3_642) + $signed(buffer_3_643); // @[Modules.scala 56:109:@14684.4]
  assign _T_66681 = _T_66680[10:0]; // @[Modules.scala 56:109:@14685.4]
  assign buffer_3_713 = $signed(_T_66681); // @[Modules.scala 56:109:@14686.4]
  assign _T_66683 = $signed(buffer_3_644) + $signed(buffer_3_645); // @[Modules.scala 56:109:@14688.4]
  assign _T_66684 = _T_66683[10:0]; // @[Modules.scala 56:109:@14689.4]
  assign buffer_3_714 = $signed(_T_66684); // @[Modules.scala 56:109:@14690.4]
  assign _T_66686 = $signed(buffer_3_646) + $signed(buffer_3_647); // @[Modules.scala 56:109:@14692.4]
  assign _T_66687 = _T_66686[10:0]; // @[Modules.scala 56:109:@14693.4]
  assign buffer_3_715 = $signed(_T_66687); // @[Modules.scala 56:109:@14694.4]
  assign _T_66689 = $signed(buffer_3_648) + $signed(buffer_3_649); // @[Modules.scala 56:109:@14696.4]
  assign _T_66690 = _T_66689[10:0]; // @[Modules.scala 56:109:@14697.4]
  assign buffer_3_716 = $signed(_T_66690); // @[Modules.scala 56:109:@14698.4]
  assign _T_66692 = $signed(buffer_3_650) + $signed(buffer_3_651); // @[Modules.scala 56:109:@14700.4]
  assign _T_66693 = _T_66692[10:0]; // @[Modules.scala 56:109:@14701.4]
  assign buffer_3_717 = $signed(_T_66693); // @[Modules.scala 56:109:@14702.4]
  assign _T_66695 = $signed(buffer_3_652) + $signed(buffer_3_653); // @[Modules.scala 56:109:@14704.4]
  assign _T_66696 = _T_66695[10:0]; // @[Modules.scala 56:109:@14705.4]
  assign buffer_3_718 = $signed(_T_66696); // @[Modules.scala 56:109:@14706.4]
  assign _T_66698 = $signed(buffer_3_654) + $signed(buffer_3_655); // @[Modules.scala 56:109:@14708.4]
  assign _T_66699 = _T_66698[10:0]; // @[Modules.scala 56:109:@14709.4]
  assign buffer_3_719 = $signed(_T_66699); // @[Modules.scala 56:109:@14710.4]
  assign _T_66701 = $signed(buffer_3_656) + $signed(buffer_3_657); // @[Modules.scala 56:109:@14712.4]
  assign _T_66702 = _T_66701[10:0]; // @[Modules.scala 56:109:@14713.4]
  assign buffer_3_720 = $signed(_T_66702); // @[Modules.scala 56:109:@14714.4]
  assign _T_66704 = $signed(buffer_3_658) + $signed(buffer_3_659); // @[Modules.scala 56:109:@14716.4]
  assign _T_66705 = _T_66704[10:0]; // @[Modules.scala 56:109:@14717.4]
  assign buffer_3_721 = $signed(_T_66705); // @[Modules.scala 56:109:@14718.4]
  assign _T_66707 = $signed(buffer_3_660) + $signed(buffer_3_661); // @[Modules.scala 56:109:@14720.4]
  assign _T_66708 = _T_66707[10:0]; // @[Modules.scala 56:109:@14721.4]
  assign buffer_3_722 = $signed(_T_66708); // @[Modules.scala 56:109:@14722.4]
  assign _T_66710 = $signed(buffer_3_662) + $signed(buffer_3_663); // @[Modules.scala 56:109:@14724.4]
  assign _T_66711 = _T_66710[10:0]; // @[Modules.scala 56:109:@14725.4]
  assign buffer_3_723 = $signed(_T_66711); // @[Modules.scala 56:109:@14726.4]
  assign _T_66713 = $signed(buffer_3_664) + $signed(buffer_3_665); // @[Modules.scala 56:109:@14728.4]
  assign _T_66714 = _T_66713[10:0]; // @[Modules.scala 56:109:@14729.4]
  assign buffer_3_724 = $signed(_T_66714); // @[Modules.scala 56:109:@14730.4]
  assign _T_66716 = $signed(buffer_3_666) + $signed(buffer_3_667); // @[Modules.scala 56:109:@14732.4]
  assign _T_66717 = _T_66716[10:0]; // @[Modules.scala 56:109:@14733.4]
  assign buffer_3_725 = $signed(_T_66717); // @[Modules.scala 56:109:@14734.4]
  assign _T_66719 = $signed(buffer_3_668) + $signed(buffer_3_669); // @[Modules.scala 56:109:@14736.4]
  assign _T_66720 = _T_66719[10:0]; // @[Modules.scala 56:109:@14737.4]
  assign buffer_3_726 = $signed(_T_66720); // @[Modules.scala 56:109:@14738.4]
  assign _T_66722 = $signed(buffer_3_670) + $signed(buffer_3_671); // @[Modules.scala 56:109:@14740.4]
  assign _T_66723 = _T_66722[10:0]; // @[Modules.scala 56:109:@14741.4]
  assign buffer_3_727 = $signed(_T_66723); // @[Modules.scala 56:109:@14742.4]
  assign _T_66725 = $signed(buffer_3_672) + $signed(buffer_3_673); // @[Modules.scala 56:109:@14744.4]
  assign _T_66726 = _T_66725[10:0]; // @[Modules.scala 56:109:@14745.4]
  assign buffer_3_728 = $signed(_T_66726); // @[Modules.scala 56:109:@14746.4]
  assign _T_66728 = $signed(buffer_3_674) + $signed(buffer_3_675); // @[Modules.scala 56:109:@14748.4]
  assign _T_66729 = _T_66728[10:0]; // @[Modules.scala 56:109:@14749.4]
  assign buffer_3_729 = $signed(_T_66729); // @[Modules.scala 56:109:@14750.4]
  assign _T_66731 = $signed(buffer_3_676) + $signed(buffer_3_677); // @[Modules.scala 56:109:@14752.4]
  assign _T_66732 = _T_66731[10:0]; // @[Modules.scala 56:109:@14753.4]
  assign buffer_3_730 = $signed(_T_66732); // @[Modules.scala 56:109:@14754.4]
  assign _T_66734 = $signed(buffer_3_678) + $signed(buffer_3_679); // @[Modules.scala 56:109:@14756.4]
  assign _T_66735 = _T_66734[10:0]; // @[Modules.scala 56:109:@14757.4]
  assign buffer_3_731 = $signed(_T_66735); // @[Modules.scala 56:109:@14758.4]
  assign _T_66737 = $signed(buffer_3_680) + $signed(buffer_3_681); // @[Modules.scala 56:109:@14760.4]
  assign _T_66738 = _T_66737[10:0]; // @[Modules.scala 56:109:@14761.4]
  assign buffer_3_732 = $signed(_T_66738); // @[Modules.scala 56:109:@14762.4]
  assign _T_66740 = $signed(buffer_3_682) + $signed(buffer_3_683); // @[Modules.scala 56:109:@14764.4]
  assign _T_66741 = _T_66740[10:0]; // @[Modules.scala 56:109:@14765.4]
  assign buffer_3_733 = $signed(_T_66741); // @[Modules.scala 56:109:@14766.4]
  assign _T_66743 = $signed(buffer_3_684) + $signed(buffer_3_685); // @[Modules.scala 56:109:@14768.4]
  assign _T_66744 = _T_66743[10:0]; // @[Modules.scala 56:109:@14769.4]
  assign buffer_3_734 = $signed(_T_66744); // @[Modules.scala 56:109:@14770.4]
  assign _T_66746 = $signed(buffer_3_686) + $signed(buffer_3_687); // @[Modules.scala 63:156:@14773.4]
  assign _T_66747 = _T_66746[10:0]; // @[Modules.scala 63:156:@14774.4]
  assign buffer_3_736 = $signed(_T_66747); // @[Modules.scala 63:156:@14775.4]
  assign _T_66749 = $signed(buffer_3_736) + $signed(buffer_3_688); // @[Modules.scala 63:156:@14777.4]
  assign _T_66750 = _T_66749[10:0]; // @[Modules.scala 63:156:@14778.4]
  assign buffer_3_737 = $signed(_T_66750); // @[Modules.scala 63:156:@14779.4]
  assign _T_66752 = $signed(buffer_3_737) + $signed(buffer_3_689); // @[Modules.scala 63:156:@14781.4]
  assign _T_66753 = _T_66752[10:0]; // @[Modules.scala 63:156:@14782.4]
  assign buffer_3_738 = $signed(_T_66753); // @[Modules.scala 63:156:@14783.4]
  assign _T_66755 = $signed(buffer_3_738) + $signed(buffer_3_690); // @[Modules.scala 63:156:@14785.4]
  assign _T_66756 = _T_66755[10:0]; // @[Modules.scala 63:156:@14786.4]
  assign buffer_3_739 = $signed(_T_66756); // @[Modules.scala 63:156:@14787.4]
  assign _T_66758 = $signed(buffer_3_739) + $signed(buffer_3_691); // @[Modules.scala 63:156:@14789.4]
  assign _T_66759 = _T_66758[10:0]; // @[Modules.scala 63:156:@14790.4]
  assign buffer_3_740 = $signed(_T_66759); // @[Modules.scala 63:156:@14791.4]
  assign _T_66761 = $signed(buffer_3_740) + $signed(buffer_3_692); // @[Modules.scala 63:156:@14793.4]
  assign _T_66762 = _T_66761[10:0]; // @[Modules.scala 63:156:@14794.4]
  assign buffer_3_741 = $signed(_T_66762); // @[Modules.scala 63:156:@14795.4]
  assign _T_66764 = $signed(buffer_3_741) + $signed(buffer_3_693); // @[Modules.scala 63:156:@14797.4]
  assign _T_66765 = _T_66764[10:0]; // @[Modules.scala 63:156:@14798.4]
  assign buffer_3_742 = $signed(_T_66765); // @[Modules.scala 63:156:@14799.4]
  assign _T_66767 = $signed(buffer_3_742) + $signed(buffer_3_694); // @[Modules.scala 63:156:@14801.4]
  assign _T_66768 = _T_66767[10:0]; // @[Modules.scala 63:156:@14802.4]
  assign buffer_3_743 = $signed(_T_66768); // @[Modules.scala 63:156:@14803.4]
  assign _T_66770 = $signed(buffer_3_743) + $signed(buffer_3_695); // @[Modules.scala 63:156:@14805.4]
  assign _T_66771 = _T_66770[10:0]; // @[Modules.scala 63:156:@14806.4]
  assign buffer_3_744 = $signed(_T_66771); // @[Modules.scala 63:156:@14807.4]
  assign _T_66773 = $signed(buffer_3_744) + $signed(buffer_3_696); // @[Modules.scala 63:156:@14809.4]
  assign _T_66774 = _T_66773[10:0]; // @[Modules.scala 63:156:@14810.4]
  assign buffer_3_745 = $signed(_T_66774); // @[Modules.scala 63:156:@14811.4]
  assign _T_66776 = $signed(buffer_3_745) + $signed(buffer_3_697); // @[Modules.scala 63:156:@14813.4]
  assign _T_66777 = _T_66776[10:0]; // @[Modules.scala 63:156:@14814.4]
  assign buffer_3_746 = $signed(_T_66777); // @[Modules.scala 63:156:@14815.4]
  assign _T_66779 = $signed(buffer_3_746) + $signed(buffer_3_698); // @[Modules.scala 63:156:@14817.4]
  assign _T_66780 = _T_66779[10:0]; // @[Modules.scala 63:156:@14818.4]
  assign buffer_3_747 = $signed(_T_66780); // @[Modules.scala 63:156:@14819.4]
  assign _T_66782 = $signed(buffer_3_747) + $signed(buffer_3_699); // @[Modules.scala 63:156:@14821.4]
  assign _T_66783 = _T_66782[10:0]; // @[Modules.scala 63:156:@14822.4]
  assign buffer_3_748 = $signed(_T_66783); // @[Modules.scala 63:156:@14823.4]
  assign _T_66785 = $signed(buffer_3_748) + $signed(buffer_3_700); // @[Modules.scala 63:156:@14825.4]
  assign _T_66786 = _T_66785[10:0]; // @[Modules.scala 63:156:@14826.4]
  assign buffer_3_749 = $signed(_T_66786); // @[Modules.scala 63:156:@14827.4]
  assign _T_66788 = $signed(buffer_3_749) + $signed(buffer_3_701); // @[Modules.scala 63:156:@14829.4]
  assign _T_66789 = _T_66788[10:0]; // @[Modules.scala 63:156:@14830.4]
  assign buffer_3_750 = $signed(_T_66789); // @[Modules.scala 63:156:@14831.4]
  assign _T_66791 = $signed(buffer_3_750) + $signed(buffer_3_702); // @[Modules.scala 63:156:@14833.4]
  assign _T_66792 = _T_66791[10:0]; // @[Modules.scala 63:156:@14834.4]
  assign buffer_3_751 = $signed(_T_66792); // @[Modules.scala 63:156:@14835.4]
  assign _T_66794 = $signed(buffer_3_751) + $signed(buffer_3_703); // @[Modules.scala 63:156:@14837.4]
  assign _T_66795 = _T_66794[10:0]; // @[Modules.scala 63:156:@14838.4]
  assign buffer_3_752 = $signed(_T_66795); // @[Modules.scala 63:156:@14839.4]
  assign _T_66797 = $signed(buffer_3_752) + $signed(buffer_3_704); // @[Modules.scala 63:156:@14841.4]
  assign _T_66798 = _T_66797[10:0]; // @[Modules.scala 63:156:@14842.4]
  assign buffer_3_753 = $signed(_T_66798); // @[Modules.scala 63:156:@14843.4]
  assign _T_66800 = $signed(buffer_3_753) + $signed(buffer_3_705); // @[Modules.scala 63:156:@14845.4]
  assign _T_66801 = _T_66800[10:0]; // @[Modules.scala 63:156:@14846.4]
  assign buffer_3_754 = $signed(_T_66801); // @[Modules.scala 63:156:@14847.4]
  assign _T_66803 = $signed(buffer_3_754) + $signed(buffer_3_706); // @[Modules.scala 63:156:@14849.4]
  assign _T_66804 = _T_66803[10:0]; // @[Modules.scala 63:156:@14850.4]
  assign buffer_3_755 = $signed(_T_66804); // @[Modules.scala 63:156:@14851.4]
  assign _T_66806 = $signed(buffer_3_755) + $signed(buffer_3_707); // @[Modules.scala 63:156:@14853.4]
  assign _T_66807 = _T_66806[10:0]; // @[Modules.scala 63:156:@14854.4]
  assign buffer_3_756 = $signed(_T_66807); // @[Modules.scala 63:156:@14855.4]
  assign _T_66809 = $signed(buffer_3_756) + $signed(buffer_3_708); // @[Modules.scala 63:156:@14857.4]
  assign _T_66810 = _T_66809[10:0]; // @[Modules.scala 63:156:@14858.4]
  assign buffer_3_757 = $signed(_T_66810); // @[Modules.scala 63:156:@14859.4]
  assign _T_66812 = $signed(buffer_3_757) + $signed(buffer_3_709); // @[Modules.scala 63:156:@14861.4]
  assign _T_66813 = _T_66812[10:0]; // @[Modules.scala 63:156:@14862.4]
  assign buffer_3_758 = $signed(_T_66813); // @[Modules.scala 63:156:@14863.4]
  assign _T_66815 = $signed(buffer_3_758) + $signed(buffer_3_710); // @[Modules.scala 63:156:@14865.4]
  assign _T_66816 = _T_66815[10:0]; // @[Modules.scala 63:156:@14866.4]
  assign buffer_3_759 = $signed(_T_66816); // @[Modules.scala 63:156:@14867.4]
  assign _T_66818 = $signed(buffer_3_759) + $signed(buffer_3_711); // @[Modules.scala 63:156:@14869.4]
  assign _T_66819 = _T_66818[10:0]; // @[Modules.scala 63:156:@14870.4]
  assign buffer_3_760 = $signed(_T_66819); // @[Modules.scala 63:156:@14871.4]
  assign _T_66821 = $signed(buffer_3_760) + $signed(buffer_3_712); // @[Modules.scala 63:156:@14873.4]
  assign _T_66822 = _T_66821[10:0]; // @[Modules.scala 63:156:@14874.4]
  assign buffer_3_761 = $signed(_T_66822); // @[Modules.scala 63:156:@14875.4]
  assign _T_66824 = $signed(buffer_3_761) + $signed(buffer_3_713); // @[Modules.scala 63:156:@14877.4]
  assign _T_66825 = _T_66824[10:0]; // @[Modules.scala 63:156:@14878.4]
  assign buffer_3_762 = $signed(_T_66825); // @[Modules.scala 63:156:@14879.4]
  assign _T_66827 = $signed(buffer_3_762) + $signed(buffer_3_714); // @[Modules.scala 63:156:@14881.4]
  assign _T_66828 = _T_66827[10:0]; // @[Modules.scala 63:156:@14882.4]
  assign buffer_3_763 = $signed(_T_66828); // @[Modules.scala 63:156:@14883.4]
  assign _T_66830 = $signed(buffer_3_763) + $signed(buffer_3_715); // @[Modules.scala 63:156:@14885.4]
  assign _T_66831 = _T_66830[10:0]; // @[Modules.scala 63:156:@14886.4]
  assign buffer_3_764 = $signed(_T_66831); // @[Modules.scala 63:156:@14887.4]
  assign _T_66833 = $signed(buffer_3_764) + $signed(buffer_3_716); // @[Modules.scala 63:156:@14889.4]
  assign _T_66834 = _T_66833[10:0]; // @[Modules.scala 63:156:@14890.4]
  assign buffer_3_765 = $signed(_T_66834); // @[Modules.scala 63:156:@14891.4]
  assign _T_66836 = $signed(buffer_3_765) + $signed(buffer_3_717); // @[Modules.scala 63:156:@14893.4]
  assign _T_66837 = _T_66836[10:0]; // @[Modules.scala 63:156:@14894.4]
  assign buffer_3_766 = $signed(_T_66837); // @[Modules.scala 63:156:@14895.4]
  assign _T_66839 = $signed(buffer_3_766) + $signed(buffer_3_718); // @[Modules.scala 63:156:@14897.4]
  assign _T_66840 = _T_66839[10:0]; // @[Modules.scala 63:156:@14898.4]
  assign buffer_3_767 = $signed(_T_66840); // @[Modules.scala 63:156:@14899.4]
  assign _T_66842 = $signed(buffer_3_767) + $signed(buffer_3_719); // @[Modules.scala 63:156:@14901.4]
  assign _T_66843 = _T_66842[10:0]; // @[Modules.scala 63:156:@14902.4]
  assign buffer_3_768 = $signed(_T_66843); // @[Modules.scala 63:156:@14903.4]
  assign _T_66845 = $signed(buffer_3_768) + $signed(buffer_3_720); // @[Modules.scala 63:156:@14905.4]
  assign _T_66846 = _T_66845[10:0]; // @[Modules.scala 63:156:@14906.4]
  assign buffer_3_769 = $signed(_T_66846); // @[Modules.scala 63:156:@14907.4]
  assign _T_66848 = $signed(buffer_3_769) + $signed(buffer_3_721); // @[Modules.scala 63:156:@14909.4]
  assign _T_66849 = _T_66848[10:0]; // @[Modules.scala 63:156:@14910.4]
  assign buffer_3_770 = $signed(_T_66849); // @[Modules.scala 63:156:@14911.4]
  assign _T_66851 = $signed(buffer_3_770) + $signed(buffer_3_722); // @[Modules.scala 63:156:@14913.4]
  assign _T_66852 = _T_66851[10:0]; // @[Modules.scala 63:156:@14914.4]
  assign buffer_3_771 = $signed(_T_66852); // @[Modules.scala 63:156:@14915.4]
  assign _T_66854 = $signed(buffer_3_771) + $signed(buffer_3_723); // @[Modules.scala 63:156:@14917.4]
  assign _T_66855 = _T_66854[10:0]; // @[Modules.scala 63:156:@14918.4]
  assign buffer_3_772 = $signed(_T_66855); // @[Modules.scala 63:156:@14919.4]
  assign _T_66857 = $signed(buffer_3_772) + $signed(buffer_3_724); // @[Modules.scala 63:156:@14921.4]
  assign _T_66858 = _T_66857[10:0]; // @[Modules.scala 63:156:@14922.4]
  assign buffer_3_773 = $signed(_T_66858); // @[Modules.scala 63:156:@14923.4]
  assign _T_66860 = $signed(buffer_3_773) + $signed(buffer_3_725); // @[Modules.scala 63:156:@14925.4]
  assign _T_66861 = _T_66860[10:0]; // @[Modules.scala 63:156:@14926.4]
  assign buffer_3_774 = $signed(_T_66861); // @[Modules.scala 63:156:@14927.4]
  assign _T_66863 = $signed(buffer_3_774) + $signed(buffer_3_726); // @[Modules.scala 63:156:@14929.4]
  assign _T_66864 = _T_66863[10:0]; // @[Modules.scala 63:156:@14930.4]
  assign buffer_3_775 = $signed(_T_66864); // @[Modules.scala 63:156:@14931.4]
  assign _T_66866 = $signed(buffer_3_775) + $signed(buffer_3_727); // @[Modules.scala 63:156:@14933.4]
  assign _T_66867 = _T_66866[10:0]; // @[Modules.scala 63:156:@14934.4]
  assign buffer_3_776 = $signed(_T_66867); // @[Modules.scala 63:156:@14935.4]
  assign _T_66869 = $signed(buffer_3_776) + $signed(buffer_3_728); // @[Modules.scala 63:156:@14937.4]
  assign _T_66870 = _T_66869[10:0]; // @[Modules.scala 63:156:@14938.4]
  assign buffer_3_777 = $signed(_T_66870); // @[Modules.scala 63:156:@14939.4]
  assign _T_66872 = $signed(buffer_3_777) + $signed(buffer_3_729); // @[Modules.scala 63:156:@14941.4]
  assign _T_66873 = _T_66872[10:0]; // @[Modules.scala 63:156:@14942.4]
  assign buffer_3_778 = $signed(_T_66873); // @[Modules.scala 63:156:@14943.4]
  assign _T_66875 = $signed(buffer_3_778) + $signed(buffer_3_730); // @[Modules.scala 63:156:@14945.4]
  assign _T_66876 = _T_66875[10:0]; // @[Modules.scala 63:156:@14946.4]
  assign buffer_3_779 = $signed(_T_66876); // @[Modules.scala 63:156:@14947.4]
  assign _T_66878 = $signed(buffer_3_779) + $signed(buffer_3_731); // @[Modules.scala 63:156:@14949.4]
  assign _T_66879 = _T_66878[10:0]; // @[Modules.scala 63:156:@14950.4]
  assign buffer_3_780 = $signed(_T_66879); // @[Modules.scala 63:156:@14951.4]
  assign _T_66881 = $signed(buffer_3_780) + $signed(buffer_3_732); // @[Modules.scala 63:156:@14953.4]
  assign _T_66882 = _T_66881[10:0]; // @[Modules.scala 63:156:@14954.4]
  assign buffer_3_781 = $signed(_T_66882); // @[Modules.scala 63:156:@14955.4]
  assign _T_66884 = $signed(buffer_3_781) + $signed(buffer_3_733); // @[Modules.scala 63:156:@14957.4]
  assign _T_66885 = _T_66884[10:0]; // @[Modules.scala 63:156:@14958.4]
  assign buffer_3_782 = $signed(_T_66885); // @[Modules.scala 63:156:@14959.4]
  assign _T_66887 = $signed(buffer_3_782) + $signed(buffer_3_734); // @[Modules.scala 63:156:@14961.4]
  assign _T_66888 = _T_66887[10:0]; // @[Modules.scala 63:156:@14962.4]
  assign buffer_3_783 = $signed(_T_66888); // @[Modules.scala 63:156:@14963.4]
  assign _T_66897 = $signed(_T_54276) + $signed(io_in_3); // @[Modules.scala 43:47:@14973.4]
  assign _T_66898 = _T_66897[4:0]; // @[Modules.scala 43:47:@14974.4]
  assign _T_66899 = $signed(_T_66898); // @[Modules.scala 43:47:@14975.4]
  assign _T_66921 = $signed(_T_54304) + $signed(io_in_11); // @[Modules.scala 43:47:@14998.4]
  assign _T_66922 = _T_66921[4:0]; // @[Modules.scala 43:47:@14999.4]
  assign _T_66923 = $signed(_T_66922); // @[Modules.scala 43:47:@15000.4]
  assign _T_66935 = $signed(5'sh0) - $signed(io_in_16); // @[Modules.scala 46:37:@15013.4]
  assign _T_66936 = _T_66935[4:0]; // @[Modules.scala 46:37:@15014.4]
  assign _T_66937 = $signed(_T_66936); // @[Modules.scala 46:37:@15015.4]
  assign _T_66938 = $signed(_T_66937) - $signed(io_in_17); // @[Modules.scala 46:47:@15016.4]
  assign _T_66939 = _T_66938[4:0]; // @[Modules.scala 46:47:@15017.4]
  assign _T_66940 = $signed(_T_66939); // @[Modules.scala 46:47:@15018.4]
  assign _T_66951 = $signed(_T_54338) - $signed(io_in_23); // @[Modules.scala 46:47:@15031.4]
  assign _T_66952 = _T_66951[4:0]; // @[Modules.scala 46:47:@15032.4]
  assign _T_66953 = $signed(_T_66952); // @[Modules.scala 46:47:@15033.4]
  assign _T_66961 = $signed(_T_57601) + $signed(io_in_27); // @[Modules.scala 43:47:@15042.4]
  assign _T_66962 = _T_66961[4:0]; // @[Modules.scala 43:47:@15043.4]
  assign _T_66963 = $signed(_T_66962); // @[Modules.scala 43:47:@15044.4]
  assign _T_66968 = $signed(_T_54355) + $signed(io_in_29); // @[Modules.scala 43:47:@15049.4]
  assign _T_66969 = _T_66968[4:0]; // @[Modules.scala 43:47:@15050.4]
  assign _T_66970 = $signed(_T_66969); // @[Modules.scala 43:47:@15051.4]
  assign _T_67000 = $signed(io_in_44) + $signed(io_in_45); // @[Modules.scala 37:46:@15087.4]
  assign _T_67001 = _T_67000[4:0]; // @[Modules.scala 37:46:@15088.4]
  assign _T_67002 = $signed(_T_67001); // @[Modules.scala 37:46:@15089.4]
  assign _T_67102 = $signed(_T_64136) + $signed(io_in_89); // @[Modules.scala 43:47:@15202.4]
  assign _T_67103 = _T_67102[4:0]; // @[Modules.scala 43:47:@15203.4]
  assign _T_67104 = $signed(_T_67103); // @[Modules.scala 43:47:@15204.4]
  assign _T_67156 = $signed(_T_60905) + $signed(io_in_117); // @[Modules.scala 43:47:@15267.4]
  assign _T_67157 = _T_67156[4:0]; // @[Modules.scala 43:47:@15268.4]
  assign _T_67158 = $signed(_T_67157); // @[Modules.scala 43:47:@15269.4]
  assign _T_67163 = $signed(_T_57775) + $signed(io_in_119); // @[Modules.scala 43:47:@15274.4]
  assign _T_67164 = _T_67163[4:0]; // @[Modules.scala 43:47:@15275.4]
  assign _T_67165 = $signed(_T_67164); // @[Modules.scala 43:47:@15276.4]
  assign _T_67169 = $signed(io_in_122) - $signed(io_in_123); // @[Modules.scala 40:46:@15282.4]
  assign _T_67170 = _T_67169[4:0]; // @[Modules.scala 40:46:@15283.4]
  assign _T_67171 = $signed(_T_67170); // @[Modules.scala 40:46:@15284.4]
  assign _T_67182 = $signed(io_in_128) - $signed(io_in_129); // @[Modules.scala 40:46:@15297.4]
  assign _T_67183 = _T_67182[4:0]; // @[Modules.scala 40:46:@15298.4]
  assign _T_67184 = $signed(_T_67183); // @[Modules.scala 40:46:@15299.4]
  assign _T_67200 = $signed(5'sh0) - $signed(io_in_134); // @[Modules.scala 46:37:@15315.4]
  assign _T_67201 = _T_67200[4:0]; // @[Modules.scala 46:37:@15316.4]
  assign _T_67202 = $signed(_T_67201); // @[Modules.scala 46:37:@15317.4]
  assign _T_67203 = $signed(_T_67202) - $signed(io_in_135); // @[Modules.scala 46:47:@15318.4]
  assign _T_67204 = _T_67203[4:0]; // @[Modules.scala 46:47:@15319.4]
  assign _T_67205 = $signed(_T_67204); // @[Modules.scala 46:47:@15320.4]
  assign _T_67209 = $signed(io_in_138) + $signed(io_in_139); // @[Modules.scala 37:46:@15326.4]
  assign _T_67210 = _T_67209[4:0]; // @[Modules.scala 37:46:@15327.4]
  assign _T_67211 = $signed(_T_67210); // @[Modules.scala 37:46:@15328.4]
  assign _T_67226 = $signed(io_in_144) + $signed(io_in_145); // @[Modules.scala 37:46:@15344.4]
  assign _T_67227 = _T_67226[4:0]; // @[Modules.scala 37:46:@15345.4]
  assign _T_67228 = $signed(_T_67227); // @[Modules.scala 37:46:@15346.4]
  assign _T_67238 = $signed(io_in_152) + $signed(io_in_153); // @[Modules.scala 37:46:@15360.4]
  assign _T_67239 = _T_67238[4:0]; // @[Modules.scala 37:46:@15361.4]
  assign _T_67240 = $signed(_T_67239); // @[Modules.scala 37:46:@15362.4]
  assign _T_67244 = $signed(io_in_156) + $signed(io_in_157); // @[Modules.scala 37:46:@15368.4]
  assign _T_67245 = _T_67244[4:0]; // @[Modules.scala 37:46:@15369.4]
  assign _T_67246 = $signed(_T_67245); // @[Modules.scala 37:46:@15370.4]
  assign _T_67250 = $signed(io_in_160) - $signed(io_in_161); // @[Modules.scala 40:46:@15376.4]
  assign _T_67251 = _T_67250[4:0]; // @[Modules.scala 40:46:@15377.4]
  assign _T_67252 = $signed(_T_67251); // @[Modules.scala 40:46:@15378.4]
  assign _T_67266 = $signed(io_in_168) + $signed(io_in_169); // @[Modules.scala 37:46:@15395.4]
  assign _T_67267 = _T_67266[4:0]; // @[Modules.scala 37:46:@15396.4]
  assign _T_67268 = $signed(_T_67267); // @[Modules.scala 37:46:@15397.4]
  assign _T_67306 = $signed(_T_54781) + $signed(io_in_185); // @[Modules.scala 43:47:@15439.4]
  assign _T_67307 = _T_67306[4:0]; // @[Modules.scala 43:47:@15440.4]
  assign _T_67308 = $signed(_T_67307); // @[Modules.scala 43:47:@15441.4]
  assign _T_67312 = $signed(io_in_188) + $signed(io_in_189); // @[Modules.scala 37:46:@15447.4]
  assign _T_67313 = _T_67312[4:0]; // @[Modules.scala 37:46:@15448.4]
  assign _T_67314 = $signed(_T_67313); // @[Modules.scala 37:46:@15449.4]
  assign _T_67345 = $signed(_T_54828) + $signed(io_in_203); // @[Modules.scala 43:47:@15484.4]
  assign _T_67346 = _T_67345[4:0]; // @[Modules.scala 43:47:@15485.4]
  assign _T_67347 = $signed(_T_67346); // @[Modules.scala 43:47:@15486.4]
  assign _T_67348 = $signed(io_in_204) - $signed(io_in_205); // @[Modules.scala 40:46:@15488.4]
  assign _T_67349 = _T_67348[4:0]; // @[Modules.scala 40:46:@15489.4]
  assign _T_67350 = $signed(_T_67349); // @[Modules.scala 40:46:@15490.4]
  assign _T_67362 = $signed(5'sh0) - $signed(io_in_210); // @[Modules.scala 46:37:@15503.4]
  assign _T_67363 = _T_67362[4:0]; // @[Modules.scala 46:37:@15504.4]
  assign _T_67364 = $signed(_T_67363); // @[Modules.scala 46:37:@15505.4]
  assign _T_67365 = $signed(_T_67364) - $signed(io_in_211); // @[Modules.scala 46:47:@15506.4]
  assign _T_67366 = _T_67365[4:0]; // @[Modules.scala 46:47:@15507.4]
  assign _T_67367 = $signed(_T_67366); // @[Modules.scala 46:47:@15508.4]
  assign _T_67372 = $signed(_T_58016) - $signed(io_in_213); // @[Modules.scala 46:47:@15513.4]
  assign _T_67373 = _T_67372[4:0]; // @[Modules.scala 46:47:@15514.4]
  assign _T_67374 = $signed(_T_67373); // @[Modules.scala 46:47:@15515.4]
  assign _T_67412 = $signed(_T_54911) + $signed(io_in_229); // @[Modules.scala 43:47:@15557.4]
  assign _T_67413 = _T_67412[4:0]; // @[Modules.scala 43:47:@15558.4]
  assign _T_67414 = $signed(_T_67413); // @[Modules.scala 43:47:@15559.4]
  assign _T_67422 = $signed(io_in_232) + $signed(io_in_233); // @[Modules.scala 37:46:@15568.4]
  assign _T_67423 = _T_67422[4:0]; // @[Modules.scala 37:46:@15569.4]
  assign _T_67424 = $signed(_T_67423); // @[Modules.scala 37:46:@15570.4]
  assign _T_67453 = $signed(_T_54960) + $signed(io_in_243); // @[Modules.scala 43:47:@15600.4]
  assign _T_67454 = _T_67453[4:0]; // @[Modules.scala 43:47:@15601.4]
  assign _T_67455 = $signed(_T_67454); // @[Modules.scala 43:47:@15602.4]
  assign _T_67456 = $signed(io_in_244) + $signed(io_in_245); // @[Modules.scala 37:46:@15604.4]
  assign _T_67457 = _T_67456[4:0]; // @[Modules.scala 37:46:@15605.4]
  assign _T_67458 = $signed(_T_67457); // @[Modules.scala 37:46:@15606.4]
  assign _T_67486 = $signed(_T_55009) + $signed(io_in_257); // @[Modules.scala 43:47:@15637.4]
  assign _T_67487 = _T_67486[4:0]; // @[Modules.scala 43:47:@15638.4]
  assign _T_67488 = $signed(_T_67487); // @[Modules.scala 43:47:@15639.4]
  assign _T_67489 = $signed(io_in_258) + $signed(io_in_259); // @[Modules.scala 37:46:@15641.4]
  assign _T_67490 = _T_67489[4:0]; // @[Modules.scala 37:46:@15642.4]
  assign _T_67491 = $signed(_T_67490); // @[Modules.scala 37:46:@15643.4]
  assign _T_67492 = $signed(io_in_260) + $signed(io_in_261); // @[Modules.scala 37:46:@15645.4]
  assign _T_67493 = _T_67492[4:0]; // @[Modules.scala 37:46:@15646.4]
  assign _T_67494 = $signed(_T_67493); // @[Modules.scala 37:46:@15647.4]
  assign _T_67594 = $signed(_T_55145) + $signed(io_in_297); // @[Modules.scala 43:47:@15753.4]
  assign _T_67595 = _T_67594[4:0]; // @[Modules.scala 43:47:@15754.4]
  assign _T_67596 = $signed(_T_67595); // @[Modules.scala 43:47:@15755.4]
  assign _T_67597 = $signed(io_in_298) + $signed(io_in_299); // @[Modules.scala 37:46:@15757.4]
  assign _T_67598 = _T_67597[4:0]; // @[Modules.scala 37:46:@15758.4]
  assign _T_67599 = $signed(_T_67598); // @[Modules.scala 37:46:@15759.4]
  assign _T_67607 = $signed(io_in_302) + $signed(io_in_303); // @[Modules.scala 37:46:@15768.4]
  assign _T_67608 = _T_67607[4:0]; // @[Modules.scala 37:46:@15769.4]
  assign _T_67609 = $signed(_T_67608); // @[Modules.scala 37:46:@15770.4]
  assign _T_67616 = $signed(io_in_308) - $signed(io_in_309); // @[Modules.scala 40:46:@15780.4]
  assign _T_67617 = _T_67616[4:0]; // @[Modules.scala 40:46:@15781.4]
  assign _T_67618 = $signed(_T_67617); // @[Modules.scala 40:46:@15782.4]
  assign _T_67623 = $signed(_T_55194) + $signed(io_in_311); // @[Modules.scala 43:47:@15787.4]
  assign _T_67624 = _T_67623[4:0]; // @[Modules.scala 43:47:@15788.4]
  assign _T_67625 = $signed(_T_67624); // @[Modules.scala 43:47:@15789.4]
  assign _T_67718 = $signed(io_in_344) - $signed(io_in_345); // @[Modules.scala 40:46:@15888.4]
  assign _T_67719 = _T_67718[4:0]; // @[Modules.scala 40:46:@15889.4]
  assign _T_67720 = $signed(_T_67719); // @[Modules.scala 40:46:@15890.4]
  assign _T_67734 = $signed(io_in_352) - $signed(io_in_353); // @[Modules.scala 40:46:@15907.4]
  assign _T_67735 = _T_67734[4:0]; // @[Modules.scala 40:46:@15908.4]
  assign _T_67736 = $signed(_T_67735); // @[Modules.scala 40:46:@15909.4]
  assign _T_67764 = $signed(io_in_364) - $signed(io_in_365); // @[Modules.scala 40:46:@15940.4]
  assign _T_67765 = _T_67764[4:0]; // @[Modules.scala 40:46:@15941.4]
  assign _T_67766 = $signed(_T_67765); // @[Modules.scala 40:46:@15942.4]
  assign _T_67781 = $signed(io_in_370) - $signed(io_in_371); // @[Modules.scala 40:46:@15958.4]
  assign _T_67782 = _T_67781[4:0]; // @[Modules.scala 40:46:@15959.4]
  assign _T_67783 = $signed(_T_67782); // @[Modules.scala 40:46:@15960.4]
  assign _T_67800 = $signed(io_in_380) - $signed(io_in_381); // @[Modules.scala 40:46:@15981.4]
  assign _T_67801 = _T_67800[4:0]; // @[Modules.scala 40:46:@15982.4]
  assign _T_67802 = $signed(_T_67801); // @[Modules.scala 40:46:@15983.4]
  assign _T_67820 = $signed(io_in_388) + $signed(io_in_389); // @[Modules.scala 37:46:@16003.4]
  assign _T_67821 = _T_67820[4:0]; // @[Modules.scala 37:46:@16004.4]
  assign _T_67822 = $signed(_T_67821); // @[Modules.scala 37:46:@16005.4]
  assign _T_67823 = $signed(io_in_390) - $signed(io_in_391); // @[Modules.scala 40:46:@16007.4]
  assign _T_67824 = _T_67823[4:0]; // @[Modules.scala 40:46:@16008.4]
  assign _T_67825 = $signed(_T_67824); // @[Modules.scala 40:46:@16009.4]
  assign _T_67826 = $signed(io_in_392) - $signed(io_in_393); // @[Modules.scala 40:46:@16011.4]
  assign _T_67827 = _T_67826[4:0]; // @[Modules.scala 40:46:@16012.4]
  assign _T_67828 = $signed(_T_67827); // @[Modules.scala 40:46:@16013.4]
  assign _T_67847 = $signed(_T_64857) + $signed(io_in_399); // @[Modules.scala 43:47:@16032.4]
  assign _T_67848 = _T_67847[4:0]; // @[Modules.scala 43:47:@16033.4]
  assign _T_67849 = $signed(_T_67848); // @[Modules.scala 43:47:@16034.4]
  assign _T_67867 = $signed(_T_58551) + $signed(io_in_407); // @[Modules.scala 43:47:@16054.4]
  assign _T_67868 = _T_67867[4:0]; // @[Modules.scala 43:47:@16055.4]
  assign _T_67869 = $signed(_T_67868); // @[Modules.scala 43:47:@16056.4]
  assign _T_67876 = $signed(io_in_412) - $signed(io_in_413); // @[Modules.scala 40:46:@16066.4]
  assign _T_67877 = _T_67876[4:0]; // @[Modules.scala 40:46:@16067.4]
  assign _T_67878 = $signed(_T_67877); // @[Modules.scala 40:46:@16068.4]
  assign _T_67882 = $signed(io_in_416) + $signed(io_in_417); // @[Modules.scala 37:46:@16074.4]
  assign _T_67883 = _T_67882[4:0]; // @[Modules.scala 37:46:@16075.4]
  assign _T_67884 = $signed(_T_67883); // @[Modules.scala 37:46:@16076.4]
  assign _T_67885 = $signed(io_in_418) - $signed(io_in_419); // @[Modules.scala 40:46:@16078.4]
  assign _T_67886 = _T_67885[4:0]; // @[Modules.scala 40:46:@16079.4]
  assign _T_67887 = $signed(_T_67886); // @[Modules.scala 40:46:@16080.4]
  assign _T_67888 = $signed(io_in_420) + $signed(io_in_421); // @[Modules.scala 37:46:@16082.4]
  assign _T_67889 = _T_67888[4:0]; // @[Modules.scala 37:46:@16083.4]
  assign _T_67890 = $signed(_T_67889); // @[Modules.scala 37:46:@16084.4]
  assign _T_67910 = $signed(io_in_432) - $signed(io_in_433); // @[Modules.scala 40:46:@16109.4]
  assign _T_67911 = _T_67910[4:0]; // @[Modules.scala 40:46:@16110.4]
  assign _T_67912 = $signed(_T_67911); // @[Modules.scala 40:46:@16111.4]
  assign _T_67916 = $signed(io_in_436) - $signed(io_in_437); // @[Modules.scala 40:46:@16117.4]
  assign _T_67917 = _T_67916[4:0]; // @[Modules.scala 40:46:@16118.4]
  assign _T_67918 = $signed(_T_67917); // @[Modules.scala 40:46:@16119.4]
  assign _T_67959 = $signed(io_in_454) - $signed(io_in_455); // @[Modules.scala 40:46:@16165.4]
  assign _T_67960 = _T_67959[4:0]; // @[Modules.scala 40:46:@16166.4]
  assign _T_67961 = $signed(_T_67960); // @[Modules.scala 40:46:@16167.4]
  assign _T_67979 = $signed(_T_58699) + $signed(io_in_463); // @[Modules.scala 43:47:@16187.4]
  assign _T_67980 = _T_67979[4:0]; // @[Modules.scala 43:47:@16188.4]
  assign _T_67981 = $signed(_T_67980); // @[Modules.scala 43:47:@16189.4]
  assign _T_68027 = $signed(_T_58763) + $signed(io_in_487); // @[Modules.scala 43:47:@16244.4]
  assign _T_68028 = _T_68027[4:0]; // @[Modules.scala 43:47:@16245.4]
  assign _T_68029 = $signed(_T_68028); // @[Modules.scala 43:47:@16246.4]
  assign _T_68044 = $signed(io_in_492) + $signed(io_in_493); // @[Modules.scala 37:46:@16262.4]
  assign _T_68045 = _T_68044[4:0]; // @[Modules.scala 37:46:@16263.4]
  assign _T_68046 = $signed(_T_68045); // @[Modules.scala 37:46:@16264.4]
  assign _T_68048 = $signed(5'sh0) - $signed(io_in_494); // @[Modules.scala 43:37:@16266.4]
  assign _T_68049 = _T_68048[4:0]; // @[Modules.scala 43:37:@16267.4]
  assign _T_68050 = $signed(_T_68049); // @[Modules.scala 43:37:@16268.4]
  assign _T_68051 = $signed(_T_68050) + $signed(io_in_495); // @[Modules.scala 43:47:@16269.4]
  assign _T_68052 = _T_68051[4:0]; // @[Modules.scala 43:47:@16270.4]
  assign _T_68053 = $signed(_T_68052); // @[Modules.scala 43:47:@16271.4]
  assign _T_68082 = $signed(io_in_512) - $signed(io_in_513); // @[Modules.scala 40:46:@16308.4]
  assign _T_68083 = _T_68082[4:0]; // @[Modules.scala 40:46:@16309.4]
  assign _T_68084 = $signed(_T_68083); // @[Modules.scala 40:46:@16310.4]
  assign _T_68085 = $signed(io_in_514) - $signed(io_in_515); // @[Modules.scala 40:46:@16312.4]
  assign _T_68086 = _T_68085[4:0]; // @[Modules.scala 40:46:@16313.4]
  assign _T_68087 = $signed(_T_68086); // @[Modules.scala 40:46:@16314.4]
  assign _T_68095 = $signed(_T_58847) + $signed(io_in_519); // @[Modules.scala 43:47:@16323.4]
  assign _T_68096 = _T_68095[4:0]; // @[Modules.scala 43:47:@16324.4]
  assign _T_68097 = $signed(_T_68096); // @[Modules.scala 43:47:@16325.4]
  assign _T_68098 = $signed(io_in_520) - $signed(io_in_521); // @[Modules.scala 40:46:@16327.4]
  assign _T_68099 = _T_68098[4:0]; // @[Modules.scala 40:46:@16328.4]
  assign _T_68100 = $signed(_T_68099); // @[Modules.scala 40:46:@16329.4]
  assign _T_68146 = $signed(io_in_544) - $signed(io_in_545); // @[Modules.scala 40:46:@16384.4]
  assign _T_68147 = _T_68146[4:0]; // @[Modules.scala 40:46:@16385.4]
  assign _T_68148 = $signed(_T_68147); // @[Modules.scala 40:46:@16386.4]
  assign _T_68149 = $signed(io_in_546) + $signed(io_in_547); // @[Modules.scala 37:46:@16388.4]
  assign _T_68150 = _T_68149[4:0]; // @[Modules.scala 37:46:@16389.4]
  assign _T_68151 = $signed(_T_68150); // @[Modules.scala 37:46:@16390.4]
  assign _T_68212 = $signed(io_in_580) + $signed(io_in_581); // @[Modules.scala 37:46:@16465.4]
  assign _T_68213 = _T_68212[4:0]; // @[Modules.scala 37:46:@16466.4]
  assign _T_68214 = $signed(_T_68213); // @[Modules.scala 37:46:@16467.4]
  assign _T_68218 = $signed(io_in_584) - $signed(io_in_585); // @[Modules.scala 40:46:@16473.4]
  assign _T_68219 = _T_68218[4:0]; // @[Modules.scala 40:46:@16474.4]
  assign _T_68220 = $signed(_T_68219); // @[Modules.scala 40:46:@16475.4]
  assign _T_68225 = $signed(_T_55868) - $signed(io_in_587); // @[Modules.scala 46:47:@16480.4]
  assign _T_68226 = _T_68225[4:0]; // @[Modules.scala 46:47:@16481.4]
  assign _T_68227 = $signed(_T_68226); // @[Modules.scala 46:47:@16482.4]
  assign _T_68268 = $signed(io_in_612) - $signed(io_in_613); // @[Modules.scala 40:46:@16535.4]
  assign _T_68269 = _T_68268[4:0]; // @[Modules.scala 40:46:@16536.4]
  assign _T_68270 = $signed(_T_68269); // @[Modules.scala 40:46:@16537.4]
  assign _T_68271 = $signed(io_in_614) + $signed(io_in_615); // @[Modules.scala 37:46:@16539.4]
  assign _T_68272 = _T_68271[4:0]; // @[Modules.scala 37:46:@16540.4]
  assign _T_68273 = $signed(_T_68272); // @[Modules.scala 37:46:@16541.4]
  assign _T_68287 = $signed(io_in_622) + $signed(io_in_623); // @[Modules.scala 37:46:@16558.4]
  assign _T_68288 = _T_68287[4:0]; // @[Modules.scala 37:46:@16559.4]
  assign _T_68289 = $signed(_T_68288); // @[Modules.scala 37:46:@16560.4]
  assign _T_68310 = $signed(_T_56005) + $signed(io_in_633); // @[Modules.scala 43:47:@16584.4]
  assign _T_68311 = _T_68310[4:0]; // @[Modules.scala 43:47:@16585.4]
  assign _T_68312 = $signed(_T_68311); // @[Modules.scala 43:47:@16586.4]
  assign _T_68346 = $signed(io_in_648) - $signed(io_in_649); // @[Modules.scala 40:46:@16625.4]
  assign _T_68347 = _T_68346[4:0]; // @[Modules.scala 40:46:@16626.4]
  assign _T_68348 = $signed(_T_68347); // @[Modules.scala 40:46:@16627.4]
  assign _T_68368 = $signed(io_in_660) - $signed(io_in_661); // @[Modules.scala 40:46:@16652.4]
  assign _T_68369 = _T_68368[4:0]; // @[Modules.scala 40:46:@16653.4]
  assign _T_68370 = $signed(_T_68369); // @[Modules.scala 40:46:@16654.4]
  assign _T_68388 = $signed(_T_59156) + $signed(io_in_669); // @[Modules.scala 43:47:@16674.4]
  assign _T_68389 = _T_68388[4:0]; // @[Modules.scala 43:47:@16675.4]
  assign _T_68390 = $signed(_T_68389); // @[Modules.scala 43:47:@16676.4]
  assign _T_68395 = $signed(_T_56118) + $signed(io_in_671); // @[Modules.scala 43:47:@16681.4]
  assign _T_68396 = _T_68395[4:0]; // @[Modules.scala 43:47:@16682.4]
  assign _T_68397 = $signed(_T_68396); // @[Modules.scala 43:47:@16683.4]
  assign _T_68398 = $signed(io_in_672) + $signed(io_in_673); // @[Modules.scala 37:46:@16685.4]
  assign _T_68399 = _T_68398[4:0]; // @[Modules.scala 37:46:@16686.4]
  assign _T_68400 = $signed(_T_68399); // @[Modules.scala 37:46:@16687.4]
  assign _T_68404 = $signed(io_in_676) - $signed(io_in_677); // @[Modules.scala 40:46:@16693.4]
  assign _T_68405 = _T_68404[4:0]; // @[Modules.scala 40:46:@16694.4]
  assign _T_68406 = $signed(_T_68405); // @[Modules.scala 40:46:@16695.4]
  assign _T_68411 = $signed(_T_62436) + $signed(io_in_679); // @[Modules.scala 43:47:@16700.4]
  assign _T_68412 = _T_68411[4:0]; // @[Modules.scala 43:47:@16701.4]
  assign _T_68413 = $signed(_T_68412); // @[Modules.scala 43:47:@16702.4]
  assign _T_68454 = $signed(_T_62483) + $signed(io_in_697); // @[Modules.scala 43:47:@16748.4]
  assign _T_68455 = _T_68454[4:0]; // @[Modules.scala 43:47:@16749.4]
  assign _T_68456 = $signed(_T_68455); // @[Modules.scala 43:47:@16750.4]
  assign _T_68457 = $signed(io_in_698) - $signed(io_in_699); // @[Modules.scala 40:46:@16752.4]
  assign _T_68458 = _T_68457[4:0]; // @[Modules.scala 40:46:@16753.4]
  assign _T_68459 = $signed(_T_68458); // @[Modules.scala 40:46:@16754.4]
  assign _T_68466 = $signed(io_in_704) - $signed(io_in_705); // @[Modules.scala 40:46:@16764.4]
  assign _T_68467 = _T_68466[4:0]; // @[Modules.scala 40:46:@16765.4]
  assign _T_68468 = $signed(_T_68467); // @[Modules.scala 40:46:@16766.4]
  assign _T_68533 = $signed(5'sh0) - $signed(io_in_724); // @[Modules.scala 46:37:@16831.4]
  assign _T_68534 = _T_68533[4:0]; // @[Modules.scala 46:37:@16832.4]
  assign _T_68535 = $signed(_T_68534); // @[Modules.scala 46:37:@16833.4]
  assign _T_68536 = $signed(_T_68535) - $signed(io_in_725); // @[Modules.scala 46:47:@16834.4]
  assign _T_68537 = _T_68536[4:0]; // @[Modules.scala 46:47:@16835.4]
  assign _T_68538 = $signed(_T_68537); // @[Modules.scala 46:47:@16836.4]
  assign _T_68539 = $signed(io_in_726) + $signed(io_in_727); // @[Modules.scala 37:46:@16838.4]
  assign _T_68540 = _T_68539[4:0]; // @[Modules.scala 37:46:@16839.4]
  assign _T_68541 = $signed(_T_68540); // @[Modules.scala 37:46:@16840.4]
  assign _T_68611 = $signed(_T_62640) - $signed(io_in_751); // @[Modules.scala 46:47:@16913.4]
  assign _T_68612 = _T_68611[4:0]; // @[Modules.scala 46:47:@16914.4]
  assign _T_68613 = $signed(_T_68612); // @[Modules.scala 46:47:@16915.4]
  assign _T_68615 = $signed(5'sh0) - $signed(io_in_752); // @[Modules.scala 43:37:@16917.4]
  assign _T_68616 = _T_68615[4:0]; // @[Modules.scala 43:37:@16918.4]
  assign _T_68617 = $signed(_T_68616); // @[Modules.scala 43:37:@16919.4]
  assign _T_68618 = $signed(_T_68617) + $signed(io_in_753); // @[Modules.scala 43:47:@16920.4]
  assign _T_68619 = _T_68618[4:0]; // @[Modules.scala 43:47:@16921.4]
  assign _T_68620 = $signed(_T_68619); // @[Modules.scala 43:47:@16922.4]
  assign _T_68659 = $signed(_T_56326) + $signed(io_in_767); // @[Modules.scala 43:47:@16963.4]
  assign _T_68660 = _T_68659[4:0]; // @[Modules.scala 43:47:@16964.4]
  assign _T_68661 = $signed(_T_68660); // @[Modules.scala 43:47:@16965.4]
  assign _T_68672 = $signed(io_in_772) - $signed(io_in_773); // @[Modules.scala 40:46:@16978.4]
  assign _T_68673 = _T_68672[4:0]; // @[Modules.scala 40:46:@16979.4]
  assign _T_68674 = $signed(_T_68673); // @[Modules.scala 40:46:@16980.4]
  assign _T_68700 = $signed(_T_56367) - $signed(io_in_781); // @[Modules.scala 46:47:@17006.4]
  assign _T_68701 = _T_68700[4:0]; // @[Modules.scala 46:47:@17007.4]
  assign _T_68702 = $signed(_T_68701); // @[Modules.scala 46:47:@17008.4]
  assign buffer_4_1 = {{6{_T_66899[4]}},_T_66899}; // @[Modules.scala 32:22:@8.4]
  assign _T_68710 = $signed(buffer_3_0) + $signed(buffer_4_1); // @[Modules.scala 50:57:@17017.4]
  assign _T_68711 = _T_68710[10:0]; // @[Modules.scala 50:57:@17018.4]
  assign buffer_4_392 = $signed(_T_68711); // @[Modules.scala 50:57:@17019.4]
  assign _T_68713 = $signed(buffer_0_2) + $signed(buffer_1_3); // @[Modules.scala 50:57:@17021.4]
  assign _T_68714 = _T_68713[10:0]; // @[Modules.scala 50:57:@17022.4]
  assign buffer_4_393 = $signed(_T_68714); // @[Modules.scala 50:57:@17023.4]
  assign buffer_4_5 = {{6{_T_66923[4]}},_T_66923}; // @[Modules.scala 32:22:@8.4]
  assign _T_68716 = $signed(buffer_3_4) + $signed(buffer_4_5); // @[Modules.scala 50:57:@17025.4]
  assign _T_68717 = _T_68716[10:0]; // @[Modules.scala 50:57:@17026.4]
  assign buffer_4_394 = $signed(_T_68717); // @[Modules.scala 50:57:@17027.4]
  assign _T_68719 = $signed(buffer_0_6) + $signed(buffer_1_7); // @[Modules.scala 50:57:@17029.4]
  assign _T_68720 = _T_68719[10:0]; // @[Modules.scala 50:57:@17030.4]
  assign buffer_4_395 = $signed(_T_68720); // @[Modules.scala 50:57:@17031.4]
  assign buffer_4_8 = {{6{_T_66940[4]}},_T_66940}; // @[Modules.scala 32:22:@8.4]
  assign _T_68722 = $signed(buffer_4_8) + $signed(buffer_1_9); // @[Modules.scala 50:57:@17033.4]
  assign _T_68723 = _T_68722[10:0]; // @[Modules.scala 50:57:@17034.4]
  assign buffer_4_396 = $signed(_T_68723); // @[Modules.scala 50:57:@17035.4]
  assign buffer_4_11 = {{6{_T_66953[4]}},_T_66953}; // @[Modules.scala 32:22:@8.4]
  assign _T_68725 = $signed(buffer_0_10) + $signed(buffer_4_11); // @[Modules.scala 50:57:@17037.4]
  assign _T_68726 = _T_68725[10:0]; // @[Modules.scala 50:57:@17038.4]
  assign buffer_4_397 = $signed(_T_68726); // @[Modules.scala 50:57:@17039.4]
  assign buffer_4_13 = {{6{_T_66963[4]}},_T_66963}; // @[Modules.scala 32:22:@8.4]
  assign _T_68728 = $signed(buffer_3_12) + $signed(buffer_4_13); // @[Modules.scala 50:57:@17041.4]
  assign _T_68729 = _T_68728[10:0]; // @[Modules.scala 50:57:@17042.4]
  assign buffer_4_398 = $signed(_T_68729); // @[Modules.scala 50:57:@17043.4]
  assign buffer_4_14 = {{6{_T_66970[4]}},_T_66970}; // @[Modules.scala 32:22:@8.4]
  assign _T_68731 = $signed(buffer_4_14) + $signed(buffer_2_15); // @[Modules.scala 50:57:@17045.4]
  assign _T_68732 = _T_68731[10:0]; // @[Modules.scala 50:57:@17046.4]
  assign buffer_4_399 = $signed(_T_68732); // @[Modules.scala 50:57:@17047.4]
  assign _T_68740 = $signed(buffer_1_20) + $signed(buffer_0_21); // @[Modules.scala 50:57:@17057.4]
  assign _T_68741 = _T_68740[10:0]; // @[Modules.scala 50:57:@17058.4]
  assign buffer_4_402 = $signed(_T_68741); // @[Modules.scala 50:57:@17059.4]
  assign buffer_4_22 = {{6{_T_67002[4]}},_T_67002}; // @[Modules.scala 32:22:@8.4]
  assign _T_68743 = $signed(buffer_4_22) + $signed(buffer_0_23); // @[Modules.scala 50:57:@17061.4]
  assign _T_68744 = _T_68743[10:0]; // @[Modules.scala 50:57:@17062.4]
  assign buffer_4_403 = $signed(_T_68744); // @[Modules.scala 50:57:@17063.4]
  assign _T_68749 = $signed(buffer_2_26) + $signed(buffer_0_27); // @[Modules.scala 50:57:@17069.4]
  assign _T_68750 = _T_68749[10:0]; // @[Modules.scala 50:57:@17070.4]
  assign buffer_4_405 = $signed(_T_68750); // @[Modules.scala 50:57:@17071.4]
  assign _T_68773 = $signed(buffer_1_42) + $signed(buffer_0_43); // @[Modules.scala 50:57:@17101.4]
  assign _T_68774 = _T_68773[10:0]; // @[Modules.scala 50:57:@17102.4]
  assign buffer_4_413 = $signed(_T_68774); // @[Modules.scala 50:57:@17103.4]
  assign buffer_4_44 = {{6{_T_67104[4]}},_T_67104}; // @[Modules.scala 32:22:@8.4]
  assign _T_68776 = $signed(buffer_4_44) + $signed(buffer_0_45); // @[Modules.scala 50:57:@17105.4]
  assign _T_68777 = _T_68776[10:0]; // @[Modules.scala 50:57:@17106.4]
  assign buffer_4_414 = $signed(_T_68777); // @[Modules.scala 50:57:@17107.4]
  assign _T_68794 = $signed(buffer_1_56) + $signed(buffer_0_57); // @[Modules.scala 50:57:@17129.4]
  assign _T_68795 = _T_68794[10:0]; // @[Modules.scala 50:57:@17130.4]
  assign buffer_4_420 = $signed(_T_68795); // @[Modules.scala 50:57:@17131.4]
  assign buffer_4_58 = {{6{_T_67158[4]}},_T_67158}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_59 = {{6{_T_67165[4]}},_T_67165}; // @[Modules.scala 32:22:@8.4]
  assign _T_68797 = $signed(buffer_4_58) + $signed(buffer_4_59); // @[Modules.scala 50:57:@17133.4]
  assign _T_68798 = _T_68797[10:0]; // @[Modules.scala 50:57:@17134.4]
  assign buffer_4_421 = $signed(_T_68798); // @[Modules.scala 50:57:@17135.4]
  assign buffer_4_61 = {{6{_T_67171[4]}},_T_67171}; // @[Modules.scala 32:22:@8.4]
  assign _T_68800 = $signed(buffer_3_60) + $signed(buffer_4_61); // @[Modules.scala 50:57:@17137.4]
  assign _T_68801 = _T_68800[10:0]; // @[Modules.scala 50:57:@17138.4]
  assign buffer_4_422 = $signed(_T_68801); // @[Modules.scala 50:57:@17139.4]
  assign _T_68803 = $signed(buffer_0_62) + $signed(buffer_3_63); // @[Modules.scala 50:57:@17141.4]
  assign _T_68804 = _T_68803[10:0]; // @[Modules.scala 50:57:@17142.4]
  assign buffer_4_423 = $signed(_T_68804); // @[Modules.scala 50:57:@17143.4]
  assign buffer_4_64 = {{6{_T_67184[4]}},_T_67184}; // @[Modules.scala 32:22:@8.4]
  assign _T_68806 = $signed(buffer_4_64) + $signed(buffer_2_65); // @[Modules.scala 50:57:@17145.4]
  assign _T_68807 = _T_68806[10:0]; // @[Modules.scala 50:57:@17146.4]
  assign buffer_4_424 = $signed(_T_68807); // @[Modules.scala 50:57:@17147.4]
  assign buffer_4_67 = {{6{_T_67205[4]}},_T_67205}; // @[Modules.scala 32:22:@8.4]
  assign _T_68809 = $signed(buffer_3_66) + $signed(buffer_4_67); // @[Modules.scala 50:57:@17149.4]
  assign _T_68810 = _T_68809[10:0]; // @[Modules.scala 50:57:@17150.4]
  assign buffer_4_425 = $signed(_T_68810); // @[Modules.scala 50:57:@17151.4]
  assign buffer_4_69 = {{6{_T_67211[4]}},_T_67211}; // @[Modules.scala 32:22:@8.4]
  assign _T_68812 = $signed(buffer_1_68) + $signed(buffer_4_69); // @[Modules.scala 50:57:@17153.4]
  assign _T_68813 = _T_68812[10:0]; // @[Modules.scala 50:57:@17154.4]
  assign buffer_4_426 = $signed(_T_68813); // @[Modules.scala 50:57:@17155.4]
  assign _T_68815 = $signed(buffer_2_70) + $signed(buffer_0_71); // @[Modules.scala 50:57:@17157.4]
  assign _T_68816 = _T_68815[10:0]; // @[Modules.scala 50:57:@17158.4]
  assign buffer_4_427 = $signed(_T_68816); // @[Modules.scala 50:57:@17159.4]
  assign buffer_4_72 = {{6{_T_67228[4]}},_T_67228}; // @[Modules.scala 32:22:@8.4]
  assign _T_68818 = $signed(buffer_4_72) + $signed(buffer_0_73); // @[Modules.scala 50:57:@17161.4]
  assign _T_68819 = _T_68818[10:0]; // @[Modules.scala 50:57:@17162.4]
  assign buffer_4_428 = $signed(_T_68819); // @[Modules.scala 50:57:@17163.4]
  assign buffer_4_76 = {{6{_T_67240[4]}},_T_67240}; // @[Modules.scala 32:22:@8.4]
  assign _T_68824 = $signed(buffer_4_76) + $signed(buffer_3_77); // @[Modules.scala 50:57:@17169.4]
  assign _T_68825 = _T_68824[10:0]; // @[Modules.scala 50:57:@17170.4]
  assign buffer_4_430 = $signed(_T_68825); // @[Modules.scala 50:57:@17171.4]
  assign buffer_4_78 = {{6{_T_67246[4]}},_T_67246}; // @[Modules.scala 32:22:@8.4]
  assign _T_68827 = $signed(buffer_4_78) + $signed(buffer_3_79); // @[Modules.scala 50:57:@17173.4]
  assign _T_68828 = _T_68827[10:0]; // @[Modules.scala 50:57:@17174.4]
  assign buffer_4_431 = $signed(_T_68828); // @[Modules.scala 50:57:@17175.4]
  assign buffer_4_80 = {{6{_T_67252[4]}},_T_67252}; // @[Modules.scala 32:22:@8.4]
  assign _T_68830 = $signed(buffer_4_80) + $signed(buffer_1_81); // @[Modules.scala 50:57:@17177.4]
  assign _T_68831 = _T_68830[10:0]; // @[Modules.scala 50:57:@17178.4]
  assign buffer_4_432 = $signed(_T_68831); // @[Modules.scala 50:57:@17179.4]
  assign buffer_4_84 = {{6{_T_67268[4]}},_T_67268}; // @[Modules.scala 32:22:@8.4]
  assign _T_68836 = $signed(buffer_4_84) + $signed(buffer_0_85); // @[Modules.scala 50:57:@17185.4]
  assign _T_68837 = _T_68836[10:0]; // @[Modules.scala 50:57:@17186.4]
  assign buffer_4_434 = $signed(_T_68837); // @[Modules.scala 50:57:@17187.4]
  assign buffer_4_92 = {{6{_T_67308[4]}},_T_67308}; // @[Modules.scala 32:22:@8.4]
  assign _T_68848 = $signed(buffer_4_92) + $signed(buffer_0_93); // @[Modules.scala 50:57:@17201.4]
  assign _T_68849 = _T_68848[10:0]; // @[Modules.scala 50:57:@17202.4]
  assign buffer_4_438 = $signed(_T_68849); // @[Modules.scala 50:57:@17203.4]
  assign buffer_4_94 = {{6{_T_67314[4]}},_T_67314}; // @[Modules.scala 32:22:@8.4]
  assign _T_68851 = $signed(buffer_4_94) + $signed(buffer_2_95); // @[Modules.scala 50:57:@17205.4]
  assign _T_68852 = _T_68851[10:0]; // @[Modules.scala 50:57:@17206.4]
  assign buffer_4_439 = $signed(_T_68852); // @[Modules.scala 50:57:@17207.4]
  assign _T_68857 = $signed(buffer_1_98) + $signed(buffer_2_99); // @[Modules.scala 50:57:@17213.4]
  assign _T_68858 = _T_68857[10:0]; // @[Modules.scala 50:57:@17214.4]
  assign buffer_4_441 = $signed(_T_68858); // @[Modules.scala 50:57:@17215.4]
  assign buffer_4_101 = {{6{_T_67347[4]}},_T_67347}; // @[Modules.scala 32:22:@8.4]
  assign _T_68860 = $signed(buffer_1_100) + $signed(buffer_4_101); // @[Modules.scala 50:57:@17217.4]
  assign _T_68861 = _T_68860[10:0]; // @[Modules.scala 50:57:@17218.4]
  assign buffer_4_442 = $signed(_T_68861); // @[Modules.scala 50:57:@17219.4]
  assign buffer_4_102 = {{6{_T_67350[4]}},_T_67350}; // @[Modules.scala 32:22:@8.4]
  assign _T_68863 = $signed(buffer_4_102) + $signed(buffer_1_103); // @[Modules.scala 50:57:@17221.4]
  assign _T_68864 = _T_68863[10:0]; // @[Modules.scala 50:57:@17222.4]
  assign buffer_4_443 = $signed(_T_68864); // @[Modules.scala 50:57:@17223.4]
  assign buffer_4_105 = {{6{_T_67367[4]}},_T_67367}; // @[Modules.scala 32:22:@8.4]
  assign _T_68866 = $signed(buffer_2_104) + $signed(buffer_4_105); // @[Modules.scala 50:57:@17225.4]
  assign _T_68867 = _T_68866[10:0]; // @[Modules.scala 50:57:@17226.4]
  assign buffer_4_444 = $signed(_T_68867); // @[Modules.scala 50:57:@17227.4]
  assign buffer_4_106 = {{6{_T_67374[4]}},_T_67374}; // @[Modules.scala 32:22:@8.4]
  assign _T_68869 = $signed(buffer_4_106) + $signed(buffer_0_107); // @[Modules.scala 50:57:@17229.4]
  assign _T_68870 = _T_68869[10:0]; // @[Modules.scala 50:57:@17230.4]
  assign buffer_4_445 = $signed(_T_68870); // @[Modules.scala 50:57:@17231.4]
  assign buffer_4_114 = {{6{_T_67414[4]}},_T_67414}; // @[Modules.scala 32:22:@8.4]
  assign _T_68881 = $signed(buffer_4_114) + $signed(buffer_0_115); // @[Modules.scala 50:57:@17245.4]
  assign _T_68882 = _T_68881[10:0]; // @[Modules.scala 50:57:@17246.4]
  assign buffer_4_449 = $signed(_T_68882); // @[Modules.scala 50:57:@17247.4]
  assign buffer_4_116 = {{6{_T_67424[4]}},_T_67424}; // @[Modules.scala 32:22:@8.4]
  assign _T_68884 = $signed(buffer_4_116) + $signed(buffer_3_117); // @[Modules.scala 50:57:@17249.4]
  assign _T_68885 = _T_68884[10:0]; // @[Modules.scala 50:57:@17250.4]
  assign buffer_4_450 = $signed(_T_68885); // @[Modules.scala 50:57:@17251.4]
  assign buffer_4_121 = {{6{_T_67455[4]}},_T_67455}; // @[Modules.scala 32:22:@8.4]
  assign _T_68890 = $signed(buffer_0_120) + $signed(buffer_4_121); // @[Modules.scala 50:57:@17257.4]
  assign _T_68891 = _T_68890[10:0]; // @[Modules.scala 50:57:@17258.4]
  assign buffer_4_452 = $signed(_T_68891); // @[Modules.scala 50:57:@17259.4]
  assign buffer_4_122 = {{6{_T_67458[4]}},_T_67458}; // @[Modules.scala 32:22:@8.4]
  assign _T_68893 = $signed(buffer_4_122) + $signed(buffer_3_123); // @[Modules.scala 50:57:@17261.4]
  assign _T_68894 = _T_68893[10:0]; // @[Modules.scala 50:57:@17262.4]
  assign buffer_4_453 = $signed(_T_68894); // @[Modules.scala 50:57:@17263.4]
  assign buffer_4_128 = {{6{_T_67488[4]}},_T_67488}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_129 = {{6{_T_67491[4]}},_T_67491}; // @[Modules.scala 32:22:@8.4]
  assign _T_68902 = $signed(buffer_4_128) + $signed(buffer_4_129); // @[Modules.scala 50:57:@17273.4]
  assign _T_68903 = _T_68902[10:0]; // @[Modules.scala 50:57:@17274.4]
  assign buffer_4_456 = $signed(_T_68903); // @[Modules.scala 50:57:@17275.4]
  assign buffer_4_130 = {{6{_T_67494[4]}},_T_67494}; // @[Modules.scala 32:22:@8.4]
  assign _T_68905 = $signed(buffer_4_130) + $signed(buffer_0_131); // @[Modules.scala 50:57:@17277.4]
  assign _T_68906 = _T_68905[10:0]; // @[Modules.scala 50:57:@17278.4]
  assign buffer_4_457 = $signed(_T_68906); // @[Modules.scala 50:57:@17279.4]
  assign _T_68920 = $signed(buffer_1_140) + $signed(buffer_0_141); // @[Modules.scala 50:57:@17297.4]
  assign _T_68921 = _T_68920[10:0]; // @[Modules.scala 50:57:@17298.4]
  assign buffer_4_462 = $signed(_T_68921); // @[Modules.scala 50:57:@17299.4]
  assign _T_68923 = $signed(buffer_3_142) + $signed(buffer_2_143); // @[Modules.scala 50:57:@17301.4]
  assign _T_68924 = _T_68923[10:0]; // @[Modules.scala 50:57:@17302.4]
  assign buffer_4_463 = $signed(_T_68924); // @[Modules.scala 50:57:@17303.4]
  assign buffer_4_148 = {{6{_T_67596[4]}},_T_67596}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_149 = {{6{_T_67599[4]}},_T_67599}; // @[Modules.scala 32:22:@8.4]
  assign _T_68932 = $signed(buffer_4_148) + $signed(buffer_4_149); // @[Modules.scala 50:57:@17313.4]
  assign _T_68933 = _T_68932[10:0]; // @[Modules.scala 50:57:@17314.4]
  assign buffer_4_466 = $signed(_T_68933); // @[Modules.scala 50:57:@17315.4]
  assign buffer_4_151 = {{6{_T_67609[4]}},_T_67609}; // @[Modules.scala 32:22:@8.4]
  assign _T_68935 = $signed(buffer_0_150) + $signed(buffer_4_151); // @[Modules.scala 50:57:@17317.4]
  assign _T_68936 = _T_68935[10:0]; // @[Modules.scala 50:57:@17318.4]
  assign buffer_4_467 = $signed(_T_68936); // @[Modules.scala 50:57:@17319.4]
  assign buffer_4_154 = {{6{_T_67618[4]}},_T_67618}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_155 = {{6{_T_67625[4]}},_T_67625}; // @[Modules.scala 32:22:@8.4]
  assign _T_68941 = $signed(buffer_4_154) + $signed(buffer_4_155); // @[Modules.scala 50:57:@17325.4]
  assign _T_68942 = _T_68941[10:0]; // @[Modules.scala 50:57:@17326.4]
  assign buffer_4_469 = $signed(_T_68942); // @[Modules.scala 50:57:@17327.4]
  assign _T_68950 = $signed(buffer_2_160) + $signed(buffer_0_161); // @[Modules.scala 50:57:@17337.4]
  assign _T_68951 = _T_68950[10:0]; // @[Modules.scala 50:57:@17338.4]
  assign buffer_4_472 = $signed(_T_68951); // @[Modules.scala 50:57:@17339.4]
  assign _T_68959 = $signed(buffer_1_166) + $signed(buffer_3_167); // @[Modules.scala 50:57:@17349.4]
  assign _T_68960 = _T_68959[10:0]; // @[Modules.scala 50:57:@17350.4]
  assign buffer_4_475 = $signed(_T_68960); // @[Modules.scala 50:57:@17351.4]
  assign buffer_4_172 = {{6{_T_67720[4]}},_T_67720}; // @[Modules.scala 32:22:@8.4]
  assign _T_68968 = $signed(buffer_4_172) + $signed(buffer_0_173); // @[Modules.scala 50:57:@17361.4]
  assign _T_68969 = _T_68968[10:0]; // @[Modules.scala 50:57:@17362.4]
  assign buffer_4_478 = $signed(_T_68969); // @[Modules.scala 50:57:@17363.4]
  assign buffer_4_176 = {{6{_T_67736[4]}},_T_67736}; // @[Modules.scala 32:22:@8.4]
  assign _T_68974 = $signed(buffer_4_176) + $signed(buffer_1_177); // @[Modules.scala 50:57:@17369.4]
  assign _T_68975 = _T_68974[10:0]; // @[Modules.scala 50:57:@17370.4]
  assign buffer_4_480 = $signed(_T_68975); // @[Modules.scala 50:57:@17371.4]
  assign _T_68980 = $signed(buffer_1_180) + $signed(buffer_2_181); // @[Modules.scala 50:57:@17377.4]
  assign _T_68981 = _T_68980[10:0]; // @[Modules.scala 50:57:@17378.4]
  assign buffer_4_482 = $signed(_T_68981); // @[Modules.scala 50:57:@17379.4]
  assign buffer_4_182 = {{6{_T_67766[4]}},_T_67766}; // @[Modules.scala 32:22:@8.4]
  assign _T_68983 = $signed(buffer_4_182) + $signed(buffer_0_183); // @[Modules.scala 50:57:@17381.4]
  assign _T_68984 = _T_68983[10:0]; // @[Modules.scala 50:57:@17382.4]
  assign buffer_4_483 = $signed(_T_68984); // @[Modules.scala 50:57:@17383.4]
  assign buffer_4_185 = {{6{_T_67783[4]}},_T_67783}; // @[Modules.scala 32:22:@8.4]
  assign _T_68986 = $signed(buffer_3_184) + $signed(buffer_4_185); // @[Modules.scala 50:57:@17385.4]
  assign _T_68987 = _T_68986[10:0]; // @[Modules.scala 50:57:@17386.4]
  assign buffer_4_484 = $signed(_T_68987); // @[Modules.scala 50:57:@17387.4]
  assign buffer_4_190 = {{6{_T_67802[4]}},_T_67802}; // @[Modules.scala 32:22:@8.4]
  assign _T_68995 = $signed(buffer_4_190) + $signed(buffer_1_191); // @[Modules.scala 50:57:@17397.4]
  assign _T_68996 = _T_68995[10:0]; // @[Modules.scala 50:57:@17398.4]
  assign buffer_4_487 = $signed(_T_68996); // @[Modules.scala 50:57:@17399.4]
  assign _T_68998 = $signed(buffer_3_192) + $signed(buffer_0_193); // @[Modules.scala 50:57:@17401.4]
  assign _T_68999 = _T_68998[10:0]; // @[Modules.scala 50:57:@17402.4]
  assign buffer_4_488 = $signed(_T_68999); // @[Modules.scala 50:57:@17403.4]
  assign buffer_4_194 = {{6{_T_67822[4]}},_T_67822}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_195 = {{6{_T_67825[4]}},_T_67825}; // @[Modules.scala 32:22:@8.4]
  assign _T_69001 = $signed(buffer_4_194) + $signed(buffer_4_195); // @[Modules.scala 50:57:@17405.4]
  assign _T_69002 = _T_69001[10:0]; // @[Modules.scala 50:57:@17406.4]
  assign buffer_4_489 = $signed(_T_69002); // @[Modules.scala 50:57:@17407.4]
  assign buffer_4_196 = {{6{_T_67828[4]}},_T_67828}; // @[Modules.scala 32:22:@8.4]
  assign _T_69004 = $signed(buffer_4_196) + $signed(buffer_0_197); // @[Modules.scala 50:57:@17409.4]
  assign _T_69005 = _T_69004[10:0]; // @[Modules.scala 50:57:@17410.4]
  assign buffer_4_490 = $signed(_T_69005); // @[Modules.scala 50:57:@17411.4]
  assign buffer_4_199 = {{6{_T_67849[4]}},_T_67849}; // @[Modules.scala 32:22:@8.4]
  assign _T_69007 = $signed(buffer_1_198) + $signed(buffer_4_199); // @[Modules.scala 50:57:@17413.4]
  assign _T_69008 = _T_69007[10:0]; // @[Modules.scala 50:57:@17414.4]
  assign buffer_4_491 = $signed(_T_69008); // @[Modules.scala 50:57:@17415.4]
  assign _T_69010 = $signed(buffer_3_200) + $signed(buffer_0_201); // @[Modules.scala 50:57:@17417.4]
  assign _T_69011 = _T_69010[10:0]; // @[Modules.scala 50:57:@17418.4]
  assign buffer_4_492 = $signed(_T_69011); // @[Modules.scala 50:57:@17419.4]
  assign buffer_4_203 = {{6{_T_67869[4]}},_T_67869}; // @[Modules.scala 32:22:@8.4]
  assign _T_69013 = $signed(buffer_0_202) + $signed(buffer_4_203); // @[Modules.scala 50:57:@17421.4]
  assign _T_69014 = _T_69013[10:0]; // @[Modules.scala 50:57:@17422.4]
  assign buffer_4_493 = $signed(_T_69014); // @[Modules.scala 50:57:@17423.4]
  assign _T_69016 = $signed(buffer_0_204) + $signed(buffer_3_205); // @[Modules.scala 50:57:@17425.4]
  assign _T_69017 = _T_69016[10:0]; // @[Modules.scala 50:57:@17426.4]
  assign buffer_4_494 = $signed(_T_69017); // @[Modules.scala 50:57:@17427.4]
  assign buffer_4_206 = {{6{_T_67878[4]}},_T_67878}; // @[Modules.scala 32:22:@8.4]
  assign _T_69019 = $signed(buffer_4_206) + $signed(buffer_0_207); // @[Modules.scala 50:57:@17429.4]
  assign _T_69020 = _T_69019[10:0]; // @[Modules.scala 50:57:@17430.4]
  assign buffer_4_495 = $signed(_T_69020); // @[Modules.scala 50:57:@17431.4]
  assign buffer_4_208 = {{6{_T_67884[4]}},_T_67884}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_209 = {{6{_T_67887[4]}},_T_67887}; // @[Modules.scala 32:22:@8.4]
  assign _T_69022 = $signed(buffer_4_208) + $signed(buffer_4_209); // @[Modules.scala 50:57:@17433.4]
  assign _T_69023 = _T_69022[10:0]; // @[Modules.scala 50:57:@17434.4]
  assign buffer_4_496 = $signed(_T_69023); // @[Modules.scala 50:57:@17435.4]
  assign buffer_4_210 = {{6{_T_67890[4]}},_T_67890}; // @[Modules.scala 32:22:@8.4]
  assign _T_69025 = $signed(buffer_4_210) + $signed(buffer_2_211); // @[Modules.scala 50:57:@17437.4]
  assign _T_69026 = _T_69025[10:0]; // @[Modules.scala 50:57:@17438.4]
  assign buffer_4_497 = $signed(_T_69026); // @[Modules.scala 50:57:@17439.4]
  assign buffer_4_216 = {{6{_T_67912[4]}},_T_67912}; // @[Modules.scala 32:22:@8.4]
  assign _T_69034 = $signed(buffer_4_216) + $signed(buffer_0_217); // @[Modules.scala 50:57:@17449.4]
  assign _T_69035 = _T_69034[10:0]; // @[Modules.scala 50:57:@17450.4]
  assign buffer_4_500 = $signed(_T_69035); // @[Modules.scala 50:57:@17451.4]
  assign buffer_4_218 = {{6{_T_67918[4]}},_T_67918}; // @[Modules.scala 32:22:@8.4]
  assign _T_69037 = $signed(buffer_4_218) + $signed(buffer_1_219); // @[Modules.scala 50:57:@17453.4]
  assign _T_69038 = _T_69037[10:0]; // @[Modules.scala 50:57:@17454.4]
  assign buffer_4_501 = $signed(_T_69038); // @[Modules.scala 50:57:@17455.4]
  assign _T_69040 = $signed(buffer_3_220) + $signed(buffer_1_221); // @[Modules.scala 50:57:@17457.4]
  assign _T_69041 = _T_69040[10:0]; // @[Modules.scala 50:57:@17458.4]
  assign buffer_4_502 = $signed(_T_69041); // @[Modules.scala 50:57:@17459.4]
  assign buffer_4_227 = {{6{_T_67961[4]}},_T_67961}; // @[Modules.scala 32:22:@8.4]
  assign _T_69049 = $signed(buffer_0_226) + $signed(buffer_4_227); // @[Modules.scala 50:57:@17469.4]
  assign _T_69050 = _T_69049[10:0]; // @[Modules.scala 50:57:@17470.4]
  assign buffer_4_505 = $signed(_T_69050); // @[Modules.scala 50:57:@17471.4]
  assign buffer_4_231 = {{6{_T_67981[4]}},_T_67981}; // @[Modules.scala 32:22:@8.4]
  assign _T_69055 = $signed(buffer_2_230) + $signed(buffer_4_231); // @[Modules.scala 50:57:@17477.4]
  assign _T_69056 = _T_69055[10:0]; // @[Modules.scala 50:57:@17478.4]
  assign buffer_4_507 = $signed(_T_69056); // @[Modules.scala 50:57:@17479.4]
  assign _T_69058 = $signed(buffer_2_232) + $signed(buffer_1_233); // @[Modules.scala 50:57:@17481.4]
  assign _T_69059 = _T_69058[10:0]; // @[Modules.scala 50:57:@17482.4]
  assign buffer_4_508 = $signed(_T_69059); // @[Modules.scala 50:57:@17483.4]
  assign _T_69067 = $signed(buffer_2_238) + $signed(buffer_1_239); // @[Modules.scala 50:57:@17493.4]
  assign _T_69068 = _T_69067[10:0]; // @[Modules.scala 50:57:@17494.4]
  assign buffer_4_511 = $signed(_T_69068); // @[Modules.scala 50:57:@17495.4]
  assign _T_69070 = $signed(buffer_3_240) + $signed(buffer_0_241); // @[Modules.scala 50:57:@17497.4]
  assign _T_69071 = _T_69070[10:0]; // @[Modules.scala 50:57:@17498.4]
  assign buffer_4_512 = $signed(_T_69071); // @[Modules.scala 50:57:@17499.4]
  assign buffer_4_243 = {{6{_T_68029[4]}},_T_68029}; // @[Modules.scala 32:22:@8.4]
  assign _T_69073 = $signed(buffer_0_242) + $signed(buffer_4_243); // @[Modules.scala 50:57:@17501.4]
  assign _T_69074 = _T_69073[10:0]; // @[Modules.scala 50:57:@17502.4]
  assign buffer_4_513 = $signed(_T_69074); // @[Modules.scala 50:57:@17503.4]
  assign buffer_4_246 = {{6{_T_68046[4]}},_T_68046}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_247 = {{6{_T_68053[4]}},_T_68053}; // @[Modules.scala 32:22:@8.4]
  assign _T_69079 = $signed(buffer_4_246) + $signed(buffer_4_247); // @[Modules.scala 50:57:@17509.4]
  assign _T_69080 = _T_69079[10:0]; // @[Modules.scala 50:57:@17510.4]
  assign buffer_4_515 = $signed(_T_69080); // @[Modules.scala 50:57:@17511.4]
  assign _T_69088 = $signed(buffer_0_252) + $signed(buffer_1_253); // @[Modules.scala 50:57:@17521.4]
  assign _T_69089 = _T_69088[10:0]; // @[Modules.scala 50:57:@17522.4]
  assign buffer_4_518 = $signed(_T_69089); // @[Modules.scala 50:57:@17523.4]
  assign buffer_4_256 = {{6{_T_68084[4]}},_T_68084}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_257 = {{6{_T_68087[4]}},_T_68087}; // @[Modules.scala 32:22:@8.4]
  assign _T_69094 = $signed(buffer_4_256) + $signed(buffer_4_257); // @[Modules.scala 50:57:@17529.4]
  assign _T_69095 = _T_69094[10:0]; // @[Modules.scala 50:57:@17530.4]
  assign buffer_4_520 = $signed(_T_69095); // @[Modules.scala 50:57:@17531.4]
  assign buffer_4_259 = {{6{_T_68097[4]}},_T_68097}; // @[Modules.scala 32:22:@8.4]
  assign _T_69097 = $signed(buffer_0_258) + $signed(buffer_4_259); // @[Modules.scala 50:57:@17533.4]
  assign _T_69098 = _T_69097[10:0]; // @[Modules.scala 50:57:@17534.4]
  assign buffer_4_521 = $signed(_T_69098); // @[Modules.scala 50:57:@17535.4]
  assign buffer_4_260 = {{6{_T_68100[4]}},_T_68100}; // @[Modules.scala 32:22:@8.4]
  assign _T_69100 = $signed(buffer_4_260) + $signed(buffer_1_261); // @[Modules.scala 50:57:@17537.4]
  assign _T_69101 = _T_69100[10:0]; // @[Modules.scala 50:57:@17538.4]
  assign buffer_4_522 = $signed(_T_69101); // @[Modules.scala 50:57:@17539.4]
  assign _T_69103 = $signed(buffer_1_262) + $signed(buffer_0_263); // @[Modules.scala 50:57:@17541.4]
  assign _T_69104 = _T_69103[10:0]; // @[Modules.scala 50:57:@17542.4]
  assign buffer_4_523 = $signed(_T_69104); // @[Modules.scala 50:57:@17543.4]
  assign _T_69109 = $signed(buffer_2_266) + $signed(buffer_0_267); // @[Modules.scala 50:57:@17549.4]
  assign _T_69110 = _T_69109[10:0]; // @[Modules.scala 50:57:@17550.4]
  assign buffer_4_525 = $signed(_T_69110); // @[Modules.scala 50:57:@17551.4]
  assign buffer_4_272 = {{6{_T_68148[4]}},_T_68148}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_273 = {{6{_T_68151[4]}},_T_68151}; // @[Modules.scala 32:22:@8.4]
  assign _T_69118 = $signed(buffer_4_272) + $signed(buffer_4_273); // @[Modules.scala 50:57:@17561.4]
  assign _T_69119 = _T_69118[10:0]; // @[Modules.scala 50:57:@17562.4]
  assign buffer_4_528 = $signed(_T_69119); // @[Modules.scala 50:57:@17563.4]
  assign _T_69127 = $signed(buffer_3_278) + $signed(buffer_1_279); // @[Modules.scala 50:57:@17573.4]
  assign _T_69128 = _T_69127[10:0]; // @[Modules.scala 50:57:@17574.4]
  assign buffer_4_531 = $signed(_T_69128); // @[Modules.scala 50:57:@17575.4]
  assign _T_69139 = $signed(buffer_1_286) + $signed(buffer_0_287); // @[Modules.scala 50:57:@17589.4]
  assign _T_69140 = _T_69139[10:0]; // @[Modules.scala 50:57:@17590.4]
  assign buffer_4_535 = $signed(_T_69140); // @[Modules.scala 50:57:@17591.4]
  assign buffer_4_290 = {{6{_T_68214[4]}},_T_68214}; // @[Modules.scala 32:22:@8.4]
  assign _T_69145 = $signed(buffer_4_290) + $signed(buffer_3_291); // @[Modules.scala 50:57:@17597.4]
  assign _T_69146 = _T_69145[10:0]; // @[Modules.scala 50:57:@17598.4]
  assign buffer_4_537 = $signed(_T_69146); // @[Modules.scala 50:57:@17599.4]
  assign buffer_4_292 = {{6{_T_68220[4]}},_T_68220}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_293 = {{6{_T_68227[4]}},_T_68227}; // @[Modules.scala 32:22:@8.4]
  assign _T_69148 = $signed(buffer_4_292) + $signed(buffer_4_293); // @[Modules.scala 50:57:@17601.4]
  assign _T_69149 = _T_69148[10:0]; // @[Modules.scala 50:57:@17602.4]
  assign buffer_4_538 = $signed(_T_69149); // @[Modules.scala 50:57:@17603.4]
  assign _T_69151 = $signed(buffer_0_294) + $signed(buffer_1_295); // @[Modules.scala 50:57:@17605.4]
  assign _T_69152 = _T_69151[10:0]; // @[Modules.scala 50:57:@17606.4]
  assign buffer_4_539 = $signed(_T_69152); // @[Modules.scala 50:57:@17607.4]
  assign _T_69157 = $signed(buffer_2_298) + $signed(buffer_1_299); // @[Modules.scala 50:57:@17613.4]
  assign _T_69158 = _T_69157[10:0]; // @[Modules.scala 50:57:@17614.4]
  assign buffer_4_541 = $signed(_T_69158); // @[Modules.scala 50:57:@17615.4]
  assign _T_69166 = $signed(buffer_2_304) + $signed(buffer_3_305); // @[Modules.scala 50:57:@17625.4]
  assign _T_69167 = _T_69166[10:0]; // @[Modules.scala 50:57:@17626.4]
  assign buffer_4_544 = $signed(_T_69167); // @[Modules.scala 50:57:@17627.4]
  assign buffer_4_306 = {{6{_T_68270[4]}},_T_68270}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_307 = {{6{_T_68273[4]}},_T_68273}; // @[Modules.scala 32:22:@8.4]
  assign _T_69169 = $signed(buffer_4_306) + $signed(buffer_4_307); // @[Modules.scala 50:57:@17629.4]
  assign _T_69170 = _T_69169[10:0]; // @[Modules.scala 50:57:@17630.4]
  assign buffer_4_545 = $signed(_T_69170); // @[Modules.scala 50:57:@17631.4]
  assign buffer_4_311 = {{6{_T_68289[4]}},_T_68289}; // @[Modules.scala 32:22:@8.4]
  assign _T_69175 = $signed(buffer_3_310) + $signed(buffer_4_311); // @[Modules.scala 50:57:@17637.4]
  assign _T_69176 = _T_69175[10:0]; // @[Modules.scala 50:57:@17638.4]
  assign buffer_4_547 = $signed(_T_69176); // @[Modules.scala 50:57:@17639.4]
  assign _T_69178 = $signed(buffer_0_312) + $signed(buffer_1_313); // @[Modules.scala 50:57:@17641.4]
  assign _T_69179 = _T_69178[10:0]; // @[Modules.scala 50:57:@17642.4]
  assign buffer_4_548 = $signed(_T_69179); // @[Modules.scala 50:57:@17643.4]
  assign buffer_4_316 = {{6{_T_68312[4]}},_T_68312}; // @[Modules.scala 32:22:@8.4]
  assign _T_69184 = $signed(buffer_4_316) + $signed(buffer_2_317); // @[Modules.scala 50:57:@17649.4]
  assign _T_69185 = _T_69184[10:0]; // @[Modules.scala 50:57:@17650.4]
  assign buffer_4_550 = $signed(_T_69185); // @[Modules.scala 50:57:@17651.4]
  assign _T_69190 = $signed(buffer_1_320) + $signed(buffer_0_321); // @[Modules.scala 50:57:@17657.4]
  assign _T_69191 = _T_69190[10:0]; // @[Modules.scala 50:57:@17658.4]
  assign buffer_4_552 = $signed(_T_69191); // @[Modules.scala 50:57:@17659.4]
  assign buffer_4_324 = {{6{_T_68348[4]}},_T_68348}; // @[Modules.scala 32:22:@8.4]
  assign _T_69196 = $signed(buffer_4_324) + $signed(buffer_0_325); // @[Modules.scala 50:57:@17665.4]
  assign _T_69197 = _T_69196[10:0]; // @[Modules.scala 50:57:@17666.4]
  assign buffer_4_554 = $signed(_T_69197); // @[Modules.scala 50:57:@17667.4]
  assign buffer_4_330 = {{6{_T_68370[4]}},_T_68370}; // @[Modules.scala 32:22:@8.4]
  assign _T_69205 = $signed(buffer_4_330) + $signed(buffer_1_331); // @[Modules.scala 50:57:@17677.4]
  assign _T_69206 = _T_69205[10:0]; // @[Modules.scala 50:57:@17678.4]
  assign buffer_4_557 = $signed(_T_69206); // @[Modules.scala 50:57:@17679.4]
  assign _T_69208 = $signed(buffer_0_332) + $signed(buffer_1_333); // @[Modules.scala 50:57:@17681.4]
  assign _T_69209 = _T_69208[10:0]; // @[Modules.scala 50:57:@17682.4]
  assign buffer_4_558 = $signed(_T_69209); // @[Modules.scala 50:57:@17683.4]
  assign buffer_4_334 = {{6{_T_68390[4]}},_T_68390}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_335 = {{6{_T_68397[4]}},_T_68397}; // @[Modules.scala 32:22:@8.4]
  assign _T_69211 = $signed(buffer_4_334) + $signed(buffer_4_335); // @[Modules.scala 50:57:@17685.4]
  assign _T_69212 = _T_69211[10:0]; // @[Modules.scala 50:57:@17686.4]
  assign buffer_4_559 = $signed(_T_69212); // @[Modules.scala 50:57:@17687.4]
  assign buffer_4_336 = {{6{_T_68400[4]}},_T_68400}; // @[Modules.scala 32:22:@8.4]
  assign _T_69214 = $signed(buffer_4_336) + $signed(buffer_1_337); // @[Modules.scala 50:57:@17689.4]
  assign _T_69215 = _T_69214[10:0]; // @[Modules.scala 50:57:@17690.4]
  assign buffer_4_560 = $signed(_T_69215); // @[Modules.scala 50:57:@17691.4]
  assign buffer_4_338 = {{6{_T_68406[4]}},_T_68406}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_339 = {{6{_T_68413[4]}},_T_68413}; // @[Modules.scala 32:22:@8.4]
  assign _T_69217 = $signed(buffer_4_338) + $signed(buffer_4_339); // @[Modules.scala 50:57:@17693.4]
  assign _T_69218 = _T_69217[10:0]; // @[Modules.scala 50:57:@17694.4]
  assign buffer_4_561 = $signed(_T_69218); // @[Modules.scala 50:57:@17695.4]
  assign _T_69223 = $signed(buffer_1_342) + $signed(buffer_3_343); // @[Modules.scala 50:57:@17701.4]
  assign _T_69224 = _T_69223[10:0]; // @[Modules.scala 50:57:@17702.4]
  assign buffer_4_563 = $signed(_T_69224); // @[Modules.scala 50:57:@17703.4]
  assign _T_69226 = $signed(buffer_0_344) + $signed(buffer_3_345); // @[Modules.scala 50:57:@17705.4]
  assign _T_69227 = _T_69226[10:0]; // @[Modules.scala 50:57:@17706.4]
  assign buffer_4_564 = $signed(_T_69227); // @[Modules.scala 50:57:@17707.4]
  assign buffer_4_348 = {{6{_T_68456[4]}},_T_68456}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_349 = {{6{_T_68459[4]}},_T_68459}; // @[Modules.scala 32:22:@8.4]
  assign _T_69232 = $signed(buffer_4_348) + $signed(buffer_4_349); // @[Modules.scala 50:57:@17713.4]
  assign _T_69233 = _T_69232[10:0]; // @[Modules.scala 50:57:@17714.4]
  assign buffer_4_566 = $signed(_T_69233); // @[Modules.scala 50:57:@17715.4]
  assign buffer_4_352 = {{6{_T_68468[4]}},_T_68468}; // @[Modules.scala 32:22:@8.4]
  assign _T_69238 = $signed(buffer_4_352) + $signed(buffer_2_353); // @[Modules.scala 50:57:@17721.4]
  assign _T_69239 = _T_69238[10:0]; // @[Modules.scala 50:57:@17722.4]
  assign buffer_4_568 = $signed(_T_69239); // @[Modules.scala 50:57:@17723.4]
  assign buffer_4_362 = {{6{_T_68538[4]}},_T_68538}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_363 = {{6{_T_68541[4]}},_T_68541}; // @[Modules.scala 32:22:@8.4]
  assign _T_69253 = $signed(buffer_4_362) + $signed(buffer_4_363); // @[Modules.scala 50:57:@17741.4]
  assign _T_69254 = _T_69253[10:0]; // @[Modules.scala 50:57:@17742.4]
  assign buffer_4_573 = $signed(_T_69254); // @[Modules.scala 50:57:@17743.4]
  assign buffer_4_375 = {{6{_T_68613[4]}},_T_68613}; // @[Modules.scala 32:22:@8.4]
  assign _T_69271 = $signed(buffer_3_374) + $signed(buffer_4_375); // @[Modules.scala 50:57:@17765.4]
  assign _T_69272 = _T_69271[10:0]; // @[Modules.scala 50:57:@17766.4]
  assign buffer_4_579 = $signed(_T_69272); // @[Modules.scala 50:57:@17767.4]
  assign buffer_4_376 = {{6{_T_68620[4]}},_T_68620}; // @[Modules.scala 32:22:@8.4]
  assign _T_69274 = $signed(buffer_4_376) + $signed(buffer_3_377); // @[Modules.scala 50:57:@17769.4]
  assign _T_69275 = _T_69274[10:0]; // @[Modules.scala 50:57:@17770.4]
  assign buffer_4_580 = $signed(_T_69275); // @[Modules.scala 50:57:@17771.4]
  assign _T_69277 = $signed(buffer_1_378) + $signed(buffer_0_379); // @[Modules.scala 50:57:@17773.4]
  assign _T_69278 = _T_69277[10:0]; // @[Modules.scala 50:57:@17774.4]
  assign buffer_4_581 = $signed(_T_69278); // @[Modules.scala 50:57:@17775.4]
  assign _T_69280 = $signed(buffer_1_380) + $signed(buffer_0_381); // @[Modules.scala 50:57:@17777.4]
  assign _T_69281 = _T_69280[10:0]; // @[Modules.scala 50:57:@17778.4]
  assign buffer_4_582 = $signed(_T_69281); // @[Modules.scala 50:57:@17779.4]
  assign buffer_4_383 = {{6{_T_68661[4]}},_T_68661}; // @[Modules.scala 32:22:@8.4]
  assign _T_69283 = $signed(buffer_0_382) + $signed(buffer_4_383); // @[Modules.scala 50:57:@17781.4]
  assign _T_69284 = _T_69283[10:0]; // @[Modules.scala 50:57:@17782.4]
  assign buffer_4_583 = $signed(_T_69284); // @[Modules.scala 50:57:@17783.4]
  assign _T_69286 = $signed(buffer_0_384) + $signed(buffer_1_385); // @[Modules.scala 50:57:@17785.4]
  assign _T_69287 = _T_69286[10:0]; // @[Modules.scala 50:57:@17786.4]
  assign buffer_4_584 = $signed(_T_69287); // @[Modules.scala 50:57:@17787.4]
  assign buffer_4_386 = {{6{_T_68674[4]}},_T_68674}; // @[Modules.scala 32:22:@8.4]
  assign _T_69289 = $signed(buffer_4_386) + $signed(buffer_0_387); // @[Modules.scala 50:57:@17789.4]
  assign _T_69290 = _T_69289[10:0]; // @[Modules.scala 50:57:@17790.4]
  assign buffer_4_585 = $signed(_T_69290); // @[Modules.scala 50:57:@17791.4]
  assign buffer_4_390 = {{6{_T_68702[4]}},_T_68702}; // @[Modules.scala 32:22:@8.4]
  assign _T_69295 = $signed(buffer_4_390) + $signed(buffer_2_391); // @[Modules.scala 50:57:@17797.4]
  assign _T_69296 = _T_69295[10:0]; // @[Modules.scala 50:57:@17798.4]
  assign buffer_4_587 = $signed(_T_69296); // @[Modules.scala 50:57:@17799.4]
  assign _T_69298 = $signed(buffer_4_392) + $signed(buffer_4_393); // @[Modules.scala 53:83:@17801.4]
  assign _T_69299 = _T_69298[10:0]; // @[Modules.scala 53:83:@17802.4]
  assign buffer_4_588 = $signed(_T_69299); // @[Modules.scala 53:83:@17803.4]
  assign _T_69301 = $signed(buffer_4_394) + $signed(buffer_4_395); // @[Modules.scala 53:83:@17805.4]
  assign _T_69302 = _T_69301[10:0]; // @[Modules.scala 53:83:@17806.4]
  assign buffer_4_589 = $signed(_T_69302); // @[Modules.scala 53:83:@17807.4]
  assign _T_69304 = $signed(buffer_4_396) + $signed(buffer_4_397); // @[Modules.scala 53:83:@17809.4]
  assign _T_69305 = _T_69304[10:0]; // @[Modules.scala 53:83:@17810.4]
  assign buffer_4_590 = $signed(_T_69305); // @[Modules.scala 53:83:@17811.4]
  assign _T_69307 = $signed(buffer_4_398) + $signed(buffer_4_399); // @[Modules.scala 53:83:@17813.4]
  assign _T_69308 = _T_69307[10:0]; // @[Modules.scala 53:83:@17814.4]
  assign buffer_4_591 = $signed(_T_69308); // @[Modules.scala 53:83:@17815.4]
  assign _T_69310 = $signed(buffer_0_400) + $signed(buffer_1_401); // @[Modules.scala 53:83:@17817.4]
  assign _T_69311 = _T_69310[10:0]; // @[Modules.scala 53:83:@17818.4]
  assign buffer_4_592 = $signed(_T_69311); // @[Modules.scala 53:83:@17819.4]
  assign _T_69313 = $signed(buffer_4_402) + $signed(buffer_4_403); // @[Modules.scala 53:83:@17821.4]
  assign _T_69314 = _T_69313[10:0]; // @[Modules.scala 53:83:@17822.4]
  assign buffer_4_593 = $signed(_T_69314); // @[Modules.scala 53:83:@17823.4]
  assign _T_69316 = $signed(buffer_1_404) + $signed(buffer_4_405); // @[Modules.scala 53:83:@17825.4]
  assign _T_69317 = _T_69316[10:0]; // @[Modules.scala 53:83:@17826.4]
  assign buffer_4_594 = $signed(_T_69317); // @[Modules.scala 53:83:@17827.4]
  assign _T_69319 = $signed(buffer_2_406) + $signed(buffer_0_407); // @[Modules.scala 53:83:@17829.4]
  assign _T_69320 = _T_69319[10:0]; // @[Modules.scala 53:83:@17830.4]
  assign buffer_4_595 = $signed(_T_69320); // @[Modules.scala 53:83:@17831.4]
  assign _T_69328 = $signed(buffer_2_412) + $signed(buffer_4_413); // @[Modules.scala 53:83:@17841.4]
  assign _T_69329 = _T_69328[10:0]; // @[Modules.scala 53:83:@17842.4]
  assign buffer_4_598 = $signed(_T_69329); // @[Modules.scala 53:83:@17843.4]
  assign _T_69331 = $signed(buffer_4_414) + $signed(buffer_1_415); // @[Modules.scala 53:83:@17845.4]
  assign _T_69332 = _T_69331[10:0]; // @[Modules.scala 53:83:@17846.4]
  assign buffer_4_599 = $signed(_T_69332); // @[Modules.scala 53:83:@17847.4]
  assign _T_69340 = $signed(buffer_4_420) + $signed(buffer_4_421); // @[Modules.scala 53:83:@17857.4]
  assign _T_69341 = _T_69340[10:0]; // @[Modules.scala 53:83:@17858.4]
  assign buffer_4_602 = $signed(_T_69341); // @[Modules.scala 53:83:@17859.4]
  assign _T_69343 = $signed(buffer_4_422) + $signed(buffer_4_423); // @[Modules.scala 53:83:@17861.4]
  assign _T_69344 = _T_69343[10:0]; // @[Modules.scala 53:83:@17862.4]
  assign buffer_4_603 = $signed(_T_69344); // @[Modules.scala 53:83:@17863.4]
  assign _T_69346 = $signed(buffer_4_424) + $signed(buffer_4_425); // @[Modules.scala 53:83:@17865.4]
  assign _T_69347 = _T_69346[10:0]; // @[Modules.scala 53:83:@17866.4]
  assign buffer_4_604 = $signed(_T_69347); // @[Modules.scala 53:83:@17867.4]
  assign _T_69349 = $signed(buffer_4_426) + $signed(buffer_4_427); // @[Modules.scala 53:83:@17869.4]
  assign _T_69350 = _T_69349[10:0]; // @[Modules.scala 53:83:@17870.4]
  assign buffer_4_605 = $signed(_T_69350); // @[Modules.scala 53:83:@17871.4]
  assign _T_69352 = $signed(buffer_4_428) + $signed(buffer_3_429); // @[Modules.scala 53:83:@17873.4]
  assign _T_69353 = _T_69352[10:0]; // @[Modules.scala 53:83:@17874.4]
  assign buffer_4_606 = $signed(_T_69353); // @[Modules.scala 53:83:@17875.4]
  assign _T_69355 = $signed(buffer_4_430) + $signed(buffer_4_431); // @[Modules.scala 53:83:@17877.4]
  assign _T_69356 = _T_69355[10:0]; // @[Modules.scala 53:83:@17878.4]
  assign buffer_4_607 = $signed(_T_69356); // @[Modules.scala 53:83:@17879.4]
  assign _T_69358 = $signed(buffer_4_432) + $signed(buffer_2_433); // @[Modules.scala 53:83:@17881.4]
  assign _T_69359 = _T_69358[10:0]; // @[Modules.scala 53:83:@17882.4]
  assign buffer_4_608 = $signed(_T_69359); // @[Modules.scala 53:83:@17883.4]
  assign _T_69361 = $signed(buffer_4_434) + $signed(buffer_3_435); // @[Modules.scala 53:83:@17885.4]
  assign _T_69362 = _T_69361[10:0]; // @[Modules.scala 53:83:@17886.4]
  assign buffer_4_609 = $signed(_T_69362); // @[Modules.scala 53:83:@17887.4]
  assign _T_69364 = $signed(buffer_1_436) + $signed(buffer_0_437); // @[Modules.scala 53:83:@17889.4]
  assign _T_69365 = _T_69364[10:0]; // @[Modules.scala 53:83:@17890.4]
  assign buffer_4_610 = $signed(_T_69365); // @[Modules.scala 53:83:@17891.4]
  assign _T_69367 = $signed(buffer_4_438) + $signed(buffer_4_439); // @[Modules.scala 53:83:@17893.4]
  assign _T_69368 = _T_69367[10:0]; // @[Modules.scala 53:83:@17894.4]
  assign buffer_4_611 = $signed(_T_69368); // @[Modules.scala 53:83:@17895.4]
  assign _T_69370 = $signed(buffer_2_440) + $signed(buffer_4_441); // @[Modules.scala 53:83:@17897.4]
  assign _T_69371 = _T_69370[10:0]; // @[Modules.scala 53:83:@17898.4]
  assign buffer_4_612 = $signed(_T_69371); // @[Modules.scala 53:83:@17899.4]
  assign _T_69373 = $signed(buffer_4_442) + $signed(buffer_4_443); // @[Modules.scala 53:83:@17901.4]
  assign _T_69374 = _T_69373[10:0]; // @[Modules.scala 53:83:@17902.4]
  assign buffer_4_613 = $signed(_T_69374); // @[Modules.scala 53:83:@17903.4]
  assign _T_69376 = $signed(buffer_4_444) + $signed(buffer_4_445); // @[Modules.scala 53:83:@17905.4]
  assign _T_69377 = _T_69376[10:0]; // @[Modules.scala 53:83:@17906.4]
  assign buffer_4_614 = $signed(_T_69377); // @[Modules.scala 53:83:@17907.4]
  assign _T_69382 = $signed(buffer_1_448) + $signed(buffer_4_449); // @[Modules.scala 53:83:@17913.4]
  assign _T_69383 = _T_69382[10:0]; // @[Modules.scala 53:83:@17914.4]
  assign buffer_4_616 = $signed(_T_69383); // @[Modules.scala 53:83:@17915.4]
  assign _T_69385 = $signed(buffer_4_450) + $signed(buffer_1_451); // @[Modules.scala 53:83:@17917.4]
  assign _T_69386 = _T_69385[10:0]; // @[Modules.scala 53:83:@17918.4]
  assign buffer_4_617 = $signed(_T_69386); // @[Modules.scala 53:83:@17919.4]
  assign _T_69388 = $signed(buffer_4_452) + $signed(buffer_4_453); // @[Modules.scala 53:83:@17921.4]
  assign _T_69389 = _T_69388[10:0]; // @[Modules.scala 53:83:@17922.4]
  assign buffer_4_618 = $signed(_T_69389); // @[Modules.scala 53:83:@17923.4]
  assign _T_69394 = $signed(buffer_4_456) + $signed(buffer_4_457); // @[Modules.scala 53:83:@17929.4]
  assign _T_69395 = _T_69394[10:0]; // @[Modules.scala 53:83:@17930.4]
  assign buffer_4_620 = $signed(_T_69395); // @[Modules.scala 53:83:@17931.4]
  assign _T_69403 = $signed(buffer_4_462) + $signed(buffer_4_463); // @[Modules.scala 53:83:@17941.4]
  assign _T_69404 = _T_69403[10:0]; // @[Modules.scala 53:83:@17942.4]
  assign buffer_4_623 = $signed(_T_69404); // @[Modules.scala 53:83:@17943.4]
  assign _T_69409 = $signed(buffer_4_466) + $signed(buffer_4_467); // @[Modules.scala 53:83:@17949.4]
  assign _T_69410 = _T_69409[10:0]; // @[Modules.scala 53:83:@17950.4]
  assign buffer_4_625 = $signed(_T_69410); // @[Modules.scala 53:83:@17951.4]
  assign _T_69412 = $signed(buffer_1_468) + $signed(buffer_4_469); // @[Modules.scala 53:83:@17953.4]
  assign _T_69413 = _T_69412[10:0]; // @[Modules.scala 53:83:@17954.4]
  assign buffer_4_626 = $signed(_T_69413); // @[Modules.scala 53:83:@17955.4]
  assign _T_69415 = $signed(buffer_3_470) + $signed(buffer_1_471); // @[Modules.scala 53:83:@17957.4]
  assign _T_69416 = _T_69415[10:0]; // @[Modules.scala 53:83:@17958.4]
  assign buffer_4_627 = $signed(_T_69416); // @[Modules.scala 53:83:@17959.4]
  assign _T_69418 = $signed(buffer_4_472) + $signed(buffer_1_473); // @[Modules.scala 53:83:@17961.4]
  assign _T_69419 = _T_69418[10:0]; // @[Modules.scala 53:83:@17962.4]
  assign buffer_4_628 = $signed(_T_69419); // @[Modules.scala 53:83:@17963.4]
  assign _T_69421 = $signed(buffer_1_474) + $signed(buffer_4_475); // @[Modules.scala 53:83:@17965.4]
  assign _T_69422 = _T_69421[10:0]; // @[Modules.scala 53:83:@17966.4]
  assign buffer_4_629 = $signed(_T_69422); // @[Modules.scala 53:83:@17967.4]
  assign _T_69424 = $signed(buffer_0_476) + $signed(buffer_3_477); // @[Modules.scala 53:83:@17969.4]
  assign _T_69425 = _T_69424[10:0]; // @[Modules.scala 53:83:@17970.4]
  assign buffer_4_630 = $signed(_T_69425); // @[Modules.scala 53:83:@17971.4]
  assign _T_69427 = $signed(buffer_4_478) + $signed(buffer_1_479); // @[Modules.scala 53:83:@17973.4]
  assign _T_69428 = _T_69427[10:0]; // @[Modules.scala 53:83:@17974.4]
  assign buffer_4_631 = $signed(_T_69428); // @[Modules.scala 53:83:@17975.4]
  assign _T_69430 = $signed(buffer_4_480) + $signed(buffer_1_481); // @[Modules.scala 53:83:@17977.4]
  assign _T_69431 = _T_69430[10:0]; // @[Modules.scala 53:83:@17978.4]
  assign buffer_4_632 = $signed(_T_69431); // @[Modules.scala 53:83:@17979.4]
  assign _T_69433 = $signed(buffer_4_482) + $signed(buffer_4_483); // @[Modules.scala 53:83:@17981.4]
  assign _T_69434 = _T_69433[10:0]; // @[Modules.scala 53:83:@17982.4]
  assign buffer_4_633 = $signed(_T_69434); // @[Modules.scala 53:83:@17983.4]
  assign _T_69436 = $signed(buffer_4_484) + $signed(buffer_0_485); // @[Modules.scala 53:83:@17985.4]
  assign _T_69437 = _T_69436[10:0]; // @[Modules.scala 53:83:@17986.4]
  assign buffer_4_634 = $signed(_T_69437); // @[Modules.scala 53:83:@17987.4]
  assign _T_69439 = $signed(buffer_1_486) + $signed(buffer_4_487); // @[Modules.scala 53:83:@17989.4]
  assign _T_69440 = _T_69439[10:0]; // @[Modules.scala 53:83:@17990.4]
  assign buffer_4_635 = $signed(_T_69440); // @[Modules.scala 53:83:@17991.4]
  assign _T_69442 = $signed(buffer_4_488) + $signed(buffer_4_489); // @[Modules.scala 53:83:@17993.4]
  assign _T_69443 = _T_69442[10:0]; // @[Modules.scala 53:83:@17994.4]
  assign buffer_4_636 = $signed(_T_69443); // @[Modules.scala 53:83:@17995.4]
  assign _T_69445 = $signed(buffer_4_490) + $signed(buffer_4_491); // @[Modules.scala 53:83:@17997.4]
  assign _T_69446 = _T_69445[10:0]; // @[Modules.scala 53:83:@17998.4]
  assign buffer_4_637 = $signed(_T_69446); // @[Modules.scala 53:83:@17999.4]
  assign _T_69448 = $signed(buffer_4_492) + $signed(buffer_4_493); // @[Modules.scala 53:83:@18001.4]
  assign _T_69449 = _T_69448[10:0]; // @[Modules.scala 53:83:@18002.4]
  assign buffer_4_638 = $signed(_T_69449); // @[Modules.scala 53:83:@18003.4]
  assign _T_69451 = $signed(buffer_4_494) + $signed(buffer_4_495); // @[Modules.scala 53:83:@18005.4]
  assign _T_69452 = _T_69451[10:0]; // @[Modules.scala 53:83:@18006.4]
  assign buffer_4_639 = $signed(_T_69452); // @[Modules.scala 53:83:@18007.4]
  assign _T_69454 = $signed(buffer_4_496) + $signed(buffer_4_497); // @[Modules.scala 53:83:@18009.4]
  assign _T_69455 = _T_69454[10:0]; // @[Modules.scala 53:83:@18010.4]
  assign buffer_4_640 = $signed(_T_69455); // @[Modules.scala 53:83:@18011.4]
  assign _T_69457 = $signed(buffer_3_498) + $signed(buffer_0_499); // @[Modules.scala 53:83:@18013.4]
  assign _T_69458 = _T_69457[10:0]; // @[Modules.scala 53:83:@18014.4]
  assign buffer_4_641 = $signed(_T_69458); // @[Modules.scala 53:83:@18015.4]
  assign _T_69460 = $signed(buffer_4_500) + $signed(buffer_4_501); // @[Modules.scala 53:83:@18017.4]
  assign _T_69461 = _T_69460[10:0]; // @[Modules.scala 53:83:@18018.4]
  assign buffer_4_642 = $signed(_T_69461); // @[Modules.scala 53:83:@18019.4]
  assign _T_69463 = $signed(buffer_4_502) + $signed(buffer_3_503); // @[Modules.scala 53:83:@18021.4]
  assign _T_69464 = _T_69463[10:0]; // @[Modules.scala 53:83:@18022.4]
  assign buffer_4_643 = $signed(_T_69464); // @[Modules.scala 53:83:@18023.4]
  assign _T_69466 = $signed(buffer_1_504) + $signed(buffer_4_505); // @[Modules.scala 53:83:@18025.4]
  assign _T_69467 = _T_69466[10:0]; // @[Modules.scala 53:83:@18026.4]
  assign buffer_4_644 = $signed(_T_69467); // @[Modules.scala 53:83:@18027.4]
  assign _T_69469 = $signed(buffer_1_506) + $signed(buffer_4_507); // @[Modules.scala 53:83:@18029.4]
  assign _T_69470 = _T_69469[10:0]; // @[Modules.scala 53:83:@18030.4]
  assign buffer_4_645 = $signed(_T_69470); // @[Modules.scala 53:83:@18031.4]
  assign _T_69472 = $signed(buffer_4_508) + $signed(buffer_1_509); // @[Modules.scala 53:83:@18033.4]
  assign _T_69473 = _T_69472[10:0]; // @[Modules.scala 53:83:@18034.4]
  assign buffer_4_646 = $signed(_T_69473); // @[Modules.scala 53:83:@18035.4]
  assign _T_69475 = $signed(buffer_3_510) + $signed(buffer_4_511); // @[Modules.scala 53:83:@18037.4]
  assign _T_69476 = _T_69475[10:0]; // @[Modules.scala 53:83:@18038.4]
  assign buffer_4_647 = $signed(_T_69476); // @[Modules.scala 53:83:@18039.4]
  assign _T_69478 = $signed(buffer_4_512) + $signed(buffer_4_513); // @[Modules.scala 53:83:@18041.4]
  assign _T_69479 = _T_69478[10:0]; // @[Modules.scala 53:83:@18042.4]
  assign buffer_4_648 = $signed(_T_69479); // @[Modules.scala 53:83:@18043.4]
  assign _T_69481 = $signed(buffer_1_514) + $signed(buffer_4_515); // @[Modules.scala 53:83:@18045.4]
  assign _T_69482 = _T_69481[10:0]; // @[Modules.scala 53:83:@18046.4]
  assign buffer_4_649 = $signed(_T_69482); // @[Modules.scala 53:83:@18047.4]
  assign _T_69487 = $signed(buffer_4_518) + $signed(buffer_3_519); // @[Modules.scala 53:83:@18053.4]
  assign _T_69488 = _T_69487[10:0]; // @[Modules.scala 53:83:@18054.4]
  assign buffer_4_651 = $signed(_T_69488); // @[Modules.scala 53:83:@18055.4]
  assign _T_69490 = $signed(buffer_4_520) + $signed(buffer_4_521); // @[Modules.scala 53:83:@18057.4]
  assign _T_69491 = _T_69490[10:0]; // @[Modules.scala 53:83:@18058.4]
  assign buffer_4_652 = $signed(_T_69491); // @[Modules.scala 53:83:@18059.4]
  assign _T_69493 = $signed(buffer_4_522) + $signed(buffer_4_523); // @[Modules.scala 53:83:@18061.4]
  assign _T_69494 = _T_69493[10:0]; // @[Modules.scala 53:83:@18062.4]
  assign buffer_4_653 = $signed(_T_69494); // @[Modules.scala 53:83:@18063.4]
  assign _T_69496 = $signed(buffer_0_524) + $signed(buffer_4_525); // @[Modules.scala 53:83:@18065.4]
  assign _T_69497 = _T_69496[10:0]; // @[Modules.scala 53:83:@18066.4]
  assign buffer_4_654 = $signed(_T_69497); // @[Modules.scala 53:83:@18067.4]
  assign _T_69502 = $signed(buffer_4_528) + $signed(buffer_1_529); // @[Modules.scala 53:83:@18073.4]
  assign _T_69503 = _T_69502[10:0]; // @[Modules.scala 53:83:@18074.4]
  assign buffer_4_656 = $signed(_T_69503); // @[Modules.scala 53:83:@18075.4]
  assign _T_69505 = $signed(buffer_3_530) + $signed(buffer_4_531); // @[Modules.scala 53:83:@18077.4]
  assign _T_69506 = _T_69505[10:0]; // @[Modules.scala 53:83:@18078.4]
  assign buffer_4_657 = $signed(_T_69506); // @[Modules.scala 53:83:@18079.4]
  assign _T_69508 = $signed(buffer_1_532) + $signed(buffer_3_533); // @[Modules.scala 53:83:@18081.4]
  assign _T_69509 = _T_69508[10:0]; // @[Modules.scala 53:83:@18082.4]
  assign buffer_4_658 = $signed(_T_69509); // @[Modules.scala 53:83:@18083.4]
  assign _T_69511 = $signed(buffer_1_534) + $signed(buffer_4_535); // @[Modules.scala 53:83:@18085.4]
  assign _T_69512 = _T_69511[10:0]; // @[Modules.scala 53:83:@18086.4]
  assign buffer_4_659 = $signed(_T_69512); // @[Modules.scala 53:83:@18087.4]
  assign _T_69514 = $signed(buffer_2_536) + $signed(buffer_4_537); // @[Modules.scala 53:83:@18089.4]
  assign _T_69515 = _T_69514[10:0]; // @[Modules.scala 53:83:@18090.4]
  assign buffer_4_660 = $signed(_T_69515); // @[Modules.scala 53:83:@18091.4]
  assign _T_69517 = $signed(buffer_4_538) + $signed(buffer_4_539); // @[Modules.scala 53:83:@18093.4]
  assign _T_69518 = _T_69517[10:0]; // @[Modules.scala 53:83:@18094.4]
  assign buffer_4_661 = $signed(_T_69518); // @[Modules.scala 53:83:@18095.4]
  assign _T_69520 = $signed(buffer_3_540) + $signed(buffer_4_541); // @[Modules.scala 53:83:@18097.4]
  assign _T_69521 = _T_69520[10:0]; // @[Modules.scala 53:83:@18098.4]
  assign buffer_4_662 = $signed(_T_69521); // @[Modules.scala 53:83:@18099.4]
  assign _T_69526 = $signed(buffer_4_544) + $signed(buffer_4_545); // @[Modules.scala 53:83:@18105.4]
  assign _T_69527 = _T_69526[10:0]; // @[Modules.scala 53:83:@18106.4]
  assign buffer_4_664 = $signed(_T_69527); // @[Modules.scala 53:83:@18107.4]
  assign _T_69529 = $signed(buffer_0_546) + $signed(buffer_4_547); // @[Modules.scala 53:83:@18109.4]
  assign _T_69530 = _T_69529[10:0]; // @[Modules.scala 53:83:@18110.4]
  assign buffer_4_665 = $signed(_T_69530); // @[Modules.scala 53:83:@18111.4]
  assign _T_69532 = $signed(buffer_4_548) + $signed(buffer_1_549); // @[Modules.scala 53:83:@18113.4]
  assign _T_69533 = _T_69532[10:0]; // @[Modules.scala 53:83:@18114.4]
  assign buffer_4_666 = $signed(_T_69533); // @[Modules.scala 53:83:@18115.4]
  assign _T_69535 = $signed(buffer_4_550) + $signed(buffer_3_551); // @[Modules.scala 53:83:@18117.4]
  assign _T_69536 = _T_69535[10:0]; // @[Modules.scala 53:83:@18118.4]
  assign buffer_4_667 = $signed(_T_69536); // @[Modules.scala 53:83:@18119.4]
  assign _T_69538 = $signed(buffer_4_552) + $signed(buffer_0_553); // @[Modules.scala 53:83:@18121.4]
  assign _T_69539 = _T_69538[10:0]; // @[Modules.scala 53:83:@18122.4]
  assign buffer_4_668 = $signed(_T_69539); // @[Modules.scala 53:83:@18123.4]
  assign _T_69541 = $signed(buffer_4_554) + $signed(buffer_1_555); // @[Modules.scala 53:83:@18125.4]
  assign _T_69542 = _T_69541[10:0]; // @[Modules.scala 53:83:@18126.4]
  assign buffer_4_669 = $signed(_T_69542); // @[Modules.scala 53:83:@18127.4]
  assign _T_69544 = $signed(buffer_1_556) + $signed(buffer_4_557); // @[Modules.scala 53:83:@18129.4]
  assign _T_69545 = _T_69544[10:0]; // @[Modules.scala 53:83:@18130.4]
  assign buffer_4_670 = $signed(_T_69545); // @[Modules.scala 53:83:@18131.4]
  assign _T_69547 = $signed(buffer_4_558) + $signed(buffer_4_559); // @[Modules.scala 53:83:@18133.4]
  assign _T_69548 = _T_69547[10:0]; // @[Modules.scala 53:83:@18134.4]
  assign buffer_4_671 = $signed(_T_69548); // @[Modules.scala 53:83:@18135.4]
  assign _T_69550 = $signed(buffer_4_560) + $signed(buffer_4_561); // @[Modules.scala 53:83:@18137.4]
  assign _T_69551 = _T_69550[10:0]; // @[Modules.scala 53:83:@18138.4]
  assign buffer_4_672 = $signed(_T_69551); // @[Modules.scala 53:83:@18139.4]
  assign _T_69553 = $signed(buffer_3_562) + $signed(buffer_4_563); // @[Modules.scala 53:83:@18141.4]
  assign _T_69554 = _T_69553[10:0]; // @[Modules.scala 53:83:@18142.4]
  assign buffer_4_673 = $signed(_T_69554); // @[Modules.scala 53:83:@18143.4]
  assign _T_69556 = $signed(buffer_4_564) + $signed(buffer_3_565); // @[Modules.scala 53:83:@18145.4]
  assign _T_69557 = _T_69556[10:0]; // @[Modules.scala 53:83:@18146.4]
  assign buffer_4_674 = $signed(_T_69557); // @[Modules.scala 53:83:@18147.4]
  assign _T_69559 = $signed(buffer_4_566) + $signed(buffer_1_567); // @[Modules.scala 53:83:@18149.4]
  assign _T_69560 = _T_69559[10:0]; // @[Modules.scala 53:83:@18150.4]
  assign buffer_4_675 = $signed(_T_69560); // @[Modules.scala 53:83:@18151.4]
  assign _T_69562 = $signed(buffer_4_568) + $signed(buffer_2_569); // @[Modules.scala 53:83:@18153.4]
  assign _T_69563 = _T_69562[10:0]; // @[Modules.scala 53:83:@18154.4]
  assign buffer_4_676 = $signed(_T_69563); // @[Modules.scala 53:83:@18155.4]
  assign _T_69568 = $signed(buffer_3_572) + $signed(buffer_4_573); // @[Modules.scala 53:83:@18161.4]
  assign _T_69569 = _T_69568[10:0]; // @[Modules.scala 53:83:@18162.4]
  assign buffer_4_678 = $signed(_T_69569); // @[Modules.scala 53:83:@18163.4]
  assign _T_69571 = $signed(buffer_3_574) + $signed(buffer_2_575); // @[Modules.scala 53:83:@18165.4]
  assign _T_69572 = _T_69571[10:0]; // @[Modules.scala 53:83:@18166.4]
  assign buffer_4_679 = $signed(_T_69572); // @[Modules.scala 53:83:@18167.4]
  assign _T_69577 = $signed(buffer_0_578) + $signed(buffer_4_579); // @[Modules.scala 53:83:@18173.4]
  assign _T_69578 = _T_69577[10:0]; // @[Modules.scala 53:83:@18174.4]
  assign buffer_4_681 = $signed(_T_69578); // @[Modules.scala 53:83:@18175.4]
  assign _T_69580 = $signed(buffer_4_580) + $signed(buffer_4_581); // @[Modules.scala 53:83:@18177.4]
  assign _T_69581 = _T_69580[10:0]; // @[Modules.scala 53:83:@18178.4]
  assign buffer_4_682 = $signed(_T_69581); // @[Modules.scala 53:83:@18179.4]
  assign _T_69583 = $signed(buffer_4_582) + $signed(buffer_4_583); // @[Modules.scala 53:83:@18181.4]
  assign _T_69584 = _T_69583[10:0]; // @[Modules.scala 53:83:@18182.4]
  assign buffer_4_683 = $signed(_T_69584); // @[Modules.scala 53:83:@18183.4]
  assign _T_69586 = $signed(buffer_4_584) + $signed(buffer_4_585); // @[Modules.scala 53:83:@18185.4]
  assign _T_69587 = _T_69586[10:0]; // @[Modules.scala 53:83:@18186.4]
  assign buffer_4_684 = $signed(_T_69587); // @[Modules.scala 53:83:@18187.4]
  assign _T_69589 = $signed(buffer_1_586) + $signed(buffer_4_587); // @[Modules.scala 53:83:@18189.4]
  assign _T_69590 = _T_69589[10:0]; // @[Modules.scala 53:83:@18190.4]
  assign buffer_4_685 = $signed(_T_69590); // @[Modules.scala 53:83:@18191.4]
  assign _T_69592 = $signed(buffer_4_588) + $signed(buffer_4_589); // @[Modules.scala 56:109:@18193.4]
  assign _T_69593 = _T_69592[10:0]; // @[Modules.scala 56:109:@18194.4]
  assign buffer_4_686 = $signed(_T_69593); // @[Modules.scala 56:109:@18195.4]
  assign _T_69595 = $signed(buffer_4_590) + $signed(buffer_4_591); // @[Modules.scala 56:109:@18197.4]
  assign _T_69596 = _T_69595[10:0]; // @[Modules.scala 56:109:@18198.4]
  assign buffer_4_687 = $signed(_T_69596); // @[Modules.scala 56:109:@18199.4]
  assign _T_69598 = $signed(buffer_4_592) + $signed(buffer_4_593); // @[Modules.scala 56:109:@18201.4]
  assign _T_69599 = _T_69598[10:0]; // @[Modules.scala 56:109:@18202.4]
  assign buffer_4_688 = $signed(_T_69599); // @[Modules.scala 56:109:@18203.4]
  assign _T_69601 = $signed(buffer_4_594) + $signed(buffer_4_595); // @[Modules.scala 56:109:@18205.4]
  assign _T_69602 = _T_69601[10:0]; // @[Modules.scala 56:109:@18206.4]
  assign buffer_4_689 = $signed(_T_69602); // @[Modules.scala 56:109:@18207.4]
  assign _T_69607 = $signed(buffer_4_598) + $signed(buffer_4_599); // @[Modules.scala 56:109:@18213.4]
  assign _T_69608 = _T_69607[10:0]; // @[Modules.scala 56:109:@18214.4]
  assign buffer_4_691 = $signed(_T_69608); // @[Modules.scala 56:109:@18215.4]
  assign _T_69613 = $signed(buffer_4_602) + $signed(buffer_4_603); // @[Modules.scala 56:109:@18221.4]
  assign _T_69614 = _T_69613[10:0]; // @[Modules.scala 56:109:@18222.4]
  assign buffer_4_693 = $signed(_T_69614); // @[Modules.scala 56:109:@18223.4]
  assign _T_69616 = $signed(buffer_4_604) + $signed(buffer_4_605); // @[Modules.scala 56:109:@18225.4]
  assign _T_69617 = _T_69616[10:0]; // @[Modules.scala 56:109:@18226.4]
  assign buffer_4_694 = $signed(_T_69617); // @[Modules.scala 56:109:@18227.4]
  assign _T_69619 = $signed(buffer_4_606) + $signed(buffer_4_607); // @[Modules.scala 56:109:@18229.4]
  assign _T_69620 = _T_69619[10:0]; // @[Modules.scala 56:109:@18230.4]
  assign buffer_4_695 = $signed(_T_69620); // @[Modules.scala 56:109:@18231.4]
  assign _T_69622 = $signed(buffer_4_608) + $signed(buffer_4_609); // @[Modules.scala 56:109:@18233.4]
  assign _T_69623 = _T_69622[10:0]; // @[Modules.scala 56:109:@18234.4]
  assign buffer_4_696 = $signed(_T_69623); // @[Modules.scala 56:109:@18235.4]
  assign _T_69625 = $signed(buffer_4_610) + $signed(buffer_4_611); // @[Modules.scala 56:109:@18237.4]
  assign _T_69626 = _T_69625[10:0]; // @[Modules.scala 56:109:@18238.4]
  assign buffer_4_697 = $signed(_T_69626); // @[Modules.scala 56:109:@18239.4]
  assign _T_69628 = $signed(buffer_4_612) + $signed(buffer_4_613); // @[Modules.scala 56:109:@18241.4]
  assign _T_69629 = _T_69628[10:0]; // @[Modules.scala 56:109:@18242.4]
  assign buffer_4_698 = $signed(_T_69629); // @[Modules.scala 56:109:@18243.4]
  assign _T_69631 = $signed(buffer_4_614) + $signed(buffer_2_615); // @[Modules.scala 56:109:@18245.4]
  assign _T_69632 = _T_69631[10:0]; // @[Modules.scala 56:109:@18246.4]
  assign buffer_4_699 = $signed(_T_69632); // @[Modules.scala 56:109:@18247.4]
  assign _T_69634 = $signed(buffer_4_616) + $signed(buffer_4_617); // @[Modules.scala 56:109:@18249.4]
  assign _T_69635 = _T_69634[10:0]; // @[Modules.scala 56:109:@18250.4]
  assign buffer_4_700 = $signed(_T_69635); // @[Modules.scala 56:109:@18251.4]
  assign _T_69637 = $signed(buffer_4_618) + $signed(buffer_2_619); // @[Modules.scala 56:109:@18253.4]
  assign _T_69638 = _T_69637[10:0]; // @[Modules.scala 56:109:@18254.4]
  assign buffer_4_701 = $signed(_T_69638); // @[Modules.scala 56:109:@18255.4]
  assign _T_69640 = $signed(buffer_4_620) + $signed(buffer_0_621); // @[Modules.scala 56:109:@18257.4]
  assign _T_69641 = _T_69640[10:0]; // @[Modules.scala 56:109:@18258.4]
  assign buffer_4_702 = $signed(_T_69641); // @[Modules.scala 56:109:@18259.4]
  assign _T_69643 = $signed(buffer_3_622) + $signed(buffer_4_623); // @[Modules.scala 56:109:@18261.4]
  assign _T_69644 = _T_69643[10:0]; // @[Modules.scala 56:109:@18262.4]
  assign buffer_4_703 = $signed(_T_69644); // @[Modules.scala 56:109:@18263.4]
  assign _T_69646 = $signed(buffer_0_624) + $signed(buffer_4_625); // @[Modules.scala 56:109:@18265.4]
  assign _T_69647 = _T_69646[10:0]; // @[Modules.scala 56:109:@18266.4]
  assign buffer_4_704 = $signed(_T_69647); // @[Modules.scala 56:109:@18267.4]
  assign _T_69649 = $signed(buffer_4_626) + $signed(buffer_4_627); // @[Modules.scala 56:109:@18269.4]
  assign _T_69650 = _T_69649[10:0]; // @[Modules.scala 56:109:@18270.4]
  assign buffer_4_705 = $signed(_T_69650); // @[Modules.scala 56:109:@18271.4]
  assign _T_69652 = $signed(buffer_4_628) + $signed(buffer_4_629); // @[Modules.scala 56:109:@18273.4]
  assign _T_69653 = _T_69652[10:0]; // @[Modules.scala 56:109:@18274.4]
  assign buffer_4_706 = $signed(_T_69653); // @[Modules.scala 56:109:@18275.4]
  assign _T_69655 = $signed(buffer_4_630) + $signed(buffer_4_631); // @[Modules.scala 56:109:@18277.4]
  assign _T_69656 = _T_69655[10:0]; // @[Modules.scala 56:109:@18278.4]
  assign buffer_4_707 = $signed(_T_69656); // @[Modules.scala 56:109:@18279.4]
  assign _T_69658 = $signed(buffer_4_632) + $signed(buffer_4_633); // @[Modules.scala 56:109:@18281.4]
  assign _T_69659 = _T_69658[10:0]; // @[Modules.scala 56:109:@18282.4]
  assign buffer_4_708 = $signed(_T_69659); // @[Modules.scala 56:109:@18283.4]
  assign _T_69661 = $signed(buffer_4_634) + $signed(buffer_4_635); // @[Modules.scala 56:109:@18285.4]
  assign _T_69662 = _T_69661[10:0]; // @[Modules.scala 56:109:@18286.4]
  assign buffer_4_709 = $signed(_T_69662); // @[Modules.scala 56:109:@18287.4]
  assign _T_69664 = $signed(buffer_4_636) + $signed(buffer_4_637); // @[Modules.scala 56:109:@18289.4]
  assign _T_69665 = _T_69664[10:0]; // @[Modules.scala 56:109:@18290.4]
  assign buffer_4_710 = $signed(_T_69665); // @[Modules.scala 56:109:@18291.4]
  assign _T_69667 = $signed(buffer_4_638) + $signed(buffer_4_639); // @[Modules.scala 56:109:@18293.4]
  assign _T_69668 = _T_69667[10:0]; // @[Modules.scala 56:109:@18294.4]
  assign buffer_4_711 = $signed(_T_69668); // @[Modules.scala 56:109:@18295.4]
  assign _T_69670 = $signed(buffer_4_640) + $signed(buffer_4_641); // @[Modules.scala 56:109:@18297.4]
  assign _T_69671 = _T_69670[10:0]; // @[Modules.scala 56:109:@18298.4]
  assign buffer_4_712 = $signed(_T_69671); // @[Modules.scala 56:109:@18299.4]
  assign _T_69673 = $signed(buffer_4_642) + $signed(buffer_4_643); // @[Modules.scala 56:109:@18301.4]
  assign _T_69674 = _T_69673[10:0]; // @[Modules.scala 56:109:@18302.4]
  assign buffer_4_713 = $signed(_T_69674); // @[Modules.scala 56:109:@18303.4]
  assign _T_69676 = $signed(buffer_4_644) + $signed(buffer_4_645); // @[Modules.scala 56:109:@18305.4]
  assign _T_69677 = _T_69676[10:0]; // @[Modules.scala 56:109:@18306.4]
  assign buffer_4_714 = $signed(_T_69677); // @[Modules.scala 56:109:@18307.4]
  assign _T_69679 = $signed(buffer_4_646) + $signed(buffer_4_647); // @[Modules.scala 56:109:@18309.4]
  assign _T_69680 = _T_69679[10:0]; // @[Modules.scala 56:109:@18310.4]
  assign buffer_4_715 = $signed(_T_69680); // @[Modules.scala 56:109:@18311.4]
  assign _T_69682 = $signed(buffer_4_648) + $signed(buffer_4_649); // @[Modules.scala 56:109:@18313.4]
  assign _T_69683 = _T_69682[10:0]; // @[Modules.scala 56:109:@18314.4]
  assign buffer_4_716 = $signed(_T_69683); // @[Modules.scala 56:109:@18315.4]
  assign _T_69685 = $signed(buffer_3_650) + $signed(buffer_4_651); // @[Modules.scala 56:109:@18317.4]
  assign _T_69686 = _T_69685[10:0]; // @[Modules.scala 56:109:@18318.4]
  assign buffer_4_717 = $signed(_T_69686); // @[Modules.scala 56:109:@18319.4]
  assign _T_69688 = $signed(buffer_4_652) + $signed(buffer_4_653); // @[Modules.scala 56:109:@18321.4]
  assign _T_69689 = _T_69688[10:0]; // @[Modules.scala 56:109:@18322.4]
  assign buffer_4_718 = $signed(_T_69689); // @[Modules.scala 56:109:@18323.4]
  assign _T_69691 = $signed(buffer_4_654) + $signed(buffer_1_655); // @[Modules.scala 56:109:@18325.4]
  assign _T_69692 = _T_69691[10:0]; // @[Modules.scala 56:109:@18326.4]
  assign buffer_4_719 = $signed(_T_69692); // @[Modules.scala 56:109:@18327.4]
  assign _T_69694 = $signed(buffer_4_656) + $signed(buffer_4_657); // @[Modules.scala 56:109:@18329.4]
  assign _T_69695 = _T_69694[10:0]; // @[Modules.scala 56:109:@18330.4]
  assign buffer_4_720 = $signed(_T_69695); // @[Modules.scala 56:109:@18331.4]
  assign _T_69697 = $signed(buffer_4_658) + $signed(buffer_4_659); // @[Modules.scala 56:109:@18333.4]
  assign _T_69698 = _T_69697[10:0]; // @[Modules.scala 56:109:@18334.4]
  assign buffer_4_721 = $signed(_T_69698); // @[Modules.scala 56:109:@18335.4]
  assign _T_69700 = $signed(buffer_4_660) + $signed(buffer_4_661); // @[Modules.scala 56:109:@18337.4]
  assign _T_69701 = _T_69700[10:0]; // @[Modules.scala 56:109:@18338.4]
  assign buffer_4_722 = $signed(_T_69701); // @[Modules.scala 56:109:@18339.4]
  assign _T_69703 = $signed(buffer_4_662) + $signed(buffer_0_663); // @[Modules.scala 56:109:@18341.4]
  assign _T_69704 = _T_69703[10:0]; // @[Modules.scala 56:109:@18342.4]
  assign buffer_4_723 = $signed(_T_69704); // @[Modules.scala 56:109:@18343.4]
  assign _T_69706 = $signed(buffer_4_664) + $signed(buffer_4_665); // @[Modules.scala 56:109:@18345.4]
  assign _T_69707 = _T_69706[10:0]; // @[Modules.scala 56:109:@18346.4]
  assign buffer_4_724 = $signed(_T_69707); // @[Modules.scala 56:109:@18347.4]
  assign _T_69709 = $signed(buffer_4_666) + $signed(buffer_4_667); // @[Modules.scala 56:109:@18349.4]
  assign _T_69710 = _T_69709[10:0]; // @[Modules.scala 56:109:@18350.4]
  assign buffer_4_725 = $signed(_T_69710); // @[Modules.scala 56:109:@18351.4]
  assign _T_69712 = $signed(buffer_4_668) + $signed(buffer_4_669); // @[Modules.scala 56:109:@18353.4]
  assign _T_69713 = _T_69712[10:0]; // @[Modules.scala 56:109:@18354.4]
  assign buffer_4_726 = $signed(_T_69713); // @[Modules.scala 56:109:@18355.4]
  assign _T_69715 = $signed(buffer_4_670) + $signed(buffer_4_671); // @[Modules.scala 56:109:@18357.4]
  assign _T_69716 = _T_69715[10:0]; // @[Modules.scala 56:109:@18358.4]
  assign buffer_4_727 = $signed(_T_69716); // @[Modules.scala 56:109:@18359.4]
  assign _T_69718 = $signed(buffer_4_672) + $signed(buffer_4_673); // @[Modules.scala 56:109:@18361.4]
  assign _T_69719 = _T_69718[10:0]; // @[Modules.scala 56:109:@18362.4]
  assign buffer_4_728 = $signed(_T_69719); // @[Modules.scala 56:109:@18363.4]
  assign _T_69721 = $signed(buffer_4_674) + $signed(buffer_4_675); // @[Modules.scala 56:109:@18365.4]
  assign _T_69722 = _T_69721[10:0]; // @[Modules.scala 56:109:@18366.4]
  assign buffer_4_729 = $signed(_T_69722); // @[Modules.scala 56:109:@18367.4]
  assign _T_69724 = $signed(buffer_4_676) + $signed(buffer_2_677); // @[Modules.scala 56:109:@18369.4]
  assign _T_69725 = _T_69724[10:0]; // @[Modules.scala 56:109:@18370.4]
  assign buffer_4_730 = $signed(_T_69725); // @[Modules.scala 56:109:@18371.4]
  assign _T_69727 = $signed(buffer_4_678) + $signed(buffer_4_679); // @[Modules.scala 56:109:@18373.4]
  assign _T_69728 = _T_69727[10:0]; // @[Modules.scala 56:109:@18374.4]
  assign buffer_4_731 = $signed(_T_69728); // @[Modules.scala 56:109:@18375.4]
  assign _T_69730 = $signed(buffer_1_680) + $signed(buffer_4_681); // @[Modules.scala 56:109:@18377.4]
  assign _T_69731 = _T_69730[10:0]; // @[Modules.scala 56:109:@18378.4]
  assign buffer_4_732 = $signed(_T_69731); // @[Modules.scala 56:109:@18379.4]
  assign _T_69733 = $signed(buffer_4_682) + $signed(buffer_4_683); // @[Modules.scala 56:109:@18381.4]
  assign _T_69734 = _T_69733[10:0]; // @[Modules.scala 56:109:@18382.4]
  assign buffer_4_733 = $signed(_T_69734); // @[Modules.scala 56:109:@18383.4]
  assign _T_69736 = $signed(buffer_4_684) + $signed(buffer_4_685); // @[Modules.scala 56:109:@18385.4]
  assign _T_69737 = _T_69736[10:0]; // @[Modules.scala 56:109:@18386.4]
  assign buffer_4_734 = $signed(_T_69737); // @[Modules.scala 56:109:@18387.4]
  assign _T_69739 = $signed(buffer_4_686) + $signed(buffer_4_687); // @[Modules.scala 63:156:@18390.4]
  assign _T_69740 = _T_69739[10:0]; // @[Modules.scala 63:156:@18391.4]
  assign buffer_4_736 = $signed(_T_69740); // @[Modules.scala 63:156:@18392.4]
  assign _T_69742 = $signed(buffer_4_736) + $signed(buffer_4_688); // @[Modules.scala 63:156:@18394.4]
  assign _T_69743 = _T_69742[10:0]; // @[Modules.scala 63:156:@18395.4]
  assign buffer_4_737 = $signed(_T_69743); // @[Modules.scala 63:156:@18396.4]
  assign _T_69745 = $signed(buffer_4_737) + $signed(buffer_4_689); // @[Modules.scala 63:156:@18398.4]
  assign _T_69746 = _T_69745[10:0]; // @[Modules.scala 63:156:@18399.4]
  assign buffer_4_738 = $signed(_T_69746); // @[Modules.scala 63:156:@18400.4]
  assign _T_69748 = $signed(buffer_4_738) + $signed(buffer_1_690); // @[Modules.scala 63:156:@18402.4]
  assign _T_69749 = _T_69748[10:0]; // @[Modules.scala 63:156:@18403.4]
  assign buffer_4_739 = $signed(_T_69749); // @[Modules.scala 63:156:@18404.4]
  assign _T_69751 = $signed(buffer_4_739) + $signed(buffer_4_691); // @[Modules.scala 63:156:@18406.4]
  assign _T_69752 = _T_69751[10:0]; // @[Modules.scala 63:156:@18407.4]
  assign buffer_4_740 = $signed(_T_69752); // @[Modules.scala 63:156:@18408.4]
  assign _T_69754 = $signed(buffer_4_740) + $signed(buffer_1_692); // @[Modules.scala 63:156:@18410.4]
  assign _T_69755 = _T_69754[10:0]; // @[Modules.scala 63:156:@18411.4]
  assign buffer_4_741 = $signed(_T_69755); // @[Modules.scala 63:156:@18412.4]
  assign _T_69757 = $signed(buffer_4_741) + $signed(buffer_4_693); // @[Modules.scala 63:156:@18414.4]
  assign _T_69758 = _T_69757[10:0]; // @[Modules.scala 63:156:@18415.4]
  assign buffer_4_742 = $signed(_T_69758); // @[Modules.scala 63:156:@18416.4]
  assign _T_69760 = $signed(buffer_4_742) + $signed(buffer_4_694); // @[Modules.scala 63:156:@18418.4]
  assign _T_69761 = _T_69760[10:0]; // @[Modules.scala 63:156:@18419.4]
  assign buffer_4_743 = $signed(_T_69761); // @[Modules.scala 63:156:@18420.4]
  assign _T_69763 = $signed(buffer_4_743) + $signed(buffer_4_695); // @[Modules.scala 63:156:@18422.4]
  assign _T_69764 = _T_69763[10:0]; // @[Modules.scala 63:156:@18423.4]
  assign buffer_4_744 = $signed(_T_69764); // @[Modules.scala 63:156:@18424.4]
  assign _T_69766 = $signed(buffer_4_744) + $signed(buffer_4_696); // @[Modules.scala 63:156:@18426.4]
  assign _T_69767 = _T_69766[10:0]; // @[Modules.scala 63:156:@18427.4]
  assign buffer_4_745 = $signed(_T_69767); // @[Modules.scala 63:156:@18428.4]
  assign _T_69769 = $signed(buffer_4_745) + $signed(buffer_4_697); // @[Modules.scala 63:156:@18430.4]
  assign _T_69770 = _T_69769[10:0]; // @[Modules.scala 63:156:@18431.4]
  assign buffer_4_746 = $signed(_T_69770); // @[Modules.scala 63:156:@18432.4]
  assign _T_69772 = $signed(buffer_4_746) + $signed(buffer_4_698); // @[Modules.scala 63:156:@18434.4]
  assign _T_69773 = _T_69772[10:0]; // @[Modules.scala 63:156:@18435.4]
  assign buffer_4_747 = $signed(_T_69773); // @[Modules.scala 63:156:@18436.4]
  assign _T_69775 = $signed(buffer_4_747) + $signed(buffer_4_699); // @[Modules.scala 63:156:@18438.4]
  assign _T_69776 = _T_69775[10:0]; // @[Modules.scala 63:156:@18439.4]
  assign buffer_4_748 = $signed(_T_69776); // @[Modules.scala 63:156:@18440.4]
  assign _T_69778 = $signed(buffer_4_748) + $signed(buffer_4_700); // @[Modules.scala 63:156:@18442.4]
  assign _T_69779 = _T_69778[10:0]; // @[Modules.scala 63:156:@18443.4]
  assign buffer_4_749 = $signed(_T_69779); // @[Modules.scala 63:156:@18444.4]
  assign _T_69781 = $signed(buffer_4_749) + $signed(buffer_4_701); // @[Modules.scala 63:156:@18446.4]
  assign _T_69782 = _T_69781[10:0]; // @[Modules.scala 63:156:@18447.4]
  assign buffer_4_750 = $signed(_T_69782); // @[Modules.scala 63:156:@18448.4]
  assign _T_69784 = $signed(buffer_4_750) + $signed(buffer_4_702); // @[Modules.scala 63:156:@18450.4]
  assign _T_69785 = _T_69784[10:0]; // @[Modules.scala 63:156:@18451.4]
  assign buffer_4_751 = $signed(_T_69785); // @[Modules.scala 63:156:@18452.4]
  assign _T_69787 = $signed(buffer_4_751) + $signed(buffer_4_703); // @[Modules.scala 63:156:@18454.4]
  assign _T_69788 = _T_69787[10:0]; // @[Modules.scala 63:156:@18455.4]
  assign buffer_4_752 = $signed(_T_69788); // @[Modules.scala 63:156:@18456.4]
  assign _T_69790 = $signed(buffer_4_752) + $signed(buffer_4_704); // @[Modules.scala 63:156:@18458.4]
  assign _T_69791 = _T_69790[10:0]; // @[Modules.scala 63:156:@18459.4]
  assign buffer_4_753 = $signed(_T_69791); // @[Modules.scala 63:156:@18460.4]
  assign _T_69793 = $signed(buffer_4_753) + $signed(buffer_4_705); // @[Modules.scala 63:156:@18462.4]
  assign _T_69794 = _T_69793[10:0]; // @[Modules.scala 63:156:@18463.4]
  assign buffer_4_754 = $signed(_T_69794); // @[Modules.scala 63:156:@18464.4]
  assign _T_69796 = $signed(buffer_4_754) + $signed(buffer_4_706); // @[Modules.scala 63:156:@18466.4]
  assign _T_69797 = _T_69796[10:0]; // @[Modules.scala 63:156:@18467.4]
  assign buffer_4_755 = $signed(_T_69797); // @[Modules.scala 63:156:@18468.4]
  assign _T_69799 = $signed(buffer_4_755) + $signed(buffer_4_707); // @[Modules.scala 63:156:@18470.4]
  assign _T_69800 = _T_69799[10:0]; // @[Modules.scala 63:156:@18471.4]
  assign buffer_4_756 = $signed(_T_69800); // @[Modules.scala 63:156:@18472.4]
  assign _T_69802 = $signed(buffer_4_756) + $signed(buffer_4_708); // @[Modules.scala 63:156:@18474.4]
  assign _T_69803 = _T_69802[10:0]; // @[Modules.scala 63:156:@18475.4]
  assign buffer_4_757 = $signed(_T_69803); // @[Modules.scala 63:156:@18476.4]
  assign _T_69805 = $signed(buffer_4_757) + $signed(buffer_4_709); // @[Modules.scala 63:156:@18478.4]
  assign _T_69806 = _T_69805[10:0]; // @[Modules.scala 63:156:@18479.4]
  assign buffer_4_758 = $signed(_T_69806); // @[Modules.scala 63:156:@18480.4]
  assign _T_69808 = $signed(buffer_4_758) + $signed(buffer_4_710); // @[Modules.scala 63:156:@18482.4]
  assign _T_69809 = _T_69808[10:0]; // @[Modules.scala 63:156:@18483.4]
  assign buffer_4_759 = $signed(_T_69809); // @[Modules.scala 63:156:@18484.4]
  assign _T_69811 = $signed(buffer_4_759) + $signed(buffer_4_711); // @[Modules.scala 63:156:@18486.4]
  assign _T_69812 = _T_69811[10:0]; // @[Modules.scala 63:156:@18487.4]
  assign buffer_4_760 = $signed(_T_69812); // @[Modules.scala 63:156:@18488.4]
  assign _T_69814 = $signed(buffer_4_760) + $signed(buffer_4_712); // @[Modules.scala 63:156:@18490.4]
  assign _T_69815 = _T_69814[10:0]; // @[Modules.scala 63:156:@18491.4]
  assign buffer_4_761 = $signed(_T_69815); // @[Modules.scala 63:156:@18492.4]
  assign _T_69817 = $signed(buffer_4_761) + $signed(buffer_4_713); // @[Modules.scala 63:156:@18494.4]
  assign _T_69818 = _T_69817[10:0]; // @[Modules.scala 63:156:@18495.4]
  assign buffer_4_762 = $signed(_T_69818); // @[Modules.scala 63:156:@18496.4]
  assign _T_69820 = $signed(buffer_4_762) + $signed(buffer_4_714); // @[Modules.scala 63:156:@18498.4]
  assign _T_69821 = _T_69820[10:0]; // @[Modules.scala 63:156:@18499.4]
  assign buffer_4_763 = $signed(_T_69821); // @[Modules.scala 63:156:@18500.4]
  assign _T_69823 = $signed(buffer_4_763) + $signed(buffer_4_715); // @[Modules.scala 63:156:@18502.4]
  assign _T_69824 = _T_69823[10:0]; // @[Modules.scala 63:156:@18503.4]
  assign buffer_4_764 = $signed(_T_69824); // @[Modules.scala 63:156:@18504.4]
  assign _T_69826 = $signed(buffer_4_764) + $signed(buffer_4_716); // @[Modules.scala 63:156:@18506.4]
  assign _T_69827 = _T_69826[10:0]; // @[Modules.scala 63:156:@18507.4]
  assign buffer_4_765 = $signed(_T_69827); // @[Modules.scala 63:156:@18508.4]
  assign _T_69829 = $signed(buffer_4_765) + $signed(buffer_4_717); // @[Modules.scala 63:156:@18510.4]
  assign _T_69830 = _T_69829[10:0]; // @[Modules.scala 63:156:@18511.4]
  assign buffer_4_766 = $signed(_T_69830); // @[Modules.scala 63:156:@18512.4]
  assign _T_69832 = $signed(buffer_4_766) + $signed(buffer_4_718); // @[Modules.scala 63:156:@18514.4]
  assign _T_69833 = _T_69832[10:0]; // @[Modules.scala 63:156:@18515.4]
  assign buffer_4_767 = $signed(_T_69833); // @[Modules.scala 63:156:@18516.4]
  assign _T_69835 = $signed(buffer_4_767) + $signed(buffer_4_719); // @[Modules.scala 63:156:@18518.4]
  assign _T_69836 = _T_69835[10:0]; // @[Modules.scala 63:156:@18519.4]
  assign buffer_4_768 = $signed(_T_69836); // @[Modules.scala 63:156:@18520.4]
  assign _T_69838 = $signed(buffer_4_768) + $signed(buffer_4_720); // @[Modules.scala 63:156:@18522.4]
  assign _T_69839 = _T_69838[10:0]; // @[Modules.scala 63:156:@18523.4]
  assign buffer_4_769 = $signed(_T_69839); // @[Modules.scala 63:156:@18524.4]
  assign _T_69841 = $signed(buffer_4_769) + $signed(buffer_4_721); // @[Modules.scala 63:156:@18526.4]
  assign _T_69842 = _T_69841[10:0]; // @[Modules.scala 63:156:@18527.4]
  assign buffer_4_770 = $signed(_T_69842); // @[Modules.scala 63:156:@18528.4]
  assign _T_69844 = $signed(buffer_4_770) + $signed(buffer_4_722); // @[Modules.scala 63:156:@18530.4]
  assign _T_69845 = _T_69844[10:0]; // @[Modules.scala 63:156:@18531.4]
  assign buffer_4_771 = $signed(_T_69845); // @[Modules.scala 63:156:@18532.4]
  assign _T_69847 = $signed(buffer_4_771) + $signed(buffer_4_723); // @[Modules.scala 63:156:@18534.4]
  assign _T_69848 = _T_69847[10:0]; // @[Modules.scala 63:156:@18535.4]
  assign buffer_4_772 = $signed(_T_69848); // @[Modules.scala 63:156:@18536.4]
  assign _T_69850 = $signed(buffer_4_772) + $signed(buffer_4_724); // @[Modules.scala 63:156:@18538.4]
  assign _T_69851 = _T_69850[10:0]; // @[Modules.scala 63:156:@18539.4]
  assign buffer_4_773 = $signed(_T_69851); // @[Modules.scala 63:156:@18540.4]
  assign _T_69853 = $signed(buffer_4_773) + $signed(buffer_4_725); // @[Modules.scala 63:156:@18542.4]
  assign _T_69854 = _T_69853[10:0]; // @[Modules.scala 63:156:@18543.4]
  assign buffer_4_774 = $signed(_T_69854); // @[Modules.scala 63:156:@18544.4]
  assign _T_69856 = $signed(buffer_4_774) + $signed(buffer_4_726); // @[Modules.scala 63:156:@18546.4]
  assign _T_69857 = _T_69856[10:0]; // @[Modules.scala 63:156:@18547.4]
  assign buffer_4_775 = $signed(_T_69857); // @[Modules.scala 63:156:@18548.4]
  assign _T_69859 = $signed(buffer_4_775) + $signed(buffer_4_727); // @[Modules.scala 63:156:@18550.4]
  assign _T_69860 = _T_69859[10:0]; // @[Modules.scala 63:156:@18551.4]
  assign buffer_4_776 = $signed(_T_69860); // @[Modules.scala 63:156:@18552.4]
  assign _T_69862 = $signed(buffer_4_776) + $signed(buffer_4_728); // @[Modules.scala 63:156:@18554.4]
  assign _T_69863 = _T_69862[10:0]; // @[Modules.scala 63:156:@18555.4]
  assign buffer_4_777 = $signed(_T_69863); // @[Modules.scala 63:156:@18556.4]
  assign _T_69865 = $signed(buffer_4_777) + $signed(buffer_4_729); // @[Modules.scala 63:156:@18558.4]
  assign _T_69866 = _T_69865[10:0]; // @[Modules.scala 63:156:@18559.4]
  assign buffer_4_778 = $signed(_T_69866); // @[Modules.scala 63:156:@18560.4]
  assign _T_69868 = $signed(buffer_4_778) + $signed(buffer_4_730); // @[Modules.scala 63:156:@18562.4]
  assign _T_69869 = _T_69868[10:0]; // @[Modules.scala 63:156:@18563.4]
  assign buffer_4_779 = $signed(_T_69869); // @[Modules.scala 63:156:@18564.4]
  assign _T_69871 = $signed(buffer_4_779) + $signed(buffer_4_731); // @[Modules.scala 63:156:@18566.4]
  assign _T_69872 = _T_69871[10:0]; // @[Modules.scala 63:156:@18567.4]
  assign buffer_4_780 = $signed(_T_69872); // @[Modules.scala 63:156:@18568.4]
  assign _T_69874 = $signed(buffer_4_780) + $signed(buffer_4_732); // @[Modules.scala 63:156:@18570.4]
  assign _T_69875 = _T_69874[10:0]; // @[Modules.scala 63:156:@18571.4]
  assign buffer_4_781 = $signed(_T_69875); // @[Modules.scala 63:156:@18572.4]
  assign _T_69877 = $signed(buffer_4_781) + $signed(buffer_4_733); // @[Modules.scala 63:156:@18574.4]
  assign _T_69878 = _T_69877[10:0]; // @[Modules.scala 63:156:@18575.4]
  assign buffer_4_782 = $signed(_T_69878); // @[Modules.scala 63:156:@18576.4]
  assign _T_69880 = $signed(buffer_4_782) + $signed(buffer_4_734); // @[Modules.scala 63:156:@18578.4]
  assign _T_69881 = _T_69880[10:0]; // @[Modules.scala 63:156:@18579.4]
  assign buffer_4_783 = $signed(_T_69881); // @[Modules.scala 63:156:@18580.4]
  assign _T_69930 = $signed(5'sh0) - $signed(io_in_20); // @[Modules.scala 43:37:@18635.4]
  assign _T_69931 = _T_69930[4:0]; // @[Modules.scala 43:37:@18636.4]
  assign _T_69932 = $signed(_T_69931); // @[Modules.scala 43:37:@18637.4]
  assign _T_69933 = $signed(_T_69932) + $signed(io_in_21); // @[Modules.scala 43:47:@18638.4]
  assign _T_69934 = _T_69933[4:0]; // @[Modules.scala 43:47:@18639.4]
  assign _T_69935 = $signed(_T_69934); // @[Modules.scala 43:47:@18640.4]
  assign _T_69967 = $signed(_T_60707) + $signed(io_in_33); // @[Modules.scala 43:47:@18674.4]
  assign _T_69968 = _T_69967[4:0]; // @[Modules.scala 43:47:@18675.4]
  assign _T_69969 = $signed(_T_69968); // @[Modules.scala 43:47:@18676.4]
  assign _T_70002 = $signed(_T_54400) + $signed(io_in_43); // @[Modules.scala 43:47:@18709.4]
  assign _T_70003 = _T_70002[4:0]; // @[Modules.scala 43:47:@18710.4]
  assign _T_70004 = $signed(_T_70003); // @[Modules.scala 43:47:@18711.4]
  assign _T_70095 = $signed(_T_54493) + $signed(io_in_73); // @[Modules.scala 43:47:@18805.4]
  assign _T_70096 = _T_70095[4:0]; // @[Modules.scala 43:47:@18806.4]
  assign _T_70097 = $signed(_T_70096); // @[Modules.scala 43:47:@18807.4]
  assign _T_70125 = $signed(io_in_84) + $signed(io_in_85); // @[Modules.scala 37:46:@18838.4]
  assign _T_70126 = _T_70125[4:0]; // @[Modules.scala 37:46:@18839.4]
  assign _T_70127 = $signed(_T_70126); // @[Modules.scala 37:46:@18840.4]
  assign _T_70202 = $signed(io_in_114) - $signed(io_in_115); // @[Modules.scala 40:46:@18922.4]
  assign _T_70203 = _T_70202[4:0]; // @[Modules.scala 40:46:@18923.4]
  assign _T_70204 = $signed(_T_70203); // @[Modules.scala 40:46:@18924.4]
  assign _T_70205 = $signed(io_in_116) + $signed(io_in_117); // @[Modules.scala 37:46:@18926.4]
  assign _T_70206 = _T_70205[4:0]; // @[Modules.scala 37:46:@18927.4]
  assign _T_70207 = $signed(_T_70206); // @[Modules.scala 37:46:@18928.4]
  assign _T_70233 = $signed(io_in_132) - $signed(io_in_133); // @[Modules.scala 40:46:@18961.4]
  assign _T_70234 = _T_70233[4:0]; // @[Modules.scala 40:46:@18962.4]
  assign _T_70235 = $signed(_T_70234); // @[Modules.scala 40:46:@18963.4]
  assign _T_70244 = $signed(5'sh0) - $signed(io_in_136); // @[Modules.scala 43:37:@18972.4]
  assign _T_70245 = _T_70244[4:0]; // @[Modules.scala 43:37:@18973.4]
  assign _T_70246 = $signed(_T_70245); // @[Modules.scala 43:37:@18974.4]
  assign _T_70247 = $signed(_T_70246) + $signed(io_in_137); // @[Modules.scala 43:47:@18975.4]
  assign _T_70248 = _T_70247[4:0]; // @[Modules.scala 43:47:@18976.4]
  assign _T_70249 = $signed(_T_70248); // @[Modules.scala 43:47:@18977.4]
  assign _T_70260 = $signed(io_in_142) + $signed(io_in_143); // @[Modules.scala 37:46:@18990.4]
  assign _T_70261 = _T_70260[4:0]; // @[Modules.scala 37:46:@18991.4]
  assign _T_70262 = $signed(_T_70261); // @[Modules.scala 37:46:@18992.4]
  assign _T_70270 = $signed(_T_57853) + $signed(io_in_147); // @[Modules.scala 43:47:@19001.4]
  assign _T_70271 = _T_70270[4:0]; // @[Modules.scala 43:47:@19002.4]
  assign _T_70272 = $signed(_T_70271); // @[Modules.scala 43:47:@19003.4]
  assign _T_70299 = $signed(_T_54709) + $signed(io_in_161); // @[Modules.scala 43:47:@19035.4]
  assign _T_70300 = _T_70299[4:0]; // @[Modules.scala 43:47:@19036.4]
  assign _T_70301 = $signed(_T_70300); // @[Modules.scala 43:47:@19037.4]
  assign _T_70306 = $signed(_T_57897) - $signed(io_in_163); // @[Modules.scala 46:47:@19042.4]
  assign _T_70307 = _T_70306[4:0]; // @[Modules.scala 46:47:@19043.4]
  assign _T_70308 = $signed(_T_70307); // @[Modules.scala 46:47:@19044.4]
  assign _T_70313 = $signed(_T_57904) + $signed(io_in_165); // @[Modules.scala 43:47:@19049.4]
  assign _T_70314 = _T_70313[4:0]; // @[Modules.scala 43:47:@19050.4]
  assign _T_70315 = $signed(_T_70314); // @[Modules.scala 43:47:@19051.4]
  assign _T_70316 = $signed(io_in_166) - $signed(io_in_167); // @[Modules.scala 40:46:@19053.4]
  assign _T_70317 = _T_70316[4:0]; // @[Modules.scala 40:46:@19054.4]
  assign _T_70318 = $signed(_T_70317); // @[Modules.scala 40:46:@19055.4]
  assign _T_70332 = $signed(io_in_174) - $signed(io_in_175); // @[Modules.scala 40:46:@19072.4]
  assign _T_70333 = _T_70332[4:0]; // @[Modules.scala 40:46:@19073.4]
  assign _T_70334 = $signed(_T_70333); // @[Modules.scala 40:46:@19074.4]
  assign _T_70344 = $signed(io_in_182) + $signed(io_in_183); // @[Modules.scala 37:46:@19088.4]
  assign _T_70345 = _T_70344[4:0]; // @[Modules.scala 37:46:@19089.4]
  assign _T_70346 = $signed(_T_70345); // @[Modules.scala 37:46:@19090.4]
  assign _T_70347 = $signed(io_in_184) + $signed(io_in_185); // @[Modules.scala 37:46:@19092.4]
  assign _T_70348 = _T_70347[4:0]; // @[Modules.scala 37:46:@19093.4]
  assign _T_70349 = $signed(_T_70348); // @[Modules.scala 37:46:@19094.4]
  assign _T_70360 = $signed(_T_57959) - $signed(io_in_191); // @[Modules.scala 46:47:@19107.4]
  assign _T_70361 = _T_70360[4:0]; // @[Modules.scala 46:47:@19108.4]
  assign _T_70362 = $signed(_T_70361); // @[Modules.scala 46:47:@19109.4]
  assign _T_70390 = $signed(io_in_202) - $signed(io_in_203); // @[Modules.scala 40:46:@19140.4]
  assign _T_70391 = _T_70390[4:0]; // @[Modules.scala 40:46:@19141.4]
  assign _T_70392 = $signed(_T_70391); // @[Modules.scala 40:46:@19142.4]
  assign _T_70419 = $signed(io_in_216) - $signed(io_in_217); // @[Modules.scala 40:46:@19174.4]
  assign _T_70420 = _T_70419[4:0]; // @[Modules.scala 40:46:@19175.4]
  assign _T_70421 = $signed(_T_70420); // @[Modules.scala 40:46:@19176.4]
  assign _T_70436 = $signed(io_in_222) - $signed(io_in_223); // @[Modules.scala 40:46:@19192.4]
  assign _T_70437 = _T_70436[4:0]; // @[Modules.scala 40:46:@19193.4]
  assign _T_70438 = $signed(_T_70437); // @[Modules.scala 40:46:@19194.4]
  assign _T_70450 = $signed(_T_54904) + $signed(io_in_227); // @[Modules.scala 43:47:@19206.4]
  assign _T_70451 = _T_70450[4:0]; // @[Modules.scala 43:47:@19207.4]
  assign _T_70452 = $signed(_T_70451); // @[Modules.scala 43:47:@19208.4]
  assign _T_70456 = $signed(io_in_230) + $signed(io_in_231); // @[Modules.scala 37:46:@19214.4]
  assign _T_70457 = _T_70456[4:0]; // @[Modules.scala 37:46:@19215.4]
  assign _T_70458 = $signed(_T_70457); // @[Modules.scala 37:46:@19216.4]
  assign _T_70497 = $signed(io_in_252) - $signed(io_in_253); // @[Modules.scala 40:46:@19264.4]
  assign _T_70498 = _T_70497[4:0]; // @[Modules.scala 40:46:@19265.4]
  assign _T_70499 = $signed(_T_70498); // @[Modules.scala 40:46:@19266.4]
  assign _T_70535 = $signed(_T_55033) + $signed(io_in_265); // @[Modules.scala 43:47:@19303.4]
  assign _T_70536 = _T_70535[4:0]; // @[Modules.scala 43:47:@19304.4]
  assign _T_70537 = $signed(_T_70536); // @[Modules.scala 43:47:@19305.4]
  assign _T_70544 = $signed(io_in_270) - $signed(io_in_271); // @[Modules.scala 40:46:@19315.4]
  assign _T_70545 = _T_70544[4:0]; // @[Modules.scala 40:46:@19316.4]
  assign _T_70546 = $signed(_T_70545); // @[Modules.scala 40:46:@19317.4]
  assign _T_70547 = $signed(io_in_272) - $signed(io_in_273); // @[Modules.scala 40:46:@19319.4]
  assign _T_70548 = _T_70547[4:0]; // @[Modules.scala 40:46:@19320.4]
  assign _T_70549 = $signed(_T_70548); // @[Modules.scala 40:46:@19321.4]
  assign _T_70550 = $signed(io_in_274) - $signed(io_in_275); // @[Modules.scala 40:46:@19323.4]
  assign _T_70551 = _T_70550[4:0]; // @[Modules.scala 40:46:@19324.4]
  assign _T_70552 = $signed(_T_70551); // @[Modules.scala 40:46:@19325.4]
  assign _T_70560 = $signed(io_in_278) - $signed(io_in_279); // @[Modules.scala 40:46:@19334.4]
  assign _T_70561 = _T_70560[4:0]; // @[Modules.scala 40:46:@19335.4]
  assign _T_70562 = $signed(_T_70561); // @[Modules.scala 40:46:@19336.4]
  assign _T_70563 = $signed(io_in_280) - $signed(io_in_281); // @[Modules.scala 40:46:@19338.4]
  assign _T_70564 = _T_70563[4:0]; // @[Modules.scala 40:46:@19339.4]
  assign _T_70565 = $signed(_T_70564); // @[Modules.scala 40:46:@19340.4]
  assign _T_70580 = $signed(io_in_286) - $signed(io_in_287); // @[Modules.scala 40:46:@19356.4]
  assign _T_70581 = _T_70580[4:0]; // @[Modules.scala 40:46:@19357.4]
  assign _T_70582 = $signed(_T_70581); // @[Modules.scala 40:46:@19358.4]
  assign _T_70604 = $signed(io_in_294) + $signed(io_in_295); // @[Modules.scala 37:46:@19381.4]
  assign _T_70605 = _T_70604[4:0]; // @[Modules.scala 37:46:@19382.4]
  assign _T_70606 = $signed(_T_70605); // @[Modules.scala 37:46:@19383.4]
  assign _T_70607 = $signed(io_in_296) - $signed(io_in_297); // @[Modules.scala 40:46:@19385.4]
  assign _T_70608 = _T_70607[4:0]; // @[Modules.scala 40:46:@19386.4]
  assign _T_70609 = $signed(_T_70608); // @[Modules.scala 40:46:@19387.4]
  assign _T_70613 = $signed(io_in_300) + $signed(io_in_301); // @[Modules.scala 37:46:@19393.4]
  assign _T_70614 = _T_70613[4:0]; // @[Modules.scala 37:46:@19394.4]
  assign _T_70615 = $signed(_T_70614); // @[Modules.scala 37:46:@19395.4]
  assign _T_70616 = $signed(io_in_302) - $signed(io_in_303); // @[Modules.scala 40:46:@19397.4]
  assign _T_70617 = _T_70616[4:0]; // @[Modules.scala 40:46:@19398.4]
  assign _T_70618 = $signed(_T_70617); // @[Modules.scala 40:46:@19399.4]
  assign _T_70630 = $signed(_T_55180) + $signed(io_in_307); // @[Modules.scala 43:47:@19411.4]
  assign _T_70631 = _T_70630[4:0]; // @[Modules.scala 43:47:@19412.4]
  assign _T_70632 = $signed(_T_70631); // @[Modules.scala 43:47:@19413.4]
  assign _T_70678 = $signed(io_in_322) + $signed(io_in_323); // @[Modules.scala 37:46:@19461.4]
  assign _T_70679 = _T_70678[4:0]; // @[Modules.scala 37:46:@19462.4]
  assign _T_70680 = $signed(_T_70679); // @[Modules.scala 37:46:@19463.4]
  assign _T_70681 = $signed(io_in_324) - $signed(io_in_325); // @[Modules.scala 40:46:@19465.4]
  assign _T_70682 = _T_70681[4:0]; // @[Modules.scala 40:46:@19466.4]
  assign _T_70683 = $signed(_T_70682); // @[Modules.scala 40:46:@19467.4]
  assign _T_70684 = $signed(io_in_326) + $signed(io_in_327); // @[Modules.scala 37:46:@19469.4]
  assign _T_70685 = _T_70684[4:0]; // @[Modules.scala 37:46:@19470.4]
  assign _T_70686 = $signed(_T_70685); // @[Modules.scala 37:46:@19471.4]
  assign _T_70690 = $signed(io_in_330) + $signed(io_in_331); // @[Modules.scala 37:46:@19477.4]
  assign _T_70691 = _T_70690[4:0]; // @[Modules.scala 37:46:@19478.4]
  assign _T_70692 = $signed(_T_70691); // @[Modules.scala 37:46:@19479.4]
  assign _T_70703 = $signed(io_in_336) + $signed(io_in_337); // @[Modules.scala 37:46:@19492.4]
  assign _T_70704 = _T_70703[4:0]; // @[Modules.scala 37:46:@19493.4]
  assign _T_70705 = $signed(_T_70704); // @[Modules.scala 37:46:@19494.4]
  assign _T_70710 = $signed(_T_55276) + $signed(io_in_339); // @[Modules.scala 43:47:@19499.4]
  assign _T_70711 = _T_70710[4:0]; // @[Modules.scala 43:47:@19500.4]
  assign _T_70712 = $signed(_T_70711); // @[Modules.scala 43:47:@19501.4]
  assign _T_70713 = $signed(io_in_340) - $signed(io_in_341); // @[Modules.scala 40:46:@19503.4]
  assign _T_70714 = _T_70713[4:0]; // @[Modules.scala 40:46:@19504.4]
  assign _T_70715 = $signed(_T_70714); // @[Modules.scala 40:46:@19505.4]
  assign _T_70754 = $signed(_T_58417) + $signed(io_in_355); // @[Modules.scala 43:47:@19546.4]
  assign _T_70755 = _T_70754[4:0]; // @[Modules.scala 43:47:@19547.4]
  assign _T_70756 = $signed(_T_70755); // @[Modules.scala 43:47:@19548.4]
  assign _T_70757 = $signed(io_in_356) - $signed(io_in_357); // @[Modules.scala 40:46:@19550.4]
  assign _T_70758 = _T_70757[4:0]; // @[Modules.scala 40:46:@19551.4]
  assign _T_70759 = $signed(_T_70758); // @[Modules.scala 40:46:@19552.4]
  assign _T_70788 = $signed(_T_55338) + $signed(io_in_367); // @[Modules.scala 43:47:@19582.4]
  assign _T_70789 = _T_70788[4:0]; // @[Modules.scala 43:47:@19583.4]
  assign _T_70790 = $signed(_T_70789); // @[Modules.scala 43:47:@19584.4]
  assign _T_70805 = $signed(io_in_372) - $signed(io_in_373); // @[Modules.scala 40:46:@19600.4]
  assign _T_70806 = _T_70805[4:0]; // @[Modules.scala 40:46:@19601.4]
  assign _T_70807 = $signed(_T_70806); // @[Modules.scala 40:46:@19602.4]
  assign _T_70812 = $signed(_T_64785) - $signed(io_in_375); // @[Modules.scala 46:47:@19607.4]
  assign _T_70813 = _T_70812[4:0]; // @[Modules.scala 46:47:@19608.4]
  assign _T_70814 = $signed(_T_70813); // @[Modules.scala 46:47:@19609.4]
  assign _T_70819 = $signed(_T_64792) + $signed(io_in_377); // @[Modules.scala 43:47:@19614.4]
  assign _T_70820 = _T_70819[4:0]; // @[Modules.scala 43:47:@19615.4]
  assign _T_70821 = $signed(_T_70820); // @[Modules.scala 43:47:@19616.4]
  assign _T_70849 = $signed(_T_61669) + $signed(io_in_389); // @[Modules.scala 43:47:@19647.4]
  assign _T_70850 = _T_70849[4:0]; // @[Modules.scala 43:47:@19648.4]
  assign _T_70851 = $signed(_T_70850); // @[Modules.scala 43:47:@19649.4]
  assign _T_70866 = $signed(_T_55396) + $signed(io_in_395); // @[Modules.scala 43:47:@19665.4]
  assign _T_70867 = _T_70866[4:0]; // @[Modules.scala 43:47:@19666.4]
  assign _T_70868 = $signed(_T_70867); // @[Modules.scala 43:47:@19667.4]
  assign _T_70887 = $signed(_T_64864) - $signed(io_in_401); // @[Modules.scala 46:47:@19686.4]
  assign _T_70888 = _T_70887[4:0]; // @[Modules.scala 46:47:@19687.4]
  assign _T_70889 = $signed(_T_70888); // @[Modules.scala 46:47:@19688.4]
  assign _T_70891 = $signed(5'sh0) - $signed(io_in_402); // @[Modules.scala 46:37:@19690.4]
  assign _T_70892 = _T_70891[4:0]; // @[Modules.scala 46:37:@19691.4]
  assign _T_70893 = $signed(_T_70892); // @[Modules.scala 46:37:@19692.4]
  assign _T_70894 = $signed(_T_70893) - $signed(io_in_403); // @[Modules.scala 46:47:@19693.4]
  assign _T_70895 = _T_70894[4:0]; // @[Modules.scala 46:47:@19694.4]
  assign _T_70896 = $signed(_T_70895); // @[Modules.scala 46:47:@19695.4]
  assign _T_70937 = $signed(_T_55443) - $signed(io_in_421); // @[Modules.scala 46:47:@19741.4]
  assign _T_70938 = _T_70937[4:0]; // @[Modules.scala 46:47:@19742.4]
  assign _T_70939 = $signed(_T_70938); // @[Modules.scala 46:47:@19743.4]
  assign _T_70944 = $signed(_T_55450) + $signed(io_in_423); // @[Modules.scala 43:47:@19748.4]
  assign _T_70945 = _T_70944[4:0]; // @[Modules.scala 43:47:@19749.4]
  assign _T_70946 = $signed(_T_70945); // @[Modules.scala 43:47:@19750.4]
  assign _T_70947 = $signed(io_in_424) - $signed(io_in_425); // @[Modules.scala 40:46:@19752.4]
  assign _T_70948 = _T_70947[4:0]; // @[Modules.scala 40:46:@19753.4]
  assign _T_70949 = $signed(_T_70948); // @[Modules.scala 40:46:@19754.4]
  assign _T_70958 = $signed(5'sh0) - $signed(io_in_428); // @[Modules.scala 46:37:@19763.4]
  assign _T_70959 = _T_70958[4:0]; // @[Modules.scala 46:37:@19764.4]
  assign _T_70960 = $signed(_T_70959); // @[Modules.scala 46:37:@19765.4]
  assign _T_70961 = $signed(_T_70960) - $signed(io_in_429); // @[Modules.scala 46:47:@19766.4]
  assign _T_70962 = _T_70961[4:0]; // @[Modules.scala 46:47:@19767.4]
  assign _T_70963 = $signed(_T_70962); // @[Modules.scala 46:47:@19768.4]
  assign _T_70981 = $signed(_T_58628) + $signed(io_in_437); // @[Modules.scala 43:47:@19788.4]
  assign _T_70982 = _T_70981[4:0]; // @[Modules.scala 43:47:@19789.4]
  assign _T_70983 = $signed(_T_70982); // @[Modules.scala 43:47:@19790.4]
  assign _T_71009 = $signed(_T_55495) + $signed(io_in_445); // @[Modules.scala 43:47:@19816.4]
  assign _T_71010 = _T_71009[4:0]; // @[Modules.scala 43:47:@19817.4]
  assign _T_71011 = $signed(_T_71010); // @[Modules.scala 43:47:@19818.4]
  assign _T_71044 = $signed(io_in_462) - $signed(io_in_463); // @[Modules.scala 40:46:@19858.4]
  assign _T_71045 = _T_71044[4:0]; // @[Modules.scala 40:46:@19859.4]
  assign _T_71046 = $signed(_T_71045); // @[Modules.scala 40:46:@19860.4]
  assign _T_71047 = $signed(io_in_464) - $signed(io_in_465); // @[Modules.scala 40:46:@19862.4]
  assign _T_71048 = _T_71047[4:0]; // @[Modules.scala 40:46:@19863.4]
  assign _T_71049 = $signed(_T_71048); // @[Modules.scala 40:46:@19864.4]
  assign _T_71054 = $signed(_T_58713) - $signed(io_in_467); // @[Modules.scala 46:47:@19869.4]
  assign _T_71055 = _T_71054[4:0]; // @[Modules.scala 46:47:@19870.4]
  assign _T_71056 = $signed(_T_71055); // @[Modules.scala 46:47:@19871.4]
  assign _T_71075 = $signed(_T_55557) + $signed(io_in_473); // @[Modules.scala 43:47:@19890.4]
  assign _T_71076 = _T_71075[4:0]; // @[Modules.scala 43:47:@19891.4]
  assign _T_71077 = $signed(_T_71076); // @[Modules.scala 43:47:@19892.4]
  assign _T_71101 = $signed(io_in_484) - $signed(io_in_485); // @[Modules.scala 40:46:@19920.4]
  assign _T_71102 = _T_71101[4:0]; // @[Modules.scala 40:46:@19921.4]
  assign _T_71103 = $signed(_T_71102); // @[Modules.scala 40:46:@19922.4]
  assign _T_71160 = $signed(io_in_510) - $signed(io_in_511); // @[Modules.scala 40:46:@19987.4]
  assign _T_71161 = _T_71160[4:0]; // @[Modules.scala 40:46:@19988.4]
  assign _T_71162 = $signed(_T_71161); // @[Modules.scala 40:46:@19989.4]
  assign _T_71167 = $signed(_T_58830) + $signed(io_in_513); // @[Modules.scala 43:47:@19994.4]
  assign _T_71168 = _T_71167[4:0]; // @[Modules.scala 43:47:@19995.4]
  assign _T_71169 = $signed(_T_71168); // @[Modules.scala 43:47:@19996.4]
  assign _T_71215 = $signed(io_in_536) - $signed(io_in_537); // @[Modules.scala 40:46:@20051.4]
  assign _T_71216 = _T_71215[4:0]; // @[Modules.scala 40:46:@20052.4]
  assign _T_71217 = $signed(_T_71216); // @[Modules.scala 40:46:@20053.4]
  assign _T_71222 = $signed(_T_55728) + $signed(io_in_539); // @[Modules.scala 43:47:@20058.4]
  assign _T_71223 = _T_71222[4:0]; // @[Modules.scala 43:47:@20059.4]
  assign _T_71224 = $signed(_T_71223); // @[Modules.scala 43:47:@20060.4]
  assign _T_71229 = $signed(_T_55735) + $signed(io_in_541); // @[Modules.scala 43:47:@20065.4]
  assign _T_71230 = _T_71229[4:0]; // @[Modules.scala 43:47:@20066.4]
  assign _T_71231 = $signed(_T_71230); // @[Modules.scala 43:47:@20067.4]
  assign _T_71270 = $signed(_T_55776) + $signed(io_in_555); // @[Modules.scala 43:47:@20108.4]
  assign _T_71271 = _T_71270[4:0]; // @[Modules.scala 43:47:@20109.4]
  assign _T_71272 = $signed(_T_71271); // @[Modules.scala 43:47:@20110.4]
  assign _T_71276 = $signed(io_in_558) + $signed(io_in_559); // @[Modules.scala 37:46:@20116.4]
  assign _T_71277 = _T_71276[4:0]; // @[Modules.scala 37:46:@20117.4]
  assign _T_71278 = $signed(_T_71277); // @[Modules.scala 37:46:@20118.4]
  assign _T_71290 = $signed(_T_55800) + $signed(io_in_563); // @[Modules.scala 43:47:@20130.4]
  assign _T_71291 = _T_71290[4:0]; // @[Modules.scala 43:47:@20131.4]
  assign _T_71292 = $signed(_T_71291); // @[Modules.scala 43:47:@20132.4]
  assign _T_71293 = $signed(io_in_564) - $signed(io_in_565); // @[Modules.scala 40:46:@20134.4]
  assign _T_71294 = _T_71293[4:0]; // @[Modules.scala 40:46:@20135.4]
  assign _T_71295 = $signed(_T_71294); // @[Modules.scala 40:46:@20136.4]
  assign _T_71310 = $signed(_T_55828) - $signed(io_in_571); // @[Modules.scala 46:47:@20152.4]
  assign _T_71311 = _T_71310[4:0]; // @[Modules.scala 46:47:@20153.4]
  assign _T_71312 = $signed(_T_71311); // @[Modules.scala 46:47:@20154.4]
  assign _T_71324 = $signed(_T_55842) - $signed(io_in_575); // @[Modules.scala 46:47:@20166.4]
  assign _T_71325 = _T_71324[4:0]; // @[Modules.scala 46:47:@20167.4]
  assign _T_71326 = $signed(_T_71325); // @[Modules.scala 46:47:@20168.4]
  assign _T_71328 = $signed(5'sh0) - $signed(io_in_576); // @[Modules.scala 46:37:@20170.4]
  assign _T_71329 = _T_71328[4:0]; // @[Modules.scala 46:37:@20171.4]
  assign _T_71330 = $signed(_T_71329); // @[Modules.scala 46:37:@20172.4]
  assign _T_71331 = $signed(_T_71330) - $signed(io_in_577); // @[Modules.scala 46:47:@20173.4]
  assign _T_71332 = _T_71331[4:0]; // @[Modules.scala 46:47:@20174.4]
  assign _T_71333 = $signed(_T_71332); // @[Modules.scala 46:47:@20175.4]
  assign _T_71335 = $signed(5'sh0) - $signed(io_in_578); // @[Modules.scala 43:37:@20177.4]
  assign _T_71336 = _T_71335[4:0]; // @[Modules.scala 43:37:@20178.4]
  assign _T_71337 = $signed(_T_71336); // @[Modules.scala 43:37:@20179.4]
  assign _T_71338 = $signed(_T_71337) + $signed(io_in_579); // @[Modules.scala 43:47:@20180.4]
  assign _T_71339 = _T_71338[4:0]; // @[Modules.scala 43:47:@20181.4]
  assign _T_71340 = $signed(_T_71339); // @[Modules.scala 43:47:@20182.4]
  assign _T_71345 = $signed(_T_62197) + $signed(io_in_581); // @[Modules.scala 43:47:@20187.4]
  assign _T_71346 = _T_71345[4:0]; // @[Modules.scala 43:47:@20188.4]
  assign _T_71347 = $signed(_T_71346); // @[Modules.scala 43:47:@20189.4]
  assign _T_71352 = $signed(_T_55858) + $signed(io_in_583); // @[Modules.scala 43:47:@20194.4]
  assign _T_71353 = _T_71352[4:0]; // @[Modules.scala 43:47:@20195.4]
  assign _T_71354 = $signed(_T_71353); // @[Modules.scala 43:47:@20196.4]
  assign _T_71391 = $signed(_T_62251) - $signed(io_in_601); // @[Modules.scala 46:47:@20239.4]
  assign _T_71392 = _T_71391[4:0]; // @[Modules.scala 46:47:@20240.4]
  assign _T_71393 = $signed(_T_71392); // @[Modules.scala 46:47:@20241.4]
  assign _T_71401 = $signed(io_in_604) - $signed(io_in_605); // @[Modules.scala 40:46:@20250.4]
  assign _T_71402 = _T_71401[4:0]; // @[Modules.scala 40:46:@20251.4]
  assign _T_71403 = $signed(_T_71402); // @[Modules.scala 40:46:@20252.4]
  assign _T_71446 = $signed(io_in_626) - $signed(io_in_627); // @[Modules.scala 40:46:@20303.4]
  assign _T_71447 = _T_71446[4:0]; // @[Modules.scala 40:46:@20304.4]
  assign _T_71448 = $signed(_T_71447); // @[Modules.scala 40:46:@20305.4]
  assign _T_71449 = $signed(io_in_628) - $signed(io_in_629); // @[Modules.scala 40:46:@20307.4]
  assign _T_71450 = _T_71449[4:0]; // @[Modules.scala 40:46:@20308.4]
  assign _T_71451 = $signed(_T_71450); // @[Modules.scala 40:46:@20309.4]
  assign _T_71479 = $signed(io_in_640) - $signed(io_in_641); // @[Modules.scala 40:46:@20340.4]
  assign _T_71480 = _T_71479[4:0]; // @[Modules.scala 40:46:@20341.4]
  assign _T_71481 = $signed(_T_71480); // @[Modules.scala 40:46:@20342.4]
  assign _T_71505 = $signed(io_in_652) - $signed(io_in_653); // @[Modules.scala 40:46:@20370.4]
  assign _T_71506 = _T_71505[4:0]; // @[Modules.scala 40:46:@20371.4]
  assign _T_71507 = $signed(_T_71506); // @[Modules.scala 40:46:@20372.4]
  assign _T_71519 = $signed(_T_56081) + $signed(io_in_657); // @[Modules.scala 43:47:@20384.4]
  assign _T_71520 = _T_71519[4:0]; // @[Modules.scala 43:47:@20385.4]
  assign _T_71521 = $signed(_T_71520); // @[Modules.scala 43:47:@20386.4]
  assign _T_71522 = $signed(io_in_658) - $signed(io_in_659); // @[Modules.scala 40:46:@20388.4]
  assign _T_71523 = _T_71522[4:0]; // @[Modules.scala 40:46:@20389.4]
  assign _T_71524 = $signed(_T_71523); // @[Modules.scala 40:46:@20390.4]
  assign _T_71539 = $signed(_T_59142) + $signed(io_in_665); // @[Modules.scala 43:47:@20406.4]
  assign _T_71540 = _T_71539[4:0]; // @[Modules.scala 43:47:@20407.4]
  assign _T_71541 = $signed(_T_71540); // @[Modules.scala 43:47:@20408.4]
  assign _T_71568 = $signed(io_in_678) - $signed(io_in_679); // @[Modules.scala 40:46:@20440.4]
  assign _T_71569 = _T_71568[4:0]; // @[Modules.scala 40:46:@20441.4]
  assign _T_71570 = $signed(_T_71569); // @[Modules.scala 40:46:@20442.4]
  assign _T_71571 = $signed(io_in_680) - $signed(io_in_681); // @[Modules.scala 40:46:@20444.4]
  assign _T_71572 = _T_71571[4:0]; // @[Modules.scala 40:46:@20445.4]
  assign _T_71573 = $signed(_T_71572); // @[Modules.scala 40:46:@20446.4]
  assign _T_71578 = $signed(_T_62450) + $signed(io_in_683); // @[Modules.scala 43:47:@20451.4]
  assign _T_71579 = _T_71578[4:0]; // @[Modules.scala 43:47:@20452.4]
  assign _T_71580 = $signed(_T_71579); // @[Modules.scala 43:47:@20453.4]
  assign _T_71592 = $signed(_T_56154) + $signed(io_in_687); // @[Modules.scala 43:47:@20465.4]
  assign _T_71593 = _T_71592[4:0]; // @[Modules.scala 43:47:@20466.4]
  assign _T_71594 = $signed(_T_71593); // @[Modules.scala 43:47:@20467.4]
  assign _T_71613 = $signed(io_in_700) - $signed(io_in_701); // @[Modules.scala 40:46:@20493.4]
  assign _T_71614 = _T_71613[4:0]; // @[Modules.scala 40:46:@20494.4]
  assign _T_71615 = $signed(_T_71614); // @[Modules.scala 40:46:@20495.4]
  assign _T_71620 = $signed(_T_65557) - $signed(io_in_703); // @[Modules.scala 46:47:@20500.4]
  assign _T_71621 = _T_71620[4:0]; // @[Modules.scala 46:47:@20501.4]
  assign _T_71622 = $signed(_T_71621); // @[Modules.scala 46:47:@20502.4]
  assign _T_71627 = $signed(_T_62507) + $signed(io_in_705); // @[Modules.scala 43:47:@20507.4]
  assign _T_71628 = _T_71627[4:0]; // @[Modules.scala 43:47:@20508.4]
  assign _T_71629 = $signed(_T_71628); // @[Modules.scala 43:47:@20509.4]
  assign _T_71654 = $signed(io_in_722) - $signed(io_in_723); // @[Modules.scala 40:46:@20543.4]
  assign _T_71655 = _T_71654[4:0]; // @[Modules.scala 40:46:@20544.4]
  assign _T_71656 = $signed(_T_71655); // @[Modules.scala 40:46:@20545.4]
  assign _T_71676 = $signed(io_in_734) - $signed(io_in_735); // @[Modules.scala 40:46:@20570.4]
  assign _T_71677 = _T_71676[4:0]; // @[Modules.scala 40:46:@20571.4]
  assign _T_71678 = $signed(_T_71677); // @[Modules.scala 40:46:@20572.4]
  assign _T_71688 = $signed(io_in_742) + $signed(io_in_743); // @[Modules.scala 37:46:@20586.4]
  assign _T_71689 = _T_71688[4:0]; // @[Modules.scala 37:46:@20587.4]
  assign _T_71690 = $signed(_T_71689); // @[Modules.scala 37:46:@20588.4]
  assign _T_71700 = $signed(io_in_750) + $signed(io_in_751); // @[Modules.scala 37:46:@20602.4]
  assign _T_71701 = _T_71700[4:0]; // @[Modules.scala 37:46:@20603.4]
  assign _T_71702 = $signed(_T_71701); // @[Modules.scala 37:46:@20604.4]
  assign _T_71720 = $signed(5'sh0) - $signed(io_in_760); // @[Modules.scala 46:37:@20625.4]
  assign _T_71721 = _T_71720[4:0]; // @[Modules.scala 46:37:@20626.4]
  assign _T_71722 = $signed(_T_71721); // @[Modules.scala 46:37:@20627.4]
  assign _T_71723 = $signed(_T_71722) - $signed(io_in_761); // @[Modules.scala 46:47:@20628.4]
  assign _T_71724 = _T_71723[4:0]; // @[Modules.scala 46:47:@20629.4]
  assign _T_71725 = $signed(_T_71724); // @[Modules.scala 46:47:@20630.4]
  assign _T_71740 = $signed(io_in_766) - $signed(io_in_767); // @[Modules.scala 40:46:@20646.4]
  assign _T_71741 = _T_71740[4:0]; // @[Modules.scala 40:46:@20647.4]
  assign _T_71742 = $signed(_T_71741); // @[Modules.scala 40:46:@20648.4]
  assign _T_71758 = $signed(io_in_778) + $signed(io_in_779); // @[Modules.scala 37:46:@20670.4]
  assign _T_71759 = _T_71758[4:0]; // @[Modules.scala 37:46:@20671.4]
  assign _T_71760 = $signed(_T_71759); // @[Modules.scala 37:46:@20672.4]
  assign _T_71767 = $signed(buffer_1_0) + $signed(buffer_3_1); // @[Modules.scala 50:57:@20682.4]
  assign _T_71768 = _T_71767[10:0]; // @[Modules.scala 50:57:@20683.4]
  assign buffer_5_392 = $signed(_T_71768); // @[Modules.scala 50:57:@20684.4]
  assign _T_71770 = $signed(buffer_2_2) + $signed(buffer_1_3); // @[Modules.scala 50:57:@20686.4]
  assign _T_71771 = _T_71770[10:0]; // @[Modules.scala 50:57:@20687.4]
  assign buffer_5_393 = $signed(_T_71771); // @[Modules.scala 50:57:@20688.4]
  assign _T_71773 = $signed(buffer_0_4) + $signed(buffer_3_5); // @[Modules.scala 50:57:@20690.4]
  assign _T_71774 = _T_71773[10:0]; // @[Modules.scala 50:57:@20691.4]
  assign buffer_5_394 = $signed(_T_71774); // @[Modules.scala 50:57:@20692.4]
  assign buffer_5_10 = {{6{_T_69935[4]}},_T_69935}; // @[Modules.scala 32:22:@8.4]
  assign _T_71782 = $signed(buffer_5_10) + $signed(buffer_4_11); // @[Modules.scala 50:57:@20702.4]
  assign _T_71783 = _T_71782[10:0]; // @[Modules.scala 50:57:@20703.4]
  assign buffer_5_397 = $signed(_T_71783); // @[Modules.scala 50:57:@20704.4]
  assign _T_71788 = $signed(buffer_0_14) + $signed(buffer_1_15); // @[Modules.scala 50:57:@20710.4]
  assign _T_71789 = _T_71788[10:0]; // @[Modules.scala 50:57:@20711.4]
  assign buffer_5_399 = $signed(_T_71789); // @[Modules.scala 50:57:@20712.4]
  assign buffer_5_16 = {{6{_T_69969[4]}},_T_69969}; // @[Modules.scala 32:22:@8.4]
  assign _T_71791 = $signed(buffer_5_16) + $signed(buffer_0_17); // @[Modules.scala 50:57:@20714.4]
  assign _T_71792 = _T_71791[10:0]; // @[Modules.scala 50:57:@20715.4]
  assign buffer_5_400 = $signed(_T_71792); // @[Modules.scala 50:57:@20716.4]
  assign buffer_5_21 = {{6{_T_70004[4]}},_T_70004}; // @[Modules.scala 32:22:@8.4]
  assign _T_71797 = $signed(buffer_0_20) + $signed(buffer_5_21); // @[Modules.scala 50:57:@20722.4]
  assign _T_71798 = _T_71797[10:0]; // @[Modules.scala 50:57:@20723.4]
  assign buffer_5_402 = $signed(_T_71798); // @[Modules.scala 50:57:@20724.4]
  assign _T_71809 = $signed(buffer_0_28) + $signed(buffer_2_29); // @[Modules.scala 50:57:@20738.4]
  assign _T_71810 = _T_71809[10:0]; // @[Modules.scala 50:57:@20739.4]
  assign buffer_5_406 = $signed(_T_71810); // @[Modules.scala 50:57:@20740.4]
  assign _T_71818 = $signed(buffer_0_34) + $signed(buffer_2_35); // @[Modules.scala 50:57:@20750.4]
  assign _T_71819 = _T_71818[10:0]; // @[Modules.scala 50:57:@20751.4]
  assign buffer_5_409 = $signed(_T_71819); // @[Modules.scala 50:57:@20752.4]
  assign buffer_5_36 = {{6{_T_70097[4]}},_T_70097}; // @[Modules.scala 32:22:@8.4]
  assign _T_71821 = $signed(buffer_5_36) + $signed(buffer_3_37); // @[Modules.scala 50:57:@20754.4]
  assign _T_71822 = _T_71821[10:0]; // @[Modules.scala 50:57:@20755.4]
  assign buffer_5_410 = $signed(_T_71822); // @[Modules.scala 50:57:@20756.4]
  assign _T_71827 = $signed(buffer_1_40) + $signed(buffer_0_41); // @[Modules.scala 50:57:@20762.4]
  assign _T_71828 = _T_71827[10:0]; // @[Modules.scala 50:57:@20763.4]
  assign buffer_5_412 = $signed(_T_71828); // @[Modules.scala 50:57:@20764.4]
  assign buffer_5_42 = {{6{_T_70127[4]}},_T_70127}; // @[Modules.scala 32:22:@8.4]
  assign _T_71830 = $signed(buffer_5_42) + $signed(buffer_0_43); // @[Modules.scala 50:57:@20766.4]
  assign _T_71831 = _T_71830[10:0]; // @[Modules.scala 50:57:@20767.4]
  assign buffer_5_413 = $signed(_T_71831); // @[Modules.scala 50:57:@20768.4]
  assign _T_71842 = $signed(buffer_2_50) + $signed(buffer_3_51); // @[Modules.scala 50:57:@20782.4]
  assign _T_71843 = _T_71842[10:0]; // @[Modules.scala 50:57:@20783.4]
  assign buffer_5_417 = $signed(_T_71843); // @[Modules.scala 50:57:@20784.4]
  assign _T_71848 = $signed(buffer_3_54) + $signed(buffer_2_55); // @[Modules.scala 50:57:@20790.4]
  assign _T_71849 = _T_71848[10:0]; // @[Modules.scala 50:57:@20791.4]
  assign buffer_5_419 = $signed(_T_71849); // @[Modules.scala 50:57:@20792.4]
  assign buffer_5_57 = {{6{_T_70204[4]}},_T_70204}; // @[Modules.scala 32:22:@8.4]
  assign _T_71851 = $signed(buffer_0_56) + $signed(buffer_5_57); // @[Modules.scala 50:57:@20794.4]
  assign _T_71852 = _T_71851[10:0]; // @[Modules.scala 50:57:@20795.4]
  assign buffer_5_420 = $signed(_T_71852); // @[Modules.scala 50:57:@20796.4]
  assign buffer_5_58 = {{6{_T_70207[4]}},_T_70207}; // @[Modules.scala 32:22:@8.4]
  assign _T_71854 = $signed(buffer_5_58) + $signed(buffer_0_59); // @[Modules.scala 50:57:@20798.4]
  assign _T_71855 = _T_71854[10:0]; // @[Modules.scala 50:57:@20799.4]
  assign buffer_5_421 = $signed(_T_71855); // @[Modules.scala 50:57:@20800.4]
  assign _T_71863 = $signed(buffer_1_64) + $signed(buffer_2_65); // @[Modules.scala 50:57:@20810.4]
  assign _T_71864 = _T_71863[10:0]; // @[Modules.scala 50:57:@20811.4]
  assign buffer_5_424 = $signed(_T_71864); // @[Modules.scala 50:57:@20812.4]
  assign buffer_5_66 = {{6{_T_70235[4]}},_T_70235}; // @[Modules.scala 32:22:@8.4]
  assign _T_71866 = $signed(buffer_5_66) + $signed(buffer_4_67); // @[Modules.scala 50:57:@20814.4]
  assign _T_71867 = _T_71866[10:0]; // @[Modules.scala 50:57:@20815.4]
  assign buffer_5_425 = $signed(_T_71867); // @[Modules.scala 50:57:@20816.4]
  assign buffer_5_68 = {{6{_T_70249[4]}},_T_70249}; // @[Modules.scala 32:22:@8.4]
  assign _T_71869 = $signed(buffer_5_68) + $signed(buffer_3_69); // @[Modules.scala 50:57:@20818.4]
  assign _T_71870 = _T_71869[10:0]; // @[Modules.scala 50:57:@20819.4]
  assign buffer_5_426 = $signed(_T_71870); // @[Modules.scala 50:57:@20820.4]
  assign buffer_5_71 = {{6{_T_70262[4]}},_T_70262}; // @[Modules.scala 32:22:@8.4]
  assign _T_71872 = $signed(buffer_2_70) + $signed(buffer_5_71); // @[Modules.scala 50:57:@20822.4]
  assign _T_71873 = _T_71872[10:0]; // @[Modules.scala 50:57:@20823.4]
  assign buffer_5_427 = $signed(_T_71873); // @[Modules.scala 50:57:@20824.4]
  assign buffer_5_73 = {{6{_T_70272[4]}},_T_70272}; // @[Modules.scala 32:22:@8.4]
  assign _T_71875 = $signed(buffer_4_72) + $signed(buffer_5_73); // @[Modules.scala 50:57:@20826.4]
  assign _T_71876 = _T_71875[10:0]; // @[Modules.scala 50:57:@20827.4]
  assign buffer_5_428 = $signed(_T_71876); // @[Modules.scala 50:57:@20828.4]
  assign buffer_5_80 = {{6{_T_70301[4]}},_T_70301}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_81 = {{6{_T_70308[4]}},_T_70308}; // @[Modules.scala 32:22:@8.4]
  assign _T_71887 = $signed(buffer_5_80) + $signed(buffer_5_81); // @[Modules.scala 50:57:@20842.4]
  assign _T_71888 = _T_71887[10:0]; // @[Modules.scala 50:57:@20843.4]
  assign buffer_5_432 = $signed(_T_71888); // @[Modules.scala 50:57:@20844.4]
  assign buffer_5_82 = {{6{_T_70315[4]}},_T_70315}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_83 = {{6{_T_70318[4]}},_T_70318}; // @[Modules.scala 32:22:@8.4]
  assign _T_71890 = $signed(buffer_5_82) + $signed(buffer_5_83); // @[Modules.scala 50:57:@20846.4]
  assign _T_71891 = _T_71890[10:0]; // @[Modules.scala 50:57:@20847.4]
  assign buffer_5_433 = $signed(_T_71891); // @[Modules.scala 50:57:@20848.4]
  assign _T_71893 = $signed(buffer_0_84) + $signed(buffer_1_85); // @[Modules.scala 50:57:@20850.4]
  assign _T_71894 = _T_71893[10:0]; // @[Modules.scala 50:57:@20851.4]
  assign buffer_5_434 = $signed(_T_71894); // @[Modules.scala 50:57:@20852.4]
  assign buffer_5_87 = {{6{_T_70334[4]}},_T_70334}; // @[Modules.scala 32:22:@8.4]
  assign _T_71896 = $signed(buffer_3_86) + $signed(buffer_5_87); // @[Modules.scala 50:57:@20854.4]
  assign _T_71897 = _T_71896[10:0]; // @[Modules.scala 50:57:@20855.4]
  assign buffer_5_435 = $signed(_T_71897); // @[Modules.scala 50:57:@20856.4]
  assign buffer_5_91 = {{6{_T_70346[4]}},_T_70346}; // @[Modules.scala 32:22:@8.4]
  assign _T_71902 = $signed(buffer_3_90) + $signed(buffer_5_91); // @[Modules.scala 50:57:@20862.4]
  assign _T_71903 = _T_71902[10:0]; // @[Modules.scala 50:57:@20863.4]
  assign buffer_5_437 = $signed(_T_71903); // @[Modules.scala 50:57:@20864.4]
  assign buffer_5_92 = {{6{_T_70349[4]}},_T_70349}; // @[Modules.scala 32:22:@8.4]
  assign _T_71905 = $signed(buffer_5_92) + $signed(buffer_3_93); // @[Modules.scala 50:57:@20866.4]
  assign _T_71906 = _T_71905[10:0]; // @[Modules.scala 50:57:@20867.4]
  assign buffer_5_438 = $signed(_T_71906); // @[Modules.scala 50:57:@20868.4]
  assign buffer_5_95 = {{6{_T_70362[4]}},_T_70362}; // @[Modules.scala 32:22:@8.4]
  assign _T_71908 = $signed(buffer_1_94) + $signed(buffer_5_95); // @[Modules.scala 50:57:@20870.4]
  assign _T_71909 = _T_71908[10:0]; // @[Modules.scala 50:57:@20871.4]
  assign buffer_5_439 = $signed(_T_71909); // @[Modules.scala 50:57:@20872.4]
  assign _T_71911 = $signed(buffer_1_96) + $signed(buffer_0_97); // @[Modules.scala 50:57:@20874.4]
  assign _T_71912 = _T_71911[10:0]; // @[Modules.scala 50:57:@20875.4]
  assign buffer_5_440 = $signed(_T_71912); // @[Modules.scala 50:57:@20876.4]
  assign buffer_5_101 = {{6{_T_70392[4]}},_T_70392}; // @[Modules.scala 32:22:@8.4]
  assign _T_71917 = $signed(buffer_3_100) + $signed(buffer_5_101); // @[Modules.scala 50:57:@20882.4]
  assign _T_71918 = _T_71917[10:0]; // @[Modules.scala 50:57:@20883.4]
  assign buffer_5_442 = $signed(_T_71918); // @[Modules.scala 50:57:@20884.4]
  assign _T_71920 = $signed(buffer_4_102) + $signed(buffer_0_103); // @[Modules.scala 50:57:@20886.4]
  assign _T_71921 = _T_71920[10:0]; // @[Modules.scala 50:57:@20887.4]
  assign buffer_5_443 = $signed(_T_71921); // @[Modules.scala 50:57:@20888.4]
  assign _T_71923 = $signed(buffer_3_104) + $signed(buffer_0_105); // @[Modules.scala 50:57:@20890.4]
  assign _T_71924 = _T_71923[10:0]; // @[Modules.scala 50:57:@20891.4]
  assign buffer_5_444 = $signed(_T_71924); // @[Modules.scala 50:57:@20892.4]
  assign _T_71926 = $signed(buffer_3_106) + $signed(buffer_1_107); // @[Modules.scala 50:57:@20894.4]
  assign _T_71927 = _T_71926[10:0]; // @[Modules.scala 50:57:@20895.4]
  assign buffer_5_445 = $signed(_T_71927); // @[Modules.scala 50:57:@20896.4]
  assign buffer_5_108 = {{6{_T_70421[4]}},_T_70421}; // @[Modules.scala 32:22:@8.4]
  assign _T_71929 = $signed(buffer_5_108) + $signed(buffer_0_109); // @[Modules.scala 50:57:@20898.4]
  assign _T_71930 = _T_71929[10:0]; // @[Modules.scala 50:57:@20899.4]
  assign buffer_5_446 = $signed(_T_71930); // @[Modules.scala 50:57:@20900.4]
  assign buffer_5_111 = {{6{_T_70438[4]}},_T_70438}; // @[Modules.scala 32:22:@8.4]
  assign _T_71932 = $signed(buffer_0_110) + $signed(buffer_5_111); // @[Modules.scala 50:57:@20902.4]
  assign _T_71933 = _T_71932[10:0]; // @[Modules.scala 50:57:@20903.4]
  assign buffer_5_447 = $signed(_T_71933); // @[Modules.scala 50:57:@20904.4]
  assign buffer_5_113 = {{6{_T_70452[4]}},_T_70452}; // @[Modules.scala 32:22:@8.4]
  assign _T_71935 = $signed(buffer_0_112) + $signed(buffer_5_113); // @[Modules.scala 50:57:@20906.4]
  assign _T_71936 = _T_71935[10:0]; // @[Modules.scala 50:57:@20907.4]
  assign buffer_5_448 = $signed(_T_71936); // @[Modules.scala 50:57:@20908.4]
  assign buffer_5_115 = {{6{_T_70458[4]}},_T_70458}; // @[Modules.scala 32:22:@8.4]
  assign _T_71938 = $signed(buffer_3_114) + $signed(buffer_5_115); // @[Modules.scala 50:57:@20910.4]
  assign _T_71939 = _T_71938[10:0]; // @[Modules.scala 50:57:@20911.4]
  assign buffer_5_449 = $signed(_T_71939); // @[Modules.scala 50:57:@20912.4]
  assign _T_71950 = $signed(buffer_4_122) + $signed(buffer_0_123); // @[Modules.scala 50:57:@20926.4]
  assign _T_71951 = _T_71950[10:0]; // @[Modules.scala 50:57:@20927.4]
  assign buffer_5_453 = $signed(_T_71951); // @[Modules.scala 50:57:@20928.4]
  assign _T_71953 = $signed(buffer_0_124) + $signed(buffer_1_125); // @[Modules.scala 50:57:@20930.4]
  assign _T_71954 = _T_71953[10:0]; // @[Modules.scala 50:57:@20931.4]
  assign buffer_5_454 = $signed(_T_71954); // @[Modules.scala 50:57:@20932.4]
  assign buffer_5_126 = {{6{_T_70499[4]}},_T_70499}; // @[Modules.scala 32:22:@8.4]
  assign _T_71956 = $signed(buffer_5_126) + $signed(buffer_0_127); // @[Modules.scala 50:57:@20934.4]
  assign _T_71957 = _T_71956[10:0]; // @[Modules.scala 50:57:@20935.4]
  assign buffer_5_455 = $signed(_T_71957); // @[Modules.scala 50:57:@20936.4]
  assign _T_71962 = $signed(buffer_2_130) + $signed(buffer_1_131); // @[Modules.scala 50:57:@20942.4]
  assign _T_71963 = _T_71962[10:0]; // @[Modules.scala 50:57:@20943.4]
  assign buffer_5_457 = $signed(_T_71963); // @[Modules.scala 50:57:@20944.4]
  assign buffer_5_132 = {{6{_T_70537[4]}},_T_70537}; // @[Modules.scala 32:22:@8.4]
  assign _T_71965 = $signed(buffer_5_132) + $signed(buffer_1_133); // @[Modules.scala 50:57:@20946.4]
  assign _T_71966 = _T_71965[10:0]; // @[Modules.scala 50:57:@20947.4]
  assign buffer_5_458 = $signed(_T_71966); // @[Modules.scala 50:57:@20948.4]
  assign buffer_5_135 = {{6{_T_70546[4]}},_T_70546}; // @[Modules.scala 32:22:@8.4]
  assign _T_71968 = $signed(buffer_3_134) + $signed(buffer_5_135); // @[Modules.scala 50:57:@20950.4]
  assign _T_71969 = _T_71968[10:0]; // @[Modules.scala 50:57:@20951.4]
  assign buffer_5_459 = $signed(_T_71969); // @[Modules.scala 50:57:@20952.4]
  assign buffer_5_136 = {{6{_T_70549[4]}},_T_70549}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_137 = {{6{_T_70552[4]}},_T_70552}; // @[Modules.scala 32:22:@8.4]
  assign _T_71971 = $signed(buffer_5_136) + $signed(buffer_5_137); // @[Modules.scala 50:57:@20954.4]
  assign _T_71972 = _T_71971[10:0]; // @[Modules.scala 50:57:@20955.4]
  assign buffer_5_460 = $signed(_T_71972); // @[Modules.scala 50:57:@20956.4]
  assign buffer_5_139 = {{6{_T_70562[4]}},_T_70562}; // @[Modules.scala 32:22:@8.4]
  assign _T_71974 = $signed(buffer_0_138) + $signed(buffer_5_139); // @[Modules.scala 50:57:@20958.4]
  assign _T_71975 = _T_71974[10:0]; // @[Modules.scala 50:57:@20959.4]
  assign buffer_5_461 = $signed(_T_71975); // @[Modules.scala 50:57:@20960.4]
  assign buffer_5_140 = {{6{_T_70565[4]}},_T_70565}; // @[Modules.scala 32:22:@8.4]
  assign _T_71977 = $signed(buffer_5_140) + $signed(buffer_0_141); // @[Modules.scala 50:57:@20962.4]
  assign _T_71978 = _T_71977[10:0]; // @[Modules.scala 50:57:@20963.4]
  assign buffer_5_462 = $signed(_T_71978); // @[Modules.scala 50:57:@20964.4]
  assign buffer_5_143 = {{6{_T_70582[4]}},_T_70582}; // @[Modules.scala 32:22:@8.4]
  assign _T_71980 = $signed(buffer_0_142) + $signed(buffer_5_143); // @[Modules.scala 50:57:@20966.4]
  assign _T_71981 = _T_71980[10:0]; // @[Modules.scala 50:57:@20967.4]
  assign buffer_5_463 = $signed(_T_71981); // @[Modules.scala 50:57:@20968.4]
  assign buffer_5_147 = {{6{_T_70606[4]}},_T_70606}; // @[Modules.scala 32:22:@8.4]
  assign _T_71986 = $signed(buffer_0_146) + $signed(buffer_5_147); // @[Modules.scala 50:57:@20974.4]
  assign _T_71987 = _T_71986[10:0]; // @[Modules.scala 50:57:@20975.4]
  assign buffer_5_465 = $signed(_T_71987); // @[Modules.scala 50:57:@20976.4]
  assign buffer_5_148 = {{6{_T_70609[4]}},_T_70609}; // @[Modules.scala 32:22:@8.4]
  assign _T_71989 = $signed(buffer_5_148) + $signed(buffer_4_149); // @[Modules.scala 50:57:@20978.4]
  assign _T_71990 = _T_71989[10:0]; // @[Modules.scala 50:57:@20979.4]
  assign buffer_5_466 = $signed(_T_71990); // @[Modules.scala 50:57:@20980.4]
  assign buffer_5_150 = {{6{_T_70615[4]}},_T_70615}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_151 = {{6{_T_70618[4]}},_T_70618}; // @[Modules.scala 32:22:@8.4]
  assign _T_71992 = $signed(buffer_5_150) + $signed(buffer_5_151); // @[Modules.scala 50:57:@20982.4]
  assign _T_71993 = _T_71992[10:0]; // @[Modules.scala 50:57:@20983.4]
  assign buffer_5_467 = $signed(_T_71993); // @[Modules.scala 50:57:@20984.4]
  assign buffer_5_153 = {{6{_T_70632[4]}},_T_70632}; // @[Modules.scala 32:22:@8.4]
  assign _T_71995 = $signed(buffer_0_152) + $signed(buffer_5_153); // @[Modules.scala 50:57:@20986.4]
  assign _T_71996 = _T_71995[10:0]; // @[Modules.scala 50:57:@20987.4]
  assign buffer_5_468 = $signed(_T_71996); // @[Modules.scala 50:57:@20988.4]
  assign _T_71998 = $signed(buffer_4_154) + $signed(buffer_0_155); // @[Modules.scala 50:57:@20990.4]
  assign _T_71999 = _T_71998[10:0]; // @[Modules.scala 50:57:@20991.4]
  assign buffer_5_469 = $signed(_T_71999); // @[Modules.scala 50:57:@20992.4]
  assign buffer_5_161 = {{6{_T_70680[4]}},_T_70680}; // @[Modules.scala 32:22:@8.4]
  assign _T_72007 = $signed(buffer_0_160) + $signed(buffer_5_161); // @[Modules.scala 50:57:@21002.4]
  assign _T_72008 = _T_72007[10:0]; // @[Modules.scala 50:57:@21003.4]
  assign buffer_5_472 = $signed(_T_72008); // @[Modules.scala 50:57:@21004.4]
  assign buffer_5_162 = {{6{_T_70683[4]}},_T_70683}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_163 = {{6{_T_70686[4]}},_T_70686}; // @[Modules.scala 32:22:@8.4]
  assign _T_72010 = $signed(buffer_5_162) + $signed(buffer_5_163); // @[Modules.scala 50:57:@21006.4]
  assign _T_72011 = _T_72010[10:0]; // @[Modules.scala 50:57:@21007.4]
  assign buffer_5_473 = $signed(_T_72011); // @[Modules.scala 50:57:@21008.4]
  assign buffer_5_165 = {{6{_T_70692[4]}},_T_70692}; // @[Modules.scala 32:22:@8.4]
  assign _T_72013 = $signed(buffer_0_164) + $signed(buffer_5_165); // @[Modules.scala 50:57:@21010.4]
  assign _T_72014 = _T_72013[10:0]; // @[Modules.scala 50:57:@21011.4]
  assign buffer_5_474 = $signed(_T_72014); // @[Modules.scala 50:57:@21012.4]
  assign buffer_5_168 = {{6{_T_70705[4]}},_T_70705}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_169 = {{6{_T_70712[4]}},_T_70712}; // @[Modules.scala 32:22:@8.4]
  assign _T_72019 = $signed(buffer_5_168) + $signed(buffer_5_169); // @[Modules.scala 50:57:@21018.4]
  assign _T_72020 = _T_72019[10:0]; // @[Modules.scala 50:57:@21019.4]
  assign buffer_5_476 = $signed(_T_72020); // @[Modules.scala 50:57:@21020.4]
  assign buffer_5_170 = {{6{_T_70715[4]}},_T_70715}; // @[Modules.scala 32:22:@8.4]
  assign _T_72022 = $signed(buffer_5_170) + $signed(buffer_3_171); // @[Modules.scala 50:57:@21022.4]
  assign _T_72023 = _T_72022[10:0]; // @[Modules.scala 50:57:@21023.4]
  assign buffer_5_477 = $signed(_T_72023); // @[Modules.scala 50:57:@21024.4]
  assign _T_72028 = $signed(buffer_3_174) + $signed(buffer_0_175); // @[Modules.scala 50:57:@21030.4]
  assign _T_72029 = _T_72028[10:0]; // @[Modules.scala 50:57:@21031.4]
  assign buffer_5_479 = $signed(_T_72029); // @[Modules.scala 50:57:@21032.4]
  assign buffer_5_177 = {{6{_T_70756[4]}},_T_70756}; // @[Modules.scala 32:22:@8.4]
  assign _T_72031 = $signed(buffer_0_176) + $signed(buffer_5_177); // @[Modules.scala 50:57:@21034.4]
  assign _T_72032 = _T_72031[10:0]; // @[Modules.scala 50:57:@21035.4]
  assign buffer_5_480 = $signed(_T_72032); // @[Modules.scala 50:57:@21036.4]
  assign buffer_5_178 = {{6{_T_70759[4]}},_T_70759}; // @[Modules.scala 32:22:@8.4]
  assign _T_72034 = $signed(buffer_5_178) + $signed(buffer_2_179); // @[Modules.scala 50:57:@21038.4]
  assign _T_72035 = _T_72034[10:0]; // @[Modules.scala 50:57:@21039.4]
  assign buffer_5_481 = $signed(_T_72035); // @[Modules.scala 50:57:@21040.4]
  assign buffer_5_183 = {{6{_T_70790[4]}},_T_70790}; // @[Modules.scala 32:22:@8.4]
  assign _T_72040 = $signed(buffer_0_182) + $signed(buffer_5_183); // @[Modules.scala 50:57:@21046.4]
  assign _T_72041 = _T_72040[10:0]; // @[Modules.scala 50:57:@21047.4]
  assign buffer_5_483 = $signed(_T_72041); // @[Modules.scala 50:57:@21048.4]
  assign buffer_5_186 = {{6{_T_70807[4]}},_T_70807}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_187 = {{6{_T_70814[4]}},_T_70814}; // @[Modules.scala 32:22:@8.4]
  assign _T_72046 = $signed(buffer_5_186) + $signed(buffer_5_187); // @[Modules.scala 50:57:@21054.4]
  assign _T_72047 = _T_72046[10:0]; // @[Modules.scala 50:57:@21055.4]
  assign buffer_5_485 = $signed(_T_72047); // @[Modules.scala 50:57:@21056.4]
  assign buffer_5_188 = {{6{_T_70821[4]}},_T_70821}; // @[Modules.scala 32:22:@8.4]
  assign _T_72049 = $signed(buffer_5_188) + $signed(buffer_0_189); // @[Modules.scala 50:57:@21058.4]
  assign _T_72050 = _T_72049[10:0]; // @[Modules.scala 50:57:@21059.4]
  assign buffer_5_486 = $signed(_T_72050); // @[Modules.scala 50:57:@21060.4]
  assign buffer_5_194 = {{6{_T_70851[4]}},_T_70851}; // @[Modules.scala 32:22:@8.4]
  assign _T_72058 = $signed(buffer_5_194) + $signed(buffer_3_195); // @[Modules.scala 50:57:@21070.4]
  assign _T_72059 = _T_72058[10:0]; // @[Modules.scala 50:57:@21071.4]
  assign buffer_5_489 = $signed(_T_72059); // @[Modules.scala 50:57:@21072.4]
  assign buffer_5_197 = {{6{_T_70868[4]}},_T_70868}; // @[Modules.scala 32:22:@8.4]
  assign _T_72061 = $signed(buffer_0_196) + $signed(buffer_5_197); // @[Modules.scala 50:57:@21074.4]
  assign _T_72062 = _T_72061[10:0]; // @[Modules.scala 50:57:@21075.4]
  assign buffer_5_490 = $signed(_T_72062); // @[Modules.scala 50:57:@21076.4]
  assign buffer_5_200 = {{6{_T_70889[4]}},_T_70889}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_201 = {{6{_T_70896[4]}},_T_70896}; // @[Modules.scala 32:22:@8.4]
  assign _T_72067 = $signed(buffer_5_200) + $signed(buffer_5_201); // @[Modules.scala 50:57:@21082.4]
  assign _T_72068 = _T_72067[10:0]; // @[Modules.scala 50:57:@21083.4]
  assign buffer_5_492 = $signed(_T_72068); // @[Modules.scala 50:57:@21084.4]
  assign _T_72079 = $signed(buffer_2_208) + $signed(buffer_3_209); // @[Modules.scala 50:57:@21098.4]
  assign _T_72080 = _T_72079[10:0]; // @[Modules.scala 50:57:@21099.4]
  assign buffer_5_496 = $signed(_T_72080); // @[Modules.scala 50:57:@21100.4]
  assign buffer_5_210 = {{6{_T_70939[4]}},_T_70939}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_211 = {{6{_T_70946[4]}},_T_70946}; // @[Modules.scala 32:22:@8.4]
  assign _T_72082 = $signed(buffer_5_210) + $signed(buffer_5_211); // @[Modules.scala 50:57:@21102.4]
  assign _T_72083 = _T_72082[10:0]; // @[Modules.scala 50:57:@21103.4]
  assign buffer_5_497 = $signed(_T_72083); // @[Modules.scala 50:57:@21104.4]
  assign buffer_5_212 = {{6{_T_70949[4]}},_T_70949}; // @[Modules.scala 32:22:@8.4]
  assign _T_72085 = $signed(buffer_5_212) + $signed(buffer_3_213); // @[Modules.scala 50:57:@21106.4]
  assign _T_72086 = _T_72085[10:0]; // @[Modules.scala 50:57:@21107.4]
  assign buffer_5_498 = $signed(_T_72086); // @[Modules.scala 50:57:@21108.4]
  assign buffer_5_214 = {{6{_T_70963[4]}},_T_70963}; // @[Modules.scala 32:22:@8.4]
  assign _T_72088 = $signed(buffer_5_214) + $signed(buffer_2_215); // @[Modules.scala 50:57:@21110.4]
  assign _T_72089 = _T_72088[10:0]; // @[Modules.scala 50:57:@21111.4]
  assign buffer_5_499 = $signed(_T_72089); // @[Modules.scala 50:57:@21112.4]
  assign buffer_5_218 = {{6{_T_70983[4]}},_T_70983}; // @[Modules.scala 32:22:@8.4]
  assign _T_72094 = $signed(buffer_5_218) + $signed(buffer_2_219); // @[Modules.scala 50:57:@21118.4]
  assign _T_72095 = _T_72094[10:0]; // @[Modules.scala 50:57:@21119.4]
  assign buffer_5_501 = $signed(_T_72095); // @[Modules.scala 50:57:@21120.4]
  assign _T_72097 = $signed(buffer_2_220) + $signed(buffer_3_221); // @[Modules.scala 50:57:@21122.4]
  assign _T_72098 = _T_72097[10:0]; // @[Modules.scala 50:57:@21123.4]
  assign buffer_5_502 = $signed(_T_72098); // @[Modules.scala 50:57:@21124.4]
  assign buffer_5_222 = {{6{_T_71011[4]}},_T_71011}; // @[Modules.scala 32:22:@8.4]
  assign _T_72100 = $signed(buffer_5_222) + $signed(buffer_3_223); // @[Modules.scala 50:57:@21126.4]
  assign _T_72101 = _T_72100[10:0]; // @[Modules.scala 50:57:@21127.4]
  assign buffer_5_503 = $signed(_T_72101); // @[Modules.scala 50:57:@21128.4]
  assign _T_72106 = $signed(buffer_3_226) + $signed(buffer_1_227); // @[Modules.scala 50:57:@21134.4]
  assign _T_72107 = _T_72106[10:0]; // @[Modules.scala 50:57:@21135.4]
  assign buffer_5_505 = $signed(_T_72107); // @[Modules.scala 50:57:@21136.4]
  assign buffer_5_231 = {{6{_T_71046[4]}},_T_71046}; // @[Modules.scala 32:22:@8.4]
  assign _T_72112 = $signed(buffer_2_230) + $signed(buffer_5_231); // @[Modules.scala 50:57:@21142.4]
  assign _T_72113 = _T_72112[10:0]; // @[Modules.scala 50:57:@21143.4]
  assign buffer_5_507 = $signed(_T_72113); // @[Modules.scala 50:57:@21144.4]
  assign buffer_5_232 = {{6{_T_71049[4]}},_T_71049}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_233 = {{6{_T_71056[4]}},_T_71056}; // @[Modules.scala 32:22:@8.4]
  assign _T_72115 = $signed(buffer_5_232) + $signed(buffer_5_233); // @[Modules.scala 50:57:@21146.4]
  assign _T_72116 = _T_72115[10:0]; // @[Modules.scala 50:57:@21147.4]
  assign buffer_5_508 = $signed(_T_72116); // @[Modules.scala 50:57:@21148.4]
  assign _T_72118 = $signed(buffer_2_234) + $signed(buffer_0_235); // @[Modules.scala 50:57:@21150.4]
  assign _T_72119 = _T_72118[10:0]; // @[Modules.scala 50:57:@21151.4]
  assign buffer_5_509 = $signed(_T_72119); // @[Modules.scala 50:57:@21152.4]
  assign buffer_5_236 = {{6{_T_71077[4]}},_T_71077}; // @[Modules.scala 32:22:@8.4]
  assign _T_72121 = $signed(buffer_5_236) + $signed(buffer_3_237); // @[Modules.scala 50:57:@21154.4]
  assign _T_72122 = _T_72121[10:0]; // @[Modules.scala 50:57:@21155.4]
  assign buffer_5_510 = $signed(_T_72122); // @[Modules.scala 50:57:@21156.4]
  assign _T_72127 = $signed(buffer_3_240) + $signed(buffer_2_241); // @[Modules.scala 50:57:@21162.4]
  assign _T_72128 = _T_72127[10:0]; // @[Modules.scala 50:57:@21163.4]
  assign buffer_5_512 = $signed(_T_72128); // @[Modules.scala 50:57:@21164.4]
  assign buffer_5_242 = {{6{_T_71103[4]}},_T_71103}; // @[Modules.scala 32:22:@8.4]
  assign _T_72130 = $signed(buffer_5_242) + $signed(buffer_1_243); // @[Modules.scala 50:57:@21166.4]
  assign _T_72131 = _T_72130[10:0]; // @[Modules.scala 50:57:@21167.4]
  assign buffer_5_513 = $signed(_T_72131); // @[Modules.scala 50:57:@21168.4]
  assign _T_72136 = $signed(buffer_1_246) + $signed(buffer_4_247); // @[Modules.scala 50:57:@21174.4]
  assign _T_72137 = _T_72136[10:0]; // @[Modules.scala 50:57:@21175.4]
  assign buffer_5_515 = $signed(_T_72137); // @[Modules.scala 50:57:@21176.4]
  assign _T_72139 = $signed(buffer_0_248) + $signed(buffer_2_249); // @[Modules.scala 50:57:@21178.4]
  assign _T_72140 = _T_72139[10:0]; // @[Modules.scala 50:57:@21179.4]
  assign buffer_5_516 = $signed(_T_72140); // @[Modules.scala 50:57:@21180.4]
  assign buffer_5_255 = {{6{_T_71162[4]}},_T_71162}; // @[Modules.scala 32:22:@8.4]
  assign _T_72148 = $signed(buffer_3_254) + $signed(buffer_5_255); // @[Modules.scala 50:57:@21190.4]
  assign _T_72149 = _T_72148[10:0]; // @[Modules.scala 50:57:@21191.4]
  assign buffer_5_519 = $signed(_T_72149); // @[Modules.scala 50:57:@21192.4]
  assign buffer_5_256 = {{6{_T_71169[4]}},_T_71169}; // @[Modules.scala 32:22:@8.4]
  assign _T_72151 = $signed(buffer_5_256) + $signed(buffer_0_257); // @[Modules.scala 50:57:@21194.4]
  assign _T_72152 = _T_72151[10:0]; // @[Modules.scala 50:57:@21195.4]
  assign buffer_5_520 = $signed(_T_72152); // @[Modules.scala 50:57:@21196.4]
  assign _T_72154 = $signed(buffer_2_258) + $signed(buffer_0_259); // @[Modules.scala 50:57:@21198.4]
  assign _T_72155 = _T_72154[10:0]; // @[Modules.scala 50:57:@21199.4]
  assign buffer_5_521 = $signed(_T_72155); // @[Modules.scala 50:57:@21200.4]
  assign _T_72157 = $signed(buffer_1_260) + $signed(buffer_0_261); // @[Modules.scala 50:57:@21202.4]
  assign _T_72158 = _T_72157[10:0]; // @[Modules.scala 50:57:@21203.4]
  assign buffer_5_522 = $signed(_T_72158); // @[Modules.scala 50:57:@21204.4]
  assign buffer_5_268 = {{6{_T_71217[4]}},_T_71217}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_269 = {{6{_T_71224[4]}},_T_71224}; // @[Modules.scala 32:22:@8.4]
  assign _T_72169 = $signed(buffer_5_268) + $signed(buffer_5_269); // @[Modules.scala 50:57:@21218.4]
  assign _T_72170 = _T_72169[10:0]; // @[Modules.scala 50:57:@21219.4]
  assign buffer_5_526 = $signed(_T_72170); // @[Modules.scala 50:57:@21220.4]
  assign buffer_5_270 = {{6{_T_71231[4]}},_T_71231}; // @[Modules.scala 32:22:@8.4]
  assign _T_72172 = $signed(buffer_5_270) + $signed(buffer_3_271); // @[Modules.scala 50:57:@21222.4]
  assign _T_72173 = _T_72172[10:0]; // @[Modules.scala 50:57:@21223.4]
  assign buffer_5_527 = $signed(_T_72173); // @[Modules.scala 50:57:@21224.4]
  assign _T_72175 = $signed(buffer_0_272) + $signed(buffer_1_273); // @[Modules.scala 50:57:@21226.4]
  assign _T_72176 = _T_72175[10:0]; // @[Modules.scala 50:57:@21227.4]
  assign buffer_5_528 = $signed(_T_72176); // @[Modules.scala 50:57:@21228.4]
  assign _T_72178 = $signed(buffer_2_274) + $signed(buffer_1_275); // @[Modules.scala 50:57:@21230.4]
  assign _T_72179 = _T_72178[10:0]; // @[Modules.scala 50:57:@21231.4]
  assign buffer_5_529 = $signed(_T_72179); // @[Modules.scala 50:57:@21232.4]
  assign buffer_5_277 = {{6{_T_71272[4]}},_T_71272}; // @[Modules.scala 32:22:@8.4]
  assign _T_72181 = $signed(buffer_0_276) + $signed(buffer_5_277); // @[Modules.scala 50:57:@21234.4]
  assign _T_72182 = _T_72181[10:0]; // @[Modules.scala 50:57:@21235.4]
  assign buffer_5_530 = $signed(_T_72182); // @[Modules.scala 50:57:@21236.4]
  assign buffer_5_279 = {{6{_T_71278[4]}},_T_71278}; // @[Modules.scala 32:22:@8.4]
  assign _T_72184 = $signed(buffer_3_278) + $signed(buffer_5_279); // @[Modules.scala 50:57:@21238.4]
  assign _T_72185 = _T_72184[10:0]; // @[Modules.scala 50:57:@21239.4]
  assign buffer_5_531 = $signed(_T_72185); // @[Modules.scala 50:57:@21240.4]
  assign buffer_5_281 = {{6{_T_71292[4]}},_T_71292}; // @[Modules.scala 32:22:@8.4]
  assign _T_72187 = $signed(buffer_0_280) + $signed(buffer_5_281); // @[Modules.scala 50:57:@21242.4]
  assign _T_72188 = _T_72187[10:0]; // @[Modules.scala 50:57:@21243.4]
  assign buffer_5_532 = $signed(_T_72188); // @[Modules.scala 50:57:@21244.4]
  assign buffer_5_282 = {{6{_T_71295[4]}},_T_71295}; // @[Modules.scala 32:22:@8.4]
  assign _T_72190 = $signed(buffer_5_282) + $signed(buffer_3_283); // @[Modules.scala 50:57:@21246.4]
  assign _T_72191 = _T_72190[10:0]; // @[Modules.scala 50:57:@21247.4]
  assign buffer_5_533 = $signed(_T_72191); // @[Modules.scala 50:57:@21248.4]
  assign buffer_5_285 = {{6{_T_71312[4]}},_T_71312}; // @[Modules.scala 32:22:@8.4]
  assign _T_72193 = $signed(buffer_0_284) + $signed(buffer_5_285); // @[Modules.scala 50:57:@21250.4]
  assign _T_72194 = _T_72193[10:0]; // @[Modules.scala 50:57:@21251.4]
  assign buffer_5_534 = $signed(_T_72194); // @[Modules.scala 50:57:@21252.4]
  assign buffer_5_287 = {{6{_T_71326[4]}},_T_71326}; // @[Modules.scala 32:22:@8.4]
  assign _T_72196 = $signed(buffer_2_286) + $signed(buffer_5_287); // @[Modules.scala 50:57:@21254.4]
  assign _T_72197 = _T_72196[10:0]; // @[Modules.scala 50:57:@21255.4]
  assign buffer_5_535 = $signed(_T_72197); // @[Modules.scala 50:57:@21256.4]
  assign buffer_5_288 = {{6{_T_71333[4]}},_T_71333}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_289 = {{6{_T_71340[4]}},_T_71340}; // @[Modules.scala 32:22:@8.4]
  assign _T_72199 = $signed(buffer_5_288) + $signed(buffer_5_289); // @[Modules.scala 50:57:@21258.4]
  assign _T_72200 = _T_72199[10:0]; // @[Modules.scala 50:57:@21259.4]
  assign buffer_5_536 = $signed(_T_72200); // @[Modules.scala 50:57:@21260.4]
  assign buffer_5_290 = {{6{_T_71347[4]}},_T_71347}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_291 = {{6{_T_71354[4]}},_T_71354}; // @[Modules.scala 32:22:@8.4]
  assign _T_72202 = $signed(buffer_5_290) + $signed(buffer_5_291); // @[Modules.scala 50:57:@21262.4]
  assign _T_72203 = _T_72202[10:0]; // @[Modules.scala 50:57:@21263.4]
  assign buffer_5_537 = $signed(_T_72203); // @[Modules.scala 50:57:@21264.4]
  assign _T_72214 = $signed(buffer_2_298) + $signed(buffer_0_299); // @[Modules.scala 50:57:@21278.4]
  assign _T_72215 = _T_72214[10:0]; // @[Modules.scala 50:57:@21279.4]
  assign buffer_5_541 = $signed(_T_72215); // @[Modules.scala 50:57:@21280.4]
  assign buffer_5_300 = {{6{_T_71393[4]}},_T_71393}; // @[Modules.scala 32:22:@8.4]
  assign _T_72217 = $signed(buffer_5_300) + $signed(buffer_3_301); // @[Modules.scala 50:57:@21282.4]
  assign _T_72218 = _T_72217[10:0]; // @[Modules.scala 50:57:@21283.4]
  assign buffer_5_542 = $signed(_T_72218); // @[Modules.scala 50:57:@21284.4]
  assign buffer_5_302 = {{6{_T_71403[4]}},_T_71403}; // @[Modules.scala 32:22:@8.4]
  assign _T_72220 = $signed(buffer_5_302) + $signed(buffer_0_303); // @[Modules.scala 50:57:@21286.4]
  assign _T_72221 = _T_72220[10:0]; // @[Modules.scala 50:57:@21287.4]
  assign buffer_5_543 = $signed(_T_72221); // @[Modules.scala 50:57:@21288.4]
  assign buffer_5_313 = {{6{_T_71448[4]}},_T_71448}; // @[Modules.scala 32:22:@8.4]
  assign _T_72235 = $signed(buffer_0_312) + $signed(buffer_5_313); // @[Modules.scala 50:57:@21306.4]
  assign _T_72236 = _T_72235[10:0]; // @[Modules.scala 50:57:@21307.4]
  assign buffer_5_548 = $signed(_T_72236); // @[Modules.scala 50:57:@21308.4]
  assign buffer_5_314 = {{6{_T_71451[4]}},_T_71451}; // @[Modules.scala 32:22:@8.4]
  assign _T_72238 = $signed(buffer_5_314) + $signed(buffer_3_315); // @[Modules.scala 50:57:@21310.4]
  assign _T_72239 = _T_72238[10:0]; // @[Modules.scala 50:57:@21311.4]
  assign buffer_5_549 = $signed(_T_72239); // @[Modules.scala 50:57:@21312.4]
  assign _T_72241 = $signed(buffer_3_316) + $signed(buffer_0_317); // @[Modules.scala 50:57:@21314.4]
  assign _T_72242 = _T_72241[10:0]; // @[Modules.scala 50:57:@21315.4]
  assign buffer_5_550 = $signed(_T_72242); // @[Modules.scala 50:57:@21316.4]
  assign buffer_5_320 = {{6{_T_71481[4]}},_T_71481}; // @[Modules.scala 32:22:@8.4]
  assign _T_72247 = $signed(buffer_5_320) + $signed(buffer_0_321); // @[Modules.scala 50:57:@21322.4]
  assign _T_72248 = _T_72247[10:0]; // @[Modules.scala 50:57:@21323.4]
  assign buffer_5_552 = $signed(_T_72248); // @[Modules.scala 50:57:@21324.4]
  assign _T_72253 = $signed(buffer_4_324) + $signed(buffer_1_325); // @[Modules.scala 50:57:@21330.4]
  assign _T_72254 = _T_72253[10:0]; // @[Modules.scala 50:57:@21331.4]
  assign buffer_5_554 = $signed(_T_72254); // @[Modules.scala 50:57:@21332.4]
  assign buffer_5_326 = {{6{_T_71507[4]}},_T_71507}; // @[Modules.scala 32:22:@8.4]
  assign _T_72256 = $signed(buffer_5_326) + $signed(buffer_0_327); // @[Modules.scala 50:57:@21334.4]
  assign _T_72257 = _T_72256[10:0]; // @[Modules.scala 50:57:@21335.4]
  assign buffer_5_555 = $signed(_T_72257); // @[Modules.scala 50:57:@21336.4]
  assign buffer_5_328 = {{6{_T_71521[4]}},_T_71521}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_329 = {{6{_T_71524[4]}},_T_71524}; // @[Modules.scala 32:22:@8.4]
  assign _T_72259 = $signed(buffer_5_328) + $signed(buffer_5_329); // @[Modules.scala 50:57:@21338.4]
  assign _T_72260 = _T_72259[10:0]; // @[Modules.scala 50:57:@21339.4]
  assign buffer_5_556 = $signed(_T_72260); // @[Modules.scala 50:57:@21340.4]
  assign _T_72262 = $signed(buffer_2_330) + $signed(buffer_0_331); // @[Modules.scala 50:57:@21342.4]
  assign _T_72263 = _T_72262[10:0]; // @[Modules.scala 50:57:@21343.4]
  assign buffer_5_557 = $signed(_T_72263); // @[Modules.scala 50:57:@21344.4]
  assign buffer_5_332 = {{6{_T_71541[4]}},_T_71541}; // @[Modules.scala 32:22:@8.4]
  assign _T_72265 = $signed(buffer_5_332) + $signed(buffer_0_333); // @[Modules.scala 50:57:@21346.4]
  assign _T_72266 = _T_72265[10:0]; // @[Modules.scala 50:57:@21347.4]
  assign buffer_5_558 = $signed(_T_72266); // @[Modules.scala 50:57:@21348.4]
  assign _T_72271 = $signed(buffer_0_336) + $signed(buffer_1_337); // @[Modules.scala 50:57:@21354.4]
  assign _T_72272 = _T_72271[10:0]; // @[Modules.scala 50:57:@21355.4]
  assign buffer_5_560 = $signed(_T_72272); // @[Modules.scala 50:57:@21356.4]
  assign buffer_5_339 = {{6{_T_71570[4]}},_T_71570}; // @[Modules.scala 32:22:@8.4]
  assign _T_72274 = $signed(buffer_0_338) + $signed(buffer_5_339); // @[Modules.scala 50:57:@21358.4]
  assign _T_72275 = _T_72274[10:0]; // @[Modules.scala 50:57:@21359.4]
  assign buffer_5_561 = $signed(_T_72275); // @[Modules.scala 50:57:@21360.4]
  assign buffer_5_340 = {{6{_T_71573[4]}},_T_71573}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_341 = {{6{_T_71580[4]}},_T_71580}; // @[Modules.scala 32:22:@8.4]
  assign _T_72277 = $signed(buffer_5_340) + $signed(buffer_5_341); // @[Modules.scala 50:57:@21362.4]
  assign _T_72278 = _T_72277[10:0]; // @[Modules.scala 50:57:@21363.4]
  assign buffer_5_562 = $signed(_T_72278); // @[Modules.scala 50:57:@21364.4]
  assign buffer_5_343 = {{6{_T_71594[4]}},_T_71594}; // @[Modules.scala 32:22:@8.4]
  assign _T_72280 = $signed(buffer_3_342) + $signed(buffer_5_343); // @[Modules.scala 50:57:@21366.4]
  assign _T_72281 = _T_72280[10:0]; // @[Modules.scala 50:57:@21367.4]
  assign buffer_5_563 = $signed(_T_72281); // @[Modules.scala 50:57:@21368.4]
  assign _T_72289 = $signed(buffer_1_348) + $signed(buffer_3_349); // @[Modules.scala 50:57:@21378.4]
  assign _T_72290 = _T_72289[10:0]; // @[Modules.scala 50:57:@21379.4]
  assign buffer_5_566 = $signed(_T_72290); // @[Modules.scala 50:57:@21380.4]
  assign buffer_5_350 = {{6{_T_71615[4]}},_T_71615}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_351 = {{6{_T_71622[4]}},_T_71622}; // @[Modules.scala 32:22:@8.4]
  assign _T_72292 = $signed(buffer_5_350) + $signed(buffer_5_351); // @[Modules.scala 50:57:@21382.4]
  assign _T_72293 = _T_72292[10:0]; // @[Modules.scala 50:57:@21383.4]
  assign buffer_5_567 = $signed(_T_72293); // @[Modules.scala 50:57:@21384.4]
  assign buffer_5_352 = {{6{_T_71629[4]}},_T_71629}; // @[Modules.scala 32:22:@8.4]
  assign _T_72295 = $signed(buffer_5_352) + $signed(buffer_0_353); // @[Modules.scala 50:57:@21386.4]
  assign _T_72296 = _T_72295[10:0]; // @[Modules.scala 50:57:@21387.4]
  assign buffer_5_568 = $signed(_T_72296); // @[Modules.scala 50:57:@21388.4]
  assign buffer_5_361 = {{6{_T_71656[4]}},_T_71656}; // @[Modules.scala 32:22:@8.4]
  assign _T_72307 = $signed(buffer_0_360) + $signed(buffer_5_361); // @[Modules.scala 50:57:@21402.4]
  assign _T_72308 = _T_72307[10:0]; // @[Modules.scala 50:57:@21403.4]
  assign buffer_5_572 = $signed(_T_72308); // @[Modules.scala 50:57:@21404.4]
  assign buffer_5_367 = {{6{_T_71678[4]}},_T_71678}; // @[Modules.scala 32:22:@8.4]
  assign _T_72316 = $signed(buffer_0_366) + $signed(buffer_5_367); // @[Modules.scala 50:57:@21414.4]
  assign _T_72317 = _T_72316[10:0]; // @[Modules.scala 50:57:@21415.4]
  assign buffer_5_575 = $signed(_T_72317); // @[Modules.scala 50:57:@21416.4]
  assign buffer_5_371 = {{6{_T_71690[4]}},_T_71690}; // @[Modules.scala 32:22:@8.4]
  assign _T_72322 = $signed(buffer_3_370) + $signed(buffer_5_371); // @[Modules.scala 50:57:@21422.4]
  assign _T_72323 = _T_72322[10:0]; // @[Modules.scala 50:57:@21423.4]
  assign buffer_5_577 = $signed(_T_72323); // @[Modules.scala 50:57:@21424.4]
  assign buffer_5_375 = {{6{_T_71702[4]}},_T_71702}; // @[Modules.scala 32:22:@8.4]
  assign _T_72328 = $signed(buffer_0_374) + $signed(buffer_5_375); // @[Modules.scala 50:57:@21430.4]
  assign _T_72329 = _T_72328[10:0]; // @[Modules.scala 50:57:@21431.4]
  assign buffer_5_579 = $signed(_T_72329); // @[Modules.scala 50:57:@21432.4]
  assign buffer_5_380 = {{6{_T_71725[4]}},_T_71725}; // @[Modules.scala 32:22:@8.4]
  assign _T_72337 = $signed(buffer_5_380) + $signed(buffer_0_381); // @[Modules.scala 50:57:@21442.4]
  assign _T_72338 = _T_72337[10:0]; // @[Modules.scala 50:57:@21443.4]
  assign buffer_5_582 = $signed(_T_72338); // @[Modules.scala 50:57:@21444.4]
  assign buffer_5_383 = {{6{_T_71742[4]}},_T_71742}; // @[Modules.scala 32:22:@8.4]
  assign _T_72340 = $signed(buffer_0_382) + $signed(buffer_5_383); // @[Modules.scala 50:57:@21446.4]
  assign _T_72341 = _T_72340[10:0]; // @[Modules.scala 50:57:@21447.4]
  assign buffer_5_583 = $signed(_T_72341); // @[Modules.scala 50:57:@21448.4]
  assign buffer_5_389 = {{6{_T_71760[4]}},_T_71760}; // @[Modules.scala 32:22:@8.4]
  assign _T_72349 = $signed(buffer_0_388) + $signed(buffer_5_389); // @[Modules.scala 50:57:@21458.4]
  assign _T_72350 = _T_72349[10:0]; // @[Modules.scala 50:57:@21459.4]
  assign buffer_5_586 = $signed(_T_72350); // @[Modules.scala 50:57:@21460.4]
  assign _T_72355 = $signed(buffer_5_392) + $signed(buffer_5_393); // @[Modules.scala 53:83:@21466.4]
  assign _T_72356 = _T_72355[10:0]; // @[Modules.scala 53:83:@21467.4]
  assign buffer_5_588 = $signed(_T_72356); // @[Modules.scala 53:83:@21468.4]
  assign _T_72358 = $signed(buffer_5_394) + $signed(buffer_4_395); // @[Modules.scala 53:83:@21470.4]
  assign _T_72359 = _T_72358[10:0]; // @[Modules.scala 53:83:@21471.4]
  assign buffer_5_589 = $signed(_T_72359); // @[Modules.scala 53:83:@21472.4]
  assign _T_72361 = $signed(buffer_0_396) + $signed(buffer_5_397); // @[Modules.scala 53:83:@21474.4]
  assign _T_72362 = _T_72361[10:0]; // @[Modules.scala 53:83:@21475.4]
  assign buffer_5_590 = $signed(_T_72362); // @[Modules.scala 53:83:@21476.4]
  assign _T_72364 = $signed(buffer_4_398) + $signed(buffer_5_399); // @[Modules.scala 53:83:@21478.4]
  assign _T_72365 = _T_72364[10:0]; // @[Modules.scala 53:83:@21479.4]
  assign buffer_5_591 = $signed(_T_72365); // @[Modules.scala 53:83:@21480.4]
  assign _T_72367 = $signed(buffer_5_400) + $signed(buffer_0_401); // @[Modules.scala 53:83:@21482.4]
  assign _T_72368 = _T_72367[10:0]; // @[Modules.scala 53:83:@21483.4]
  assign buffer_5_592 = $signed(_T_72368); // @[Modules.scala 53:83:@21484.4]
  assign _T_72370 = $signed(buffer_5_402) + $signed(buffer_4_403); // @[Modules.scala 53:83:@21486.4]
  assign _T_72371 = _T_72370[10:0]; // @[Modules.scala 53:83:@21487.4]
  assign buffer_5_593 = $signed(_T_72371); // @[Modules.scala 53:83:@21488.4]
  assign _T_72373 = $signed(buffer_0_404) + $signed(buffer_4_405); // @[Modules.scala 53:83:@21490.4]
  assign _T_72374 = _T_72373[10:0]; // @[Modules.scala 53:83:@21491.4]
  assign buffer_5_594 = $signed(_T_72374); // @[Modules.scala 53:83:@21492.4]
  assign _T_72376 = $signed(buffer_5_406) + $signed(buffer_3_407); // @[Modules.scala 53:83:@21494.4]
  assign _T_72377 = _T_72376[10:0]; // @[Modules.scala 53:83:@21495.4]
  assign buffer_5_595 = $signed(_T_72377); // @[Modules.scala 53:83:@21496.4]
  assign _T_72379 = $signed(buffer_3_408) + $signed(buffer_5_409); // @[Modules.scala 53:83:@21498.4]
  assign _T_72380 = _T_72379[10:0]; // @[Modules.scala 53:83:@21499.4]
  assign buffer_5_596 = $signed(_T_72380); // @[Modules.scala 53:83:@21500.4]
  assign _T_72382 = $signed(buffer_5_410) + $signed(buffer_3_411); // @[Modules.scala 53:83:@21502.4]
  assign _T_72383 = _T_72382[10:0]; // @[Modules.scala 53:83:@21503.4]
  assign buffer_5_597 = $signed(_T_72383); // @[Modules.scala 53:83:@21504.4]
  assign _T_72385 = $signed(buffer_5_412) + $signed(buffer_5_413); // @[Modules.scala 53:83:@21506.4]
  assign _T_72386 = _T_72385[10:0]; // @[Modules.scala 53:83:@21507.4]
  assign buffer_5_598 = $signed(_T_72386); // @[Modules.scala 53:83:@21508.4]
  assign _T_72391 = $signed(buffer_3_416) + $signed(buffer_5_417); // @[Modules.scala 53:83:@21514.4]
  assign _T_72392 = _T_72391[10:0]; // @[Modules.scala 53:83:@21515.4]
  assign buffer_5_600 = $signed(_T_72392); // @[Modules.scala 53:83:@21516.4]
  assign _T_72394 = $signed(buffer_3_418) + $signed(buffer_5_419); // @[Modules.scala 53:83:@21518.4]
  assign _T_72395 = _T_72394[10:0]; // @[Modules.scala 53:83:@21519.4]
  assign buffer_5_601 = $signed(_T_72395); // @[Modules.scala 53:83:@21520.4]
  assign _T_72397 = $signed(buffer_5_420) + $signed(buffer_5_421); // @[Modules.scala 53:83:@21522.4]
  assign _T_72398 = _T_72397[10:0]; // @[Modules.scala 53:83:@21523.4]
  assign buffer_5_602 = $signed(_T_72398); // @[Modules.scala 53:83:@21524.4]
  assign _T_72403 = $signed(buffer_5_424) + $signed(buffer_5_425); // @[Modules.scala 53:83:@21530.4]
  assign _T_72404 = _T_72403[10:0]; // @[Modules.scala 53:83:@21531.4]
  assign buffer_5_604 = $signed(_T_72404); // @[Modules.scala 53:83:@21532.4]
  assign _T_72406 = $signed(buffer_5_426) + $signed(buffer_5_427); // @[Modules.scala 53:83:@21534.4]
  assign _T_72407 = _T_72406[10:0]; // @[Modules.scala 53:83:@21535.4]
  assign buffer_5_605 = $signed(_T_72407); // @[Modules.scala 53:83:@21536.4]
  assign _T_72409 = $signed(buffer_5_428) + $signed(buffer_3_429); // @[Modules.scala 53:83:@21538.4]
  assign _T_72410 = _T_72409[10:0]; // @[Modules.scala 53:83:@21539.4]
  assign buffer_5_606 = $signed(_T_72410); // @[Modules.scala 53:83:@21540.4]
  assign _T_72412 = $signed(buffer_4_430) + $signed(buffer_1_431); // @[Modules.scala 53:83:@21542.4]
  assign _T_72413 = _T_72412[10:0]; // @[Modules.scala 53:83:@21543.4]
  assign buffer_5_607 = $signed(_T_72413); // @[Modules.scala 53:83:@21544.4]
  assign _T_72415 = $signed(buffer_5_432) + $signed(buffer_5_433); // @[Modules.scala 53:83:@21546.4]
  assign _T_72416 = _T_72415[10:0]; // @[Modules.scala 53:83:@21547.4]
  assign buffer_5_608 = $signed(_T_72416); // @[Modules.scala 53:83:@21548.4]
  assign _T_72418 = $signed(buffer_5_434) + $signed(buffer_5_435); // @[Modules.scala 53:83:@21550.4]
  assign _T_72419 = _T_72418[10:0]; // @[Modules.scala 53:83:@21551.4]
  assign buffer_5_609 = $signed(_T_72419); // @[Modules.scala 53:83:@21552.4]
  assign _T_72421 = $signed(buffer_3_436) + $signed(buffer_5_437); // @[Modules.scala 53:83:@21554.4]
  assign _T_72422 = _T_72421[10:0]; // @[Modules.scala 53:83:@21555.4]
  assign buffer_5_610 = $signed(_T_72422); // @[Modules.scala 53:83:@21556.4]
  assign _T_72424 = $signed(buffer_5_438) + $signed(buffer_5_439); // @[Modules.scala 53:83:@21558.4]
  assign _T_72425 = _T_72424[10:0]; // @[Modules.scala 53:83:@21559.4]
  assign buffer_5_611 = $signed(_T_72425); // @[Modules.scala 53:83:@21560.4]
  assign _T_72427 = $signed(buffer_5_440) + $signed(buffer_3_441); // @[Modules.scala 53:83:@21562.4]
  assign _T_72428 = _T_72427[10:0]; // @[Modules.scala 53:83:@21563.4]
  assign buffer_5_612 = $signed(_T_72428); // @[Modules.scala 53:83:@21564.4]
  assign _T_72430 = $signed(buffer_5_442) + $signed(buffer_5_443); // @[Modules.scala 53:83:@21566.4]
  assign _T_72431 = _T_72430[10:0]; // @[Modules.scala 53:83:@21567.4]
  assign buffer_5_613 = $signed(_T_72431); // @[Modules.scala 53:83:@21568.4]
  assign _T_72433 = $signed(buffer_5_444) + $signed(buffer_5_445); // @[Modules.scala 53:83:@21570.4]
  assign _T_72434 = _T_72433[10:0]; // @[Modules.scala 53:83:@21571.4]
  assign buffer_5_614 = $signed(_T_72434); // @[Modules.scala 53:83:@21572.4]
  assign _T_72436 = $signed(buffer_5_446) + $signed(buffer_5_447); // @[Modules.scala 53:83:@21574.4]
  assign _T_72437 = _T_72436[10:0]; // @[Modules.scala 53:83:@21575.4]
  assign buffer_5_615 = $signed(_T_72437); // @[Modules.scala 53:83:@21576.4]
  assign _T_72439 = $signed(buffer_5_448) + $signed(buffer_5_449); // @[Modules.scala 53:83:@21578.4]
  assign _T_72440 = _T_72439[10:0]; // @[Modules.scala 53:83:@21579.4]
  assign buffer_5_616 = $signed(_T_72440); // @[Modules.scala 53:83:@21580.4]
  assign _T_72442 = $signed(buffer_4_450) + $signed(buffer_3_451); // @[Modules.scala 53:83:@21582.4]
  assign _T_72443 = _T_72442[10:0]; // @[Modules.scala 53:83:@21583.4]
  assign buffer_5_617 = $signed(_T_72443); // @[Modules.scala 53:83:@21584.4]
  assign _T_72445 = $signed(buffer_3_452) + $signed(buffer_5_453); // @[Modules.scala 53:83:@21586.4]
  assign _T_72446 = _T_72445[10:0]; // @[Modules.scala 53:83:@21587.4]
  assign buffer_5_618 = $signed(_T_72446); // @[Modules.scala 53:83:@21588.4]
  assign _T_72448 = $signed(buffer_5_454) + $signed(buffer_5_455); // @[Modules.scala 53:83:@21590.4]
  assign _T_72449 = _T_72448[10:0]; // @[Modules.scala 53:83:@21591.4]
  assign buffer_5_619 = $signed(_T_72449); // @[Modules.scala 53:83:@21592.4]
  assign _T_72451 = $signed(buffer_3_456) + $signed(buffer_5_457); // @[Modules.scala 53:83:@21594.4]
  assign _T_72452 = _T_72451[10:0]; // @[Modules.scala 53:83:@21595.4]
  assign buffer_5_620 = $signed(_T_72452); // @[Modules.scala 53:83:@21596.4]
  assign _T_72454 = $signed(buffer_5_458) + $signed(buffer_5_459); // @[Modules.scala 53:83:@21598.4]
  assign _T_72455 = _T_72454[10:0]; // @[Modules.scala 53:83:@21599.4]
  assign buffer_5_621 = $signed(_T_72455); // @[Modules.scala 53:83:@21600.4]
  assign _T_72457 = $signed(buffer_5_460) + $signed(buffer_5_461); // @[Modules.scala 53:83:@21602.4]
  assign _T_72458 = _T_72457[10:0]; // @[Modules.scala 53:83:@21603.4]
  assign buffer_5_622 = $signed(_T_72458); // @[Modules.scala 53:83:@21604.4]
  assign _T_72460 = $signed(buffer_5_462) + $signed(buffer_5_463); // @[Modules.scala 53:83:@21606.4]
  assign _T_72461 = _T_72460[10:0]; // @[Modules.scala 53:83:@21607.4]
  assign buffer_5_623 = $signed(_T_72461); // @[Modules.scala 53:83:@21608.4]
  assign _T_72463 = $signed(buffer_3_464) + $signed(buffer_5_465); // @[Modules.scala 53:83:@21610.4]
  assign _T_72464 = _T_72463[10:0]; // @[Modules.scala 53:83:@21611.4]
  assign buffer_5_624 = $signed(_T_72464); // @[Modules.scala 53:83:@21612.4]
  assign _T_72466 = $signed(buffer_5_466) + $signed(buffer_5_467); // @[Modules.scala 53:83:@21614.4]
  assign _T_72467 = _T_72466[10:0]; // @[Modules.scala 53:83:@21615.4]
  assign buffer_5_625 = $signed(_T_72467); // @[Modules.scala 53:83:@21616.4]
  assign _T_72469 = $signed(buffer_5_468) + $signed(buffer_5_469); // @[Modules.scala 53:83:@21618.4]
  assign _T_72470 = _T_72469[10:0]; // @[Modules.scala 53:83:@21619.4]
  assign buffer_5_626 = $signed(_T_72470); // @[Modules.scala 53:83:@21620.4]
  assign _T_72475 = $signed(buffer_5_472) + $signed(buffer_5_473); // @[Modules.scala 53:83:@21626.4]
  assign _T_72476 = _T_72475[10:0]; // @[Modules.scala 53:83:@21627.4]
  assign buffer_5_628 = $signed(_T_72476); // @[Modules.scala 53:83:@21628.4]
  assign _T_72478 = $signed(buffer_5_474) + $signed(buffer_3_475); // @[Modules.scala 53:83:@21630.4]
  assign _T_72479 = _T_72478[10:0]; // @[Modules.scala 53:83:@21631.4]
  assign buffer_5_629 = $signed(_T_72479); // @[Modules.scala 53:83:@21632.4]
  assign _T_72481 = $signed(buffer_5_476) + $signed(buffer_5_477); // @[Modules.scala 53:83:@21634.4]
  assign _T_72482 = _T_72481[10:0]; // @[Modules.scala 53:83:@21635.4]
  assign buffer_5_630 = $signed(_T_72482); // @[Modules.scala 53:83:@21636.4]
  assign _T_72484 = $signed(buffer_3_478) + $signed(buffer_5_479); // @[Modules.scala 53:83:@21638.4]
  assign _T_72485 = _T_72484[10:0]; // @[Modules.scala 53:83:@21639.4]
  assign buffer_5_631 = $signed(_T_72485); // @[Modules.scala 53:83:@21640.4]
  assign _T_72487 = $signed(buffer_5_480) + $signed(buffer_5_481); // @[Modules.scala 53:83:@21642.4]
  assign _T_72488 = _T_72487[10:0]; // @[Modules.scala 53:83:@21643.4]
  assign buffer_5_632 = $signed(_T_72488); // @[Modules.scala 53:83:@21644.4]
  assign _T_72490 = $signed(buffer_2_482) + $signed(buffer_5_483); // @[Modules.scala 53:83:@21646.4]
  assign _T_72491 = _T_72490[10:0]; // @[Modules.scala 53:83:@21647.4]
  assign buffer_5_633 = $signed(_T_72491); // @[Modules.scala 53:83:@21648.4]
  assign _T_72493 = $signed(buffer_3_484) + $signed(buffer_5_485); // @[Modules.scala 53:83:@21650.4]
  assign _T_72494 = _T_72493[10:0]; // @[Modules.scala 53:83:@21651.4]
  assign buffer_5_634 = $signed(_T_72494); // @[Modules.scala 53:83:@21652.4]
  assign _T_72496 = $signed(buffer_5_486) + $signed(buffer_0_487); // @[Modules.scala 53:83:@21654.4]
  assign _T_72497 = _T_72496[10:0]; // @[Modules.scala 53:83:@21655.4]
  assign buffer_5_635 = $signed(_T_72497); // @[Modules.scala 53:83:@21656.4]
  assign _T_72499 = $signed(buffer_3_488) + $signed(buffer_5_489); // @[Modules.scala 53:83:@21658.4]
  assign _T_72500 = _T_72499[10:0]; // @[Modules.scala 53:83:@21659.4]
  assign buffer_5_636 = $signed(_T_72500); // @[Modules.scala 53:83:@21660.4]
  assign _T_72502 = $signed(buffer_5_490) + $signed(buffer_3_491); // @[Modules.scala 53:83:@21662.4]
  assign _T_72503 = _T_72502[10:0]; // @[Modules.scala 53:83:@21663.4]
  assign buffer_5_637 = $signed(_T_72503); // @[Modules.scala 53:83:@21664.4]
  assign _T_72505 = $signed(buffer_5_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@21666.4]
  assign _T_72506 = _T_72505[10:0]; // @[Modules.scala 53:83:@21667.4]
  assign buffer_5_638 = $signed(_T_72506); // @[Modules.scala 53:83:@21668.4]
  assign _T_72508 = $signed(buffer_4_494) + $signed(buffer_3_495); // @[Modules.scala 53:83:@21670.4]
  assign _T_72509 = _T_72508[10:0]; // @[Modules.scala 53:83:@21671.4]
  assign buffer_5_639 = $signed(_T_72509); // @[Modules.scala 53:83:@21672.4]
  assign _T_72511 = $signed(buffer_5_496) + $signed(buffer_5_497); // @[Modules.scala 53:83:@21674.4]
  assign _T_72512 = _T_72511[10:0]; // @[Modules.scala 53:83:@21675.4]
  assign buffer_5_640 = $signed(_T_72512); // @[Modules.scala 53:83:@21676.4]
  assign _T_72514 = $signed(buffer_5_498) + $signed(buffer_5_499); // @[Modules.scala 53:83:@21678.4]
  assign _T_72515 = _T_72514[10:0]; // @[Modules.scala 53:83:@21679.4]
  assign buffer_5_641 = $signed(_T_72515); // @[Modules.scala 53:83:@21680.4]
  assign _T_72517 = $signed(buffer_0_500) + $signed(buffer_5_501); // @[Modules.scala 53:83:@21682.4]
  assign _T_72518 = _T_72517[10:0]; // @[Modules.scala 53:83:@21683.4]
  assign buffer_5_642 = $signed(_T_72518); // @[Modules.scala 53:83:@21684.4]
  assign _T_72520 = $signed(buffer_5_502) + $signed(buffer_5_503); // @[Modules.scala 53:83:@21686.4]
  assign _T_72521 = _T_72520[10:0]; // @[Modules.scala 53:83:@21687.4]
  assign buffer_5_643 = $signed(_T_72521); // @[Modules.scala 53:83:@21688.4]
  assign _T_72523 = $signed(buffer_3_504) + $signed(buffer_5_505); // @[Modules.scala 53:83:@21690.4]
  assign _T_72524 = _T_72523[10:0]; // @[Modules.scala 53:83:@21691.4]
  assign buffer_5_644 = $signed(_T_72524); // @[Modules.scala 53:83:@21692.4]
  assign _T_72526 = $signed(buffer_1_506) + $signed(buffer_5_507); // @[Modules.scala 53:83:@21694.4]
  assign _T_72527 = _T_72526[10:0]; // @[Modules.scala 53:83:@21695.4]
  assign buffer_5_645 = $signed(_T_72527); // @[Modules.scala 53:83:@21696.4]
  assign _T_72529 = $signed(buffer_5_508) + $signed(buffer_5_509); // @[Modules.scala 53:83:@21698.4]
  assign _T_72530 = _T_72529[10:0]; // @[Modules.scala 53:83:@21699.4]
  assign buffer_5_646 = $signed(_T_72530); // @[Modules.scala 53:83:@21700.4]
  assign _T_72532 = $signed(buffer_5_510) + $signed(buffer_3_511); // @[Modules.scala 53:83:@21702.4]
  assign _T_72533 = _T_72532[10:0]; // @[Modules.scala 53:83:@21703.4]
  assign buffer_5_647 = $signed(_T_72533); // @[Modules.scala 53:83:@21704.4]
  assign _T_72535 = $signed(buffer_5_512) + $signed(buffer_5_513); // @[Modules.scala 53:83:@21706.4]
  assign _T_72536 = _T_72535[10:0]; // @[Modules.scala 53:83:@21707.4]
  assign buffer_5_648 = $signed(_T_72536); // @[Modules.scala 53:83:@21708.4]
  assign _T_72538 = $signed(buffer_2_514) + $signed(buffer_5_515); // @[Modules.scala 53:83:@21710.4]
  assign _T_72539 = _T_72538[10:0]; // @[Modules.scala 53:83:@21711.4]
  assign buffer_5_649 = $signed(_T_72539); // @[Modules.scala 53:83:@21712.4]
  assign _T_72541 = $signed(buffer_5_516) + $signed(buffer_3_517); // @[Modules.scala 53:83:@21714.4]
  assign _T_72542 = _T_72541[10:0]; // @[Modules.scala 53:83:@21715.4]
  assign buffer_5_650 = $signed(_T_72542); // @[Modules.scala 53:83:@21716.4]
  assign _T_72544 = $signed(buffer_3_518) + $signed(buffer_5_519); // @[Modules.scala 53:83:@21718.4]
  assign _T_72545 = _T_72544[10:0]; // @[Modules.scala 53:83:@21719.4]
  assign buffer_5_651 = $signed(_T_72545); // @[Modules.scala 53:83:@21720.4]
  assign _T_72547 = $signed(buffer_5_520) + $signed(buffer_5_521); // @[Modules.scala 53:83:@21722.4]
  assign _T_72548 = _T_72547[10:0]; // @[Modules.scala 53:83:@21723.4]
  assign buffer_5_652 = $signed(_T_72548); // @[Modules.scala 53:83:@21724.4]
  assign _T_72550 = $signed(buffer_5_522) + $signed(buffer_1_523); // @[Modules.scala 53:83:@21726.4]
  assign _T_72551 = _T_72550[10:0]; // @[Modules.scala 53:83:@21727.4]
  assign buffer_5_653 = $signed(_T_72551); // @[Modules.scala 53:83:@21728.4]
  assign _T_72553 = $signed(buffer_3_524) + $signed(buffer_4_525); // @[Modules.scala 53:83:@21730.4]
  assign _T_72554 = _T_72553[10:0]; // @[Modules.scala 53:83:@21731.4]
  assign buffer_5_654 = $signed(_T_72554); // @[Modules.scala 53:83:@21732.4]
  assign _T_72556 = $signed(buffer_5_526) + $signed(buffer_5_527); // @[Modules.scala 53:83:@21734.4]
  assign _T_72557 = _T_72556[10:0]; // @[Modules.scala 53:83:@21735.4]
  assign buffer_5_655 = $signed(_T_72557); // @[Modules.scala 53:83:@21736.4]
  assign _T_72559 = $signed(buffer_5_528) + $signed(buffer_5_529); // @[Modules.scala 53:83:@21738.4]
  assign _T_72560 = _T_72559[10:0]; // @[Modules.scala 53:83:@21739.4]
  assign buffer_5_656 = $signed(_T_72560); // @[Modules.scala 53:83:@21740.4]
  assign _T_72562 = $signed(buffer_5_530) + $signed(buffer_5_531); // @[Modules.scala 53:83:@21742.4]
  assign _T_72563 = _T_72562[10:0]; // @[Modules.scala 53:83:@21743.4]
  assign buffer_5_657 = $signed(_T_72563); // @[Modules.scala 53:83:@21744.4]
  assign _T_72565 = $signed(buffer_5_532) + $signed(buffer_5_533); // @[Modules.scala 53:83:@21746.4]
  assign _T_72566 = _T_72565[10:0]; // @[Modules.scala 53:83:@21747.4]
  assign buffer_5_658 = $signed(_T_72566); // @[Modules.scala 53:83:@21748.4]
  assign _T_72568 = $signed(buffer_5_534) + $signed(buffer_5_535); // @[Modules.scala 53:83:@21750.4]
  assign _T_72569 = _T_72568[10:0]; // @[Modules.scala 53:83:@21751.4]
  assign buffer_5_659 = $signed(_T_72569); // @[Modules.scala 53:83:@21752.4]
  assign _T_72571 = $signed(buffer_5_536) + $signed(buffer_5_537); // @[Modules.scala 53:83:@21754.4]
  assign _T_72572 = _T_72571[10:0]; // @[Modules.scala 53:83:@21755.4]
  assign buffer_5_660 = $signed(_T_72572); // @[Modules.scala 53:83:@21756.4]
  assign _T_72574 = $signed(buffer_3_538) + $signed(buffer_4_539); // @[Modules.scala 53:83:@21758.4]
  assign _T_72575 = _T_72574[10:0]; // @[Modules.scala 53:83:@21759.4]
  assign buffer_5_661 = $signed(_T_72575); // @[Modules.scala 53:83:@21760.4]
  assign _T_72577 = $signed(buffer_1_540) + $signed(buffer_5_541); // @[Modules.scala 53:83:@21762.4]
  assign _T_72578 = _T_72577[10:0]; // @[Modules.scala 53:83:@21763.4]
  assign buffer_5_662 = $signed(_T_72578); // @[Modules.scala 53:83:@21764.4]
  assign _T_72580 = $signed(buffer_5_542) + $signed(buffer_5_543); // @[Modules.scala 53:83:@21766.4]
  assign _T_72581 = _T_72580[10:0]; // @[Modules.scala 53:83:@21767.4]
  assign buffer_5_663 = $signed(_T_72581); // @[Modules.scala 53:83:@21768.4]
  assign _T_72583 = $signed(buffer_2_544) + $signed(buffer_0_545); // @[Modules.scala 53:83:@21770.4]
  assign _T_72584 = _T_72583[10:0]; // @[Modules.scala 53:83:@21771.4]
  assign buffer_5_664 = $signed(_T_72584); // @[Modules.scala 53:83:@21772.4]
  assign _T_72586 = $signed(buffer_1_546) + $signed(buffer_4_547); // @[Modules.scala 53:83:@21774.4]
  assign _T_72587 = _T_72586[10:0]; // @[Modules.scala 53:83:@21775.4]
  assign buffer_5_665 = $signed(_T_72587); // @[Modules.scala 53:83:@21776.4]
  assign _T_72589 = $signed(buffer_5_548) + $signed(buffer_5_549); // @[Modules.scala 53:83:@21778.4]
  assign _T_72590 = _T_72589[10:0]; // @[Modules.scala 53:83:@21779.4]
  assign buffer_5_666 = $signed(_T_72590); // @[Modules.scala 53:83:@21780.4]
  assign _T_72592 = $signed(buffer_5_550) + $signed(buffer_0_551); // @[Modules.scala 53:83:@21782.4]
  assign _T_72593 = _T_72592[10:0]; // @[Modules.scala 53:83:@21783.4]
  assign buffer_5_667 = $signed(_T_72593); // @[Modules.scala 53:83:@21784.4]
  assign _T_72595 = $signed(buffer_5_552) + $signed(buffer_1_553); // @[Modules.scala 53:83:@21786.4]
  assign _T_72596 = _T_72595[10:0]; // @[Modules.scala 53:83:@21787.4]
  assign buffer_5_668 = $signed(_T_72596); // @[Modules.scala 53:83:@21788.4]
  assign _T_72598 = $signed(buffer_5_554) + $signed(buffer_5_555); // @[Modules.scala 53:83:@21790.4]
  assign _T_72599 = _T_72598[10:0]; // @[Modules.scala 53:83:@21791.4]
  assign buffer_5_669 = $signed(_T_72599); // @[Modules.scala 53:83:@21792.4]
  assign _T_72601 = $signed(buffer_5_556) + $signed(buffer_5_557); // @[Modules.scala 53:83:@21794.4]
  assign _T_72602 = _T_72601[10:0]; // @[Modules.scala 53:83:@21795.4]
  assign buffer_5_670 = $signed(_T_72602); // @[Modules.scala 53:83:@21796.4]
  assign _T_72604 = $signed(buffer_5_558) + $signed(buffer_0_559); // @[Modules.scala 53:83:@21798.4]
  assign _T_72605 = _T_72604[10:0]; // @[Modules.scala 53:83:@21799.4]
  assign buffer_5_671 = $signed(_T_72605); // @[Modules.scala 53:83:@21800.4]
  assign _T_72607 = $signed(buffer_5_560) + $signed(buffer_5_561); // @[Modules.scala 53:83:@21802.4]
  assign _T_72608 = _T_72607[10:0]; // @[Modules.scala 53:83:@21803.4]
  assign buffer_5_672 = $signed(_T_72608); // @[Modules.scala 53:83:@21804.4]
  assign _T_72610 = $signed(buffer_5_562) + $signed(buffer_5_563); // @[Modules.scala 53:83:@21806.4]
  assign _T_72611 = _T_72610[10:0]; // @[Modules.scala 53:83:@21807.4]
  assign buffer_5_673 = $signed(_T_72611); // @[Modules.scala 53:83:@21808.4]
  assign _T_72616 = $signed(buffer_5_566) + $signed(buffer_5_567); // @[Modules.scala 53:83:@21814.4]
  assign _T_72617 = _T_72616[10:0]; // @[Modules.scala 53:83:@21815.4]
  assign buffer_5_675 = $signed(_T_72617); // @[Modules.scala 53:83:@21816.4]
  assign _T_72619 = $signed(buffer_5_568) + $signed(buffer_3_569); // @[Modules.scala 53:83:@21818.4]
  assign _T_72620 = _T_72619[10:0]; // @[Modules.scala 53:83:@21819.4]
  assign buffer_5_676 = $signed(_T_72620); // @[Modules.scala 53:83:@21820.4]
  assign _T_72625 = $signed(buffer_5_572) + $signed(buffer_0_573); // @[Modules.scala 53:83:@21826.4]
  assign _T_72626 = _T_72625[10:0]; // @[Modules.scala 53:83:@21827.4]
  assign buffer_5_678 = $signed(_T_72626); // @[Modules.scala 53:83:@21828.4]
  assign _T_72628 = $signed(buffer_2_574) + $signed(buffer_5_575); // @[Modules.scala 53:83:@21830.4]
  assign _T_72629 = _T_72628[10:0]; // @[Modules.scala 53:83:@21831.4]
  assign buffer_5_679 = $signed(_T_72629); // @[Modules.scala 53:83:@21832.4]
  assign _T_72631 = $signed(buffer_3_576) + $signed(buffer_5_577); // @[Modules.scala 53:83:@21834.4]
  assign _T_72632 = _T_72631[10:0]; // @[Modules.scala 53:83:@21835.4]
  assign buffer_5_680 = $signed(_T_72632); // @[Modules.scala 53:83:@21836.4]
  assign _T_72634 = $signed(buffer_3_578) + $signed(buffer_5_579); // @[Modules.scala 53:83:@21838.4]
  assign _T_72635 = _T_72634[10:0]; // @[Modules.scala 53:83:@21839.4]
  assign buffer_5_681 = $signed(_T_72635); // @[Modules.scala 53:83:@21840.4]
  assign _T_72637 = $signed(buffer_3_580) + $signed(buffer_1_581); // @[Modules.scala 53:83:@21842.4]
  assign _T_72638 = _T_72637[10:0]; // @[Modules.scala 53:83:@21843.4]
  assign buffer_5_682 = $signed(_T_72638); // @[Modules.scala 53:83:@21844.4]
  assign _T_72640 = $signed(buffer_5_582) + $signed(buffer_5_583); // @[Modules.scala 53:83:@21846.4]
  assign _T_72641 = _T_72640[10:0]; // @[Modules.scala 53:83:@21847.4]
  assign buffer_5_683 = $signed(_T_72641); // @[Modules.scala 53:83:@21848.4]
  assign _T_72646 = $signed(buffer_5_586) + $signed(buffer_3_587); // @[Modules.scala 53:83:@21854.4]
  assign _T_72647 = _T_72646[10:0]; // @[Modules.scala 53:83:@21855.4]
  assign buffer_5_685 = $signed(_T_72647); // @[Modules.scala 53:83:@21856.4]
  assign _T_72649 = $signed(buffer_5_588) + $signed(buffer_5_589); // @[Modules.scala 56:109:@21858.4]
  assign _T_72650 = _T_72649[10:0]; // @[Modules.scala 56:109:@21859.4]
  assign buffer_5_686 = $signed(_T_72650); // @[Modules.scala 56:109:@21860.4]
  assign _T_72652 = $signed(buffer_5_590) + $signed(buffer_5_591); // @[Modules.scala 56:109:@21862.4]
  assign _T_72653 = _T_72652[10:0]; // @[Modules.scala 56:109:@21863.4]
  assign buffer_5_687 = $signed(_T_72653); // @[Modules.scala 56:109:@21864.4]
  assign _T_72655 = $signed(buffer_5_592) + $signed(buffer_5_593); // @[Modules.scala 56:109:@21866.4]
  assign _T_72656 = _T_72655[10:0]; // @[Modules.scala 56:109:@21867.4]
  assign buffer_5_688 = $signed(_T_72656); // @[Modules.scala 56:109:@21868.4]
  assign _T_72658 = $signed(buffer_5_594) + $signed(buffer_5_595); // @[Modules.scala 56:109:@21870.4]
  assign _T_72659 = _T_72658[10:0]; // @[Modules.scala 56:109:@21871.4]
  assign buffer_5_689 = $signed(_T_72659); // @[Modules.scala 56:109:@21872.4]
  assign _T_72661 = $signed(buffer_5_596) + $signed(buffer_5_597); // @[Modules.scala 56:109:@21874.4]
  assign _T_72662 = _T_72661[10:0]; // @[Modules.scala 56:109:@21875.4]
  assign buffer_5_690 = $signed(_T_72662); // @[Modules.scala 56:109:@21876.4]
  assign _T_72664 = $signed(buffer_5_598) + $signed(buffer_0_599); // @[Modules.scala 56:109:@21878.4]
  assign _T_72665 = _T_72664[10:0]; // @[Modules.scala 56:109:@21879.4]
  assign buffer_5_691 = $signed(_T_72665); // @[Modules.scala 56:109:@21880.4]
  assign _T_72667 = $signed(buffer_5_600) + $signed(buffer_5_601); // @[Modules.scala 56:109:@21882.4]
  assign _T_72668 = _T_72667[10:0]; // @[Modules.scala 56:109:@21883.4]
  assign buffer_5_692 = $signed(_T_72668); // @[Modules.scala 56:109:@21884.4]
  assign _T_72670 = $signed(buffer_5_602) + $signed(buffer_3_603); // @[Modules.scala 56:109:@21886.4]
  assign _T_72671 = _T_72670[10:0]; // @[Modules.scala 56:109:@21887.4]
  assign buffer_5_693 = $signed(_T_72671); // @[Modules.scala 56:109:@21888.4]
  assign _T_72673 = $signed(buffer_5_604) + $signed(buffer_5_605); // @[Modules.scala 56:109:@21890.4]
  assign _T_72674 = _T_72673[10:0]; // @[Modules.scala 56:109:@21891.4]
  assign buffer_5_694 = $signed(_T_72674); // @[Modules.scala 56:109:@21892.4]
  assign _T_72676 = $signed(buffer_5_606) + $signed(buffer_5_607); // @[Modules.scala 56:109:@21894.4]
  assign _T_72677 = _T_72676[10:0]; // @[Modules.scala 56:109:@21895.4]
  assign buffer_5_695 = $signed(_T_72677); // @[Modules.scala 56:109:@21896.4]
  assign _T_72679 = $signed(buffer_5_608) + $signed(buffer_5_609); // @[Modules.scala 56:109:@21898.4]
  assign _T_72680 = _T_72679[10:0]; // @[Modules.scala 56:109:@21899.4]
  assign buffer_5_696 = $signed(_T_72680); // @[Modules.scala 56:109:@21900.4]
  assign _T_72682 = $signed(buffer_5_610) + $signed(buffer_5_611); // @[Modules.scala 56:109:@21902.4]
  assign _T_72683 = _T_72682[10:0]; // @[Modules.scala 56:109:@21903.4]
  assign buffer_5_697 = $signed(_T_72683); // @[Modules.scala 56:109:@21904.4]
  assign _T_72685 = $signed(buffer_5_612) + $signed(buffer_5_613); // @[Modules.scala 56:109:@21906.4]
  assign _T_72686 = _T_72685[10:0]; // @[Modules.scala 56:109:@21907.4]
  assign buffer_5_698 = $signed(_T_72686); // @[Modules.scala 56:109:@21908.4]
  assign _T_72688 = $signed(buffer_5_614) + $signed(buffer_5_615); // @[Modules.scala 56:109:@21910.4]
  assign _T_72689 = _T_72688[10:0]; // @[Modules.scala 56:109:@21911.4]
  assign buffer_5_699 = $signed(_T_72689); // @[Modules.scala 56:109:@21912.4]
  assign _T_72691 = $signed(buffer_5_616) + $signed(buffer_5_617); // @[Modules.scala 56:109:@21914.4]
  assign _T_72692 = _T_72691[10:0]; // @[Modules.scala 56:109:@21915.4]
  assign buffer_5_700 = $signed(_T_72692); // @[Modules.scala 56:109:@21916.4]
  assign _T_72694 = $signed(buffer_5_618) + $signed(buffer_5_619); // @[Modules.scala 56:109:@21918.4]
  assign _T_72695 = _T_72694[10:0]; // @[Modules.scala 56:109:@21919.4]
  assign buffer_5_701 = $signed(_T_72695); // @[Modules.scala 56:109:@21920.4]
  assign _T_72697 = $signed(buffer_5_620) + $signed(buffer_5_621); // @[Modules.scala 56:109:@21922.4]
  assign _T_72698 = _T_72697[10:0]; // @[Modules.scala 56:109:@21923.4]
  assign buffer_5_702 = $signed(_T_72698); // @[Modules.scala 56:109:@21924.4]
  assign _T_72700 = $signed(buffer_5_622) + $signed(buffer_5_623); // @[Modules.scala 56:109:@21926.4]
  assign _T_72701 = _T_72700[10:0]; // @[Modules.scala 56:109:@21927.4]
  assign buffer_5_703 = $signed(_T_72701); // @[Modules.scala 56:109:@21928.4]
  assign _T_72703 = $signed(buffer_5_624) + $signed(buffer_5_625); // @[Modules.scala 56:109:@21930.4]
  assign _T_72704 = _T_72703[10:0]; // @[Modules.scala 56:109:@21931.4]
  assign buffer_5_704 = $signed(_T_72704); // @[Modules.scala 56:109:@21932.4]
  assign _T_72706 = $signed(buffer_5_626) + $signed(buffer_3_627); // @[Modules.scala 56:109:@21934.4]
  assign _T_72707 = _T_72706[10:0]; // @[Modules.scala 56:109:@21935.4]
  assign buffer_5_705 = $signed(_T_72707); // @[Modules.scala 56:109:@21936.4]
  assign _T_72709 = $signed(buffer_5_628) + $signed(buffer_5_629); // @[Modules.scala 56:109:@21938.4]
  assign _T_72710 = _T_72709[10:0]; // @[Modules.scala 56:109:@21939.4]
  assign buffer_5_706 = $signed(_T_72710); // @[Modules.scala 56:109:@21940.4]
  assign _T_72712 = $signed(buffer_5_630) + $signed(buffer_5_631); // @[Modules.scala 56:109:@21942.4]
  assign _T_72713 = _T_72712[10:0]; // @[Modules.scala 56:109:@21943.4]
  assign buffer_5_707 = $signed(_T_72713); // @[Modules.scala 56:109:@21944.4]
  assign _T_72715 = $signed(buffer_5_632) + $signed(buffer_5_633); // @[Modules.scala 56:109:@21946.4]
  assign _T_72716 = _T_72715[10:0]; // @[Modules.scala 56:109:@21947.4]
  assign buffer_5_708 = $signed(_T_72716); // @[Modules.scala 56:109:@21948.4]
  assign _T_72718 = $signed(buffer_5_634) + $signed(buffer_5_635); // @[Modules.scala 56:109:@21950.4]
  assign _T_72719 = _T_72718[10:0]; // @[Modules.scala 56:109:@21951.4]
  assign buffer_5_709 = $signed(_T_72719); // @[Modules.scala 56:109:@21952.4]
  assign _T_72721 = $signed(buffer_5_636) + $signed(buffer_5_637); // @[Modules.scala 56:109:@21954.4]
  assign _T_72722 = _T_72721[10:0]; // @[Modules.scala 56:109:@21955.4]
  assign buffer_5_710 = $signed(_T_72722); // @[Modules.scala 56:109:@21956.4]
  assign _T_72724 = $signed(buffer_5_638) + $signed(buffer_5_639); // @[Modules.scala 56:109:@21958.4]
  assign _T_72725 = _T_72724[10:0]; // @[Modules.scala 56:109:@21959.4]
  assign buffer_5_711 = $signed(_T_72725); // @[Modules.scala 56:109:@21960.4]
  assign _T_72727 = $signed(buffer_5_640) + $signed(buffer_5_641); // @[Modules.scala 56:109:@21962.4]
  assign _T_72728 = _T_72727[10:0]; // @[Modules.scala 56:109:@21963.4]
  assign buffer_5_712 = $signed(_T_72728); // @[Modules.scala 56:109:@21964.4]
  assign _T_72730 = $signed(buffer_5_642) + $signed(buffer_5_643); // @[Modules.scala 56:109:@21966.4]
  assign _T_72731 = _T_72730[10:0]; // @[Modules.scala 56:109:@21967.4]
  assign buffer_5_713 = $signed(_T_72731); // @[Modules.scala 56:109:@21968.4]
  assign _T_72733 = $signed(buffer_5_644) + $signed(buffer_5_645); // @[Modules.scala 56:109:@21970.4]
  assign _T_72734 = _T_72733[10:0]; // @[Modules.scala 56:109:@21971.4]
  assign buffer_5_714 = $signed(_T_72734); // @[Modules.scala 56:109:@21972.4]
  assign _T_72736 = $signed(buffer_5_646) + $signed(buffer_5_647); // @[Modules.scala 56:109:@21974.4]
  assign _T_72737 = _T_72736[10:0]; // @[Modules.scala 56:109:@21975.4]
  assign buffer_5_715 = $signed(_T_72737); // @[Modules.scala 56:109:@21976.4]
  assign _T_72739 = $signed(buffer_5_648) + $signed(buffer_5_649); // @[Modules.scala 56:109:@21978.4]
  assign _T_72740 = _T_72739[10:0]; // @[Modules.scala 56:109:@21979.4]
  assign buffer_5_716 = $signed(_T_72740); // @[Modules.scala 56:109:@21980.4]
  assign _T_72742 = $signed(buffer_5_650) + $signed(buffer_5_651); // @[Modules.scala 56:109:@21982.4]
  assign _T_72743 = _T_72742[10:0]; // @[Modules.scala 56:109:@21983.4]
  assign buffer_5_717 = $signed(_T_72743); // @[Modules.scala 56:109:@21984.4]
  assign _T_72745 = $signed(buffer_5_652) + $signed(buffer_5_653); // @[Modules.scala 56:109:@21986.4]
  assign _T_72746 = _T_72745[10:0]; // @[Modules.scala 56:109:@21987.4]
  assign buffer_5_718 = $signed(_T_72746); // @[Modules.scala 56:109:@21988.4]
  assign _T_72748 = $signed(buffer_5_654) + $signed(buffer_5_655); // @[Modules.scala 56:109:@21990.4]
  assign _T_72749 = _T_72748[10:0]; // @[Modules.scala 56:109:@21991.4]
  assign buffer_5_719 = $signed(_T_72749); // @[Modules.scala 56:109:@21992.4]
  assign _T_72751 = $signed(buffer_5_656) + $signed(buffer_5_657); // @[Modules.scala 56:109:@21994.4]
  assign _T_72752 = _T_72751[10:0]; // @[Modules.scala 56:109:@21995.4]
  assign buffer_5_720 = $signed(_T_72752); // @[Modules.scala 56:109:@21996.4]
  assign _T_72754 = $signed(buffer_5_658) + $signed(buffer_5_659); // @[Modules.scala 56:109:@21998.4]
  assign _T_72755 = _T_72754[10:0]; // @[Modules.scala 56:109:@21999.4]
  assign buffer_5_721 = $signed(_T_72755); // @[Modules.scala 56:109:@22000.4]
  assign _T_72757 = $signed(buffer_5_660) + $signed(buffer_5_661); // @[Modules.scala 56:109:@22002.4]
  assign _T_72758 = _T_72757[10:0]; // @[Modules.scala 56:109:@22003.4]
  assign buffer_5_722 = $signed(_T_72758); // @[Modules.scala 56:109:@22004.4]
  assign _T_72760 = $signed(buffer_5_662) + $signed(buffer_5_663); // @[Modules.scala 56:109:@22006.4]
  assign _T_72761 = _T_72760[10:0]; // @[Modules.scala 56:109:@22007.4]
  assign buffer_5_723 = $signed(_T_72761); // @[Modules.scala 56:109:@22008.4]
  assign _T_72763 = $signed(buffer_5_664) + $signed(buffer_5_665); // @[Modules.scala 56:109:@22010.4]
  assign _T_72764 = _T_72763[10:0]; // @[Modules.scala 56:109:@22011.4]
  assign buffer_5_724 = $signed(_T_72764); // @[Modules.scala 56:109:@22012.4]
  assign _T_72766 = $signed(buffer_5_666) + $signed(buffer_5_667); // @[Modules.scala 56:109:@22014.4]
  assign _T_72767 = _T_72766[10:0]; // @[Modules.scala 56:109:@22015.4]
  assign buffer_5_725 = $signed(_T_72767); // @[Modules.scala 56:109:@22016.4]
  assign _T_72769 = $signed(buffer_5_668) + $signed(buffer_5_669); // @[Modules.scala 56:109:@22018.4]
  assign _T_72770 = _T_72769[10:0]; // @[Modules.scala 56:109:@22019.4]
  assign buffer_5_726 = $signed(_T_72770); // @[Modules.scala 56:109:@22020.4]
  assign _T_72772 = $signed(buffer_5_670) + $signed(buffer_5_671); // @[Modules.scala 56:109:@22022.4]
  assign _T_72773 = _T_72772[10:0]; // @[Modules.scala 56:109:@22023.4]
  assign buffer_5_727 = $signed(_T_72773); // @[Modules.scala 56:109:@22024.4]
  assign _T_72775 = $signed(buffer_5_672) + $signed(buffer_5_673); // @[Modules.scala 56:109:@22026.4]
  assign _T_72776 = _T_72775[10:0]; // @[Modules.scala 56:109:@22027.4]
  assign buffer_5_728 = $signed(_T_72776); // @[Modules.scala 56:109:@22028.4]
  assign _T_72778 = $signed(buffer_0_674) + $signed(buffer_5_675); // @[Modules.scala 56:109:@22030.4]
  assign _T_72779 = _T_72778[10:0]; // @[Modules.scala 56:109:@22031.4]
  assign buffer_5_729 = $signed(_T_72779); // @[Modules.scala 56:109:@22032.4]
  assign _T_72781 = $signed(buffer_5_676) + $signed(buffer_0_677); // @[Modules.scala 56:109:@22034.4]
  assign _T_72782 = _T_72781[10:0]; // @[Modules.scala 56:109:@22035.4]
  assign buffer_5_730 = $signed(_T_72782); // @[Modules.scala 56:109:@22036.4]
  assign _T_72784 = $signed(buffer_5_678) + $signed(buffer_5_679); // @[Modules.scala 56:109:@22038.4]
  assign _T_72785 = _T_72784[10:0]; // @[Modules.scala 56:109:@22039.4]
  assign buffer_5_731 = $signed(_T_72785); // @[Modules.scala 56:109:@22040.4]
  assign _T_72787 = $signed(buffer_5_680) + $signed(buffer_5_681); // @[Modules.scala 56:109:@22042.4]
  assign _T_72788 = _T_72787[10:0]; // @[Modules.scala 56:109:@22043.4]
  assign buffer_5_732 = $signed(_T_72788); // @[Modules.scala 56:109:@22044.4]
  assign _T_72790 = $signed(buffer_5_682) + $signed(buffer_5_683); // @[Modules.scala 56:109:@22046.4]
  assign _T_72791 = _T_72790[10:0]; // @[Modules.scala 56:109:@22047.4]
  assign buffer_5_733 = $signed(_T_72791); // @[Modules.scala 56:109:@22048.4]
  assign _T_72793 = $signed(buffer_3_684) + $signed(buffer_5_685); // @[Modules.scala 56:109:@22050.4]
  assign _T_72794 = _T_72793[10:0]; // @[Modules.scala 56:109:@22051.4]
  assign buffer_5_734 = $signed(_T_72794); // @[Modules.scala 56:109:@22052.4]
  assign _T_72796 = $signed(buffer_5_686) + $signed(buffer_5_687); // @[Modules.scala 63:156:@22055.4]
  assign _T_72797 = _T_72796[10:0]; // @[Modules.scala 63:156:@22056.4]
  assign buffer_5_736 = $signed(_T_72797); // @[Modules.scala 63:156:@22057.4]
  assign _T_72799 = $signed(buffer_5_736) + $signed(buffer_5_688); // @[Modules.scala 63:156:@22059.4]
  assign _T_72800 = _T_72799[10:0]; // @[Modules.scala 63:156:@22060.4]
  assign buffer_5_737 = $signed(_T_72800); // @[Modules.scala 63:156:@22061.4]
  assign _T_72802 = $signed(buffer_5_737) + $signed(buffer_5_689); // @[Modules.scala 63:156:@22063.4]
  assign _T_72803 = _T_72802[10:0]; // @[Modules.scala 63:156:@22064.4]
  assign buffer_5_738 = $signed(_T_72803); // @[Modules.scala 63:156:@22065.4]
  assign _T_72805 = $signed(buffer_5_738) + $signed(buffer_5_690); // @[Modules.scala 63:156:@22067.4]
  assign _T_72806 = _T_72805[10:0]; // @[Modules.scala 63:156:@22068.4]
  assign buffer_5_739 = $signed(_T_72806); // @[Modules.scala 63:156:@22069.4]
  assign _T_72808 = $signed(buffer_5_739) + $signed(buffer_5_691); // @[Modules.scala 63:156:@22071.4]
  assign _T_72809 = _T_72808[10:0]; // @[Modules.scala 63:156:@22072.4]
  assign buffer_5_740 = $signed(_T_72809); // @[Modules.scala 63:156:@22073.4]
  assign _T_72811 = $signed(buffer_5_740) + $signed(buffer_5_692); // @[Modules.scala 63:156:@22075.4]
  assign _T_72812 = _T_72811[10:0]; // @[Modules.scala 63:156:@22076.4]
  assign buffer_5_741 = $signed(_T_72812); // @[Modules.scala 63:156:@22077.4]
  assign _T_72814 = $signed(buffer_5_741) + $signed(buffer_5_693); // @[Modules.scala 63:156:@22079.4]
  assign _T_72815 = _T_72814[10:0]; // @[Modules.scala 63:156:@22080.4]
  assign buffer_5_742 = $signed(_T_72815); // @[Modules.scala 63:156:@22081.4]
  assign _T_72817 = $signed(buffer_5_742) + $signed(buffer_5_694); // @[Modules.scala 63:156:@22083.4]
  assign _T_72818 = _T_72817[10:0]; // @[Modules.scala 63:156:@22084.4]
  assign buffer_5_743 = $signed(_T_72818); // @[Modules.scala 63:156:@22085.4]
  assign _T_72820 = $signed(buffer_5_743) + $signed(buffer_5_695); // @[Modules.scala 63:156:@22087.4]
  assign _T_72821 = _T_72820[10:0]; // @[Modules.scala 63:156:@22088.4]
  assign buffer_5_744 = $signed(_T_72821); // @[Modules.scala 63:156:@22089.4]
  assign _T_72823 = $signed(buffer_5_744) + $signed(buffer_5_696); // @[Modules.scala 63:156:@22091.4]
  assign _T_72824 = _T_72823[10:0]; // @[Modules.scala 63:156:@22092.4]
  assign buffer_5_745 = $signed(_T_72824); // @[Modules.scala 63:156:@22093.4]
  assign _T_72826 = $signed(buffer_5_745) + $signed(buffer_5_697); // @[Modules.scala 63:156:@22095.4]
  assign _T_72827 = _T_72826[10:0]; // @[Modules.scala 63:156:@22096.4]
  assign buffer_5_746 = $signed(_T_72827); // @[Modules.scala 63:156:@22097.4]
  assign _T_72829 = $signed(buffer_5_746) + $signed(buffer_5_698); // @[Modules.scala 63:156:@22099.4]
  assign _T_72830 = _T_72829[10:0]; // @[Modules.scala 63:156:@22100.4]
  assign buffer_5_747 = $signed(_T_72830); // @[Modules.scala 63:156:@22101.4]
  assign _T_72832 = $signed(buffer_5_747) + $signed(buffer_5_699); // @[Modules.scala 63:156:@22103.4]
  assign _T_72833 = _T_72832[10:0]; // @[Modules.scala 63:156:@22104.4]
  assign buffer_5_748 = $signed(_T_72833); // @[Modules.scala 63:156:@22105.4]
  assign _T_72835 = $signed(buffer_5_748) + $signed(buffer_5_700); // @[Modules.scala 63:156:@22107.4]
  assign _T_72836 = _T_72835[10:0]; // @[Modules.scala 63:156:@22108.4]
  assign buffer_5_749 = $signed(_T_72836); // @[Modules.scala 63:156:@22109.4]
  assign _T_72838 = $signed(buffer_5_749) + $signed(buffer_5_701); // @[Modules.scala 63:156:@22111.4]
  assign _T_72839 = _T_72838[10:0]; // @[Modules.scala 63:156:@22112.4]
  assign buffer_5_750 = $signed(_T_72839); // @[Modules.scala 63:156:@22113.4]
  assign _T_72841 = $signed(buffer_5_750) + $signed(buffer_5_702); // @[Modules.scala 63:156:@22115.4]
  assign _T_72842 = _T_72841[10:0]; // @[Modules.scala 63:156:@22116.4]
  assign buffer_5_751 = $signed(_T_72842); // @[Modules.scala 63:156:@22117.4]
  assign _T_72844 = $signed(buffer_5_751) + $signed(buffer_5_703); // @[Modules.scala 63:156:@22119.4]
  assign _T_72845 = _T_72844[10:0]; // @[Modules.scala 63:156:@22120.4]
  assign buffer_5_752 = $signed(_T_72845); // @[Modules.scala 63:156:@22121.4]
  assign _T_72847 = $signed(buffer_5_752) + $signed(buffer_5_704); // @[Modules.scala 63:156:@22123.4]
  assign _T_72848 = _T_72847[10:0]; // @[Modules.scala 63:156:@22124.4]
  assign buffer_5_753 = $signed(_T_72848); // @[Modules.scala 63:156:@22125.4]
  assign _T_72850 = $signed(buffer_5_753) + $signed(buffer_5_705); // @[Modules.scala 63:156:@22127.4]
  assign _T_72851 = _T_72850[10:0]; // @[Modules.scala 63:156:@22128.4]
  assign buffer_5_754 = $signed(_T_72851); // @[Modules.scala 63:156:@22129.4]
  assign _T_72853 = $signed(buffer_5_754) + $signed(buffer_5_706); // @[Modules.scala 63:156:@22131.4]
  assign _T_72854 = _T_72853[10:0]; // @[Modules.scala 63:156:@22132.4]
  assign buffer_5_755 = $signed(_T_72854); // @[Modules.scala 63:156:@22133.4]
  assign _T_72856 = $signed(buffer_5_755) + $signed(buffer_5_707); // @[Modules.scala 63:156:@22135.4]
  assign _T_72857 = _T_72856[10:0]; // @[Modules.scala 63:156:@22136.4]
  assign buffer_5_756 = $signed(_T_72857); // @[Modules.scala 63:156:@22137.4]
  assign _T_72859 = $signed(buffer_5_756) + $signed(buffer_5_708); // @[Modules.scala 63:156:@22139.4]
  assign _T_72860 = _T_72859[10:0]; // @[Modules.scala 63:156:@22140.4]
  assign buffer_5_757 = $signed(_T_72860); // @[Modules.scala 63:156:@22141.4]
  assign _T_72862 = $signed(buffer_5_757) + $signed(buffer_5_709); // @[Modules.scala 63:156:@22143.4]
  assign _T_72863 = _T_72862[10:0]; // @[Modules.scala 63:156:@22144.4]
  assign buffer_5_758 = $signed(_T_72863); // @[Modules.scala 63:156:@22145.4]
  assign _T_72865 = $signed(buffer_5_758) + $signed(buffer_5_710); // @[Modules.scala 63:156:@22147.4]
  assign _T_72866 = _T_72865[10:0]; // @[Modules.scala 63:156:@22148.4]
  assign buffer_5_759 = $signed(_T_72866); // @[Modules.scala 63:156:@22149.4]
  assign _T_72868 = $signed(buffer_5_759) + $signed(buffer_5_711); // @[Modules.scala 63:156:@22151.4]
  assign _T_72869 = _T_72868[10:0]; // @[Modules.scala 63:156:@22152.4]
  assign buffer_5_760 = $signed(_T_72869); // @[Modules.scala 63:156:@22153.4]
  assign _T_72871 = $signed(buffer_5_760) + $signed(buffer_5_712); // @[Modules.scala 63:156:@22155.4]
  assign _T_72872 = _T_72871[10:0]; // @[Modules.scala 63:156:@22156.4]
  assign buffer_5_761 = $signed(_T_72872); // @[Modules.scala 63:156:@22157.4]
  assign _T_72874 = $signed(buffer_5_761) + $signed(buffer_5_713); // @[Modules.scala 63:156:@22159.4]
  assign _T_72875 = _T_72874[10:0]; // @[Modules.scala 63:156:@22160.4]
  assign buffer_5_762 = $signed(_T_72875); // @[Modules.scala 63:156:@22161.4]
  assign _T_72877 = $signed(buffer_5_762) + $signed(buffer_5_714); // @[Modules.scala 63:156:@22163.4]
  assign _T_72878 = _T_72877[10:0]; // @[Modules.scala 63:156:@22164.4]
  assign buffer_5_763 = $signed(_T_72878); // @[Modules.scala 63:156:@22165.4]
  assign _T_72880 = $signed(buffer_5_763) + $signed(buffer_5_715); // @[Modules.scala 63:156:@22167.4]
  assign _T_72881 = _T_72880[10:0]; // @[Modules.scala 63:156:@22168.4]
  assign buffer_5_764 = $signed(_T_72881); // @[Modules.scala 63:156:@22169.4]
  assign _T_72883 = $signed(buffer_5_764) + $signed(buffer_5_716); // @[Modules.scala 63:156:@22171.4]
  assign _T_72884 = _T_72883[10:0]; // @[Modules.scala 63:156:@22172.4]
  assign buffer_5_765 = $signed(_T_72884); // @[Modules.scala 63:156:@22173.4]
  assign _T_72886 = $signed(buffer_5_765) + $signed(buffer_5_717); // @[Modules.scala 63:156:@22175.4]
  assign _T_72887 = _T_72886[10:0]; // @[Modules.scala 63:156:@22176.4]
  assign buffer_5_766 = $signed(_T_72887); // @[Modules.scala 63:156:@22177.4]
  assign _T_72889 = $signed(buffer_5_766) + $signed(buffer_5_718); // @[Modules.scala 63:156:@22179.4]
  assign _T_72890 = _T_72889[10:0]; // @[Modules.scala 63:156:@22180.4]
  assign buffer_5_767 = $signed(_T_72890); // @[Modules.scala 63:156:@22181.4]
  assign _T_72892 = $signed(buffer_5_767) + $signed(buffer_5_719); // @[Modules.scala 63:156:@22183.4]
  assign _T_72893 = _T_72892[10:0]; // @[Modules.scala 63:156:@22184.4]
  assign buffer_5_768 = $signed(_T_72893); // @[Modules.scala 63:156:@22185.4]
  assign _T_72895 = $signed(buffer_5_768) + $signed(buffer_5_720); // @[Modules.scala 63:156:@22187.4]
  assign _T_72896 = _T_72895[10:0]; // @[Modules.scala 63:156:@22188.4]
  assign buffer_5_769 = $signed(_T_72896); // @[Modules.scala 63:156:@22189.4]
  assign _T_72898 = $signed(buffer_5_769) + $signed(buffer_5_721); // @[Modules.scala 63:156:@22191.4]
  assign _T_72899 = _T_72898[10:0]; // @[Modules.scala 63:156:@22192.4]
  assign buffer_5_770 = $signed(_T_72899); // @[Modules.scala 63:156:@22193.4]
  assign _T_72901 = $signed(buffer_5_770) + $signed(buffer_5_722); // @[Modules.scala 63:156:@22195.4]
  assign _T_72902 = _T_72901[10:0]; // @[Modules.scala 63:156:@22196.4]
  assign buffer_5_771 = $signed(_T_72902); // @[Modules.scala 63:156:@22197.4]
  assign _T_72904 = $signed(buffer_5_771) + $signed(buffer_5_723); // @[Modules.scala 63:156:@22199.4]
  assign _T_72905 = _T_72904[10:0]; // @[Modules.scala 63:156:@22200.4]
  assign buffer_5_772 = $signed(_T_72905); // @[Modules.scala 63:156:@22201.4]
  assign _T_72907 = $signed(buffer_5_772) + $signed(buffer_5_724); // @[Modules.scala 63:156:@22203.4]
  assign _T_72908 = _T_72907[10:0]; // @[Modules.scala 63:156:@22204.4]
  assign buffer_5_773 = $signed(_T_72908); // @[Modules.scala 63:156:@22205.4]
  assign _T_72910 = $signed(buffer_5_773) + $signed(buffer_5_725); // @[Modules.scala 63:156:@22207.4]
  assign _T_72911 = _T_72910[10:0]; // @[Modules.scala 63:156:@22208.4]
  assign buffer_5_774 = $signed(_T_72911); // @[Modules.scala 63:156:@22209.4]
  assign _T_72913 = $signed(buffer_5_774) + $signed(buffer_5_726); // @[Modules.scala 63:156:@22211.4]
  assign _T_72914 = _T_72913[10:0]; // @[Modules.scala 63:156:@22212.4]
  assign buffer_5_775 = $signed(_T_72914); // @[Modules.scala 63:156:@22213.4]
  assign _T_72916 = $signed(buffer_5_775) + $signed(buffer_5_727); // @[Modules.scala 63:156:@22215.4]
  assign _T_72917 = _T_72916[10:0]; // @[Modules.scala 63:156:@22216.4]
  assign buffer_5_776 = $signed(_T_72917); // @[Modules.scala 63:156:@22217.4]
  assign _T_72919 = $signed(buffer_5_776) + $signed(buffer_5_728); // @[Modules.scala 63:156:@22219.4]
  assign _T_72920 = _T_72919[10:0]; // @[Modules.scala 63:156:@22220.4]
  assign buffer_5_777 = $signed(_T_72920); // @[Modules.scala 63:156:@22221.4]
  assign _T_72922 = $signed(buffer_5_777) + $signed(buffer_5_729); // @[Modules.scala 63:156:@22223.4]
  assign _T_72923 = _T_72922[10:0]; // @[Modules.scala 63:156:@22224.4]
  assign buffer_5_778 = $signed(_T_72923); // @[Modules.scala 63:156:@22225.4]
  assign _T_72925 = $signed(buffer_5_778) + $signed(buffer_5_730); // @[Modules.scala 63:156:@22227.4]
  assign _T_72926 = _T_72925[10:0]; // @[Modules.scala 63:156:@22228.4]
  assign buffer_5_779 = $signed(_T_72926); // @[Modules.scala 63:156:@22229.4]
  assign _T_72928 = $signed(buffer_5_779) + $signed(buffer_5_731); // @[Modules.scala 63:156:@22231.4]
  assign _T_72929 = _T_72928[10:0]; // @[Modules.scala 63:156:@22232.4]
  assign buffer_5_780 = $signed(_T_72929); // @[Modules.scala 63:156:@22233.4]
  assign _T_72931 = $signed(buffer_5_780) + $signed(buffer_5_732); // @[Modules.scala 63:156:@22235.4]
  assign _T_72932 = _T_72931[10:0]; // @[Modules.scala 63:156:@22236.4]
  assign buffer_5_781 = $signed(_T_72932); // @[Modules.scala 63:156:@22237.4]
  assign _T_72934 = $signed(buffer_5_781) + $signed(buffer_5_733); // @[Modules.scala 63:156:@22239.4]
  assign _T_72935 = _T_72934[10:0]; // @[Modules.scala 63:156:@22240.4]
  assign buffer_5_782 = $signed(_T_72935); // @[Modules.scala 63:156:@22241.4]
  assign _T_72937 = $signed(buffer_5_782) + $signed(buffer_5_734); // @[Modules.scala 63:156:@22243.4]
  assign _T_72938 = _T_72937[10:0]; // @[Modules.scala 63:156:@22244.4]
  assign buffer_5_783 = $signed(_T_72938); // @[Modules.scala 63:156:@22245.4]
  assign _T_73239 = $signed(5'sh0) - $signed(io_in_100); // @[Modules.scala 46:37:@22559.4]
  assign _T_73240 = _T_73239[4:0]; // @[Modules.scala 46:37:@22560.4]
  assign _T_73241 = $signed(_T_73240); // @[Modules.scala 46:37:@22561.4]
  assign _T_73242 = $signed(_T_73241) - $signed(io_in_101); // @[Modules.scala 46:47:@22562.4]
  assign _T_73243 = _T_73242[4:0]; // @[Modules.scala 46:47:@22563.4]
  assign _T_73244 = $signed(_T_73243); // @[Modules.scala 46:47:@22564.4]
  assign _T_73259 = $signed(io_in_106) - $signed(io_in_107); // @[Modules.scala 40:46:@22580.4]
  assign _T_73260 = _T_73259[4:0]; // @[Modules.scala 40:46:@22581.4]
  assign _T_73261 = $signed(_T_73260); // @[Modules.scala 40:46:@22582.4]
  assign _T_73328 = $signed(_T_54625) - $signed(io_in_129); // @[Modules.scala 46:47:@22651.4]
  assign _T_73329 = _T_73328[4:0]; // @[Modules.scala 46:47:@22652.4]
  assign _T_73330 = $signed(_T_73329); // @[Modules.scala 46:47:@22653.4]
  assign _T_73375 = $signed(io_in_146) - $signed(io_in_147); // @[Modules.scala 40:46:@22702.4]
  assign _T_73376 = _T_73375[4:0]; // @[Modules.scala 40:46:@22703.4]
  assign _T_73377 = $signed(_T_73376); // @[Modules.scala 40:46:@22704.4]
  assign _T_73382 = $signed(_T_61005) + $signed(io_in_149); // @[Modules.scala 43:47:@22709.4]
  assign _T_73383 = _T_73382[4:0]; // @[Modules.scala 43:47:@22710.4]
  assign _T_73384 = $signed(_T_73383); // @[Modules.scala 43:47:@22711.4]
  assign _T_73437 = $signed(_T_54722) - $signed(io_in_167); // @[Modules.scala 46:47:@22766.4]
  assign _T_73438 = _T_73437[4:0]; // @[Modules.scala 46:47:@22767.4]
  assign _T_73439 = $signed(_T_73438); // @[Modules.scala 46:47:@22768.4]
  assign _T_73454 = $signed(_T_61069) + $signed(io_in_173); // @[Modules.scala 43:47:@22784.4]
  assign _T_73455 = _T_73454[4:0]; // @[Modules.scala 43:47:@22785.4]
  assign _T_73456 = $signed(_T_73455); // @[Modules.scala 43:47:@22786.4]
  assign _T_73490 = $signed(_T_54791) + $signed(io_in_189); // @[Modules.scala 43:47:@22825.4]
  assign _T_73491 = _T_73490[4:0]; // @[Modules.scala 43:47:@22826.4]
  assign _T_73492 = $signed(_T_73491); // @[Modules.scala 43:47:@22827.4]
  assign _T_73507 = $signed(io_in_194) - $signed(io_in_195); // @[Modules.scala 40:46:@22843.4]
  assign _T_73508 = _T_73507[4:0]; // @[Modules.scala 40:46:@22844.4]
  assign _T_73509 = $signed(_T_73508); // @[Modules.scala 40:46:@22845.4]
  assign _T_73514 = $signed(_T_64354) - $signed(io_in_197); // @[Modules.scala 46:47:@22850.4]
  assign _T_73515 = _T_73514[4:0]; // @[Modules.scala 46:47:@22851.4]
  assign _T_73516 = $signed(_T_73515); // @[Modules.scala 46:47:@22852.4]
  assign _T_73530 = $signed(io_in_204) + $signed(io_in_205); // @[Modules.scala 37:46:@22869.4]
  assign _T_73531 = _T_73530[4:0]; // @[Modules.scala 37:46:@22870.4]
  assign _T_73532 = $signed(_T_73531); // @[Modules.scala 37:46:@22871.4]
  assign _T_73549 = $signed(io_in_214) - $signed(io_in_215); // @[Modules.scala 40:46:@22892.4]
  assign _T_73550 = _T_73549[4:0]; // @[Modules.scala 40:46:@22893.4]
  assign _T_73551 = $signed(_T_73550); // @[Modules.scala 40:46:@22894.4]
  assign _T_73608 = $signed(_T_54953) + $signed(io_in_241); // @[Modules.scala 43:47:@22959.4]
  assign _T_73609 = _T_73608[4:0]; // @[Modules.scala 43:47:@22960.4]
  assign _T_73610 = $signed(_T_73609); // @[Modules.scala 43:47:@22961.4]
  assign _T_73611 = $signed(io_in_242) - $signed(io_in_243); // @[Modules.scala 40:46:@22963.4]
  assign _T_73612 = _T_73611[4:0]; // @[Modules.scala 40:46:@22964.4]
  assign _T_73613 = $signed(_T_73612); // @[Modules.scala 40:46:@22965.4]
  assign _T_73617 = $signed(io_in_246) - $signed(io_in_247); // @[Modules.scala 40:46:@22971.4]
  assign _T_73618 = _T_73617[4:0]; // @[Modules.scala 40:46:@22972.4]
  assign _T_73619 = $signed(_T_73618); // @[Modules.scala 40:46:@22973.4]
  assign _T_73651 = $signed(io_in_258) - $signed(io_in_259); // @[Modules.scala 40:46:@23007.4]
  assign _T_73652 = _T_73651[4:0]; // @[Modules.scala 40:46:@23008.4]
  assign _T_73653 = $signed(_T_73652); // @[Modules.scala 40:46:@23009.4]
  assign _T_73657 = $signed(io_in_262) + $signed(io_in_263); // @[Modules.scala 37:46:@23015.4]
  assign _T_73658 = _T_73657[4:0]; // @[Modules.scala 37:46:@23016.4]
  assign _T_73659 = $signed(_T_73658); // @[Modules.scala 37:46:@23017.4]
  assign _T_73727 = $signed(io_in_290) - $signed(io_in_291); // @[Modules.scala 40:46:@23092.4]
  assign _T_73728 = _T_73727[4:0]; // @[Modules.scala 40:46:@23093.4]
  assign _T_73729 = $signed(_T_73728); // @[Modules.scala 40:46:@23094.4]
  assign _T_73750 = $signed(_T_55159) + $signed(io_in_301); // @[Modules.scala 43:47:@23118.4]
  assign _T_73751 = _T_73750[4:0]; // @[Modules.scala 43:47:@23119.4]
  assign _T_73752 = $signed(_T_73751); // @[Modules.scala 43:47:@23120.4]
  assign _T_73792 = $signed(_T_55201) + $signed(io_in_313); // @[Modules.scala 43:47:@23160.4]
  assign _T_73793 = _T_73792[4:0]; // @[Modules.scala 43:47:@23161.4]
  assign _T_73794 = $signed(_T_73793); // @[Modules.scala 43:47:@23162.4]
  assign _T_73806 = $signed(_T_58324) + $signed(io_in_317); // @[Modules.scala 43:47:@23174.4]
  assign _T_73807 = _T_73806[4:0]; // @[Modules.scala 43:47:@23175.4]
  assign _T_73808 = $signed(_T_73807); // @[Modules.scala 43:47:@23176.4]
  assign _T_73819 = $signed(_T_55228) + $signed(io_in_323); // @[Modules.scala 43:47:@23189.4]
  assign _T_73820 = _T_73819[4:0]; // @[Modules.scala 43:47:@23190.4]
  assign _T_73821 = $signed(_T_73820); // @[Modules.scala 43:47:@23191.4]
  assign _T_73822 = $signed(io_in_324) + $signed(io_in_325); // @[Modules.scala 37:46:@23193.4]
  assign _T_73823 = _T_73822[4:0]; // @[Modules.scala 37:46:@23194.4]
  assign _T_73824 = $signed(_T_73823); // @[Modules.scala 37:46:@23195.4]
  assign _T_73849 = $signed(_T_55266) - $signed(io_in_335); // @[Modules.scala 46:47:@23222.4]
  assign _T_73850 = _T_73849[4:0]; // @[Modules.scala 46:47:@23223.4]
  assign _T_73851 = $signed(_T_73850); // @[Modules.scala 46:47:@23224.4]
  assign _T_73859 = $signed(io_in_338) + $signed(io_in_339); // @[Modules.scala 37:46:@23233.4]
  assign _T_73860 = _T_73859[4:0]; // @[Modules.scala 37:46:@23234.4]
  assign _T_73861 = $signed(_T_73860); // @[Modules.scala 37:46:@23235.4]
  assign _T_73862 = $signed(io_in_340) + $signed(io_in_341); // @[Modules.scala 37:46:@23237.4]
  assign _T_73863 = _T_73862[4:0]; // @[Modules.scala 37:46:@23238.4]
  assign _T_73864 = $signed(_T_73863); // @[Modules.scala 37:46:@23239.4]
  assign _T_73869 = $signed(_T_64681) + $signed(io_in_343); // @[Modules.scala 43:47:@23244.4]
  assign _T_73870 = _T_73869[4:0]; // @[Modules.scala 43:47:@23245.4]
  assign _T_73871 = $signed(_T_73870); // @[Modules.scala 43:47:@23246.4]
  assign _T_73879 = $signed(_T_64695) + $signed(io_in_347); // @[Modules.scala 43:47:@23255.4]
  assign _T_73880 = _T_73879[4:0]; // @[Modules.scala 43:47:@23256.4]
  assign _T_73881 = $signed(_T_73880); // @[Modules.scala 43:47:@23257.4]
  assign _T_73893 = $signed(_T_58403) + $signed(io_in_351); // @[Modules.scala 43:47:@23269.4]
  assign _T_73894 = _T_73893[4:0]; // @[Modules.scala 43:47:@23270.4]
  assign _T_73895 = $signed(_T_73894); // @[Modules.scala 43:47:@23271.4]
  assign _T_73906 = $signed(_T_58424) + $signed(io_in_357); // @[Modules.scala 43:47:@23284.4]
  assign _T_73907 = _T_73906[4:0]; // @[Modules.scala 43:47:@23285.4]
  assign _T_73908 = $signed(_T_73907); // @[Modules.scala 43:47:@23286.4]
  assign _T_73909 = $signed(io_in_358) - $signed(io_in_359); // @[Modules.scala 40:46:@23288.4]
  assign _T_73910 = _T_73909[4:0]; // @[Modules.scala 40:46:@23289.4]
  assign _T_73911 = $signed(_T_73910); // @[Modules.scala 40:46:@23290.4]
  assign _T_73959 = $signed(_T_58481) + $signed(io_in_379); // @[Modules.scala 43:47:@23343.4]
  assign _T_73960 = _T_73959[4:0]; // @[Modules.scala 43:47:@23344.4]
  assign _T_73961 = $signed(_T_73960); // @[Modules.scala 43:47:@23345.4]
  assign _T_73992 = $signed(_T_55389) + $signed(io_in_393); // @[Modules.scala 43:47:@23380.4]
  assign _T_73993 = _T_73992[4:0]; // @[Modules.scala 43:47:@23381.4]
  assign _T_73994 = $signed(_T_73993); // @[Modules.scala 43:47:@23382.4]
  assign _T_74045 = $signed(io_in_414) - $signed(io_in_415); // @[Modules.scala 40:46:@23439.4]
  assign _T_74046 = _T_74045[4:0]; // @[Modules.scala 40:46:@23440.4]
  assign _T_74047 = $signed(_T_74046); // @[Modules.scala 40:46:@23441.4]
  assign _T_74079 = $signed(io_in_426) - $signed(io_in_427); // @[Modules.scala 40:46:@23475.4]
  assign _T_74080 = _T_74079[4:0]; // @[Modules.scala 40:46:@23476.4]
  assign _T_74081 = $signed(_T_74080); // @[Modules.scala 40:46:@23477.4]
  assign _T_74082 = $signed(io_in_428) - $signed(io_in_429); // @[Modules.scala 40:46:@23479.4]
  assign _T_74083 = _T_74082[4:0]; // @[Modules.scala 40:46:@23480.4]
  assign _T_74084 = $signed(_T_74083); // @[Modules.scala 40:46:@23481.4]
  assign _T_74089 = $signed(_T_61764) + $signed(io_in_431); // @[Modules.scala 43:47:@23486.4]
  assign _T_74090 = _T_74089[4:0]; // @[Modules.scala 43:47:@23487.4]
  assign _T_74091 = $signed(_T_74090); // @[Modules.scala 43:47:@23488.4]
  assign _T_74099 = $signed(_T_58621) + $signed(io_in_435); // @[Modules.scala 43:47:@23497.4]
  assign _T_74100 = _T_74099[4:0]; // @[Modules.scala 43:47:@23498.4]
  assign _T_74101 = $signed(_T_74100); // @[Modules.scala 43:47:@23499.4]
  assign _T_74105 = $signed(io_in_438) + $signed(io_in_439); // @[Modules.scala 37:46:@23505.4]
  assign _T_74106 = _T_74105[4:0]; // @[Modules.scala 37:46:@23506.4]
  assign _T_74107 = $signed(_T_74106); // @[Modules.scala 37:46:@23507.4]
  assign _T_74111 = $signed(io_in_442) - $signed(io_in_443); // @[Modules.scala 40:46:@23513.4]
  assign _T_74112 = _T_74111[4:0]; // @[Modules.scala 40:46:@23514.4]
  assign _T_74113 = $signed(_T_74112); // @[Modules.scala 40:46:@23515.4]
  assign _T_74151 = $signed(_T_61846) + $signed(io_in_459); // @[Modules.scala 43:47:@23557.4]
  assign _T_74152 = _T_74151[4:0]; // @[Modules.scala 43:47:@23558.4]
  assign _T_74153 = $signed(_T_74152); // @[Modules.scala 43:47:@23559.4]
  assign _T_74167 = $signed(io_in_466) - $signed(io_in_467); // @[Modules.scala 40:46:@23576.4]
  assign _T_74168 = _T_74167[4:0]; // @[Modules.scala 40:46:@23577.4]
  assign _T_74169 = $signed(_T_74168); // @[Modules.scala 40:46:@23578.4]
  assign _T_74173 = $signed(io_in_470) - $signed(io_in_471); // @[Modules.scala 40:46:@23584.4]
  assign _T_74174 = _T_74173[4:0]; // @[Modules.scala 40:46:@23585.4]
  assign _T_74175 = $signed(_T_74174); // @[Modules.scala 40:46:@23586.4]
  assign _T_74211 = $signed(_T_61906) + $signed(io_in_483); // @[Modules.scala 43:47:@23623.4]
  assign _T_74212 = _T_74211[4:0]; // @[Modules.scala 43:47:@23624.4]
  assign _T_74213 = $signed(_T_74212); // @[Modules.scala 43:47:@23625.4]
  assign _T_74260 = $signed(io_in_504) + $signed(io_in_505); // @[Modules.scala 37:46:@23679.4]
  assign _T_74261 = _T_74260[4:0]; // @[Modules.scala 37:46:@23680.4]
  assign _T_74262 = $signed(_T_74261); // @[Modules.scala 37:46:@23681.4]
  assign _T_74263 = $signed(io_in_506) - $signed(io_in_507); // @[Modules.scala 40:46:@23683.4]
  assign _T_74264 = _T_74263[4:0]; // @[Modules.scala 40:46:@23684.4]
  assign _T_74265 = $signed(_T_74264); // @[Modules.scala 40:46:@23685.4]
  assign _T_74315 = $signed(_T_55684) - $signed(io_in_523); // @[Modules.scala 46:47:@23736.4]
  assign _T_74316 = _T_74315[4:0]; // @[Modules.scala 46:47:@23737.4]
  assign _T_74317 = $signed(_T_74316); // @[Modules.scala 46:47:@23738.4]
  assign _T_74417 = $signed(5'sh0) - $signed(io_in_552); // @[Modules.scala 46:37:@23838.4]
  assign _T_74418 = _T_74417[4:0]; // @[Modules.scala 46:37:@23839.4]
  assign _T_74419 = $signed(_T_74418); // @[Modules.scala 46:37:@23840.4]
  assign _T_74420 = $signed(_T_74419) - $signed(io_in_553); // @[Modules.scala 46:47:@23841.4]
  assign _T_74421 = _T_74420[4:0]; // @[Modules.scala 46:47:@23842.4]
  assign _T_74422 = $signed(_T_74421); // @[Modules.scala 46:47:@23843.4]
  assign _T_74511 = $signed(_T_71337) - $signed(io_in_579); // @[Modules.scala 46:47:@23932.4]
  assign _T_74512 = _T_74511[4:0]; // @[Modules.scala 46:47:@23933.4]
  assign _T_74513 = $signed(_T_74512); // @[Modules.scala 46:47:@23934.4]
  assign _T_74542 = $signed(io_in_588) + $signed(io_in_589); // @[Modules.scala 37:46:@23964.4]
  assign _T_74543 = _T_74542[4:0]; // @[Modules.scala 37:46:@23965.4]
  assign _T_74544 = $signed(_T_74543); // @[Modules.scala 37:46:@23966.4]
  assign _T_74598 = $signed(_T_62261) - $signed(io_in_605); // @[Modules.scala 46:47:@24020.4]
  assign _T_74599 = _T_74598[4:0]; // @[Modules.scala 46:47:@24021.4]
  assign _T_74600 = $signed(_T_74599); // @[Modules.scala 46:47:@24022.4]
  assign _T_74626 = $signed(_T_59036) + $signed(io_in_613); // @[Modules.scala 43:47:@24048.4]
  assign _T_74627 = _T_74626[4:0]; // @[Modules.scala 43:47:@24049.4]
  assign _T_74628 = $signed(_T_74627); // @[Modules.scala 43:47:@24050.4]
  assign _T_74664 = $signed(_T_55977) + $signed(io_in_625); // @[Modules.scala 43:47:@24087.4]
  assign _T_74665 = _T_74664[4:0]; // @[Modules.scala 43:47:@24088.4]
  assign _T_74666 = $signed(_T_74665); // @[Modules.scala 43:47:@24089.4]
  assign _T_74681 = $signed(_T_55998) + $signed(io_in_631); // @[Modules.scala 43:47:@24105.4]
  assign _T_74682 = _T_74681[4:0]; // @[Modules.scala 43:47:@24106.4]
  assign _T_74683 = $signed(_T_74682); // @[Modules.scala 43:47:@24107.4]
  assign _T_74709 = $signed(_T_56026) - $signed(io_in_639); // @[Modules.scala 46:47:@24133.4]
  assign _T_74710 = _T_74709[4:0]; // @[Modules.scala 46:47:@24134.4]
  assign _T_74711 = $signed(_T_74710); // @[Modules.scala 46:47:@24135.4]
  assign _T_74730 = $signed(5'sh0) - $signed(io_in_646); // @[Modules.scala 46:37:@24155.4]
  assign _T_74731 = _T_74730[4:0]; // @[Modules.scala 46:37:@24156.4]
  assign _T_74732 = $signed(_T_74731); // @[Modules.scala 46:37:@24157.4]
  assign _T_74733 = $signed(_T_74732) - $signed(io_in_647); // @[Modules.scala 46:47:@24158.4]
  assign _T_74734 = _T_74733[4:0]; // @[Modules.scala 46:47:@24159.4]
  assign _T_74735 = $signed(_T_74734); // @[Modules.scala 46:47:@24160.4]
  assign _T_74749 = $signed(io_in_654) - $signed(io_in_655); // @[Modules.scala 40:46:@24177.4]
  assign _T_74750 = _T_74749[4:0]; // @[Modules.scala 40:46:@24178.4]
  assign _T_74751 = $signed(_T_74750); // @[Modules.scala 40:46:@24179.4]
  assign _T_74815 = $signed(_T_65483) - $signed(io_in_675); // @[Modules.scala 46:47:@24244.4]
  assign _T_74816 = _T_74815[4:0]; // @[Modules.scala 46:47:@24245.4]
  assign _T_74817 = $signed(_T_74816); // @[Modules.scala 46:47:@24246.4]
  assign _T_74927 = $signed(io_in_714) - $signed(io_in_715); // @[Modules.scala 40:46:@24363.4]
  assign _T_74928 = _T_74927[4:0]; // @[Modules.scala 40:46:@24364.4]
  assign _T_74929 = $signed(_T_74928); // @[Modules.scala 40:46:@24365.4]
  assign _T_74941 = $signed(_T_59275) + $signed(io_in_719); // @[Modules.scala 43:47:@24377.4]
  assign _T_74942 = _T_74941[4:0]; // @[Modules.scala 43:47:@24378.4]
  assign _T_74943 = $signed(_T_74942); // @[Modules.scala 43:47:@24379.4]
  assign _T_75056 = $signed(_T_59402) + $signed(io_in_769); // @[Modules.scala 43:47:@24507.4]
  assign _T_75057 = _T_75056[4:0]; // @[Modules.scala 43:47:@24508.4]
  assign _T_75058 = $signed(_T_75057); // @[Modules.scala 43:47:@24509.4]
  assign _T_75080 = $signed(_T_59430) + $signed(io_in_777); // @[Modules.scala 43:47:@24532.4]
  assign _T_75081 = _T_75080[4:0]; // @[Modules.scala 43:47:@24533.4]
  assign _T_75082 = $signed(_T_75081); // @[Modules.scala 43:47:@24534.4]
  assign _T_75103 = $signed(buffer_0_2) + $signed(buffer_2_3); // @[Modules.scala 50:57:@24558.4]
  assign _T_75104 = _T_75103[10:0]; // @[Modules.scala 50:57:@24559.4]
  assign buffer_6_393 = $signed(_T_75104); // @[Modules.scala 50:57:@24560.4]
  assign _T_75106 = $signed(buffer_2_4) + $signed(buffer_3_5); // @[Modules.scala 50:57:@24562.4]
  assign _T_75107 = _T_75106[10:0]; // @[Modules.scala 50:57:@24563.4]
  assign buffer_6_394 = $signed(_T_75107); // @[Modules.scala 50:57:@24564.4]
  assign _T_75139 = $signed(buffer_3_26) + $signed(buffer_0_27); // @[Modules.scala 50:57:@24606.4]
  assign _T_75140 = _T_75139[10:0]; // @[Modules.scala 50:57:@24607.4]
  assign buffer_6_405 = $signed(_T_75140); // @[Modules.scala 50:57:@24608.4]
  assign _T_75142 = $signed(buffer_2_28) + $signed(buffer_3_29); // @[Modules.scala 50:57:@24610.4]
  assign _T_75143 = _T_75142[10:0]; // @[Modules.scala 50:57:@24611.4]
  assign buffer_6_406 = $signed(_T_75143); // @[Modules.scala 50:57:@24612.4]
  assign _T_75163 = $signed(buffer_5_42) + $signed(buffer_3_43); // @[Modules.scala 50:57:@24638.4]
  assign _T_75164 = _T_75163[10:0]; // @[Modules.scala 50:57:@24639.4]
  assign buffer_6_413 = $signed(_T_75164); // @[Modules.scala 50:57:@24640.4]
  assign _T_75169 = $signed(buffer_3_46) + $signed(buffer_2_47); // @[Modules.scala 50:57:@24646.4]
  assign _T_75170 = _T_75169[10:0]; // @[Modules.scala 50:57:@24647.4]
  assign buffer_6_415 = $signed(_T_75170); // @[Modules.scala 50:57:@24648.4]
  assign buffer_6_50 = {{6{_T_73244[4]}},_T_73244}; // @[Modules.scala 32:22:@8.4]
  assign _T_75175 = $signed(buffer_6_50) + $signed(buffer_3_51); // @[Modules.scala 50:57:@24654.4]
  assign _T_75176 = _T_75175[10:0]; // @[Modules.scala 50:57:@24655.4]
  assign buffer_6_417 = $signed(_T_75176); // @[Modules.scala 50:57:@24656.4]
  assign buffer_6_53 = {{6{_T_73261[4]}},_T_73261}; // @[Modules.scala 32:22:@8.4]
  assign _T_75178 = $signed(buffer_3_52) + $signed(buffer_6_53); // @[Modules.scala 50:57:@24658.4]
  assign _T_75179 = _T_75178[10:0]; // @[Modules.scala 50:57:@24659.4]
  assign buffer_6_418 = $signed(_T_75179); // @[Modules.scala 50:57:@24660.4]
  assign _T_75181 = $signed(buffer_2_54) + $signed(buffer_0_55); // @[Modules.scala 50:57:@24662.4]
  assign _T_75182 = _T_75181[10:0]; // @[Modules.scala 50:57:@24663.4]
  assign buffer_6_419 = $signed(_T_75182); // @[Modules.scala 50:57:@24664.4]
  assign buffer_6_64 = {{6{_T_73330[4]}},_T_73330}; // @[Modules.scala 32:22:@8.4]
  assign _T_75196 = $signed(buffer_6_64) + $signed(buffer_2_65); // @[Modules.scala 50:57:@24682.4]
  assign _T_75197 = _T_75196[10:0]; // @[Modules.scala 50:57:@24683.4]
  assign buffer_6_424 = $signed(_T_75197); // @[Modules.scala 50:57:@24684.4]
  assign buffer_6_73 = {{6{_T_73377[4]}},_T_73377}; // @[Modules.scala 32:22:@8.4]
  assign _T_75208 = $signed(buffer_3_72) + $signed(buffer_6_73); // @[Modules.scala 50:57:@24698.4]
  assign _T_75209 = _T_75208[10:0]; // @[Modules.scala 50:57:@24699.4]
  assign buffer_6_428 = $signed(_T_75209); // @[Modules.scala 50:57:@24700.4]
  assign buffer_6_74 = {{6{_T_73384[4]}},_T_73384}; // @[Modules.scala 32:22:@8.4]
  assign _T_75211 = $signed(buffer_6_74) + $signed(buffer_0_75); // @[Modules.scala 50:57:@24702.4]
  assign _T_75212 = _T_75211[10:0]; // @[Modules.scala 50:57:@24703.4]
  assign buffer_6_429 = $signed(_T_75212); // @[Modules.scala 50:57:@24704.4]
  assign buffer_6_83 = {{6{_T_73439[4]}},_T_73439}; // @[Modules.scala 32:22:@8.4]
  assign _T_75223 = $signed(buffer_2_82) + $signed(buffer_6_83); // @[Modules.scala 50:57:@24718.4]
  assign _T_75224 = _T_75223[10:0]; // @[Modules.scala 50:57:@24719.4]
  assign buffer_6_433 = $signed(_T_75224); // @[Modules.scala 50:57:@24720.4]
  assign buffer_6_86 = {{6{_T_73456[4]}},_T_73456}; // @[Modules.scala 32:22:@8.4]
  assign _T_75229 = $signed(buffer_6_86) + $signed(buffer_1_87); // @[Modules.scala 50:57:@24726.4]
  assign _T_75230 = _T_75229[10:0]; // @[Modules.scala 50:57:@24727.4]
  assign buffer_6_435 = $signed(_T_75230); // @[Modules.scala 50:57:@24728.4]
  assign _T_75232 = $signed(buffer_0_88) + $signed(buffer_1_89); // @[Modules.scala 50:57:@24730.4]
  assign _T_75233 = _T_75232[10:0]; // @[Modules.scala 50:57:@24731.4]
  assign buffer_6_436 = $signed(_T_75233); // @[Modules.scala 50:57:@24732.4]
  assign buffer_6_94 = {{6{_T_73492[4]}},_T_73492}; // @[Modules.scala 32:22:@8.4]
  assign _T_75241 = $signed(buffer_6_94) + $signed(buffer_5_95); // @[Modules.scala 50:57:@24742.4]
  assign _T_75242 = _T_75241[10:0]; // @[Modules.scala 50:57:@24743.4]
  assign buffer_6_439 = $signed(_T_75242); // @[Modules.scala 50:57:@24744.4]
  assign buffer_6_97 = {{6{_T_73509[4]}},_T_73509}; // @[Modules.scala 32:22:@8.4]
  assign _T_75244 = $signed(buffer_1_96) + $signed(buffer_6_97); // @[Modules.scala 50:57:@24746.4]
  assign _T_75245 = _T_75244[10:0]; // @[Modules.scala 50:57:@24747.4]
  assign buffer_6_440 = $signed(_T_75245); // @[Modules.scala 50:57:@24748.4]
  assign buffer_6_98 = {{6{_T_73516[4]}},_T_73516}; // @[Modules.scala 32:22:@8.4]
  assign _T_75247 = $signed(buffer_6_98) + $signed(buffer_3_99); // @[Modules.scala 50:57:@24750.4]
  assign _T_75248 = _T_75247[10:0]; // @[Modules.scala 50:57:@24751.4]
  assign buffer_6_441 = $signed(_T_75248); // @[Modules.scala 50:57:@24752.4]
  assign _T_75250 = $signed(buffer_3_100) + $signed(buffer_4_101); // @[Modules.scala 50:57:@24754.4]
  assign _T_75251 = _T_75250[10:0]; // @[Modules.scala 50:57:@24755.4]
  assign buffer_6_442 = $signed(_T_75251); // @[Modules.scala 50:57:@24756.4]
  assign buffer_6_102 = {{6{_T_73532[4]}},_T_73532}; // @[Modules.scala 32:22:@8.4]
  assign _T_75253 = $signed(buffer_6_102) + $signed(buffer_3_103); // @[Modules.scala 50:57:@24758.4]
  assign _T_75254 = _T_75253[10:0]; // @[Modules.scala 50:57:@24759.4]
  assign buffer_6_443 = $signed(_T_75254); // @[Modules.scala 50:57:@24760.4]
  assign _T_75256 = $signed(buffer_3_104) + $signed(buffer_4_105); // @[Modules.scala 50:57:@24762.4]
  assign _T_75257 = _T_75256[10:0]; // @[Modules.scala 50:57:@24763.4]
  assign buffer_6_444 = $signed(_T_75257); // @[Modules.scala 50:57:@24764.4]
  assign buffer_6_107 = {{6{_T_73551[4]}},_T_73551}; // @[Modules.scala 32:22:@8.4]
  assign _T_75259 = $signed(buffer_3_106) + $signed(buffer_6_107); // @[Modules.scala 50:57:@24766.4]
  assign _T_75260 = _T_75259[10:0]; // @[Modules.scala 50:57:@24767.4]
  assign buffer_6_445 = $signed(_T_75260); // @[Modules.scala 50:57:@24768.4]
  assign _T_75262 = $signed(buffer_5_108) + $signed(buffer_3_109); // @[Modules.scala 50:57:@24770.4]
  assign _T_75263 = _T_75262[10:0]; // @[Modules.scala 50:57:@24771.4]
  assign buffer_6_446 = $signed(_T_75263); // @[Modules.scala 50:57:@24772.4]
  assign _T_75268 = $signed(buffer_0_112) + $signed(buffer_3_113); // @[Modules.scala 50:57:@24778.4]
  assign _T_75269 = _T_75268[10:0]; // @[Modules.scala 50:57:@24779.4]
  assign buffer_6_448 = $signed(_T_75269); // @[Modules.scala 50:57:@24780.4]
  assign _T_75274 = $signed(buffer_3_116) + $signed(buffer_2_117); // @[Modules.scala 50:57:@24786.4]
  assign _T_75275 = _T_75274[10:0]; // @[Modules.scala 50:57:@24787.4]
  assign buffer_6_450 = $signed(_T_75275); // @[Modules.scala 50:57:@24788.4]
  assign buffer_6_120 = {{6{_T_73610[4]}},_T_73610}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_121 = {{6{_T_73613[4]}},_T_73613}; // @[Modules.scala 32:22:@8.4]
  assign _T_75280 = $signed(buffer_6_120) + $signed(buffer_6_121); // @[Modules.scala 50:57:@24794.4]
  assign _T_75281 = _T_75280[10:0]; // @[Modules.scala 50:57:@24795.4]
  assign buffer_6_452 = $signed(_T_75281); // @[Modules.scala 50:57:@24796.4]
  assign buffer_6_123 = {{6{_T_73619[4]}},_T_73619}; // @[Modules.scala 32:22:@8.4]
  assign _T_75283 = $signed(buffer_3_122) + $signed(buffer_6_123); // @[Modules.scala 50:57:@24798.4]
  assign _T_75284 = _T_75283[10:0]; // @[Modules.scala 50:57:@24799.4]
  assign buffer_6_453 = $signed(_T_75284); // @[Modules.scala 50:57:@24800.4]
  assign _T_75289 = $signed(buffer_0_126) + $signed(buffer_3_127); // @[Modules.scala 50:57:@24806.4]
  assign _T_75290 = _T_75289[10:0]; // @[Modules.scala 50:57:@24807.4]
  assign buffer_6_455 = $signed(_T_75290); // @[Modules.scala 50:57:@24808.4]
  assign buffer_6_129 = {{6{_T_73653[4]}},_T_73653}; // @[Modules.scala 32:22:@8.4]
  assign _T_75292 = $signed(buffer_4_128) + $signed(buffer_6_129); // @[Modules.scala 50:57:@24810.4]
  assign _T_75293 = _T_75292[10:0]; // @[Modules.scala 50:57:@24811.4]
  assign buffer_6_456 = $signed(_T_75293); // @[Modules.scala 50:57:@24812.4]
  assign buffer_6_131 = {{6{_T_73659[4]}},_T_73659}; // @[Modules.scala 32:22:@8.4]
  assign _T_75295 = $signed(buffer_4_130) + $signed(buffer_6_131); // @[Modules.scala 50:57:@24814.4]
  assign _T_75296 = _T_75295[10:0]; // @[Modules.scala 50:57:@24815.4]
  assign buffer_6_457 = $signed(_T_75296); // @[Modules.scala 50:57:@24816.4]
  assign _T_75304 = $signed(buffer_5_136) + $signed(buffer_0_137); // @[Modules.scala 50:57:@24826.4]
  assign _T_75305 = _T_75304[10:0]; // @[Modules.scala 50:57:@24827.4]
  assign buffer_6_460 = $signed(_T_75305); // @[Modules.scala 50:57:@24828.4]
  assign _T_75310 = $signed(buffer_0_140) + $signed(buffer_3_141); // @[Modules.scala 50:57:@24834.4]
  assign _T_75311 = _T_75310[10:0]; // @[Modules.scala 50:57:@24835.4]
  assign buffer_6_462 = $signed(_T_75311); // @[Modules.scala 50:57:@24836.4]
  assign buffer_6_145 = {{6{_T_73729[4]}},_T_73729}; // @[Modules.scala 32:22:@8.4]
  assign _T_75316 = $signed(buffer_0_144) + $signed(buffer_6_145); // @[Modules.scala 50:57:@24842.4]
  assign _T_75317 = _T_75316[10:0]; // @[Modules.scala 50:57:@24843.4]
  assign buffer_6_464 = $signed(_T_75317); // @[Modules.scala 50:57:@24844.4]
  assign _T_75319 = $signed(buffer_1_146) + $signed(buffer_3_147); // @[Modules.scala 50:57:@24846.4]
  assign _T_75320 = _T_75319[10:0]; // @[Modules.scala 50:57:@24847.4]
  assign buffer_6_465 = $signed(_T_75320); // @[Modules.scala 50:57:@24848.4]
  assign _T_75322 = $signed(buffer_3_148) + $signed(buffer_4_149); // @[Modules.scala 50:57:@24850.4]
  assign _T_75323 = _T_75322[10:0]; // @[Modules.scala 50:57:@24851.4]
  assign buffer_6_466 = $signed(_T_75323); // @[Modules.scala 50:57:@24852.4]
  assign buffer_6_150 = {{6{_T_73752[4]}},_T_73752}; // @[Modules.scala 32:22:@8.4]
  assign _T_75325 = $signed(buffer_6_150) + $signed(buffer_0_151); // @[Modules.scala 50:57:@24854.4]
  assign _T_75326 = _T_75325[10:0]; // @[Modules.scala 50:57:@24855.4]
  assign buffer_6_467 = $signed(_T_75326); // @[Modules.scala 50:57:@24856.4]
  assign _T_75331 = $signed(buffer_3_154) + $signed(buffer_4_155); // @[Modules.scala 50:57:@24862.4]
  assign _T_75332 = _T_75331[10:0]; // @[Modules.scala 50:57:@24863.4]
  assign buffer_6_469 = $signed(_T_75332); // @[Modules.scala 50:57:@24864.4]
  assign buffer_6_156 = {{6{_T_73794[4]}},_T_73794}; // @[Modules.scala 32:22:@8.4]
  assign _T_75334 = $signed(buffer_6_156) + $signed(buffer_0_157); // @[Modules.scala 50:57:@24866.4]
  assign _T_75335 = _T_75334[10:0]; // @[Modules.scala 50:57:@24867.4]
  assign buffer_6_470 = $signed(_T_75335); // @[Modules.scala 50:57:@24868.4]
  assign buffer_6_158 = {{6{_T_73808[4]}},_T_73808}; // @[Modules.scala 32:22:@8.4]
  assign _T_75337 = $signed(buffer_6_158) + $signed(buffer_0_159); // @[Modules.scala 50:57:@24870.4]
  assign _T_75338 = _T_75337[10:0]; // @[Modules.scala 50:57:@24871.4]
  assign buffer_6_471 = $signed(_T_75338); // @[Modules.scala 50:57:@24872.4]
  assign buffer_6_161 = {{6{_T_73821[4]}},_T_73821}; // @[Modules.scala 32:22:@8.4]
  assign _T_75340 = $signed(buffer_2_160) + $signed(buffer_6_161); // @[Modules.scala 50:57:@24874.4]
  assign _T_75341 = _T_75340[10:0]; // @[Modules.scala 50:57:@24875.4]
  assign buffer_6_472 = $signed(_T_75341); // @[Modules.scala 50:57:@24876.4]
  assign buffer_6_162 = {{6{_T_73824[4]}},_T_73824}; // @[Modules.scala 32:22:@8.4]
  assign _T_75343 = $signed(buffer_6_162) + $signed(buffer_5_163); // @[Modules.scala 50:57:@24878.4]
  assign _T_75344 = _T_75343[10:0]; // @[Modules.scala 50:57:@24879.4]
  assign buffer_6_473 = $signed(_T_75344); // @[Modules.scala 50:57:@24880.4]
  assign buffer_6_167 = {{6{_T_73851[4]}},_T_73851}; // @[Modules.scala 32:22:@8.4]
  assign _T_75349 = $signed(buffer_0_166) + $signed(buffer_6_167); // @[Modules.scala 50:57:@24886.4]
  assign _T_75350 = _T_75349[10:0]; // @[Modules.scala 50:57:@24887.4]
  assign buffer_6_475 = $signed(_T_75350); // @[Modules.scala 50:57:@24888.4]
  assign buffer_6_169 = {{6{_T_73861[4]}},_T_73861}; // @[Modules.scala 32:22:@8.4]
  assign _T_75352 = $signed(buffer_3_168) + $signed(buffer_6_169); // @[Modules.scala 50:57:@24890.4]
  assign _T_75353 = _T_75352[10:0]; // @[Modules.scala 50:57:@24891.4]
  assign buffer_6_476 = $signed(_T_75353); // @[Modules.scala 50:57:@24892.4]
  assign buffer_6_170 = {{6{_T_73864[4]}},_T_73864}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_171 = {{6{_T_73871[4]}},_T_73871}; // @[Modules.scala 32:22:@8.4]
  assign _T_75355 = $signed(buffer_6_170) + $signed(buffer_6_171); // @[Modules.scala 50:57:@24894.4]
  assign _T_75356 = _T_75355[10:0]; // @[Modules.scala 50:57:@24895.4]
  assign buffer_6_477 = $signed(_T_75356); // @[Modules.scala 50:57:@24896.4]
  assign buffer_6_173 = {{6{_T_73881[4]}},_T_73881}; // @[Modules.scala 32:22:@8.4]
  assign _T_75358 = $signed(buffer_0_172) + $signed(buffer_6_173); // @[Modules.scala 50:57:@24898.4]
  assign _T_75359 = _T_75358[10:0]; // @[Modules.scala 50:57:@24899.4]
  assign buffer_6_478 = $signed(_T_75359); // @[Modules.scala 50:57:@24900.4]
  assign buffer_6_175 = {{6{_T_73895[4]}},_T_73895}; // @[Modules.scala 32:22:@8.4]
  assign _T_75361 = $signed(buffer_3_174) + $signed(buffer_6_175); // @[Modules.scala 50:57:@24902.4]
  assign _T_75362 = _T_75361[10:0]; // @[Modules.scala 50:57:@24903.4]
  assign buffer_6_479 = $signed(_T_75362); // @[Modules.scala 50:57:@24904.4]
  assign buffer_6_178 = {{6{_T_73908[4]}},_T_73908}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_179 = {{6{_T_73911[4]}},_T_73911}; // @[Modules.scala 32:22:@8.4]
  assign _T_75367 = $signed(buffer_6_178) + $signed(buffer_6_179); // @[Modules.scala 50:57:@24910.4]
  assign _T_75368 = _T_75367[10:0]; // @[Modules.scala 50:57:@24911.4]
  assign buffer_6_481 = $signed(_T_75368); // @[Modules.scala 50:57:@24912.4]
  assign _T_75373 = $signed(buffer_4_182) + $signed(buffer_5_183); // @[Modules.scala 50:57:@24918.4]
  assign _T_75374 = _T_75373[10:0]; // @[Modules.scala 50:57:@24919.4]
  assign buffer_6_483 = $signed(_T_75374); // @[Modules.scala 50:57:@24920.4]
  assign _T_75379 = $signed(buffer_5_186) + $signed(buffer_0_187); // @[Modules.scala 50:57:@24926.4]
  assign _T_75380 = _T_75379[10:0]; // @[Modules.scala 50:57:@24927.4]
  assign buffer_6_485 = $signed(_T_75380); // @[Modules.scala 50:57:@24928.4]
  assign buffer_6_189 = {{6{_T_73961[4]}},_T_73961}; // @[Modules.scala 32:22:@8.4]
  assign _T_75382 = $signed(buffer_3_188) + $signed(buffer_6_189); // @[Modules.scala 50:57:@24930.4]
  assign _T_75383 = _T_75382[10:0]; // @[Modules.scala 50:57:@24931.4]
  assign buffer_6_486 = $signed(_T_75383); // @[Modules.scala 50:57:@24932.4]
  assign buffer_6_196 = {{6{_T_73994[4]}},_T_73994}; // @[Modules.scala 32:22:@8.4]
  assign _T_75394 = $signed(buffer_6_196) + $signed(buffer_5_197); // @[Modules.scala 50:57:@24946.4]
  assign _T_75395 = _T_75394[10:0]; // @[Modules.scala 50:57:@24947.4]
  assign buffer_6_490 = $signed(_T_75395); // @[Modules.scala 50:57:@24948.4]
  assign _T_75400 = $signed(buffer_3_200) + $signed(buffer_5_201); // @[Modules.scala 50:57:@24954.4]
  assign _T_75401 = _T_75400[10:0]; // @[Modules.scala 50:57:@24955.4]
  assign buffer_6_492 = $signed(_T_75401); // @[Modules.scala 50:57:@24956.4]
  assign _T_75403 = $signed(buffer_3_202) + $signed(buffer_4_203); // @[Modules.scala 50:57:@24958.4]
  assign _T_75404 = _T_75403[10:0]; // @[Modules.scala 50:57:@24959.4]
  assign buffer_6_493 = $signed(_T_75404); // @[Modules.scala 50:57:@24960.4]
  assign buffer_6_207 = {{6{_T_74047[4]}},_T_74047}; // @[Modules.scala 32:22:@8.4]
  assign _T_75409 = $signed(buffer_4_206) + $signed(buffer_6_207); // @[Modules.scala 50:57:@24966.4]
  assign _T_75410 = _T_75409[10:0]; // @[Modules.scala 50:57:@24967.4]
  assign buffer_6_495 = $signed(_T_75410); // @[Modules.scala 50:57:@24968.4]
  assign _T_75412 = $signed(buffer_3_208) + $signed(buffer_0_209); // @[Modules.scala 50:57:@24970.4]
  assign _T_75413 = _T_75412[10:0]; // @[Modules.scala 50:57:@24971.4]
  assign buffer_6_496 = $signed(_T_75413); // @[Modules.scala 50:57:@24972.4]
  assign _T_75415 = $signed(buffer_0_210) + $signed(buffer_5_211); // @[Modules.scala 50:57:@24974.4]
  assign _T_75416 = _T_75415[10:0]; // @[Modules.scala 50:57:@24975.4]
  assign buffer_6_497 = $signed(_T_75416); // @[Modules.scala 50:57:@24976.4]
  assign buffer_6_213 = {{6{_T_74081[4]}},_T_74081}; // @[Modules.scala 32:22:@8.4]
  assign _T_75418 = $signed(buffer_3_212) + $signed(buffer_6_213); // @[Modules.scala 50:57:@24978.4]
  assign _T_75419 = _T_75418[10:0]; // @[Modules.scala 50:57:@24979.4]
  assign buffer_6_498 = $signed(_T_75419); // @[Modules.scala 50:57:@24980.4]
  assign buffer_6_214 = {{6{_T_74084[4]}},_T_74084}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_215 = {{6{_T_74091[4]}},_T_74091}; // @[Modules.scala 32:22:@8.4]
  assign _T_75421 = $signed(buffer_6_214) + $signed(buffer_6_215); // @[Modules.scala 50:57:@24982.4]
  assign _T_75422 = _T_75421[10:0]; // @[Modules.scala 50:57:@24983.4]
  assign buffer_6_499 = $signed(_T_75422); // @[Modules.scala 50:57:@24984.4]
  assign buffer_6_217 = {{6{_T_74101[4]}},_T_74101}; // @[Modules.scala 32:22:@8.4]
  assign _T_75424 = $signed(buffer_4_216) + $signed(buffer_6_217); // @[Modules.scala 50:57:@24986.4]
  assign _T_75425 = _T_75424[10:0]; // @[Modules.scala 50:57:@24987.4]
  assign buffer_6_500 = $signed(_T_75425); // @[Modules.scala 50:57:@24988.4]
  assign buffer_6_219 = {{6{_T_74107[4]}},_T_74107}; // @[Modules.scala 32:22:@8.4]
  assign _T_75427 = $signed(buffer_0_218) + $signed(buffer_6_219); // @[Modules.scala 50:57:@24990.4]
  assign _T_75428 = _T_75427[10:0]; // @[Modules.scala 50:57:@24991.4]
  assign buffer_6_501 = $signed(_T_75428); // @[Modules.scala 50:57:@24992.4]
  assign buffer_6_221 = {{6{_T_74113[4]}},_T_74113}; // @[Modules.scala 32:22:@8.4]
  assign _T_75430 = $signed(buffer_0_220) + $signed(buffer_6_221); // @[Modules.scala 50:57:@24994.4]
  assign _T_75431 = _T_75430[10:0]; // @[Modules.scala 50:57:@24995.4]
  assign buffer_6_502 = $signed(_T_75431); // @[Modules.scala 50:57:@24996.4]
  assign _T_75436 = $signed(buffer_3_224) + $signed(buffer_0_225); // @[Modules.scala 50:57:@25002.4]
  assign _T_75437 = _T_75436[10:0]; // @[Modules.scala 50:57:@25003.4]
  assign buffer_6_504 = $signed(_T_75437); // @[Modules.scala 50:57:@25004.4]
  assign buffer_6_229 = {{6{_T_74153[4]}},_T_74153}; // @[Modules.scala 32:22:@8.4]
  assign _T_75442 = $signed(buffer_2_228) + $signed(buffer_6_229); // @[Modules.scala 50:57:@25010.4]
  assign _T_75443 = _T_75442[10:0]; // @[Modules.scala 50:57:@25011.4]
  assign buffer_6_506 = $signed(_T_75443); // @[Modules.scala 50:57:@25012.4]
  assign _T_75445 = $signed(buffer_1_230) + $signed(buffer_0_231); // @[Modules.scala 50:57:@25014.4]
  assign _T_75446 = _T_75445[10:0]; // @[Modules.scala 50:57:@25015.4]
  assign buffer_6_507 = $signed(_T_75446); // @[Modules.scala 50:57:@25016.4]
  assign buffer_6_233 = {{6{_T_74169[4]}},_T_74169}; // @[Modules.scala 32:22:@8.4]
  assign _T_75448 = $signed(buffer_0_232) + $signed(buffer_6_233); // @[Modules.scala 50:57:@25018.4]
  assign _T_75449 = _T_75448[10:0]; // @[Modules.scala 50:57:@25019.4]
  assign buffer_6_508 = $signed(_T_75449); // @[Modules.scala 50:57:@25020.4]
  assign buffer_6_235 = {{6{_T_74175[4]}},_T_74175}; // @[Modules.scala 32:22:@8.4]
  assign _T_75451 = $signed(buffer_0_234) + $signed(buffer_6_235); // @[Modules.scala 50:57:@25022.4]
  assign _T_75452 = _T_75451[10:0]; // @[Modules.scala 50:57:@25023.4]
  assign buffer_6_509 = $signed(_T_75452); // @[Modules.scala 50:57:@25024.4]
  assign _T_75457 = $signed(buffer_1_238) + $signed(buffer_0_239); // @[Modules.scala 50:57:@25030.4]
  assign _T_75458 = _T_75457[10:0]; // @[Modules.scala 50:57:@25031.4]
  assign buffer_6_511 = $signed(_T_75458); // @[Modules.scala 50:57:@25032.4]
  assign buffer_6_241 = {{6{_T_74213[4]}},_T_74213}; // @[Modules.scala 32:22:@8.4]
  assign _T_75460 = $signed(buffer_0_240) + $signed(buffer_6_241); // @[Modules.scala 50:57:@25034.4]
  assign _T_75461 = _T_75460[10:0]; // @[Modules.scala 50:57:@25035.4]
  assign buffer_6_512 = $signed(_T_75461); // @[Modules.scala 50:57:@25036.4]
  assign _T_75463 = $signed(buffer_5_242) + $signed(buffer_0_243); // @[Modules.scala 50:57:@25038.4]
  assign _T_75464 = _T_75463[10:0]; // @[Modules.scala 50:57:@25039.4]
  assign buffer_6_513 = $signed(_T_75464); // @[Modules.scala 50:57:@25040.4]
  assign _T_75469 = $signed(buffer_4_246) + $signed(buffer_0_247); // @[Modules.scala 50:57:@25046.4]
  assign _T_75470 = _T_75469[10:0]; // @[Modules.scala 50:57:@25047.4]
  assign buffer_6_515 = $signed(_T_75470); // @[Modules.scala 50:57:@25048.4]
  assign buffer_6_252 = {{6{_T_74262[4]}},_T_74262}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_253 = {{6{_T_74265[4]}},_T_74265}; // @[Modules.scala 32:22:@8.4]
  assign _T_75478 = $signed(buffer_6_252) + $signed(buffer_6_253); // @[Modules.scala 50:57:@25058.4]
  assign _T_75479 = _T_75478[10:0]; // @[Modules.scala 50:57:@25059.4]
  assign buffer_6_518 = $signed(_T_75479); // @[Modules.scala 50:57:@25060.4]
  assign _T_75487 = $signed(buffer_1_258) + $signed(buffer_0_259); // @[Modules.scala 50:57:@25070.4]
  assign _T_75488 = _T_75487[10:0]; // @[Modules.scala 50:57:@25071.4]
  assign buffer_6_521 = $signed(_T_75488); // @[Modules.scala 50:57:@25072.4]
  assign buffer_6_261 = {{6{_T_74317[4]}},_T_74317}; // @[Modules.scala 32:22:@8.4]
  assign _T_75490 = $signed(buffer_2_260) + $signed(buffer_6_261); // @[Modules.scala 50:57:@25074.4]
  assign _T_75491 = _T_75490[10:0]; // @[Modules.scala 50:57:@25075.4]
  assign buffer_6_522 = $signed(_T_75491); // @[Modules.scala 50:57:@25076.4]
  assign _T_75505 = $signed(buffer_0_270) + $signed(buffer_3_271); // @[Modules.scala 50:57:@25094.4]
  assign _T_75506 = _T_75505[10:0]; // @[Modules.scala 50:57:@25095.4]
  assign buffer_6_527 = $signed(_T_75506); // @[Modules.scala 50:57:@25096.4]
  assign buffer_6_276 = {{6{_T_74422[4]}},_T_74422}; // @[Modules.scala 32:22:@8.4]
  assign _T_75514 = $signed(buffer_6_276) + $signed(buffer_0_277); // @[Modules.scala 50:57:@25106.4]
  assign _T_75515 = _T_75514[10:0]; // @[Modules.scala 50:57:@25107.4]
  assign buffer_6_530 = $signed(_T_75515); // @[Modules.scala 50:57:@25108.4]
  assign buffer_6_289 = {{6{_T_74513[4]}},_T_74513}; // @[Modules.scala 32:22:@8.4]
  assign _T_75532 = $signed(buffer_5_288) + $signed(buffer_6_289); // @[Modules.scala 50:57:@25130.4]
  assign _T_75533 = _T_75532[10:0]; // @[Modules.scala 50:57:@25131.4]
  assign buffer_6_536 = $signed(_T_75533); // @[Modules.scala 50:57:@25132.4]
  assign _T_75538 = $signed(buffer_1_292) + $signed(buffer_4_293); // @[Modules.scala 50:57:@25138.4]
  assign _T_75539 = _T_75538[10:0]; // @[Modules.scala 50:57:@25139.4]
  assign buffer_6_538 = $signed(_T_75539); // @[Modules.scala 50:57:@25140.4]
  assign buffer_6_294 = {{6{_T_74544[4]}},_T_74544}; // @[Modules.scala 32:22:@8.4]
  assign _T_75541 = $signed(buffer_6_294) + $signed(buffer_0_295); // @[Modules.scala 50:57:@25142.4]
  assign _T_75542 = _T_75541[10:0]; // @[Modules.scala 50:57:@25143.4]
  assign buffer_6_539 = $signed(_T_75542); // @[Modules.scala 50:57:@25144.4]
  assign buffer_6_302 = {{6{_T_74600[4]}},_T_74600}; // @[Modules.scala 32:22:@8.4]
  assign _T_75553 = $signed(buffer_6_302) + $signed(buffer_2_303); // @[Modules.scala 50:57:@25158.4]
  assign _T_75554 = _T_75553[10:0]; // @[Modules.scala 50:57:@25159.4]
  assign buffer_6_543 = $signed(_T_75554); // @[Modules.scala 50:57:@25160.4]
  assign buffer_6_306 = {{6{_T_74628[4]}},_T_74628}; // @[Modules.scala 32:22:@8.4]
  assign _T_75559 = $signed(buffer_6_306) + $signed(buffer_0_307); // @[Modules.scala 50:57:@25166.4]
  assign _T_75560 = _T_75559[10:0]; // @[Modules.scala 50:57:@25167.4]
  assign buffer_6_545 = $signed(_T_75560); // @[Modules.scala 50:57:@25168.4]
  assign buffer_6_312 = {{6{_T_74666[4]}},_T_74666}; // @[Modules.scala 32:22:@8.4]
  assign _T_75568 = $signed(buffer_6_312) + $signed(buffer_0_313); // @[Modules.scala 50:57:@25178.4]
  assign _T_75569 = _T_75568[10:0]; // @[Modules.scala 50:57:@25179.4]
  assign buffer_6_548 = $signed(_T_75569); // @[Modules.scala 50:57:@25180.4]
  assign buffer_6_315 = {{6{_T_74683[4]}},_T_74683}; // @[Modules.scala 32:22:@8.4]
  assign _T_75571 = $signed(buffer_5_314) + $signed(buffer_6_315); // @[Modules.scala 50:57:@25182.4]
  assign _T_75572 = _T_75571[10:0]; // @[Modules.scala 50:57:@25183.4]
  assign buffer_6_549 = $signed(_T_75572); // @[Modules.scala 50:57:@25184.4]
  assign buffer_6_319 = {{6{_T_74711[4]}},_T_74711}; // @[Modules.scala 32:22:@8.4]
  assign _T_75577 = $signed(buffer_0_318) + $signed(buffer_6_319); // @[Modules.scala 50:57:@25190.4]
  assign _T_75578 = _T_75577[10:0]; // @[Modules.scala 50:57:@25191.4]
  assign buffer_6_551 = $signed(_T_75578); // @[Modules.scala 50:57:@25192.4]
  assign buffer_6_323 = {{6{_T_74735[4]}},_T_74735}; // @[Modules.scala 32:22:@8.4]
  assign _T_75583 = $signed(buffer_1_322) + $signed(buffer_6_323); // @[Modules.scala 50:57:@25198.4]
  assign _T_75584 = _T_75583[10:0]; // @[Modules.scala 50:57:@25199.4]
  assign buffer_6_553 = $signed(_T_75584); // @[Modules.scala 50:57:@25200.4]
  assign _T_75586 = $signed(buffer_0_324) + $signed(buffer_1_325); // @[Modules.scala 50:57:@25202.4]
  assign _T_75587 = _T_75586[10:0]; // @[Modules.scala 50:57:@25203.4]
  assign buffer_6_554 = $signed(_T_75587); // @[Modules.scala 50:57:@25204.4]
  assign buffer_6_327 = {{6{_T_74751[4]}},_T_74751}; // @[Modules.scala 32:22:@8.4]
  assign _T_75589 = $signed(buffer_5_326) + $signed(buffer_6_327); // @[Modules.scala 50:57:@25206.4]
  assign _T_75590 = _T_75589[10:0]; // @[Modules.scala 50:57:@25207.4]
  assign buffer_6_555 = $signed(_T_75590); // @[Modules.scala 50:57:@25208.4]
  assign _T_75601 = $signed(buffer_1_334) + $signed(buffer_4_335); // @[Modules.scala 50:57:@25222.4]
  assign _T_75602 = _T_75601[10:0]; // @[Modules.scala 50:57:@25223.4]
  assign buffer_6_559 = $signed(_T_75602); // @[Modules.scala 50:57:@25224.4]
  assign buffer_6_337 = {{6{_T_74817[4]}},_T_74817}; // @[Modules.scala 32:22:@8.4]
  assign _T_75604 = $signed(buffer_4_336) + $signed(buffer_6_337); // @[Modules.scala 50:57:@25226.4]
  assign _T_75605 = _T_75604[10:0]; // @[Modules.scala 50:57:@25227.4]
  assign buffer_6_560 = $signed(_T_75605); // @[Modules.scala 50:57:@25228.4]
  assign _T_75616 = $signed(buffer_2_344) + $signed(buffer_3_345); // @[Modules.scala 50:57:@25242.4]
  assign _T_75617 = _T_75616[10:0]; // @[Modules.scala 50:57:@25243.4]
  assign buffer_6_564 = $signed(_T_75617); // @[Modules.scala 50:57:@25244.4]
  assign _T_75619 = $signed(buffer_0_346) + $signed(buffer_1_347); // @[Modules.scala 50:57:@25246.4]
  assign _T_75620 = _T_75619[10:0]; // @[Modules.scala 50:57:@25247.4]
  assign buffer_6_565 = $signed(_T_75620); // @[Modules.scala 50:57:@25248.4]
  assign _T_75631 = $signed(buffer_0_354) + $signed(buffer_1_355); // @[Modules.scala 50:57:@25262.4]
  assign _T_75632 = _T_75631[10:0]; // @[Modules.scala 50:57:@25263.4]
  assign buffer_6_569 = $signed(_T_75632); // @[Modules.scala 50:57:@25264.4]
  assign buffer_6_357 = {{6{_T_74929[4]}},_T_74929}; // @[Modules.scala 32:22:@8.4]
  assign _T_75634 = $signed(buffer_1_356) + $signed(buffer_6_357); // @[Modules.scala 50:57:@25266.4]
  assign _T_75635 = _T_75634[10:0]; // @[Modules.scala 50:57:@25267.4]
  assign buffer_6_570 = $signed(_T_75635); // @[Modules.scala 50:57:@25268.4]
  assign buffer_6_359 = {{6{_T_74943[4]}},_T_74943}; // @[Modules.scala 32:22:@8.4]
  assign _T_75637 = $signed(buffer_2_358) + $signed(buffer_6_359); // @[Modules.scala 50:57:@25270.4]
  assign _T_75638 = _T_75637[10:0]; // @[Modules.scala 50:57:@25271.4]
  assign buffer_6_571 = $signed(_T_75638); // @[Modules.scala 50:57:@25272.4]
  assign _T_75643 = $signed(buffer_4_362) + $signed(buffer_0_363); // @[Modules.scala 50:57:@25278.4]
  assign _T_75644 = _T_75643[10:0]; // @[Modules.scala 50:57:@25279.4]
  assign buffer_6_573 = $signed(_T_75644); // @[Modules.scala 50:57:@25280.4]
  assign _T_75646 = $signed(buffer_0_364) + $signed(buffer_2_365); // @[Modules.scala 50:57:@25282.4]
  assign _T_75647 = _T_75646[10:0]; // @[Modules.scala 50:57:@25283.4]
  assign buffer_6_574 = $signed(_T_75647); // @[Modules.scala 50:57:@25284.4]
  assign _T_75661 = $signed(buffer_0_374) + $signed(buffer_4_375); // @[Modules.scala 50:57:@25302.4]
  assign _T_75662 = _T_75661[10:0]; // @[Modules.scala 50:57:@25303.4]
  assign buffer_6_579 = $signed(_T_75662); // @[Modules.scala 50:57:@25304.4]
  assign buffer_6_384 = {{6{_T_75058[4]}},_T_75058}; // @[Modules.scala 32:22:@8.4]
  assign _T_75676 = $signed(buffer_6_384) + $signed(buffer_3_385); // @[Modules.scala 50:57:@25322.4]
  assign _T_75677 = _T_75676[10:0]; // @[Modules.scala 50:57:@25323.4]
  assign buffer_6_584 = $signed(_T_75677); // @[Modules.scala 50:57:@25324.4]
  assign buffer_6_388 = {{6{_T_75082[4]}},_T_75082}; // @[Modules.scala 32:22:@8.4]
  assign _T_75682 = $signed(buffer_6_388) + $signed(buffer_5_389); // @[Modules.scala 50:57:@25330.4]
  assign _T_75683 = _T_75682[10:0]; // @[Modules.scala 50:57:@25331.4]
  assign buffer_6_586 = $signed(_T_75683); // @[Modules.scala 50:57:@25332.4]
  assign _T_75688 = $signed(buffer_0_392) + $signed(buffer_6_393); // @[Modules.scala 53:83:@25338.4]
  assign _T_75689 = _T_75688[10:0]; // @[Modules.scala 53:83:@25339.4]
  assign buffer_6_588 = $signed(_T_75689); // @[Modules.scala 53:83:@25340.4]
  assign _T_75691 = $signed(buffer_6_394) + $signed(buffer_0_395); // @[Modules.scala 53:83:@25342.4]
  assign _T_75692 = _T_75691[10:0]; // @[Modules.scala 53:83:@25343.4]
  assign buffer_6_589 = $signed(_T_75692); // @[Modules.scala 53:83:@25344.4]
  assign _T_75694 = $signed(buffer_1_396) + $signed(buffer_4_397); // @[Modules.scala 53:83:@25346.4]
  assign _T_75695 = _T_75694[10:0]; // @[Modules.scala 53:83:@25347.4]
  assign buffer_6_590 = $signed(_T_75695); // @[Modules.scala 53:83:@25348.4]
  assign _T_75697 = $signed(buffer_1_398) + $signed(buffer_0_399); // @[Modules.scala 53:83:@25350.4]
  assign _T_75698 = _T_75697[10:0]; // @[Modules.scala 53:83:@25351.4]
  assign buffer_6_591 = $signed(_T_75698); // @[Modules.scala 53:83:@25352.4]
  assign _T_75700 = $signed(buffer_3_400) + $signed(buffer_0_401); // @[Modules.scala 53:83:@25354.4]
  assign _T_75701 = _T_75700[10:0]; // @[Modules.scala 53:83:@25355.4]
  assign buffer_6_592 = $signed(_T_75701); // @[Modules.scala 53:83:@25356.4]
  assign _T_75706 = $signed(buffer_0_404) + $signed(buffer_6_405); // @[Modules.scala 53:83:@25362.4]
  assign _T_75707 = _T_75706[10:0]; // @[Modules.scala 53:83:@25363.4]
  assign buffer_6_594 = $signed(_T_75707); // @[Modules.scala 53:83:@25364.4]
  assign _T_75709 = $signed(buffer_6_406) + $signed(buffer_0_407); // @[Modules.scala 53:83:@25366.4]
  assign _T_75710 = _T_75709[10:0]; // @[Modules.scala 53:83:@25367.4]
  assign buffer_6_595 = $signed(_T_75710); // @[Modules.scala 53:83:@25368.4]
  assign _T_75718 = $signed(buffer_2_412) + $signed(buffer_6_413); // @[Modules.scala 53:83:@25378.4]
  assign _T_75719 = _T_75718[10:0]; // @[Modules.scala 53:83:@25379.4]
  assign buffer_6_598 = $signed(_T_75719); // @[Modules.scala 53:83:@25380.4]
  assign _T_75721 = $signed(buffer_3_414) + $signed(buffer_6_415); // @[Modules.scala 53:83:@25382.4]
  assign _T_75722 = _T_75721[10:0]; // @[Modules.scala 53:83:@25383.4]
  assign buffer_6_599 = $signed(_T_75722); // @[Modules.scala 53:83:@25384.4]
  assign _T_75724 = $signed(buffer_2_416) + $signed(buffer_6_417); // @[Modules.scala 53:83:@25386.4]
  assign _T_75725 = _T_75724[10:0]; // @[Modules.scala 53:83:@25387.4]
  assign buffer_6_600 = $signed(_T_75725); // @[Modules.scala 53:83:@25388.4]
  assign _T_75727 = $signed(buffer_6_418) + $signed(buffer_6_419); // @[Modules.scala 53:83:@25390.4]
  assign _T_75728 = _T_75727[10:0]; // @[Modules.scala 53:83:@25391.4]
  assign buffer_6_601 = $signed(_T_75728); // @[Modules.scala 53:83:@25392.4]
  assign _T_75730 = $signed(buffer_5_420) + $signed(buffer_2_421); // @[Modules.scala 53:83:@25394.4]
  assign _T_75731 = _T_75730[10:0]; // @[Modules.scala 53:83:@25395.4]
  assign buffer_6_602 = $signed(_T_75731); // @[Modules.scala 53:83:@25396.4]
  assign _T_75736 = $signed(buffer_6_424) + $signed(buffer_0_425); // @[Modules.scala 53:83:@25402.4]
  assign _T_75737 = _T_75736[10:0]; // @[Modules.scala 53:83:@25403.4]
  assign buffer_6_604 = $signed(_T_75737); // @[Modules.scala 53:83:@25404.4]
  assign _T_75739 = $signed(buffer_0_426) + $signed(buffer_4_427); // @[Modules.scala 53:83:@25406.4]
  assign _T_75740 = _T_75739[10:0]; // @[Modules.scala 53:83:@25407.4]
  assign buffer_6_605 = $signed(_T_75740); // @[Modules.scala 53:83:@25408.4]
  assign _T_75742 = $signed(buffer_6_428) + $signed(buffer_6_429); // @[Modules.scala 53:83:@25410.4]
  assign _T_75743 = _T_75742[10:0]; // @[Modules.scala 53:83:@25411.4]
  assign buffer_6_606 = $signed(_T_75743); // @[Modules.scala 53:83:@25412.4]
  assign _T_75748 = $signed(buffer_0_432) + $signed(buffer_6_433); // @[Modules.scala 53:83:@25418.4]
  assign _T_75749 = _T_75748[10:0]; // @[Modules.scala 53:83:@25419.4]
  assign buffer_6_608 = $signed(_T_75749); // @[Modules.scala 53:83:@25420.4]
  assign _T_75751 = $signed(buffer_2_434) + $signed(buffer_6_435); // @[Modules.scala 53:83:@25422.4]
  assign _T_75752 = _T_75751[10:0]; // @[Modules.scala 53:83:@25423.4]
  assign buffer_6_609 = $signed(_T_75752); // @[Modules.scala 53:83:@25424.4]
  assign _T_75754 = $signed(buffer_6_436) + $signed(buffer_1_437); // @[Modules.scala 53:83:@25426.4]
  assign _T_75755 = _T_75754[10:0]; // @[Modules.scala 53:83:@25427.4]
  assign buffer_6_610 = $signed(_T_75755); // @[Modules.scala 53:83:@25428.4]
  assign _T_75757 = $signed(buffer_3_438) + $signed(buffer_6_439); // @[Modules.scala 53:83:@25430.4]
  assign _T_75758 = _T_75757[10:0]; // @[Modules.scala 53:83:@25431.4]
  assign buffer_6_611 = $signed(_T_75758); // @[Modules.scala 53:83:@25432.4]
  assign _T_75760 = $signed(buffer_6_440) + $signed(buffer_6_441); // @[Modules.scala 53:83:@25434.4]
  assign _T_75761 = _T_75760[10:0]; // @[Modules.scala 53:83:@25435.4]
  assign buffer_6_612 = $signed(_T_75761); // @[Modules.scala 53:83:@25436.4]
  assign _T_75763 = $signed(buffer_6_442) + $signed(buffer_6_443); // @[Modules.scala 53:83:@25438.4]
  assign _T_75764 = _T_75763[10:0]; // @[Modules.scala 53:83:@25439.4]
  assign buffer_6_613 = $signed(_T_75764); // @[Modules.scala 53:83:@25440.4]
  assign _T_75766 = $signed(buffer_6_444) + $signed(buffer_6_445); // @[Modules.scala 53:83:@25442.4]
  assign _T_75767 = _T_75766[10:0]; // @[Modules.scala 53:83:@25443.4]
  assign buffer_6_614 = $signed(_T_75767); // @[Modules.scala 53:83:@25444.4]
  assign _T_75769 = $signed(buffer_6_446) + $signed(buffer_5_447); // @[Modules.scala 53:83:@25446.4]
  assign _T_75770 = _T_75769[10:0]; // @[Modules.scala 53:83:@25447.4]
  assign buffer_6_615 = $signed(_T_75770); // @[Modules.scala 53:83:@25448.4]
  assign _T_75772 = $signed(buffer_6_448) + $signed(buffer_3_449); // @[Modules.scala 53:83:@25450.4]
  assign _T_75773 = _T_75772[10:0]; // @[Modules.scala 53:83:@25451.4]
  assign buffer_6_616 = $signed(_T_75773); // @[Modules.scala 53:83:@25452.4]
  assign _T_75775 = $signed(buffer_6_450) + $signed(buffer_3_451); // @[Modules.scala 53:83:@25454.4]
  assign _T_75776 = _T_75775[10:0]; // @[Modules.scala 53:83:@25455.4]
  assign buffer_6_617 = $signed(_T_75776); // @[Modules.scala 53:83:@25456.4]
  assign _T_75778 = $signed(buffer_6_452) + $signed(buffer_6_453); // @[Modules.scala 53:83:@25458.4]
  assign _T_75779 = _T_75778[10:0]; // @[Modules.scala 53:83:@25459.4]
  assign buffer_6_618 = $signed(_T_75779); // @[Modules.scala 53:83:@25460.4]
  assign _T_75781 = $signed(buffer_0_454) + $signed(buffer_6_455); // @[Modules.scala 53:83:@25462.4]
  assign _T_75782 = _T_75781[10:0]; // @[Modules.scala 53:83:@25463.4]
  assign buffer_6_619 = $signed(_T_75782); // @[Modules.scala 53:83:@25464.4]
  assign _T_75784 = $signed(buffer_6_456) + $signed(buffer_6_457); // @[Modules.scala 53:83:@25466.4]
  assign _T_75785 = _T_75784[10:0]; // @[Modules.scala 53:83:@25467.4]
  assign buffer_6_620 = $signed(_T_75785); // @[Modules.scala 53:83:@25468.4]
  assign _T_75790 = $signed(buffer_6_460) + $signed(buffer_0_461); // @[Modules.scala 53:83:@25474.4]
  assign _T_75791 = _T_75790[10:0]; // @[Modules.scala 53:83:@25475.4]
  assign buffer_6_622 = $signed(_T_75791); // @[Modules.scala 53:83:@25476.4]
  assign _T_75793 = $signed(buffer_6_462) + $signed(buffer_0_463); // @[Modules.scala 53:83:@25478.4]
  assign _T_75794 = _T_75793[10:0]; // @[Modules.scala 53:83:@25479.4]
  assign buffer_6_623 = $signed(_T_75794); // @[Modules.scala 53:83:@25480.4]
  assign _T_75796 = $signed(buffer_6_464) + $signed(buffer_6_465); // @[Modules.scala 53:83:@25482.4]
  assign _T_75797 = _T_75796[10:0]; // @[Modules.scala 53:83:@25483.4]
  assign buffer_6_624 = $signed(_T_75797); // @[Modules.scala 53:83:@25484.4]
  assign _T_75799 = $signed(buffer_6_466) + $signed(buffer_6_467); // @[Modules.scala 53:83:@25486.4]
  assign _T_75800 = _T_75799[10:0]; // @[Modules.scala 53:83:@25487.4]
  assign buffer_6_625 = $signed(_T_75800); // @[Modules.scala 53:83:@25488.4]
  assign _T_75802 = $signed(buffer_0_468) + $signed(buffer_6_469); // @[Modules.scala 53:83:@25490.4]
  assign _T_75803 = _T_75802[10:0]; // @[Modules.scala 53:83:@25491.4]
  assign buffer_6_626 = $signed(_T_75803); // @[Modules.scala 53:83:@25492.4]
  assign _T_75805 = $signed(buffer_6_470) + $signed(buffer_6_471); // @[Modules.scala 53:83:@25494.4]
  assign _T_75806 = _T_75805[10:0]; // @[Modules.scala 53:83:@25495.4]
  assign buffer_6_627 = $signed(_T_75806); // @[Modules.scala 53:83:@25496.4]
  assign _T_75808 = $signed(buffer_6_472) + $signed(buffer_6_473); // @[Modules.scala 53:83:@25498.4]
  assign _T_75809 = _T_75808[10:0]; // @[Modules.scala 53:83:@25499.4]
  assign buffer_6_628 = $signed(_T_75809); // @[Modules.scala 53:83:@25500.4]
  assign _T_75811 = $signed(buffer_0_474) + $signed(buffer_6_475); // @[Modules.scala 53:83:@25502.4]
  assign _T_75812 = _T_75811[10:0]; // @[Modules.scala 53:83:@25503.4]
  assign buffer_6_629 = $signed(_T_75812); // @[Modules.scala 53:83:@25504.4]
  assign _T_75814 = $signed(buffer_6_476) + $signed(buffer_6_477); // @[Modules.scala 53:83:@25506.4]
  assign _T_75815 = _T_75814[10:0]; // @[Modules.scala 53:83:@25507.4]
  assign buffer_6_630 = $signed(_T_75815); // @[Modules.scala 53:83:@25508.4]
  assign _T_75817 = $signed(buffer_6_478) + $signed(buffer_6_479); // @[Modules.scala 53:83:@25510.4]
  assign _T_75818 = _T_75817[10:0]; // @[Modules.scala 53:83:@25511.4]
  assign buffer_6_631 = $signed(_T_75818); // @[Modules.scala 53:83:@25512.4]
  assign _T_75820 = $signed(buffer_0_480) + $signed(buffer_6_481); // @[Modules.scala 53:83:@25514.4]
  assign _T_75821 = _T_75820[10:0]; // @[Modules.scala 53:83:@25515.4]
  assign buffer_6_632 = $signed(_T_75821); // @[Modules.scala 53:83:@25516.4]
  assign _T_75823 = $signed(buffer_0_482) + $signed(buffer_6_483); // @[Modules.scala 53:83:@25518.4]
  assign _T_75824 = _T_75823[10:0]; // @[Modules.scala 53:83:@25519.4]
  assign buffer_6_633 = $signed(_T_75824); // @[Modules.scala 53:83:@25520.4]
  assign _T_75826 = $signed(buffer_0_484) + $signed(buffer_6_485); // @[Modules.scala 53:83:@25522.4]
  assign _T_75827 = _T_75826[10:0]; // @[Modules.scala 53:83:@25523.4]
  assign buffer_6_634 = $signed(_T_75827); // @[Modules.scala 53:83:@25524.4]
  assign _T_75829 = $signed(buffer_6_486) + $signed(buffer_0_487); // @[Modules.scala 53:83:@25526.4]
  assign _T_75830 = _T_75829[10:0]; // @[Modules.scala 53:83:@25527.4]
  assign buffer_6_635 = $signed(_T_75830); // @[Modules.scala 53:83:@25528.4]
  assign _T_75832 = $signed(buffer_2_488) + $signed(buffer_5_489); // @[Modules.scala 53:83:@25530.4]
  assign _T_75833 = _T_75832[10:0]; // @[Modules.scala 53:83:@25531.4]
  assign buffer_6_636 = $signed(_T_75833); // @[Modules.scala 53:83:@25532.4]
  assign _T_75835 = $signed(buffer_6_490) + $signed(buffer_0_491); // @[Modules.scala 53:83:@25534.4]
  assign _T_75836 = _T_75835[10:0]; // @[Modules.scala 53:83:@25535.4]
  assign buffer_6_637 = $signed(_T_75836); // @[Modules.scala 53:83:@25536.4]
  assign _T_75838 = $signed(buffer_6_492) + $signed(buffer_6_493); // @[Modules.scala 53:83:@25538.4]
  assign _T_75839 = _T_75838[10:0]; // @[Modules.scala 53:83:@25539.4]
  assign buffer_6_638 = $signed(_T_75839); // @[Modules.scala 53:83:@25540.4]
  assign _T_75841 = $signed(buffer_0_494) + $signed(buffer_6_495); // @[Modules.scala 53:83:@25542.4]
  assign _T_75842 = _T_75841[10:0]; // @[Modules.scala 53:83:@25543.4]
  assign buffer_6_639 = $signed(_T_75842); // @[Modules.scala 53:83:@25544.4]
  assign _T_75844 = $signed(buffer_6_496) + $signed(buffer_6_497); // @[Modules.scala 53:83:@25546.4]
  assign _T_75845 = _T_75844[10:0]; // @[Modules.scala 53:83:@25547.4]
  assign buffer_6_640 = $signed(_T_75845); // @[Modules.scala 53:83:@25548.4]
  assign _T_75847 = $signed(buffer_6_498) + $signed(buffer_6_499); // @[Modules.scala 53:83:@25550.4]
  assign _T_75848 = _T_75847[10:0]; // @[Modules.scala 53:83:@25551.4]
  assign buffer_6_641 = $signed(_T_75848); // @[Modules.scala 53:83:@25552.4]
  assign _T_75850 = $signed(buffer_6_500) + $signed(buffer_6_501); // @[Modules.scala 53:83:@25554.4]
  assign _T_75851 = _T_75850[10:0]; // @[Modules.scala 53:83:@25555.4]
  assign buffer_6_642 = $signed(_T_75851); // @[Modules.scala 53:83:@25556.4]
  assign _T_75853 = $signed(buffer_6_502) + $signed(buffer_0_503); // @[Modules.scala 53:83:@25558.4]
  assign _T_75854 = _T_75853[10:0]; // @[Modules.scala 53:83:@25559.4]
  assign buffer_6_643 = $signed(_T_75854); // @[Modules.scala 53:83:@25560.4]
  assign _T_75856 = $signed(buffer_6_504) + $signed(buffer_3_505); // @[Modules.scala 53:83:@25562.4]
  assign _T_75857 = _T_75856[10:0]; // @[Modules.scala 53:83:@25563.4]
  assign buffer_6_644 = $signed(_T_75857); // @[Modules.scala 53:83:@25564.4]
  assign _T_75859 = $signed(buffer_6_506) + $signed(buffer_6_507); // @[Modules.scala 53:83:@25566.4]
  assign _T_75860 = _T_75859[10:0]; // @[Modules.scala 53:83:@25567.4]
  assign buffer_6_645 = $signed(_T_75860); // @[Modules.scala 53:83:@25568.4]
  assign _T_75862 = $signed(buffer_6_508) + $signed(buffer_6_509); // @[Modules.scala 53:83:@25570.4]
  assign _T_75863 = _T_75862[10:0]; // @[Modules.scala 53:83:@25571.4]
  assign buffer_6_646 = $signed(_T_75863); // @[Modules.scala 53:83:@25572.4]
  assign _T_75865 = $signed(buffer_0_510) + $signed(buffer_6_511); // @[Modules.scala 53:83:@25574.4]
  assign _T_75866 = _T_75865[10:0]; // @[Modules.scala 53:83:@25575.4]
  assign buffer_6_647 = $signed(_T_75866); // @[Modules.scala 53:83:@25576.4]
  assign _T_75868 = $signed(buffer_6_512) + $signed(buffer_6_513); // @[Modules.scala 53:83:@25578.4]
  assign _T_75869 = _T_75868[10:0]; // @[Modules.scala 53:83:@25579.4]
  assign buffer_6_648 = $signed(_T_75869); // @[Modules.scala 53:83:@25580.4]
  assign _T_75871 = $signed(buffer_2_514) + $signed(buffer_6_515); // @[Modules.scala 53:83:@25582.4]
  assign _T_75872 = _T_75871[10:0]; // @[Modules.scala 53:83:@25583.4]
  assign buffer_6_649 = $signed(_T_75872); // @[Modules.scala 53:83:@25584.4]
  assign _T_75874 = $signed(buffer_5_516) + $signed(buffer_0_517); // @[Modules.scala 53:83:@25586.4]
  assign _T_75875 = _T_75874[10:0]; // @[Modules.scala 53:83:@25587.4]
  assign buffer_6_650 = $signed(_T_75875); // @[Modules.scala 53:83:@25588.4]
  assign _T_75877 = $signed(buffer_6_518) + $signed(buffer_0_519); // @[Modules.scala 53:83:@25590.4]
  assign _T_75878 = _T_75877[10:0]; // @[Modules.scala 53:83:@25591.4]
  assign buffer_6_651 = $signed(_T_75878); // @[Modules.scala 53:83:@25592.4]
  assign _T_75880 = $signed(buffer_3_520) + $signed(buffer_6_521); // @[Modules.scala 53:83:@25594.4]
  assign _T_75881 = _T_75880[10:0]; // @[Modules.scala 53:83:@25595.4]
  assign buffer_6_652 = $signed(_T_75881); // @[Modules.scala 53:83:@25596.4]
  assign _T_75883 = $signed(buffer_6_522) + $signed(buffer_2_523); // @[Modules.scala 53:83:@25598.4]
  assign _T_75884 = _T_75883[10:0]; // @[Modules.scala 53:83:@25599.4]
  assign buffer_6_653 = $signed(_T_75884); // @[Modules.scala 53:83:@25600.4]
  assign _T_75889 = $signed(buffer_0_526) + $signed(buffer_6_527); // @[Modules.scala 53:83:@25606.4]
  assign _T_75890 = _T_75889[10:0]; // @[Modules.scala 53:83:@25607.4]
  assign buffer_6_655 = $signed(_T_75890); // @[Modules.scala 53:83:@25608.4]
  assign _T_75892 = $signed(buffer_0_528) + $signed(buffer_3_529); // @[Modules.scala 53:83:@25610.4]
  assign _T_75893 = _T_75892[10:0]; // @[Modules.scala 53:83:@25611.4]
  assign buffer_6_656 = $signed(_T_75893); // @[Modules.scala 53:83:@25612.4]
  assign _T_75895 = $signed(buffer_6_530) + $signed(buffer_2_531); // @[Modules.scala 53:83:@25614.4]
  assign _T_75896 = _T_75895[10:0]; // @[Modules.scala 53:83:@25615.4]
  assign buffer_6_657 = $signed(_T_75896); // @[Modules.scala 53:83:@25616.4]
  assign _T_75904 = $signed(buffer_6_536) + $signed(buffer_2_537); // @[Modules.scala 53:83:@25626.4]
  assign _T_75905 = _T_75904[10:0]; // @[Modules.scala 53:83:@25627.4]
  assign buffer_6_660 = $signed(_T_75905); // @[Modules.scala 53:83:@25628.4]
  assign _T_75907 = $signed(buffer_6_538) + $signed(buffer_6_539); // @[Modules.scala 53:83:@25630.4]
  assign _T_75908 = _T_75907[10:0]; // @[Modules.scala 53:83:@25631.4]
  assign buffer_6_661 = $signed(_T_75908); // @[Modules.scala 53:83:@25632.4]
  assign _T_75913 = $signed(buffer_5_542) + $signed(buffer_6_543); // @[Modules.scala 53:83:@25638.4]
  assign _T_75914 = _T_75913[10:0]; // @[Modules.scala 53:83:@25639.4]
  assign buffer_6_663 = $signed(_T_75914); // @[Modules.scala 53:83:@25640.4]
  assign _T_75916 = $signed(buffer_0_544) + $signed(buffer_6_545); // @[Modules.scala 53:83:@25642.4]
  assign _T_75917 = _T_75916[10:0]; // @[Modules.scala 53:83:@25643.4]
  assign buffer_6_664 = $signed(_T_75917); // @[Modules.scala 53:83:@25644.4]
  assign _T_75922 = $signed(buffer_6_548) + $signed(buffer_6_549); // @[Modules.scala 53:83:@25650.4]
  assign _T_75923 = _T_75922[10:0]; // @[Modules.scala 53:83:@25651.4]
  assign buffer_6_666 = $signed(_T_75923); // @[Modules.scala 53:83:@25652.4]
  assign _T_75925 = $signed(buffer_0_550) + $signed(buffer_6_551); // @[Modules.scala 53:83:@25654.4]
  assign _T_75926 = _T_75925[10:0]; // @[Modules.scala 53:83:@25655.4]
  assign buffer_6_667 = $signed(_T_75926); // @[Modules.scala 53:83:@25656.4]
  assign _T_75928 = $signed(buffer_0_552) + $signed(buffer_6_553); // @[Modules.scala 53:83:@25658.4]
  assign _T_75929 = _T_75928[10:0]; // @[Modules.scala 53:83:@25659.4]
  assign buffer_6_668 = $signed(_T_75929); // @[Modules.scala 53:83:@25660.4]
  assign _T_75931 = $signed(buffer_6_554) + $signed(buffer_6_555); // @[Modules.scala 53:83:@25662.4]
  assign _T_75932 = _T_75931[10:0]; // @[Modules.scala 53:83:@25663.4]
  assign buffer_6_669 = $signed(_T_75932); // @[Modules.scala 53:83:@25664.4]
  assign _T_75934 = $signed(buffer_0_556) + $signed(buffer_3_557); // @[Modules.scala 53:83:@25666.4]
  assign _T_75935 = _T_75934[10:0]; // @[Modules.scala 53:83:@25667.4]
  assign buffer_6_670 = $signed(_T_75935); // @[Modules.scala 53:83:@25668.4]
  assign _T_75937 = $signed(buffer_1_558) + $signed(buffer_6_559); // @[Modules.scala 53:83:@25670.4]
  assign _T_75938 = _T_75937[10:0]; // @[Modules.scala 53:83:@25671.4]
  assign buffer_6_671 = $signed(_T_75938); // @[Modules.scala 53:83:@25672.4]
  assign _T_75940 = $signed(buffer_6_560) + $signed(buffer_5_561); // @[Modules.scala 53:83:@25674.4]
  assign _T_75941 = _T_75940[10:0]; // @[Modules.scala 53:83:@25675.4]
  assign buffer_6_672 = $signed(_T_75941); // @[Modules.scala 53:83:@25676.4]
  assign _T_75943 = $signed(buffer_2_562) + $signed(buffer_0_563); // @[Modules.scala 53:83:@25678.4]
  assign _T_75944 = _T_75943[10:0]; // @[Modules.scala 53:83:@25679.4]
  assign buffer_6_673 = $signed(_T_75944); // @[Modules.scala 53:83:@25680.4]
  assign _T_75946 = $signed(buffer_6_564) + $signed(buffer_6_565); // @[Modules.scala 53:83:@25682.4]
  assign _T_75947 = _T_75946[10:0]; // @[Modules.scala 53:83:@25683.4]
  assign buffer_6_674 = $signed(_T_75947); // @[Modules.scala 53:83:@25684.4]
  assign _T_75949 = $signed(buffer_2_566) + $signed(buffer_3_567); // @[Modules.scala 53:83:@25686.4]
  assign _T_75950 = _T_75949[10:0]; // @[Modules.scala 53:83:@25687.4]
  assign buffer_6_675 = $signed(_T_75950); // @[Modules.scala 53:83:@25688.4]
  assign _T_75952 = $signed(buffer_0_568) + $signed(buffer_6_569); // @[Modules.scala 53:83:@25690.4]
  assign _T_75953 = _T_75952[10:0]; // @[Modules.scala 53:83:@25691.4]
  assign buffer_6_676 = $signed(_T_75953); // @[Modules.scala 53:83:@25692.4]
  assign _T_75955 = $signed(buffer_6_570) + $signed(buffer_6_571); // @[Modules.scala 53:83:@25694.4]
  assign _T_75956 = _T_75955[10:0]; // @[Modules.scala 53:83:@25695.4]
  assign buffer_6_677 = $signed(_T_75956); // @[Modules.scala 53:83:@25696.4]
  assign _T_75958 = $signed(buffer_0_572) + $signed(buffer_6_573); // @[Modules.scala 53:83:@25698.4]
  assign _T_75959 = _T_75958[10:0]; // @[Modules.scala 53:83:@25699.4]
  assign buffer_6_678 = $signed(_T_75959); // @[Modules.scala 53:83:@25700.4]
  assign _T_75961 = $signed(buffer_6_574) + $signed(buffer_0_575); // @[Modules.scala 53:83:@25702.4]
  assign _T_75962 = _T_75961[10:0]; // @[Modules.scala 53:83:@25703.4]
  assign buffer_6_679 = $signed(_T_75962); // @[Modules.scala 53:83:@25704.4]
  assign _T_75967 = $signed(buffer_3_578) + $signed(buffer_6_579); // @[Modules.scala 53:83:@25710.4]
  assign _T_75968 = _T_75967[10:0]; // @[Modules.scala 53:83:@25711.4]
  assign buffer_6_681 = $signed(_T_75968); // @[Modules.scala 53:83:@25712.4]
  assign _T_75970 = $signed(buffer_3_580) + $signed(buffer_4_581); // @[Modules.scala 53:83:@25714.4]
  assign _T_75971 = _T_75970[10:0]; // @[Modules.scala 53:83:@25715.4]
  assign buffer_6_682 = $signed(_T_75971); // @[Modules.scala 53:83:@25716.4]
  assign _T_75973 = $signed(buffer_5_582) + $signed(buffer_0_583); // @[Modules.scala 53:83:@25718.4]
  assign _T_75974 = _T_75973[10:0]; // @[Modules.scala 53:83:@25719.4]
  assign buffer_6_683 = $signed(_T_75974); // @[Modules.scala 53:83:@25720.4]
  assign _T_75976 = $signed(buffer_6_584) + $signed(buffer_0_585); // @[Modules.scala 53:83:@25722.4]
  assign _T_75977 = _T_75976[10:0]; // @[Modules.scala 53:83:@25723.4]
  assign buffer_6_684 = $signed(_T_75977); // @[Modules.scala 53:83:@25724.4]
  assign _T_75979 = $signed(buffer_6_586) + $signed(buffer_4_587); // @[Modules.scala 53:83:@25726.4]
  assign _T_75980 = _T_75979[10:0]; // @[Modules.scala 53:83:@25727.4]
  assign buffer_6_685 = $signed(_T_75980); // @[Modules.scala 53:83:@25728.4]
  assign _T_75982 = $signed(buffer_6_588) + $signed(buffer_6_589); // @[Modules.scala 56:109:@25730.4]
  assign _T_75983 = _T_75982[10:0]; // @[Modules.scala 56:109:@25731.4]
  assign buffer_6_686 = $signed(_T_75983); // @[Modules.scala 56:109:@25732.4]
  assign _T_75985 = $signed(buffer_6_590) + $signed(buffer_6_591); // @[Modules.scala 56:109:@25734.4]
  assign _T_75986 = _T_75985[10:0]; // @[Modules.scala 56:109:@25735.4]
  assign buffer_6_687 = $signed(_T_75986); // @[Modules.scala 56:109:@25736.4]
  assign _T_75988 = $signed(buffer_6_592) + $signed(buffer_0_593); // @[Modules.scala 56:109:@25738.4]
  assign _T_75989 = _T_75988[10:0]; // @[Modules.scala 56:109:@25739.4]
  assign buffer_6_688 = $signed(_T_75989); // @[Modules.scala 56:109:@25740.4]
  assign _T_75991 = $signed(buffer_6_594) + $signed(buffer_6_595); // @[Modules.scala 56:109:@25742.4]
  assign _T_75992 = _T_75991[10:0]; // @[Modules.scala 56:109:@25743.4]
  assign buffer_6_689 = $signed(_T_75992); // @[Modules.scala 56:109:@25744.4]
  assign _T_75997 = $signed(buffer_6_598) + $signed(buffer_6_599); // @[Modules.scala 56:109:@25750.4]
  assign _T_75998 = _T_75997[10:0]; // @[Modules.scala 56:109:@25751.4]
  assign buffer_6_691 = $signed(_T_75998); // @[Modules.scala 56:109:@25752.4]
  assign _T_76000 = $signed(buffer_6_600) + $signed(buffer_6_601); // @[Modules.scala 56:109:@25754.4]
  assign _T_76001 = _T_76000[10:0]; // @[Modules.scala 56:109:@25755.4]
  assign buffer_6_692 = $signed(_T_76001); // @[Modules.scala 56:109:@25756.4]
  assign _T_76003 = $signed(buffer_6_602) + $signed(buffer_0_603); // @[Modules.scala 56:109:@25758.4]
  assign _T_76004 = _T_76003[10:0]; // @[Modules.scala 56:109:@25759.4]
  assign buffer_6_693 = $signed(_T_76004); // @[Modules.scala 56:109:@25760.4]
  assign _T_76006 = $signed(buffer_6_604) + $signed(buffer_6_605); // @[Modules.scala 56:109:@25762.4]
  assign _T_76007 = _T_76006[10:0]; // @[Modules.scala 56:109:@25763.4]
  assign buffer_6_694 = $signed(_T_76007); // @[Modules.scala 56:109:@25764.4]
  assign _T_76009 = $signed(buffer_6_606) + $signed(buffer_0_607); // @[Modules.scala 56:109:@25766.4]
  assign _T_76010 = _T_76009[10:0]; // @[Modules.scala 56:109:@25767.4]
  assign buffer_6_695 = $signed(_T_76010); // @[Modules.scala 56:109:@25768.4]
  assign _T_76012 = $signed(buffer_6_608) + $signed(buffer_6_609); // @[Modules.scala 56:109:@25770.4]
  assign _T_76013 = _T_76012[10:0]; // @[Modules.scala 56:109:@25771.4]
  assign buffer_6_696 = $signed(_T_76013); // @[Modules.scala 56:109:@25772.4]
  assign _T_76015 = $signed(buffer_6_610) + $signed(buffer_6_611); // @[Modules.scala 56:109:@25774.4]
  assign _T_76016 = _T_76015[10:0]; // @[Modules.scala 56:109:@25775.4]
  assign buffer_6_697 = $signed(_T_76016); // @[Modules.scala 56:109:@25776.4]
  assign _T_76018 = $signed(buffer_6_612) + $signed(buffer_6_613); // @[Modules.scala 56:109:@25778.4]
  assign _T_76019 = _T_76018[10:0]; // @[Modules.scala 56:109:@25779.4]
  assign buffer_6_698 = $signed(_T_76019); // @[Modules.scala 56:109:@25780.4]
  assign _T_76021 = $signed(buffer_6_614) + $signed(buffer_6_615); // @[Modules.scala 56:109:@25782.4]
  assign _T_76022 = _T_76021[10:0]; // @[Modules.scala 56:109:@25783.4]
  assign buffer_6_699 = $signed(_T_76022); // @[Modules.scala 56:109:@25784.4]
  assign _T_76024 = $signed(buffer_6_616) + $signed(buffer_6_617); // @[Modules.scala 56:109:@25786.4]
  assign _T_76025 = _T_76024[10:0]; // @[Modules.scala 56:109:@25787.4]
  assign buffer_6_700 = $signed(_T_76025); // @[Modules.scala 56:109:@25788.4]
  assign _T_76027 = $signed(buffer_6_618) + $signed(buffer_6_619); // @[Modules.scala 56:109:@25790.4]
  assign _T_76028 = _T_76027[10:0]; // @[Modules.scala 56:109:@25791.4]
  assign buffer_6_701 = $signed(_T_76028); // @[Modules.scala 56:109:@25792.4]
  assign _T_76030 = $signed(buffer_6_620) + $signed(buffer_3_621); // @[Modules.scala 56:109:@25794.4]
  assign _T_76031 = _T_76030[10:0]; // @[Modules.scala 56:109:@25795.4]
  assign buffer_6_702 = $signed(_T_76031); // @[Modules.scala 56:109:@25796.4]
  assign _T_76033 = $signed(buffer_6_622) + $signed(buffer_6_623); // @[Modules.scala 56:109:@25798.4]
  assign _T_76034 = _T_76033[10:0]; // @[Modules.scala 56:109:@25799.4]
  assign buffer_6_703 = $signed(_T_76034); // @[Modules.scala 56:109:@25800.4]
  assign _T_76036 = $signed(buffer_6_624) + $signed(buffer_6_625); // @[Modules.scala 56:109:@25802.4]
  assign _T_76037 = _T_76036[10:0]; // @[Modules.scala 56:109:@25803.4]
  assign buffer_6_704 = $signed(_T_76037); // @[Modules.scala 56:109:@25804.4]
  assign _T_76039 = $signed(buffer_6_626) + $signed(buffer_6_627); // @[Modules.scala 56:109:@25806.4]
  assign _T_76040 = _T_76039[10:0]; // @[Modules.scala 56:109:@25807.4]
  assign buffer_6_705 = $signed(_T_76040); // @[Modules.scala 56:109:@25808.4]
  assign _T_76042 = $signed(buffer_6_628) + $signed(buffer_6_629); // @[Modules.scala 56:109:@25810.4]
  assign _T_76043 = _T_76042[10:0]; // @[Modules.scala 56:109:@25811.4]
  assign buffer_6_706 = $signed(_T_76043); // @[Modules.scala 56:109:@25812.4]
  assign _T_76045 = $signed(buffer_6_630) + $signed(buffer_6_631); // @[Modules.scala 56:109:@25814.4]
  assign _T_76046 = _T_76045[10:0]; // @[Modules.scala 56:109:@25815.4]
  assign buffer_6_707 = $signed(_T_76046); // @[Modules.scala 56:109:@25816.4]
  assign _T_76048 = $signed(buffer_6_632) + $signed(buffer_6_633); // @[Modules.scala 56:109:@25818.4]
  assign _T_76049 = _T_76048[10:0]; // @[Modules.scala 56:109:@25819.4]
  assign buffer_6_708 = $signed(_T_76049); // @[Modules.scala 56:109:@25820.4]
  assign _T_76051 = $signed(buffer_6_634) + $signed(buffer_6_635); // @[Modules.scala 56:109:@25822.4]
  assign _T_76052 = _T_76051[10:0]; // @[Modules.scala 56:109:@25823.4]
  assign buffer_6_709 = $signed(_T_76052); // @[Modules.scala 56:109:@25824.4]
  assign _T_76054 = $signed(buffer_6_636) + $signed(buffer_6_637); // @[Modules.scala 56:109:@25826.4]
  assign _T_76055 = _T_76054[10:0]; // @[Modules.scala 56:109:@25827.4]
  assign buffer_6_710 = $signed(_T_76055); // @[Modules.scala 56:109:@25828.4]
  assign _T_76057 = $signed(buffer_6_638) + $signed(buffer_6_639); // @[Modules.scala 56:109:@25830.4]
  assign _T_76058 = _T_76057[10:0]; // @[Modules.scala 56:109:@25831.4]
  assign buffer_6_711 = $signed(_T_76058); // @[Modules.scala 56:109:@25832.4]
  assign _T_76060 = $signed(buffer_6_640) + $signed(buffer_6_641); // @[Modules.scala 56:109:@25834.4]
  assign _T_76061 = _T_76060[10:0]; // @[Modules.scala 56:109:@25835.4]
  assign buffer_6_712 = $signed(_T_76061); // @[Modules.scala 56:109:@25836.4]
  assign _T_76063 = $signed(buffer_6_642) + $signed(buffer_6_643); // @[Modules.scala 56:109:@25838.4]
  assign _T_76064 = _T_76063[10:0]; // @[Modules.scala 56:109:@25839.4]
  assign buffer_6_713 = $signed(_T_76064); // @[Modules.scala 56:109:@25840.4]
  assign _T_76066 = $signed(buffer_6_644) + $signed(buffer_6_645); // @[Modules.scala 56:109:@25842.4]
  assign _T_76067 = _T_76066[10:0]; // @[Modules.scala 56:109:@25843.4]
  assign buffer_6_714 = $signed(_T_76067); // @[Modules.scala 56:109:@25844.4]
  assign _T_76069 = $signed(buffer_6_646) + $signed(buffer_6_647); // @[Modules.scala 56:109:@25846.4]
  assign _T_76070 = _T_76069[10:0]; // @[Modules.scala 56:109:@25847.4]
  assign buffer_6_715 = $signed(_T_76070); // @[Modules.scala 56:109:@25848.4]
  assign _T_76072 = $signed(buffer_6_648) + $signed(buffer_6_649); // @[Modules.scala 56:109:@25850.4]
  assign _T_76073 = _T_76072[10:0]; // @[Modules.scala 56:109:@25851.4]
  assign buffer_6_716 = $signed(_T_76073); // @[Modules.scala 56:109:@25852.4]
  assign _T_76075 = $signed(buffer_6_650) + $signed(buffer_6_651); // @[Modules.scala 56:109:@25854.4]
  assign _T_76076 = _T_76075[10:0]; // @[Modules.scala 56:109:@25855.4]
  assign buffer_6_717 = $signed(_T_76076); // @[Modules.scala 56:109:@25856.4]
  assign _T_76078 = $signed(buffer_6_652) + $signed(buffer_6_653); // @[Modules.scala 56:109:@25858.4]
  assign _T_76079 = _T_76078[10:0]; // @[Modules.scala 56:109:@25859.4]
  assign buffer_6_718 = $signed(_T_76079); // @[Modules.scala 56:109:@25860.4]
  assign _T_76081 = $signed(buffer_2_654) + $signed(buffer_6_655); // @[Modules.scala 56:109:@25862.4]
  assign _T_76082 = _T_76081[10:0]; // @[Modules.scala 56:109:@25863.4]
  assign buffer_6_719 = $signed(_T_76082); // @[Modules.scala 56:109:@25864.4]
  assign _T_76084 = $signed(buffer_6_656) + $signed(buffer_6_657); // @[Modules.scala 56:109:@25866.4]
  assign _T_76085 = _T_76084[10:0]; // @[Modules.scala 56:109:@25867.4]
  assign buffer_6_720 = $signed(_T_76085); // @[Modules.scala 56:109:@25868.4]
  assign _T_76087 = $signed(buffer_0_658) + $signed(buffer_5_659); // @[Modules.scala 56:109:@25870.4]
  assign _T_76088 = _T_76087[10:0]; // @[Modules.scala 56:109:@25871.4]
  assign buffer_6_721 = $signed(_T_76088); // @[Modules.scala 56:109:@25872.4]
  assign _T_76090 = $signed(buffer_6_660) + $signed(buffer_6_661); // @[Modules.scala 56:109:@25874.4]
  assign _T_76091 = _T_76090[10:0]; // @[Modules.scala 56:109:@25875.4]
  assign buffer_6_722 = $signed(_T_76091); // @[Modules.scala 56:109:@25876.4]
  assign _T_76093 = $signed(buffer_0_662) + $signed(buffer_6_663); // @[Modules.scala 56:109:@25878.4]
  assign _T_76094 = _T_76093[10:0]; // @[Modules.scala 56:109:@25879.4]
  assign buffer_6_723 = $signed(_T_76094); // @[Modules.scala 56:109:@25880.4]
  assign _T_76096 = $signed(buffer_6_664) + $signed(buffer_2_665); // @[Modules.scala 56:109:@25882.4]
  assign _T_76097 = _T_76096[10:0]; // @[Modules.scala 56:109:@25883.4]
  assign buffer_6_724 = $signed(_T_76097); // @[Modules.scala 56:109:@25884.4]
  assign _T_76099 = $signed(buffer_6_666) + $signed(buffer_6_667); // @[Modules.scala 56:109:@25886.4]
  assign _T_76100 = _T_76099[10:0]; // @[Modules.scala 56:109:@25887.4]
  assign buffer_6_725 = $signed(_T_76100); // @[Modules.scala 56:109:@25888.4]
  assign _T_76102 = $signed(buffer_6_668) + $signed(buffer_6_669); // @[Modules.scala 56:109:@25890.4]
  assign _T_76103 = _T_76102[10:0]; // @[Modules.scala 56:109:@25891.4]
  assign buffer_6_726 = $signed(_T_76103); // @[Modules.scala 56:109:@25892.4]
  assign _T_76105 = $signed(buffer_6_670) + $signed(buffer_6_671); // @[Modules.scala 56:109:@25894.4]
  assign _T_76106 = _T_76105[10:0]; // @[Modules.scala 56:109:@25895.4]
  assign buffer_6_727 = $signed(_T_76106); // @[Modules.scala 56:109:@25896.4]
  assign _T_76108 = $signed(buffer_6_672) + $signed(buffer_6_673); // @[Modules.scala 56:109:@25898.4]
  assign _T_76109 = _T_76108[10:0]; // @[Modules.scala 56:109:@25899.4]
  assign buffer_6_728 = $signed(_T_76109); // @[Modules.scala 56:109:@25900.4]
  assign _T_76111 = $signed(buffer_6_674) + $signed(buffer_6_675); // @[Modules.scala 56:109:@25902.4]
  assign _T_76112 = _T_76111[10:0]; // @[Modules.scala 56:109:@25903.4]
  assign buffer_6_729 = $signed(_T_76112); // @[Modules.scala 56:109:@25904.4]
  assign _T_76114 = $signed(buffer_6_676) + $signed(buffer_6_677); // @[Modules.scala 56:109:@25906.4]
  assign _T_76115 = _T_76114[10:0]; // @[Modules.scala 56:109:@25907.4]
  assign buffer_6_730 = $signed(_T_76115); // @[Modules.scala 56:109:@25908.4]
  assign _T_76117 = $signed(buffer_6_678) + $signed(buffer_6_679); // @[Modules.scala 56:109:@25910.4]
  assign _T_76118 = _T_76117[10:0]; // @[Modules.scala 56:109:@25911.4]
  assign buffer_6_731 = $signed(_T_76118); // @[Modules.scala 56:109:@25912.4]
  assign _T_76120 = $signed(buffer_5_680) + $signed(buffer_6_681); // @[Modules.scala 56:109:@25914.4]
  assign _T_76121 = _T_76120[10:0]; // @[Modules.scala 56:109:@25915.4]
  assign buffer_6_732 = $signed(_T_76121); // @[Modules.scala 56:109:@25916.4]
  assign _T_76123 = $signed(buffer_6_682) + $signed(buffer_6_683); // @[Modules.scala 56:109:@25918.4]
  assign _T_76124 = _T_76123[10:0]; // @[Modules.scala 56:109:@25919.4]
  assign buffer_6_733 = $signed(_T_76124); // @[Modules.scala 56:109:@25920.4]
  assign _T_76126 = $signed(buffer_6_684) + $signed(buffer_6_685); // @[Modules.scala 56:109:@25922.4]
  assign _T_76127 = _T_76126[10:0]; // @[Modules.scala 56:109:@25923.4]
  assign buffer_6_734 = $signed(_T_76127); // @[Modules.scala 56:109:@25924.4]
  assign _T_76129 = $signed(buffer_6_686) + $signed(buffer_6_687); // @[Modules.scala 63:156:@25927.4]
  assign _T_76130 = _T_76129[10:0]; // @[Modules.scala 63:156:@25928.4]
  assign buffer_6_736 = $signed(_T_76130); // @[Modules.scala 63:156:@25929.4]
  assign _T_76132 = $signed(buffer_6_736) + $signed(buffer_6_688); // @[Modules.scala 63:156:@25931.4]
  assign _T_76133 = _T_76132[10:0]; // @[Modules.scala 63:156:@25932.4]
  assign buffer_6_737 = $signed(_T_76133); // @[Modules.scala 63:156:@25933.4]
  assign _T_76135 = $signed(buffer_6_737) + $signed(buffer_6_689); // @[Modules.scala 63:156:@25935.4]
  assign _T_76136 = _T_76135[10:0]; // @[Modules.scala 63:156:@25936.4]
  assign buffer_6_738 = $signed(_T_76136); // @[Modules.scala 63:156:@25937.4]
  assign _T_76138 = $signed(buffer_6_738) + $signed(buffer_3_690); // @[Modules.scala 63:156:@25939.4]
  assign _T_76139 = _T_76138[10:0]; // @[Modules.scala 63:156:@25940.4]
  assign buffer_6_739 = $signed(_T_76139); // @[Modules.scala 63:156:@25941.4]
  assign _T_76141 = $signed(buffer_6_739) + $signed(buffer_6_691); // @[Modules.scala 63:156:@25943.4]
  assign _T_76142 = _T_76141[10:0]; // @[Modules.scala 63:156:@25944.4]
  assign buffer_6_740 = $signed(_T_76142); // @[Modules.scala 63:156:@25945.4]
  assign _T_76144 = $signed(buffer_6_740) + $signed(buffer_6_692); // @[Modules.scala 63:156:@25947.4]
  assign _T_76145 = _T_76144[10:0]; // @[Modules.scala 63:156:@25948.4]
  assign buffer_6_741 = $signed(_T_76145); // @[Modules.scala 63:156:@25949.4]
  assign _T_76147 = $signed(buffer_6_741) + $signed(buffer_6_693); // @[Modules.scala 63:156:@25951.4]
  assign _T_76148 = _T_76147[10:0]; // @[Modules.scala 63:156:@25952.4]
  assign buffer_6_742 = $signed(_T_76148); // @[Modules.scala 63:156:@25953.4]
  assign _T_76150 = $signed(buffer_6_742) + $signed(buffer_6_694); // @[Modules.scala 63:156:@25955.4]
  assign _T_76151 = _T_76150[10:0]; // @[Modules.scala 63:156:@25956.4]
  assign buffer_6_743 = $signed(_T_76151); // @[Modules.scala 63:156:@25957.4]
  assign _T_76153 = $signed(buffer_6_743) + $signed(buffer_6_695); // @[Modules.scala 63:156:@25959.4]
  assign _T_76154 = _T_76153[10:0]; // @[Modules.scala 63:156:@25960.4]
  assign buffer_6_744 = $signed(_T_76154); // @[Modules.scala 63:156:@25961.4]
  assign _T_76156 = $signed(buffer_6_744) + $signed(buffer_6_696); // @[Modules.scala 63:156:@25963.4]
  assign _T_76157 = _T_76156[10:0]; // @[Modules.scala 63:156:@25964.4]
  assign buffer_6_745 = $signed(_T_76157); // @[Modules.scala 63:156:@25965.4]
  assign _T_76159 = $signed(buffer_6_745) + $signed(buffer_6_697); // @[Modules.scala 63:156:@25967.4]
  assign _T_76160 = _T_76159[10:0]; // @[Modules.scala 63:156:@25968.4]
  assign buffer_6_746 = $signed(_T_76160); // @[Modules.scala 63:156:@25969.4]
  assign _T_76162 = $signed(buffer_6_746) + $signed(buffer_6_698); // @[Modules.scala 63:156:@25971.4]
  assign _T_76163 = _T_76162[10:0]; // @[Modules.scala 63:156:@25972.4]
  assign buffer_6_747 = $signed(_T_76163); // @[Modules.scala 63:156:@25973.4]
  assign _T_76165 = $signed(buffer_6_747) + $signed(buffer_6_699); // @[Modules.scala 63:156:@25975.4]
  assign _T_76166 = _T_76165[10:0]; // @[Modules.scala 63:156:@25976.4]
  assign buffer_6_748 = $signed(_T_76166); // @[Modules.scala 63:156:@25977.4]
  assign _T_76168 = $signed(buffer_6_748) + $signed(buffer_6_700); // @[Modules.scala 63:156:@25979.4]
  assign _T_76169 = _T_76168[10:0]; // @[Modules.scala 63:156:@25980.4]
  assign buffer_6_749 = $signed(_T_76169); // @[Modules.scala 63:156:@25981.4]
  assign _T_76171 = $signed(buffer_6_749) + $signed(buffer_6_701); // @[Modules.scala 63:156:@25983.4]
  assign _T_76172 = _T_76171[10:0]; // @[Modules.scala 63:156:@25984.4]
  assign buffer_6_750 = $signed(_T_76172); // @[Modules.scala 63:156:@25985.4]
  assign _T_76174 = $signed(buffer_6_750) + $signed(buffer_6_702); // @[Modules.scala 63:156:@25987.4]
  assign _T_76175 = _T_76174[10:0]; // @[Modules.scala 63:156:@25988.4]
  assign buffer_6_751 = $signed(_T_76175); // @[Modules.scala 63:156:@25989.4]
  assign _T_76177 = $signed(buffer_6_751) + $signed(buffer_6_703); // @[Modules.scala 63:156:@25991.4]
  assign _T_76178 = _T_76177[10:0]; // @[Modules.scala 63:156:@25992.4]
  assign buffer_6_752 = $signed(_T_76178); // @[Modules.scala 63:156:@25993.4]
  assign _T_76180 = $signed(buffer_6_752) + $signed(buffer_6_704); // @[Modules.scala 63:156:@25995.4]
  assign _T_76181 = _T_76180[10:0]; // @[Modules.scala 63:156:@25996.4]
  assign buffer_6_753 = $signed(_T_76181); // @[Modules.scala 63:156:@25997.4]
  assign _T_76183 = $signed(buffer_6_753) + $signed(buffer_6_705); // @[Modules.scala 63:156:@25999.4]
  assign _T_76184 = _T_76183[10:0]; // @[Modules.scala 63:156:@26000.4]
  assign buffer_6_754 = $signed(_T_76184); // @[Modules.scala 63:156:@26001.4]
  assign _T_76186 = $signed(buffer_6_754) + $signed(buffer_6_706); // @[Modules.scala 63:156:@26003.4]
  assign _T_76187 = _T_76186[10:0]; // @[Modules.scala 63:156:@26004.4]
  assign buffer_6_755 = $signed(_T_76187); // @[Modules.scala 63:156:@26005.4]
  assign _T_76189 = $signed(buffer_6_755) + $signed(buffer_6_707); // @[Modules.scala 63:156:@26007.4]
  assign _T_76190 = _T_76189[10:0]; // @[Modules.scala 63:156:@26008.4]
  assign buffer_6_756 = $signed(_T_76190); // @[Modules.scala 63:156:@26009.4]
  assign _T_76192 = $signed(buffer_6_756) + $signed(buffer_6_708); // @[Modules.scala 63:156:@26011.4]
  assign _T_76193 = _T_76192[10:0]; // @[Modules.scala 63:156:@26012.4]
  assign buffer_6_757 = $signed(_T_76193); // @[Modules.scala 63:156:@26013.4]
  assign _T_76195 = $signed(buffer_6_757) + $signed(buffer_6_709); // @[Modules.scala 63:156:@26015.4]
  assign _T_76196 = _T_76195[10:0]; // @[Modules.scala 63:156:@26016.4]
  assign buffer_6_758 = $signed(_T_76196); // @[Modules.scala 63:156:@26017.4]
  assign _T_76198 = $signed(buffer_6_758) + $signed(buffer_6_710); // @[Modules.scala 63:156:@26019.4]
  assign _T_76199 = _T_76198[10:0]; // @[Modules.scala 63:156:@26020.4]
  assign buffer_6_759 = $signed(_T_76199); // @[Modules.scala 63:156:@26021.4]
  assign _T_76201 = $signed(buffer_6_759) + $signed(buffer_6_711); // @[Modules.scala 63:156:@26023.4]
  assign _T_76202 = _T_76201[10:0]; // @[Modules.scala 63:156:@26024.4]
  assign buffer_6_760 = $signed(_T_76202); // @[Modules.scala 63:156:@26025.4]
  assign _T_76204 = $signed(buffer_6_760) + $signed(buffer_6_712); // @[Modules.scala 63:156:@26027.4]
  assign _T_76205 = _T_76204[10:0]; // @[Modules.scala 63:156:@26028.4]
  assign buffer_6_761 = $signed(_T_76205); // @[Modules.scala 63:156:@26029.4]
  assign _T_76207 = $signed(buffer_6_761) + $signed(buffer_6_713); // @[Modules.scala 63:156:@26031.4]
  assign _T_76208 = _T_76207[10:0]; // @[Modules.scala 63:156:@26032.4]
  assign buffer_6_762 = $signed(_T_76208); // @[Modules.scala 63:156:@26033.4]
  assign _T_76210 = $signed(buffer_6_762) + $signed(buffer_6_714); // @[Modules.scala 63:156:@26035.4]
  assign _T_76211 = _T_76210[10:0]; // @[Modules.scala 63:156:@26036.4]
  assign buffer_6_763 = $signed(_T_76211); // @[Modules.scala 63:156:@26037.4]
  assign _T_76213 = $signed(buffer_6_763) + $signed(buffer_6_715); // @[Modules.scala 63:156:@26039.4]
  assign _T_76214 = _T_76213[10:0]; // @[Modules.scala 63:156:@26040.4]
  assign buffer_6_764 = $signed(_T_76214); // @[Modules.scala 63:156:@26041.4]
  assign _T_76216 = $signed(buffer_6_764) + $signed(buffer_6_716); // @[Modules.scala 63:156:@26043.4]
  assign _T_76217 = _T_76216[10:0]; // @[Modules.scala 63:156:@26044.4]
  assign buffer_6_765 = $signed(_T_76217); // @[Modules.scala 63:156:@26045.4]
  assign _T_76219 = $signed(buffer_6_765) + $signed(buffer_6_717); // @[Modules.scala 63:156:@26047.4]
  assign _T_76220 = _T_76219[10:0]; // @[Modules.scala 63:156:@26048.4]
  assign buffer_6_766 = $signed(_T_76220); // @[Modules.scala 63:156:@26049.4]
  assign _T_76222 = $signed(buffer_6_766) + $signed(buffer_6_718); // @[Modules.scala 63:156:@26051.4]
  assign _T_76223 = _T_76222[10:0]; // @[Modules.scala 63:156:@26052.4]
  assign buffer_6_767 = $signed(_T_76223); // @[Modules.scala 63:156:@26053.4]
  assign _T_76225 = $signed(buffer_6_767) + $signed(buffer_6_719); // @[Modules.scala 63:156:@26055.4]
  assign _T_76226 = _T_76225[10:0]; // @[Modules.scala 63:156:@26056.4]
  assign buffer_6_768 = $signed(_T_76226); // @[Modules.scala 63:156:@26057.4]
  assign _T_76228 = $signed(buffer_6_768) + $signed(buffer_6_720); // @[Modules.scala 63:156:@26059.4]
  assign _T_76229 = _T_76228[10:0]; // @[Modules.scala 63:156:@26060.4]
  assign buffer_6_769 = $signed(_T_76229); // @[Modules.scala 63:156:@26061.4]
  assign _T_76231 = $signed(buffer_6_769) + $signed(buffer_6_721); // @[Modules.scala 63:156:@26063.4]
  assign _T_76232 = _T_76231[10:0]; // @[Modules.scala 63:156:@26064.4]
  assign buffer_6_770 = $signed(_T_76232); // @[Modules.scala 63:156:@26065.4]
  assign _T_76234 = $signed(buffer_6_770) + $signed(buffer_6_722); // @[Modules.scala 63:156:@26067.4]
  assign _T_76235 = _T_76234[10:0]; // @[Modules.scala 63:156:@26068.4]
  assign buffer_6_771 = $signed(_T_76235); // @[Modules.scala 63:156:@26069.4]
  assign _T_76237 = $signed(buffer_6_771) + $signed(buffer_6_723); // @[Modules.scala 63:156:@26071.4]
  assign _T_76238 = _T_76237[10:0]; // @[Modules.scala 63:156:@26072.4]
  assign buffer_6_772 = $signed(_T_76238); // @[Modules.scala 63:156:@26073.4]
  assign _T_76240 = $signed(buffer_6_772) + $signed(buffer_6_724); // @[Modules.scala 63:156:@26075.4]
  assign _T_76241 = _T_76240[10:0]; // @[Modules.scala 63:156:@26076.4]
  assign buffer_6_773 = $signed(_T_76241); // @[Modules.scala 63:156:@26077.4]
  assign _T_76243 = $signed(buffer_6_773) + $signed(buffer_6_725); // @[Modules.scala 63:156:@26079.4]
  assign _T_76244 = _T_76243[10:0]; // @[Modules.scala 63:156:@26080.4]
  assign buffer_6_774 = $signed(_T_76244); // @[Modules.scala 63:156:@26081.4]
  assign _T_76246 = $signed(buffer_6_774) + $signed(buffer_6_726); // @[Modules.scala 63:156:@26083.4]
  assign _T_76247 = _T_76246[10:0]; // @[Modules.scala 63:156:@26084.4]
  assign buffer_6_775 = $signed(_T_76247); // @[Modules.scala 63:156:@26085.4]
  assign _T_76249 = $signed(buffer_6_775) + $signed(buffer_6_727); // @[Modules.scala 63:156:@26087.4]
  assign _T_76250 = _T_76249[10:0]; // @[Modules.scala 63:156:@26088.4]
  assign buffer_6_776 = $signed(_T_76250); // @[Modules.scala 63:156:@26089.4]
  assign _T_76252 = $signed(buffer_6_776) + $signed(buffer_6_728); // @[Modules.scala 63:156:@26091.4]
  assign _T_76253 = _T_76252[10:0]; // @[Modules.scala 63:156:@26092.4]
  assign buffer_6_777 = $signed(_T_76253); // @[Modules.scala 63:156:@26093.4]
  assign _T_76255 = $signed(buffer_6_777) + $signed(buffer_6_729); // @[Modules.scala 63:156:@26095.4]
  assign _T_76256 = _T_76255[10:0]; // @[Modules.scala 63:156:@26096.4]
  assign buffer_6_778 = $signed(_T_76256); // @[Modules.scala 63:156:@26097.4]
  assign _T_76258 = $signed(buffer_6_778) + $signed(buffer_6_730); // @[Modules.scala 63:156:@26099.4]
  assign _T_76259 = _T_76258[10:0]; // @[Modules.scala 63:156:@26100.4]
  assign buffer_6_779 = $signed(_T_76259); // @[Modules.scala 63:156:@26101.4]
  assign _T_76261 = $signed(buffer_6_779) + $signed(buffer_6_731); // @[Modules.scala 63:156:@26103.4]
  assign _T_76262 = _T_76261[10:0]; // @[Modules.scala 63:156:@26104.4]
  assign buffer_6_780 = $signed(_T_76262); // @[Modules.scala 63:156:@26105.4]
  assign _T_76264 = $signed(buffer_6_780) + $signed(buffer_6_732); // @[Modules.scala 63:156:@26107.4]
  assign _T_76265 = _T_76264[10:0]; // @[Modules.scala 63:156:@26108.4]
  assign buffer_6_781 = $signed(_T_76265); // @[Modules.scala 63:156:@26109.4]
  assign _T_76267 = $signed(buffer_6_781) + $signed(buffer_6_733); // @[Modules.scala 63:156:@26111.4]
  assign _T_76268 = _T_76267[10:0]; // @[Modules.scala 63:156:@26112.4]
  assign buffer_6_782 = $signed(_T_76268); // @[Modules.scala 63:156:@26113.4]
  assign _T_76270 = $signed(buffer_6_782) + $signed(buffer_6_734); // @[Modules.scala 63:156:@26115.4]
  assign _T_76271 = _T_76270[10:0]; // @[Modules.scala 63:156:@26116.4]
  assign buffer_6_783 = $signed(_T_76271); // @[Modules.scala 63:156:@26117.4]
  assign _T_76273 = $signed(io_in_0) + $signed(io_in_1); // @[Modules.scala 37:46:@26120.4]
  assign _T_76274 = _T_76273[4:0]; // @[Modules.scala 37:46:@26121.4]
  assign _T_76275 = $signed(_T_76274); // @[Modules.scala 37:46:@26122.4]
  assign _T_76317 = $signed(_T_66937) + $signed(io_in_17); // @[Modules.scala 43:47:@26167.4]
  assign _T_76318 = _T_76317[4:0]; // @[Modules.scala 43:47:@26168.4]
  assign _T_76319 = $signed(_T_76318); // @[Modules.scala 43:47:@26169.4]
  assign _T_76331 = $signed(_T_69932) - $signed(io_in_21); // @[Modules.scala 46:47:@26181.4]
  assign _T_76332 = _T_76331[4:0]; // @[Modules.scala 46:47:@26182.4]
  assign _T_76333 = $signed(_T_76332); // @[Modules.scala 46:47:@26183.4]
  assign _T_76372 = $signed(_T_54372) + $signed(io_in_35); // @[Modules.scala 43:47:@26224.4]
  assign _T_76373 = _T_76372[4:0]; // @[Modules.scala 43:47:@26225.4]
  assign _T_76374 = $signed(_T_76373); // @[Modules.scala 43:47:@26226.4]
  assign _T_76410 = $signed(io_in_54) + $signed(io_in_55); // @[Modules.scala 37:46:@26270.4]
  assign _T_76411 = _T_76410[4:0]; // @[Modules.scala 37:46:@26271.4]
  assign _T_76412 = $signed(_T_76411); // @[Modules.scala 37:46:@26272.4]
  assign _T_76562 = $signed(io_in_126) - $signed(io_in_127); // @[Modules.scala 40:46:@26447.4]
  assign _T_76563 = _T_76562[4:0]; // @[Modules.scala 40:46:@26448.4]
  assign _T_76564 = $signed(_T_76563); // @[Modules.scala 40:46:@26449.4]
  assign _T_76625 = $signed(io_in_152) - $signed(io_in_153); // @[Modules.scala 40:46:@26517.4]
  assign _T_76626 = _T_76625[4:0]; // @[Modules.scala 40:46:@26518.4]
  assign _T_76627 = $signed(_T_76626); // @[Modules.scala 40:46:@26519.4]
  assign _T_76666 = $signed(_T_54746) + $signed(io_in_175); // @[Modules.scala 43:47:@26567.4]
  assign _T_76667 = _T_76666[4:0]; // @[Modules.scala 43:47:@26568.4]
  assign _T_76668 = $signed(_T_76667); // @[Modules.scala 43:47:@26569.4]
  assign _T_76680 = $signed(_T_54760) + $signed(io_in_179); // @[Modules.scala 43:47:@26581.4]
  assign _T_76681 = _T_76680[4:0]; // @[Modules.scala 43:47:@26582.4]
  assign _T_76682 = $signed(_T_76681); // @[Modules.scala 43:47:@26583.4]
  assign _T_76781 = $signed(io_in_216) + $signed(io_in_217); // @[Modules.scala 37:46:@26690.4]
  assign _T_76782 = _T_76781[4:0]; // @[Modules.scala 37:46:@26691.4]
  assign _T_76783 = $signed(_T_76782); // @[Modules.scala 37:46:@26692.4]
  assign _T_76825 = $signed(_T_54925) + $signed(io_in_233); // @[Modules.scala 43:47:@26737.4]
  assign _T_76826 = _T_76825[4:0]; // @[Modules.scala 43:47:@26738.4]
  assign _T_76827 = $signed(_T_76826); // @[Modules.scala 43:47:@26739.4]
  assign _T_76828 = $signed(io_in_234) - $signed(io_in_235); // @[Modules.scala 40:46:@26741.4]
  assign _T_76829 = _T_76828[4:0]; // @[Modules.scala 40:46:@26742.4]
  assign _T_76830 = $signed(_T_76829); // @[Modules.scala 40:46:@26743.4]
  assign _T_76945 = $signed(_T_55061) + $signed(io_in_273); // @[Modules.scala 43:47:@26862.4]
  assign _T_76946 = _T_76945[4:0]; // @[Modules.scala 43:47:@26863.4]
  assign _T_76947 = $signed(_T_76946); // @[Modules.scala 43:47:@26864.4]
  assign _T_76971 = $signed(io_in_284) + $signed(io_in_285); // @[Modules.scala 37:46:@26892.4]
  assign _T_76972 = _T_76971[4:0]; // @[Modules.scala 37:46:@26893.4]
  assign _T_76973 = $signed(_T_76972); // @[Modules.scala 37:46:@26894.4]
  assign _T_76974 = $signed(io_in_286) + $signed(io_in_287); // @[Modules.scala 37:46:@26896.4]
  assign _T_76975 = _T_76974[4:0]; // @[Modules.scala 37:46:@26897.4]
  assign _T_76976 = $signed(_T_76975); // @[Modules.scala 37:46:@26898.4]
  assign _T_76977 = $signed(io_in_288) - $signed(io_in_289); // @[Modules.scala 40:46:@26900.4]
  assign _T_76978 = _T_76977[4:0]; // @[Modules.scala 40:46:@26901.4]
  assign _T_76979 = $signed(_T_76978); // @[Modules.scala 40:46:@26902.4]
  assign _T_76983 = $signed(io_in_292) - $signed(io_in_293); // @[Modules.scala 40:46:@26908.4]
  assign _T_76984 = _T_76983[4:0]; // @[Modules.scala 40:46:@26909.4]
  assign _T_76985 = $signed(_T_76984); // @[Modules.scala 40:46:@26910.4]
  assign _T_77041 = $signed(io_in_312) + $signed(io_in_313); // @[Modules.scala 37:46:@26969.4]
  assign _T_77042 = _T_77041[4:0]; // @[Modules.scala 37:46:@26970.4]
  assign _T_77043 = $signed(_T_77042); // @[Modules.scala 37:46:@26971.4]
  assign _T_77117 = $signed(_T_64664) - $signed(io_in_337); // @[Modules.scala 46:47:@27047.4]
  assign _T_77118 = _T_77117[4:0]; // @[Modules.scala 46:47:@27048.4]
  assign _T_77119 = $signed(_T_77118); // @[Modules.scala 46:47:@27049.4]
  assign _T_77191 = $signed(io_in_364) + $signed(io_in_365); // @[Modules.scala 37:46:@27127.4]
  assign _T_77192 = _T_77191[4:0]; // @[Modules.scala 37:46:@27128.4]
  assign _T_77193 = $signed(_T_77192); // @[Modules.scala 37:46:@27129.4]
  assign _T_77234 = $signed(_T_58495) + $signed(io_in_383); // @[Modules.scala 43:47:@27175.4]
  assign _T_77235 = _T_77234[4:0]; // @[Modules.scala 43:47:@27176.4]
  assign _T_77236 = $signed(_T_77235); // @[Modules.scala 43:47:@27177.4]
  assign _T_77271 = $signed(io_in_396) - $signed(io_in_397); // @[Modules.scala 40:46:@27215.4]
  assign _T_77272 = _T_77271[4:0]; // @[Modules.scala 40:46:@27216.4]
  assign _T_77273 = $signed(_T_77272); // @[Modules.scala 40:46:@27217.4]
  assign _T_77274 = $signed(io_in_398) - $signed(io_in_399); // @[Modules.scala 40:46:@27219.4]
  assign _T_77275 = _T_77274[4:0]; // @[Modules.scala 40:46:@27220.4]
  assign _T_77276 = $signed(_T_77275); // @[Modules.scala 40:46:@27221.4]
  assign _T_77389 = $signed(_T_58658) - $signed(io_in_449); // @[Modules.scala 46:47:@27349.4]
  assign _T_77390 = _T_77389[4:0]; // @[Modules.scala 46:47:@27350.4]
  assign _T_77391 = $signed(_T_77390); // @[Modules.scala 46:47:@27351.4]
  assign _T_77396 = $signed(_T_55512) + $signed(io_in_451); // @[Modules.scala 43:47:@27356.4]
  assign _T_77397 = _T_77396[4:0]; // @[Modules.scala 43:47:@27357.4]
  assign _T_77398 = $signed(_T_77397); // @[Modules.scala 43:47:@27358.4]
  assign _T_77443 = $signed(_T_61869) + $signed(io_in_469); // @[Modules.scala 43:47:@27407.4]
  assign _T_77444 = _T_77443[4:0]; // @[Modules.scala 43:47:@27408.4]
  assign _T_77445 = $signed(_T_77444); // @[Modules.scala 43:47:@27409.4]
  assign _T_77467 = $signed(5'sh0) - $signed(io_in_478); // @[Modules.scala 46:37:@27433.4]
  assign _T_77468 = _T_77467[4:0]; // @[Modules.scala 46:37:@27434.4]
  assign _T_77469 = $signed(_T_77468); // @[Modules.scala 46:37:@27435.4]
  assign _T_77470 = $signed(_T_77469) - $signed(io_in_479); // @[Modules.scala 46:47:@27436.4]
  assign _T_77471 = _T_77470[4:0]; // @[Modules.scala 46:47:@27437.4]
  assign _T_77472 = $signed(_T_77471); // @[Modules.scala 46:47:@27438.4]
  assign _T_77473 = $signed(io_in_480) - $signed(io_in_481); // @[Modules.scala 40:46:@27440.4]
  assign _T_77474 = _T_77473[4:0]; // @[Modules.scala 40:46:@27441.4]
  assign _T_77475 = $signed(_T_77474); // @[Modules.scala 40:46:@27442.4]
  assign _T_77502 = $signed(_T_68050) - $signed(io_in_495); // @[Modules.scala 46:47:@27474.4]
  assign _T_77503 = _T_77502[4:0]; // @[Modules.scala 46:47:@27475.4]
  assign _T_77504 = $signed(_T_77503); // @[Modules.scala 46:47:@27476.4]
  assign _T_77522 = $signed(io_in_502) - $signed(io_in_503); // @[Modules.scala 40:46:@27496.4]
  assign _T_77523 = _T_77522[4:0]; // @[Modules.scala 40:46:@27497.4]
  assign _T_77524 = $signed(_T_77523); // @[Modules.scala 40:46:@27498.4]
  assign _T_77567 = $signed(io_in_524) - $signed(io_in_525); // @[Modules.scala 40:46:@27549.4]
  assign _T_77568 = _T_77567[4:0]; // @[Modules.scala 40:46:@27550.4]
  assign _T_77569 = $signed(_T_77568); // @[Modules.scala 40:46:@27551.4]
  assign _T_77574 = $signed(_T_62028) + $signed(io_in_527); // @[Modules.scala 43:47:@27556.4]
  assign _T_77575 = _T_77574[4:0]; // @[Modules.scala 43:47:@27557.4]
  assign _T_77576 = $signed(_T_77575); // @[Modules.scala 43:47:@27558.4]
  assign _T_77604 = $signed(io_in_538) - $signed(io_in_539); // @[Modules.scala 40:46:@27589.4]
  assign _T_77605 = _T_77604[4:0]; // @[Modules.scala 40:46:@27590.4]
  assign _T_77606 = $signed(_T_77605); // @[Modules.scala 40:46:@27591.4]
  assign _T_77629 = $signed(_T_74419) + $signed(io_in_553); // @[Modules.scala 43:47:@27620.4]
  assign _T_77630 = _T_77629[4:0]; // @[Modules.scala 43:47:@27621.4]
  assign _T_77631 = $signed(_T_77630); // @[Modules.scala 43:47:@27622.4]
  assign _T_77692 = $signed(io_in_586) - $signed(io_in_587); // @[Modules.scala 40:46:@27697.4]
  assign _T_77693 = _T_77692[4:0]; // @[Modules.scala 40:46:@27698.4]
  assign _T_77694 = $signed(_T_77693); // @[Modules.scala 40:46:@27699.4]
  assign _T_77730 = $signed(_T_55910) + $signed(io_in_599); // @[Modules.scala 43:47:@27736.4]
  assign _T_77731 = _T_77730[4:0]; // @[Modules.scala 43:47:@27737.4]
  assign _T_77732 = $signed(_T_77731); // @[Modules.scala 43:47:@27738.4]
  assign _T_77744 = $signed(_T_65323) + $signed(io_in_603); // @[Modules.scala 43:47:@27750.4]
  assign _T_77745 = _T_77744[4:0]; // @[Modules.scala 43:47:@27751.4]
  assign _T_77746 = $signed(_T_77745); // @[Modules.scala 43:47:@27752.4]
  assign _T_77774 = $signed(_T_55946) - $signed(io_in_615); // @[Modules.scala 46:47:@27783.4]
  assign _T_77775 = _T_77774[4:0]; // @[Modules.scala 46:47:@27784.4]
  assign _T_77776 = $signed(_T_77775); // @[Modules.scala 46:47:@27785.4]
  assign _T_77794 = $signed(io_in_622) - $signed(io_in_623); // @[Modules.scala 40:46:@27805.4]
  assign _T_77795 = _T_77794[4:0]; // @[Modules.scala 40:46:@27806.4]
  assign _T_77796 = $signed(_T_77795); // @[Modules.scala 40:46:@27807.4]
  assign _T_77960 = $signed(_T_65519) + $signed(io_in_691); // @[Modules.scala 43:47:@27989.4]
  assign _T_77961 = _T_77960[4:0]; // @[Modules.scala 43:47:@27990.4]
  assign _T_77962 = $signed(_T_77961); // @[Modules.scala 43:47:@27991.4]
  assign _T_78189 = $signed(_T_71722) + $signed(io_in_761); // @[Modules.scala 43:47:@28222.4]
  assign _T_78190 = _T_78189[4:0]; // @[Modules.scala 43:47:@28223.4]
  assign _T_78191 = $signed(_T_78190); // @[Modules.scala 43:47:@28224.4]
  assign _T_78255 = $signed(io_in_780) + $signed(io_in_781); // @[Modules.scala 37:46:@28289.4]
  assign _T_78256 = _T_78255[4:0]; // @[Modules.scala 37:46:@28290.4]
  assign _T_78257 = $signed(_T_78256); // @[Modules.scala 37:46:@28291.4]
  assign buffer_7_0 = {{6{_T_76275[4]}},_T_76275}; // @[Modules.scala 32:22:@8.4]
  assign _T_78265 = $signed(buffer_7_0) + $signed(buffer_0_1); // @[Modules.scala 50:57:@28300.4]
  assign _T_78266 = _T_78265[10:0]; // @[Modules.scala 50:57:@28301.4]
  assign buffer_7_392 = $signed(_T_78266); // @[Modules.scala 50:57:@28302.4]
  assign _T_78268 = $signed(buffer_2_2) + $signed(buffer_0_3); // @[Modules.scala 50:57:@28304.4]
  assign _T_78269 = _T_78268[10:0]; // @[Modules.scala 50:57:@28305.4]
  assign buffer_7_393 = $signed(_T_78269); // @[Modules.scala 50:57:@28306.4]
  assign buffer_7_8 = {{6{_T_76319[4]}},_T_76319}; // @[Modules.scala 32:22:@8.4]
  assign _T_78277 = $signed(buffer_7_8) + $signed(buffer_2_9); // @[Modules.scala 50:57:@28316.4]
  assign _T_78278 = _T_78277[10:0]; // @[Modules.scala 50:57:@28317.4]
  assign buffer_7_396 = $signed(_T_78278); // @[Modules.scala 50:57:@28318.4]
  assign buffer_7_10 = {{6{_T_76333[4]}},_T_76333}; // @[Modules.scala 32:22:@8.4]
  assign _T_78280 = $signed(buffer_7_10) + $signed(buffer_0_11); // @[Modules.scala 50:57:@28320.4]
  assign _T_78281 = _T_78280[10:0]; // @[Modules.scala 50:57:@28321.4]
  assign buffer_7_397 = $signed(_T_78281); // @[Modules.scala 50:57:@28322.4]
  assign _T_78286 = $signed(buffer_1_14) + $signed(buffer_3_15); // @[Modules.scala 50:57:@28328.4]
  assign _T_78287 = _T_78286[10:0]; // @[Modules.scala 50:57:@28329.4]
  assign buffer_7_399 = $signed(_T_78287); // @[Modules.scala 50:57:@28330.4]
  assign buffer_7_17 = {{6{_T_76374[4]}},_T_76374}; // @[Modules.scala 32:22:@8.4]
  assign _T_78289 = $signed(buffer_5_16) + $signed(buffer_7_17); // @[Modules.scala 50:57:@28332.4]
  assign _T_78290 = _T_78289[10:0]; // @[Modules.scala 50:57:@28333.4]
  assign buffer_7_400 = $signed(_T_78290); // @[Modules.scala 50:57:@28334.4]
  assign buffer_7_27 = {{6{_T_76412[4]}},_T_76412}; // @[Modules.scala 32:22:@8.4]
  assign _T_78304 = $signed(buffer_3_26) + $signed(buffer_7_27); // @[Modules.scala 50:57:@28352.4]
  assign _T_78305 = _T_78304[10:0]; // @[Modules.scala 50:57:@28353.4]
  assign buffer_7_405 = $signed(_T_78305); // @[Modules.scala 50:57:@28354.4]
  assign _T_78310 = $signed(buffer_3_30) + $signed(buffer_1_31); // @[Modules.scala 50:57:@28360.4]
  assign _T_78311 = _T_78310[10:0]; // @[Modules.scala 50:57:@28361.4]
  assign buffer_7_407 = $signed(_T_78311); // @[Modules.scala 50:57:@28362.4]
  assign _T_78337 = $signed(buffer_2_48) + $signed(buffer_0_49); // @[Modules.scala 50:57:@28396.4]
  assign _T_78338 = _T_78337[10:0]; // @[Modules.scala 50:57:@28397.4]
  assign buffer_7_416 = $signed(_T_78338); // @[Modules.scala 50:57:@28398.4]
  assign _T_78352 = $signed(buffer_4_58) + $signed(buffer_0_59); // @[Modules.scala 50:57:@28416.4]
  assign _T_78353 = _T_78352[10:0]; // @[Modules.scala 50:57:@28417.4]
  assign buffer_7_421 = $signed(_T_78353); // @[Modules.scala 50:57:@28418.4]
  assign _T_78355 = $signed(buffer_3_60) + $signed(buffer_0_61); // @[Modules.scala 50:57:@28420.4]
  assign _T_78356 = _T_78355[10:0]; // @[Modules.scala 50:57:@28421.4]
  assign buffer_7_422 = $signed(_T_78356); // @[Modules.scala 50:57:@28422.4]
  assign buffer_7_63 = {{6{_T_76564[4]}},_T_76564}; // @[Modules.scala 32:22:@8.4]
  assign _T_78358 = $signed(buffer_0_62) + $signed(buffer_7_63); // @[Modules.scala 50:57:@28424.4]
  assign _T_78359 = _T_78358[10:0]; // @[Modules.scala 50:57:@28425.4]
  assign buffer_7_423 = $signed(_T_78359); // @[Modules.scala 50:57:@28426.4]
  assign _T_78364 = $signed(buffer_3_66) + $signed(buffer_0_67); // @[Modules.scala 50:57:@28432.4]
  assign _T_78365 = _T_78364[10:0]; // @[Modules.scala 50:57:@28433.4]
  assign buffer_7_425 = $signed(_T_78365); // @[Modules.scala 50:57:@28434.4]
  assign _T_78373 = $signed(buffer_1_72) + $signed(buffer_5_73); // @[Modules.scala 50:57:@28444.4]
  assign _T_78374 = _T_78373[10:0]; // @[Modules.scala 50:57:@28445.4]
  assign buffer_7_428 = $signed(_T_78374); // @[Modules.scala 50:57:@28446.4]
  assign _T_78376 = $signed(buffer_6_74) + $signed(buffer_1_75); // @[Modules.scala 50:57:@28448.4]
  assign _T_78377 = _T_78376[10:0]; // @[Modules.scala 50:57:@28449.4]
  assign buffer_7_429 = $signed(_T_78377); // @[Modules.scala 50:57:@28450.4]
  assign buffer_7_76 = {{6{_T_76627[4]}},_T_76627}; // @[Modules.scala 32:22:@8.4]
  assign _T_78379 = $signed(buffer_7_76) + $signed(buffer_3_77); // @[Modules.scala 50:57:@28452.4]
  assign _T_78380 = _T_78379[10:0]; // @[Modules.scala 50:57:@28453.4]
  assign buffer_7_430 = $signed(_T_78380); // @[Modules.scala 50:57:@28454.4]
  assign buffer_7_87 = {{6{_T_76668[4]}},_T_76668}; // @[Modules.scala 32:22:@8.4]
  assign _T_78394 = $signed(buffer_3_86) + $signed(buffer_7_87); // @[Modules.scala 50:57:@28472.4]
  assign _T_78395 = _T_78394[10:0]; // @[Modules.scala 50:57:@28473.4]
  assign buffer_7_435 = $signed(_T_78395); // @[Modules.scala 50:57:@28474.4]
  assign buffer_7_89 = {{6{_T_76682[4]}},_T_76682}; // @[Modules.scala 32:22:@8.4]
  assign _T_78397 = $signed(buffer_0_88) + $signed(buffer_7_89); // @[Modules.scala 50:57:@28476.4]
  assign _T_78398 = _T_78397[10:0]; // @[Modules.scala 50:57:@28477.4]
  assign buffer_7_436 = $signed(_T_78398); // @[Modules.scala 50:57:@28478.4]
  assign _T_78406 = $signed(buffer_6_94) + $signed(buffer_2_95); // @[Modules.scala 50:57:@28488.4]
  assign _T_78407 = _T_78406[10:0]; // @[Modules.scala 50:57:@28489.4]
  assign buffer_7_439 = $signed(_T_78407); // @[Modules.scala 50:57:@28490.4]
  assign buffer_7_108 = {{6{_T_76783[4]}},_T_76783}; // @[Modules.scala 32:22:@8.4]
  assign _T_78427 = $signed(buffer_7_108) + $signed(buffer_2_109); // @[Modules.scala 50:57:@28516.4]
  assign _T_78428 = _T_78427[10:0]; // @[Modules.scala 50:57:@28517.4]
  assign buffer_7_446 = $signed(_T_78428); // @[Modules.scala 50:57:@28518.4]
  assign _T_78436 = $signed(buffer_0_114) + $signed(buffer_3_115); // @[Modules.scala 50:57:@28528.4]
  assign _T_78437 = _T_78436[10:0]; // @[Modules.scala 50:57:@28529.4]
  assign buffer_7_449 = $signed(_T_78437); // @[Modules.scala 50:57:@28530.4]
  assign buffer_7_116 = {{6{_T_76827[4]}},_T_76827}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_117 = {{6{_T_76830[4]}},_T_76830}; // @[Modules.scala 32:22:@8.4]
  assign _T_78439 = $signed(buffer_7_116) + $signed(buffer_7_117); // @[Modules.scala 50:57:@28532.4]
  assign _T_78440 = _T_78439[10:0]; // @[Modules.scala 50:57:@28533.4]
  assign buffer_7_450 = $signed(_T_78440); // @[Modules.scala 50:57:@28534.4]
  assign _T_78448 = $signed(buffer_3_122) + $signed(buffer_1_123); // @[Modules.scala 50:57:@28544.4]
  assign _T_78449 = _T_78448[10:0]; // @[Modules.scala 50:57:@28545.4]
  assign buffer_7_453 = $signed(_T_78449); // @[Modules.scala 50:57:@28546.4]
  assign _T_78466 = $signed(buffer_0_134) + $signed(buffer_5_135); // @[Modules.scala 50:57:@28568.4]
  assign _T_78467 = _T_78466[10:0]; // @[Modules.scala 50:57:@28569.4]
  assign buffer_7_459 = $signed(_T_78467); // @[Modules.scala 50:57:@28570.4]
  assign buffer_7_136 = {{6{_T_76947[4]}},_T_76947}; // @[Modules.scala 32:22:@8.4]
  assign _T_78469 = $signed(buffer_7_136) + $signed(buffer_3_137); // @[Modules.scala 50:57:@28572.4]
  assign _T_78470 = _T_78469[10:0]; // @[Modules.scala 50:57:@28573.4]
  assign buffer_7_460 = $signed(_T_78470); // @[Modules.scala 50:57:@28574.4]
  assign buffer_7_142 = {{6{_T_76973[4]}},_T_76973}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_143 = {{6{_T_76976[4]}},_T_76976}; // @[Modules.scala 32:22:@8.4]
  assign _T_78478 = $signed(buffer_7_142) + $signed(buffer_7_143); // @[Modules.scala 50:57:@28584.4]
  assign _T_78479 = _T_78478[10:0]; // @[Modules.scala 50:57:@28585.4]
  assign buffer_7_463 = $signed(_T_78479); // @[Modules.scala 50:57:@28586.4]
  assign buffer_7_144 = {{6{_T_76979[4]}},_T_76979}; // @[Modules.scala 32:22:@8.4]
  assign _T_78481 = $signed(buffer_7_144) + $signed(buffer_6_145); // @[Modules.scala 50:57:@28588.4]
  assign _T_78482 = _T_78481[10:0]; // @[Modules.scala 50:57:@28589.4]
  assign buffer_7_464 = $signed(_T_78482); // @[Modules.scala 50:57:@28590.4]
  assign buffer_7_146 = {{6{_T_76985[4]}},_T_76985}; // @[Modules.scala 32:22:@8.4]
  assign _T_78484 = $signed(buffer_7_146) + $signed(buffer_0_147); // @[Modules.scala 50:57:@28592.4]
  assign _T_78485 = _T_78484[10:0]; // @[Modules.scala 50:57:@28593.4]
  assign buffer_7_465 = $signed(_T_78485); // @[Modules.scala 50:57:@28594.4]
  assign buffer_7_156 = {{6{_T_77043[4]}},_T_77043}; // @[Modules.scala 32:22:@8.4]
  assign _T_78499 = $signed(buffer_7_156) + $signed(buffer_0_157); // @[Modules.scala 50:57:@28612.4]
  assign _T_78500 = _T_78499[10:0]; // @[Modules.scala 50:57:@28613.4]
  assign buffer_7_470 = $signed(_T_78500); // @[Modules.scala 50:57:@28614.4]
  assign _T_78502 = $signed(buffer_6_158) + $signed(buffer_3_159); // @[Modules.scala 50:57:@28616.4]
  assign _T_78503 = _T_78502[10:0]; // @[Modules.scala 50:57:@28617.4]
  assign buffer_7_471 = $signed(_T_78503); // @[Modules.scala 50:57:@28618.4]
  assign buffer_7_168 = {{6{_T_77119[4]}},_T_77119}; // @[Modules.scala 32:22:@8.4]
  assign _T_78517 = $signed(buffer_7_168) + $signed(buffer_0_169); // @[Modules.scala 50:57:@28636.4]
  assign _T_78518 = _T_78517[10:0]; // @[Modules.scala 50:57:@28637.4]
  assign buffer_7_476 = $signed(_T_78518); // @[Modules.scala 50:57:@28638.4]
  assign _T_78532 = $signed(buffer_6_178) + $signed(buffer_2_179); // @[Modules.scala 50:57:@28656.4]
  assign _T_78533 = _T_78532[10:0]; // @[Modules.scala 50:57:@28657.4]
  assign buffer_7_481 = $signed(_T_78533); // @[Modules.scala 50:57:@28658.4]
  assign buffer_7_182 = {{6{_T_77193[4]}},_T_77193}; // @[Modules.scala 32:22:@8.4]
  assign _T_78538 = $signed(buffer_7_182) + $signed(buffer_5_183); // @[Modules.scala 50:57:@28664.4]
  assign _T_78539 = _T_78538[10:0]; // @[Modules.scala 50:57:@28665.4]
  assign buffer_7_483 = $signed(_T_78539); // @[Modules.scala 50:57:@28666.4]
  assign buffer_7_191 = {{6{_T_77236[4]}},_T_77236}; // @[Modules.scala 32:22:@8.4]
  assign _T_78550 = $signed(buffer_1_190) + $signed(buffer_7_191); // @[Modules.scala 50:57:@28680.4]
  assign _T_78551 = _T_78550[10:0]; // @[Modules.scala 50:57:@28681.4]
  assign buffer_7_487 = $signed(_T_78551); // @[Modules.scala 50:57:@28682.4]
  assign _T_78559 = $signed(buffer_4_196) + $signed(buffer_5_197); // @[Modules.scala 50:57:@28692.4]
  assign _T_78560 = _T_78559[10:0]; // @[Modules.scala 50:57:@28693.4]
  assign buffer_7_490 = $signed(_T_78560); // @[Modules.scala 50:57:@28694.4]
  assign buffer_7_198 = {{6{_T_77273[4]}},_T_77273}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_199 = {{6{_T_77276[4]}},_T_77276}; // @[Modules.scala 32:22:@8.4]
  assign _T_78562 = $signed(buffer_7_198) + $signed(buffer_7_199); // @[Modules.scala 50:57:@28696.4]
  assign _T_78563 = _T_78562[10:0]; // @[Modules.scala 50:57:@28697.4]
  assign buffer_7_491 = $signed(_T_78563); // @[Modules.scala 50:57:@28698.4]
  assign _T_78565 = $signed(buffer_5_200) + $signed(buffer_0_201); // @[Modules.scala 50:57:@28700.4]
  assign _T_78566 = _T_78565[10:0]; // @[Modules.scala 50:57:@28701.4]
  assign buffer_7_492 = $signed(_T_78566); // @[Modules.scala 50:57:@28702.4]
  assign _T_78571 = $signed(buffer_1_204) + $signed(buffer_3_205); // @[Modules.scala 50:57:@28708.4]
  assign _T_78572 = _T_78571[10:0]; // @[Modules.scala 50:57:@28709.4]
  assign buffer_7_494 = $signed(_T_78572); // @[Modules.scala 50:57:@28710.4]
  assign _T_78580 = $signed(buffer_3_210) + $signed(buffer_5_211); // @[Modules.scala 50:57:@28720.4]
  assign _T_78581 = _T_78580[10:0]; // @[Modules.scala 50:57:@28721.4]
  assign buffer_7_497 = $signed(_T_78581); // @[Modules.scala 50:57:@28722.4]
  assign _T_78583 = $signed(buffer_3_212) + $signed(buffer_0_213); // @[Modules.scala 50:57:@28724.4]
  assign _T_78584 = _T_78583[10:0]; // @[Modules.scala 50:57:@28725.4]
  assign buffer_7_498 = $signed(_T_78584); // @[Modules.scala 50:57:@28726.4]
  assign _T_78586 = $signed(buffer_0_214) + $signed(buffer_6_215); // @[Modules.scala 50:57:@28728.4]
  assign _T_78587 = _T_78586[10:0]; // @[Modules.scala 50:57:@28729.4]
  assign buffer_7_499 = $signed(_T_78587); // @[Modules.scala 50:57:@28730.4]
  assign _T_78592 = $signed(buffer_4_218) + $signed(buffer_0_219); // @[Modules.scala 50:57:@28736.4]
  assign _T_78593 = _T_78592[10:0]; // @[Modules.scala 50:57:@28737.4]
  assign buffer_7_501 = $signed(_T_78593); // @[Modules.scala 50:57:@28738.4]
  assign buffer_7_224 = {{6{_T_77391[4]}},_T_77391}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_225 = {{6{_T_77398[4]}},_T_77398}; // @[Modules.scala 32:22:@8.4]
  assign _T_78601 = $signed(buffer_7_224) + $signed(buffer_7_225); // @[Modules.scala 50:57:@28748.4]
  assign _T_78602 = _T_78601[10:0]; // @[Modules.scala 50:57:@28749.4]
  assign buffer_7_504 = $signed(_T_78602); // @[Modules.scala 50:57:@28750.4]
  assign _T_78607 = $signed(buffer_3_228) + $signed(buffer_0_229); // @[Modules.scala 50:57:@28756.4]
  assign _T_78608 = _T_78607[10:0]; // @[Modules.scala 50:57:@28757.4]
  assign buffer_7_506 = $signed(_T_78608); // @[Modules.scala 50:57:@28758.4]
  assign buffer_7_234 = {{6{_T_77445[4]}},_T_77445}; // @[Modules.scala 32:22:@8.4]
  assign _T_78616 = $signed(buffer_7_234) + $signed(buffer_0_235); // @[Modules.scala 50:57:@28768.4]
  assign _T_78617 = _T_78616[10:0]; // @[Modules.scala 50:57:@28769.4]
  assign buffer_7_509 = $signed(_T_78617); // @[Modules.scala 50:57:@28770.4]
  assign buffer_7_239 = {{6{_T_77472[4]}},_T_77472}; // @[Modules.scala 32:22:@8.4]
  assign _T_78622 = $signed(buffer_0_238) + $signed(buffer_7_239); // @[Modules.scala 50:57:@28776.4]
  assign _T_78623 = _T_78622[10:0]; // @[Modules.scala 50:57:@28777.4]
  assign buffer_7_511 = $signed(_T_78623); // @[Modules.scala 50:57:@28778.4]
  assign buffer_7_240 = {{6{_T_77475[4]}},_T_77475}; // @[Modules.scala 32:22:@8.4]
  assign _T_78625 = $signed(buffer_7_240) + $signed(buffer_0_241); // @[Modules.scala 50:57:@28780.4]
  assign _T_78626 = _T_78625[10:0]; // @[Modules.scala 50:57:@28781.4]
  assign buffer_7_512 = $signed(_T_78626); // @[Modules.scala 50:57:@28782.4]
  assign buffer_7_247 = {{6{_T_77504[4]}},_T_77504}; // @[Modules.scala 32:22:@8.4]
  assign _T_78634 = $signed(buffer_0_246) + $signed(buffer_7_247); // @[Modules.scala 50:57:@28792.4]
  assign _T_78635 = _T_78634[10:0]; // @[Modules.scala 50:57:@28793.4]
  assign buffer_7_515 = $signed(_T_78635); // @[Modules.scala 50:57:@28794.4]
  assign buffer_7_251 = {{6{_T_77524[4]}},_T_77524}; // @[Modules.scala 32:22:@8.4]
  assign _T_78640 = $signed(buffer_3_250) + $signed(buffer_7_251); // @[Modules.scala 50:57:@28800.4]
  assign _T_78641 = _T_78640[10:0]; // @[Modules.scala 50:57:@28801.4]
  assign buffer_7_517 = $signed(_T_78641); // @[Modules.scala 50:57:@28802.4]
  assign _T_78655 = $signed(buffer_2_260) + $signed(buffer_1_261); // @[Modules.scala 50:57:@28820.4]
  assign _T_78656 = _T_78655[10:0]; // @[Modules.scala 50:57:@28821.4]
  assign buffer_7_522 = $signed(_T_78656); // @[Modules.scala 50:57:@28822.4]
  assign buffer_7_262 = {{6{_T_77569[4]}},_T_77569}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_263 = {{6{_T_77576[4]}},_T_77576}; // @[Modules.scala 32:22:@8.4]
  assign _T_78658 = $signed(buffer_7_262) + $signed(buffer_7_263); // @[Modules.scala 50:57:@28824.4]
  assign _T_78659 = _T_78658[10:0]; // @[Modules.scala 50:57:@28825.4]
  assign buffer_7_523 = $signed(_T_78659); // @[Modules.scala 50:57:@28826.4]
  assign buffer_7_269 = {{6{_T_77606[4]}},_T_77606}; // @[Modules.scala 32:22:@8.4]
  assign _T_78667 = $signed(buffer_0_268) + $signed(buffer_7_269); // @[Modules.scala 50:57:@28836.4]
  assign _T_78668 = _T_78667[10:0]; // @[Modules.scala 50:57:@28837.4]
  assign buffer_7_526 = $signed(_T_78668); // @[Modules.scala 50:57:@28838.4]
  assign _T_78673 = $signed(buffer_1_272) + $signed(buffer_4_273); // @[Modules.scala 50:57:@28844.4]
  assign _T_78674 = _T_78673[10:0]; // @[Modules.scala 50:57:@28845.4]
  assign buffer_7_528 = $signed(_T_78674); // @[Modules.scala 50:57:@28846.4]
  assign _T_78676 = $signed(buffer_1_274) + $signed(buffer_0_275); // @[Modules.scala 50:57:@28848.4]
  assign _T_78677 = _T_78676[10:0]; // @[Modules.scala 50:57:@28849.4]
  assign buffer_7_529 = $signed(_T_78677); // @[Modules.scala 50:57:@28850.4]
  assign buffer_7_276 = {{6{_T_77631[4]}},_T_77631}; // @[Modules.scala 32:22:@8.4]
  assign _T_78679 = $signed(buffer_7_276) + $signed(buffer_3_277); // @[Modules.scala 50:57:@28852.4]
  assign _T_78680 = _T_78679[10:0]; // @[Modules.scala 50:57:@28853.4]
  assign buffer_7_530 = $signed(_T_78680); // @[Modules.scala 50:57:@28854.4]
  assign _T_78688 = $signed(buffer_0_282) + $signed(buffer_3_283); // @[Modules.scala 50:57:@28864.4]
  assign _T_78689 = _T_78688[10:0]; // @[Modules.scala 50:57:@28865.4]
  assign buffer_7_533 = $signed(_T_78689); // @[Modules.scala 50:57:@28866.4]
  assign buffer_7_293 = {{6{_T_77694[4]}},_T_77694}; // @[Modules.scala 32:22:@8.4]
  assign _T_78703 = $signed(buffer_4_292) + $signed(buffer_7_293); // @[Modules.scala 50:57:@28884.4]
  assign _T_78704 = _T_78703[10:0]; // @[Modules.scala 50:57:@28885.4]
  assign buffer_7_538 = $signed(_T_78704); // @[Modules.scala 50:57:@28886.4]
  assign _T_78706 = $signed(buffer_1_294) + $signed(buffer_0_295); // @[Modules.scala 50:57:@28888.4]
  assign _T_78707 = _T_78706[10:0]; // @[Modules.scala 50:57:@28889.4]
  assign buffer_7_539 = $signed(_T_78707); // @[Modules.scala 50:57:@28890.4]
  assign buffer_7_299 = {{6{_T_77732[4]}},_T_77732}; // @[Modules.scala 32:22:@8.4]
  assign _T_78712 = $signed(buffer_2_298) + $signed(buffer_7_299); // @[Modules.scala 50:57:@28896.4]
  assign _T_78713 = _T_78712[10:0]; // @[Modules.scala 50:57:@28897.4]
  assign buffer_7_541 = $signed(_T_78713); // @[Modules.scala 50:57:@28898.4]
  assign buffer_7_301 = {{6{_T_77746[4]}},_T_77746}; // @[Modules.scala 32:22:@8.4]
  assign _T_78715 = $signed(buffer_2_300) + $signed(buffer_7_301); // @[Modules.scala 50:57:@28900.4]
  assign _T_78716 = _T_78715[10:0]; // @[Modules.scala 50:57:@28901.4]
  assign buffer_7_542 = $signed(_T_78716); // @[Modules.scala 50:57:@28902.4]
  assign buffer_7_307 = {{6{_T_77776[4]}},_T_77776}; // @[Modules.scala 32:22:@8.4]
  assign _T_78724 = $signed(buffer_4_306) + $signed(buffer_7_307); // @[Modules.scala 50:57:@28912.4]
  assign _T_78725 = _T_78724[10:0]; // @[Modules.scala 50:57:@28913.4]
  assign buffer_7_545 = $signed(_T_78725); // @[Modules.scala 50:57:@28914.4]
  assign _T_78727 = $signed(buffer_1_308) + $signed(buffer_2_309); // @[Modules.scala 50:57:@28916.4]
  assign _T_78728 = _T_78727[10:0]; // @[Modules.scala 50:57:@28917.4]
  assign buffer_7_546 = $signed(_T_78728); // @[Modules.scala 50:57:@28918.4]
  assign buffer_7_311 = {{6{_T_77796[4]}},_T_77796}; // @[Modules.scala 32:22:@8.4]
  assign _T_78730 = $signed(buffer_3_310) + $signed(buffer_7_311); // @[Modules.scala 50:57:@28920.4]
  assign _T_78731 = _T_78730[10:0]; // @[Modules.scala 50:57:@28921.4]
  assign buffer_7_547 = $signed(_T_78731); // @[Modules.scala 50:57:@28922.4]
  assign _T_78733 = $signed(buffer_6_312) + $signed(buffer_3_313); // @[Modules.scala 50:57:@28924.4]
  assign _T_78734 = _T_78733[10:0]; // @[Modules.scala 50:57:@28925.4]
  assign buffer_7_548 = $signed(_T_78734); // @[Modules.scala 50:57:@28926.4]
  assign _T_78739 = $signed(buffer_0_316) + $signed(buffer_2_317); // @[Modules.scala 50:57:@28932.4]
  assign _T_78740 = _T_78739[10:0]; // @[Modules.scala 50:57:@28933.4]
  assign buffer_7_550 = $signed(_T_78740); // @[Modules.scala 50:57:@28934.4]
  assign _T_78748 = $signed(buffer_2_322) + $signed(buffer_6_323); // @[Modules.scala 50:57:@28944.4]
  assign _T_78749 = _T_78748[10:0]; // @[Modules.scala 50:57:@28945.4]
  assign buffer_7_553 = $signed(_T_78749); // @[Modules.scala 50:57:@28946.4]
  assign _T_78757 = $signed(buffer_0_328) + $signed(buffer_5_329); // @[Modules.scala 50:57:@28956.4]
  assign _T_78758 = _T_78757[10:0]; // @[Modules.scala 50:57:@28957.4]
  assign buffer_7_556 = $signed(_T_78758); // @[Modules.scala 50:57:@28958.4]
  assign _T_78763 = $signed(buffer_0_332) + $signed(buffer_3_333); // @[Modules.scala 50:57:@28964.4]
  assign _T_78764 = _T_78763[10:0]; // @[Modules.scala 50:57:@28965.4]
  assign buffer_7_558 = $signed(_T_78764); // @[Modules.scala 50:57:@28966.4]
  assign _T_78766 = $signed(buffer_0_334) + $signed(buffer_2_335); // @[Modules.scala 50:57:@28968.4]
  assign _T_78767 = _T_78766[10:0]; // @[Modules.scala 50:57:@28969.4]
  assign buffer_7_559 = $signed(_T_78767); // @[Modules.scala 50:57:@28970.4]
  assign _T_78769 = $signed(buffer_4_336) + $signed(buffer_0_337); // @[Modules.scala 50:57:@28972.4]
  assign _T_78770 = _T_78769[10:0]; // @[Modules.scala 50:57:@28973.4]
  assign buffer_7_560 = $signed(_T_78770); // @[Modules.scala 50:57:@28974.4]
  assign _T_78778 = $signed(buffer_2_342) + $signed(buffer_3_343); // @[Modules.scala 50:57:@28984.4]
  assign _T_78779 = _T_78778[10:0]; // @[Modules.scala 50:57:@28985.4]
  assign buffer_7_563 = $signed(_T_78779); // @[Modules.scala 50:57:@28986.4]
  assign buffer_7_345 = {{6{_T_77962[4]}},_T_77962}; // @[Modules.scala 32:22:@8.4]
  assign _T_78781 = $signed(buffer_3_344) + $signed(buffer_7_345); // @[Modules.scala 50:57:@28988.4]
  assign _T_78782 = _T_78781[10:0]; // @[Modules.scala 50:57:@28989.4]
  assign buffer_7_564 = $signed(_T_78782); // @[Modules.scala 50:57:@28990.4]
  assign _T_78787 = $signed(buffer_4_348) + $signed(buffer_1_349); // @[Modules.scala 50:57:@28996.4]
  assign _T_78788 = _T_78787[10:0]; // @[Modules.scala 50:57:@28997.4]
  assign buffer_7_566 = $signed(_T_78788); // @[Modules.scala 50:57:@28998.4]
  assign _T_78790 = $signed(buffer_2_350) + $signed(buffer_5_351); // @[Modules.scala 50:57:@29000.4]
  assign _T_78791 = _T_78790[10:0]; // @[Modules.scala 50:57:@29001.4]
  assign buffer_7_567 = $signed(_T_78791); // @[Modules.scala 50:57:@29002.4]
  assign _T_78808 = $signed(buffer_4_362) + $signed(buffer_1_363); // @[Modules.scala 50:57:@29024.4]
  assign _T_78809 = _T_78808[10:0]; // @[Modules.scala 50:57:@29025.4]
  assign buffer_7_573 = $signed(_T_78809); // @[Modules.scala 50:57:@29026.4]
  assign _T_78829 = $signed(buffer_4_376) + $signed(buffer_0_377); // @[Modules.scala 50:57:@29052.4]
  assign _T_78830 = _T_78829[10:0]; // @[Modules.scala 50:57:@29053.4]
  assign buffer_7_580 = $signed(_T_78830); // @[Modules.scala 50:57:@29054.4]
  assign buffer_7_380 = {{6{_T_78191[4]}},_T_78191}; // @[Modules.scala 32:22:@8.4]
  assign _T_78835 = $signed(buffer_7_380) + $signed(buffer_0_381); // @[Modules.scala 50:57:@29060.4]
  assign _T_78836 = _T_78835[10:0]; // @[Modules.scala 50:57:@29061.4]
  assign buffer_7_582 = $signed(_T_78836); // @[Modules.scala 50:57:@29062.4]
  assign buffer_7_390 = {{6{_T_78257[4]}},_T_78257}; // @[Modules.scala 32:22:@8.4]
  assign _T_78850 = $signed(buffer_7_390) + $signed(buffer_2_391); // @[Modules.scala 50:57:@29080.4]
  assign _T_78851 = _T_78850[10:0]; // @[Modules.scala 50:57:@29081.4]
  assign buffer_7_587 = $signed(_T_78851); // @[Modules.scala 50:57:@29082.4]
  assign _T_78853 = $signed(buffer_7_392) + $signed(buffer_7_393); // @[Modules.scala 53:83:@29084.4]
  assign _T_78854 = _T_78853[10:0]; // @[Modules.scala 53:83:@29085.4]
  assign buffer_7_588 = $signed(_T_78854); // @[Modules.scala 53:83:@29086.4]
  assign _T_78859 = $signed(buffer_7_396) + $signed(buffer_7_397); // @[Modules.scala 53:83:@29092.4]
  assign _T_78860 = _T_78859[10:0]; // @[Modules.scala 53:83:@29093.4]
  assign buffer_7_590 = $signed(_T_78860); // @[Modules.scala 53:83:@29094.4]
  assign _T_78862 = $signed(buffer_2_398) + $signed(buffer_7_399); // @[Modules.scala 53:83:@29096.4]
  assign _T_78863 = _T_78862[10:0]; // @[Modules.scala 53:83:@29097.4]
  assign buffer_7_591 = $signed(_T_78863); // @[Modules.scala 53:83:@29098.4]
  assign _T_78865 = $signed(buffer_7_400) + $signed(buffer_1_401); // @[Modules.scala 53:83:@29100.4]
  assign _T_78866 = _T_78865[10:0]; // @[Modules.scala 53:83:@29101.4]
  assign buffer_7_592 = $signed(_T_78866); // @[Modules.scala 53:83:@29102.4]
  assign _T_78868 = $signed(buffer_2_402) + $signed(buffer_4_403); // @[Modules.scala 53:83:@29104.4]
  assign _T_78869 = _T_78868[10:0]; // @[Modules.scala 53:83:@29105.4]
  assign buffer_7_593 = $signed(_T_78869); // @[Modules.scala 53:83:@29106.4]
  assign _T_78871 = $signed(buffer_1_404) + $signed(buffer_7_405); // @[Modules.scala 53:83:@29108.4]
  assign _T_78872 = _T_78871[10:0]; // @[Modules.scala 53:83:@29109.4]
  assign buffer_7_594 = $signed(_T_78872); // @[Modules.scala 53:83:@29110.4]
  assign _T_78874 = $signed(buffer_0_406) + $signed(buffer_7_407); // @[Modules.scala 53:83:@29112.4]
  assign _T_78875 = _T_78874[10:0]; // @[Modules.scala 53:83:@29113.4]
  assign buffer_7_595 = $signed(_T_78875); // @[Modules.scala 53:83:@29114.4]
  assign _T_78883 = $signed(buffer_3_412) + $signed(buffer_1_413); // @[Modules.scala 53:83:@29124.4]
  assign _T_78884 = _T_78883[10:0]; // @[Modules.scala 53:83:@29125.4]
  assign buffer_7_598 = $signed(_T_78884); // @[Modules.scala 53:83:@29126.4]
  assign _T_78886 = $signed(buffer_2_414) + $signed(buffer_1_415); // @[Modules.scala 53:83:@29128.4]
  assign _T_78887 = _T_78886[10:0]; // @[Modules.scala 53:83:@29129.4]
  assign buffer_7_599 = $signed(_T_78887); // @[Modules.scala 53:83:@29130.4]
  assign _T_78889 = $signed(buffer_7_416) + $signed(buffer_2_417); // @[Modules.scala 53:83:@29132.4]
  assign _T_78890 = _T_78889[10:0]; // @[Modules.scala 53:83:@29133.4]
  assign buffer_7_600 = $signed(_T_78890); // @[Modules.scala 53:83:@29134.4]
  assign _T_78892 = $signed(buffer_0_418) + $signed(buffer_6_419); // @[Modules.scala 53:83:@29136.4]
  assign _T_78893 = _T_78892[10:0]; // @[Modules.scala 53:83:@29137.4]
  assign buffer_7_601 = $signed(_T_78893); // @[Modules.scala 53:83:@29138.4]
  assign _T_78895 = $signed(buffer_0_420) + $signed(buffer_7_421); // @[Modules.scala 53:83:@29140.4]
  assign _T_78896 = _T_78895[10:0]; // @[Modules.scala 53:83:@29141.4]
  assign buffer_7_602 = $signed(_T_78896); // @[Modules.scala 53:83:@29142.4]
  assign _T_78898 = $signed(buffer_7_422) + $signed(buffer_7_423); // @[Modules.scala 53:83:@29144.4]
  assign _T_78899 = _T_78898[10:0]; // @[Modules.scala 53:83:@29145.4]
  assign buffer_7_603 = $signed(_T_78899); // @[Modules.scala 53:83:@29146.4]
  assign _T_78901 = $signed(buffer_4_424) + $signed(buffer_7_425); // @[Modules.scala 53:83:@29148.4]
  assign _T_78902 = _T_78901[10:0]; // @[Modules.scala 53:83:@29149.4]
  assign buffer_7_604 = $signed(_T_78902); // @[Modules.scala 53:83:@29150.4]
  assign _T_78904 = $signed(buffer_4_426) + $signed(buffer_2_427); // @[Modules.scala 53:83:@29152.4]
  assign _T_78905 = _T_78904[10:0]; // @[Modules.scala 53:83:@29153.4]
  assign buffer_7_605 = $signed(_T_78905); // @[Modules.scala 53:83:@29154.4]
  assign _T_78907 = $signed(buffer_7_428) + $signed(buffer_7_429); // @[Modules.scala 53:83:@29156.4]
  assign _T_78908 = _T_78907[10:0]; // @[Modules.scala 53:83:@29157.4]
  assign buffer_7_606 = $signed(_T_78908); // @[Modules.scala 53:83:@29158.4]
  assign _T_78910 = $signed(buffer_7_430) + $signed(buffer_4_431); // @[Modules.scala 53:83:@29160.4]
  assign _T_78911 = _T_78910[10:0]; // @[Modules.scala 53:83:@29161.4]
  assign buffer_7_607 = $signed(_T_78911); // @[Modules.scala 53:83:@29162.4]
  assign _T_78916 = $signed(buffer_2_434) + $signed(buffer_7_435); // @[Modules.scala 53:83:@29168.4]
  assign _T_78917 = _T_78916[10:0]; // @[Modules.scala 53:83:@29169.4]
  assign buffer_7_609 = $signed(_T_78917); // @[Modules.scala 53:83:@29170.4]
  assign _T_78919 = $signed(buffer_7_436) + $signed(buffer_0_437); // @[Modules.scala 53:83:@29172.4]
  assign _T_78920 = _T_78919[10:0]; // @[Modules.scala 53:83:@29173.4]
  assign buffer_7_610 = $signed(_T_78920); // @[Modules.scala 53:83:@29174.4]
  assign _T_78922 = $signed(buffer_2_438) + $signed(buffer_7_439); // @[Modules.scala 53:83:@29176.4]
  assign _T_78923 = _T_78922[10:0]; // @[Modules.scala 53:83:@29177.4]
  assign buffer_7_611 = $signed(_T_78923); // @[Modules.scala 53:83:@29178.4]
  assign _T_78925 = $signed(buffer_2_440) + $signed(buffer_0_441); // @[Modules.scala 53:83:@29180.4]
  assign _T_78926 = _T_78925[10:0]; // @[Modules.scala 53:83:@29181.4]
  assign buffer_7_612 = $signed(_T_78926); // @[Modules.scala 53:83:@29182.4]
  assign _T_78928 = $signed(buffer_1_442) + $signed(buffer_5_443); // @[Modules.scala 53:83:@29184.4]
  assign _T_78929 = _T_78928[10:0]; // @[Modules.scala 53:83:@29185.4]
  assign buffer_7_613 = $signed(_T_78929); // @[Modules.scala 53:83:@29186.4]
  assign _T_78934 = $signed(buffer_7_446) + $signed(buffer_2_447); // @[Modules.scala 53:83:@29192.4]
  assign _T_78935 = _T_78934[10:0]; // @[Modules.scala 53:83:@29193.4]
  assign buffer_7_615 = $signed(_T_78935); // @[Modules.scala 53:83:@29194.4]
  assign _T_78937 = $signed(buffer_0_448) + $signed(buffer_7_449); // @[Modules.scala 53:83:@29196.4]
  assign _T_78938 = _T_78937[10:0]; // @[Modules.scala 53:83:@29197.4]
  assign buffer_7_616 = $signed(_T_78938); // @[Modules.scala 53:83:@29198.4]
  assign _T_78940 = $signed(buffer_7_450) + $signed(buffer_1_451); // @[Modules.scala 53:83:@29200.4]
  assign _T_78941 = _T_78940[10:0]; // @[Modules.scala 53:83:@29201.4]
  assign buffer_7_617 = $signed(_T_78941); // @[Modules.scala 53:83:@29202.4]
  assign _T_78943 = $signed(buffer_4_452) + $signed(buffer_7_453); // @[Modules.scala 53:83:@29204.4]
  assign _T_78944 = _T_78943[10:0]; // @[Modules.scala 53:83:@29205.4]
  assign buffer_7_618 = $signed(_T_78944); // @[Modules.scala 53:83:@29206.4]
  assign _T_78952 = $signed(buffer_0_458) + $signed(buffer_7_459); // @[Modules.scala 53:83:@29216.4]
  assign _T_78953 = _T_78952[10:0]; // @[Modules.scala 53:83:@29217.4]
  assign buffer_7_621 = $signed(_T_78953); // @[Modules.scala 53:83:@29218.4]
  assign _T_78955 = $signed(buffer_7_460) + $signed(buffer_1_461); // @[Modules.scala 53:83:@29220.4]
  assign _T_78956 = _T_78955[10:0]; // @[Modules.scala 53:83:@29221.4]
  assign buffer_7_622 = $signed(_T_78956); // @[Modules.scala 53:83:@29222.4]
  assign _T_78958 = $signed(buffer_0_462) + $signed(buffer_7_463); // @[Modules.scala 53:83:@29224.4]
  assign _T_78959 = _T_78958[10:0]; // @[Modules.scala 53:83:@29225.4]
  assign buffer_7_623 = $signed(_T_78959); // @[Modules.scala 53:83:@29226.4]
  assign _T_78961 = $signed(buffer_7_464) + $signed(buffer_7_465); // @[Modules.scala 53:83:@29228.4]
  assign _T_78962 = _T_78961[10:0]; // @[Modules.scala 53:83:@29229.4]
  assign buffer_7_624 = $signed(_T_78962); // @[Modules.scala 53:83:@29230.4]
  assign _T_78970 = $signed(buffer_7_470) + $signed(buffer_7_471); // @[Modules.scala 53:83:@29240.4]
  assign _T_78971 = _T_78970[10:0]; // @[Modules.scala 53:83:@29241.4]
  assign buffer_7_627 = $signed(_T_78971); // @[Modules.scala 53:83:@29242.4]
  assign _T_78979 = $signed(buffer_7_476) + $signed(buffer_6_477); // @[Modules.scala 53:83:@29252.4]
  assign _T_78980 = _T_78979[10:0]; // @[Modules.scala 53:83:@29253.4]
  assign buffer_7_630 = $signed(_T_78980); // @[Modules.scala 53:83:@29254.4]
  assign _T_78985 = $signed(buffer_1_480) + $signed(buffer_7_481); // @[Modules.scala 53:83:@29260.4]
  assign _T_78986 = _T_78985[10:0]; // @[Modules.scala 53:83:@29261.4]
  assign buffer_7_632 = $signed(_T_78986); // @[Modules.scala 53:83:@29262.4]
  assign _T_78988 = $signed(buffer_2_482) + $signed(buffer_7_483); // @[Modules.scala 53:83:@29264.4]
  assign _T_78989 = _T_78988[10:0]; // @[Modules.scala 53:83:@29265.4]
  assign buffer_7_633 = $signed(_T_78989); // @[Modules.scala 53:83:@29266.4]
  assign _T_78994 = $signed(buffer_0_486) + $signed(buffer_7_487); // @[Modules.scala 53:83:@29272.4]
  assign _T_78995 = _T_78994[10:0]; // @[Modules.scala 53:83:@29273.4]
  assign buffer_7_635 = $signed(_T_78995); // @[Modules.scala 53:83:@29274.4]
  assign _T_79000 = $signed(buffer_7_490) + $signed(buffer_7_491); // @[Modules.scala 53:83:@29280.4]
  assign _T_79001 = _T_79000[10:0]; // @[Modules.scala 53:83:@29281.4]
  assign buffer_7_637 = $signed(_T_79001); // @[Modules.scala 53:83:@29282.4]
  assign _T_79003 = $signed(buffer_7_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@29284.4]
  assign _T_79004 = _T_79003[10:0]; // @[Modules.scala 53:83:@29285.4]
  assign buffer_7_638 = $signed(_T_79004); // @[Modules.scala 53:83:@29286.4]
  assign _T_79006 = $signed(buffer_7_494) + $signed(buffer_3_495); // @[Modules.scala 53:83:@29288.4]
  assign _T_79007 = _T_79006[10:0]; // @[Modules.scala 53:83:@29289.4]
  assign buffer_7_639 = $signed(_T_79007); // @[Modules.scala 53:83:@29290.4]
  assign _T_79009 = $signed(buffer_5_496) + $signed(buffer_7_497); // @[Modules.scala 53:83:@29292.4]
  assign _T_79010 = _T_79009[10:0]; // @[Modules.scala 53:83:@29293.4]
  assign buffer_7_640 = $signed(_T_79010); // @[Modules.scala 53:83:@29294.4]
  assign _T_79012 = $signed(buffer_7_498) + $signed(buffer_7_499); // @[Modules.scala 53:83:@29296.4]
  assign _T_79013 = _T_79012[10:0]; // @[Modules.scala 53:83:@29297.4]
  assign buffer_7_641 = $signed(_T_79013); // @[Modules.scala 53:83:@29298.4]
  assign _T_79015 = $signed(buffer_0_500) + $signed(buffer_7_501); // @[Modules.scala 53:83:@29300.4]
  assign _T_79016 = _T_79015[10:0]; // @[Modules.scala 53:83:@29301.4]
  assign buffer_7_642 = $signed(_T_79016); // @[Modules.scala 53:83:@29302.4]
  assign _T_79018 = $signed(buffer_3_502) + $signed(buffer_5_503); // @[Modules.scala 53:83:@29304.4]
  assign _T_79019 = _T_79018[10:0]; // @[Modules.scala 53:83:@29305.4]
  assign buffer_7_643 = $signed(_T_79019); // @[Modules.scala 53:83:@29306.4]
  assign _T_79021 = $signed(buffer_7_504) + $signed(buffer_1_505); // @[Modules.scala 53:83:@29308.4]
  assign _T_79022 = _T_79021[10:0]; // @[Modules.scala 53:83:@29309.4]
  assign buffer_7_644 = $signed(_T_79022); // @[Modules.scala 53:83:@29310.4]
  assign _T_79024 = $signed(buffer_7_506) + $signed(buffer_2_507); // @[Modules.scala 53:83:@29312.4]
  assign _T_79025 = _T_79024[10:0]; // @[Modules.scala 53:83:@29313.4]
  assign buffer_7_645 = $signed(_T_79025); // @[Modules.scala 53:83:@29314.4]
  assign _T_79027 = $signed(buffer_5_508) + $signed(buffer_7_509); // @[Modules.scala 53:83:@29316.4]
  assign _T_79028 = _T_79027[10:0]; // @[Modules.scala 53:83:@29317.4]
  assign buffer_7_646 = $signed(_T_79028); // @[Modules.scala 53:83:@29318.4]
  assign _T_79030 = $signed(buffer_3_510) + $signed(buffer_7_511); // @[Modules.scala 53:83:@29320.4]
  assign _T_79031 = _T_79030[10:0]; // @[Modules.scala 53:83:@29321.4]
  assign buffer_7_647 = $signed(_T_79031); // @[Modules.scala 53:83:@29322.4]
  assign _T_79033 = $signed(buffer_7_512) + $signed(buffer_2_513); // @[Modules.scala 53:83:@29324.4]
  assign _T_79034 = _T_79033[10:0]; // @[Modules.scala 53:83:@29325.4]
  assign buffer_7_648 = $signed(_T_79034); // @[Modules.scala 53:83:@29326.4]
  assign _T_79036 = $signed(buffer_2_514) + $signed(buffer_7_515); // @[Modules.scala 53:83:@29328.4]
  assign _T_79037 = _T_79036[10:0]; // @[Modules.scala 53:83:@29329.4]
  assign buffer_7_649 = $signed(_T_79037); // @[Modules.scala 53:83:@29330.4]
  assign _T_79039 = $signed(buffer_5_516) + $signed(buffer_7_517); // @[Modules.scala 53:83:@29332.4]
  assign _T_79040 = _T_79039[10:0]; // @[Modules.scala 53:83:@29333.4]
  assign buffer_7_650 = $signed(_T_79040); // @[Modules.scala 53:83:@29334.4]
  assign _T_79042 = $signed(buffer_2_518) + $signed(buffer_3_519); // @[Modules.scala 53:83:@29336.4]
  assign _T_79043 = _T_79042[10:0]; // @[Modules.scala 53:83:@29337.4]
  assign buffer_7_651 = $signed(_T_79043); // @[Modules.scala 53:83:@29338.4]
  assign _T_79045 = $signed(buffer_0_520) + $signed(buffer_5_521); // @[Modules.scala 53:83:@29340.4]
  assign _T_79046 = _T_79045[10:0]; // @[Modules.scala 53:83:@29341.4]
  assign buffer_7_652 = $signed(_T_79046); // @[Modules.scala 53:83:@29342.4]
  assign _T_79048 = $signed(buffer_7_522) + $signed(buffer_7_523); // @[Modules.scala 53:83:@29344.4]
  assign _T_79049 = _T_79048[10:0]; // @[Modules.scala 53:83:@29345.4]
  assign buffer_7_653 = $signed(_T_79049); // @[Modules.scala 53:83:@29346.4]
  assign _T_79051 = $signed(buffer_3_524) + $signed(buffer_2_525); // @[Modules.scala 53:83:@29348.4]
  assign _T_79052 = _T_79051[10:0]; // @[Modules.scala 53:83:@29349.4]
  assign buffer_7_654 = $signed(_T_79052); // @[Modules.scala 53:83:@29350.4]
  assign _T_79054 = $signed(buffer_7_526) + $signed(buffer_1_527); // @[Modules.scala 53:83:@29352.4]
  assign _T_79055 = _T_79054[10:0]; // @[Modules.scala 53:83:@29353.4]
  assign buffer_7_655 = $signed(_T_79055); // @[Modules.scala 53:83:@29354.4]
  assign _T_79057 = $signed(buffer_7_528) + $signed(buffer_7_529); // @[Modules.scala 53:83:@29356.4]
  assign _T_79058 = _T_79057[10:0]; // @[Modules.scala 53:83:@29357.4]
  assign buffer_7_656 = $signed(_T_79058); // @[Modules.scala 53:83:@29358.4]
  assign _T_79060 = $signed(buffer_7_530) + $signed(buffer_5_531); // @[Modules.scala 53:83:@29360.4]
  assign _T_79061 = _T_79060[10:0]; // @[Modules.scala 53:83:@29361.4]
  assign buffer_7_657 = $signed(_T_79061); // @[Modules.scala 53:83:@29362.4]
  assign _T_79063 = $signed(buffer_2_532) + $signed(buffer_7_533); // @[Modules.scala 53:83:@29364.4]
  assign _T_79064 = _T_79063[10:0]; // @[Modules.scala 53:83:@29365.4]
  assign buffer_7_658 = $signed(_T_79064); // @[Modules.scala 53:83:@29366.4]
  assign _T_79069 = $signed(buffer_2_536) + $signed(buffer_3_537); // @[Modules.scala 53:83:@29372.4]
  assign _T_79070 = _T_79069[10:0]; // @[Modules.scala 53:83:@29373.4]
  assign buffer_7_660 = $signed(_T_79070); // @[Modules.scala 53:83:@29374.4]
  assign _T_79072 = $signed(buffer_7_538) + $signed(buffer_7_539); // @[Modules.scala 53:83:@29376.4]
  assign _T_79073 = _T_79072[10:0]; // @[Modules.scala 53:83:@29377.4]
  assign buffer_7_661 = $signed(_T_79073); // @[Modules.scala 53:83:@29378.4]
  assign _T_79075 = $signed(buffer_2_540) + $signed(buffer_7_541); // @[Modules.scala 53:83:@29380.4]
  assign _T_79076 = _T_79075[10:0]; // @[Modules.scala 53:83:@29381.4]
  assign buffer_7_662 = $signed(_T_79076); // @[Modules.scala 53:83:@29382.4]
  assign _T_79078 = $signed(buffer_7_542) + $signed(buffer_3_543); // @[Modules.scala 53:83:@29384.4]
  assign _T_79079 = _T_79078[10:0]; // @[Modules.scala 53:83:@29385.4]
  assign buffer_7_663 = $signed(_T_79079); // @[Modules.scala 53:83:@29386.4]
  assign _T_79081 = $signed(buffer_3_544) + $signed(buffer_7_545); // @[Modules.scala 53:83:@29388.4]
  assign _T_79082 = _T_79081[10:0]; // @[Modules.scala 53:83:@29389.4]
  assign buffer_7_664 = $signed(_T_79082); // @[Modules.scala 53:83:@29390.4]
  assign _T_79084 = $signed(buffer_7_546) + $signed(buffer_7_547); // @[Modules.scala 53:83:@29392.4]
  assign _T_79085 = _T_79084[10:0]; // @[Modules.scala 53:83:@29393.4]
  assign buffer_7_665 = $signed(_T_79085); // @[Modules.scala 53:83:@29394.4]
  assign _T_79087 = $signed(buffer_7_548) + $signed(buffer_0_549); // @[Modules.scala 53:83:@29396.4]
  assign _T_79088 = _T_79087[10:0]; // @[Modules.scala 53:83:@29397.4]
  assign buffer_7_666 = $signed(_T_79088); // @[Modules.scala 53:83:@29398.4]
  assign _T_79090 = $signed(buffer_7_550) + $signed(buffer_3_551); // @[Modules.scala 53:83:@29400.4]
  assign _T_79091 = _T_79090[10:0]; // @[Modules.scala 53:83:@29401.4]
  assign buffer_7_667 = $signed(_T_79091); // @[Modules.scala 53:83:@29402.4]
  assign _T_79093 = $signed(buffer_3_552) + $signed(buffer_7_553); // @[Modules.scala 53:83:@29404.4]
  assign _T_79094 = _T_79093[10:0]; // @[Modules.scala 53:83:@29405.4]
  assign buffer_7_668 = $signed(_T_79094); // @[Modules.scala 53:83:@29406.4]
  assign _T_79096 = $signed(buffer_0_554) + $signed(buffer_5_555); // @[Modules.scala 53:83:@29408.4]
  assign _T_79097 = _T_79096[10:0]; // @[Modules.scala 53:83:@29409.4]
  assign buffer_7_669 = $signed(_T_79097); // @[Modules.scala 53:83:@29410.4]
  assign _T_79099 = $signed(buffer_7_556) + $signed(buffer_4_557); // @[Modules.scala 53:83:@29412.4]
  assign _T_79100 = _T_79099[10:0]; // @[Modules.scala 53:83:@29413.4]
  assign buffer_7_670 = $signed(_T_79100); // @[Modules.scala 53:83:@29414.4]
  assign _T_79102 = $signed(buffer_7_558) + $signed(buffer_7_559); // @[Modules.scala 53:83:@29416.4]
  assign _T_79103 = _T_79102[10:0]; // @[Modules.scala 53:83:@29417.4]
  assign buffer_7_671 = $signed(_T_79103); // @[Modules.scala 53:83:@29418.4]
  assign _T_79105 = $signed(buffer_7_560) + $signed(buffer_2_561); // @[Modules.scala 53:83:@29420.4]
  assign _T_79106 = _T_79105[10:0]; // @[Modules.scala 53:83:@29421.4]
  assign buffer_7_672 = $signed(_T_79106); // @[Modules.scala 53:83:@29422.4]
  assign _T_79108 = $signed(buffer_2_562) + $signed(buffer_7_563); // @[Modules.scala 53:83:@29424.4]
  assign _T_79109 = _T_79108[10:0]; // @[Modules.scala 53:83:@29425.4]
  assign buffer_7_673 = $signed(_T_79109); // @[Modules.scala 53:83:@29426.4]
  assign _T_79111 = $signed(buffer_7_564) + $signed(buffer_3_565); // @[Modules.scala 53:83:@29428.4]
  assign _T_79112 = _T_79111[10:0]; // @[Modules.scala 53:83:@29429.4]
  assign buffer_7_674 = $signed(_T_79112); // @[Modules.scala 53:83:@29430.4]
  assign _T_79114 = $signed(buffer_7_566) + $signed(buffer_7_567); // @[Modules.scala 53:83:@29432.4]
  assign _T_79115 = _T_79114[10:0]; // @[Modules.scala 53:83:@29433.4]
  assign buffer_7_675 = $signed(_T_79115); // @[Modules.scala 53:83:@29434.4]
  assign _T_79123 = $signed(buffer_3_572) + $signed(buffer_7_573); // @[Modules.scala 53:83:@29444.4]
  assign _T_79124 = _T_79123[10:0]; // @[Modules.scala 53:83:@29445.4]
  assign buffer_7_678 = $signed(_T_79124); // @[Modules.scala 53:83:@29446.4]
  assign _T_79135 = $signed(buffer_7_580) + $signed(buffer_1_581); // @[Modules.scala 53:83:@29460.4]
  assign _T_79136 = _T_79135[10:0]; // @[Modules.scala 53:83:@29461.4]
  assign buffer_7_682 = $signed(_T_79136); // @[Modules.scala 53:83:@29462.4]
  assign _T_79138 = $signed(buffer_7_582) + $signed(buffer_4_583); // @[Modules.scala 53:83:@29464.4]
  assign _T_79139 = _T_79138[10:0]; // @[Modules.scala 53:83:@29465.4]
  assign buffer_7_683 = $signed(_T_79139); // @[Modules.scala 53:83:@29466.4]
  assign _T_79144 = $signed(buffer_1_586) + $signed(buffer_7_587); // @[Modules.scala 53:83:@29472.4]
  assign _T_79145 = _T_79144[10:0]; // @[Modules.scala 53:83:@29473.4]
  assign buffer_7_685 = $signed(_T_79145); // @[Modules.scala 53:83:@29474.4]
  assign _T_79147 = $signed(buffer_7_588) + $signed(buffer_2_589); // @[Modules.scala 56:109:@29476.4]
  assign _T_79148 = _T_79147[10:0]; // @[Modules.scala 56:109:@29477.4]
  assign buffer_7_686 = $signed(_T_79148); // @[Modules.scala 56:109:@29478.4]
  assign _T_79150 = $signed(buffer_7_590) + $signed(buffer_7_591); // @[Modules.scala 56:109:@29480.4]
  assign _T_79151 = _T_79150[10:0]; // @[Modules.scala 56:109:@29481.4]
  assign buffer_7_687 = $signed(_T_79151); // @[Modules.scala 56:109:@29482.4]
  assign _T_79153 = $signed(buffer_7_592) + $signed(buffer_7_593); // @[Modules.scala 56:109:@29484.4]
  assign _T_79154 = _T_79153[10:0]; // @[Modules.scala 56:109:@29485.4]
  assign buffer_7_688 = $signed(_T_79154); // @[Modules.scala 56:109:@29486.4]
  assign _T_79156 = $signed(buffer_7_594) + $signed(buffer_7_595); // @[Modules.scala 56:109:@29488.4]
  assign _T_79157 = _T_79156[10:0]; // @[Modules.scala 56:109:@29489.4]
  assign buffer_7_689 = $signed(_T_79157); // @[Modules.scala 56:109:@29490.4]
  assign _T_79162 = $signed(buffer_7_598) + $signed(buffer_7_599); // @[Modules.scala 56:109:@29496.4]
  assign _T_79163 = _T_79162[10:0]; // @[Modules.scala 56:109:@29497.4]
  assign buffer_7_691 = $signed(_T_79163); // @[Modules.scala 56:109:@29498.4]
  assign _T_79165 = $signed(buffer_7_600) + $signed(buffer_7_601); // @[Modules.scala 56:109:@29500.4]
  assign _T_79166 = _T_79165[10:0]; // @[Modules.scala 56:109:@29501.4]
  assign buffer_7_692 = $signed(_T_79166); // @[Modules.scala 56:109:@29502.4]
  assign _T_79168 = $signed(buffer_7_602) + $signed(buffer_7_603); // @[Modules.scala 56:109:@29504.4]
  assign _T_79169 = _T_79168[10:0]; // @[Modules.scala 56:109:@29505.4]
  assign buffer_7_693 = $signed(_T_79169); // @[Modules.scala 56:109:@29506.4]
  assign _T_79171 = $signed(buffer_7_604) + $signed(buffer_7_605); // @[Modules.scala 56:109:@29508.4]
  assign _T_79172 = _T_79171[10:0]; // @[Modules.scala 56:109:@29509.4]
  assign buffer_7_694 = $signed(_T_79172); // @[Modules.scala 56:109:@29510.4]
  assign _T_79174 = $signed(buffer_7_606) + $signed(buffer_7_607); // @[Modules.scala 56:109:@29512.4]
  assign _T_79175 = _T_79174[10:0]; // @[Modules.scala 56:109:@29513.4]
  assign buffer_7_695 = $signed(_T_79175); // @[Modules.scala 56:109:@29514.4]
  assign _T_79177 = $signed(buffer_2_608) + $signed(buffer_7_609); // @[Modules.scala 56:109:@29516.4]
  assign _T_79178 = _T_79177[10:0]; // @[Modules.scala 56:109:@29517.4]
  assign buffer_7_696 = $signed(_T_79178); // @[Modules.scala 56:109:@29518.4]
  assign _T_79180 = $signed(buffer_7_610) + $signed(buffer_7_611); // @[Modules.scala 56:109:@29520.4]
  assign _T_79181 = _T_79180[10:0]; // @[Modules.scala 56:109:@29521.4]
  assign buffer_7_697 = $signed(_T_79181); // @[Modules.scala 56:109:@29522.4]
  assign _T_79183 = $signed(buffer_7_612) + $signed(buffer_7_613); // @[Modules.scala 56:109:@29524.4]
  assign _T_79184 = _T_79183[10:0]; // @[Modules.scala 56:109:@29525.4]
  assign buffer_7_698 = $signed(_T_79184); // @[Modules.scala 56:109:@29526.4]
  assign _T_79186 = $signed(buffer_4_614) + $signed(buffer_7_615); // @[Modules.scala 56:109:@29528.4]
  assign _T_79187 = _T_79186[10:0]; // @[Modules.scala 56:109:@29529.4]
  assign buffer_7_699 = $signed(_T_79187); // @[Modules.scala 56:109:@29530.4]
  assign _T_79189 = $signed(buffer_7_616) + $signed(buffer_7_617); // @[Modules.scala 56:109:@29532.4]
  assign _T_79190 = _T_79189[10:0]; // @[Modules.scala 56:109:@29533.4]
  assign buffer_7_700 = $signed(_T_79190); // @[Modules.scala 56:109:@29534.4]
  assign _T_79192 = $signed(buffer_7_618) + $signed(buffer_2_619); // @[Modules.scala 56:109:@29536.4]
  assign _T_79193 = _T_79192[10:0]; // @[Modules.scala 56:109:@29537.4]
  assign buffer_7_701 = $signed(_T_79193); // @[Modules.scala 56:109:@29538.4]
  assign _T_79195 = $signed(buffer_2_620) + $signed(buffer_7_621); // @[Modules.scala 56:109:@29540.4]
  assign _T_79196 = _T_79195[10:0]; // @[Modules.scala 56:109:@29541.4]
  assign buffer_7_702 = $signed(_T_79196); // @[Modules.scala 56:109:@29542.4]
  assign _T_79198 = $signed(buffer_7_622) + $signed(buffer_7_623); // @[Modules.scala 56:109:@29544.4]
  assign _T_79199 = _T_79198[10:0]; // @[Modules.scala 56:109:@29545.4]
  assign buffer_7_703 = $signed(_T_79199); // @[Modules.scala 56:109:@29546.4]
  assign _T_79201 = $signed(buffer_7_624) + $signed(buffer_0_625); // @[Modules.scala 56:109:@29548.4]
  assign _T_79202 = _T_79201[10:0]; // @[Modules.scala 56:109:@29549.4]
  assign buffer_7_704 = $signed(_T_79202); // @[Modules.scala 56:109:@29550.4]
  assign _T_79204 = $signed(buffer_1_626) + $signed(buffer_7_627); // @[Modules.scala 56:109:@29552.4]
  assign _T_79205 = _T_79204[10:0]; // @[Modules.scala 56:109:@29553.4]
  assign buffer_7_705 = $signed(_T_79205); // @[Modules.scala 56:109:@29554.4]
  assign _T_79207 = $signed(buffer_4_628) + $signed(buffer_2_629); // @[Modules.scala 56:109:@29556.4]
  assign _T_79208 = _T_79207[10:0]; // @[Modules.scala 56:109:@29557.4]
  assign buffer_7_706 = $signed(_T_79208); // @[Modules.scala 56:109:@29558.4]
  assign _T_79210 = $signed(buffer_7_630) + $signed(buffer_1_631); // @[Modules.scala 56:109:@29560.4]
  assign _T_79211 = _T_79210[10:0]; // @[Modules.scala 56:109:@29561.4]
  assign buffer_7_707 = $signed(_T_79211); // @[Modules.scala 56:109:@29562.4]
  assign _T_79213 = $signed(buffer_7_632) + $signed(buffer_7_633); // @[Modules.scala 56:109:@29564.4]
  assign _T_79214 = _T_79213[10:0]; // @[Modules.scala 56:109:@29565.4]
  assign buffer_7_708 = $signed(_T_79214); // @[Modules.scala 56:109:@29566.4]
  assign _T_79216 = $signed(buffer_4_634) + $signed(buffer_7_635); // @[Modules.scala 56:109:@29568.4]
  assign _T_79217 = _T_79216[10:0]; // @[Modules.scala 56:109:@29569.4]
  assign buffer_7_709 = $signed(_T_79217); // @[Modules.scala 56:109:@29570.4]
  assign _T_79219 = $signed(buffer_3_636) + $signed(buffer_7_637); // @[Modules.scala 56:109:@29572.4]
  assign _T_79220 = _T_79219[10:0]; // @[Modules.scala 56:109:@29573.4]
  assign buffer_7_710 = $signed(_T_79220); // @[Modules.scala 56:109:@29574.4]
  assign _T_79222 = $signed(buffer_7_638) + $signed(buffer_7_639); // @[Modules.scala 56:109:@29576.4]
  assign _T_79223 = _T_79222[10:0]; // @[Modules.scala 56:109:@29577.4]
  assign buffer_7_711 = $signed(_T_79223); // @[Modules.scala 56:109:@29578.4]
  assign _T_79225 = $signed(buffer_7_640) + $signed(buffer_7_641); // @[Modules.scala 56:109:@29580.4]
  assign _T_79226 = _T_79225[10:0]; // @[Modules.scala 56:109:@29581.4]
  assign buffer_7_712 = $signed(_T_79226); // @[Modules.scala 56:109:@29582.4]
  assign _T_79228 = $signed(buffer_7_642) + $signed(buffer_7_643); // @[Modules.scala 56:109:@29584.4]
  assign _T_79229 = _T_79228[10:0]; // @[Modules.scala 56:109:@29585.4]
  assign buffer_7_713 = $signed(_T_79229); // @[Modules.scala 56:109:@29586.4]
  assign _T_79231 = $signed(buffer_7_644) + $signed(buffer_7_645); // @[Modules.scala 56:109:@29588.4]
  assign _T_79232 = _T_79231[10:0]; // @[Modules.scala 56:109:@29589.4]
  assign buffer_7_714 = $signed(_T_79232); // @[Modules.scala 56:109:@29590.4]
  assign _T_79234 = $signed(buffer_7_646) + $signed(buffer_7_647); // @[Modules.scala 56:109:@29592.4]
  assign _T_79235 = _T_79234[10:0]; // @[Modules.scala 56:109:@29593.4]
  assign buffer_7_715 = $signed(_T_79235); // @[Modules.scala 56:109:@29594.4]
  assign _T_79237 = $signed(buffer_7_648) + $signed(buffer_7_649); // @[Modules.scala 56:109:@29596.4]
  assign _T_79238 = _T_79237[10:0]; // @[Modules.scala 56:109:@29597.4]
  assign buffer_7_716 = $signed(_T_79238); // @[Modules.scala 56:109:@29598.4]
  assign _T_79240 = $signed(buffer_7_650) + $signed(buffer_7_651); // @[Modules.scala 56:109:@29600.4]
  assign _T_79241 = _T_79240[10:0]; // @[Modules.scala 56:109:@29601.4]
  assign buffer_7_717 = $signed(_T_79241); // @[Modules.scala 56:109:@29602.4]
  assign _T_79243 = $signed(buffer_7_652) + $signed(buffer_7_653); // @[Modules.scala 56:109:@29604.4]
  assign _T_79244 = _T_79243[10:0]; // @[Modules.scala 56:109:@29605.4]
  assign buffer_7_718 = $signed(_T_79244); // @[Modules.scala 56:109:@29606.4]
  assign _T_79246 = $signed(buffer_7_654) + $signed(buffer_7_655); // @[Modules.scala 56:109:@29608.4]
  assign _T_79247 = _T_79246[10:0]; // @[Modules.scala 56:109:@29609.4]
  assign buffer_7_719 = $signed(_T_79247); // @[Modules.scala 56:109:@29610.4]
  assign _T_79249 = $signed(buffer_7_656) + $signed(buffer_7_657); // @[Modules.scala 56:109:@29612.4]
  assign _T_79250 = _T_79249[10:0]; // @[Modules.scala 56:109:@29613.4]
  assign buffer_7_720 = $signed(_T_79250); // @[Modules.scala 56:109:@29614.4]
  assign _T_79252 = $signed(buffer_7_658) + $signed(buffer_3_659); // @[Modules.scala 56:109:@29616.4]
  assign _T_79253 = _T_79252[10:0]; // @[Modules.scala 56:109:@29617.4]
  assign buffer_7_721 = $signed(_T_79253); // @[Modules.scala 56:109:@29618.4]
  assign _T_79255 = $signed(buffer_7_660) + $signed(buffer_7_661); // @[Modules.scala 56:109:@29620.4]
  assign _T_79256 = _T_79255[10:0]; // @[Modules.scala 56:109:@29621.4]
  assign buffer_7_722 = $signed(_T_79256); // @[Modules.scala 56:109:@29622.4]
  assign _T_79258 = $signed(buffer_7_662) + $signed(buffer_7_663); // @[Modules.scala 56:109:@29624.4]
  assign _T_79259 = _T_79258[10:0]; // @[Modules.scala 56:109:@29625.4]
  assign buffer_7_723 = $signed(_T_79259); // @[Modules.scala 56:109:@29626.4]
  assign _T_79261 = $signed(buffer_7_664) + $signed(buffer_7_665); // @[Modules.scala 56:109:@29628.4]
  assign _T_79262 = _T_79261[10:0]; // @[Modules.scala 56:109:@29629.4]
  assign buffer_7_724 = $signed(_T_79262); // @[Modules.scala 56:109:@29630.4]
  assign _T_79264 = $signed(buffer_7_666) + $signed(buffer_7_667); // @[Modules.scala 56:109:@29632.4]
  assign _T_79265 = _T_79264[10:0]; // @[Modules.scala 56:109:@29633.4]
  assign buffer_7_725 = $signed(_T_79265); // @[Modules.scala 56:109:@29634.4]
  assign _T_79267 = $signed(buffer_7_668) + $signed(buffer_7_669); // @[Modules.scala 56:109:@29636.4]
  assign _T_79268 = _T_79267[10:0]; // @[Modules.scala 56:109:@29637.4]
  assign buffer_7_726 = $signed(_T_79268); // @[Modules.scala 56:109:@29638.4]
  assign _T_79270 = $signed(buffer_7_670) + $signed(buffer_7_671); // @[Modules.scala 56:109:@29640.4]
  assign _T_79271 = _T_79270[10:0]; // @[Modules.scala 56:109:@29641.4]
  assign buffer_7_727 = $signed(_T_79271); // @[Modules.scala 56:109:@29642.4]
  assign _T_79273 = $signed(buffer_7_672) + $signed(buffer_7_673); // @[Modules.scala 56:109:@29644.4]
  assign _T_79274 = _T_79273[10:0]; // @[Modules.scala 56:109:@29645.4]
  assign buffer_7_728 = $signed(_T_79274); // @[Modules.scala 56:109:@29646.4]
  assign _T_79276 = $signed(buffer_7_674) + $signed(buffer_7_675); // @[Modules.scala 56:109:@29648.4]
  assign _T_79277 = _T_79276[10:0]; // @[Modules.scala 56:109:@29649.4]
  assign buffer_7_729 = $signed(_T_79277); // @[Modules.scala 56:109:@29650.4]
  assign _T_79282 = $signed(buffer_7_678) + $signed(buffer_1_679); // @[Modules.scala 56:109:@29656.4]
  assign _T_79283 = _T_79282[10:0]; // @[Modules.scala 56:109:@29657.4]
  assign buffer_7_731 = $signed(_T_79283); // @[Modules.scala 56:109:@29658.4]
  assign _T_79288 = $signed(buffer_7_682) + $signed(buffer_7_683); // @[Modules.scala 56:109:@29664.4]
  assign _T_79289 = _T_79288[10:0]; // @[Modules.scala 56:109:@29665.4]
  assign buffer_7_733 = $signed(_T_79289); // @[Modules.scala 56:109:@29666.4]
  assign _T_79291 = $signed(buffer_1_684) + $signed(buffer_7_685); // @[Modules.scala 56:109:@29668.4]
  assign _T_79292 = _T_79291[10:0]; // @[Modules.scala 56:109:@29669.4]
  assign buffer_7_734 = $signed(_T_79292); // @[Modules.scala 56:109:@29670.4]
  assign _T_79294 = $signed(buffer_7_686) + $signed(buffer_7_687); // @[Modules.scala 63:156:@29673.4]
  assign _T_79295 = _T_79294[10:0]; // @[Modules.scala 63:156:@29674.4]
  assign buffer_7_736 = $signed(_T_79295); // @[Modules.scala 63:156:@29675.4]
  assign _T_79297 = $signed(buffer_7_736) + $signed(buffer_7_688); // @[Modules.scala 63:156:@29677.4]
  assign _T_79298 = _T_79297[10:0]; // @[Modules.scala 63:156:@29678.4]
  assign buffer_7_737 = $signed(_T_79298); // @[Modules.scala 63:156:@29679.4]
  assign _T_79300 = $signed(buffer_7_737) + $signed(buffer_7_689); // @[Modules.scala 63:156:@29681.4]
  assign _T_79301 = _T_79300[10:0]; // @[Modules.scala 63:156:@29682.4]
  assign buffer_7_738 = $signed(_T_79301); // @[Modules.scala 63:156:@29683.4]
  assign _T_79303 = $signed(buffer_7_738) + $signed(buffer_1_690); // @[Modules.scala 63:156:@29685.4]
  assign _T_79304 = _T_79303[10:0]; // @[Modules.scala 63:156:@29686.4]
  assign buffer_7_739 = $signed(_T_79304); // @[Modules.scala 63:156:@29687.4]
  assign _T_79306 = $signed(buffer_7_739) + $signed(buffer_7_691); // @[Modules.scala 63:156:@29689.4]
  assign _T_79307 = _T_79306[10:0]; // @[Modules.scala 63:156:@29690.4]
  assign buffer_7_740 = $signed(_T_79307); // @[Modules.scala 63:156:@29691.4]
  assign _T_79309 = $signed(buffer_7_740) + $signed(buffer_7_692); // @[Modules.scala 63:156:@29693.4]
  assign _T_79310 = _T_79309[10:0]; // @[Modules.scala 63:156:@29694.4]
  assign buffer_7_741 = $signed(_T_79310); // @[Modules.scala 63:156:@29695.4]
  assign _T_79312 = $signed(buffer_7_741) + $signed(buffer_7_693); // @[Modules.scala 63:156:@29697.4]
  assign _T_79313 = _T_79312[10:0]; // @[Modules.scala 63:156:@29698.4]
  assign buffer_7_742 = $signed(_T_79313); // @[Modules.scala 63:156:@29699.4]
  assign _T_79315 = $signed(buffer_7_742) + $signed(buffer_7_694); // @[Modules.scala 63:156:@29701.4]
  assign _T_79316 = _T_79315[10:0]; // @[Modules.scala 63:156:@29702.4]
  assign buffer_7_743 = $signed(_T_79316); // @[Modules.scala 63:156:@29703.4]
  assign _T_79318 = $signed(buffer_7_743) + $signed(buffer_7_695); // @[Modules.scala 63:156:@29705.4]
  assign _T_79319 = _T_79318[10:0]; // @[Modules.scala 63:156:@29706.4]
  assign buffer_7_744 = $signed(_T_79319); // @[Modules.scala 63:156:@29707.4]
  assign _T_79321 = $signed(buffer_7_744) + $signed(buffer_7_696); // @[Modules.scala 63:156:@29709.4]
  assign _T_79322 = _T_79321[10:0]; // @[Modules.scala 63:156:@29710.4]
  assign buffer_7_745 = $signed(_T_79322); // @[Modules.scala 63:156:@29711.4]
  assign _T_79324 = $signed(buffer_7_745) + $signed(buffer_7_697); // @[Modules.scala 63:156:@29713.4]
  assign _T_79325 = _T_79324[10:0]; // @[Modules.scala 63:156:@29714.4]
  assign buffer_7_746 = $signed(_T_79325); // @[Modules.scala 63:156:@29715.4]
  assign _T_79327 = $signed(buffer_7_746) + $signed(buffer_7_698); // @[Modules.scala 63:156:@29717.4]
  assign _T_79328 = _T_79327[10:0]; // @[Modules.scala 63:156:@29718.4]
  assign buffer_7_747 = $signed(_T_79328); // @[Modules.scala 63:156:@29719.4]
  assign _T_79330 = $signed(buffer_7_747) + $signed(buffer_7_699); // @[Modules.scala 63:156:@29721.4]
  assign _T_79331 = _T_79330[10:0]; // @[Modules.scala 63:156:@29722.4]
  assign buffer_7_748 = $signed(_T_79331); // @[Modules.scala 63:156:@29723.4]
  assign _T_79333 = $signed(buffer_7_748) + $signed(buffer_7_700); // @[Modules.scala 63:156:@29725.4]
  assign _T_79334 = _T_79333[10:0]; // @[Modules.scala 63:156:@29726.4]
  assign buffer_7_749 = $signed(_T_79334); // @[Modules.scala 63:156:@29727.4]
  assign _T_79336 = $signed(buffer_7_749) + $signed(buffer_7_701); // @[Modules.scala 63:156:@29729.4]
  assign _T_79337 = _T_79336[10:0]; // @[Modules.scala 63:156:@29730.4]
  assign buffer_7_750 = $signed(_T_79337); // @[Modules.scala 63:156:@29731.4]
  assign _T_79339 = $signed(buffer_7_750) + $signed(buffer_7_702); // @[Modules.scala 63:156:@29733.4]
  assign _T_79340 = _T_79339[10:0]; // @[Modules.scala 63:156:@29734.4]
  assign buffer_7_751 = $signed(_T_79340); // @[Modules.scala 63:156:@29735.4]
  assign _T_79342 = $signed(buffer_7_751) + $signed(buffer_7_703); // @[Modules.scala 63:156:@29737.4]
  assign _T_79343 = _T_79342[10:0]; // @[Modules.scala 63:156:@29738.4]
  assign buffer_7_752 = $signed(_T_79343); // @[Modules.scala 63:156:@29739.4]
  assign _T_79345 = $signed(buffer_7_752) + $signed(buffer_7_704); // @[Modules.scala 63:156:@29741.4]
  assign _T_79346 = _T_79345[10:0]; // @[Modules.scala 63:156:@29742.4]
  assign buffer_7_753 = $signed(_T_79346); // @[Modules.scala 63:156:@29743.4]
  assign _T_79348 = $signed(buffer_7_753) + $signed(buffer_7_705); // @[Modules.scala 63:156:@29745.4]
  assign _T_79349 = _T_79348[10:0]; // @[Modules.scala 63:156:@29746.4]
  assign buffer_7_754 = $signed(_T_79349); // @[Modules.scala 63:156:@29747.4]
  assign _T_79351 = $signed(buffer_7_754) + $signed(buffer_7_706); // @[Modules.scala 63:156:@29749.4]
  assign _T_79352 = _T_79351[10:0]; // @[Modules.scala 63:156:@29750.4]
  assign buffer_7_755 = $signed(_T_79352); // @[Modules.scala 63:156:@29751.4]
  assign _T_79354 = $signed(buffer_7_755) + $signed(buffer_7_707); // @[Modules.scala 63:156:@29753.4]
  assign _T_79355 = _T_79354[10:0]; // @[Modules.scala 63:156:@29754.4]
  assign buffer_7_756 = $signed(_T_79355); // @[Modules.scala 63:156:@29755.4]
  assign _T_79357 = $signed(buffer_7_756) + $signed(buffer_7_708); // @[Modules.scala 63:156:@29757.4]
  assign _T_79358 = _T_79357[10:0]; // @[Modules.scala 63:156:@29758.4]
  assign buffer_7_757 = $signed(_T_79358); // @[Modules.scala 63:156:@29759.4]
  assign _T_79360 = $signed(buffer_7_757) + $signed(buffer_7_709); // @[Modules.scala 63:156:@29761.4]
  assign _T_79361 = _T_79360[10:0]; // @[Modules.scala 63:156:@29762.4]
  assign buffer_7_758 = $signed(_T_79361); // @[Modules.scala 63:156:@29763.4]
  assign _T_79363 = $signed(buffer_7_758) + $signed(buffer_7_710); // @[Modules.scala 63:156:@29765.4]
  assign _T_79364 = _T_79363[10:0]; // @[Modules.scala 63:156:@29766.4]
  assign buffer_7_759 = $signed(_T_79364); // @[Modules.scala 63:156:@29767.4]
  assign _T_79366 = $signed(buffer_7_759) + $signed(buffer_7_711); // @[Modules.scala 63:156:@29769.4]
  assign _T_79367 = _T_79366[10:0]; // @[Modules.scala 63:156:@29770.4]
  assign buffer_7_760 = $signed(_T_79367); // @[Modules.scala 63:156:@29771.4]
  assign _T_79369 = $signed(buffer_7_760) + $signed(buffer_7_712); // @[Modules.scala 63:156:@29773.4]
  assign _T_79370 = _T_79369[10:0]; // @[Modules.scala 63:156:@29774.4]
  assign buffer_7_761 = $signed(_T_79370); // @[Modules.scala 63:156:@29775.4]
  assign _T_79372 = $signed(buffer_7_761) + $signed(buffer_7_713); // @[Modules.scala 63:156:@29777.4]
  assign _T_79373 = _T_79372[10:0]; // @[Modules.scala 63:156:@29778.4]
  assign buffer_7_762 = $signed(_T_79373); // @[Modules.scala 63:156:@29779.4]
  assign _T_79375 = $signed(buffer_7_762) + $signed(buffer_7_714); // @[Modules.scala 63:156:@29781.4]
  assign _T_79376 = _T_79375[10:0]; // @[Modules.scala 63:156:@29782.4]
  assign buffer_7_763 = $signed(_T_79376); // @[Modules.scala 63:156:@29783.4]
  assign _T_79378 = $signed(buffer_7_763) + $signed(buffer_7_715); // @[Modules.scala 63:156:@29785.4]
  assign _T_79379 = _T_79378[10:0]; // @[Modules.scala 63:156:@29786.4]
  assign buffer_7_764 = $signed(_T_79379); // @[Modules.scala 63:156:@29787.4]
  assign _T_79381 = $signed(buffer_7_764) + $signed(buffer_7_716); // @[Modules.scala 63:156:@29789.4]
  assign _T_79382 = _T_79381[10:0]; // @[Modules.scala 63:156:@29790.4]
  assign buffer_7_765 = $signed(_T_79382); // @[Modules.scala 63:156:@29791.4]
  assign _T_79384 = $signed(buffer_7_765) + $signed(buffer_7_717); // @[Modules.scala 63:156:@29793.4]
  assign _T_79385 = _T_79384[10:0]; // @[Modules.scala 63:156:@29794.4]
  assign buffer_7_766 = $signed(_T_79385); // @[Modules.scala 63:156:@29795.4]
  assign _T_79387 = $signed(buffer_7_766) + $signed(buffer_7_718); // @[Modules.scala 63:156:@29797.4]
  assign _T_79388 = _T_79387[10:0]; // @[Modules.scala 63:156:@29798.4]
  assign buffer_7_767 = $signed(_T_79388); // @[Modules.scala 63:156:@29799.4]
  assign _T_79390 = $signed(buffer_7_767) + $signed(buffer_7_719); // @[Modules.scala 63:156:@29801.4]
  assign _T_79391 = _T_79390[10:0]; // @[Modules.scala 63:156:@29802.4]
  assign buffer_7_768 = $signed(_T_79391); // @[Modules.scala 63:156:@29803.4]
  assign _T_79393 = $signed(buffer_7_768) + $signed(buffer_7_720); // @[Modules.scala 63:156:@29805.4]
  assign _T_79394 = _T_79393[10:0]; // @[Modules.scala 63:156:@29806.4]
  assign buffer_7_769 = $signed(_T_79394); // @[Modules.scala 63:156:@29807.4]
  assign _T_79396 = $signed(buffer_7_769) + $signed(buffer_7_721); // @[Modules.scala 63:156:@29809.4]
  assign _T_79397 = _T_79396[10:0]; // @[Modules.scala 63:156:@29810.4]
  assign buffer_7_770 = $signed(_T_79397); // @[Modules.scala 63:156:@29811.4]
  assign _T_79399 = $signed(buffer_7_770) + $signed(buffer_7_722); // @[Modules.scala 63:156:@29813.4]
  assign _T_79400 = _T_79399[10:0]; // @[Modules.scala 63:156:@29814.4]
  assign buffer_7_771 = $signed(_T_79400); // @[Modules.scala 63:156:@29815.4]
  assign _T_79402 = $signed(buffer_7_771) + $signed(buffer_7_723); // @[Modules.scala 63:156:@29817.4]
  assign _T_79403 = _T_79402[10:0]; // @[Modules.scala 63:156:@29818.4]
  assign buffer_7_772 = $signed(_T_79403); // @[Modules.scala 63:156:@29819.4]
  assign _T_79405 = $signed(buffer_7_772) + $signed(buffer_7_724); // @[Modules.scala 63:156:@29821.4]
  assign _T_79406 = _T_79405[10:0]; // @[Modules.scala 63:156:@29822.4]
  assign buffer_7_773 = $signed(_T_79406); // @[Modules.scala 63:156:@29823.4]
  assign _T_79408 = $signed(buffer_7_773) + $signed(buffer_7_725); // @[Modules.scala 63:156:@29825.4]
  assign _T_79409 = _T_79408[10:0]; // @[Modules.scala 63:156:@29826.4]
  assign buffer_7_774 = $signed(_T_79409); // @[Modules.scala 63:156:@29827.4]
  assign _T_79411 = $signed(buffer_7_774) + $signed(buffer_7_726); // @[Modules.scala 63:156:@29829.4]
  assign _T_79412 = _T_79411[10:0]; // @[Modules.scala 63:156:@29830.4]
  assign buffer_7_775 = $signed(_T_79412); // @[Modules.scala 63:156:@29831.4]
  assign _T_79414 = $signed(buffer_7_775) + $signed(buffer_7_727); // @[Modules.scala 63:156:@29833.4]
  assign _T_79415 = _T_79414[10:0]; // @[Modules.scala 63:156:@29834.4]
  assign buffer_7_776 = $signed(_T_79415); // @[Modules.scala 63:156:@29835.4]
  assign _T_79417 = $signed(buffer_7_776) + $signed(buffer_7_728); // @[Modules.scala 63:156:@29837.4]
  assign _T_79418 = _T_79417[10:0]; // @[Modules.scala 63:156:@29838.4]
  assign buffer_7_777 = $signed(_T_79418); // @[Modules.scala 63:156:@29839.4]
  assign _T_79420 = $signed(buffer_7_777) + $signed(buffer_7_729); // @[Modules.scala 63:156:@29841.4]
  assign _T_79421 = _T_79420[10:0]; // @[Modules.scala 63:156:@29842.4]
  assign buffer_7_778 = $signed(_T_79421); // @[Modules.scala 63:156:@29843.4]
  assign _T_79423 = $signed(buffer_7_778) + $signed(buffer_2_730); // @[Modules.scala 63:156:@29845.4]
  assign _T_79424 = _T_79423[10:0]; // @[Modules.scala 63:156:@29846.4]
  assign buffer_7_779 = $signed(_T_79424); // @[Modules.scala 63:156:@29847.4]
  assign _T_79426 = $signed(buffer_7_779) + $signed(buffer_7_731); // @[Modules.scala 63:156:@29849.4]
  assign _T_79427 = _T_79426[10:0]; // @[Modules.scala 63:156:@29850.4]
  assign buffer_7_780 = $signed(_T_79427); // @[Modules.scala 63:156:@29851.4]
  assign _T_79429 = $signed(buffer_7_780) + $signed(buffer_4_732); // @[Modules.scala 63:156:@29853.4]
  assign _T_79430 = _T_79429[10:0]; // @[Modules.scala 63:156:@29854.4]
  assign buffer_7_781 = $signed(_T_79430); // @[Modules.scala 63:156:@29855.4]
  assign _T_79432 = $signed(buffer_7_781) + $signed(buffer_7_733); // @[Modules.scala 63:156:@29857.4]
  assign _T_79433 = _T_79432[10:0]; // @[Modules.scala 63:156:@29858.4]
  assign buffer_7_782 = $signed(_T_79433); // @[Modules.scala 63:156:@29859.4]
  assign _T_79435 = $signed(buffer_7_782) + $signed(buffer_7_734); // @[Modules.scala 63:156:@29861.4]
  assign _T_79436 = _T_79435[10:0]; // @[Modules.scala 63:156:@29862.4]
  assign buffer_7_783 = $signed(_T_79436); // @[Modules.scala 63:156:@29863.4]
  assign _T_79763 = $signed(_T_60884) + $signed(io_in_111); // @[Modules.scala 43:47:@30206.4]
  assign _T_79764 = _T_79763[4:0]; // @[Modules.scala 43:47:@30207.4]
  assign _T_79765 = $signed(_T_79764); // @[Modules.scala 43:47:@30208.4]
  assign _T_79786 = $signed(_T_54597) + $signed(io_in_121); // @[Modules.scala 43:47:@30232.4]
  assign _T_79787 = _T_79786[4:0]; // @[Modules.scala 43:47:@30233.4]
  assign _T_79788 = $signed(_T_79787); // @[Modules.scala 43:47:@30234.4]
  assign _T_79793 = $signed(_T_54604) + $signed(io_in_123); // @[Modules.scala 43:47:@30239.4]
  assign _T_79794 = _T_79793[4:0]; // @[Modules.scala 43:47:@30240.4]
  assign _T_79795 = $signed(_T_79794); // @[Modules.scala 43:47:@30241.4]
  assign _T_79800 = $signed(_T_54611) + $signed(io_in_125); // @[Modules.scala 43:47:@30246.4]
  assign _T_79801 = _T_79800[4:0]; // @[Modules.scala 43:47:@30247.4]
  assign _T_79802 = $signed(_T_79801); // @[Modules.scala 43:47:@30248.4]
  assign _T_79838 = $signed(_T_70246) - $signed(io_in_137); // @[Modules.scala 46:47:@30285.4]
  assign _T_79839 = _T_79838[4:0]; // @[Modules.scala 46:47:@30286.4]
  assign _T_79840 = $signed(_T_79839); // @[Modules.scala 46:47:@30287.4]
  assign _T_79958 = $signed(io_in_192) - $signed(io_in_193); // @[Modules.scala 40:46:@30424.4]
  assign _T_79959 = _T_79958[4:0]; // @[Modules.scala 40:46:@30425.4]
  assign _T_79960 = $signed(_T_79959); // @[Modules.scala 40:46:@30426.4]
  assign _T_80042 = $signed(_T_54897) + $signed(io_in_225); // @[Modules.scala 43:47:@30515.4]
  assign _T_80043 = _T_80042[4:0]; // @[Modules.scala 43:47:@30516.4]
  assign _T_80044 = $signed(_T_80043); // @[Modules.scala 43:47:@30517.4]
  assign _T_80051 = $signed(io_in_230) - $signed(io_in_231); // @[Modules.scala 40:46:@30527.4]
  assign _T_80052 = _T_80051[4:0]; // @[Modules.scala 40:46:@30528.4]
  assign _T_80053 = $signed(_T_80052); // @[Modules.scala 40:46:@30529.4]
  assign _T_80068 = $signed(io_in_236) - $signed(io_in_237); // @[Modules.scala 40:46:@30545.4]
  assign _T_80069 = _T_80068[4:0]; // @[Modules.scala 40:46:@30546.4]
  assign _T_80070 = $signed(_T_80069); // @[Modules.scala 40:46:@30547.4]
  assign _T_80111 = $signed(io_in_254) - $signed(io_in_255); // @[Modules.scala 40:46:@30593.4]
  assign _T_80112 = _T_80111[4:0]; // @[Modules.scala 40:46:@30594.4]
  assign _T_80113 = $signed(_T_80112); // @[Modules.scala 40:46:@30595.4]
  assign _T_80114 = $signed(io_in_256) - $signed(io_in_257); // @[Modules.scala 40:46:@30597.4]
  assign _T_80115 = _T_80114[4:0]; // @[Modules.scala 40:46:@30598.4]
  assign _T_80116 = $signed(_T_80115); // @[Modules.scala 40:46:@30599.4]
  assign _T_80181 = $signed(io_in_282) - $signed(io_in_283); // @[Modules.scala 40:46:@30670.4]
  assign _T_80182 = _T_80181[4:0]; // @[Modules.scala 40:46:@30671.4]
  assign _T_80183 = $signed(_T_80182); // @[Modules.scala 40:46:@30672.4]
  assign _T_80417 = $signed(io_in_362) + $signed(io_in_363); // @[Modules.scala 37:46:@30917.4]
  assign _T_80418 = _T_80417[4:0]; // @[Modules.scala 37:46:@30918.4]
  assign _T_80419 = $signed(_T_80418); // @[Modules.scala 37:46:@30919.4]
  assign _T_80453 = $signed(io_in_378) - $signed(io_in_379); // @[Modules.scala 40:46:@30958.4]
  assign _T_80454 = _T_80453[4:0]; // @[Modules.scala 40:46:@30959.4]
  assign _T_80455 = $signed(_T_80454); // @[Modules.scala 40:46:@30960.4]
  assign _T_80470 = $signed(io_in_384) - $signed(io_in_385); // @[Modules.scala 40:46:@30976.4]
  assign _T_80471 = _T_80470[4:0]; // @[Modules.scala 40:46:@30977.4]
  assign _T_80472 = $signed(_T_80471); // @[Modules.scala 40:46:@30978.4]
  assign _T_80497 = $signed(io_in_394) + $signed(io_in_395); // @[Modules.scala 37:46:@31005.4]
  assign _T_80498 = _T_80497[4:0]; // @[Modules.scala 37:46:@31006.4]
  assign _T_80499 = $signed(_T_80498); // @[Modules.scala 37:46:@31007.4]
  assign _T_80522 = $signed(_T_64888) + $signed(io_in_409); // @[Modules.scala 43:47:@31036.4]
  assign _T_80523 = _T_80522[4:0]; // @[Modules.scala 43:47:@31037.4]
  assign _T_80524 = $signed(_T_80523); // @[Modules.scala 43:47:@31038.4]
  assign _T_80671 = $signed(_T_77469) + $signed(io_in_479); // @[Modules.scala 43:47:@31209.4]
  assign _T_80672 = _T_80671[4:0]; // @[Modules.scala 43:47:@31210.4]
  assign _T_80673 = $signed(_T_80672); // @[Modules.scala 43:47:@31211.4]
  assign _T_80710 = $signed(_T_55613) + $signed(io_in_497); // @[Modules.scala 43:47:@31254.4]
  assign _T_80711 = _T_80710[4:0]; // @[Modules.scala 43:47:@31255.4]
  assign _T_80712 = $signed(_T_80711); // @[Modules.scala 43:47:@31256.4]
  assign _T_80740 = $signed(_T_55651) + $signed(io_in_509); // @[Modules.scala 43:47:@31287.4]
  assign _T_80741 = _T_80740[4:0]; // @[Modules.scala 43:47:@31288.4]
  assign _T_80742 = $signed(_T_80741); // @[Modules.scala 43:47:@31289.4]
  assign _T_80890 = $signed(_T_55821) + $signed(io_in_569); // @[Modules.scala 43:47:@31452.4]
  assign _T_80891 = _T_80890[4:0]; // @[Modules.scala 43:47:@31453.4]
  assign _T_80892 = $signed(_T_80891); // @[Modules.scala 43:47:@31454.4]
  assign _T_80952 = $signed(_T_55903) + $signed(io_in_597); // @[Modules.scala 43:47:@31523.4]
  assign _T_80953 = _T_80952[4:0]; // @[Modules.scala 43:47:@31524.4]
  assign _T_80954 = $signed(_T_80953); // @[Modules.scala 43:47:@31525.4]
  assign _T_80987 = $signed(_T_62268) + $signed(io_in_607); // @[Modules.scala 43:47:@31558.4]
  assign _T_80988 = _T_80987[4:0]; // @[Modules.scala 43:47:@31559.4]
  assign _T_80989 = $signed(_T_80988); // @[Modules.scala 43:47:@31560.4]
  assign _T_81023 = $signed(_T_55970) + $signed(io_in_623); // @[Modules.scala 43:47:@31599.4]
  assign _T_81024 = _T_81023[4:0]; // @[Modules.scala 43:47:@31600.4]
  assign _T_81025 = $signed(_T_81024); // @[Modules.scala 43:47:@31601.4]
  assign _T_81095 = $signed(_T_56074) + $signed(io_in_655); // @[Modules.scala 43:47:@31681.4]
  assign _T_81096 = _T_81095[4:0]; // @[Modules.scala 43:47:@31682.4]
  assign _T_81097 = $signed(_T_81096); // @[Modules.scala 43:47:@31683.4]
  assign _T_81410 = $signed(_T_68617) - $signed(io_in_753); // @[Modules.scala 46:47:@32003.4]
  assign _T_81411 = _T_81410[4:0]; // @[Modules.scala 46:47:@32004.4]
  assign _T_81412 = $signed(_T_81411); // @[Modules.scala 46:47:@32005.4]
  assign _T_81427 = $signed(_T_56302) + $signed(io_in_759); // @[Modules.scala 43:47:@32021.4]
  assign _T_81428 = _T_81427[4:0]; // @[Modules.scala 43:47:@32022.4]
  assign _T_81429 = $signed(_T_81428); // @[Modules.scala 43:47:@32023.4]
  assign _T_81440 = $signed(io_in_764) - $signed(io_in_765); // @[Modules.scala 40:46:@32036.4]
  assign _T_81441 = _T_81440[4:0]; // @[Modules.scala 40:46:@32037.4]
  assign _T_81442 = $signed(_T_81441); // @[Modules.scala 40:46:@32038.4]
  assign _T_81504 = $signed(buffer_1_4) + $signed(buffer_2_5); // @[Modules.scala 50:57:@32105.4]
  assign _T_81505 = _T_81504[10:0]; // @[Modules.scala 50:57:@32106.4]
  assign buffer_8_394 = $signed(_T_81505); // @[Modules.scala 50:57:@32107.4]
  assign _T_81513 = $signed(buffer_0_10) + $signed(buffer_2_11); // @[Modules.scala 50:57:@32117.4]
  assign _T_81514 = _T_81513[10:0]; // @[Modules.scala 50:57:@32118.4]
  assign buffer_8_397 = $signed(_T_81514); // @[Modules.scala 50:57:@32119.4]
  assign _T_81519 = $signed(buffer_3_14) + $signed(buffer_0_15); // @[Modules.scala 50:57:@32125.4]
  assign _T_81520 = _T_81519[10:0]; // @[Modules.scala 50:57:@32126.4]
  assign buffer_8_399 = $signed(_T_81520); // @[Modules.scala 50:57:@32127.4]
  assign _T_81522 = $signed(buffer_2_16) + $signed(buffer_0_17); // @[Modules.scala 50:57:@32129.4]
  assign _T_81523 = _T_81522[10:0]; // @[Modules.scala 50:57:@32130.4]
  assign buffer_8_400 = $signed(_T_81523); // @[Modules.scala 50:57:@32131.4]
  assign _T_81564 = $signed(buffer_4_44) + $signed(buffer_3_45); // @[Modules.scala 50:57:@32185.4]
  assign _T_81565 = _T_81564[10:0]; // @[Modules.scala 50:57:@32186.4]
  assign buffer_8_414 = $signed(_T_81565); // @[Modules.scala 50:57:@32187.4]
  assign buffer_8_55 = {{6{_T_79765[4]}},_T_79765}; // @[Modules.scala 32:22:@8.4]
  assign _T_81579 = $signed(buffer_2_54) + $signed(buffer_8_55); // @[Modules.scala 50:57:@32205.4]
  assign _T_81580 = _T_81579[10:0]; // @[Modules.scala 50:57:@32206.4]
  assign buffer_8_419 = $signed(_T_81580); // @[Modules.scala 50:57:@32207.4]
  assign _T_81582 = $signed(buffer_1_56) + $signed(buffer_3_57); // @[Modules.scala 50:57:@32209.4]
  assign _T_81583 = _T_81582[10:0]; // @[Modules.scala 50:57:@32210.4]
  assign buffer_8_420 = $signed(_T_81583); // @[Modules.scala 50:57:@32211.4]
  assign buffer_8_60 = {{6{_T_79788[4]}},_T_79788}; // @[Modules.scala 32:22:@8.4]
  assign buffer_8_61 = {{6{_T_79795[4]}},_T_79795}; // @[Modules.scala 32:22:@8.4]
  assign _T_81588 = $signed(buffer_8_60) + $signed(buffer_8_61); // @[Modules.scala 50:57:@32217.4]
  assign _T_81589 = _T_81588[10:0]; // @[Modules.scala 50:57:@32218.4]
  assign buffer_8_422 = $signed(_T_81589); // @[Modules.scala 50:57:@32219.4]
  assign buffer_8_62 = {{6{_T_79802[4]}},_T_79802}; // @[Modules.scala 32:22:@8.4]
  assign _T_81591 = $signed(buffer_8_62) + $signed(buffer_7_63); // @[Modules.scala 50:57:@32221.4]
  assign _T_81592 = _T_81591[10:0]; // @[Modules.scala 50:57:@32222.4]
  assign buffer_8_423 = $signed(_T_81592); // @[Modules.scala 50:57:@32223.4]
  assign buffer_8_68 = {{6{_T_79840[4]}},_T_79840}; // @[Modules.scala 32:22:@8.4]
  assign _T_81600 = $signed(buffer_8_68) + $signed(buffer_0_69); // @[Modules.scala 50:57:@32233.4]
  assign _T_81601 = _T_81600[10:0]; // @[Modules.scala 50:57:@32234.4]
  assign buffer_8_426 = $signed(_T_81601); // @[Modules.scala 50:57:@32235.4]
  assign _T_81603 = $signed(buffer_0_70) + $signed(buffer_5_71); // @[Modules.scala 50:57:@32237.4]
  assign _T_81604 = _T_81603[10:0]; // @[Modules.scala 50:57:@32238.4]
  assign buffer_8_427 = $signed(_T_81604); // @[Modules.scala 50:57:@32239.4]
  assign _T_81621 = $signed(buffer_0_82) + $signed(buffer_6_83); // @[Modules.scala 50:57:@32261.4]
  assign _T_81622 = _T_81621[10:0]; // @[Modules.scala 50:57:@32262.4]
  assign buffer_8_433 = $signed(_T_81622); // @[Modules.scala 50:57:@32263.4]
  assign buffer_8_96 = {{6{_T_79960[4]}},_T_79960}; // @[Modules.scala 32:22:@8.4]
  assign _T_81642 = $signed(buffer_8_96) + $signed(buffer_6_97); // @[Modules.scala 50:57:@32289.4]
  assign _T_81643 = _T_81642[10:0]; // @[Modules.scala 50:57:@32290.4]
  assign buffer_8_440 = $signed(_T_81643); // @[Modules.scala 50:57:@32291.4]
  assign _T_81651 = $signed(buffer_6_102) + $signed(buffer_1_103); // @[Modules.scala 50:57:@32301.4]
  assign _T_81652 = _T_81651[10:0]; // @[Modules.scala 50:57:@32302.4]
  assign buffer_8_443 = $signed(_T_81652); // @[Modules.scala 50:57:@32303.4]
  assign _T_81657 = $signed(buffer_4_106) + $signed(buffer_1_107); // @[Modules.scala 50:57:@32309.4]
  assign _T_81658 = _T_81657[10:0]; // @[Modules.scala 50:57:@32310.4]
  assign buffer_8_445 = $signed(_T_81658); // @[Modules.scala 50:57:@32311.4]
  assign buffer_8_112 = {{6{_T_80044[4]}},_T_80044}; // @[Modules.scala 32:22:@8.4]
  assign _T_81666 = $signed(buffer_8_112) + $signed(buffer_3_113); // @[Modules.scala 50:57:@32321.4]
  assign _T_81667 = _T_81666[10:0]; // @[Modules.scala 50:57:@32322.4]
  assign buffer_8_448 = $signed(_T_81667); // @[Modules.scala 50:57:@32323.4]
  assign buffer_8_115 = {{6{_T_80053[4]}},_T_80053}; // @[Modules.scala 32:22:@8.4]
  assign _T_81669 = $signed(buffer_3_114) + $signed(buffer_8_115); // @[Modules.scala 50:57:@32325.4]
  assign _T_81670 = _T_81669[10:0]; // @[Modules.scala 50:57:@32326.4]
  assign buffer_8_449 = $signed(_T_81670); // @[Modules.scala 50:57:@32327.4]
  assign buffer_8_118 = {{6{_T_80070[4]}},_T_80070}; // @[Modules.scala 32:22:@8.4]
  assign _T_81675 = $signed(buffer_8_118) + $signed(buffer_0_119); // @[Modules.scala 50:57:@32333.4]
  assign _T_81676 = _T_81675[10:0]; // @[Modules.scala 50:57:@32334.4]
  assign buffer_8_451 = $signed(_T_81676); // @[Modules.scala 50:57:@32335.4]
  assign _T_81678 = $signed(buffer_0_120) + $signed(buffer_3_121); // @[Modules.scala 50:57:@32337.4]
  assign _T_81679 = _T_81678[10:0]; // @[Modules.scala 50:57:@32338.4]
  assign buffer_8_452 = $signed(_T_81679); // @[Modules.scala 50:57:@32339.4]
  assign _T_81681 = $signed(buffer_4_122) + $signed(buffer_6_123); // @[Modules.scala 50:57:@32341.4]
  assign _T_81682 = _T_81681[10:0]; // @[Modules.scala 50:57:@32342.4]
  assign buffer_8_453 = $signed(_T_81682); // @[Modules.scala 50:57:@32343.4]
  assign buffer_8_127 = {{6{_T_80113[4]}},_T_80113}; // @[Modules.scala 32:22:@8.4]
  assign _T_81687 = $signed(buffer_5_126) + $signed(buffer_8_127); // @[Modules.scala 50:57:@32349.4]
  assign _T_81688 = _T_81687[10:0]; // @[Modules.scala 50:57:@32350.4]
  assign buffer_8_455 = $signed(_T_81688); // @[Modules.scala 50:57:@32351.4]
  assign buffer_8_128 = {{6{_T_80116[4]}},_T_80116}; // @[Modules.scala 32:22:@8.4]
  assign _T_81690 = $signed(buffer_8_128) + $signed(buffer_0_129); // @[Modules.scala 50:57:@32353.4]
  assign _T_81691 = _T_81690[10:0]; // @[Modules.scala 50:57:@32354.4]
  assign buffer_8_456 = $signed(_T_81691); // @[Modules.scala 50:57:@32355.4]
  assign _T_81693 = $signed(buffer_0_130) + $signed(buffer_1_131); // @[Modules.scala 50:57:@32357.4]
  assign _T_81694 = _T_81693[10:0]; // @[Modules.scala 50:57:@32358.4]
  assign buffer_8_457 = $signed(_T_81694); // @[Modules.scala 50:57:@32359.4]
  assign _T_81702 = $signed(buffer_3_136) + $signed(buffer_5_137); // @[Modules.scala 50:57:@32369.4]
  assign _T_81703 = _T_81702[10:0]; // @[Modules.scala 50:57:@32370.4]
  assign buffer_8_460 = $signed(_T_81703); // @[Modules.scala 50:57:@32371.4]
  assign buffer_8_141 = {{6{_T_80183[4]}},_T_80183}; // @[Modules.scala 32:22:@8.4]
  assign _T_81708 = $signed(buffer_5_140) + $signed(buffer_8_141); // @[Modules.scala 50:57:@32377.4]
  assign _T_81709 = _T_81708[10:0]; // @[Modules.scala 50:57:@32378.4]
  assign buffer_8_462 = $signed(_T_81709); // @[Modules.scala 50:57:@32379.4]
  assign _T_81729 = $signed(buffer_4_154) + $signed(buffer_3_155); // @[Modules.scala 50:57:@32405.4]
  assign _T_81730 = _T_81729[10:0]; // @[Modules.scala 50:57:@32406.4]
  assign buffer_8_469 = $signed(_T_81730); // @[Modules.scala 50:57:@32407.4]
  assign _T_81741 = $signed(buffer_6_162) + $signed(buffer_0_163); // @[Modules.scala 50:57:@32421.4]
  assign _T_81742 = _T_81741[10:0]; // @[Modules.scala 50:57:@32422.4]
  assign buffer_8_473 = $signed(_T_81742); // @[Modules.scala 50:57:@32423.4]
  assign _T_81750 = $signed(buffer_0_168) + $signed(buffer_5_169); // @[Modules.scala 50:57:@32433.4]
  assign _T_81751 = _T_81750[10:0]; // @[Modules.scala 50:57:@32434.4]
  assign buffer_8_476 = $signed(_T_81751); // @[Modules.scala 50:57:@32435.4]
  assign _T_81762 = $signed(buffer_1_176) + $signed(buffer_5_177); // @[Modules.scala 50:57:@32449.4]
  assign _T_81763 = _T_81762[10:0]; // @[Modules.scala 50:57:@32450.4]
  assign buffer_8_480 = $signed(_T_81763); // @[Modules.scala 50:57:@32451.4]
  assign buffer_8_181 = {{6{_T_80419[4]}},_T_80419}; // @[Modules.scala 32:22:@8.4]
  assign _T_81768 = $signed(buffer_0_180) + $signed(buffer_8_181); // @[Modules.scala 50:57:@32457.4]
  assign _T_81769 = _T_81768[10:0]; // @[Modules.scala 50:57:@32458.4]
  assign buffer_8_482 = $signed(_T_81769); // @[Modules.scala 50:57:@32459.4]
  assign buffer_8_189 = {{6{_T_80455[4]}},_T_80455}; // @[Modules.scala 32:22:@8.4]
  assign _T_81780 = $signed(buffer_0_188) + $signed(buffer_8_189); // @[Modules.scala 50:57:@32473.4]
  assign _T_81781 = _T_81780[10:0]; // @[Modules.scala 50:57:@32474.4]
  assign buffer_8_486 = $signed(_T_81781); // @[Modules.scala 50:57:@32475.4]
  assign buffer_8_192 = {{6{_T_80472[4]}},_T_80472}; // @[Modules.scala 32:22:@8.4]
  assign _T_81786 = $signed(buffer_8_192) + $signed(buffer_2_193); // @[Modules.scala 50:57:@32481.4]
  assign _T_81787 = _T_81786[10:0]; // @[Modules.scala 50:57:@32482.4]
  assign buffer_8_488 = $signed(_T_81787); // @[Modules.scala 50:57:@32483.4]
  assign buffer_8_197 = {{6{_T_80499[4]}},_T_80499}; // @[Modules.scala 32:22:@8.4]
  assign _T_81792 = $signed(buffer_6_196) + $signed(buffer_8_197); // @[Modules.scala 50:57:@32489.4]
  assign _T_81793 = _T_81792[10:0]; // @[Modules.scala 50:57:@32490.4]
  assign buffer_8_490 = $signed(_T_81793); // @[Modules.scala 50:57:@32491.4]
  assign _T_81798 = $signed(buffer_0_200) + $signed(buffer_3_201); // @[Modules.scala 50:57:@32497.4]
  assign _T_81799 = _T_81798[10:0]; // @[Modules.scala 50:57:@32498.4]
  assign buffer_8_492 = $signed(_T_81799); // @[Modules.scala 50:57:@32499.4]
  assign buffer_8_204 = {{6{_T_80524[4]}},_T_80524}; // @[Modules.scala 32:22:@8.4]
  assign _T_81804 = $signed(buffer_8_204) + $signed(buffer_0_205); // @[Modules.scala 50:57:@32505.4]
  assign _T_81805 = _T_81804[10:0]; // @[Modules.scala 50:57:@32506.4]
  assign buffer_8_494 = $signed(_T_81805); // @[Modules.scala 50:57:@32507.4]
  assign _T_81807 = $signed(buffer_4_206) + $signed(buffer_3_207); // @[Modules.scala 50:57:@32509.4]
  assign _T_81808 = _T_81807[10:0]; // @[Modules.scala 50:57:@32510.4]
  assign buffer_8_495 = $signed(_T_81808); // @[Modules.scala 50:57:@32511.4]
  assign _T_81828 = $signed(buffer_2_220) + $signed(buffer_6_221); // @[Modules.scala 50:57:@32537.4]
  assign _T_81829 = _T_81828[10:0]; // @[Modules.scala 50:57:@32538.4]
  assign buffer_8_502 = $signed(_T_81829); // @[Modules.scala 50:57:@32539.4]
  assign _T_81831 = $signed(buffer_0_222) + $signed(buffer_3_223); // @[Modules.scala 50:57:@32541.4]
  assign _T_81832 = _T_81831[10:0]; // @[Modules.scala 50:57:@32542.4]
  assign buffer_8_503 = $signed(_T_81832); // @[Modules.scala 50:57:@32543.4]
  assign _T_81834 = $signed(buffer_3_224) + $signed(buffer_7_225); // @[Modules.scala 50:57:@32545.4]
  assign _T_81835 = _T_81834[10:0]; // @[Modules.scala 50:57:@32546.4]
  assign buffer_8_504 = $signed(_T_81835); // @[Modules.scala 50:57:@32547.4]
  assign buffer_8_239 = {{6{_T_80673[4]}},_T_80673}; // @[Modules.scala 32:22:@8.4]
  assign _T_81855 = $signed(buffer_2_238) + $signed(buffer_8_239); // @[Modules.scala 50:57:@32573.4]
  assign _T_81856 = _T_81855[10:0]; // @[Modules.scala 50:57:@32574.4]
  assign buffer_8_511 = $signed(_T_81856); // @[Modules.scala 50:57:@32575.4]
  assign _T_81867 = $signed(buffer_4_246) + $signed(buffer_7_247); // @[Modules.scala 50:57:@32589.4]
  assign _T_81868 = _T_81867[10:0]; // @[Modules.scala 50:57:@32590.4]
  assign buffer_8_515 = $signed(_T_81868); // @[Modules.scala 50:57:@32591.4]
  assign buffer_8_248 = {{6{_T_80712[4]}},_T_80712}; // @[Modules.scala 32:22:@8.4]
  assign _T_81870 = $signed(buffer_8_248) + $signed(buffer_0_249); // @[Modules.scala 50:57:@32593.4]
  assign _T_81871 = _T_81870[10:0]; // @[Modules.scala 50:57:@32594.4]
  assign buffer_8_516 = $signed(_T_81871); // @[Modules.scala 50:57:@32595.4]
  assign _T_81876 = $signed(buffer_1_252) + $signed(buffer_0_253); // @[Modules.scala 50:57:@32601.4]
  assign _T_81877 = _T_81876[10:0]; // @[Modules.scala 50:57:@32602.4]
  assign buffer_8_518 = $signed(_T_81877); // @[Modules.scala 50:57:@32603.4]
  assign buffer_8_254 = {{6{_T_80742[4]}},_T_80742}; // @[Modules.scala 32:22:@8.4]
  assign _T_81879 = $signed(buffer_8_254) + $signed(buffer_1_255); // @[Modules.scala 50:57:@32605.4]
  assign _T_81880 = _T_81879[10:0]; // @[Modules.scala 50:57:@32606.4]
  assign buffer_8_519 = $signed(_T_81880); // @[Modules.scala 50:57:@32607.4]
  assign _T_81897 = $signed(buffer_2_266) + $signed(buffer_1_267); // @[Modules.scala 50:57:@32629.4]
  assign _T_81898 = _T_81897[10:0]; // @[Modules.scala 50:57:@32630.4]
  assign buffer_8_525 = $signed(_T_81898); // @[Modules.scala 50:57:@32631.4]
  assign _T_81900 = $signed(buffer_1_268) + $signed(buffer_7_269); // @[Modules.scala 50:57:@32633.4]
  assign _T_81901 = _T_81900[10:0]; // @[Modules.scala 50:57:@32634.4]
  assign buffer_8_526 = $signed(_T_81901); // @[Modules.scala 50:57:@32635.4]
  assign _T_81906 = $signed(buffer_2_272) + $signed(buffer_3_273); // @[Modules.scala 50:57:@32641.4]
  assign _T_81907 = _T_81906[10:0]; // @[Modules.scala 50:57:@32642.4]
  assign buffer_8_528 = $signed(_T_81907); // @[Modules.scala 50:57:@32643.4]
  assign _T_81912 = $signed(buffer_7_276) + $signed(buffer_5_277); // @[Modules.scala 50:57:@32649.4]
  assign _T_81913 = _T_81912[10:0]; // @[Modules.scala 50:57:@32650.4]
  assign buffer_8_530 = $signed(_T_81913); // @[Modules.scala 50:57:@32651.4]
  assign _T_81918 = $signed(buffer_0_280) + $signed(buffer_1_281); // @[Modules.scala 50:57:@32657.4]
  assign _T_81919 = _T_81918[10:0]; // @[Modules.scala 50:57:@32658.4]
  assign buffer_8_532 = $signed(_T_81919); // @[Modules.scala 50:57:@32659.4]
  assign _T_81921 = $signed(buffer_5_282) + $signed(buffer_1_283); // @[Modules.scala 50:57:@32661.4]
  assign _T_81922 = _T_81921[10:0]; // @[Modules.scala 50:57:@32662.4]
  assign buffer_8_533 = $signed(_T_81922); // @[Modules.scala 50:57:@32663.4]
  assign buffer_8_284 = {{6{_T_80892[4]}},_T_80892}; // @[Modules.scala 32:22:@8.4]
  assign _T_81924 = $signed(buffer_8_284) + $signed(buffer_5_285); // @[Modules.scala 50:57:@32665.4]
  assign _T_81925 = _T_81924[10:0]; // @[Modules.scala 50:57:@32666.4]
  assign buffer_8_534 = $signed(_T_81925); // @[Modules.scala 50:57:@32667.4]
  assign _T_81936 = $signed(buffer_0_292) + $signed(buffer_7_293); // @[Modules.scala 50:57:@32681.4]
  assign _T_81937 = _T_81936[10:0]; // @[Modules.scala 50:57:@32682.4]
  assign buffer_8_538 = $signed(_T_81937); // @[Modules.scala 50:57:@32683.4]
  assign buffer_8_298 = {{6{_T_80954[4]}},_T_80954}; // @[Modules.scala 32:22:@8.4]
  assign _T_81945 = $signed(buffer_8_298) + $signed(buffer_0_299); // @[Modules.scala 50:57:@32693.4]
  assign _T_81946 = _T_81945[10:0]; // @[Modules.scala 50:57:@32694.4]
  assign buffer_8_541 = $signed(_T_81946); // @[Modules.scala 50:57:@32695.4]
  assign _T_81948 = $signed(buffer_5_300) + $signed(buffer_7_301); // @[Modules.scala 50:57:@32697.4]
  assign _T_81949 = _T_81948[10:0]; // @[Modules.scala 50:57:@32698.4]
  assign buffer_8_542 = $signed(_T_81949); // @[Modules.scala 50:57:@32699.4]
  assign buffer_8_303 = {{6{_T_80989[4]}},_T_80989}; // @[Modules.scala 32:22:@8.4]
  assign _T_81951 = $signed(buffer_6_302) + $signed(buffer_8_303); // @[Modules.scala 50:57:@32701.4]
  assign _T_81952 = _T_81951[10:0]; // @[Modules.scala 50:57:@32702.4]
  assign buffer_8_543 = $signed(_T_81952); // @[Modules.scala 50:57:@32703.4]
  assign buffer_8_311 = {{6{_T_81025[4]}},_T_81025}; // @[Modules.scala 32:22:@8.4]
  assign _T_81963 = $signed(buffer_3_310) + $signed(buffer_8_311); // @[Modules.scala 50:57:@32717.4]
  assign _T_81964 = _T_81963[10:0]; // @[Modules.scala 50:57:@32718.4]
  assign buffer_8_547 = $signed(_T_81964); // @[Modules.scala 50:57:@32719.4]
  assign _T_81966 = $signed(buffer_1_312) + $signed(buffer_0_313); // @[Modules.scala 50:57:@32721.4]
  assign _T_81967 = _T_81966[10:0]; // @[Modules.scala 50:57:@32722.4]
  assign buffer_8_548 = $signed(_T_81967); // @[Modules.scala 50:57:@32723.4]
  assign _T_81969 = $signed(buffer_0_314) + $signed(buffer_6_315); // @[Modules.scala 50:57:@32725.4]
  assign _T_81970 = _T_81969[10:0]; // @[Modules.scala 50:57:@32726.4]
  assign buffer_8_549 = $signed(_T_81970); // @[Modules.scala 50:57:@32727.4]
  assign _T_81984 = $signed(buffer_1_324) + $signed(buffer_2_325); // @[Modules.scala 50:57:@32745.4]
  assign _T_81985 = _T_81984[10:0]; // @[Modules.scala 50:57:@32746.4]
  assign buffer_8_554 = $signed(_T_81985); // @[Modules.scala 50:57:@32747.4]
  assign buffer_8_327 = {{6{_T_81097[4]}},_T_81097}; // @[Modules.scala 32:22:@8.4]
  assign _T_81987 = $signed(buffer_3_326) + $signed(buffer_8_327); // @[Modules.scala 50:57:@32749.4]
  assign _T_81988 = _T_81987[10:0]; // @[Modules.scala 50:57:@32750.4]
  assign buffer_8_555 = $signed(_T_81988); // @[Modules.scala 50:57:@32751.4]
  assign _T_81993 = $signed(buffer_4_330) + $signed(buffer_0_331); // @[Modules.scala 50:57:@32757.4]
  assign _T_81994 = _T_81993[10:0]; // @[Modules.scala 50:57:@32758.4]
  assign buffer_8_557 = $signed(_T_81994); // @[Modules.scala 50:57:@32759.4]
  assign _T_81999 = $signed(buffer_4_334) + $signed(buffer_3_335); // @[Modules.scala 50:57:@32765.4]
  assign _T_82000 = _T_81999[10:0]; // @[Modules.scala 50:57:@32766.4]
  assign buffer_8_559 = $signed(_T_82000); // @[Modules.scala 50:57:@32767.4]
  assign _T_82005 = $signed(buffer_4_338) + $signed(buffer_2_339); // @[Modules.scala 50:57:@32773.4]
  assign _T_82006 = _T_82005[10:0]; // @[Modules.scala 50:57:@32774.4]
  assign buffer_8_561 = $signed(_T_82006); // @[Modules.scala 50:57:@32775.4]
  assign _T_82023 = $signed(buffer_5_350) + $signed(buffer_3_351); // @[Modules.scala 50:57:@32797.4]
  assign _T_82024 = _T_82023[10:0]; // @[Modules.scala 50:57:@32798.4]
  assign buffer_8_567 = $signed(_T_82024); // @[Modules.scala 50:57:@32799.4]
  assign buffer_8_376 = {{6{_T_81412[4]}},_T_81412}; // @[Modules.scala 32:22:@8.4]
  assign _T_82062 = $signed(buffer_8_376) + $signed(buffer_3_377); // @[Modules.scala 50:57:@32849.4]
  assign _T_82063 = _T_82062[10:0]; // @[Modules.scala 50:57:@32850.4]
  assign buffer_8_580 = $signed(_T_82063); // @[Modules.scala 50:57:@32851.4]
  assign buffer_8_379 = {{6{_T_81429[4]}},_T_81429}; // @[Modules.scala 32:22:@8.4]
  assign _T_82065 = $signed(buffer_1_378) + $signed(buffer_8_379); // @[Modules.scala 50:57:@32853.4]
  assign _T_82066 = _T_82065[10:0]; // @[Modules.scala 50:57:@32854.4]
  assign buffer_8_581 = $signed(_T_82066); // @[Modules.scala 50:57:@32855.4]
  assign buffer_8_382 = {{6{_T_81442[4]}},_T_81442}; // @[Modules.scala 32:22:@8.4]
  assign _T_82071 = $signed(buffer_8_382) + $signed(buffer_0_383); // @[Modules.scala 50:57:@32861.4]
  assign _T_82072 = _T_82071[10:0]; // @[Modules.scala 50:57:@32862.4]
  assign buffer_8_583 = $signed(_T_82072); // @[Modules.scala 50:57:@32863.4]
  assign _T_82080 = $signed(buffer_1_388) + $signed(buffer_5_389); // @[Modules.scala 50:57:@32873.4]
  assign _T_82081 = _T_82080[10:0]; // @[Modules.scala 50:57:@32874.4]
  assign buffer_8_586 = $signed(_T_82081); // @[Modules.scala 50:57:@32875.4]
  assign _T_82089 = $signed(buffer_8_394) + $signed(buffer_4_395); // @[Modules.scala 53:83:@32885.4]
  assign _T_82090 = _T_82089[10:0]; // @[Modules.scala 53:83:@32886.4]
  assign buffer_8_589 = $signed(_T_82090); // @[Modules.scala 53:83:@32887.4]
  assign _T_82092 = $signed(buffer_3_396) + $signed(buffer_8_397); // @[Modules.scala 53:83:@32889.4]
  assign _T_82093 = _T_82092[10:0]; // @[Modules.scala 53:83:@32890.4]
  assign buffer_8_590 = $signed(_T_82093); // @[Modules.scala 53:83:@32891.4]
  assign _T_82095 = $signed(buffer_3_398) + $signed(buffer_8_399); // @[Modules.scala 53:83:@32893.4]
  assign _T_82096 = _T_82095[10:0]; // @[Modules.scala 53:83:@32894.4]
  assign buffer_8_591 = $signed(_T_82096); // @[Modules.scala 53:83:@32895.4]
  assign _T_82098 = $signed(buffer_8_400) + $signed(buffer_0_401); // @[Modules.scala 53:83:@32897.4]
  assign _T_82099 = _T_82098[10:0]; // @[Modules.scala 53:83:@32898.4]
  assign buffer_8_592 = $signed(_T_82099); // @[Modules.scala 53:83:@32899.4]
  assign _T_82104 = $signed(buffer_0_404) + $signed(buffer_7_405); // @[Modules.scala 53:83:@32905.4]
  assign _T_82105 = _T_82104[10:0]; // @[Modules.scala 53:83:@32906.4]
  assign buffer_8_594 = $signed(_T_82105); // @[Modules.scala 53:83:@32907.4]
  assign _T_82116 = $signed(buffer_0_412) + $signed(buffer_6_413); // @[Modules.scala 53:83:@32921.4]
  assign _T_82117 = _T_82116[10:0]; // @[Modules.scala 53:83:@32922.4]
  assign buffer_8_598 = $signed(_T_82117); // @[Modules.scala 53:83:@32923.4]
  assign _T_82119 = $signed(buffer_8_414) + $signed(buffer_6_415); // @[Modules.scala 53:83:@32925.4]
  assign _T_82120 = _T_82119[10:0]; // @[Modules.scala 53:83:@32926.4]
  assign buffer_8_599 = $signed(_T_82120); // @[Modules.scala 53:83:@32927.4]
  assign _T_82125 = $signed(buffer_3_418) + $signed(buffer_8_419); // @[Modules.scala 53:83:@32933.4]
  assign _T_82126 = _T_82125[10:0]; // @[Modules.scala 53:83:@32934.4]
  assign buffer_8_601 = $signed(_T_82126); // @[Modules.scala 53:83:@32935.4]
  assign _T_82128 = $signed(buffer_8_420) + $signed(buffer_5_421); // @[Modules.scala 53:83:@32937.4]
  assign _T_82129 = _T_82128[10:0]; // @[Modules.scala 53:83:@32938.4]
  assign buffer_8_602 = $signed(_T_82129); // @[Modules.scala 53:83:@32939.4]
  assign _T_82131 = $signed(buffer_8_422) + $signed(buffer_8_423); // @[Modules.scala 53:83:@32941.4]
  assign _T_82132 = _T_82131[10:0]; // @[Modules.scala 53:83:@32942.4]
  assign buffer_8_603 = $signed(_T_82132); // @[Modules.scala 53:83:@32943.4]
  assign _T_82134 = $signed(buffer_6_424) + $signed(buffer_4_425); // @[Modules.scala 53:83:@32945.4]
  assign _T_82135 = _T_82134[10:0]; // @[Modules.scala 53:83:@32946.4]
  assign buffer_8_604 = $signed(_T_82135); // @[Modules.scala 53:83:@32947.4]
  assign _T_82137 = $signed(buffer_8_426) + $signed(buffer_8_427); // @[Modules.scala 53:83:@32949.4]
  assign _T_82138 = _T_82137[10:0]; // @[Modules.scala 53:83:@32950.4]
  assign buffer_8_605 = $signed(_T_82138); // @[Modules.scala 53:83:@32951.4]
  assign _T_82146 = $signed(buffer_1_432) + $signed(buffer_8_433); // @[Modules.scala 53:83:@32961.4]
  assign _T_82147 = _T_82146[10:0]; // @[Modules.scala 53:83:@32962.4]
  assign buffer_8_608 = $signed(_T_82147); // @[Modules.scala 53:83:@32963.4]
  assign _T_82152 = $signed(buffer_3_436) + $signed(buffer_0_437); // @[Modules.scala 53:83:@32969.4]
  assign _T_82153 = _T_82152[10:0]; // @[Modules.scala 53:83:@32970.4]
  assign buffer_8_610 = $signed(_T_82153); // @[Modules.scala 53:83:@32971.4]
  assign _T_82155 = $signed(buffer_2_438) + $signed(buffer_4_439); // @[Modules.scala 53:83:@32973.4]
  assign _T_82156 = _T_82155[10:0]; // @[Modules.scala 53:83:@32974.4]
  assign buffer_8_611 = $signed(_T_82156); // @[Modules.scala 53:83:@32975.4]
  assign _T_82158 = $signed(buffer_8_440) + $signed(buffer_3_441); // @[Modules.scala 53:83:@32977.4]
  assign _T_82159 = _T_82158[10:0]; // @[Modules.scala 53:83:@32978.4]
  assign buffer_8_612 = $signed(_T_82159); // @[Modules.scala 53:83:@32979.4]
  assign _T_82161 = $signed(buffer_3_442) + $signed(buffer_8_443); // @[Modules.scala 53:83:@32981.4]
  assign _T_82162 = _T_82161[10:0]; // @[Modules.scala 53:83:@32982.4]
  assign buffer_8_613 = $signed(_T_82162); // @[Modules.scala 53:83:@32983.4]
  assign _T_82164 = $signed(buffer_4_444) + $signed(buffer_8_445); // @[Modules.scala 53:83:@32985.4]
  assign _T_82165 = _T_82164[10:0]; // @[Modules.scala 53:83:@32986.4]
  assign buffer_8_614 = $signed(_T_82165); // @[Modules.scala 53:83:@32987.4]
  assign _T_82167 = $signed(buffer_2_446) + $signed(buffer_0_447); // @[Modules.scala 53:83:@32989.4]
  assign _T_82168 = _T_82167[10:0]; // @[Modules.scala 53:83:@32990.4]
  assign buffer_8_615 = $signed(_T_82168); // @[Modules.scala 53:83:@32991.4]
  assign _T_82170 = $signed(buffer_8_448) + $signed(buffer_8_449); // @[Modules.scala 53:83:@32993.4]
  assign _T_82171 = _T_82170[10:0]; // @[Modules.scala 53:83:@32994.4]
  assign buffer_8_616 = $signed(_T_82171); // @[Modules.scala 53:83:@32995.4]
  assign _T_82173 = $signed(buffer_0_450) + $signed(buffer_8_451); // @[Modules.scala 53:83:@32997.4]
  assign _T_82174 = _T_82173[10:0]; // @[Modules.scala 53:83:@32998.4]
  assign buffer_8_617 = $signed(_T_82174); // @[Modules.scala 53:83:@32999.4]
  assign _T_82176 = $signed(buffer_8_452) + $signed(buffer_8_453); // @[Modules.scala 53:83:@33001.4]
  assign _T_82177 = _T_82176[10:0]; // @[Modules.scala 53:83:@33002.4]
  assign buffer_8_618 = $signed(_T_82177); // @[Modules.scala 53:83:@33003.4]
  assign _T_82179 = $signed(buffer_0_454) + $signed(buffer_8_455); // @[Modules.scala 53:83:@33005.4]
  assign _T_82180 = _T_82179[10:0]; // @[Modules.scala 53:83:@33006.4]
  assign buffer_8_619 = $signed(_T_82180); // @[Modules.scala 53:83:@33007.4]
  assign _T_82182 = $signed(buffer_8_456) + $signed(buffer_8_457); // @[Modules.scala 53:83:@33009.4]
  assign _T_82183 = _T_82182[10:0]; // @[Modules.scala 53:83:@33010.4]
  assign buffer_8_620 = $signed(_T_82183); // @[Modules.scala 53:83:@33011.4]
  assign _T_82185 = $signed(buffer_0_458) + $signed(buffer_5_459); // @[Modules.scala 53:83:@33013.4]
  assign _T_82186 = _T_82185[10:0]; // @[Modules.scala 53:83:@33014.4]
  assign buffer_8_621 = $signed(_T_82186); // @[Modules.scala 53:83:@33015.4]
  assign _T_82188 = $signed(buffer_8_460) + $signed(buffer_0_461); // @[Modules.scala 53:83:@33017.4]
  assign _T_82189 = _T_82188[10:0]; // @[Modules.scala 53:83:@33018.4]
  assign buffer_8_622 = $signed(_T_82189); // @[Modules.scala 53:83:@33019.4]
  assign _T_82191 = $signed(buffer_8_462) + $signed(buffer_0_463); // @[Modules.scala 53:83:@33021.4]
  assign _T_82192 = _T_82191[10:0]; // @[Modules.scala 53:83:@33022.4]
  assign buffer_8_623 = $signed(_T_82192); // @[Modules.scala 53:83:@33023.4]
  assign _T_82197 = $signed(buffer_3_466) + $signed(buffer_0_467); // @[Modules.scala 53:83:@33029.4]
  assign _T_82198 = _T_82197[10:0]; // @[Modules.scala 53:83:@33030.4]
  assign buffer_8_625 = $signed(_T_82198); // @[Modules.scala 53:83:@33031.4]
  assign _T_82200 = $signed(buffer_5_468) + $signed(buffer_8_469); // @[Modules.scala 53:83:@33033.4]
  assign _T_82201 = _T_82200[10:0]; // @[Modules.scala 53:83:@33034.4]
  assign buffer_8_626 = $signed(_T_82201); // @[Modules.scala 53:83:@33035.4]
  assign _T_82206 = $signed(buffer_5_472) + $signed(buffer_8_473); // @[Modules.scala 53:83:@33041.4]
  assign _T_82207 = _T_82206[10:0]; // @[Modules.scala 53:83:@33042.4]
  assign buffer_8_628 = $signed(_T_82207); // @[Modules.scala 53:83:@33043.4]
  assign _T_82209 = $signed(buffer_2_474) + $signed(buffer_0_475); // @[Modules.scala 53:83:@33045.4]
  assign _T_82210 = _T_82209[10:0]; // @[Modules.scala 53:83:@33046.4]
  assign buffer_8_629 = $signed(_T_82210); // @[Modules.scala 53:83:@33047.4]
  assign _T_82212 = $signed(buffer_8_476) + $signed(buffer_3_477); // @[Modules.scala 53:83:@33049.4]
  assign _T_82213 = _T_82212[10:0]; // @[Modules.scala 53:83:@33050.4]
  assign buffer_8_630 = $signed(_T_82213); // @[Modules.scala 53:83:@33051.4]
  assign _T_82218 = $signed(buffer_8_480) + $signed(buffer_5_481); // @[Modules.scala 53:83:@33057.4]
  assign _T_82219 = _T_82218[10:0]; // @[Modules.scala 53:83:@33058.4]
  assign buffer_8_632 = $signed(_T_82219); // @[Modules.scala 53:83:@33059.4]
  assign _T_82221 = $signed(buffer_8_482) + $signed(buffer_4_483); // @[Modules.scala 53:83:@33061.4]
  assign _T_82222 = _T_82221[10:0]; // @[Modules.scala 53:83:@33062.4]
  assign buffer_8_633 = $signed(_T_82222); // @[Modules.scala 53:83:@33063.4]
  assign _T_82224 = $signed(buffer_3_484) + $signed(buffer_0_485); // @[Modules.scala 53:83:@33065.4]
  assign _T_82225 = _T_82224[10:0]; // @[Modules.scala 53:83:@33066.4]
  assign buffer_8_634 = $signed(_T_82225); // @[Modules.scala 53:83:@33067.4]
  assign _T_82227 = $signed(buffer_8_486) + $signed(buffer_1_487); // @[Modules.scala 53:83:@33069.4]
  assign _T_82228 = _T_82227[10:0]; // @[Modules.scala 53:83:@33070.4]
  assign buffer_8_635 = $signed(_T_82228); // @[Modules.scala 53:83:@33071.4]
  assign _T_82230 = $signed(buffer_8_488) + $signed(buffer_5_489); // @[Modules.scala 53:83:@33073.4]
  assign _T_82231 = _T_82230[10:0]; // @[Modules.scala 53:83:@33074.4]
  assign buffer_8_636 = $signed(_T_82231); // @[Modules.scala 53:83:@33075.4]
  assign _T_82233 = $signed(buffer_8_490) + $signed(buffer_0_491); // @[Modules.scala 53:83:@33077.4]
  assign _T_82234 = _T_82233[10:0]; // @[Modules.scala 53:83:@33078.4]
  assign buffer_8_637 = $signed(_T_82234); // @[Modules.scala 53:83:@33079.4]
  assign _T_82236 = $signed(buffer_8_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@33081.4]
  assign _T_82237 = _T_82236[10:0]; // @[Modules.scala 53:83:@33082.4]
  assign buffer_8_638 = $signed(_T_82237); // @[Modules.scala 53:83:@33083.4]
  assign _T_82239 = $signed(buffer_8_494) + $signed(buffer_8_495); // @[Modules.scala 53:83:@33085.4]
  assign _T_82240 = _T_82239[10:0]; // @[Modules.scala 53:83:@33086.4]
  assign buffer_8_639 = $signed(_T_82240); // @[Modules.scala 53:83:@33087.4]
  assign _T_82245 = $signed(buffer_7_498) + $signed(buffer_2_499); // @[Modules.scala 53:83:@33093.4]
  assign _T_82246 = _T_82245[10:0]; // @[Modules.scala 53:83:@33094.4]
  assign buffer_8_641 = $signed(_T_82246); // @[Modules.scala 53:83:@33095.4]
  assign _T_82248 = $signed(buffer_0_500) + $signed(buffer_6_501); // @[Modules.scala 53:83:@33097.4]
  assign _T_82249 = _T_82248[10:0]; // @[Modules.scala 53:83:@33098.4]
  assign buffer_8_642 = $signed(_T_82249); // @[Modules.scala 53:83:@33099.4]
  assign _T_82251 = $signed(buffer_8_502) + $signed(buffer_8_503); // @[Modules.scala 53:83:@33101.4]
  assign _T_82252 = _T_82251[10:0]; // @[Modules.scala 53:83:@33102.4]
  assign buffer_8_643 = $signed(_T_82252); // @[Modules.scala 53:83:@33103.4]
  assign _T_82254 = $signed(buffer_8_504) + $signed(buffer_3_505); // @[Modules.scala 53:83:@33105.4]
  assign _T_82255 = _T_82254[10:0]; // @[Modules.scala 53:83:@33106.4]
  assign buffer_8_644 = $signed(_T_82255); // @[Modules.scala 53:83:@33107.4]
  assign _T_82260 = $signed(buffer_0_508) + $signed(buffer_7_509); // @[Modules.scala 53:83:@33113.4]
  assign _T_82261 = _T_82260[10:0]; // @[Modules.scala 53:83:@33114.4]
  assign buffer_8_646 = $signed(_T_82261); // @[Modules.scala 53:83:@33115.4]
  assign _T_82263 = $signed(buffer_5_510) + $signed(buffer_8_511); // @[Modules.scala 53:83:@33117.4]
  assign _T_82264 = _T_82263[10:0]; // @[Modules.scala 53:83:@33118.4]
  assign buffer_8_647 = $signed(_T_82264); // @[Modules.scala 53:83:@33119.4]
  assign _T_82266 = $signed(buffer_4_512) + $signed(buffer_5_513); // @[Modules.scala 53:83:@33121.4]
  assign _T_82267 = _T_82266[10:0]; // @[Modules.scala 53:83:@33122.4]
  assign buffer_8_648 = $signed(_T_82267); // @[Modules.scala 53:83:@33123.4]
  assign _T_82269 = $signed(buffer_2_514) + $signed(buffer_8_515); // @[Modules.scala 53:83:@33125.4]
  assign _T_82270 = _T_82269[10:0]; // @[Modules.scala 53:83:@33126.4]
  assign buffer_8_649 = $signed(_T_82270); // @[Modules.scala 53:83:@33127.4]
  assign _T_82272 = $signed(buffer_8_516) + $signed(buffer_3_517); // @[Modules.scala 53:83:@33129.4]
  assign _T_82273 = _T_82272[10:0]; // @[Modules.scala 53:83:@33130.4]
  assign buffer_8_650 = $signed(_T_82273); // @[Modules.scala 53:83:@33131.4]
  assign _T_82275 = $signed(buffer_8_518) + $signed(buffer_8_519); // @[Modules.scala 53:83:@33133.4]
  assign _T_82276 = _T_82275[10:0]; // @[Modules.scala 53:83:@33134.4]
  assign buffer_8_651 = $signed(_T_82276); // @[Modules.scala 53:83:@33135.4]
  assign _T_82278 = $signed(buffer_3_520) + $signed(buffer_5_521); // @[Modules.scala 53:83:@33137.4]
  assign _T_82279 = _T_82278[10:0]; // @[Modules.scala 53:83:@33138.4]
  assign buffer_8_652 = $signed(_T_82279); // @[Modules.scala 53:83:@33139.4]
  assign _T_82281 = $signed(buffer_6_522) + $signed(buffer_7_523); // @[Modules.scala 53:83:@33141.4]
  assign _T_82282 = _T_82281[10:0]; // @[Modules.scala 53:83:@33142.4]
  assign buffer_8_653 = $signed(_T_82282); // @[Modules.scala 53:83:@33143.4]
  assign _T_82284 = $signed(buffer_3_524) + $signed(buffer_8_525); // @[Modules.scala 53:83:@33145.4]
  assign _T_82285 = _T_82284[10:0]; // @[Modules.scala 53:83:@33146.4]
  assign buffer_8_654 = $signed(_T_82285); // @[Modules.scala 53:83:@33147.4]
  assign _T_82287 = $signed(buffer_8_526) + $signed(buffer_6_527); // @[Modules.scala 53:83:@33149.4]
  assign _T_82288 = _T_82287[10:0]; // @[Modules.scala 53:83:@33150.4]
  assign buffer_8_655 = $signed(_T_82288); // @[Modules.scala 53:83:@33151.4]
  assign _T_82290 = $signed(buffer_8_528) + $signed(buffer_3_529); // @[Modules.scala 53:83:@33153.4]
  assign _T_82291 = _T_82290[10:0]; // @[Modules.scala 53:83:@33154.4]
  assign buffer_8_656 = $signed(_T_82291); // @[Modules.scala 53:83:@33155.4]
  assign _T_82293 = $signed(buffer_8_530) + $signed(buffer_5_531); // @[Modules.scala 53:83:@33157.4]
  assign _T_82294 = _T_82293[10:0]; // @[Modules.scala 53:83:@33158.4]
  assign buffer_8_657 = $signed(_T_82294); // @[Modules.scala 53:83:@33159.4]
  assign _T_82296 = $signed(buffer_8_532) + $signed(buffer_8_533); // @[Modules.scala 53:83:@33161.4]
  assign _T_82297 = _T_82296[10:0]; // @[Modules.scala 53:83:@33162.4]
  assign buffer_8_658 = $signed(_T_82297); // @[Modules.scala 53:83:@33163.4]
  assign _T_82299 = $signed(buffer_8_534) + $signed(buffer_5_535); // @[Modules.scala 53:83:@33165.4]
  assign _T_82300 = _T_82299[10:0]; // @[Modules.scala 53:83:@33166.4]
  assign buffer_8_659 = $signed(_T_82300); // @[Modules.scala 53:83:@33167.4]
  assign _T_82302 = $signed(buffer_0_536) + $signed(buffer_4_537); // @[Modules.scala 53:83:@33169.4]
  assign _T_82303 = _T_82302[10:0]; // @[Modules.scala 53:83:@33170.4]
  assign buffer_8_660 = $signed(_T_82303); // @[Modules.scala 53:83:@33171.4]
  assign _T_82305 = $signed(buffer_8_538) + $signed(buffer_1_539); // @[Modules.scala 53:83:@33173.4]
  assign _T_82306 = _T_82305[10:0]; // @[Modules.scala 53:83:@33174.4]
  assign buffer_8_661 = $signed(_T_82306); // @[Modules.scala 53:83:@33175.4]
  assign _T_82308 = $signed(buffer_1_540) + $signed(buffer_8_541); // @[Modules.scala 53:83:@33177.4]
  assign _T_82309 = _T_82308[10:0]; // @[Modules.scala 53:83:@33178.4]
  assign buffer_8_662 = $signed(_T_82309); // @[Modules.scala 53:83:@33179.4]
  assign _T_82311 = $signed(buffer_8_542) + $signed(buffer_8_543); // @[Modules.scala 53:83:@33181.4]
  assign _T_82312 = _T_82311[10:0]; // @[Modules.scala 53:83:@33182.4]
  assign buffer_8_663 = $signed(_T_82312); // @[Modules.scala 53:83:@33183.4]
  assign _T_82317 = $signed(buffer_1_546) + $signed(buffer_8_547); // @[Modules.scala 53:83:@33189.4]
  assign _T_82318 = _T_82317[10:0]; // @[Modules.scala 53:83:@33190.4]
  assign buffer_8_665 = $signed(_T_82318); // @[Modules.scala 53:83:@33191.4]
  assign _T_82320 = $signed(buffer_8_548) + $signed(buffer_8_549); // @[Modules.scala 53:83:@33193.4]
  assign _T_82321 = _T_82320[10:0]; // @[Modules.scala 53:83:@33194.4]
  assign buffer_8_666 = $signed(_T_82321); // @[Modules.scala 53:83:@33195.4]
  assign _T_82329 = $signed(buffer_8_554) + $signed(buffer_8_555); // @[Modules.scala 53:83:@33205.4]
  assign _T_82330 = _T_82329[10:0]; // @[Modules.scala 53:83:@33206.4]
  assign buffer_8_669 = $signed(_T_82330); // @[Modules.scala 53:83:@33207.4]
  assign _T_82332 = $signed(buffer_0_556) + $signed(buffer_8_557); // @[Modules.scala 53:83:@33209.4]
  assign _T_82333 = _T_82332[10:0]; // @[Modules.scala 53:83:@33210.4]
  assign buffer_8_670 = $signed(_T_82333); // @[Modules.scala 53:83:@33211.4]
  assign _T_82335 = $signed(buffer_1_558) + $signed(buffer_8_559); // @[Modules.scala 53:83:@33213.4]
  assign _T_82336 = _T_82335[10:0]; // @[Modules.scala 53:83:@33214.4]
  assign buffer_8_671 = $signed(_T_82336); // @[Modules.scala 53:83:@33215.4]
  assign _T_82338 = $signed(buffer_5_560) + $signed(buffer_8_561); // @[Modules.scala 53:83:@33217.4]
  assign _T_82339 = _T_82338[10:0]; // @[Modules.scala 53:83:@33218.4]
  assign buffer_8_672 = $signed(_T_82339); // @[Modules.scala 53:83:@33219.4]
  assign _T_82347 = $signed(buffer_4_566) + $signed(buffer_8_567); // @[Modules.scala 53:83:@33229.4]
  assign _T_82348 = _T_82347[10:0]; // @[Modules.scala 53:83:@33230.4]
  assign buffer_8_675 = $signed(_T_82348); // @[Modules.scala 53:83:@33231.4]
  assign _T_82368 = $signed(buffer_8_580) + $signed(buffer_8_581); // @[Modules.scala 53:83:@33257.4]
  assign _T_82369 = _T_82368[10:0]; // @[Modules.scala 53:83:@33258.4]
  assign buffer_8_682 = $signed(_T_82369); // @[Modules.scala 53:83:@33259.4]
  assign _T_82371 = $signed(buffer_4_582) + $signed(buffer_8_583); // @[Modules.scala 53:83:@33261.4]
  assign _T_82372 = _T_82371[10:0]; // @[Modules.scala 53:83:@33262.4]
  assign buffer_8_683 = $signed(_T_82372); // @[Modules.scala 53:83:@33263.4]
  assign _T_82377 = $signed(buffer_8_586) + $signed(buffer_1_587); // @[Modules.scala 53:83:@33269.4]
  assign _T_82378 = _T_82377[10:0]; // @[Modules.scala 53:83:@33270.4]
  assign buffer_8_685 = $signed(_T_82378); // @[Modules.scala 53:83:@33271.4]
  assign _T_82380 = $signed(buffer_4_588) + $signed(buffer_8_589); // @[Modules.scala 56:109:@33273.4]
  assign _T_82381 = _T_82380[10:0]; // @[Modules.scala 56:109:@33274.4]
  assign buffer_8_686 = $signed(_T_82381); // @[Modules.scala 56:109:@33275.4]
  assign _T_82383 = $signed(buffer_8_590) + $signed(buffer_8_591); // @[Modules.scala 56:109:@33277.4]
  assign _T_82384 = _T_82383[10:0]; // @[Modules.scala 56:109:@33278.4]
  assign buffer_8_687 = $signed(_T_82384); // @[Modules.scala 56:109:@33279.4]
  assign _T_82386 = $signed(buffer_8_592) + $signed(buffer_0_593); // @[Modules.scala 56:109:@33281.4]
  assign _T_82387 = _T_82386[10:0]; // @[Modules.scala 56:109:@33282.4]
  assign buffer_8_688 = $signed(_T_82387); // @[Modules.scala 56:109:@33283.4]
  assign _T_82389 = $signed(buffer_8_594) + $signed(buffer_0_595); // @[Modules.scala 56:109:@33285.4]
  assign _T_82390 = _T_82389[10:0]; // @[Modules.scala 56:109:@33286.4]
  assign buffer_8_689 = $signed(_T_82390); // @[Modules.scala 56:109:@33287.4]
  assign _T_82395 = $signed(buffer_8_598) + $signed(buffer_8_599); // @[Modules.scala 56:109:@33293.4]
  assign _T_82396 = _T_82395[10:0]; // @[Modules.scala 56:109:@33294.4]
  assign buffer_8_691 = $signed(_T_82396); // @[Modules.scala 56:109:@33295.4]
  assign _T_82398 = $signed(buffer_6_600) + $signed(buffer_8_601); // @[Modules.scala 56:109:@33297.4]
  assign _T_82399 = _T_82398[10:0]; // @[Modules.scala 56:109:@33298.4]
  assign buffer_8_692 = $signed(_T_82399); // @[Modules.scala 56:109:@33299.4]
  assign _T_82401 = $signed(buffer_8_602) + $signed(buffer_8_603); // @[Modules.scala 56:109:@33301.4]
  assign _T_82402 = _T_82401[10:0]; // @[Modules.scala 56:109:@33302.4]
  assign buffer_8_693 = $signed(_T_82402); // @[Modules.scala 56:109:@33303.4]
  assign _T_82404 = $signed(buffer_8_604) + $signed(buffer_8_605); // @[Modules.scala 56:109:@33305.4]
  assign _T_82405 = _T_82404[10:0]; // @[Modules.scala 56:109:@33306.4]
  assign buffer_8_694 = $signed(_T_82405); // @[Modules.scala 56:109:@33307.4]
  assign _T_82410 = $signed(buffer_8_608) + $signed(buffer_3_609); // @[Modules.scala 56:109:@33313.4]
  assign _T_82411 = _T_82410[10:0]; // @[Modules.scala 56:109:@33314.4]
  assign buffer_8_696 = $signed(_T_82411); // @[Modules.scala 56:109:@33315.4]
  assign _T_82413 = $signed(buffer_8_610) + $signed(buffer_8_611); // @[Modules.scala 56:109:@33317.4]
  assign _T_82414 = _T_82413[10:0]; // @[Modules.scala 56:109:@33318.4]
  assign buffer_8_697 = $signed(_T_82414); // @[Modules.scala 56:109:@33319.4]
  assign _T_82416 = $signed(buffer_8_612) + $signed(buffer_8_613); // @[Modules.scala 56:109:@33321.4]
  assign _T_82417 = _T_82416[10:0]; // @[Modules.scala 56:109:@33322.4]
  assign buffer_8_698 = $signed(_T_82417); // @[Modules.scala 56:109:@33323.4]
  assign _T_82419 = $signed(buffer_8_614) + $signed(buffer_8_615); // @[Modules.scala 56:109:@33325.4]
  assign _T_82420 = _T_82419[10:0]; // @[Modules.scala 56:109:@33326.4]
  assign buffer_8_699 = $signed(_T_82420); // @[Modules.scala 56:109:@33327.4]
  assign _T_82422 = $signed(buffer_8_616) + $signed(buffer_8_617); // @[Modules.scala 56:109:@33329.4]
  assign _T_82423 = _T_82422[10:0]; // @[Modules.scala 56:109:@33330.4]
  assign buffer_8_700 = $signed(_T_82423); // @[Modules.scala 56:109:@33331.4]
  assign _T_82425 = $signed(buffer_8_618) + $signed(buffer_8_619); // @[Modules.scala 56:109:@33333.4]
  assign _T_82426 = _T_82425[10:0]; // @[Modules.scala 56:109:@33334.4]
  assign buffer_8_701 = $signed(_T_82426); // @[Modules.scala 56:109:@33335.4]
  assign _T_82428 = $signed(buffer_8_620) + $signed(buffer_8_621); // @[Modules.scala 56:109:@33337.4]
  assign _T_82429 = _T_82428[10:0]; // @[Modules.scala 56:109:@33338.4]
  assign buffer_8_702 = $signed(_T_82429); // @[Modules.scala 56:109:@33339.4]
  assign _T_82431 = $signed(buffer_8_622) + $signed(buffer_8_623); // @[Modules.scala 56:109:@33341.4]
  assign _T_82432 = _T_82431[10:0]; // @[Modules.scala 56:109:@33342.4]
  assign buffer_8_703 = $signed(_T_82432); // @[Modules.scala 56:109:@33343.4]
  assign _T_82434 = $signed(buffer_5_624) + $signed(buffer_8_625); // @[Modules.scala 56:109:@33345.4]
  assign _T_82435 = _T_82434[10:0]; // @[Modules.scala 56:109:@33346.4]
  assign buffer_8_704 = $signed(_T_82435); // @[Modules.scala 56:109:@33347.4]
  assign _T_82437 = $signed(buffer_8_626) + $signed(buffer_3_627); // @[Modules.scala 56:109:@33349.4]
  assign _T_82438 = _T_82437[10:0]; // @[Modules.scala 56:109:@33350.4]
  assign buffer_8_705 = $signed(_T_82438); // @[Modules.scala 56:109:@33351.4]
  assign _T_82440 = $signed(buffer_8_628) + $signed(buffer_8_629); // @[Modules.scala 56:109:@33353.4]
  assign _T_82441 = _T_82440[10:0]; // @[Modules.scala 56:109:@33354.4]
  assign buffer_8_706 = $signed(_T_82441); // @[Modules.scala 56:109:@33355.4]
  assign _T_82443 = $signed(buffer_8_630) + $signed(buffer_5_631); // @[Modules.scala 56:109:@33357.4]
  assign _T_82444 = _T_82443[10:0]; // @[Modules.scala 56:109:@33358.4]
  assign buffer_8_707 = $signed(_T_82444); // @[Modules.scala 56:109:@33359.4]
  assign _T_82446 = $signed(buffer_8_632) + $signed(buffer_8_633); // @[Modules.scala 56:109:@33361.4]
  assign _T_82447 = _T_82446[10:0]; // @[Modules.scala 56:109:@33362.4]
  assign buffer_8_708 = $signed(_T_82447); // @[Modules.scala 56:109:@33363.4]
  assign _T_82449 = $signed(buffer_8_634) + $signed(buffer_8_635); // @[Modules.scala 56:109:@33365.4]
  assign _T_82450 = _T_82449[10:0]; // @[Modules.scala 56:109:@33366.4]
  assign buffer_8_709 = $signed(_T_82450); // @[Modules.scala 56:109:@33367.4]
  assign _T_82452 = $signed(buffer_8_636) + $signed(buffer_8_637); // @[Modules.scala 56:109:@33369.4]
  assign _T_82453 = _T_82452[10:0]; // @[Modules.scala 56:109:@33370.4]
  assign buffer_8_710 = $signed(_T_82453); // @[Modules.scala 56:109:@33371.4]
  assign _T_82455 = $signed(buffer_8_638) + $signed(buffer_8_639); // @[Modules.scala 56:109:@33373.4]
  assign _T_82456 = _T_82455[10:0]; // @[Modules.scala 56:109:@33374.4]
  assign buffer_8_711 = $signed(_T_82456); // @[Modules.scala 56:109:@33375.4]
  assign _T_82458 = $signed(buffer_3_640) + $signed(buffer_8_641); // @[Modules.scala 56:109:@33377.4]
  assign _T_82459 = _T_82458[10:0]; // @[Modules.scala 56:109:@33378.4]
  assign buffer_8_712 = $signed(_T_82459); // @[Modules.scala 56:109:@33379.4]
  assign _T_82461 = $signed(buffer_8_642) + $signed(buffer_8_643); // @[Modules.scala 56:109:@33381.4]
  assign _T_82462 = _T_82461[10:0]; // @[Modules.scala 56:109:@33382.4]
  assign buffer_8_713 = $signed(_T_82462); // @[Modules.scala 56:109:@33383.4]
  assign _T_82464 = $signed(buffer_8_644) + $signed(buffer_2_645); // @[Modules.scala 56:109:@33385.4]
  assign _T_82465 = _T_82464[10:0]; // @[Modules.scala 56:109:@33386.4]
  assign buffer_8_714 = $signed(_T_82465); // @[Modules.scala 56:109:@33387.4]
  assign _T_82467 = $signed(buffer_8_646) + $signed(buffer_8_647); // @[Modules.scala 56:109:@33389.4]
  assign _T_82468 = _T_82467[10:0]; // @[Modules.scala 56:109:@33390.4]
  assign buffer_8_715 = $signed(_T_82468); // @[Modules.scala 56:109:@33391.4]
  assign _T_82470 = $signed(buffer_8_648) + $signed(buffer_8_649); // @[Modules.scala 56:109:@33393.4]
  assign _T_82471 = _T_82470[10:0]; // @[Modules.scala 56:109:@33394.4]
  assign buffer_8_716 = $signed(_T_82471); // @[Modules.scala 56:109:@33395.4]
  assign _T_82473 = $signed(buffer_8_650) + $signed(buffer_8_651); // @[Modules.scala 56:109:@33397.4]
  assign _T_82474 = _T_82473[10:0]; // @[Modules.scala 56:109:@33398.4]
  assign buffer_8_717 = $signed(_T_82474); // @[Modules.scala 56:109:@33399.4]
  assign _T_82476 = $signed(buffer_8_652) + $signed(buffer_8_653); // @[Modules.scala 56:109:@33401.4]
  assign _T_82477 = _T_82476[10:0]; // @[Modules.scala 56:109:@33402.4]
  assign buffer_8_718 = $signed(_T_82477); // @[Modules.scala 56:109:@33403.4]
  assign _T_82479 = $signed(buffer_8_654) + $signed(buffer_8_655); // @[Modules.scala 56:109:@33405.4]
  assign _T_82480 = _T_82479[10:0]; // @[Modules.scala 56:109:@33406.4]
  assign buffer_8_719 = $signed(_T_82480); // @[Modules.scala 56:109:@33407.4]
  assign _T_82482 = $signed(buffer_8_656) + $signed(buffer_8_657); // @[Modules.scala 56:109:@33409.4]
  assign _T_82483 = _T_82482[10:0]; // @[Modules.scala 56:109:@33410.4]
  assign buffer_8_720 = $signed(_T_82483); // @[Modules.scala 56:109:@33411.4]
  assign _T_82485 = $signed(buffer_8_658) + $signed(buffer_8_659); // @[Modules.scala 56:109:@33413.4]
  assign _T_82486 = _T_82485[10:0]; // @[Modules.scala 56:109:@33414.4]
  assign buffer_8_721 = $signed(_T_82486); // @[Modules.scala 56:109:@33415.4]
  assign _T_82488 = $signed(buffer_8_660) + $signed(buffer_8_661); // @[Modules.scala 56:109:@33417.4]
  assign _T_82489 = _T_82488[10:0]; // @[Modules.scala 56:109:@33418.4]
  assign buffer_8_722 = $signed(_T_82489); // @[Modules.scala 56:109:@33419.4]
  assign _T_82491 = $signed(buffer_8_662) + $signed(buffer_8_663); // @[Modules.scala 56:109:@33421.4]
  assign _T_82492 = _T_82491[10:0]; // @[Modules.scala 56:109:@33422.4]
  assign buffer_8_723 = $signed(_T_82492); // @[Modules.scala 56:109:@33423.4]
  assign _T_82494 = $signed(buffer_3_664) + $signed(buffer_8_665); // @[Modules.scala 56:109:@33425.4]
  assign _T_82495 = _T_82494[10:0]; // @[Modules.scala 56:109:@33426.4]
  assign buffer_8_724 = $signed(_T_82495); // @[Modules.scala 56:109:@33427.4]
  assign _T_82497 = $signed(buffer_8_666) + $signed(buffer_4_667); // @[Modules.scala 56:109:@33429.4]
  assign _T_82498 = _T_82497[10:0]; // @[Modules.scala 56:109:@33430.4]
  assign buffer_8_725 = $signed(_T_82498); // @[Modules.scala 56:109:@33431.4]
  assign _T_82500 = $signed(buffer_3_668) + $signed(buffer_8_669); // @[Modules.scala 56:109:@33433.4]
  assign _T_82501 = _T_82500[10:0]; // @[Modules.scala 56:109:@33434.4]
  assign buffer_8_726 = $signed(_T_82501); // @[Modules.scala 56:109:@33435.4]
  assign _T_82503 = $signed(buffer_8_670) + $signed(buffer_8_671); // @[Modules.scala 56:109:@33437.4]
  assign _T_82504 = _T_82503[10:0]; // @[Modules.scala 56:109:@33438.4]
  assign buffer_8_727 = $signed(_T_82504); // @[Modules.scala 56:109:@33439.4]
  assign _T_82506 = $signed(buffer_8_672) + $signed(buffer_6_673); // @[Modules.scala 56:109:@33441.4]
  assign _T_82507 = _T_82506[10:0]; // @[Modules.scala 56:109:@33442.4]
  assign buffer_8_728 = $signed(_T_82507); // @[Modules.scala 56:109:@33443.4]
  assign _T_82509 = $signed(buffer_3_674) + $signed(buffer_8_675); // @[Modules.scala 56:109:@33445.4]
  assign _T_82510 = _T_82509[10:0]; // @[Modules.scala 56:109:@33446.4]
  assign buffer_8_729 = $signed(_T_82510); // @[Modules.scala 56:109:@33447.4]
  assign _T_82515 = $signed(buffer_4_678) + $signed(buffer_1_679); // @[Modules.scala 56:109:@33453.4]
  assign _T_82516 = _T_82515[10:0]; // @[Modules.scala 56:109:@33454.4]
  assign buffer_8_731 = $signed(_T_82516); // @[Modules.scala 56:109:@33455.4]
  assign _T_82521 = $signed(buffer_8_682) + $signed(buffer_8_683); // @[Modules.scala 56:109:@33461.4]
  assign _T_82522 = _T_82521[10:0]; // @[Modules.scala 56:109:@33462.4]
  assign buffer_8_733 = $signed(_T_82522); // @[Modules.scala 56:109:@33463.4]
  assign _T_82524 = $signed(buffer_1_684) + $signed(buffer_8_685); // @[Modules.scala 56:109:@33465.4]
  assign _T_82525 = _T_82524[10:0]; // @[Modules.scala 56:109:@33466.4]
  assign buffer_8_734 = $signed(_T_82525); // @[Modules.scala 56:109:@33467.4]
  assign _T_82527 = $signed(buffer_8_686) + $signed(buffer_8_687); // @[Modules.scala 63:156:@33470.4]
  assign _T_82528 = _T_82527[10:0]; // @[Modules.scala 63:156:@33471.4]
  assign buffer_8_736 = $signed(_T_82528); // @[Modules.scala 63:156:@33472.4]
  assign _T_82530 = $signed(buffer_8_736) + $signed(buffer_8_688); // @[Modules.scala 63:156:@33474.4]
  assign _T_82531 = _T_82530[10:0]; // @[Modules.scala 63:156:@33475.4]
  assign buffer_8_737 = $signed(_T_82531); // @[Modules.scala 63:156:@33476.4]
  assign _T_82533 = $signed(buffer_8_737) + $signed(buffer_8_689); // @[Modules.scala 63:156:@33478.4]
  assign _T_82534 = _T_82533[10:0]; // @[Modules.scala 63:156:@33479.4]
  assign buffer_8_738 = $signed(_T_82534); // @[Modules.scala 63:156:@33480.4]
  assign _T_82536 = $signed(buffer_8_738) + $signed(buffer_3_690); // @[Modules.scala 63:156:@33482.4]
  assign _T_82537 = _T_82536[10:0]; // @[Modules.scala 63:156:@33483.4]
  assign buffer_8_739 = $signed(_T_82537); // @[Modules.scala 63:156:@33484.4]
  assign _T_82539 = $signed(buffer_8_739) + $signed(buffer_8_691); // @[Modules.scala 63:156:@33486.4]
  assign _T_82540 = _T_82539[10:0]; // @[Modules.scala 63:156:@33487.4]
  assign buffer_8_740 = $signed(_T_82540); // @[Modules.scala 63:156:@33488.4]
  assign _T_82542 = $signed(buffer_8_740) + $signed(buffer_8_692); // @[Modules.scala 63:156:@33490.4]
  assign _T_82543 = _T_82542[10:0]; // @[Modules.scala 63:156:@33491.4]
  assign buffer_8_741 = $signed(_T_82543); // @[Modules.scala 63:156:@33492.4]
  assign _T_82545 = $signed(buffer_8_741) + $signed(buffer_8_693); // @[Modules.scala 63:156:@33494.4]
  assign _T_82546 = _T_82545[10:0]; // @[Modules.scala 63:156:@33495.4]
  assign buffer_8_742 = $signed(_T_82546); // @[Modules.scala 63:156:@33496.4]
  assign _T_82548 = $signed(buffer_8_742) + $signed(buffer_8_694); // @[Modules.scala 63:156:@33498.4]
  assign _T_82549 = _T_82548[10:0]; // @[Modules.scala 63:156:@33499.4]
  assign buffer_8_743 = $signed(_T_82549); // @[Modules.scala 63:156:@33500.4]
  assign _T_82551 = $signed(buffer_8_743) + $signed(buffer_4_695); // @[Modules.scala 63:156:@33502.4]
  assign _T_82552 = _T_82551[10:0]; // @[Modules.scala 63:156:@33503.4]
  assign buffer_8_744 = $signed(_T_82552); // @[Modules.scala 63:156:@33504.4]
  assign _T_82554 = $signed(buffer_8_744) + $signed(buffer_8_696); // @[Modules.scala 63:156:@33506.4]
  assign _T_82555 = _T_82554[10:0]; // @[Modules.scala 63:156:@33507.4]
  assign buffer_8_745 = $signed(_T_82555); // @[Modules.scala 63:156:@33508.4]
  assign _T_82557 = $signed(buffer_8_745) + $signed(buffer_8_697); // @[Modules.scala 63:156:@33510.4]
  assign _T_82558 = _T_82557[10:0]; // @[Modules.scala 63:156:@33511.4]
  assign buffer_8_746 = $signed(_T_82558); // @[Modules.scala 63:156:@33512.4]
  assign _T_82560 = $signed(buffer_8_746) + $signed(buffer_8_698); // @[Modules.scala 63:156:@33514.4]
  assign _T_82561 = _T_82560[10:0]; // @[Modules.scala 63:156:@33515.4]
  assign buffer_8_747 = $signed(_T_82561); // @[Modules.scala 63:156:@33516.4]
  assign _T_82563 = $signed(buffer_8_747) + $signed(buffer_8_699); // @[Modules.scala 63:156:@33518.4]
  assign _T_82564 = _T_82563[10:0]; // @[Modules.scala 63:156:@33519.4]
  assign buffer_8_748 = $signed(_T_82564); // @[Modules.scala 63:156:@33520.4]
  assign _T_82566 = $signed(buffer_8_748) + $signed(buffer_8_700); // @[Modules.scala 63:156:@33522.4]
  assign _T_82567 = _T_82566[10:0]; // @[Modules.scala 63:156:@33523.4]
  assign buffer_8_749 = $signed(_T_82567); // @[Modules.scala 63:156:@33524.4]
  assign _T_82569 = $signed(buffer_8_749) + $signed(buffer_8_701); // @[Modules.scala 63:156:@33526.4]
  assign _T_82570 = _T_82569[10:0]; // @[Modules.scala 63:156:@33527.4]
  assign buffer_8_750 = $signed(_T_82570); // @[Modules.scala 63:156:@33528.4]
  assign _T_82572 = $signed(buffer_8_750) + $signed(buffer_8_702); // @[Modules.scala 63:156:@33530.4]
  assign _T_82573 = _T_82572[10:0]; // @[Modules.scala 63:156:@33531.4]
  assign buffer_8_751 = $signed(_T_82573); // @[Modules.scala 63:156:@33532.4]
  assign _T_82575 = $signed(buffer_8_751) + $signed(buffer_8_703); // @[Modules.scala 63:156:@33534.4]
  assign _T_82576 = _T_82575[10:0]; // @[Modules.scala 63:156:@33535.4]
  assign buffer_8_752 = $signed(_T_82576); // @[Modules.scala 63:156:@33536.4]
  assign _T_82578 = $signed(buffer_8_752) + $signed(buffer_8_704); // @[Modules.scala 63:156:@33538.4]
  assign _T_82579 = _T_82578[10:0]; // @[Modules.scala 63:156:@33539.4]
  assign buffer_8_753 = $signed(_T_82579); // @[Modules.scala 63:156:@33540.4]
  assign _T_82581 = $signed(buffer_8_753) + $signed(buffer_8_705); // @[Modules.scala 63:156:@33542.4]
  assign _T_82582 = _T_82581[10:0]; // @[Modules.scala 63:156:@33543.4]
  assign buffer_8_754 = $signed(_T_82582); // @[Modules.scala 63:156:@33544.4]
  assign _T_82584 = $signed(buffer_8_754) + $signed(buffer_8_706); // @[Modules.scala 63:156:@33546.4]
  assign _T_82585 = _T_82584[10:0]; // @[Modules.scala 63:156:@33547.4]
  assign buffer_8_755 = $signed(_T_82585); // @[Modules.scala 63:156:@33548.4]
  assign _T_82587 = $signed(buffer_8_755) + $signed(buffer_8_707); // @[Modules.scala 63:156:@33550.4]
  assign _T_82588 = _T_82587[10:0]; // @[Modules.scala 63:156:@33551.4]
  assign buffer_8_756 = $signed(_T_82588); // @[Modules.scala 63:156:@33552.4]
  assign _T_82590 = $signed(buffer_8_756) + $signed(buffer_8_708); // @[Modules.scala 63:156:@33554.4]
  assign _T_82591 = _T_82590[10:0]; // @[Modules.scala 63:156:@33555.4]
  assign buffer_8_757 = $signed(_T_82591); // @[Modules.scala 63:156:@33556.4]
  assign _T_82593 = $signed(buffer_8_757) + $signed(buffer_8_709); // @[Modules.scala 63:156:@33558.4]
  assign _T_82594 = _T_82593[10:0]; // @[Modules.scala 63:156:@33559.4]
  assign buffer_8_758 = $signed(_T_82594); // @[Modules.scala 63:156:@33560.4]
  assign _T_82596 = $signed(buffer_8_758) + $signed(buffer_8_710); // @[Modules.scala 63:156:@33562.4]
  assign _T_82597 = _T_82596[10:0]; // @[Modules.scala 63:156:@33563.4]
  assign buffer_8_759 = $signed(_T_82597); // @[Modules.scala 63:156:@33564.4]
  assign _T_82599 = $signed(buffer_8_759) + $signed(buffer_8_711); // @[Modules.scala 63:156:@33566.4]
  assign _T_82600 = _T_82599[10:0]; // @[Modules.scala 63:156:@33567.4]
  assign buffer_8_760 = $signed(_T_82600); // @[Modules.scala 63:156:@33568.4]
  assign _T_82602 = $signed(buffer_8_760) + $signed(buffer_8_712); // @[Modules.scala 63:156:@33570.4]
  assign _T_82603 = _T_82602[10:0]; // @[Modules.scala 63:156:@33571.4]
  assign buffer_8_761 = $signed(_T_82603); // @[Modules.scala 63:156:@33572.4]
  assign _T_82605 = $signed(buffer_8_761) + $signed(buffer_8_713); // @[Modules.scala 63:156:@33574.4]
  assign _T_82606 = _T_82605[10:0]; // @[Modules.scala 63:156:@33575.4]
  assign buffer_8_762 = $signed(_T_82606); // @[Modules.scala 63:156:@33576.4]
  assign _T_82608 = $signed(buffer_8_762) + $signed(buffer_8_714); // @[Modules.scala 63:156:@33578.4]
  assign _T_82609 = _T_82608[10:0]; // @[Modules.scala 63:156:@33579.4]
  assign buffer_8_763 = $signed(_T_82609); // @[Modules.scala 63:156:@33580.4]
  assign _T_82611 = $signed(buffer_8_763) + $signed(buffer_8_715); // @[Modules.scala 63:156:@33582.4]
  assign _T_82612 = _T_82611[10:0]; // @[Modules.scala 63:156:@33583.4]
  assign buffer_8_764 = $signed(_T_82612); // @[Modules.scala 63:156:@33584.4]
  assign _T_82614 = $signed(buffer_8_764) + $signed(buffer_8_716); // @[Modules.scala 63:156:@33586.4]
  assign _T_82615 = _T_82614[10:0]; // @[Modules.scala 63:156:@33587.4]
  assign buffer_8_765 = $signed(_T_82615); // @[Modules.scala 63:156:@33588.4]
  assign _T_82617 = $signed(buffer_8_765) + $signed(buffer_8_717); // @[Modules.scala 63:156:@33590.4]
  assign _T_82618 = _T_82617[10:0]; // @[Modules.scala 63:156:@33591.4]
  assign buffer_8_766 = $signed(_T_82618); // @[Modules.scala 63:156:@33592.4]
  assign _T_82620 = $signed(buffer_8_766) + $signed(buffer_8_718); // @[Modules.scala 63:156:@33594.4]
  assign _T_82621 = _T_82620[10:0]; // @[Modules.scala 63:156:@33595.4]
  assign buffer_8_767 = $signed(_T_82621); // @[Modules.scala 63:156:@33596.4]
  assign _T_82623 = $signed(buffer_8_767) + $signed(buffer_8_719); // @[Modules.scala 63:156:@33598.4]
  assign _T_82624 = _T_82623[10:0]; // @[Modules.scala 63:156:@33599.4]
  assign buffer_8_768 = $signed(_T_82624); // @[Modules.scala 63:156:@33600.4]
  assign _T_82626 = $signed(buffer_8_768) + $signed(buffer_8_720); // @[Modules.scala 63:156:@33602.4]
  assign _T_82627 = _T_82626[10:0]; // @[Modules.scala 63:156:@33603.4]
  assign buffer_8_769 = $signed(_T_82627); // @[Modules.scala 63:156:@33604.4]
  assign _T_82629 = $signed(buffer_8_769) + $signed(buffer_8_721); // @[Modules.scala 63:156:@33606.4]
  assign _T_82630 = _T_82629[10:0]; // @[Modules.scala 63:156:@33607.4]
  assign buffer_8_770 = $signed(_T_82630); // @[Modules.scala 63:156:@33608.4]
  assign _T_82632 = $signed(buffer_8_770) + $signed(buffer_8_722); // @[Modules.scala 63:156:@33610.4]
  assign _T_82633 = _T_82632[10:0]; // @[Modules.scala 63:156:@33611.4]
  assign buffer_8_771 = $signed(_T_82633); // @[Modules.scala 63:156:@33612.4]
  assign _T_82635 = $signed(buffer_8_771) + $signed(buffer_8_723); // @[Modules.scala 63:156:@33614.4]
  assign _T_82636 = _T_82635[10:0]; // @[Modules.scala 63:156:@33615.4]
  assign buffer_8_772 = $signed(_T_82636); // @[Modules.scala 63:156:@33616.4]
  assign _T_82638 = $signed(buffer_8_772) + $signed(buffer_8_724); // @[Modules.scala 63:156:@33618.4]
  assign _T_82639 = _T_82638[10:0]; // @[Modules.scala 63:156:@33619.4]
  assign buffer_8_773 = $signed(_T_82639); // @[Modules.scala 63:156:@33620.4]
  assign _T_82641 = $signed(buffer_8_773) + $signed(buffer_8_725); // @[Modules.scala 63:156:@33622.4]
  assign _T_82642 = _T_82641[10:0]; // @[Modules.scala 63:156:@33623.4]
  assign buffer_8_774 = $signed(_T_82642); // @[Modules.scala 63:156:@33624.4]
  assign _T_82644 = $signed(buffer_8_774) + $signed(buffer_8_726); // @[Modules.scala 63:156:@33626.4]
  assign _T_82645 = _T_82644[10:0]; // @[Modules.scala 63:156:@33627.4]
  assign buffer_8_775 = $signed(_T_82645); // @[Modules.scala 63:156:@33628.4]
  assign _T_82647 = $signed(buffer_8_775) + $signed(buffer_8_727); // @[Modules.scala 63:156:@33630.4]
  assign _T_82648 = _T_82647[10:0]; // @[Modules.scala 63:156:@33631.4]
  assign buffer_8_776 = $signed(_T_82648); // @[Modules.scala 63:156:@33632.4]
  assign _T_82650 = $signed(buffer_8_776) + $signed(buffer_8_728); // @[Modules.scala 63:156:@33634.4]
  assign _T_82651 = _T_82650[10:0]; // @[Modules.scala 63:156:@33635.4]
  assign buffer_8_777 = $signed(_T_82651); // @[Modules.scala 63:156:@33636.4]
  assign _T_82653 = $signed(buffer_8_777) + $signed(buffer_8_729); // @[Modules.scala 63:156:@33638.4]
  assign _T_82654 = _T_82653[10:0]; // @[Modules.scala 63:156:@33639.4]
  assign buffer_8_778 = $signed(_T_82654); // @[Modules.scala 63:156:@33640.4]
  assign _T_82656 = $signed(buffer_8_778) + $signed(buffer_2_730); // @[Modules.scala 63:156:@33642.4]
  assign _T_82657 = _T_82656[10:0]; // @[Modules.scala 63:156:@33643.4]
  assign buffer_8_779 = $signed(_T_82657); // @[Modules.scala 63:156:@33644.4]
  assign _T_82659 = $signed(buffer_8_779) + $signed(buffer_8_731); // @[Modules.scala 63:156:@33646.4]
  assign _T_82660 = _T_82659[10:0]; // @[Modules.scala 63:156:@33647.4]
  assign buffer_8_780 = $signed(_T_82660); // @[Modules.scala 63:156:@33648.4]
  assign _T_82662 = $signed(buffer_8_780) + $signed(buffer_4_732); // @[Modules.scala 63:156:@33650.4]
  assign _T_82663 = _T_82662[10:0]; // @[Modules.scala 63:156:@33651.4]
  assign buffer_8_781 = $signed(_T_82663); // @[Modules.scala 63:156:@33652.4]
  assign _T_82665 = $signed(buffer_8_781) + $signed(buffer_8_733); // @[Modules.scala 63:156:@33654.4]
  assign _T_82666 = _T_82665[10:0]; // @[Modules.scala 63:156:@33655.4]
  assign buffer_8_782 = $signed(_T_82666); // @[Modules.scala 63:156:@33656.4]
  assign _T_82668 = $signed(buffer_8_782) + $signed(buffer_8_734); // @[Modules.scala 63:156:@33658.4]
  assign _T_82669 = _T_82668[10:0]; // @[Modules.scala 63:156:@33659.4]
  assign buffer_8_783 = $signed(_T_82669); // @[Modules.scala 63:156:@33660.4]
  assign _T_82678 = $signed(io_in_2) + $signed(io_in_3); // @[Modules.scala 37:46:@33670.4]
  assign _T_82679 = _T_82678[4:0]; // @[Modules.scala 37:46:@33671.4]
  assign _T_82680 = $signed(_T_82679); // @[Modules.scala 37:46:@33672.4]
  assign _T_82685 = $signed(_T_54283) - $signed(io_in_5); // @[Modules.scala 46:47:@33677.4]
  assign _T_82686 = _T_82685[4:0]; // @[Modules.scala 46:47:@33678.4]
  assign _T_82687 = $signed(_T_82686); // @[Modules.scala 46:47:@33679.4]
  assign _T_82730 = $signed(io_in_18) + $signed(io_in_19); // @[Modules.scala 37:46:@33723.4]
  assign _T_82731 = _T_82730[4:0]; // @[Modules.scala 37:46:@33724.4]
  assign _T_82732 = $signed(_T_82731); // @[Modules.scala 37:46:@33725.4]
  assign _T_82858 = $signed(_T_57701) + $signed(io_in_83); // @[Modules.scala 43:47:@33875.4]
  assign _T_82859 = _T_82858[4:0]; // @[Modules.scala 43:47:@33876.4]
  assign _T_82860 = $signed(_T_82859); // @[Modules.scala 43:47:@33877.4]
  assign _T_82996 = $signed(_T_54674) + $signed(io_in_151); // @[Modules.scala 43:47:@34038.4]
  assign _T_82997 = _T_82996[4:0]; // @[Modules.scala 43:47:@34039.4]
  assign _T_82998 = $signed(_T_82997); // @[Modules.scala 43:47:@34040.4]
  assign _T_83013 = $signed(_T_54695) + $signed(io_in_157); // @[Modules.scala 43:47:@34056.4]
  assign _T_83014 = _T_83013[4:0]; // @[Modules.scala 43:47:@34057.4]
  assign _T_83015 = $signed(_T_83014); // @[Modules.scala 43:47:@34058.4]
  assign _T_83054 = $signed(_T_54736) + $signed(io_in_171); // @[Modules.scala 43:47:@34099.4]
  assign _T_83055 = _T_83054[4:0]; // @[Modules.scala 43:47:@34100.4]
  assign _T_83056 = $signed(_T_83055); // @[Modules.scala 43:47:@34101.4]
  assign _T_83084 = $signed(_T_54774) + $signed(io_in_183); // @[Modules.scala 43:47:@34132.4]
  assign _T_83085 = _T_83084[4:0]; // @[Modules.scala 43:47:@34133.4]
  assign _T_83086 = $signed(_T_83085); // @[Modules.scala 43:47:@34134.4]
  assign _T_83197 = $signed(io_in_228) - $signed(io_in_229); // @[Modules.scala 40:46:@34257.4]
  assign _T_83198 = _T_83197[4:0]; // @[Modules.scala 40:46:@34258.4]
  assign _T_83199 = $signed(_T_83198); // @[Modules.scala 40:46:@34259.4]
  assign _T_83241 = $signed(_T_54967) + $signed(io_in_245); // @[Modules.scala 43:47:@34304.4]
  assign _T_83242 = _T_83241[4:0]; // @[Modules.scala 43:47:@34305.4]
  assign _T_83243 = $signed(_T_83242); // @[Modules.scala 43:47:@34306.4]
  assign _T_83294 = $signed(io_in_266) - $signed(io_in_267); // @[Modules.scala 40:46:@34363.4]
  assign _T_83295 = _T_83294[4:0]; // @[Modules.scala 40:46:@34364.4]
  assign _T_83296 = $signed(_T_83295); // @[Modules.scala 40:46:@34365.4]
  assign _T_83399 = $signed(io_in_304) - $signed(io_in_305); // @[Modules.scala 40:46:@34475.4]
  assign _T_83400 = _T_83399[4:0]; // @[Modules.scala 40:46:@34476.4]
  assign _T_83401 = $signed(_T_83400); // @[Modules.scala 40:46:@34477.4]
  assign _T_83415 = $signed(io_in_312) - $signed(io_in_313); // @[Modules.scala 40:46:@34494.4]
  assign _T_83416 = _T_83415[4:0]; // @[Modules.scala 40:46:@34495.4]
  assign _T_83417 = $signed(_T_83416); // @[Modules.scala 40:46:@34496.4]
  assign _T_83443 = $signed(_T_55221) + $signed(io_in_321); // @[Modules.scala 43:47:@34522.4]
  assign _T_83444 = _T_83443[4:0]; // @[Modules.scala 43:47:@34523.4]
  assign _T_83445 = $signed(_T_83444); // @[Modules.scala 43:47:@34524.4]
  assign _T_83509 = $signed(_T_64702) + $signed(io_in_349); // @[Modules.scala 43:47:@34596.4]
  assign _T_83510 = _T_83509[4:0]; // @[Modules.scala 43:47:@34597.4]
  assign _T_83511 = $signed(_T_83510); // @[Modules.scala 43:47:@34598.4]
  assign _T_83588 = $signed(io_in_382) - $signed(io_in_383); // @[Modules.scala 40:46:@34685.4]
  assign _T_83589 = _T_83588[4:0]; // @[Modules.scala 40:46:@34686.4]
  assign _T_83590 = $signed(_T_83589); // @[Modules.scala 40:46:@34687.4]
  assign _T_83635 = $signed(io_in_400) - $signed(io_in_401); // @[Modules.scala 40:46:@34736.4]
  assign _T_83636 = _T_83635[4:0]; // @[Modules.scala 40:46:@34737.4]
  assign _T_83637 = $signed(_T_83636); // @[Modules.scala 40:46:@34738.4]
  assign _T_83765 = $signed(io_in_452) - $signed(io_in_453); // @[Modules.scala 40:46:@34879.4]
  assign _T_83766 = _T_83765[4:0]; // @[Modules.scala 40:46:@34880.4]
  assign _T_83767 = $signed(_T_83766); // @[Modules.scala 40:46:@34881.4]
  assign _T_83858 = $signed(io_in_490) - $signed(io_in_491); // @[Modules.scala 40:46:@34982.4]
  assign _T_83859 = _T_83858[4:0]; // @[Modules.scala 40:46:@34983.4]
  assign _T_83860 = $signed(_T_83859); // @[Modules.scala 40:46:@34984.4]
  assign _T_84008 = $signed(_T_55814) + $signed(io_in_567); // @[Modules.scala 43:47:@35161.4]
  assign _T_84009 = _T_84008[4:0]; // @[Modules.scala 43:47:@35162.4]
  assign _T_84010 = $signed(_T_84009); // @[Modules.scala 43:47:@35163.4]
  assign _T_84067 = $signed(io_in_600) - $signed(io_in_601); // @[Modules.scala 40:46:@35235.4]
  assign _T_84068 = _T_84067[4:0]; // @[Modules.scala 40:46:@35236.4]
  assign _T_84069 = $signed(_T_84068); // @[Modules.scala 40:46:@35237.4]
  assign _T_84079 = $signed(io_in_608) - $signed(io_in_609); // @[Modules.scala 40:46:@35251.4]
  assign _T_84080 = _T_84079[4:0]; // @[Modules.scala 40:46:@35252.4]
  assign _T_84081 = $signed(_T_84080); // @[Modules.scala 40:46:@35253.4]
  assign _T_84086 = $signed(_T_55936) + $signed(io_in_611); // @[Modules.scala 43:47:@35258.4]
  assign _T_84087 = _T_84086[4:0]; // @[Modules.scala 43:47:@35259.4]
  assign _T_84088 = $signed(_T_84087); // @[Modules.scala 43:47:@35260.4]
  assign _T_84151 = $signed(_T_59094) + $signed(io_in_641); // @[Modules.scala 43:47:@35333.4]
  assign _T_84152 = _T_84151[4:0]; // @[Modules.scala 43:47:@35334.4]
  assign _T_84153 = $signed(_T_84152); // @[Modules.scala 43:47:@35335.4]
  assign _T_84261 = $signed(_T_59208) + $signed(io_in_693); // @[Modules.scala 43:47:@35461.4]
  assign _T_84262 = _T_84261[4:0]; // @[Modules.scala 43:47:@35462.4]
  assign _T_84263 = $signed(_T_84262); // @[Modules.scala 43:47:@35463.4]
  assign _T_84264 = $signed(io_in_694) - $signed(io_in_695); // @[Modules.scala 40:46:@35465.4]
  assign _T_84265 = _T_84264[4:0]; // @[Modules.scala 40:46:@35466.4]
  assign _T_84266 = $signed(_T_84265); // @[Modules.scala 40:46:@35467.4]
  assign _T_84293 = $signed(io_in_708) - $signed(io_in_709); // @[Modules.scala 40:46:@35499.4]
  assign _T_84294 = _T_84293[4:0]; // @[Modules.scala 40:46:@35500.4]
  assign _T_84295 = $signed(_T_84294); // @[Modules.scala 40:46:@35501.4]
  assign _T_84303 = $signed(io_in_712) - $signed(io_in_713); // @[Modules.scala 40:46:@35510.4]
  assign _T_84304 = _T_84303[4:0]; // @[Modules.scala 40:46:@35511.4]
  assign _T_84305 = $signed(_T_84304); // @[Modules.scala 40:46:@35512.4]
  assign _T_84317 = $signed(_T_62549) + $signed(io_in_717); // @[Modules.scala 43:47:@35524.4]
  assign _T_84318 = _T_84317[4:0]; // @[Modules.scala 43:47:@35525.4]
  assign _T_84319 = $signed(_T_84318); // @[Modules.scala 43:47:@35526.4]
  assign _T_84345 = $signed(_T_68535) + $signed(io_in_725); // @[Modules.scala 43:47:@35552.4]
  assign _T_84346 = _T_84345[4:0]; // @[Modules.scala 43:47:@35553.4]
  assign _T_84347 = $signed(_T_84346); // @[Modules.scala 43:47:@35554.4]
  assign _T_84355 = $signed(_T_59298) + $signed(io_in_729); // @[Modules.scala 43:47:@35563.4]
  assign _T_84356 = _T_84355[4:0]; // @[Modules.scala 43:47:@35564.4]
  assign _T_84357 = $signed(_T_84356); // @[Modules.scala 43:47:@35565.4]
  assign _T_84430 = $signed(_T_65659) - $signed(io_in_755); // @[Modules.scala 46:47:@35642.4]
  assign _T_84431 = _T_84430[4:0]; // @[Modules.scala 46:47:@35643.4]
  assign _T_84432 = $signed(_T_84431); // @[Modules.scala 46:47:@35644.4]
  assign _T_84436 = $signed(io_in_758) - $signed(io_in_759); // @[Modules.scala 40:46:@35650.4]
  assign _T_84437 = _T_84436[4:0]; // @[Modules.scala 40:46:@35651.4]
  assign _T_84438 = $signed(_T_84437); // @[Modules.scala 40:46:@35652.4]
  assign _T_84450 = $signed(_T_56312) + $signed(io_in_763); // @[Modules.scala 43:47:@35664.4]
  assign _T_84451 = _T_84450[4:0]; // @[Modules.scala 43:47:@35665.4]
  assign _T_84452 = $signed(_T_84451); // @[Modules.scala 43:47:@35666.4]
  assign _T_84472 = $signed(io_in_774) - $signed(io_in_775); // @[Modules.scala 40:46:@35691.4]
  assign _T_84473 = _T_84472[4:0]; // @[Modules.scala 40:46:@35692.4]
  assign _T_84474 = $signed(_T_84473); // @[Modules.scala 40:46:@35693.4]
  assign buffer_9_1 = {{6{_T_82680[4]}},_T_82680}; // @[Modules.scala 32:22:@8.4]
  assign _T_84487 = $signed(buffer_1_0) + $signed(buffer_9_1); // @[Modules.scala 50:57:@35711.4]
  assign _T_84488 = _T_84487[10:0]; // @[Modules.scala 50:57:@35712.4]
  assign buffer_9_392 = $signed(_T_84488); // @[Modules.scala 50:57:@35713.4]
  assign buffer_9_2 = {{6{_T_82687[4]}},_T_82687}; // @[Modules.scala 32:22:@8.4]
  assign _T_84490 = $signed(buffer_9_2) + $signed(buffer_0_3); // @[Modules.scala 50:57:@35715.4]
  assign _T_84491 = _T_84490[10:0]; // @[Modules.scala 50:57:@35716.4]
  assign buffer_9_393 = $signed(_T_84491); // @[Modules.scala 50:57:@35717.4]
  assign _T_84493 = $signed(buffer_3_4) + $signed(buffer_0_5); // @[Modules.scala 50:57:@35719.4]
  assign _T_84494 = _T_84493[10:0]; // @[Modules.scala 50:57:@35720.4]
  assign buffer_9_394 = $signed(_T_84494); // @[Modules.scala 50:57:@35721.4]
  assign buffer_9_9 = {{6{_T_82732[4]}},_T_82732}; // @[Modules.scala 32:22:@8.4]
  assign _T_84499 = $signed(buffer_4_8) + $signed(buffer_9_9); // @[Modules.scala 50:57:@35727.4]
  assign _T_84500 = _T_84499[10:0]; // @[Modules.scala 50:57:@35728.4]
  assign buffer_9_396 = $signed(_T_84500); // @[Modules.scala 50:57:@35729.4]
  assign _T_84505 = $signed(buffer_3_12) + $signed(buffer_1_13); // @[Modules.scala 50:57:@35735.4]
  assign _T_84506 = _T_84505[10:0]; // @[Modules.scala 50:57:@35736.4]
  assign buffer_9_398 = $signed(_T_84506); // @[Modules.scala 50:57:@35737.4]
  assign _T_84520 = $signed(buffer_4_22) + $signed(buffer_1_23); // @[Modules.scala 50:57:@35755.4]
  assign _T_84521 = _T_84520[10:0]; // @[Modules.scala 50:57:@35756.4]
  assign buffer_9_403 = $signed(_T_84521); // @[Modules.scala 50:57:@35757.4]
  assign buffer_9_41 = {{6{_T_82860[4]}},_T_82860}; // @[Modules.scala 32:22:@8.4]
  assign _T_84547 = $signed(buffer_1_40) + $signed(buffer_9_41); // @[Modules.scala 50:57:@35791.4]
  assign _T_84548 = _T_84547[10:0]; // @[Modules.scala 50:57:@35792.4]
  assign buffer_9_412 = $signed(_T_84548); // @[Modules.scala 50:57:@35793.4]
  assign _T_84571 = $signed(buffer_0_56) + $signed(buffer_3_57); // @[Modules.scala 50:57:@35823.4]
  assign _T_84572 = _T_84571[10:0]; // @[Modules.scala 50:57:@35824.4]
  assign buffer_9_420 = $signed(_T_84572); // @[Modules.scala 50:57:@35825.4]
  assign _T_84589 = $signed(buffer_8_68) + $signed(buffer_4_69); // @[Modules.scala 50:57:@35847.4]
  assign _T_84590 = _T_84589[10:0]; // @[Modules.scala 50:57:@35848.4]
  assign buffer_9_426 = $signed(_T_84590); // @[Modules.scala 50:57:@35849.4]
  assign buffer_9_75 = {{6{_T_82998[4]}},_T_82998}; // @[Modules.scala 32:22:@8.4]
  assign _T_84598 = $signed(buffer_0_74) + $signed(buffer_9_75); // @[Modules.scala 50:57:@35859.4]
  assign _T_84599 = _T_84598[10:0]; // @[Modules.scala 50:57:@35860.4]
  assign buffer_9_429 = $signed(_T_84599); // @[Modules.scala 50:57:@35861.4]
  assign _T_84601 = $signed(buffer_7_76) + $signed(buffer_0_77); // @[Modules.scala 50:57:@35863.4]
  assign _T_84602 = _T_84601[10:0]; // @[Modules.scala 50:57:@35864.4]
  assign buffer_9_430 = $signed(_T_84602); // @[Modules.scala 50:57:@35865.4]
  assign buffer_9_78 = {{6{_T_83015[4]}},_T_83015}; // @[Modules.scala 32:22:@8.4]
  assign _T_84604 = $signed(buffer_9_78) + $signed(buffer_2_79); // @[Modules.scala 50:57:@35867.4]
  assign _T_84605 = _T_84604[10:0]; // @[Modules.scala 50:57:@35868.4]
  assign buffer_9_431 = $signed(_T_84605); // @[Modules.scala 50:57:@35869.4]
  assign _T_84607 = $signed(buffer_0_80) + $signed(buffer_5_81); // @[Modules.scala 50:57:@35871.4]
  assign _T_84608 = _T_84607[10:0]; // @[Modules.scala 50:57:@35872.4]
  assign buffer_9_432 = $signed(_T_84608); // @[Modules.scala 50:57:@35873.4]
  assign buffer_9_85 = {{6{_T_83056[4]}},_T_83056}; // @[Modules.scala 32:22:@8.4]
  assign _T_84613 = $signed(buffer_4_84) + $signed(buffer_9_85); // @[Modules.scala 50:57:@35879.4]
  assign _T_84614 = _T_84613[10:0]; // @[Modules.scala 50:57:@35880.4]
  assign buffer_9_434 = $signed(_T_84614); // @[Modules.scala 50:57:@35881.4]
  assign buffer_9_91 = {{6{_T_83086[4]}},_T_83086}; // @[Modules.scala 32:22:@8.4]
  assign _T_84622 = $signed(buffer_3_90) + $signed(buffer_9_91); // @[Modules.scala 50:57:@35891.4]
  assign _T_84623 = _T_84622[10:0]; // @[Modules.scala 50:57:@35892.4]
  assign buffer_9_437 = $signed(_T_84623); // @[Modules.scala 50:57:@35893.4]
  assign _T_84628 = $signed(buffer_0_94) + $signed(buffer_5_95); // @[Modules.scala 50:57:@35899.4]
  assign _T_84629 = _T_84628[10:0]; // @[Modules.scala 50:57:@35900.4]
  assign buffer_9_439 = $signed(_T_84629); // @[Modules.scala 50:57:@35901.4]
  assign _T_84631 = $signed(buffer_1_96) + $signed(buffer_2_97); // @[Modules.scala 50:57:@35903.4]
  assign _T_84632 = _T_84631[10:0]; // @[Modules.scala 50:57:@35904.4]
  assign buffer_9_440 = $signed(_T_84632); // @[Modules.scala 50:57:@35905.4]
  assign _T_84640 = $signed(buffer_4_102) + $signed(buffer_2_103); // @[Modules.scala 50:57:@35915.4]
  assign _T_84641 = _T_84640[10:0]; // @[Modules.scala 50:57:@35916.4]
  assign buffer_9_443 = $signed(_T_84641); // @[Modules.scala 50:57:@35917.4]
  assign _T_84646 = $signed(buffer_1_106) + $signed(buffer_0_107); // @[Modules.scala 50:57:@35923.4]
  assign _T_84647 = _T_84646[10:0]; // @[Modules.scala 50:57:@35924.4]
  assign buffer_9_445 = $signed(_T_84647); // @[Modules.scala 50:57:@35925.4]
  assign _T_84649 = $signed(buffer_7_108) + $signed(buffer_0_109); // @[Modules.scala 50:57:@35927.4]
  assign _T_84650 = _T_84649[10:0]; // @[Modules.scala 50:57:@35928.4]
  assign buffer_9_446 = $signed(_T_84650); // @[Modules.scala 50:57:@35929.4]
  assign _T_84652 = $signed(buffer_0_110) + $signed(buffer_2_111); // @[Modules.scala 50:57:@35931.4]
  assign _T_84653 = _T_84652[10:0]; // @[Modules.scala 50:57:@35932.4]
  assign buffer_9_447 = $signed(_T_84653); // @[Modules.scala 50:57:@35933.4]
  assign _T_84655 = $signed(buffer_1_112) + $signed(buffer_5_113); // @[Modules.scala 50:57:@35935.4]
  assign _T_84656 = _T_84655[10:0]; // @[Modules.scala 50:57:@35936.4]
  assign buffer_9_448 = $signed(_T_84656); // @[Modules.scala 50:57:@35937.4]
  assign buffer_9_114 = {{6{_T_83199[4]}},_T_83199}; // @[Modules.scala 32:22:@8.4]
  assign _T_84658 = $signed(buffer_9_114) + $signed(buffer_8_115); // @[Modules.scala 50:57:@35939.4]
  assign _T_84659 = _T_84658[10:0]; // @[Modules.scala 50:57:@35940.4]
  assign buffer_9_449 = $signed(_T_84659); // @[Modules.scala 50:57:@35941.4]
  assign _T_84664 = $signed(buffer_0_118) + $signed(buffer_3_119); // @[Modules.scala 50:57:@35947.4]
  assign _T_84665 = _T_84664[10:0]; // @[Modules.scala 50:57:@35948.4]
  assign buffer_9_451 = $signed(_T_84665); // @[Modules.scala 50:57:@35949.4]
  assign buffer_9_122 = {{6{_T_83243[4]}},_T_83243}; // @[Modules.scala 32:22:@8.4]
  assign _T_84670 = $signed(buffer_9_122) + $signed(buffer_0_123); // @[Modules.scala 50:57:@35955.4]
  assign _T_84671 = _T_84670[10:0]; // @[Modules.scala 50:57:@35956.4]
  assign buffer_9_453 = $signed(_T_84671); // @[Modules.scala 50:57:@35957.4]
  assign _T_84679 = $signed(buffer_8_128) + $signed(buffer_4_129); // @[Modules.scala 50:57:@35967.4]
  assign _T_84680 = _T_84679[10:0]; // @[Modules.scala 50:57:@35968.4]
  assign buffer_9_456 = $signed(_T_84680); // @[Modules.scala 50:57:@35969.4]
  assign buffer_9_133 = {{6{_T_83296[4]}},_T_83296}; // @[Modules.scala 32:22:@8.4]
  assign _T_84685 = $signed(buffer_0_132) + $signed(buffer_9_133); // @[Modules.scala 50:57:@35975.4]
  assign _T_84686 = _T_84685[10:0]; // @[Modules.scala 50:57:@35976.4]
  assign buffer_9_458 = $signed(_T_84686); // @[Modules.scala 50:57:@35977.4]
  assign _T_84694 = $signed(buffer_0_138) + $signed(buffer_1_139); // @[Modules.scala 50:57:@35987.4]
  assign _T_84695 = _T_84694[10:0]; // @[Modules.scala 50:57:@35988.4]
  assign buffer_9_461 = $signed(_T_84695); // @[Modules.scala 50:57:@35989.4]
  assign _T_84697 = $signed(buffer_3_140) + $signed(buffer_1_141); // @[Modules.scala 50:57:@35991.4]
  assign _T_84698 = _T_84697[10:0]; // @[Modules.scala 50:57:@35992.4]
  assign buffer_9_462 = $signed(_T_84698); // @[Modules.scala 50:57:@35993.4]
  assign _T_84700 = $signed(buffer_3_142) + $signed(buffer_5_143); // @[Modules.scala 50:57:@35995.4]
  assign _T_84701 = _T_84700[10:0]; // @[Modules.scala 50:57:@35996.4]
  assign buffer_9_463 = $signed(_T_84701); // @[Modules.scala 50:57:@35997.4]
  assign _T_84712 = $signed(buffer_6_150) + $signed(buffer_4_151); // @[Modules.scala 50:57:@36011.4]
  assign _T_84713 = _T_84712[10:0]; // @[Modules.scala 50:57:@36012.4]
  assign buffer_9_467 = $signed(_T_84713); // @[Modules.scala 50:57:@36013.4]
  assign buffer_9_152 = {{6{_T_83401[4]}},_T_83401}; // @[Modules.scala 32:22:@8.4]
  assign _T_84715 = $signed(buffer_9_152) + $signed(buffer_5_153); // @[Modules.scala 50:57:@36015.4]
  assign _T_84716 = _T_84715[10:0]; // @[Modules.scala 50:57:@36016.4]
  assign buffer_9_468 = $signed(_T_84716); // @[Modules.scala 50:57:@36017.4]
  assign buffer_9_156 = {{6{_T_83417[4]}},_T_83417}; // @[Modules.scala 32:22:@8.4]
  assign _T_84721 = $signed(buffer_9_156) + $signed(buffer_3_157); // @[Modules.scala 50:57:@36023.4]
  assign _T_84722 = _T_84721[10:0]; // @[Modules.scala 50:57:@36024.4]
  assign buffer_9_470 = $signed(_T_84722); // @[Modules.scala 50:57:@36025.4]
  assign buffer_9_160 = {{6{_T_83445[4]}},_T_83445}; // @[Modules.scala 32:22:@8.4]
  assign _T_84727 = $signed(buffer_9_160) + $signed(buffer_5_161); // @[Modules.scala 50:57:@36031.4]
  assign _T_84728 = _T_84727[10:0]; // @[Modules.scala 50:57:@36032.4]
  assign buffer_9_472 = $signed(_T_84728); // @[Modules.scala 50:57:@36033.4]
  assign buffer_9_174 = {{6{_T_83511[4]}},_T_83511}; // @[Modules.scala 32:22:@8.4]
  assign _T_84748 = $signed(buffer_9_174) + $signed(buffer_0_175); // @[Modules.scala 50:57:@36059.4]
  assign _T_84749 = _T_84748[10:0]; // @[Modules.scala 50:57:@36060.4]
  assign buffer_9_479 = $signed(_T_84749); // @[Modules.scala 50:57:@36061.4]
  assign _T_84751 = $signed(buffer_1_176) + $signed(buffer_0_177); // @[Modules.scala 50:57:@36063.4]
  assign _T_84752 = _T_84751[10:0]; // @[Modules.scala 50:57:@36064.4]
  assign buffer_9_480 = $signed(_T_84752); // @[Modules.scala 50:57:@36065.4]
  assign _T_84754 = $signed(buffer_0_178) + $signed(buffer_2_179); // @[Modules.scala 50:57:@36067.4]
  assign _T_84755 = _T_84754[10:0]; // @[Modules.scala 50:57:@36068.4]
  assign buffer_9_481 = $signed(_T_84755); // @[Modules.scala 50:57:@36069.4]
  assign _T_84766 = $signed(buffer_3_186) + $signed(buffer_5_187); // @[Modules.scala 50:57:@36083.4]
  assign _T_84767 = _T_84766[10:0]; // @[Modules.scala 50:57:@36084.4]
  assign buffer_9_485 = $signed(_T_84767); // @[Modules.scala 50:57:@36085.4]
  assign buffer_9_191 = {{6{_T_83590[4]}},_T_83590}; // @[Modules.scala 32:22:@8.4]
  assign _T_84772 = $signed(buffer_4_190) + $signed(buffer_9_191); // @[Modules.scala 50:57:@36091.4]
  assign _T_84773 = _T_84772[10:0]; // @[Modules.scala 50:57:@36092.4]
  assign buffer_9_487 = $signed(_T_84773); // @[Modules.scala 50:57:@36093.4]
  assign _T_84778 = $signed(buffer_4_194) + $signed(buffer_3_195); // @[Modules.scala 50:57:@36099.4]
  assign _T_84779 = _T_84778[10:0]; // @[Modules.scala 50:57:@36100.4]
  assign buffer_9_489 = $signed(_T_84779); // @[Modules.scala 50:57:@36101.4]
  assign _T_84781 = $signed(buffer_6_196) + $signed(buffer_3_197); // @[Modules.scala 50:57:@36103.4]
  assign _T_84782 = _T_84781[10:0]; // @[Modules.scala 50:57:@36104.4]
  assign buffer_9_490 = $signed(_T_84782); // @[Modules.scala 50:57:@36105.4]
  assign buffer_9_200 = {{6{_T_83637[4]}},_T_83637}; // @[Modules.scala 32:22:@8.4]
  assign _T_84787 = $signed(buffer_9_200) + $signed(buffer_5_201); // @[Modules.scala 50:57:@36111.4]
  assign _T_84788 = _T_84787[10:0]; // @[Modules.scala 50:57:@36112.4]
  assign buffer_9_492 = $signed(_T_84788); // @[Modules.scala 50:57:@36113.4]
  assign _T_84805 = $signed(buffer_2_212) + $signed(buffer_1_213); // @[Modules.scala 50:57:@36135.4]
  assign _T_84806 = _T_84805[10:0]; // @[Modules.scala 50:57:@36136.4]
  assign buffer_9_498 = $signed(_T_84806); // @[Modules.scala 50:57:@36137.4]
  assign _T_84808 = $signed(buffer_5_214) + $signed(buffer_6_215); // @[Modules.scala 50:57:@36139.4]
  assign _T_84809 = _T_84808[10:0]; // @[Modules.scala 50:57:@36140.4]
  assign buffer_9_499 = $signed(_T_84809); // @[Modules.scala 50:57:@36141.4]
  assign _T_84823 = $signed(buffer_0_224) + $signed(buffer_1_225); // @[Modules.scala 50:57:@36159.4]
  assign _T_84824 = _T_84823[10:0]; // @[Modules.scala 50:57:@36160.4]
  assign buffer_9_504 = $signed(_T_84824); // @[Modules.scala 50:57:@36161.4]
  assign buffer_9_226 = {{6{_T_83767[4]}},_T_83767}; // @[Modules.scala 32:22:@8.4]
  assign _T_84826 = $signed(buffer_9_226) + $signed(buffer_1_227); // @[Modules.scala 50:57:@36163.4]
  assign _T_84827 = _T_84826[10:0]; // @[Modules.scala 50:57:@36164.4]
  assign buffer_9_505 = $signed(_T_84827); // @[Modules.scala 50:57:@36165.4]
  assign _T_84829 = $signed(buffer_3_228) + $signed(buffer_6_229); // @[Modules.scala 50:57:@36167.4]
  assign _T_84830 = _T_84829[10:0]; // @[Modules.scala 50:57:@36168.4]
  assign buffer_9_506 = $signed(_T_84830); // @[Modules.scala 50:57:@36169.4]
  assign _T_84835 = $signed(buffer_1_232) + $signed(buffer_5_233); // @[Modules.scala 50:57:@36175.4]
  assign _T_84836 = _T_84835[10:0]; // @[Modules.scala 50:57:@36176.4]
  assign buffer_9_508 = $signed(_T_84836); // @[Modules.scala 50:57:@36177.4]
  assign _T_84847 = $signed(buffer_7_240) + $signed(buffer_2_241); // @[Modules.scala 50:57:@36191.4]
  assign _T_84848 = _T_84847[10:0]; // @[Modules.scala 50:57:@36192.4]
  assign buffer_9_512 = $signed(_T_84848); // @[Modules.scala 50:57:@36193.4]
  assign buffer_9_245 = {{6{_T_83860[4]}},_T_83860}; // @[Modules.scala 32:22:@8.4]
  assign _T_84853 = $signed(buffer_2_244) + $signed(buffer_9_245); // @[Modules.scala 50:57:@36199.4]
  assign _T_84854 = _T_84853[10:0]; // @[Modules.scala 50:57:@36200.4]
  assign buffer_9_514 = $signed(_T_84854); // @[Modules.scala 50:57:@36201.4]
  assign _T_84868 = $signed(buffer_3_254) + $signed(buffer_0_255); // @[Modules.scala 50:57:@36219.4]
  assign _T_84869 = _T_84868[10:0]; // @[Modules.scala 50:57:@36220.4]
  assign buffer_9_519 = $signed(_T_84869); // @[Modules.scala 50:57:@36221.4]
  assign _T_84889 = $signed(buffer_1_268) + $signed(buffer_5_269); // @[Modules.scala 50:57:@36247.4]
  assign _T_84890 = _T_84889[10:0]; // @[Modules.scala 50:57:@36248.4]
  assign buffer_9_526 = $signed(_T_84890); // @[Modules.scala 50:57:@36249.4]
  assign buffer_9_283 = {{6{_T_84010[4]}},_T_84010}; // @[Modules.scala 32:22:@8.4]
  assign _T_84910 = $signed(buffer_1_282) + $signed(buffer_9_283); // @[Modules.scala 50:57:@36275.4]
  assign _T_84911 = _T_84910[10:0]; // @[Modules.scala 50:57:@36276.4]
  assign buffer_9_533 = $signed(_T_84911); // @[Modules.scala 50:57:@36277.4]
  assign _T_84913 = $signed(buffer_8_284) + $signed(buffer_1_285); // @[Modules.scala 50:57:@36279.4]
  assign _T_84914 = _T_84913[10:0]; // @[Modules.scala 50:57:@36280.4]
  assign buffer_9_534 = $signed(_T_84914); // @[Modules.scala 50:57:@36281.4]
  assign _T_84916 = $signed(buffer_3_286) + $signed(buffer_1_287); // @[Modules.scala 50:57:@36283.4]
  assign _T_84917 = _T_84916[10:0]; // @[Modules.scala 50:57:@36284.4]
  assign buffer_9_535 = $signed(_T_84917); // @[Modules.scala 50:57:@36285.4]
  assign _T_84934 = $signed(buffer_1_298) + $signed(buffer_2_299); // @[Modules.scala 50:57:@36307.4]
  assign _T_84935 = _T_84934[10:0]; // @[Modules.scala 50:57:@36308.4]
  assign buffer_9_541 = $signed(_T_84935); // @[Modules.scala 50:57:@36309.4]
  assign buffer_9_300 = {{6{_T_84069[4]}},_T_84069}; // @[Modules.scala 32:22:@8.4]
  assign _T_84937 = $signed(buffer_9_300) + $signed(buffer_0_301); // @[Modules.scala 50:57:@36311.4]
  assign _T_84938 = _T_84937[10:0]; // @[Modules.scala 50:57:@36312.4]
  assign buffer_9_542 = $signed(_T_84938); // @[Modules.scala 50:57:@36313.4]
  assign buffer_9_304 = {{6{_T_84081[4]}},_T_84081}; // @[Modules.scala 32:22:@8.4]
  assign buffer_9_305 = {{6{_T_84088[4]}},_T_84088}; // @[Modules.scala 32:22:@8.4]
  assign _T_84943 = $signed(buffer_9_304) + $signed(buffer_9_305); // @[Modules.scala 50:57:@36319.4]
  assign _T_84944 = _T_84943[10:0]; // @[Modules.scala 50:57:@36320.4]
  assign buffer_9_544 = $signed(_T_84944); // @[Modules.scala 50:57:@36321.4]
  assign _T_84955 = $signed(buffer_1_312) + $signed(buffer_5_313); // @[Modules.scala 50:57:@36335.4]
  assign _T_84956 = _T_84955[10:0]; // @[Modules.scala 50:57:@36336.4]
  assign buffer_9_548 = $signed(_T_84956); // @[Modules.scala 50:57:@36337.4]
  assign _T_84961 = $signed(buffer_4_316) + $signed(buffer_0_317); // @[Modules.scala 50:57:@36343.4]
  assign _T_84962 = _T_84961[10:0]; // @[Modules.scala 50:57:@36344.4]
  assign buffer_9_550 = $signed(_T_84962); // @[Modules.scala 50:57:@36345.4]
  assign _T_84964 = $signed(buffer_1_318) + $signed(buffer_0_319); // @[Modules.scala 50:57:@36347.4]
  assign _T_84965 = _T_84964[10:0]; // @[Modules.scala 50:57:@36348.4]
  assign buffer_9_551 = $signed(_T_84965); // @[Modules.scala 50:57:@36349.4]
  assign buffer_9_320 = {{6{_T_84153[4]}},_T_84153}; // @[Modules.scala 32:22:@8.4]
  assign _T_84967 = $signed(buffer_9_320) + $signed(buffer_3_321); // @[Modules.scala 50:57:@36351.4]
  assign _T_84968 = _T_84967[10:0]; // @[Modules.scala 50:57:@36352.4]
  assign buffer_9_552 = $signed(_T_84968); // @[Modules.scala 50:57:@36353.4]
  assign _T_84976 = $signed(buffer_1_326) + $signed(buffer_8_327); // @[Modules.scala 50:57:@36363.4]
  assign _T_84977 = _T_84976[10:0]; // @[Modules.scala 50:57:@36364.4]
  assign buffer_9_555 = $signed(_T_84977); // @[Modules.scala 50:57:@36365.4]
  assign _T_84985 = $signed(buffer_5_332) + $signed(buffer_1_333); // @[Modules.scala 50:57:@36375.4]
  assign _T_84986 = _T_84985[10:0]; // @[Modules.scala 50:57:@36376.4]
  assign buffer_9_558 = $signed(_T_84986); // @[Modules.scala 50:57:@36377.4]
  assign buffer_9_346 = {{6{_T_84263[4]}},_T_84263}; // @[Modules.scala 32:22:@8.4]
  assign buffer_9_347 = {{6{_T_84266[4]}},_T_84266}; // @[Modules.scala 32:22:@8.4]
  assign _T_85006 = $signed(buffer_9_346) + $signed(buffer_9_347); // @[Modules.scala 50:57:@36403.4]
  assign _T_85007 = _T_85006[10:0]; // @[Modules.scala 50:57:@36404.4]
  assign buffer_9_565 = $signed(_T_85007); // @[Modules.scala 50:57:@36405.4]
  assign _T_85009 = $signed(buffer_0_348) + $signed(buffer_3_349); // @[Modules.scala 50:57:@36407.4]
  assign _T_85010 = _T_85009[10:0]; // @[Modules.scala 50:57:@36408.4]
  assign buffer_9_566 = $signed(_T_85010); // @[Modules.scala 50:57:@36409.4]
  assign _T_85012 = $signed(buffer_5_350) + $signed(buffer_0_351); // @[Modules.scala 50:57:@36411.4]
  assign _T_85013 = _T_85012[10:0]; // @[Modules.scala 50:57:@36412.4]
  assign buffer_9_567 = $signed(_T_85013); // @[Modules.scala 50:57:@36413.4]
  assign buffer_9_354 = {{6{_T_84295[4]}},_T_84295}; // @[Modules.scala 32:22:@8.4]
  assign _T_85018 = $signed(buffer_9_354) + $signed(buffer_2_355); // @[Modules.scala 50:57:@36419.4]
  assign _T_85019 = _T_85018[10:0]; // @[Modules.scala 50:57:@36420.4]
  assign buffer_9_569 = $signed(_T_85019); // @[Modules.scala 50:57:@36421.4]
  assign buffer_9_356 = {{6{_T_84305[4]}},_T_84305}; // @[Modules.scala 32:22:@8.4]
  assign _T_85021 = $signed(buffer_9_356) + $signed(buffer_2_357); // @[Modules.scala 50:57:@36423.4]
  assign _T_85022 = _T_85021[10:0]; // @[Modules.scala 50:57:@36424.4]
  assign buffer_9_570 = $signed(_T_85022); // @[Modules.scala 50:57:@36425.4]
  assign buffer_9_358 = {{6{_T_84319[4]}},_T_84319}; // @[Modules.scala 32:22:@8.4]
  assign _T_85024 = $signed(buffer_9_358) + $signed(buffer_6_359); // @[Modules.scala 50:57:@36427.4]
  assign _T_85025 = _T_85024[10:0]; // @[Modules.scala 50:57:@36428.4]
  assign buffer_9_571 = $signed(_T_85025); // @[Modules.scala 50:57:@36429.4]
  assign buffer_9_362 = {{6{_T_84347[4]}},_T_84347}; // @[Modules.scala 32:22:@8.4]
  assign _T_85030 = $signed(buffer_9_362) + $signed(buffer_1_363); // @[Modules.scala 50:57:@36435.4]
  assign _T_85031 = _T_85030[10:0]; // @[Modules.scala 50:57:@36436.4]
  assign buffer_9_573 = $signed(_T_85031); // @[Modules.scala 50:57:@36437.4]
  assign buffer_9_364 = {{6{_T_84357[4]}},_T_84357}; // @[Modules.scala 32:22:@8.4]
  assign _T_85033 = $signed(buffer_9_364) + $signed(buffer_3_365); // @[Modules.scala 50:57:@36439.4]
  assign _T_85034 = _T_85033[10:0]; // @[Modules.scala 50:57:@36440.4]
  assign buffer_9_574 = $signed(_T_85034); // @[Modules.scala 50:57:@36441.4]
  assign _T_85045 = $signed(buffer_0_372) + $signed(buffer_3_373); // @[Modules.scala 50:57:@36455.4]
  assign _T_85046 = _T_85045[10:0]; // @[Modules.scala 50:57:@36456.4]
  assign buffer_9_578 = $signed(_T_85046); // @[Modules.scala 50:57:@36457.4]
  assign _T_85048 = $signed(buffer_0_374) + $signed(buffer_2_375); // @[Modules.scala 50:57:@36459.4]
  assign _T_85049 = _T_85048[10:0]; // @[Modules.scala 50:57:@36460.4]
  assign buffer_9_579 = $signed(_T_85049); // @[Modules.scala 50:57:@36461.4]
  assign buffer_9_377 = {{6{_T_84432[4]}},_T_84432}; // @[Modules.scala 32:22:@8.4]
  assign _T_85051 = $signed(buffer_0_376) + $signed(buffer_9_377); // @[Modules.scala 50:57:@36463.4]
  assign _T_85052 = _T_85051[10:0]; // @[Modules.scala 50:57:@36464.4]
  assign buffer_9_580 = $signed(_T_85052); // @[Modules.scala 50:57:@36465.4]
  assign buffer_9_379 = {{6{_T_84438[4]}},_T_84438}; // @[Modules.scala 32:22:@8.4]
  assign _T_85054 = $signed(buffer_3_378) + $signed(buffer_9_379); // @[Modules.scala 50:57:@36467.4]
  assign _T_85055 = _T_85054[10:0]; // @[Modules.scala 50:57:@36468.4]
  assign buffer_9_581 = $signed(_T_85055); // @[Modules.scala 50:57:@36469.4]
  assign buffer_9_381 = {{6{_T_84452[4]}},_T_84452}; // @[Modules.scala 32:22:@8.4]
  assign _T_85057 = $signed(buffer_5_380) + $signed(buffer_9_381); // @[Modules.scala 50:57:@36471.4]
  assign _T_85058 = _T_85057[10:0]; // @[Modules.scala 50:57:@36472.4]
  assign buffer_9_582 = $signed(_T_85058); // @[Modules.scala 50:57:@36473.4]
  assign _T_85060 = $signed(buffer_3_382) + $signed(buffer_4_383); // @[Modules.scala 50:57:@36475.4]
  assign _T_85061 = _T_85060[10:0]; // @[Modules.scala 50:57:@36476.4]
  assign buffer_9_583 = $signed(_T_85061); // @[Modules.scala 50:57:@36477.4]
  assign buffer_9_387 = {{6{_T_84474[4]}},_T_84474}; // @[Modules.scala 32:22:@8.4]
  assign _T_85066 = $signed(buffer_3_386) + $signed(buffer_9_387); // @[Modules.scala 50:57:@36483.4]
  assign _T_85067 = _T_85066[10:0]; // @[Modules.scala 50:57:@36484.4]
  assign buffer_9_585 = $signed(_T_85067); // @[Modules.scala 50:57:@36485.4]
  assign _T_85075 = $signed(buffer_9_392) + $signed(buffer_9_393); // @[Modules.scala 53:83:@36495.4]
  assign _T_85076 = _T_85075[10:0]; // @[Modules.scala 53:83:@36496.4]
  assign buffer_9_588 = $signed(_T_85076); // @[Modules.scala 53:83:@36497.4]
  assign _T_85078 = $signed(buffer_9_394) + $signed(buffer_0_395); // @[Modules.scala 53:83:@36499.4]
  assign _T_85079 = _T_85078[10:0]; // @[Modules.scala 53:83:@36500.4]
  assign buffer_9_589 = $signed(_T_85079); // @[Modules.scala 53:83:@36501.4]
  assign _T_85081 = $signed(buffer_9_396) + $signed(buffer_5_397); // @[Modules.scala 53:83:@36503.4]
  assign _T_85082 = _T_85081[10:0]; // @[Modules.scala 53:83:@36504.4]
  assign buffer_9_590 = $signed(_T_85082); // @[Modules.scala 53:83:@36505.4]
  assign _T_85084 = $signed(buffer_9_398) + $signed(buffer_3_399); // @[Modules.scala 53:83:@36507.4]
  assign _T_85085 = _T_85084[10:0]; // @[Modules.scala 53:83:@36508.4]
  assign buffer_9_591 = $signed(_T_85085); // @[Modules.scala 53:83:@36509.4]
  assign _T_85090 = $signed(buffer_1_402) + $signed(buffer_9_403); // @[Modules.scala 53:83:@36515.4]
  assign _T_85091 = _T_85090[10:0]; // @[Modules.scala 53:83:@36516.4]
  assign buffer_9_593 = $signed(_T_85091); // @[Modules.scala 53:83:@36517.4]
  assign _T_85093 = $signed(buffer_1_404) + $signed(buffer_6_405); // @[Modules.scala 53:83:@36519.4]
  assign _T_85094 = _T_85093[10:0]; // @[Modules.scala 53:83:@36520.4]
  assign buffer_9_594 = $signed(_T_85094); // @[Modules.scala 53:83:@36521.4]
  assign _T_85096 = $signed(buffer_2_406) + $signed(buffer_1_407); // @[Modules.scala 53:83:@36523.4]
  assign _T_85097 = _T_85096[10:0]; // @[Modules.scala 53:83:@36524.4]
  assign buffer_9_595 = $signed(_T_85097); // @[Modules.scala 53:83:@36525.4]
  assign _T_85105 = $signed(buffer_9_412) + $signed(buffer_1_413); // @[Modules.scala 53:83:@36535.4]
  assign _T_85106 = _T_85105[10:0]; // @[Modules.scala 53:83:@36536.4]
  assign buffer_9_598 = $signed(_T_85106); // @[Modules.scala 53:83:@36537.4]
  assign _T_85117 = $signed(buffer_9_420) + $signed(buffer_7_421); // @[Modules.scala 53:83:@36551.4]
  assign _T_85118 = _T_85117[10:0]; // @[Modules.scala 53:83:@36552.4]
  assign buffer_9_602 = $signed(_T_85118); // @[Modules.scala 53:83:@36553.4]
  assign _T_85123 = $signed(buffer_1_424) + $signed(buffer_4_425); // @[Modules.scala 53:83:@36559.4]
  assign _T_85124 = _T_85123[10:0]; // @[Modules.scala 53:83:@36560.4]
  assign buffer_9_604 = $signed(_T_85124); // @[Modules.scala 53:83:@36561.4]
  assign _T_85126 = $signed(buffer_9_426) + $signed(buffer_5_427); // @[Modules.scala 53:83:@36563.4]
  assign _T_85127 = _T_85126[10:0]; // @[Modules.scala 53:83:@36564.4]
  assign buffer_9_605 = $signed(_T_85127); // @[Modules.scala 53:83:@36565.4]
  assign _T_85129 = $signed(buffer_4_428) + $signed(buffer_9_429); // @[Modules.scala 53:83:@36567.4]
  assign _T_85130 = _T_85129[10:0]; // @[Modules.scala 53:83:@36568.4]
  assign buffer_9_606 = $signed(_T_85130); // @[Modules.scala 53:83:@36569.4]
  assign _T_85132 = $signed(buffer_9_430) + $signed(buffer_9_431); // @[Modules.scala 53:83:@36571.4]
  assign _T_85133 = _T_85132[10:0]; // @[Modules.scala 53:83:@36572.4]
  assign buffer_9_607 = $signed(_T_85133); // @[Modules.scala 53:83:@36573.4]
  assign _T_85135 = $signed(buffer_9_432) + $signed(buffer_1_433); // @[Modules.scala 53:83:@36575.4]
  assign _T_85136 = _T_85135[10:0]; // @[Modules.scala 53:83:@36576.4]
  assign buffer_9_608 = $signed(_T_85136); // @[Modules.scala 53:83:@36577.4]
  assign _T_85138 = $signed(buffer_9_434) + $signed(buffer_1_435); // @[Modules.scala 53:83:@36579.4]
  assign _T_85139 = _T_85138[10:0]; // @[Modules.scala 53:83:@36580.4]
  assign buffer_9_609 = $signed(_T_85139); // @[Modules.scala 53:83:@36581.4]
  assign _T_85141 = $signed(buffer_7_436) + $signed(buffer_9_437); // @[Modules.scala 53:83:@36583.4]
  assign _T_85142 = _T_85141[10:0]; // @[Modules.scala 53:83:@36584.4]
  assign buffer_9_610 = $signed(_T_85142); // @[Modules.scala 53:83:@36585.4]
  assign _T_85144 = $signed(buffer_3_438) + $signed(buffer_9_439); // @[Modules.scala 53:83:@36587.4]
  assign _T_85145 = _T_85144[10:0]; // @[Modules.scala 53:83:@36588.4]
  assign buffer_9_611 = $signed(_T_85145); // @[Modules.scala 53:83:@36589.4]
  assign _T_85147 = $signed(buffer_9_440) + $signed(buffer_1_441); // @[Modules.scala 53:83:@36591.4]
  assign _T_85148 = _T_85147[10:0]; // @[Modules.scala 53:83:@36592.4]
  assign buffer_9_612 = $signed(_T_85148); // @[Modules.scala 53:83:@36593.4]
  assign _T_85150 = $signed(buffer_5_442) + $signed(buffer_9_443); // @[Modules.scala 53:83:@36595.4]
  assign _T_85151 = _T_85150[10:0]; // @[Modules.scala 53:83:@36596.4]
  assign buffer_9_613 = $signed(_T_85151); // @[Modules.scala 53:83:@36597.4]
  assign _T_85153 = $signed(buffer_2_444) + $signed(buffer_9_445); // @[Modules.scala 53:83:@36599.4]
  assign _T_85154 = _T_85153[10:0]; // @[Modules.scala 53:83:@36600.4]
  assign buffer_9_614 = $signed(_T_85154); // @[Modules.scala 53:83:@36601.4]
  assign _T_85156 = $signed(buffer_9_446) + $signed(buffer_9_447); // @[Modules.scala 53:83:@36603.4]
  assign _T_85157 = _T_85156[10:0]; // @[Modules.scala 53:83:@36604.4]
  assign buffer_9_615 = $signed(_T_85157); // @[Modules.scala 53:83:@36605.4]
  assign _T_85159 = $signed(buffer_9_448) + $signed(buffer_9_449); // @[Modules.scala 53:83:@36607.4]
  assign _T_85160 = _T_85159[10:0]; // @[Modules.scala 53:83:@36608.4]
  assign buffer_9_616 = $signed(_T_85160); // @[Modules.scala 53:83:@36609.4]
  assign _T_85162 = $signed(buffer_7_450) + $signed(buffer_9_451); // @[Modules.scala 53:83:@36611.4]
  assign _T_85163 = _T_85162[10:0]; // @[Modules.scala 53:83:@36612.4]
  assign buffer_9_617 = $signed(_T_85163); // @[Modules.scala 53:83:@36613.4]
  assign _T_85165 = $signed(buffer_4_452) + $signed(buffer_9_453); // @[Modules.scala 53:83:@36615.4]
  assign _T_85166 = _T_85165[10:0]; // @[Modules.scala 53:83:@36616.4]
  assign buffer_9_618 = $signed(_T_85166); // @[Modules.scala 53:83:@36617.4]
  assign _T_85171 = $signed(buffer_9_456) + $signed(buffer_1_457); // @[Modules.scala 53:83:@36623.4]
  assign _T_85172 = _T_85171[10:0]; // @[Modules.scala 53:83:@36624.4]
  assign buffer_9_620 = $signed(_T_85172); // @[Modules.scala 53:83:@36625.4]
  assign _T_85174 = $signed(buffer_9_458) + $signed(buffer_0_459); // @[Modules.scala 53:83:@36627.4]
  assign _T_85175 = _T_85174[10:0]; // @[Modules.scala 53:83:@36628.4]
  assign buffer_9_621 = $signed(_T_85175); // @[Modules.scala 53:83:@36629.4]
  assign _T_85177 = $signed(buffer_0_460) + $signed(buffer_9_461); // @[Modules.scala 53:83:@36631.4]
  assign _T_85178 = _T_85177[10:0]; // @[Modules.scala 53:83:@36632.4]
  assign buffer_9_622 = $signed(_T_85178); // @[Modules.scala 53:83:@36633.4]
  assign _T_85180 = $signed(buffer_9_462) + $signed(buffer_9_463); // @[Modules.scala 53:83:@36635.4]
  assign _T_85181 = _T_85180[10:0]; // @[Modules.scala 53:83:@36636.4]
  assign buffer_9_623 = $signed(_T_85181); // @[Modules.scala 53:83:@36637.4]
  assign _T_85186 = $signed(buffer_0_466) + $signed(buffer_9_467); // @[Modules.scala 53:83:@36643.4]
  assign _T_85187 = _T_85186[10:0]; // @[Modules.scala 53:83:@36644.4]
  assign buffer_9_625 = $signed(_T_85187); // @[Modules.scala 53:83:@36645.4]
  assign _T_85189 = $signed(buffer_9_468) + $signed(buffer_8_469); // @[Modules.scala 53:83:@36647.4]
  assign _T_85190 = _T_85189[10:0]; // @[Modules.scala 53:83:@36648.4]
  assign buffer_9_626 = $signed(_T_85190); // @[Modules.scala 53:83:@36649.4]
  assign _T_85192 = $signed(buffer_9_470) + $signed(buffer_3_471); // @[Modules.scala 53:83:@36651.4]
  assign _T_85193 = _T_85192[10:0]; // @[Modules.scala 53:83:@36652.4]
  assign buffer_9_627 = $signed(_T_85193); // @[Modules.scala 53:83:@36653.4]
  assign _T_85195 = $signed(buffer_9_472) + $signed(buffer_6_473); // @[Modules.scala 53:83:@36655.4]
  assign _T_85196 = _T_85195[10:0]; // @[Modules.scala 53:83:@36656.4]
  assign buffer_9_628 = $signed(_T_85196); // @[Modules.scala 53:83:@36657.4]
  assign _T_85198 = $signed(buffer_5_474) + $signed(buffer_1_475); // @[Modules.scala 53:83:@36659.4]
  assign _T_85199 = _T_85198[10:0]; // @[Modules.scala 53:83:@36660.4]
  assign buffer_9_629 = $signed(_T_85199); // @[Modules.scala 53:83:@36661.4]
  assign _T_85204 = $signed(buffer_3_478) + $signed(buffer_9_479); // @[Modules.scala 53:83:@36667.4]
  assign _T_85205 = _T_85204[10:0]; // @[Modules.scala 53:83:@36668.4]
  assign buffer_9_631 = $signed(_T_85205); // @[Modules.scala 53:83:@36669.4]
  assign _T_85207 = $signed(buffer_9_480) + $signed(buffer_9_481); // @[Modules.scala 53:83:@36671.4]
  assign _T_85208 = _T_85207[10:0]; // @[Modules.scala 53:83:@36672.4]
  assign buffer_9_632 = $signed(_T_85208); // @[Modules.scala 53:83:@36673.4]
  assign _T_85213 = $signed(buffer_3_484) + $signed(buffer_9_485); // @[Modules.scala 53:83:@36679.4]
  assign _T_85214 = _T_85213[10:0]; // @[Modules.scala 53:83:@36680.4]
  assign buffer_9_634 = $signed(_T_85214); // @[Modules.scala 53:83:@36681.4]
  assign _T_85216 = $signed(buffer_0_486) + $signed(buffer_9_487); // @[Modules.scala 53:83:@36683.4]
  assign _T_85217 = _T_85216[10:0]; // @[Modules.scala 53:83:@36684.4]
  assign buffer_9_635 = $signed(_T_85217); // @[Modules.scala 53:83:@36685.4]
  assign _T_85219 = $signed(buffer_3_488) + $signed(buffer_9_489); // @[Modules.scala 53:83:@36687.4]
  assign _T_85220 = _T_85219[10:0]; // @[Modules.scala 53:83:@36688.4]
  assign buffer_9_636 = $signed(_T_85220); // @[Modules.scala 53:83:@36689.4]
  assign _T_85222 = $signed(buffer_9_490) + $signed(buffer_3_491); // @[Modules.scala 53:83:@36691.4]
  assign _T_85223 = _T_85222[10:0]; // @[Modules.scala 53:83:@36692.4]
  assign buffer_9_637 = $signed(_T_85223); // @[Modules.scala 53:83:@36693.4]
  assign _T_85225 = $signed(buffer_9_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@36695.4]
  assign _T_85226 = _T_85225[10:0]; // @[Modules.scala 53:83:@36696.4]
  assign buffer_9_638 = $signed(_T_85226); // @[Modules.scala 53:83:@36697.4]
  assign _T_85231 = $signed(buffer_3_496) + $signed(buffer_2_497); // @[Modules.scala 53:83:@36703.4]
  assign _T_85232 = _T_85231[10:0]; // @[Modules.scala 53:83:@36704.4]
  assign buffer_9_640 = $signed(_T_85232); // @[Modules.scala 53:83:@36705.4]
  assign _T_85234 = $signed(buffer_9_498) + $signed(buffer_9_499); // @[Modules.scala 53:83:@36707.4]
  assign _T_85235 = _T_85234[10:0]; // @[Modules.scala 53:83:@36708.4]
  assign buffer_9_641 = $signed(_T_85235); // @[Modules.scala 53:83:@36709.4]
  assign _T_85243 = $signed(buffer_9_504) + $signed(buffer_9_505); // @[Modules.scala 53:83:@36719.4]
  assign _T_85244 = _T_85243[10:0]; // @[Modules.scala 53:83:@36720.4]
  assign buffer_9_644 = $signed(_T_85244); // @[Modules.scala 53:83:@36721.4]
  assign _T_85246 = $signed(buffer_9_506) + $signed(buffer_2_507); // @[Modules.scala 53:83:@36723.4]
  assign _T_85247 = _T_85246[10:0]; // @[Modules.scala 53:83:@36724.4]
  assign buffer_9_645 = $signed(_T_85247); // @[Modules.scala 53:83:@36725.4]
  assign _T_85249 = $signed(buffer_9_508) + $signed(buffer_5_509); // @[Modules.scala 53:83:@36727.4]
  assign _T_85250 = _T_85249[10:0]; // @[Modules.scala 53:83:@36728.4]
  assign buffer_9_646 = $signed(_T_85250); // @[Modules.scala 53:83:@36729.4]
  assign _T_85255 = $signed(buffer_9_512) + $signed(buffer_2_513); // @[Modules.scala 53:83:@36735.4]
  assign _T_85256 = _T_85255[10:0]; // @[Modules.scala 53:83:@36736.4]
  assign buffer_9_648 = $signed(_T_85256); // @[Modules.scala 53:83:@36737.4]
  assign _T_85258 = $signed(buffer_9_514) + $signed(buffer_1_515); // @[Modules.scala 53:83:@36739.4]
  assign _T_85259 = _T_85258[10:0]; // @[Modules.scala 53:83:@36740.4]
  assign buffer_9_649 = $signed(_T_85259); // @[Modules.scala 53:83:@36741.4]
  assign _T_85264 = $signed(buffer_1_518) + $signed(buffer_9_519); // @[Modules.scala 53:83:@36747.4]
  assign _T_85265 = _T_85264[10:0]; // @[Modules.scala 53:83:@36748.4]
  assign buffer_9_651 = $signed(_T_85265); // @[Modules.scala 53:83:@36749.4]
  assign _T_85276 = $signed(buffer_9_526) + $signed(buffer_1_527); // @[Modules.scala 53:83:@36763.4]
  assign _T_85277 = _T_85276[10:0]; // @[Modules.scala 53:83:@36764.4]
  assign buffer_9_655 = $signed(_T_85277); // @[Modules.scala 53:83:@36765.4]
  assign _T_85285 = $signed(buffer_8_532) + $signed(buffer_9_533); // @[Modules.scala 53:83:@36775.4]
  assign _T_85286 = _T_85285[10:0]; // @[Modules.scala 53:83:@36776.4]
  assign buffer_9_658 = $signed(_T_85286); // @[Modules.scala 53:83:@36777.4]
  assign _T_85288 = $signed(buffer_9_534) + $signed(buffer_9_535); // @[Modules.scala 53:83:@36779.4]
  assign _T_85289 = _T_85288[10:0]; // @[Modules.scala 53:83:@36780.4]
  assign buffer_9_659 = $signed(_T_85289); // @[Modules.scala 53:83:@36781.4]
  assign _T_85294 = $signed(buffer_8_538) + $signed(buffer_4_539); // @[Modules.scala 53:83:@36787.4]
  assign _T_85295 = _T_85294[10:0]; // @[Modules.scala 53:83:@36788.4]
  assign buffer_9_661 = $signed(_T_85295); // @[Modules.scala 53:83:@36789.4]
  assign _T_85297 = $signed(buffer_3_540) + $signed(buffer_9_541); // @[Modules.scala 53:83:@36791.4]
  assign _T_85298 = _T_85297[10:0]; // @[Modules.scala 53:83:@36792.4]
  assign buffer_9_662 = $signed(_T_85298); // @[Modules.scala 53:83:@36793.4]
  assign _T_85300 = $signed(buffer_9_542) + $signed(buffer_0_543); // @[Modules.scala 53:83:@36795.4]
  assign _T_85301 = _T_85300[10:0]; // @[Modules.scala 53:83:@36796.4]
  assign buffer_9_663 = $signed(_T_85301); // @[Modules.scala 53:83:@36797.4]
  assign _T_85303 = $signed(buffer_9_544) + $signed(buffer_3_545); // @[Modules.scala 53:83:@36799.4]
  assign _T_85304 = _T_85303[10:0]; // @[Modules.scala 53:83:@36800.4]
  assign buffer_9_664 = $signed(_T_85304); // @[Modules.scala 53:83:@36801.4]
  assign _T_85309 = $signed(buffer_9_548) + $signed(buffer_5_549); // @[Modules.scala 53:83:@36807.4]
  assign _T_85310 = _T_85309[10:0]; // @[Modules.scala 53:83:@36808.4]
  assign buffer_9_666 = $signed(_T_85310); // @[Modules.scala 53:83:@36809.4]
  assign _T_85312 = $signed(buffer_9_550) + $signed(buffer_9_551); // @[Modules.scala 53:83:@36811.4]
  assign _T_85313 = _T_85312[10:0]; // @[Modules.scala 53:83:@36812.4]
  assign buffer_9_667 = $signed(_T_85313); // @[Modules.scala 53:83:@36813.4]
  assign _T_85315 = $signed(buffer_9_552) + $signed(buffer_1_553); // @[Modules.scala 53:83:@36815.4]
  assign _T_85316 = _T_85315[10:0]; // @[Modules.scala 53:83:@36816.4]
  assign buffer_9_668 = $signed(_T_85316); // @[Modules.scala 53:83:@36817.4]
  assign _T_85318 = $signed(buffer_1_554) + $signed(buffer_9_555); // @[Modules.scala 53:83:@36819.4]
  assign _T_85319 = _T_85318[10:0]; // @[Modules.scala 53:83:@36820.4]
  assign buffer_9_669 = $signed(_T_85319); // @[Modules.scala 53:83:@36821.4]
  assign _T_85324 = $signed(buffer_9_558) + $signed(buffer_8_559); // @[Modules.scala 53:83:@36827.4]
  assign _T_85325 = _T_85324[10:0]; // @[Modules.scala 53:83:@36828.4]
  assign buffer_9_671 = $signed(_T_85325); // @[Modules.scala 53:83:@36829.4]
  assign _T_85327 = $signed(buffer_5_560) + $signed(buffer_0_561); // @[Modules.scala 53:83:@36831.4]
  assign _T_85328 = _T_85327[10:0]; // @[Modules.scala 53:83:@36832.4]
  assign buffer_9_672 = $signed(_T_85328); // @[Modules.scala 53:83:@36833.4]
  assign _T_85333 = $signed(buffer_4_564) + $signed(buffer_9_565); // @[Modules.scala 53:83:@36839.4]
  assign _T_85334 = _T_85333[10:0]; // @[Modules.scala 53:83:@36840.4]
  assign buffer_9_674 = $signed(_T_85334); // @[Modules.scala 53:83:@36841.4]
  assign _T_85336 = $signed(buffer_9_566) + $signed(buffer_9_567); // @[Modules.scala 53:83:@36843.4]
  assign _T_85337 = _T_85336[10:0]; // @[Modules.scala 53:83:@36844.4]
  assign buffer_9_675 = $signed(_T_85337); // @[Modules.scala 53:83:@36845.4]
  assign _T_85339 = $signed(buffer_2_568) + $signed(buffer_9_569); // @[Modules.scala 53:83:@36847.4]
  assign _T_85340 = _T_85339[10:0]; // @[Modules.scala 53:83:@36848.4]
  assign buffer_9_676 = $signed(_T_85340); // @[Modules.scala 53:83:@36849.4]
  assign _T_85342 = $signed(buffer_9_570) + $signed(buffer_9_571); // @[Modules.scala 53:83:@36851.4]
  assign _T_85343 = _T_85342[10:0]; // @[Modules.scala 53:83:@36852.4]
  assign buffer_9_677 = $signed(_T_85343); // @[Modules.scala 53:83:@36853.4]
  assign _T_85345 = $signed(buffer_3_572) + $signed(buffer_9_573); // @[Modules.scala 53:83:@36855.4]
  assign _T_85346 = _T_85345[10:0]; // @[Modules.scala 53:83:@36856.4]
  assign buffer_9_678 = $signed(_T_85346); // @[Modules.scala 53:83:@36857.4]
  assign _T_85348 = $signed(buffer_9_574) + $signed(buffer_1_575); // @[Modules.scala 53:83:@36859.4]
  assign _T_85349 = _T_85348[10:0]; // @[Modules.scala 53:83:@36860.4]
  assign buffer_9_679 = $signed(_T_85349); // @[Modules.scala 53:83:@36861.4]
  assign _T_85354 = $signed(buffer_9_578) + $signed(buffer_9_579); // @[Modules.scala 53:83:@36867.4]
  assign _T_85355 = _T_85354[10:0]; // @[Modules.scala 53:83:@36868.4]
  assign buffer_9_681 = $signed(_T_85355); // @[Modules.scala 53:83:@36869.4]
  assign _T_85357 = $signed(buffer_9_580) + $signed(buffer_9_581); // @[Modules.scala 53:83:@36871.4]
  assign _T_85358 = _T_85357[10:0]; // @[Modules.scala 53:83:@36872.4]
  assign buffer_9_682 = $signed(_T_85358); // @[Modules.scala 53:83:@36873.4]
  assign _T_85360 = $signed(buffer_9_582) + $signed(buffer_9_583); // @[Modules.scala 53:83:@36875.4]
  assign _T_85361 = _T_85360[10:0]; // @[Modules.scala 53:83:@36876.4]
  assign buffer_9_683 = $signed(_T_85361); // @[Modules.scala 53:83:@36877.4]
  assign _T_85363 = $signed(buffer_3_584) + $signed(buffer_9_585); // @[Modules.scala 53:83:@36879.4]
  assign _T_85364 = _T_85363[10:0]; // @[Modules.scala 53:83:@36880.4]
  assign buffer_9_684 = $signed(_T_85364); // @[Modules.scala 53:83:@36881.4]
  assign _T_85369 = $signed(buffer_9_588) + $signed(buffer_9_589); // @[Modules.scala 56:109:@36887.4]
  assign _T_85370 = _T_85369[10:0]; // @[Modules.scala 56:109:@36888.4]
  assign buffer_9_686 = $signed(_T_85370); // @[Modules.scala 56:109:@36889.4]
  assign _T_85372 = $signed(buffer_9_590) + $signed(buffer_9_591); // @[Modules.scala 56:109:@36891.4]
  assign _T_85373 = _T_85372[10:0]; // @[Modules.scala 56:109:@36892.4]
  assign buffer_9_687 = $signed(_T_85373); // @[Modules.scala 56:109:@36893.4]
  assign _T_85375 = $signed(buffer_2_592) + $signed(buffer_9_593); // @[Modules.scala 56:109:@36895.4]
  assign _T_85376 = _T_85375[10:0]; // @[Modules.scala 56:109:@36896.4]
  assign buffer_9_688 = $signed(_T_85376); // @[Modules.scala 56:109:@36897.4]
  assign _T_85378 = $signed(buffer_9_594) + $signed(buffer_9_595); // @[Modules.scala 56:109:@36899.4]
  assign _T_85379 = _T_85378[10:0]; // @[Modules.scala 56:109:@36900.4]
  assign buffer_9_689 = $signed(_T_85379); // @[Modules.scala 56:109:@36901.4]
  assign _T_85384 = $signed(buffer_9_598) + $signed(buffer_1_599); // @[Modules.scala 56:109:@36907.4]
  assign _T_85385 = _T_85384[10:0]; // @[Modules.scala 56:109:@36908.4]
  assign buffer_9_691 = $signed(_T_85385); // @[Modules.scala 56:109:@36909.4]
  assign _T_85390 = $signed(buffer_9_602) + $signed(buffer_3_603); // @[Modules.scala 56:109:@36915.4]
  assign _T_85391 = _T_85390[10:0]; // @[Modules.scala 56:109:@36916.4]
  assign buffer_9_693 = $signed(_T_85391); // @[Modules.scala 56:109:@36917.4]
  assign _T_85393 = $signed(buffer_9_604) + $signed(buffer_9_605); // @[Modules.scala 56:109:@36919.4]
  assign _T_85394 = _T_85393[10:0]; // @[Modules.scala 56:109:@36920.4]
  assign buffer_9_694 = $signed(_T_85394); // @[Modules.scala 56:109:@36921.4]
  assign _T_85396 = $signed(buffer_9_606) + $signed(buffer_9_607); // @[Modules.scala 56:109:@36923.4]
  assign _T_85397 = _T_85396[10:0]; // @[Modules.scala 56:109:@36924.4]
  assign buffer_9_695 = $signed(_T_85397); // @[Modules.scala 56:109:@36925.4]
  assign _T_85399 = $signed(buffer_9_608) + $signed(buffer_9_609); // @[Modules.scala 56:109:@36927.4]
  assign _T_85400 = _T_85399[10:0]; // @[Modules.scala 56:109:@36928.4]
  assign buffer_9_696 = $signed(_T_85400); // @[Modules.scala 56:109:@36929.4]
  assign _T_85402 = $signed(buffer_9_610) + $signed(buffer_9_611); // @[Modules.scala 56:109:@36931.4]
  assign _T_85403 = _T_85402[10:0]; // @[Modules.scala 56:109:@36932.4]
  assign buffer_9_697 = $signed(_T_85403); // @[Modules.scala 56:109:@36933.4]
  assign _T_85405 = $signed(buffer_9_612) + $signed(buffer_9_613); // @[Modules.scala 56:109:@36935.4]
  assign _T_85406 = _T_85405[10:0]; // @[Modules.scala 56:109:@36936.4]
  assign buffer_9_698 = $signed(_T_85406); // @[Modules.scala 56:109:@36937.4]
  assign _T_85408 = $signed(buffer_9_614) + $signed(buffer_9_615); // @[Modules.scala 56:109:@36939.4]
  assign _T_85409 = _T_85408[10:0]; // @[Modules.scala 56:109:@36940.4]
  assign buffer_9_699 = $signed(_T_85409); // @[Modules.scala 56:109:@36941.4]
  assign _T_85411 = $signed(buffer_9_616) + $signed(buffer_9_617); // @[Modules.scala 56:109:@36943.4]
  assign _T_85412 = _T_85411[10:0]; // @[Modules.scala 56:109:@36944.4]
  assign buffer_9_700 = $signed(_T_85412); // @[Modules.scala 56:109:@36945.4]
  assign _T_85414 = $signed(buffer_9_618) + $signed(buffer_5_619); // @[Modules.scala 56:109:@36947.4]
  assign _T_85415 = _T_85414[10:0]; // @[Modules.scala 56:109:@36948.4]
  assign buffer_9_701 = $signed(_T_85415); // @[Modules.scala 56:109:@36949.4]
  assign _T_85417 = $signed(buffer_9_620) + $signed(buffer_9_621); // @[Modules.scala 56:109:@36951.4]
  assign _T_85418 = _T_85417[10:0]; // @[Modules.scala 56:109:@36952.4]
  assign buffer_9_702 = $signed(_T_85418); // @[Modules.scala 56:109:@36953.4]
  assign _T_85420 = $signed(buffer_9_622) + $signed(buffer_9_623); // @[Modules.scala 56:109:@36955.4]
  assign _T_85421 = _T_85420[10:0]; // @[Modules.scala 56:109:@36956.4]
  assign buffer_9_703 = $signed(_T_85421); // @[Modules.scala 56:109:@36957.4]
  assign _T_85423 = $signed(buffer_5_624) + $signed(buffer_9_625); // @[Modules.scala 56:109:@36959.4]
  assign _T_85424 = _T_85423[10:0]; // @[Modules.scala 56:109:@36960.4]
  assign buffer_9_704 = $signed(_T_85424); // @[Modules.scala 56:109:@36961.4]
  assign _T_85426 = $signed(buffer_9_626) + $signed(buffer_9_627); // @[Modules.scala 56:109:@36963.4]
  assign _T_85427 = _T_85426[10:0]; // @[Modules.scala 56:109:@36964.4]
  assign buffer_9_705 = $signed(_T_85427); // @[Modules.scala 56:109:@36965.4]
  assign _T_85429 = $signed(buffer_9_628) + $signed(buffer_9_629); // @[Modules.scala 56:109:@36967.4]
  assign _T_85430 = _T_85429[10:0]; // @[Modules.scala 56:109:@36968.4]
  assign buffer_9_706 = $signed(_T_85430); // @[Modules.scala 56:109:@36969.4]
  assign _T_85432 = $signed(buffer_8_630) + $signed(buffer_9_631); // @[Modules.scala 56:109:@36971.4]
  assign _T_85433 = _T_85432[10:0]; // @[Modules.scala 56:109:@36972.4]
  assign buffer_9_707 = $signed(_T_85433); // @[Modules.scala 56:109:@36973.4]
  assign _T_85435 = $signed(buffer_9_632) + $signed(buffer_4_633); // @[Modules.scala 56:109:@36975.4]
  assign _T_85436 = _T_85435[10:0]; // @[Modules.scala 56:109:@36976.4]
  assign buffer_9_708 = $signed(_T_85436); // @[Modules.scala 56:109:@36977.4]
  assign _T_85438 = $signed(buffer_9_634) + $signed(buffer_9_635); // @[Modules.scala 56:109:@36979.4]
  assign _T_85439 = _T_85438[10:0]; // @[Modules.scala 56:109:@36980.4]
  assign buffer_9_709 = $signed(_T_85439); // @[Modules.scala 56:109:@36981.4]
  assign _T_85441 = $signed(buffer_9_636) + $signed(buffer_9_637); // @[Modules.scala 56:109:@36983.4]
  assign _T_85442 = _T_85441[10:0]; // @[Modules.scala 56:109:@36984.4]
  assign buffer_9_710 = $signed(_T_85442); // @[Modules.scala 56:109:@36985.4]
  assign _T_85444 = $signed(buffer_9_638) + $signed(buffer_5_639); // @[Modules.scala 56:109:@36987.4]
  assign _T_85445 = _T_85444[10:0]; // @[Modules.scala 56:109:@36988.4]
  assign buffer_9_711 = $signed(_T_85445); // @[Modules.scala 56:109:@36989.4]
  assign _T_85447 = $signed(buffer_9_640) + $signed(buffer_9_641); // @[Modules.scala 56:109:@36991.4]
  assign _T_85448 = _T_85447[10:0]; // @[Modules.scala 56:109:@36992.4]
  assign buffer_9_712 = $signed(_T_85448); // @[Modules.scala 56:109:@36993.4]
  assign _T_85450 = $signed(buffer_2_642) + $signed(buffer_3_643); // @[Modules.scala 56:109:@36995.4]
  assign _T_85451 = _T_85450[10:0]; // @[Modules.scala 56:109:@36996.4]
  assign buffer_9_713 = $signed(_T_85451); // @[Modules.scala 56:109:@36997.4]
  assign _T_85453 = $signed(buffer_9_644) + $signed(buffer_9_645); // @[Modules.scala 56:109:@36999.4]
  assign _T_85454 = _T_85453[10:0]; // @[Modules.scala 56:109:@37000.4]
  assign buffer_9_714 = $signed(_T_85454); // @[Modules.scala 56:109:@37001.4]
  assign _T_85456 = $signed(buffer_9_646) + $signed(buffer_4_647); // @[Modules.scala 56:109:@37003.4]
  assign _T_85457 = _T_85456[10:0]; // @[Modules.scala 56:109:@37004.4]
  assign buffer_9_715 = $signed(_T_85457); // @[Modules.scala 56:109:@37005.4]
  assign _T_85459 = $signed(buffer_9_648) + $signed(buffer_9_649); // @[Modules.scala 56:109:@37007.4]
  assign _T_85460 = _T_85459[10:0]; // @[Modules.scala 56:109:@37008.4]
  assign buffer_9_716 = $signed(_T_85460); // @[Modules.scala 56:109:@37009.4]
  assign _T_85462 = $signed(buffer_3_650) + $signed(buffer_9_651); // @[Modules.scala 56:109:@37011.4]
  assign _T_85463 = _T_85462[10:0]; // @[Modules.scala 56:109:@37012.4]
  assign buffer_9_717 = $signed(_T_85463); // @[Modules.scala 56:109:@37013.4]
  assign _T_85465 = $signed(buffer_7_652) + $signed(buffer_3_653); // @[Modules.scala 56:109:@37015.4]
  assign _T_85466 = _T_85465[10:0]; // @[Modules.scala 56:109:@37016.4]
  assign buffer_9_718 = $signed(_T_85466); // @[Modules.scala 56:109:@37017.4]
  assign _T_85468 = $signed(buffer_8_654) + $signed(buffer_9_655); // @[Modules.scala 56:109:@37019.4]
  assign _T_85469 = _T_85468[10:0]; // @[Modules.scala 56:109:@37020.4]
  assign buffer_9_719 = $signed(_T_85469); // @[Modules.scala 56:109:@37021.4]
  assign _T_85471 = $signed(buffer_1_656) + $signed(buffer_3_657); // @[Modules.scala 56:109:@37023.4]
  assign _T_85472 = _T_85471[10:0]; // @[Modules.scala 56:109:@37024.4]
  assign buffer_9_720 = $signed(_T_85472); // @[Modules.scala 56:109:@37025.4]
  assign _T_85474 = $signed(buffer_9_658) + $signed(buffer_9_659); // @[Modules.scala 56:109:@37027.4]
  assign _T_85475 = _T_85474[10:0]; // @[Modules.scala 56:109:@37028.4]
  assign buffer_9_721 = $signed(_T_85475); // @[Modules.scala 56:109:@37029.4]
  assign _T_85477 = $signed(buffer_7_660) + $signed(buffer_9_661); // @[Modules.scala 56:109:@37031.4]
  assign _T_85478 = _T_85477[10:0]; // @[Modules.scala 56:109:@37032.4]
  assign buffer_9_722 = $signed(_T_85478); // @[Modules.scala 56:109:@37033.4]
  assign _T_85480 = $signed(buffer_9_662) + $signed(buffer_9_663); // @[Modules.scala 56:109:@37035.4]
  assign _T_85481 = _T_85480[10:0]; // @[Modules.scala 56:109:@37036.4]
  assign buffer_9_723 = $signed(_T_85481); // @[Modules.scala 56:109:@37037.4]
  assign _T_85483 = $signed(buffer_9_664) + $signed(buffer_4_665); // @[Modules.scala 56:109:@37039.4]
  assign _T_85484 = _T_85483[10:0]; // @[Modules.scala 56:109:@37040.4]
  assign buffer_9_724 = $signed(_T_85484); // @[Modules.scala 56:109:@37041.4]
  assign _T_85486 = $signed(buffer_9_666) + $signed(buffer_9_667); // @[Modules.scala 56:109:@37043.4]
  assign _T_85487 = _T_85486[10:0]; // @[Modules.scala 56:109:@37044.4]
  assign buffer_9_725 = $signed(_T_85487); // @[Modules.scala 56:109:@37045.4]
  assign _T_85489 = $signed(buffer_9_668) + $signed(buffer_9_669); // @[Modules.scala 56:109:@37047.4]
  assign _T_85490 = _T_85489[10:0]; // @[Modules.scala 56:109:@37048.4]
  assign buffer_9_726 = $signed(_T_85490); // @[Modules.scala 56:109:@37049.4]
  assign _T_85492 = $signed(buffer_4_670) + $signed(buffer_9_671); // @[Modules.scala 56:109:@37051.4]
  assign _T_85493 = _T_85492[10:0]; // @[Modules.scala 56:109:@37052.4]
  assign buffer_9_727 = $signed(_T_85493); // @[Modules.scala 56:109:@37053.4]
  assign _T_85495 = $signed(buffer_9_672) + $signed(buffer_4_673); // @[Modules.scala 56:109:@37055.4]
  assign _T_85496 = _T_85495[10:0]; // @[Modules.scala 56:109:@37056.4]
  assign buffer_9_728 = $signed(_T_85496); // @[Modules.scala 56:109:@37057.4]
  assign _T_85498 = $signed(buffer_9_674) + $signed(buffer_9_675); // @[Modules.scala 56:109:@37059.4]
  assign _T_85499 = _T_85498[10:0]; // @[Modules.scala 56:109:@37060.4]
  assign buffer_9_729 = $signed(_T_85499); // @[Modules.scala 56:109:@37061.4]
  assign _T_85501 = $signed(buffer_9_676) + $signed(buffer_9_677); // @[Modules.scala 56:109:@37063.4]
  assign _T_85502 = _T_85501[10:0]; // @[Modules.scala 56:109:@37064.4]
  assign buffer_9_730 = $signed(_T_85502); // @[Modules.scala 56:109:@37065.4]
  assign _T_85504 = $signed(buffer_9_678) + $signed(buffer_9_679); // @[Modules.scala 56:109:@37067.4]
  assign _T_85505 = _T_85504[10:0]; // @[Modules.scala 56:109:@37068.4]
  assign buffer_9_731 = $signed(_T_85505); // @[Modules.scala 56:109:@37069.4]
  assign _T_85507 = $signed(buffer_1_680) + $signed(buffer_9_681); // @[Modules.scala 56:109:@37071.4]
  assign _T_85508 = _T_85507[10:0]; // @[Modules.scala 56:109:@37072.4]
  assign buffer_9_732 = $signed(_T_85508); // @[Modules.scala 56:109:@37073.4]
  assign _T_85510 = $signed(buffer_9_682) + $signed(buffer_9_683); // @[Modules.scala 56:109:@37075.4]
  assign _T_85511 = _T_85510[10:0]; // @[Modules.scala 56:109:@37076.4]
  assign buffer_9_733 = $signed(_T_85511); // @[Modules.scala 56:109:@37077.4]
  assign _T_85513 = $signed(buffer_9_684) + $signed(buffer_5_685); // @[Modules.scala 56:109:@37079.4]
  assign _T_85514 = _T_85513[10:0]; // @[Modules.scala 56:109:@37080.4]
  assign buffer_9_734 = $signed(_T_85514); // @[Modules.scala 56:109:@37081.4]
  assign _T_85516 = $signed(buffer_9_686) + $signed(buffer_9_687); // @[Modules.scala 63:156:@37084.4]
  assign _T_85517 = _T_85516[10:0]; // @[Modules.scala 63:156:@37085.4]
  assign buffer_9_736 = $signed(_T_85517); // @[Modules.scala 63:156:@37086.4]
  assign _T_85519 = $signed(buffer_9_736) + $signed(buffer_9_688); // @[Modules.scala 63:156:@37088.4]
  assign _T_85520 = _T_85519[10:0]; // @[Modules.scala 63:156:@37089.4]
  assign buffer_9_737 = $signed(_T_85520); // @[Modules.scala 63:156:@37090.4]
  assign _T_85522 = $signed(buffer_9_737) + $signed(buffer_9_689); // @[Modules.scala 63:156:@37092.4]
  assign _T_85523 = _T_85522[10:0]; // @[Modules.scala 63:156:@37093.4]
  assign buffer_9_738 = $signed(_T_85523); // @[Modules.scala 63:156:@37094.4]
  assign _T_85525 = $signed(buffer_9_738) + $signed(buffer_1_690); // @[Modules.scala 63:156:@37096.4]
  assign _T_85526 = _T_85525[10:0]; // @[Modules.scala 63:156:@37097.4]
  assign buffer_9_739 = $signed(_T_85526); // @[Modules.scala 63:156:@37098.4]
  assign _T_85528 = $signed(buffer_9_739) + $signed(buffer_9_691); // @[Modules.scala 63:156:@37100.4]
  assign _T_85529 = _T_85528[10:0]; // @[Modules.scala 63:156:@37101.4]
  assign buffer_9_740 = $signed(_T_85529); // @[Modules.scala 63:156:@37102.4]
  assign _T_85531 = $signed(buffer_9_740) + $signed(buffer_1_692); // @[Modules.scala 63:156:@37104.4]
  assign _T_85532 = _T_85531[10:0]; // @[Modules.scala 63:156:@37105.4]
  assign buffer_9_741 = $signed(_T_85532); // @[Modules.scala 63:156:@37106.4]
  assign _T_85534 = $signed(buffer_9_741) + $signed(buffer_9_693); // @[Modules.scala 63:156:@37108.4]
  assign _T_85535 = _T_85534[10:0]; // @[Modules.scala 63:156:@37109.4]
  assign buffer_9_742 = $signed(_T_85535); // @[Modules.scala 63:156:@37110.4]
  assign _T_85537 = $signed(buffer_9_742) + $signed(buffer_9_694); // @[Modules.scala 63:156:@37112.4]
  assign _T_85538 = _T_85537[10:0]; // @[Modules.scala 63:156:@37113.4]
  assign buffer_9_743 = $signed(_T_85538); // @[Modules.scala 63:156:@37114.4]
  assign _T_85540 = $signed(buffer_9_743) + $signed(buffer_9_695); // @[Modules.scala 63:156:@37116.4]
  assign _T_85541 = _T_85540[10:0]; // @[Modules.scala 63:156:@37117.4]
  assign buffer_9_744 = $signed(_T_85541); // @[Modules.scala 63:156:@37118.4]
  assign _T_85543 = $signed(buffer_9_744) + $signed(buffer_9_696); // @[Modules.scala 63:156:@37120.4]
  assign _T_85544 = _T_85543[10:0]; // @[Modules.scala 63:156:@37121.4]
  assign buffer_9_745 = $signed(_T_85544); // @[Modules.scala 63:156:@37122.4]
  assign _T_85546 = $signed(buffer_9_745) + $signed(buffer_9_697); // @[Modules.scala 63:156:@37124.4]
  assign _T_85547 = _T_85546[10:0]; // @[Modules.scala 63:156:@37125.4]
  assign buffer_9_746 = $signed(_T_85547); // @[Modules.scala 63:156:@37126.4]
  assign _T_85549 = $signed(buffer_9_746) + $signed(buffer_9_698); // @[Modules.scala 63:156:@37128.4]
  assign _T_85550 = _T_85549[10:0]; // @[Modules.scala 63:156:@37129.4]
  assign buffer_9_747 = $signed(_T_85550); // @[Modules.scala 63:156:@37130.4]
  assign _T_85552 = $signed(buffer_9_747) + $signed(buffer_9_699); // @[Modules.scala 63:156:@37132.4]
  assign _T_85553 = _T_85552[10:0]; // @[Modules.scala 63:156:@37133.4]
  assign buffer_9_748 = $signed(_T_85553); // @[Modules.scala 63:156:@37134.4]
  assign _T_85555 = $signed(buffer_9_748) + $signed(buffer_9_700); // @[Modules.scala 63:156:@37136.4]
  assign _T_85556 = _T_85555[10:0]; // @[Modules.scala 63:156:@37137.4]
  assign buffer_9_749 = $signed(_T_85556); // @[Modules.scala 63:156:@37138.4]
  assign _T_85558 = $signed(buffer_9_749) + $signed(buffer_9_701); // @[Modules.scala 63:156:@37140.4]
  assign _T_85559 = _T_85558[10:0]; // @[Modules.scala 63:156:@37141.4]
  assign buffer_9_750 = $signed(_T_85559); // @[Modules.scala 63:156:@37142.4]
  assign _T_85561 = $signed(buffer_9_750) + $signed(buffer_9_702); // @[Modules.scala 63:156:@37144.4]
  assign _T_85562 = _T_85561[10:0]; // @[Modules.scala 63:156:@37145.4]
  assign buffer_9_751 = $signed(_T_85562); // @[Modules.scala 63:156:@37146.4]
  assign _T_85564 = $signed(buffer_9_751) + $signed(buffer_9_703); // @[Modules.scala 63:156:@37148.4]
  assign _T_85565 = _T_85564[10:0]; // @[Modules.scala 63:156:@37149.4]
  assign buffer_9_752 = $signed(_T_85565); // @[Modules.scala 63:156:@37150.4]
  assign _T_85567 = $signed(buffer_9_752) + $signed(buffer_9_704); // @[Modules.scala 63:156:@37152.4]
  assign _T_85568 = _T_85567[10:0]; // @[Modules.scala 63:156:@37153.4]
  assign buffer_9_753 = $signed(_T_85568); // @[Modules.scala 63:156:@37154.4]
  assign _T_85570 = $signed(buffer_9_753) + $signed(buffer_9_705); // @[Modules.scala 63:156:@37156.4]
  assign _T_85571 = _T_85570[10:0]; // @[Modules.scala 63:156:@37157.4]
  assign buffer_9_754 = $signed(_T_85571); // @[Modules.scala 63:156:@37158.4]
  assign _T_85573 = $signed(buffer_9_754) + $signed(buffer_9_706); // @[Modules.scala 63:156:@37160.4]
  assign _T_85574 = _T_85573[10:0]; // @[Modules.scala 63:156:@37161.4]
  assign buffer_9_755 = $signed(_T_85574); // @[Modules.scala 63:156:@37162.4]
  assign _T_85576 = $signed(buffer_9_755) + $signed(buffer_9_707); // @[Modules.scala 63:156:@37164.4]
  assign _T_85577 = _T_85576[10:0]; // @[Modules.scala 63:156:@37165.4]
  assign buffer_9_756 = $signed(_T_85577); // @[Modules.scala 63:156:@37166.4]
  assign _T_85579 = $signed(buffer_9_756) + $signed(buffer_9_708); // @[Modules.scala 63:156:@37168.4]
  assign _T_85580 = _T_85579[10:0]; // @[Modules.scala 63:156:@37169.4]
  assign buffer_9_757 = $signed(_T_85580); // @[Modules.scala 63:156:@37170.4]
  assign _T_85582 = $signed(buffer_9_757) + $signed(buffer_9_709); // @[Modules.scala 63:156:@37172.4]
  assign _T_85583 = _T_85582[10:0]; // @[Modules.scala 63:156:@37173.4]
  assign buffer_9_758 = $signed(_T_85583); // @[Modules.scala 63:156:@37174.4]
  assign _T_85585 = $signed(buffer_9_758) + $signed(buffer_9_710); // @[Modules.scala 63:156:@37176.4]
  assign _T_85586 = _T_85585[10:0]; // @[Modules.scala 63:156:@37177.4]
  assign buffer_9_759 = $signed(_T_85586); // @[Modules.scala 63:156:@37178.4]
  assign _T_85588 = $signed(buffer_9_759) + $signed(buffer_9_711); // @[Modules.scala 63:156:@37180.4]
  assign _T_85589 = _T_85588[10:0]; // @[Modules.scala 63:156:@37181.4]
  assign buffer_9_760 = $signed(_T_85589); // @[Modules.scala 63:156:@37182.4]
  assign _T_85591 = $signed(buffer_9_760) + $signed(buffer_9_712); // @[Modules.scala 63:156:@37184.4]
  assign _T_85592 = _T_85591[10:0]; // @[Modules.scala 63:156:@37185.4]
  assign buffer_9_761 = $signed(_T_85592); // @[Modules.scala 63:156:@37186.4]
  assign _T_85594 = $signed(buffer_9_761) + $signed(buffer_9_713); // @[Modules.scala 63:156:@37188.4]
  assign _T_85595 = _T_85594[10:0]; // @[Modules.scala 63:156:@37189.4]
  assign buffer_9_762 = $signed(_T_85595); // @[Modules.scala 63:156:@37190.4]
  assign _T_85597 = $signed(buffer_9_762) + $signed(buffer_9_714); // @[Modules.scala 63:156:@37192.4]
  assign _T_85598 = _T_85597[10:0]; // @[Modules.scala 63:156:@37193.4]
  assign buffer_9_763 = $signed(_T_85598); // @[Modules.scala 63:156:@37194.4]
  assign _T_85600 = $signed(buffer_9_763) + $signed(buffer_9_715); // @[Modules.scala 63:156:@37196.4]
  assign _T_85601 = _T_85600[10:0]; // @[Modules.scala 63:156:@37197.4]
  assign buffer_9_764 = $signed(_T_85601); // @[Modules.scala 63:156:@37198.4]
  assign _T_85603 = $signed(buffer_9_764) + $signed(buffer_9_716); // @[Modules.scala 63:156:@37200.4]
  assign _T_85604 = _T_85603[10:0]; // @[Modules.scala 63:156:@37201.4]
  assign buffer_9_765 = $signed(_T_85604); // @[Modules.scala 63:156:@37202.4]
  assign _T_85606 = $signed(buffer_9_765) + $signed(buffer_9_717); // @[Modules.scala 63:156:@37204.4]
  assign _T_85607 = _T_85606[10:0]; // @[Modules.scala 63:156:@37205.4]
  assign buffer_9_766 = $signed(_T_85607); // @[Modules.scala 63:156:@37206.4]
  assign _T_85609 = $signed(buffer_9_766) + $signed(buffer_9_718); // @[Modules.scala 63:156:@37208.4]
  assign _T_85610 = _T_85609[10:0]; // @[Modules.scala 63:156:@37209.4]
  assign buffer_9_767 = $signed(_T_85610); // @[Modules.scala 63:156:@37210.4]
  assign _T_85612 = $signed(buffer_9_767) + $signed(buffer_9_719); // @[Modules.scala 63:156:@37212.4]
  assign _T_85613 = _T_85612[10:0]; // @[Modules.scala 63:156:@37213.4]
  assign buffer_9_768 = $signed(_T_85613); // @[Modules.scala 63:156:@37214.4]
  assign _T_85615 = $signed(buffer_9_768) + $signed(buffer_9_720); // @[Modules.scala 63:156:@37216.4]
  assign _T_85616 = _T_85615[10:0]; // @[Modules.scala 63:156:@37217.4]
  assign buffer_9_769 = $signed(_T_85616); // @[Modules.scala 63:156:@37218.4]
  assign _T_85618 = $signed(buffer_9_769) + $signed(buffer_9_721); // @[Modules.scala 63:156:@37220.4]
  assign _T_85619 = _T_85618[10:0]; // @[Modules.scala 63:156:@37221.4]
  assign buffer_9_770 = $signed(_T_85619); // @[Modules.scala 63:156:@37222.4]
  assign _T_85621 = $signed(buffer_9_770) + $signed(buffer_9_722); // @[Modules.scala 63:156:@37224.4]
  assign _T_85622 = _T_85621[10:0]; // @[Modules.scala 63:156:@37225.4]
  assign buffer_9_771 = $signed(_T_85622); // @[Modules.scala 63:156:@37226.4]
  assign _T_85624 = $signed(buffer_9_771) + $signed(buffer_9_723); // @[Modules.scala 63:156:@37228.4]
  assign _T_85625 = _T_85624[10:0]; // @[Modules.scala 63:156:@37229.4]
  assign buffer_9_772 = $signed(_T_85625); // @[Modules.scala 63:156:@37230.4]
  assign _T_85627 = $signed(buffer_9_772) + $signed(buffer_9_724); // @[Modules.scala 63:156:@37232.4]
  assign _T_85628 = _T_85627[10:0]; // @[Modules.scala 63:156:@37233.4]
  assign buffer_9_773 = $signed(_T_85628); // @[Modules.scala 63:156:@37234.4]
  assign _T_85630 = $signed(buffer_9_773) + $signed(buffer_9_725); // @[Modules.scala 63:156:@37236.4]
  assign _T_85631 = _T_85630[10:0]; // @[Modules.scala 63:156:@37237.4]
  assign buffer_9_774 = $signed(_T_85631); // @[Modules.scala 63:156:@37238.4]
  assign _T_85633 = $signed(buffer_9_774) + $signed(buffer_9_726); // @[Modules.scala 63:156:@37240.4]
  assign _T_85634 = _T_85633[10:0]; // @[Modules.scala 63:156:@37241.4]
  assign buffer_9_775 = $signed(_T_85634); // @[Modules.scala 63:156:@37242.4]
  assign _T_85636 = $signed(buffer_9_775) + $signed(buffer_9_727); // @[Modules.scala 63:156:@37244.4]
  assign _T_85637 = _T_85636[10:0]; // @[Modules.scala 63:156:@37245.4]
  assign buffer_9_776 = $signed(_T_85637); // @[Modules.scala 63:156:@37246.4]
  assign _T_85639 = $signed(buffer_9_776) + $signed(buffer_9_728); // @[Modules.scala 63:156:@37248.4]
  assign _T_85640 = _T_85639[10:0]; // @[Modules.scala 63:156:@37249.4]
  assign buffer_9_777 = $signed(_T_85640); // @[Modules.scala 63:156:@37250.4]
  assign _T_85642 = $signed(buffer_9_777) + $signed(buffer_9_729); // @[Modules.scala 63:156:@37252.4]
  assign _T_85643 = _T_85642[10:0]; // @[Modules.scala 63:156:@37253.4]
  assign buffer_9_778 = $signed(_T_85643); // @[Modules.scala 63:156:@37254.4]
  assign _T_85645 = $signed(buffer_9_778) + $signed(buffer_9_730); // @[Modules.scala 63:156:@37256.4]
  assign _T_85646 = _T_85645[10:0]; // @[Modules.scala 63:156:@37257.4]
  assign buffer_9_779 = $signed(_T_85646); // @[Modules.scala 63:156:@37258.4]
  assign _T_85648 = $signed(buffer_9_779) + $signed(buffer_9_731); // @[Modules.scala 63:156:@37260.4]
  assign _T_85649 = _T_85648[10:0]; // @[Modules.scala 63:156:@37261.4]
  assign buffer_9_780 = $signed(_T_85649); // @[Modules.scala 63:156:@37262.4]
  assign _T_85651 = $signed(buffer_9_780) + $signed(buffer_9_732); // @[Modules.scala 63:156:@37264.4]
  assign _T_85652 = _T_85651[10:0]; // @[Modules.scala 63:156:@37265.4]
  assign buffer_9_781 = $signed(_T_85652); // @[Modules.scala 63:156:@37266.4]
  assign _T_85654 = $signed(buffer_9_781) + $signed(buffer_9_733); // @[Modules.scala 63:156:@37268.4]
  assign _T_85655 = _T_85654[10:0]; // @[Modules.scala 63:156:@37269.4]
  assign buffer_9_782 = $signed(_T_85655); // @[Modules.scala 63:156:@37270.4]
  assign _T_85657 = $signed(buffer_9_782) + $signed(buffer_9_734); // @[Modules.scala 63:156:@37272.4]
  assign _T_85658 = _T_85657[10:0]; // @[Modules.scala 63:156:@37273.4]
  assign buffer_9_783 = $signed(_T_85658); // @[Modules.scala 63:156:@37274.4]
  assign _T_85880 = $signed(io_in_112) + $signed(io_in_113); // @[Modules.scala 37:46:@37540.4]
  assign _T_85881 = _T_85880[4:0]; // @[Modules.scala 37:46:@37541.4]
  assign _T_85882 = $signed(_T_85881); // @[Modules.scala 37:46:@37542.4]
  assign _T_85959 = $signed(_T_54688) + $signed(io_in_155); // @[Modules.scala 43:47:@37636.4]
  assign _T_85960 = _T_85959[4:0]; // @[Modules.scala 43:47:@37637.4]
  assign _T_85961 = $signed(_T_85960); // @[Modules.scala 43:47:@37638.4]
  assign _T_86000 = $signed(io_in_176) - $signed(io_in_177); // @[Modules.scala 40:46:@37686.4]
  assign _T_86001 = _T_86000[4:0]; // @[Modules.scala 40:46:@37687.4]
  assign _T_86002 = $signed(_T_86001); // @[Modules.scala 40:46:@37688.4]
  assign _T_86068 = $signed(io_in_200) - $signed(io_in_201); // @[Modules.scala 40:46:@37758.4]
  assign _T_86069 = _T_86068[4:0]; // @[Modules.scala 40:46:@37759.4]
  assign _T_86070 = $signed(_T_86069); // @[Modules.scala 40:46:@37760.4]
  assign _T_86165 = $signed(io_in_238) - $signed(io_in_239); // @[Modules.scala 40:46:@37864.4]
  assign _T_86166 = _T_86165[4:0]; // @[Modules.scala 40:46:@37865.4]
  assign _T_86167 = $signed(_T_86166); // @[Modules.scala 40:46:@37866.4]
  assign _T_86386 = $signed(io_in_308) + $signed(io_in_309); // @[Modules.scala 37:46:@38091.4]
  assign _T_86387 = _T_86386[4:0]; // @[Modules.scala 37:46:@38092.4]
  assign _T_86388 = $signed(_T_86387); // @[Modules.scala 37:46:@38093.4]
  assign _T_86607 = $signed(_T_61662) + $signed(io_in_387); // @[Modules.scala 43:47:@38325.4]
  assign _T_86608 = _T_86607[4:0]; // @[Modules.scala 43:47:@38326.4]
  assign _T_86609 = $signed(_T_86608); // @[Modules.scala 43:47:@38327.4]
  assign _T_86657 = $signed(io_in_406) - $signed(io_in_407); // @[Modules.scala 40:46:@38380.4]
  assign _T_86658 = _T_86657[4:0]; // @[Modules.scala 40:46:@38381.4]
  assign _T_86659 = $signed(_T_86658); // @[Modules.scala 40:46:@38382.4]
  assign _T_86774 = $signed(_T_58692) + $signed(io_in_461); // @[Modules.scala 43:47:@38515.4]
  assign _T_86775 = _T_86774[4:0]; // @[Modules.scala 43:47:@38516.4]
  assign _T_86776 = $signed(_T_86775); // @[Modules.scala 43:47:@38517.4]
  assign _T_86873 = $signed(_T_55658) + $signed(io_in_511); // @[Modules.scala 43:47:@38633.4]
  assign _T_86874 = _T_86873[4:0]; // @[Modules.scala 43:47:@38634.4]
  assign _T_86875 = $signed(_T_86874); // @[Modules.scala 43:47:@38635.4]
  assign _T_87126 = $signed(io_in_636) - $signed(io_in_637); // @[Modules.scala 40:46:@38933.4]
  assign _T_87127 = _T_87126[4:0]; // @[Modules.scala 40:46:@38934.4]
  assign _T_87128 = $signed(_T_87127); // @[Modules.scala 40:46:@38935.4]
  assign _T_87146 = $signed(io_in_644) + $signed(io_in_645); // @[Modules.scala 37:46:@38955.4]
  assign _T_87147 = _T_87146[4:0]; // @[Modules.scala 37:46:@38956.4]
  assign _T_87148 = $signed(_T_87147); // @[Modules.scala 37:46:@38957.4]
  assign _T_87291 = $signed(io_in_706) - $signed(io_in_707); // @[Modules.scala 40:46:@39118.4]
  assign _T_87292 = _T_87291[4:0]; // @[Modules.scala 40:46:@39119.4]
  assign _T_87293 = $signed(_T_87292); // @[Modules.scala 40:46:@39120.4]
  assign _T_87380 = $signed(_T_56249) + $signed(io_in_737); // @[Modules.scala 43:47:@39211.4]
  assign _T_87381 = _T_87380[4:0]; // @[Modules.scala 43:47:@39212.4]
  assign _T_87382 = $signed(_T_87381); // @[Modules.scala 43:47:@39213.4]
  assign _T_87495 = $signed(buffer_9_2) + $signed(buffer_1_3); // @[Modules.scala 50:57:@39341.4]
  assign _T_87496 = _T_87495[10:0]; // @[Modules.scala 50:57:@39342.4]
  assign buffer_10_393 = $signed(_T_87496); // @[Modules.scala 50:57:@39343.4]
  assign _T_87498 = $signed(buffer_1_4) + $signed(buffer_3_5); // @[Modules.scala 50:57:@39345.4]
  assign _T_87499 = _T_87498[10:0]; // @[Modules.scala 50:57:@39346.4]
  assign buffer_10_394 = $signed(_T_87499); // @[Modules.scala 50:57:@39347.4]
  assign _T_87510 = $signed(buffer_0_12) + $signed(buffer_3_13); // @[Modules.scala 50:57:@39361.4]
  assign _T_87511 = _T_87510[10:0]; // @[Modules.scala 50:57:@39362.4]
  assign buffer_10_398 = $signed(_T_87511); // @[Modules.scala 50:57:@39363.4]
  assign _T_87531 = $signed(buffer_1_26) + $signed(buffer_0_27); // @[Modules.scala 50:57:@39389.4]
  assign _T_87532 = _T_87531[10:0]; // @[Modules.scala 50:57:@39390.4]
  assign buffer_10_405 = $signed(_T_87532); // @[Modules.scala 50:57:@39391.4]
  assign _T_87537 = $signed(buffer_0_30) + $signed(buffer_1_31); // @[Modules.scala 50:57:@39397.4]
  assign _T_87538 = _T_87537[10:0]; // @[Modules.scala 50:57:@39398.4]
  assign buffer_10_407 = $signed(_T_87538); // @[Modules.scala 50:57:@39399.4]
  assign _T_87555 = $signed(buffer_0_42) + $signed(buffer_1_43); // @[Modules.scala 50:57:@39421.4]
  assign _T_87556 = _T_87555[10:0]; // @[Modules.scala 50:57:@39422.4]
  assign buffer_10_413 = $signed(_T_87556); // @[Modules.scala 50:57:@39423.4]
  assign _T_87573 = $signed(buffer_0_54) + $signed(buffer_3_55); // @[Modules.scala 50:57:@39445.4]
  assign _T_87574 = _T_87573[10:0]; // @[Modules.scala 50:57:@39446.4]
  assign buffer_10_419 = $signed(_T_87574); // @[Modules.scala 50:57:@39447.4]
  assign buffer_10_56 = {{6{_T_85882[4]}},_T_85882}; // @[Modules.scala 32:22:@8.4]
  assign _T_87576 = $signed(buffer_10_56) + $signed(buffer_1_57); // @[Modules.scala 50:57:@39449.4]
  assign _T_87577 = _T_87576[10:0]; // @[Modules.scala 50:57:@39450.4]
  assign buffer_10_420 = $signed(_T_87577); // @[Modules.scala 50:57:@39451.4]
  assign _T_87588 = $signed(buffer_4_64) + $signed(buffer_1_65); // @[Modules.scala 50:57:@39465.4]
  assign _T_87589 = _T_87588[10:0]; // @[Modules.scala 50:57:@39466.4]
  assign buffer_10_424 = $signed(_T_87589); // @[Modules.scala 50:57:@39467.4]
  assign _T_87594 = $signed(buffer_5_68) + $signed(buffer_4_69); // @[Modules.scala 50:57:@39473.4]
  assign _T_87595 = _T_87594[10:0]; // @[Modules.scala 50:57:@39474.4]
  assign buffer_10_426 = $signed(_T_87595); // @[Modules.scala 50:57:@39475.4]
  assign _T_87597 = $signed(buffer_1_70) + $signed(buffer_5_71); // @[Modules.scala 50:57:@39477.4]
  assign _T_87598 = _T_87597[10:0]; // @[Modules.scala 50:57:@39478.4]
  assign buffer_10_427 = $signed(_T_87598); // @[Modules.scala 50:57:@39479.4]
  assign _T_87603 = $signed(buffer_1_74) + $signed(buffer_3_75); // @[Modules.scala 50:57:@39485.4]
  assign _T_87604 = _T_87603[10:0]; // @[Modules.scala 50:57:@39486.4]
  assign buffer_10_429 = $signed(_T_87604); // @[Modules.scala 50:57:@39487.4]
  assign buffer_10_77 = {{6{_T_85961[4]}},_T_85961}; // @[Modules.scala 32:22:@8.4]
  assign _T_87606 = $signed(buffer_4_76) + $signed(buffer_10_77); // @[Modules.scala 50:57:@39489.4]
  assign _T_87607 = _T_87606[10:0]; // @[Modules.scala 50:57:@39490.4]
  assign buffer_10_430 = $signed(_T_87607); // @[Modules.scala 50:57:@39491.4]
  assign _T_87609 = $signed(buffer_4_78) + $signed(buffer_0_79); // @[Modules.scala 50:57:@39493.4]
  assign _T_87610 = _T_87609[10:0]; // @[Modules.scala 50:57:@39494.4]
  assign buffer_10_431 = $signed(_T_87610); // @[Modules.scala 50:57:@39495.4]
  assign _T_87612 = $signed(buffer_4_80) + $signed(buffer_0_81); // @[Modules.scala 50:57:@39497.4]
  assign _T_87613 = _T_87612[10:0]; // @[Modules.scala 50:57:@39498.4]
  assign buffer_10_432 = $signed(_T_87613); // @[Modules.scala 50:57:@39499.4]
  assign _T_87615 = $signed(buffer_0_82) + $signed(buffer_1_83); // @[Modules.scala 50:57:@39501.4]
  assign _T_87616 = _T_87615[10:0]; // @[Modules.scala 50:57:@39502.4]
  assign buffer_10_433 = $signed(_T_87616); // @[Modules.scala 50:57:@39503.4]
  assign _T_87618 = $signed(buffer_4_84) + $signed(buffer_1_85); // @[Modules.scala 50:57:@39505.4]
  assign _T_87619 = _T_87618[10:0]; // @[Modules.scala 50:57:@39506.4]
  assign buffer_10_434 = $signed(_T_87619); // @[Modules.scala 50:57:@39507.4]
  assign _T_87621 = $signed(buffer_0_86) + $signed(buffer_7_87); // @[Modules.scala 50:57:@39509.4]
  assign _T_87622 = _T_87621[10:0]; // @[Modules.scala 50:57:@39510.4]
  assign buffer_10_435 = $signed(_T_87622); // @[Modules.scala 50:57:@39511.4]
  assign buffer_10_88 = {{6{_T_86002[4]}},_T_86002}; // @[Modules.scala 32:22:@8.4]
  assign _T_87624 = $signed(buffer_10_88) + $signed(buffer_7_89); // @[Modules.scala 50:57:@39513.4]
  assign _T_87625 = _T_87624[10:0]; // @[Modules.scala 50:57:@39514.4]
  assign buffer_10_436 = $signed(_T_87625); // @[Modules.scala 50:57:@39515.4]
  assign _T_87636 = $signed(buffer_0_96) + $signed(buffer_2_97); // @[Modules.scala 50:57:@39529.4]
  assign _T_87637 = _T_87636[10:0]; // @[Modules.scala 50:57:@39530.4]
  assign buffer_10_440 = $signed(_T_87637); // @[Modules.scala 50:57:@39531.4]
  assign buffer_10_100 = {{6{_T_86070[4]}},_T_86070}; // @[Modules.scala 32:22:@8.4]
  assign _T_87642 = $signed(buffer_10_100) + $signed(buffer_1_101); // @[Modules.scala 50:57:@39537.4]
  assign _T_87643 = _T_87642[10:0]; // @[Modules.scala 50:57:@39538.4]
  assign buffer_10_442 = $signed(_T_87643); // @[Modules.scala 50:57:@39539.4]
  assign _T_87645 = $signed(buffer_0_102) + $signed(buffer_1_103); // @[Modules.scala 50:57:@39541.4]
  assign _T_87646 = _T_87645[10:0]; // @[Modules.scala 50:57:@39542.4]
  assign buffer_10_443 = $signed(_T_87646); // @[Modules.scala 50:57:@39543.4]
  assign _T_87648 = $signed(buffer_2_104) + $signed(buffer_3_105); // @[Modules.scala 50:57:@39545.4]
  assign _T_87649 = _T_87648[10:0]; // @[Modules.scala 50:57:@39546.4]
  assign buffer_10_444 = $signed(_T_87649); // @[Modules.scala 50:57:@39547.4]
  assign _T_87663 = $signed(buffer_3_114) + $signed(buffer_0_115); // @[Modules.scala 50:57:@39565.4]
  assign _T_87664 = _T_87663[10:0]; // @[Modules.scala 50:57:@39566.4]
  assign buffer_10_449 = $signed(_T_87664); // @[Modules.scala 50:57:@39567.4]
  assign buffer_10_119 = {{6{_T_86167[4]}},_T_86167}; // @[Modules.scala 32:22:@8.4]
  assign _T_87669 = $signed(buffer_1_118) + $signed(buffer_10_119); // @[Modules.scala 50:57:@39573.4]
  assign _T_87670 = _T_87669[10:0]; // @[Modules.scala 50:57:@39574.4]
  assign buffer_10_451 = $signed(_T_87670); // @[Modules.scala 50:57:@39575.4]
  assign buffer_10_154 = {{6{_T_86388[4]}},_T_86388}; // @[Modules.scala 32:22:@8.4]
  assign _T_87723 = $signed(buffer_10_154) + $signed(buffer_3_155); // @[Modules.scala 50:57:@39645.4]
  assign _T_87724 = _T_87723[10:0]; // @[Modules.scala 50:57:@39646.4]
  assign buffer_10_469 = $signed(_T_87724); // @[Modules.scala 50:57:@39647.4]
  assign _T_87735 = $signed(buffer_5_162) + $signed(buffer_0_163); // @[Modules.scala 50:57:@39661.4]
  assign _T_87736 = _T_87735[10:0]; // @[Modules.scala 50:57:@39662.4]
  assign buffer_10_473 = $signed(_T_87736); // @[Modules.scala 50:57:@39663.4]
  assign _T_87741 = $signed(buffer_2_166) + $signed(buffer_0_167); // @[Modules.scala 50:57:@39669.4]
  assign _T_87742 = _T_87741[10:0]; // @[Modules.scala 50:57:@39670.4]
  assign buffer_10_475 = $signed(_T_87742); // @[Modules.scala 50:57:@39671.4]
  assign _T_87756 = $signed(buffer_0_176) + $signed(buffer_2_177); // @[Modules.scala 50:57:@39689.4]
  assign _T_87757 = _T_87756[10:0]; // @[Modules.scala 50:57:@39690.4]
  assign buffer_10_480 = $signed(_T_87757); // @[Modules.scala 50:57:@39691.4]
  assign _T_87777 = $signed(buffer_1_190) + $signed(buffer_0_191); // @[Modules.scala 50:57:@39717.4]
  assign _T_87778 = _T_87777[10:0]; // @[Modules.scala 50:57:@39718.4]
  assign buffer_10_487 = $signed(_T_87778); // @[Modules.scala 50:57:@39719.4]
  assign buffer_10_193 = {{6{_T_86609[4]}},_T_86609}; // @[Modules.scala 32:22:@8.4]
  assign _T_87780 = $signed(buffer_0_192) + $signed(buffer_10_193); // @[Modules.scala 50:57:@39721.4]
  assign _T_87781 = _T_87780[10:0]; // @[Modules.scala 50:57:@39722.4]
  assign buffer_10_488 = $signed(_T_87781); // @[Modules.scala 50:57:@39723.4]
  assign buffer_10_203 = {{6{_T_86659[4]}},_T_86659}; // @[Modules.scala 32:22:@8.4]
  assign _T_87795 = $signed(buffer_0_202) + $signed(buffer_10_203); // @[Modules.scala 50:57:@39741.4]
  assign _T_87796 = _T_87795[10:0]; // @[Modules.scala 50:57:@39742.4]
  assign buffer_10_493 = $signed(_T_87796); // @[Modules.scala 50:57:@39743.4]
  assign _T_87801 = $signed(buffer_3_206) + $signed(buffer_0_207); // @[Modules.scala 50:57:@39749.4]
  assign _T_87802 = _T_87801[10:0]; // @[Modules.scala 50:57:@39750.4]
  assign buffer_10_495 = $signed(_T_87802); // @[Modules.scala 50:57:@39751.4]
  assign _T_87804 = $signed(buffer_4_208) + $signed(buffer_3_209); // @[Modules.scala 50:57:@39753.4]
  assign _T_87805 = _T_87804[10:0]; // @[Modules.scala 50:57:@39754.4]
  assign buffer_10_496 = $signed(_T_87805); // @[Modules.scala 50:57:@39755.4]
  assign _T_87822 = $signed(buffer_1_220) + $signed(buffer_6_221); // @[Modules.scala 50:57:@39777.4]
  assign _T_87823 = _T_87822[10:0]; // @[Modules.scala 50:57:@39778.4]
  assign buffer_10_502 = $signed(_T_87823); // @[Modules.scala 50:57:@39779.4]
  assign _T_87831 = $signed(buffer_9_226) + $signed(buffer_4_227); // @[Modules.scala 50:57:@39789.4]
  assign _T_87832 = _T_87831[10:0]; // @[Modules.scala 50:57:@39790.4]
  assign buffer_10_505 = $signed(_T_87832); // @[Modules.scala 50:57:@39791.4]
  assign buffer_10_230 = {{6{_T_86776[4]}},_T_86776}; // @[Modules.scala 32:22:@8.4]
  assign _T_87837 = $signed(buffer_10_230) + $signed(buffer_5_231); // @[Modules.scala 50:57:@39797.4]
  assign _T_87838 = _T_87837[10:0]; // @[Modules.scala 50:57:@39798.4]
  assign buffer_10_507 = $signed(_T_87838); // @[Modules.scala 50:57:@39799.4]
  assign _T_87843 = $signed(buffer_1_234) + $signed(buffer_6_235); // @[Modules.scala 50:57:@39805.4]
  assign _T_87844 = _T_87843[10:0]; // @[Modules.scala 50:57:@39806.4]
  assign buffer_10_509 = $signed(_T_87844); // @[Modules.scala 50:57:@39807.4]
  assign _T_87858 = $signed(buffer_1_244) + $signed(buffer_9_245); // @[Modules.scala 50:57:@39825.4]
  assign _T_87859 = _T_87858[10:0]; // @[Modules.scala 50:57:@39826.4]
  assign buffer_10_514 = $signed(_T_87859); // @[Modules.scala 50:57:@39827.4]
  assign _T_87861 = $signed(buffer_4_246) + $signed(buffer_1_247); // @[Modules.scala 50:57:@39829.4]
  assign _T_87862 = _T_87861[10:0]; // @[Modules.scala 50:57:@39830.4]
  assign buffer_10_515 = $signed(_T_87862); // @[Modules.scala 50:57:@39831.4]
  assign buffer_10_255 = {{6{_T_86875[4]}},_T_86875}; // @[Modules.scala 32:22:@8.4]
  assign _T_87873 = $signed(buffer_1_254) + $signed(buffer_10_255); // @[Modules.scala 50:57:@39845.4]
  assign _T_87874 = _T_87873[10:0]; // @[Modules.scala 50:57:@39846.4]
  assign buffer_10_519 = $signed(_T_87874); // @[Modules.scala 50:57:@39847.4]
  assign _T_87876 = $signed(buffer_4_256) + $signed(buffer_0_257); // @[Modules.scala 50:57:@39849.4]
  assign _T_87877 = _T_87876[10:0]; // @[Modules.scala 50:57:@39850.4]
  assign buffer_10_520 = $signed(_T_87877); // @[Modules.scala 50:57:@39851.4]
  assign _T_87879 = $signed(buffer_2_258) + $signed(buffer_1_259); // @[Modules.scala 50:57:@39853.4]
  assign _T_87880 = _T_87879[10:0]; // @[Modules.scala 50:57:@39854.4]
  assign buffer_10_521 = $signed(_T_87880); // @[Modules.scala 50:57:@39855.4]
  assign _T_87897 = $signed(buffer_5_270) + $signed(buffer_1_271); // @[Modules.scala 50:57:@39877.4]
  assign _T_87898 = _T_87897[10:0]; // @[Modules.scala 50:57:@39878.4]
  assign buffer_10_527 = $signed(_T_87898); // @[Modules.scala 50:57:@39879.4]
  assign _T_87918 = $signed(buffer_1_284) + $signed(buffer_0_285); // @[Modules.scala 50:57:@39905.4]
  assign _T_87919 = _T_87918[10:0]; // @[Modules.scala 50:57:@39906.4]
  assign buffer_10_534 = $signed(_T_87919); // @[Modules.scala 50:57:@39907.4]
  assign _T_87927 = $signed(buffer_4_290) + $signed(buffer_5_291); // @[Modules.scala 50:57:@39917.4]
  assign _T_87928 = _T_87927[10:0]; // @[Modules.scala 50:57:@39918.4]
  assign buffer_10_537 = $signed(_T_87928); // @[Modules.scala 50:57:@39919.4]
  assign _T_87948 = $signed(buffer_2_304) + $signed(buffer_9_305); // @[Modules.scala 50:57:@39945.4]
  assign _T_87949 = _T_87948[10:0]; // @[Modules.scala 50:57:@39946.4]
  assign buffer_10_544 = $signed(_T_87949); // @[Modules.scala 50:57:@39947.4]
  assign _T_87951 = $signed(buffer_0_306) + $signed(buffer_4_307); // @[Modules.scala 50:57:@39949.4]
  assign _T_87952 = _T_87951[10:0]; // @[Modules.scala 50:57:@39950.4]
  assign buffer_10_545 = $signed(_T_87952); // @[Modules.scala 50:57:@39951.4]
  assign buffer_10_318 = {{6{_T_87128[4]}},_T_87128}; // @[Modules.scala 32:22:@8.4]
  assign _T_87969 = $signed(buffer_10_318) + $signed(buffer_0_319); // @[Modules.scala 50:57:@39973.4]
  assign _T_87970 = _T_87969[10:0]; // @[Modules.scala 50:57:@39974.4]
  assign buffer_10_551 = $signed(_T_87970); // @[Modules.scala 50:57:@39975.4]
  assign _T_87972 = $signed(buffer_9_320) + $signed(buffer_1_321); // @[Modules.scala 50:57:@39977.4]
  assign _T_87973 = _T_87972[10:0]; // @[Modules.scala 50:57:@39978.4]
  assign buffer_10_552 = $signed(_T_87973); // @[Modules.scala 50:57:@39979.4]
  assign buffer_10_322 = {{6{_T_87148[4]}},_T_87148}; // @[Modules.scala 32:22:@8.4]
  assign _T_87975 = $signed(buffer_10_322) + $signed(buffer_0_323); // @[Modules.scala 50:57:@39981.4]
  assign _T_87976 = _T_87975[10:0]; // @[Modules.scala 50:57:@39982.4]
  assign buffer_10_553 = $signed(_T_87976); // @[Modules.scala 50:57:@39983.4]
  assign _T_87981 = $signed(buffer_1_326) + $signed(buffer_6_327); // @[Modules.scala 50:57:@39989.4]
  assign _T_87982 = _T_87981[10:0]; // @[Modules.scala 50:57:@39990.4]
  assign buffer_10_555 = $signed(_T_87982); // @[Modules.scala 50:57:@39991.4]
  assign _T_88005 = $signed(buffer_2_342) + $signed(buffer_1_343); // @[Modules.scala 50:57:@40021.4]
  assign _T_88006 = _T_88005[10:0]; // @[Modules.scala 50:57:@40022.4]
  assign buffer_10_563 = $signed(_T_88006); // @[Modules.scala 50:57:@40023.4]
  assign buffer_10_353 = {{6{_T_87293[4]}},_T_87293}; // @[Modules.scala 32:22:@8.4]
  assign _T_88020 = $signed(buffer_2_352) + $signed(buffer_10_353); // @[Modules.scala 50:57:@40041.4]
  assign _T_88021 = _T_88020[10:0]; // @[Modules.scala 50:57:@40042.4]
  assign buffer_10_568 = $signed(_T_88021); // @[Modules.scala 50:57:@40043.4]
  assign buffer_10_368 = {{6{_T_87382[4]}},_T_87382}; // @[Modules.scala 32:22:@8.4]
  assign _T_88044 = $signed(buffer_10_368) + $signed(buffer_0_369); // @[Modules.scala 50:57:@40073.4]
  assign _T_88045 = _T_88044[10:0]; // @[Modules.scala 50:57:@40074.4]
  assign buffer_10_576 = $signed(_T_88045); // @[Modules.scala 50:57:@40075.4]
  assign _T_88056 = $signed(buffer_4_376) + $signed(buffer_9_377); // @[Modules.scala 50:57:@40089.4]
  assign _T_88057 = _T_88056[10:0]; // @[Modules.scala 50:57:@40090.4]
  assign buffer_10_580 = $signed(_T_88057); // @[Modules.scala 50:57:@40091.4]
  assign _T_88059 = $signed(buffer_3_378) + $signed(buffer_1_379); // @[Modules.scala 50:57:@40093.4]
  assign _T_88060 = _T_88059[10:0]; // @[Modules.scala 50:57:@40094.4]
  assign buffer_10_581 = $signed(_T_88060); // @[Modules.scala 50:57:@40095.4]
  assign _T_88062 = $signed(buffer_7_380) + $signed(buffer_1_381); // @[Modules.scala 50:57:@40097.4]
  assign _T_88063 = _T_88062[10:0]; // @[Modules.scala 50:57:@40098.4]
  assign buffer_10_582 = $signed(_T_88063); // @[Modules.scala 50:57:@40099.4]
  assign _T_88077 = $signed(buffer_7_390) + $signed(buffer_0_391); // @[Modules.scala 50:57:@40117.4]
  assign _T_88078 = _T_88077[10:0]; // @[Modules.scala 50:57:@40118.4]
  assign buffer_10_587 = $signed(_T_88078); // @[Modules.scala 50:57:@40119.4]
  assign _T_88080 = $signed(buffer_0_392) + $signed(buffer_10_393); // @[Modules.scala 53:83:@40121.4]
  assign _T_88081 = _T_88080[10:0]; // @[Modules.scala 53:83:@40122.4]
  assign buffer_10_588 = $signed(_T_88081); // @[Modules.scala 53:83:@40123.4]
  assign _T_88083 = $signed(buffer_10_394) + $signed(buffer_4_395); // @[Modules.scala 53:83:@40125.4]
  assign _T_88084 = _T_88083[10:0]; // @[Modules.scala 53:83:@40126.4]
  assign buffer_10_589 = $signed(_T_88084); // @[Modules.scala 53:83:@40127.4]
  assign _T_88089 = $signed(buffer_10_398) + $signed(buffer_1_399); // @[Modules.scala 53:83:@40133.4]
  assign _T_88090 = _T_88089[10:0]; // @[Modules.scala 53:83:@40134.4]
  assign buffer_10_591 = $signed(_T_88090); // @[Modules.scala 53:83:@40135.4]
  assign _T_88098 = $signed(buffer_1_404) + $signed(buffer_10_405); // @[Modules.scala 53:83:@40145.4]
  assign _T_88099 = _T_88098[10:0]; // @[Modules.scala 53:83:@40146.4]
  assign buffer_10_594 = $signed(_T_88099); // @[Modules.scala 53:83:@40147.4]
  assign _T_88101 = $signed(buffer_2_406) + $signed(buffer_10_407); // @[Modules.scala 53:83:@40149.4]
  assign _T_88102 = _T_88101[10:0]; // @[Modules.scala 53:83:@40150.4]
  assign buffer_10_595 = $signed(_T_88102); // @[Modules.scala 53:83:@40151.4]
  assign _T_88110 = $signed(buffer_9_412) + $signed(buffer_10_413); // @[Modules.scala 53:83:@40161.4]
  assign _T_88111 = _T_88110[10:0]; // @[Modules.scala 53:83:@40162.4]
  assign buffer_10_598 = $signed(_T_88111); // @[Modules.scala 53:83:@40163.4]
  assign _T_88119 = $signed(buffer_0_418) + $signed(buffer_10_419); // @[Modules.scala 53:83:@40173.4]
  assign _T_88120 = _T_88119[10:0]; // @[Modules.scala 53:83:@40174.4]
  assign buffer_10_601 = $signed(_T_88120); // @[Modules.scala 53:83:@40175.4]
  assign _T_88122 = $signed(buffer_10_420) + $signed(buffer_7_421); // @[Modules.scala 53:83:@40177.4]
  assign _T_88123 = _T_88122[10:0]; // @[Modules.scala 53:83:@40178.4]
  assign buffer_10_602 = $signed(_T_88123); // @[Modules.scala 53:83:@40179.4]
  assign _T_88125 = $signed(buffer_4_422) + $signed(buffer_3_423); // @[Modules.scala 53:83:@40181.4]
  assign _T_88126 = _T_88125[10:0]; // @[Modules.scala 53:83:@40182.4]
  assign buffer_10_603 = $signed(_T_88126); // @[Modules.scala 53:83:@40183.4]
  assign _T_88128 = $signed(buffer_10_424) + $signed(buffer_0_425); // @[Modules.scala 53:83:@40185.4]
  assign _T_88129 = _T_88128[10:0]; // @[Modules.scala 53:83:@40186.4]
  assign buffer_10_604 = $signed(_T_88129); // @[Modules.scala 53:83:@40187.4]
  assign _T_88131 = $signed(buffer_10_426) + $signed(buffer_10_427); // @[Modules.scala 53:83:@40189.4]
  assign _T_88132 = _T_88131[10:0]; // @[Modules.scala 53:83:@40190.4]
  assign buffer_10_605 = $signed(_T_88132); // @[Modules.scala 53:83:@40191.4]
  assign _T_88134 = $signed(buffer_4_428) + $signed(buffer_10_429); // @[Modules.scala 53:83:@40193.4]
  assign _T_88135 = _T_88134[10:0]; // @[Modules.scala 53:83:@40194.4]
  assign buffer_10_606 = $signed(_T_88135); // @[Modules.scala 53:83:@40195.4]
  assign _T_88137 = $signed(buffer_10_430) + $signed(buffer_10_431); // @[Modules.scala 53:83:@40197.4]
  assign _T_88138 = _T_88137[10:0]; // @[Modules.scala 53:83:@40198.4]
  assign buffer_10_607 = $signed(_T_88138); // @[Modules.scala 53:83:@40199.4]
  assign _T_88140 = $signed(buffer_10_432) + $signed(buffer_10_433); // @[Modules.scala 53:83:@40201.4]
  assign _T_88141 = _T_88140[10:0]; // @[Modules.scala 53:83:@40202.4]
  assign buffer_10_608 = $signed(_T_88141); // @[Modules.scala 53:83:@40203.4]
  assign _T_88143 = $signed(buffer_10_434) + $signed(buffer_10_435); // @[Modules.scala 53:83:@40205.4]
  assign _T_88144 = _T_88143[10:0]; // @[Modules.scala 53:83:@40206.4]
  assign buffer_10_609 = $signed(_T_88144); // @[Modules.scala 53:83:@40207.4]
  assign _T_88146 = $signed(buffer_10_436) + $signed(buffer_1_437); // @[Modules.scala 53:83:@40209.4]
  assign _T_88147 = _T_88146[10:0]; // @[Modules.scala 53:83:@40210.4]
  assign buffer_10_610 = $signed(_T_88147); // @[Modules.scala 53:83:@40211.4]
  assign _T_88149 = $signed(buffer_2_438) + $signed(buffer_9_439); // @[Modules.scala 53:83:@40213.4]
  assign _T_88150 = _T_88149[10:0]; // @[Modules.scala 53:83:@40214.4]
  assign buffer_10_611 = $signed(_T_88150); // @[Modules.scala 53:83:@40215.4]
  assign _T_88152 = $signed(buffer_10_440) + $signed(buffer_3_441); // @[Modules.scala 53:83:@40217.4]
  assign _T_88153 = _T_88152[10:0]; // @[Modules.scala 53:83:@40218.4]
  assign buffer_10_612 = $signed(_T_88153); // @[Modules.scala 53:83:@40219.4]
  assign _T_88155 = $signed(buffer_10_442) + $signed(buffer_10_443); // @[Modules.scala 53:83:@40221.4]
  assign _T_88156 = _T_88155[10:0]; // @[Modules.scala 53:83:@40222.4]
  assign buffer_10_613 = $signed(_T_88156); // @[Modules.scala 53:83:@40223.4]
  assign _T_88158 = $signed(buffer_10_444) + $signed(buffer_0_445); // @[Modules.scala 53:83:@40225.4]
  assign _T_88159 = _T_88158[10:0]; // @[Modules.scala 53:83:@40226.4]
  assign buffer_10_614 = $signed(_T_88159); // @[Modules.scala 53:83:@40227.4]
  assign _T_88161 = $signed(buffer_0_446) + $signed(buffer_5_447); // @[Modules.scala 53:83:@40229.4]
  assign _T_88162 = _T_88161[10:0]; // @[Modules.scala 53:83:@40230.4]
  assign buffer_10_615 = $signed(_T_88162); // @[Modules.scala 53:83:@40231.4]
  assign _T_88164 = $signed(buffer_3_448) + $signed(buffer_10_449); // @[Modules.scala 53:83:@40233.4]
  assign _T_88165 = _T_88164[10:0]; // @[Modules.scala 53:83:@40234.4]
  assign buffer_10_616 = $signed(_T_88165); // @[Modules.scala 53:83:@40235.4]
  assign _T_88167 = $signed(buffer_0_450) + $signed(buffer_10_451); // @[Modules.scala 53:83:@40237.4]
  assign _T_88168 = _T_88167[10:0]; // @[Modules.scala 53:83:@40238.4]
  assign buffer_10_617 = $signed(_T_88168); // @[Modules.scala 53:83:@40239.4]
  assign _T_88173 = $signed(buffer_0_454) + $signed(buffer_3_455); // @[Modules.scala 53:83:@40245.4]
  assign _T_88174 = _T_88173[10:0]; // @[Modules.scala 53:83:@40246.4]
  assign buffer_10_619 = $signed(_T_88174); // @[Modules.scala 53:83:@40247.4]
  assign _T_88176 = $signed(buffer_3_456) + $signed(buffer_8_457); // @[Modules.scala 53:83:@40249.4]
  assign _T_88177 = _T_88176[10:0]; // @[Modules.scala 53:83:@40250.4]
  assign buffer_10_620 = $signed(_T_88177); // @[Modules.scala 53:83:@40251.4]
  assign _T_88185 = $signed(buffer_9_462) + $signed(buffer_0_463); // @[Modules.scala 53:83:@40261.4]
  assign _T_88186 = _T_88185[10:0]; // @[Modules.scala 53:83:@40262.4]
  assign buffer_10_623 = $signed(_T_88186); // @[Modules.scala 53:83:@40263.4]
  assign _T_88194 = $signed(buffer_5_468) + $signed(buffer_10_469); // @[Modules.scala 53:83:@40273.4]
  assign _T_88195 = _T_88194[10:0]; // @[Modules.scala 53:83:@40274.4]
  assign buffer_10_626 = $signed(_T_88195); // @[Modules.scala 53:83:@40275.4]
  assign _T_88200 = $signed(buffer_5_472) + $signed(buffer_10_473); // @[Modules.scala 53:83:@40281.4]
  assign _T_88201 = _T_88200[10:0]; // @[Modules.scala 53:83:@40282.4]
  assign buffer_10_628 = $signed(_T_88201); // @[Modules.scala 53:83:@40283.4]
  assign _T_88203 = $signed(buffer_2_474) + $signed(buffer_10_475); // @[Modules.scala 53:83:@40285.4]
  assign _T_88204 = _T_88203[10:0]; // @[Modules.scala 53:83:@40286.4]
  assign buffer_10_629 = $signed(_T_88204); // @[Modules.scala 53:83:@40287.4]
  assign _T_88212 = $signed(buffer_10_480) + $signed(buffer_5_481); // @[Modules.scala 53:83:@40297.4]
  assign _T_88213 = _T_88212[10:0]; // @[Modules.scala 53:83:@40298.4]
  assign buffer_10_632 = $signed(_T_88213); // @[Modules.scala 53:83:@40299.4]
  assign _T_88215 = $signed(buffer_4_482) + $signed(buffer_6_483); // @[Modules.scala 53:83:@40301.4]
  assign _T_88216 = _T_88215[10:0]; // @[Modules.scala 53:83:@40302.4]
  assign buffer_10_633 = $signed(_T_88216); // @[Modules.scala 53:83:@40303.4]
  assign _T_88221 = $signed(buffer_5_486) + $signed(buffer_10_487); // @[Modules.scala 53:83:@40309.4]
  assign _T_88222 = _T_88221[10:0]; // @[Modules.scala 53:83:@40310.4]
  assign buffer_10_635 = $signed(_T_88222); // @[Modules.scala 53:83:@40311.4]
  assign _T_88224 = $signed(buffer_10_488) + $signed(buffer_9_489); // @[Modules.scala 53:83:@40313.4]
  assign _T_88225 = _T_88224[10:0]; // @[Modules.scala 53:83:@40314.4]
  assign buffer_10_636 = $signed(_T_88225); // @[Modules.scala 53:83:@40315.4]
  assign _T_88227 = $signed(buffer_7_490) + $signed(buffer_3_491); // @[Modules.scala 53:83:@40317.4]
  assign _T_88228 = _T_88227[10:0]; // @[Modules.scala 53:83:@40318.4]
  assign buffer_10_637 = $signed(_T_88228); // @[Modules.scala 53:83:@40319.4]
  assign _T_88230 = $signed(buffer_6_492) + $signed(buffer_10_493); // @[Modules.scala 53:83:@40321.4]
  assign _T_88231 = _T_88230[10:0]; // @[Modules.scala 53:83:@40322.4]
  assign buffer_10_638 = $signed(_T_88231); // @[Modules.scala 53:83:@40323.4]
  assign _T_88233 = $signed(buffer_7_494) + $signed(buffer_10_495); // @[Modules.scala 53:83:@40325.4]
  assign _T_88234 = _T_88233[10:0]; // @[Modules.scala 53:83:@40326.4]
  assign buffer_10_639 = $signed(_T_88234); // @[Modules.scala 53:83:@40327.4]
  assign _T_88236 = $signed(buffer_10_496) + $signed(buffer_3_497); // @[Modules.scala 53:83:@40329.4]
  assign _T_88237 = _T_88236[10:0]; // @[Modules.scala 53:83:@40330.4]
  assign buffer_10_640 = $signed(_T_88237); // @[Modules.scala 53:83:@40331.4]
  assign _T_88239 = $signed(buffer_9_498) + $signed(buffer_5_499); // @[Modules.scala 53:83:@40333.4]
  assign _T_88240 = _T_88239[10:0]; // @[Modules.scala 53:83:@40334.4]
  assign buffer_10_641 = $signed(_T_88240); // @[Modules.scala 53:83:@40335.4]
  assign _T_88242 = $signed(buffer_0_500) + $signed(buffer_1_501); // @[Modules.scala 53:83:@40337.4]
  assign _T_88243 = _T_88242[10:0]; // @[Modules.scala 53:83:@40338.4]
  assign buffer_10_642 = $signed(_T_88243); // @[Modules.scala 53:83:@40339.4]
  assign _T_88245 = $signed(buffer_10_502) + $signed(buffer_3_503); // @[Modules.scala 53:83:@40341.4]
  assign _T_88246 = _T_88245[10:0]; // @[Modules.scala 53:83:@40342.4]
  assign buffer_10_643 = $signed(_T_88246); // @[Modules.scala 53:83:@40343.4]
  assign _T_88248 = $signed(buffer_9_504) + $signed(buffer_10_505); // @[Modules.scala 53:83:@40345.4]
  assign _T_88249 = _T_88248[10:0]; // @[Modules.scala 53:83:@40346.4]
  assign buffer_10_644 = $signed(_T_88249); // @[Modules.scala 53:83:@40347.4]
  assign _T_88251 = $signed(buffer_1_506) + $signed(buffer_10_507); // @[Modules.scala 53:83:@40349.4]
  assign _T_88252 = _T_88251[10:0]; // @[Modules.scala 53:83:@40350.4]
  assign buffer_10_645 = $signed(_T_88252); // @[Modules.scala 53:83:@40351.4]
  assign _T_88254 = $signed(buffer_3_508) + $signed(buffer_10_509); // @[Modules.scala 53:83:@40353.4]
  assign _T_88255 = _T_88254[10:0]; // @[Modules.scala 53:83:@40354.4]
  assign buffer_10_646 = $signed(_T_88255); // @[Modules.scala 53:83:@40355.4]
  assign _T_88260 = $signed(buffer_4_512) + $signed(buffer_1_513); // @[Modules.scala 53:83:@40361.4]
  assign _T_88261 = _T_88260[10:0]; // @[Modules.scala 53:83:@40362.4]
  assign buffer_10_648 = $signed(_T_88261); // @[Modules.scala 53:83:@40363.4]
  assign _T_88263 = $signed(buffer_10_514) + $signed(buffer_10_515); // @[Modules.scala 53:83:@40365.4]
  assign _T_88264 = _T_88263[10:0]; // @[Modules.scala 53:83:@40366.4]
  assign buffer_10_649 = $signed(_T_88264); // @[Modules.scala 53:83:@40367.4]
  assign _T_88269 = $signed(buffer_4_518) + $signed(buffer_10_519); // @[Modules.scala 53:83:@40373.4]
  assign _T_88270 = _T_88269[10:0]; // @[Modules.scala 53:83:@40374.4]
  assign buffer_10_651 = $signed(_T_88270); // @[Modules.scala 53:83:@40375.4]
  assign _T_88272 = $signed(buffer_10_520) + $signed(buffer_10_521); // @[Modules.scala 53:83:@40377.4]
  assign _T_88273 = _T_88272[10:0]; // @[Modules.scala 53:83:@40378.4]
  assign buffer_10_652 = $signed(_T_88273); // @[Modules.scala 53:83:@40379.4]
  assign _T_88275 = $signed(buffer_1_522) + $signed(buffer_4_523); // @[Modules.scala 53:83:@40381.4]
  assign _T_88276 = _T_88275[10:0]; // @[Modules.scala 53:83:@40382.4]
  assign buffer_10_653 = $signed(_T_88276); // @[Modules.scala 53:83:@40383.4]
  assign _T_88281 = $signed(buffer_9_526) + $signed(buffer_10_527); // @[Modules.scala 53:83:@40389.4]
  assign _T_88282 = _T_88281[10:0]; // @[Modules.scala 53:83:@40390.4]
  assign buffer_10_655 = $signed(_T_88282); // @[Modules.scala 53:83:@40391.4]
  assign _T_88284 = $signed(buffer_7_528) + $signed(buffer_1_529); // @[Modules.scala 53:83:@40393.4]
  assign _T_88285 = _T_88284[10:0]; // @[Modules.scala 53:83:@40394.4]
  assign buffer_10_656 = $signed(_T_88285); // @[Modules.scala 53:83:@40395.4]
  assign _T_88287 = $signed(buffer_3_530) + $signed(buffer_5_531); // @[Modules.scala 53:83:@40397.4]
  assign _T_88288 = _T_88287[10:0]; // @[Modules.scala 53:83:@40398.4]
  assign buffer_10_657 = $signed(_T_88288); // @[Modules.scala 53:83:@40399.4]
  assign _T_88290 = $signed(buffer_8_532) + $signed(buffer_3_533); // @[Modules.scala 53:83:@40401.4]
  assign _T_88291 = _T_88290[10:0]; // @[Modules.scala 53:83:@40402.4]
  assign buffer_10_658 = $signed(_T_88291); // @[Modules.scala 53:83:@40403.4]
  assign _T_88293 = $signed(buffer_10_534) + $signed(buffer_5_535); // @[Modules.scala 53:83:@40405.4]
  assign _T_88294 = _T_88293[10:0]; // @[Modules.scala 53:83:@40406.4]
  assign buffer_10_659 = $signed(_T_88294); // @[Modules.scala 53:83:@40407.4]
  assign _T_88296 = $signed(buffer_2_536) + $signed(buffer_10_537); // @[Modules.scala 53:83:@40409.4]
  assign _T_88297 = _T_88296[10:0]; // @[Modules.scala 53:83:@40410.4]
  assign buffer_10_660 = $signed(_T_88297); // @[Modules.scala 53:83:@40411.4]
  assign _T_88308 = $signed(buffer_10_544) + $signed(buffer_10_545); // @[Modules.scala 53:83:@40425.4]
  assign _T_88309 = _T_88308[10:0]; // @[Modules.scala 53:83:@40426.4]
  assign buffer_10_664 = $signed(_T_88309); // @[Modules.scala 53:83:@40427.4]
  assign _T_88314 = $signed(buffer_6_548) + $signed(buffer_8_549); // @[Modules.scala 53:83:@40433.4]
  assign _T_88315 = _T_88314[10:0]; // @[Modules.scala 53:83:@40434.4]
  assign buffer_10_666 = $signed(_T_88315); // @[Modules.scala 53:83:@40435.4]
  assign _T_88317 = $signed(buffer_2_550) + $signed(buffer_10_551); // @[Modules.scala 53:83:@40437.4]
  assign _T_88318 = _T_88317[10:0]; // @[Modules.scala 53:83:@40438.4]
  assign buffer_10_667 = $signed(_T_88318); // @[Modules.scala 53:83:@40439.4]
  assign _T_88320 = $signed(buffer_10_552) + $signed(buffer_10_553); // @[Modules.scala 53:83:@40441.4]
  assign _T_88321 = _T_88320[10:0]; // @[Modules.scala 53:83:@40442.4]
  assign buffer_10_668 = $signed(_T_88321); // @[Modules.scala 53:83:@40443.4]
  assign _T_88323 = $signed(buffer_1_554) + $signed(buffer_10_555); // @[Modules.scala 53:83:@40445.4]
  assign _T_88324 = _T_88323[10:0]; // @[Modules.scala 53:83:@40446.4]
  assign buffer_10_669 = $signed(_T_88324); // @[Modules.scala 53:83:@40447.4]
  assign _T_88335 = $signed(buffer_3_562) + $signed(buffer_10_563); // @[Modules.scala 53:83:@40461.4]
  assign _T_88336 = _T_88335[10:0]; // @[Modules.scala 53:83:@40462.4]
  assign buffer_10_673 = $signed(_T_88336); // @[Modules.scala 53:83:@40463.4]
  assign _T_88344 = $signed(buffer_10_568) + $signed(buffer_2_569); // @[Modules.scala 53:83:@40473.4]
  assign _T_88345 = _T_88344[10:0]; // @[Modules.scala 53:83:@40474.4]
  assign buffer_10_676 = $signed(_T_88345); // @[Modules.scala 53:83:@40475.4]
  assign _T_88350 = $signed(buffer_3_572) + $signed(buffer_1_573); // @[Modules.scala 53:83:@40481.4]
  assign _T_88351 = _T_88350[10:0]; // @[Modules.scala 53:83:@40482.4]
  assign buffer_10_678 = $signed(_T_88351); // @[Modules.scala 53:83:@40483.4]
  assign _T_88353 = $signed(buffer_3_574) + $signed(buffer_1_575); // @[Modules.scala 53:83:@40485.4]
  assign _T_88354 = _T_88353[10:0]; // @[Modules.scala 53:83:@40486.4]
  assign buffer_10_679 = $signed(_T_88354); // @[Modules.scala 53:83:@40487.4]
  assign _T_88356 = $signed(buffer_10_576) + $signed(buffer_1_577); // @[Modules.scala 53:83:@40489.4]
  assign _T_88357 = _T_88356[10:0]; // @[Modules.scala 53:83:@40490.4]
  assign buffer_10_680 = $signed(_T_88357); // @[Modules.scala 53:83:@40491.4]
  assign _T_88362 = $signed(buffer_10_580) + $signed(buffer_10_581); // @[Modules.scala 53:83:@40497.4]
  assign _T_88363 = _T_88362[10:0]; // @[Modules.scala 53:83:@40498.4]
  assign buffer_10_682 = $signed(_T_88363); // @[Modules.scala 53:83:@40499.4]
  assign _T_88365 = $signed(buffer_10_582) + $signed(buffer_3_583); // @[Modules.scala 53:83:@40501.4]
  assign _T_88366 = _T_88365[10:0]; // @[Modules.scala 53:83:@40502.4]
  assign buffer_10_683 = $signed(_T_88366); // @[Modules.scala 53:83:@40503.4]
  assign _T_88371 = $signed(buffer_5_586) + $signed(buffer_10_587); // @[Modules.scala 53:83:@40509.4]
  assign _T_88372 = _T_88371[10:0]; // @[Modules.scala 53:83:@40510.4]
  assign buffer_10_685 = $signed(_T_88372); // @[Modules.scala 53:83:@40511.4]
  assign _T_88374 = $signed(buffer_10_588) + $signed(buffer_10_589); // @[Modules.scala 56:109:@40513.4]
  assign _T_88375 = _T_88374[10:0]; // @[Modules.scala 56:109:@40514.4]
  assign buffer_10_686 = $signed(_T_88375); // @[Modules.scala 56:109:@40515.4]
  assign _T_88377 = $signed(buffer_9_590) + $signed(buffer_10_591); // @[Modules.scala 56:109:@40517.4]
  assign _T_88378 = _T_88377[10:0]; // @[Modules.scala 56:109:@40518.4]
  assign buffer_10_687 = $signed(_T_88378); // @[Modules.scala 56:109:@40519.4]
  assign _T_88383 = $signed(buffer_10_594) + $signed(buffer_10_595); // @[Modules.scala 56:109:@40525.4]
  assign _T_88384 = _T_88383[10:0]; // @[Modules.scala 56:109:@40526.4]
  assign buffer_10_689 = $signed(_T_88384); // @[Modules.scala 56:109:@40527.4]
  assign _T_88389 = $signed(buffer_10_598) + $signed(buffer_1_599); // @[Modules.scala 56:109:@40533.4]
  assign _T_88390 = _T_88389[10:0]; // @[Modules.scala 56:109:@40534.4]
  assign buffer_10_691 = $signed(_T_88390); // @[Modules.scala 56:109:@40535.4]
  assign _T_88392 = $signed(buffer_1_600) + $signed(buffer_10_601); // @[Modules.scala 56:109:@40537.4]
  assign _T_88393 = _T_88392[10:0]; // @[Modules.scala 56:109:@40538.4]
  assign buffer_10_692 = $signed(_T_88393); // @[Modules.scala 56:109:@40539.4]
  assign _T_88395 = $signed(buffer_10_602) + $signed(buffer_10_603); // @[Modules.scala 56:109:@40541.4]
  assign _T_88396 = _T_88395[10:0]; // @[Modules.scala 56:109:@40542.4]
  assign buffer_10_693 = $signed(_T_88396); // @[Modules.scala 56:109:@40543.4]
  assign _T_88398 = $signed(buffer_10_604) + $signed(buffer_10_605); // @[Modules.scala 56:109:@40545.4]
  assign _T_88399 = _T_88398[10:0]; // @[Modules.scala 56:109:@40546.4]
  assign buffer_10_694 = $signed(_T_88399); // @[Modules.scala 56:109:@40547.4]
  assign _T_88401 = $signed(buffer_10_606) + $signed(buffer_10_607); // @[Modules.scala 56:109:@40549.4]
  assign _T_88402 = _T_88401[10:0]; // @[Modules.scala 56:109:@40550.4]
  assign buffer_10_695 = $signed(_T_88402); // @[Modules.scala 56:109:@40551.4]
  assign _T_88404 = $signed(buffer_10_608) + $signed(buffer_10_609); // @[Modules.scala 56:109:@40553.4]
  assign _T_88405 = _T_88404[10:0]; // @[Modules.scala 56:109:@40554.4]
  assign buffer_10_696 = $signed(_T_88405); // @[Modules.scala 56:109:@40555.4]
  assign _T_88407 = $signed(buffer_10_610) + $signed(buffer_10_611); // @[Modules.scala 56:109:@40557.4]
  assign _T_88408 = _T_88407[10:0]; // @[Modules.scala 56:109:@40558.4]
  assign buffer_10_697 = $signed(_T_88408); // @[Modules.scala 56:109:@40559.4]
  assign _T_88410 = $signed(buffer_10_612) + $signed(buffer_10_613); // @[Modules.scala 56:109:@40561.4]
  assign _T_88411 = _T_88410[10:0]; // @[Modules.scala 56:109:@40562.4]
  assign buffer_10_698 = $signed(_T_88411); // @[Modules.scala 56:109:@40563.4]
  assign _T_88413 = $signed(buffer_10_614) + $signed(buffer_10_615); // @[Modules.scala 56:109:@40565.4]
  assign _T_88414 = _T_88413[10:0]; // @[Modules.scala 56:109:@40566.4]
  assign buffer_10_699 = $signed(_T_88414); // @[Modules.scala 56:109:@40567.4]
  assign _T_88416 = $signed(buffer_10_616) + $signed(buffer_10_617); // @[Modules.scala 56:109:@40569.4]
  assign _T_88417 = _T_88416[10:0]; // @[Modules.scala 56:109:@40570.4]
  assign buffer_10_700 = $signed(_T_88417); // @[Modules.scala 56:109:@40571.4]
  assign _T_88419 = $signed(buffer_0_618) + $signed(buffer_10_619); // @[Modules.scala 56:109:@40573.4]
  assign _T_88420 = _T_88419[10:0]; // @[Modules.scala 56:109:@40574.4]
  assign buffer_10_701 = $signed(_T_88420); // @[Modules.scala 56:109:@40575.4]
  assign _T_88422 = $signed(buffer_10_620) + $signed(buffer_0_621); // @[Modules.scala 56:109:@40577.4]
  assign _T_88423 = _T_88422[10:0]; // @[Modules.scala 56:109:@40578.4]
  assign buffer_10_702 = $signed(_T_88423); // @[Modules.scala 56:109:@40579.4]
  assign _T_88425 = $signed(buffer_0_622) + $signed(buffer_10_623); // @[Modules.scala 56:109:@40581.4]
  assign _T_88426 = _T_88425[10:0]; // @[Modules.scala 56:109:@40582.4]
  assign buffer_10_703 = $signed(_T_88426); // @[Modules.scala 56:109:@40583.4]
  assign _T_88428 = $signed(buffer_5_624) + $signed(buffer_0_625); // @[Modules.scala 56:109:@40585.4]
  assign _T_88429 = _T_88428[10:0]; // @[Modules.scala 56:109:@40586.4]
  assign buffer_10_704 = $signed(_T_88429); // @[Modules.scala 56:109:@40587.4]
  assign _T_88431 = $signed(buffer_10_626) + $signed(buffer_3_627); // @[Modules.scala 56:109:@40589.4]
  assign _T_88432 = _T_88431[10:0]; // @[Modules.scala 56:109:@40590.4]
  assign buffer_10_705 = $signed(_T_88432); // @[Modules.scala 56:109:@40591.4]
  assign _T_88434 = $signed(buffer_10_628) + $signed(buffer_10_629); // @[Modules.scala 56:109:@40593.4]
  assign _T_88435 = _T_88434[10:0]; // @[Modules.scala 56:109:@40594.4]
  assign buffer_10_706 = $signed(_T_88435); // @[Modules.scala 56:109:@40595.4]
  assign _T_88440 = $signed(buffer_10_632) + $signed(buffer_10_633); // @[Modules.scala 56:109:@40601.4]
  assign _T_88441 = _T_88440[10:0]; // @[Modules.scala 56:109:@40602.4]
  assign buffer_10_708 = $signed(_T_88441); // @[Modules.scala 56:109:@40603.4]
  assign _T_88443 = $signed(buffer_9_634) + $signed(buffer_10_635); // @[Modules.scala 56:109:@40605.4]
  assign _T_88444 = _T_88443[10:0]; // @[Modules.scala 56:109:@40606.4]
  assign buffer_10_709 = $signed(_T_88444); // @[Modules.scala 56:109:@40607.4]
  assign _T_88446 = $signed(buffer_10_636) + $signed(buffer_10_637); // @[Modules.scala 56:109:@40609.4]
  assign _T_88447 = _T_88446[10:0]; // @[Modules.scala 56:109:@40610.4]
  assign buffer_10_710 = $signed(_T_88447); // @[Modules.scala 56:109:@40611.4]
  assign _T_88449 = $signed(buffer_10_638) + $signed(buffer_10_639); // @[Modules.scala 56:109:@40613.4]
  assign _T_88450 = _T_88449[10:0]; // @[Modules.scala 56:109:@40614.4]
  assign buffer_10_711 = $signed(_T_88450); // @[Modules.scala 56:109:@40615.4]
  assign _T_88452 = $signed(buffer_10_640) + $signed(buffer_10_641); // @[Modules.scala 56:109:@40617.4]
  assign _T_88453 = _T_88452[10:0]; // @[Modules.scala 56:109:@40618.4]
  assign buffer_10_712 = $signed(_T_88453); // @[Modules.scala 56:109:@40619.4]
  assign _T_88455 = $signed(buffer_10_642) + $signed(buffer_10_643); // @[Modules.scala 56:109:@40621.4]
  assign _T_88456 = _T_88455[10:0]; // @[Modules.scala 56:109:@40622.4]
  assign buffer_10_713 = $signed(_T_88456); // @[Modules.scala 56:109:@40623.4]
  assign _T_88458 = $signed(buffer_10_644) + $signed(buffer_10_645); // @[Modules.scala 56:109:@40625.4]
  assign _T_88459 = _T_88458[10:0]; // @[Modules.scala 56:109:@40626.4]
  assign buffer_10_714 = $signed(_T_88459); // @[Modules.scala 56:109:@40627.4]
  assign _T_88461 = $signed(buffer_10_646) + $signed(buffer_4_647); // @[Modules.scala 56:109:@40629.4]
  assign _T_88462 = _T_88461[10:0]; // @[Modules.scala 56:109:@40630.4]
  assign buffer_10_715 = $signed(_T_88462); // @[Modules.scala 56:109:@40631.4]
  assign _T_88464 = $signed(buffer_10_648) + $signed(buffer_10_649); // @[Modules.scala 56:109:@40633.4]
  assign _T_88465 = _T_88464[10:0]; // @[Modules.scala 56:109:@40634.4]
  assign buffer_10_716 = $signed(_T_88465); // @[Modules.scala 56:109:@40635.4]
  assign _T_88467 = $signed(buffer_3_650) + $signed(buffer_10_651); // @[Modules.scala 56:109:@40637.4]
  assign _T_88468 = _T_88467[10:0]; // @[Modules.scala 56:109:@40638.4]
  assign buffer_10_717 = $signed(_T_88468); // @[Modules.scala 56:109:@40639.4]
  assign _T_88470 = $signed(buffer_10_652) + $signed(buffer_10_653); // @[Modules.scala 56:109:@40641.4]
  assign _T_88471 = _T_88470[10:0]; // @[Modules.scala 56:109:@40642.4]
  assign buffer_10_718 = $signed(_T_88471); // @[Modules.scala 56:109:@40643.4]
  assign _T_88473 = $signed(buffer_8_654) + $signed(buffer_10_655); // @[Modules.scala 56:109:@40645.4]
  assign _T_88474 = _T_88473[10:0]; // @[Modules.scala 56:109:@40646.4]
  assign buffer_10_719 = $signed(_T_88474); // @[Modules.scala 56:109:@40647.4]
  assign _T_88476 = $signed(buffer_10_656) + $signed(buffer_10_657); // @[Modules.scala 56:109:@40649.4]
  assign _T_88477 = _T_88476[10:0]; // @[Modules.scala 56:109:@40650.4]
  assign buffer_10_720 = $signed(_T_88477); // @[Modules.scala 56:109:@40651.4]
  assign _T_88479 = $signed(buffer_10_658) + $signed(buffer_10_659); // @[Modules.scala 56:109:@40653.4]
  assign _T_88480 = _T_88479[10:0]; // @[Modules.scala 56:109:@40654.4]
  assign buffer_10_721 = $signed(_T_88480); // @[Modules.scala 56:109:@40655.4]
  assign _T_88482 = $signed(buffer_10_660) + $signed(buffer_3_661); // @[Modules.scala 56:109:@40657.4]
  assign _T_88483 = _T_88482[10:0]; // @[Modules.scala 56:109:@40658.4]
  assign buffer_10_722 = $signed(_T_88483); // @[Modules.scala 56:109:@40659.4]
  assign _T_88485 = $signed(buffer_4_662) + $signed(buffer_1_663); // @[Modules.scala 56:109:@40661.4]
  assign _T_88486 = _T_88485[10:0]; // @[Modules.scala 56:109:@40662.4]
  assign buffer_10_723 = $signed(_T_88486); // @[Modules.scala 56:109:@40663.4]
  assign _T_88488 = $signed(buffer_10_664) + $signed(buffer_5_665); // @[Modules.scala 56:109:@40665.4]
  assign _T_88489 = _T_88488[10:0]; // @[Modules.scala 56:109:@40666.4]
  assign buffer_10_724 = $signed(_T_88489); // @[Modules.scala 56:109:@40667.4]
  assign _T_88491 = $signed(buffer_10_666) + $signed(buffer_10_667); // @[Modules.scala 56:109:@40669.4]
  assign _T_88492 = _T_88491[10:0]; // @[Modules.scala 56:109:@40670.4]
  assign buffer_10_725 = $signed(_T_88492); // @[Modules.scala 56:109:@40671.4]
  assign _T_88494 = $signed(buffer_10_668) + $signed(buffer_10_669); // @[Modules.scala 56:109:@40673.4]
  assign _T_88495 = _T_88494[10:0]; // @[Modules.scala 56:109:@40674.4]
  assign buffer_10_726 = $signed(_T_88495); // @[Modules.scala 56:109:@40675.4]
  assign _T_88497 = $signed(buffer_6_670) + $signed(buffer_8_671); // @[Modules.scala 56:109:@40677.4]
  assign _T_88498 = _T_88497[10:0]; // @[Modules.scala 56:109:@40678.4]
  assign buffer_10_727 = $signed(_T_88498); // @[Modules.scala 56:109:@40679.4]
  assign _T_88500 = $signed(buffer_1_672) + $signed(buffer_10_673); // @[Modules.scala 56:109:@40681.4]
  assign _T_88501 = _T_88500[10:0]; // @[Modules.scala 56:109:@40682.4]
  assign buffer_10_728 = $signed(_T_88501); // @[Modules.scala 56:109:@40683.4]
  assign _T_88503 = $signed(buffer_3_674) + $signed(buffer_9_675); // @[Modules.scala 56:109:@40685.4]
  assign _T_88504 = _T_88503[10:0]; // @[Modules.scala 56:109:@40686.4]
  assign buffer_10_729 = $signed(_T_88504); // @[Modules.scala 56:109:@40687.4]
  assign _T_88506 = $signed(buffer_10_676) + $signed(buffer_2_677); // @[Modules.scala 56:109:@40689.4]
  assign _T_88507 = _T_88506[10:0]; // @[Modules.scala 56:109:@40690.4]
  assign buffer_10_730 = $signed(_T_88507); // @[Modules.scala 56:109:@40691.4]
  assign _T_88509 = $signed(buffer_10_678) + $signed(buffer_10_679); // @[Modules.scala 56:109:@40693.4]
  assign _T_88510 = _T_88509[10:0]; // @[Modules.scala 56:109:@40694.4]
  assign buffer_10_731 = $signed(_T_88510); // @[Modules.scala 56:109:@40695.4]
  assign _T_88512 = $signed(buffer_10_680) + $signed(buffer_4_681); // @[Modules.scala 56:109:@40697.4]
  assign _T_88513 = _T_88512[10:0]; // @[Modules.scala 56:109:@40698.4]
  assign buffer_10_732 = $signed(_T_88513); // @[Modules.scala 56:109:@40699.4]
  assign _T_88515 = $signed(buffer_10_682) + $signed(buffer_10_683); // @[Modules.scala 56:109:@40701.4]
  assign _T_88516 = _T_88515[10:0]; // @[Modules.scala 56:109:@40702.4]
  assign buffer_10_733 = $signed(_T_88516); // @[Modules.scala 56:109:@40703.4]
  assign _T_88518 = $signed(buffer_9_684) + $signed(buffer_10_685); // @[Modules.scala 56:109:@40705.4]
  assign _T_88519 = _T_88518[10:0]; // @[Modules.scala 56:109:@40706.4]
  assign buffer_10_734 = $signed(_T_88519); // @[Modules.scala 56:109:@40707.4]
  assign _T_88521 = $signed(buffer_10_686) + $signed(buffer_10_687); // @[Modules.scala 63:156:@40710.4]
  assign _T_88522 = _T_88521[10:0]; // @[Modules.scala 63:156:@40711.4]
  assign buffer_10_736 = $signed(_T_88522); // @[Modules.scala 63:156:@40712.4]
  assign _T_88524 = $signed(buffer_10_736) + $signed(buffer_9_688); // @[Modules.scala 63:156:@40714.4]
  assign _T_88525 = _T_88524[10:0]; // @[Modules.scala 63:156:@40715.4]
  assign buffer_10_737 = $signed(_T_88525); // @[Modules.scala 63:156:@40716.4]
  assign _T_88527 = $signed(buffer_10_737) + $signed(buffer_10_689); // @[Modules.scala 63:156:@40718.4]
  assign _T_88528 = _T_88527[10:0]; // @[Modules.scala 63:156:@40719.4]
  assign buffer_10_738 = $signed(_T_88528); // @[Modules.scala 63:156:@40720.4]
  assign _T_88530 = $signed(buffer_10_738) + $signed(buffer_1_690); // @[Modules.scala 63:156:@40722.4]
  assign _T_88531 = _T_88530[10:0]; // @[Modules.scala 63:156:@40723.4]
  assign buffer_10_739 = $signed(_T_88531); // @[Modules.scala 63:156:@40724.4]
  assign _T_88533 = $signed(buffer_10_739) + $signed(buffer_10_691); // @[Modules.scala 63:156:@40726.4]
  assign _T_88534 = _T_88533[10:0]; // @[Modules.scala 63:156:@40727.4]
  assign buffer_10_740 = $signed(_T_88534); // @[Modules.scala 63:156:@40728.4]
  assign _T_88536 = $signed(buffer_10_740) + $signed(buffer_10_692); // @[Modules.scala 63:156:@40730.4]
  assign _T_88537 = _T_88536[10:0]; // @[Modules.scala 63:156:@40731.4]
  assign buffer_10_741 = $signed(_T_88537); // @[Modules.scala 63:156:@40732.4]
  assign _T_88539 = $signed(buffer_10_741) + $signed(buffer_10_693); // @[Modules.scala 63:156:@40734.4]
  assign _T_88540 = _T_88539[10:0]; // @[Modules.scala 63:156:@40735.4]
  assign buffer_10_742 = $signed(_T_88540); // @[Modules.scala 63:156:@40736.4]
  assign _T_88542 = $signed(buffer_10_742) + $signed(buffer_10_694); // @[Modules.scala 63:156:@40738.4]
  assign _T_88543 = _T_88542[10:0]; // @[Modules.scala 63:156:@40739.4]
  assign buffer_10_743 = $signed(_T_88543); // @[Modules.scala 63:156:@40740.4]
  assign _T_88545 = $signed(buffer_10_743) + $signed(buffer_10_695); // @[Modules.scala 63:156:@40742.4]
  assign _T_88546 = _T_88545[10:0]; // @[Modules.scala 63:156:@40743.4]
  assign buffer_10_744 = $signed(_T_88546); // @[Modules.scala 63:156:@40744.4]
  assign _T_88548 = $signed(buffer_10_744) + $signed(buffer_10_696); // @[Modules.scala 63:156:@40746.4]
  assign _T_88549 = _T_88548[10:0]; // @[Modules.scala 63:156:@40747.4]
  assign buffer_10_745 = $signed(_T_88549); // @[Modules.scala 63:156:@40748.4]
  assign _T_88551 = $signed(buffer_10_745) + $signed(buffer_10_697); // @[Modules.scala 63:156:@40750.4]
  assign _T_88552 = _T_88551[10:0]; // @[Modules.scala 63:156:@40751.4]
  assign buffer_10_746 = $signed(_T_88552); // @[Modules.scala 63:156:@40752.4]
  assign _T_88554 = $signed(buffer_10_746) + $signed(buffer_10_698); // @[Modules.scala 63:156:@40754.4]
  assign _T_88555 = _T_88554[10:0]; // @[Modules.scala 63:156:@40755.4]
  assign buffer_10_747 = $signed(_T_88555); // @[Modules.scala 63:156:@40756.4]
  assign _T_88557 = $signed(buffer_10_747) + $signed(buffer_10_699); // @[Modules.scala 63:156:@40758.4]
  assign _T_88558 = _T_88557[10:0]; // @[Modules.scala 63:156:@40759.4]
  assign buffer_10_748 = $signed(_T_88558); // @[Modules.scala 63:156:@40760.4]
  assign _T_88560 = $signed(buffer_10_748) + $signed(buffer_10_700); // @[Modules.scala 63:156:@40762.4]
  assign _T_88561 = _T_88560[10:0]; // @[Modules.scala 63:156:@40763.4]
  assign buffer_10_749 = $signed(_T_88561); // @[Modules.scala 63:156:@40764.4]
  assign _T_88563 = $signed(buffer_10_749) + $signed(buffer_10_701); // @[Modules.scala 63:156:@40766.4]
  assign _T_88564 = _T_88563[10:0]; // @[Modules.scala 63:156:@40767.4]
  assign buffer_10_750 = $signed(_T_88564); // @[Modules.scala 63:156:@40768.4]
  assign _T_88566 = $signed(buffer_10_750) + $signed(buffer_10_702); // @[Modules.scala 63:156:@40770.4]
  assign _T_88567 = _T_88566[10:0]; // @[Modules.scala 63:156:@40771.4]
  assign buffer_10_751 = $signed(_T_88567); // @[Modules.scala 63:156:@40772.4]
  assign _T_88569 = $signed(buffer_10_751) + $signed(buffer_10_703); // @[Modules.scala 63:156:@40774.4]
  assign _T_88570 = _T_88569[10:0]; // @[Modules.scala 63:156:@40775.4]
  assign buffer_10_752 = $signed(_T_88570); // @[Modules.scala 63:156:@40776.4]
  assign _T_88572 = $signed(buffer_10_752) + $signed(buffer_10_704); // @[Modules.scala 63:156:@40778.4]
  assign _T_88573 = _T_88572[10:0]; // @[Modules.scala 63:156:@40779.4]
  assign buffer_10_753 = $signed(_T_88573); // @[Modules.scala 63:156:@40780.4]
  assign _T_88575 = $signed(buffer_10_753) + $signed(buffer_10_705); // @[Modules.scala 63:156:@40782.4]
  assign _T_88576 = _T_88575[10:0]; // @[Modules.scala 63:156:@40783.4]
  assign buffer_10_754 = $signed(_T_88576); // @[Modules.scala 63:156:@40784.4]
  assign _T_88578 = $signed(buffer_10_754) + $signed(buffer_10_706); // @[Modules.scala 63:156:@40786.4]
  assign _T_88579 = _T_88578[10:0]; // @[Modules.scala 63:156:@40787.4]
  assign buffer_10_755 = $signed(_T_88579); // @[Modules.scala 63:156:@40788.4]
  assign _T_88581 = $signed(buffer_10_755) + $signed(buffer_9_707); // @[Modules.scala 63:156:@40790.4]
  assign _T_88582 = _T_88581[10:0]; // @[Modules.scala 63:156:@40791.4]
  assign buffer_10_756 = $signed(_T_88582); // @[Modules.scala 63:156:@40792.4]
  assign _T_88584 = $signed(buffer_10_756) + $signed(buffer_10_708); // @[Modules.scala 63:156:@40794.4]
  assign _T_88585 = _T_88584[10:0]; // @[Modules.scala 63:156:@40795.4]
  assign buffer_10_757 = $signed(_T_88585); // @[Modules.scala 63:156:@40796.4]
  assign _T_88587 = $signed(buffer_10_757) + $signed(buffer_10_709); // @[Modules.scala 63:156:@40798.4]
  assign _T_88588 = _T_88587[10:0]; // @[Modules.scala 63:156:@40799.4]
  assign buffer_10_758 = $signed(_T_88588); // @[Modules.scala 63:156:@40800.4]
  assign _T_88590 = $signed(buffer_10_758) + $signed(buffer_10_710); // @[Modules.scala 63:156:@40802.4]
  assign _T_88591 = _T_88590[10:0]; // @[Modules.scala 63:156:@40803.4]
  assign buffer_10_759 = $signed(_T_88591); // @[Modules.scala 63:156:@40804.4]
  assign _T_88593 = $signed(buffer_10_759) + $signed(buffer_10_711); // @[Modules.scala 63:156:@40806.4]
  assign _T_88594 = _T_88593[10:0]; // @[Modules.scala 63:156:@40807.4]
  assign buffer_10_760 = $signed(_T_88594); // @[Modules.scala 63:156:@40808.4]
  assign _T_88596 = $signed(buffer_10_760) + $signed(buffer_10_712); // @[Modules.scala 63:156:@40810.4]
  assign _T_88597 = _T_88596[10:0]; // @[Modules.scala 63:156:@40811.4]
  assign buffer_10_761 = $signed(_T_88597); // @[Modules.scala 63:156:@40812.4]
  assign _T_88599 = $signed(buffer_10_761) + $signed(buffer_10_713); // @[Modules.scala 63:156:@40814.4]
  assign _T_88600 = _T_88599[10:0]; // @[Modules.scala 63:156:@40815.4]
  assign buffer_10_762 = $signed(_T_88600); // @[Modules.scala 63:156:@40816.4]
  assign _T_88602 = $signed(buffer_10_762) + $signed(buffer_10_714); // @[Modules.scala 63:156:@40818.4]
  assign _T_88603 = _T_88602[10:0]; // @[Modules.scala 63:156:@40819.4]
  assign buffer_10_763 = $signed(_T_88603); // @[Modules.scala 63:156:@40820.4]
  assign _T_88605 = $signed(buffer_10_763) + $signed(buffer_10_715); // @[Modules.scala 63:156:@40822.4]
  assign _T_88606 = _T_88605[10:0]; // @[Modules.scala 63:156:@40823.4]
  assign buffer_10_764 = $signed(_T_88606); // @[Modules.scala 63:156:@40824.4]
  assign _T_88608 = $signed(buffer_10_764) + $signed(buffer_10_716); // @[Modules.scala 63:156:@40826.4]
  assign _T_88609 = _T_88608[10:0]; // @[Modules.scala 63:156:@40827.4]
  assign buffer_10_765 = $signed(_T_88609); // @[Modules.scala 63:156:@40828.4]
  assign _T_88611 = $signed(buffer_10_765) + $signed(buffer_10_717); // @[Modules.scala 63:156:@40830.4]
  assign _T_88612 = _T_88611[10:0]; // @[Modules.scala 63:156:@40831.4]
  assign buffer_10_766 = $signed(_T_88612); // @[Modules.scala 63:156:@40832.4]
  assign _T_88614 = $signed(buffer_10_766) + $signed(buffer_10_718); // @[Modules.scala 63:156:@40834.4]
  assign _T_88615 = _T_88614[10:0]; // @[Modules.scala 63:156:@40835.4]
  assign buffer_10_767 = $signed(_T_88615); // @[Modules.scala 63:156:@40836.4]
  assign _T_88617 = $signed(buffer_10_767) + $signed(buffer_10_719); // @[Modules.scala 63:156:@40838.4]
  assign _T_88618 = _T_88617[10:0]; // @[Modules.scala 63:156:@40839.4]
  assign buffer_10_768 = $signed(_T_88618); // @[Modules.scala 63:156:@40840.4]
  assign _T_88620 = $signed(buffer_10_768) + $signed(buffer_10_720); // @[Modules.scala 63:156:@40842.4]
  assign _T_88621 = _T_88620[10:0]; // @[Modules.scala 63:156:@40843.4]
  assign buffer_10_769 = $signed(_T_88621); // @[Modules.scala 63:156:@40844.4]
  assign _T_88623 = $signed(buffer_10_769) + $signed(buffer_10_721); // @[Modules.scala 63:156:@40846.4]
  assign _T_88624 = _T_88623[10:0]; // @[Modules.scala 63:156:@40847.4]
  assign buffer_10_770 = $signed(_T_88624); // @[Modules.scala 63:156:@40848.4]
  assign _T_88626 = $signed(buffer_10_770) + $signed(buffer_10_722); // @[Modules.scala 63:156:@40850.4]
  assign _T_88627 = _T_88626[10:0]; // @[Modules.scala 63:156:@40851.4]
  assign buffer_10_771 = $signed(_T_88627); // @[Modules.scala 63:156:@40852.4]
  assign _T_88629 = $signed(buffer_10_771) + $signed(buffer_10_723); // @[Modules.scala 63:156:@40854.4]
  assign _T_88630 = _T_88629[10:0]; // @[Modules.scala 63:156:@40855.4]
  assign buffer_10_772 = $signed(_T_88630); // @[Modules.scala 63:156:@40856.4]
  assign _T_88632 = $signed(buffer_10_772) + $signed(buffer_10_724); // @[Modules.scala 63:156:@40858.4]
  assign _T_88633 = _T_88632[10:0]; // @[Modules.scala 63:156:@40859.4]
  assign buffer_10_773 = $signed(_T_88633); // @[Modules.scala 63:156:@40860.4]
  assign _T_88635 = $signed(buffer_10_773) + $signed(buffer_10_725); // @[Modules.scala 63:156:@40862.4]
  assign _T_88636 = _T_88635[10:0]; // @[Modules.scala 63:156:@40863.4]
  assign buffer_10_774 = $signed(_T_88636); // @[Modules.scala 63:156:@40864.4]
  assign _T_88638 = $signed(buffer_10_774) + $signed(buffer_10_726); // @[Modules.scala 63:156:@40866.4]
  assign _T_88639 = _T_88638[10:0]; // @[Modules.scala 63:156:@40867.4]
  assign buffer_10_775 = $signed(_T_88639); // @[Modules.scala 63:156:@40868.4]
  assign _T_88641 = $signed(buffer_10_775) + $signed(buffer_10_727); // @[Modules.scala 63:156:@40870.4]
  assign _T_88642 = _T_88641[10:0]; // @[Modules.scala 63:156:@40871.4]
  assign buffer_10_776 = $signed(_T_88642); // @[Modules.scala 63:156:@40872.4]
  assign _T_88644 = $signed(buffer_10_776) + $signed(buffer_10_728); // @[Modules.scala 63:156:@40874.4]
  assign _T_88645 = _T_88644[10:0]; // @[Modules.scala 63:156:@40875.4]
  assign buffer_10_777 = $signed(_T_88645); // @[Modules.scala 63:156:@40876.4]
  assign _T_88647 = $signed(buffer_10_777) + $signed(buffer_10_729); // @[Modules.scala 63:156:@40878.4]
  assign _T_88648 = _T_88647[10:0]; // @[Modules.scala 63:156:@40879.4]
  assign buffer_10_778 = $signed(_T_88648); // @[Modules.scala 63:156:@40880.4]
  assign _T_88650 = $signed(buffer_10_778) + $signed(buffer_10_730); // @[Modules.scala 63:156:@40882.4]
  assign _T_88651 = _T_88650[10:0]; // @[Modules.scala 63:156:@40883.4]
  assign buffer_10_779 = $signed(_T_88651); // @[Modules.scala 63:156:@40884.4]
  assign _T_88653 = $signed(buffer_10_779) + $signed(buffer_10_731); // @[Modules.scala 63:156:@40886.4]
  assign _T_88654 = _T_88653[10:0]; // @[Modules.scala 63:156:@40887.4]
  assign buffer_10_780 = $signed(_T_88654); // @[Modules.scala 63:156:@40888.4]
  assign _T_88656 = $signed(buffer_10_780) + $signed(buffer_10_732); // @[Modules.scala 63:156:@40890.4]
  assign _T_88657 = _T_88656[10:0]; // @[Modules.scala 63:156:@40891.4]
  assign buffer_10_781 = $signed(_T_88657); // @[Modules.scala 63:156:@40892.4]
  assign _T_88659 = $signed(buffer_10_781) + $signed(buffer_10_733); // @[Modules.scala 63:156:@40894.4]
  assign _T_88660 = _T_88659[10:0]; // @[Modules.scala 63:156:@40895.4]
  assign buffer_10_782 = $signed(_T_88660); // @[Modules.scala 63:156:@40896.4]
  assign _T_88662 = $signed(buffer_10_782) + $signed(buffer_10_734); // @[Modules.scala 63:156:@40898.4]
  assign _T_88663 = _T_88662[10:0]; // @[Modules.scala 63:156:@40899.4]
  assign buffer_10_783 = $signed(_T_88663); // @[Modules.scala 63:156:@40900.4]
  assign _T_88750 = $signed(_T_54386) + $signed(io_in_39); // @[Modules.scala 43:47:@41000.4]
  assign _T_88751 = _T_88750[4:0]; // @[Modules.scala 43:47:@41001.4]
  assign _T_88752 = $signed(_T_88751); // @[Modules.scala 43:47:@41002.4]
  assign _T_88759 = $signed(io_in_44) - $signed(io_in_45); // @[Modules.scala 40:46:@41012.4]
  assign _T_88760 = _T_88759[4:0]; // @[Modules.scala 40:46:@41013.4]
  assign _T_88761 = $signed(_T_88760); // @[Modules.scala 40:46:@41014.4]
  assign _T_88766 = $signed(_T_54414) + $signed(io_in_47); // @[Modules.scala 43:47:@41019.4]
  assign _T_88767 = _T_88766[4:0]; // @[Modules.scala 43:47:@41020.4]
  assign _T_88768 = $signed(_T_88767); // @[Modules.scala 43:47:@41021.4]
  assign _T_88878 = $signed(io_in_86) + $signed(io_in_87); // @[Modules.scala 37:46:@41138.4]
  assign _T_88879 = _T_88878[4:0]; // @[Modules.scala 37:46:@41139.4]
  assign _T_88880 = $signed(_T_88879); // @[Modules.scala 37:46:@41140.4]
  assign _T_89147 = $signed(_T_54767) + $signed(io_in_181); // @[Modules.scala 43:47:@41422.4]
  assign _T_89148 = _T_89147[4:0]; // @[Modules.scala 43:47:@41423.4]
  assign _T_89149 = $signed(_T_89148); // @[Modules.scala 43:47:@41424.4]
  assign _T_89220 = $signed(_T_67364) + $signed(io_in_211); // @[Modules.scala 43:47:@41503.4]
  assign _T_89221 = _T_89220[4:0]; // @[Modules.scala 43:47:@41504.4]
  assign _T_89222 = $signed(_T_89221); // @[Modules.scala 43:47:@41505.4]
  assign _T_89245 = $signed(io_in_224) - $signed(io_in_225); // @[Modules.scala 40:46:@41534.4]
  assign _T_89246 = _T_89245[4:0]; // @[Modules.scala 40:46:@41535.4]
  assign _T_89247 = $signed(_T_89246); // @[Modules.scala 40:46:@41536.4]
  assign _T_89286 = $signed(_T_54946) + $signed(io_in_239); // @[Modules.scala 43:47:@41577.4]
  assign _T_89287 = _T_89286[4:0]; // @[Modules.scala 43:47:@41578.4]
  assign _T_89288 = $signed(_T_89287); // @[Modules.scala 43:47:@41579.4]
  assign _T_89366 = $signed(_T_55054) + $signed(io_in_271); // @[Modules.scala 43:47:@41665.4]
  assign _T_89367 = _T_89366[4:0]; // @[Modules.scala 43:47:@41666.4]
  assign _T_89368 = $signed(_T_89367); // @[Modules.scala 43:47:@41667.4]
  assign _T_89604 = $signed(_T_64771) + $signed(io_in_371); // @[Modules.scala 43:47:@41931.4]
  assign _T_89605 = _T_89604[4:0]; // @[Modules.scala 43:47:@41932.4]
  assign _T_89606 = $signed(_T_89605); // @[Modules.scala 43:47:@41933.4]
  assign _T_89611 = $signed(_T_64778) + $signed(io_in_373); // @[Modules.scala 43:47:@41938.4]
  assign _T_89612 = _T_89611[4:0]; // @[Modules.scala 43:47:@41939.4]
  assign _T_89613 = $signed(_T_89612); // @[Modules.scala 43:47:@41940.4]
  assign _T_89767 = $signed(_T_70960) + $signed(io_in_429); // @[Modules.scala 43:47:@42104.4]
  assign _T_89768 = _T_89767[4:0]; // @[Modules.scala 43:47:@42105.4]
  assign _T_89769 = $signed(_T_89768); // @[Modules.scala 43:47:@42106.4]
  assign _T_89780 = $signed(io_in_434) - $signed(io_in_435); // @[Modules.scala 40:46:@42119.4]
  assign _T_89781 = _T_89780[4:0]; // @[Modules.scala 40:46:@42120.4]
  assign _T_89782 = $signed(_T_89781); // @[Modules.scala 40:46:@42121.4]
  assign _T_89832 = $signed(io_in_450) - $signed(io_in_451); // @[Modules.scala 40:46:@42172.4]
  assign _T_89833 = _T_89832[4:0]; // @[Modules.scala 40:46:@42173.4]
  assign _T_89834 = $signed(_T_89833); // @[Modules.scala 40:46:@42174.4]
  assign _T_89894 = $signed(_T_55550) + $signed(io_in_471); // @[Modules.scala 43:47:@42236.4]
  assign _T_89895 = _T_89894[4:0]; // @[Modules.scala 43:47:@42237.4]
  assign _T_89896 = $signed(_T_89895); // @[Modules.scala 43:47:@42238.4]
  assign _T_89929 = $signed(_T_55581) + $signed(io_in_481); // @[Modules.scala 43:47:@42271.4]
  assign _T_89930 = _T_89929[4:0]; // @[Modules.scala 43:47:@42272.4]
  assign _T_89931 = $signed(_T_89930); // @[Modules.scala 43:47:@42273.4]
  assign _T_89980 = $signed(_T_61942) + $signed(io_in_499); // @[Modules.scala 43:47:@42325.4]
  assign _T_89981 = _T_89980[4:0]; // @[Modules.scala 43:47:@42326.4]
  assign _T_89982 = $signed(_T_89981); // @[Modules.scala 43:47:@42327.4]
  assign _T_90031 = $signed(_T_58840) + $signed(io_in_517); // @[Modules.scala 43:47:@42379.4]
  assign _T_90032 = _T_90031[4:0]; // @[Modules.scala 43:47:@42380.4]
  assign _T_90033 = $signed(_T_90032); // @[Modules.scala 43:47:@42381.4]
  assign _T_90168 = $signed(io_in_562) - $signed(io_in_563); // @[Modules.scala 40:46:@42522.4]
  assign _T_90169 = _T_90168[4:0]; // @[Modules.scala 40:46:@42523.4]
  assign _T_90170 = $signed(_T_90169); // @[Modules.scala 40:46:@42524.4]
  assign _T_90323 = $signed(_T_55963) + $signed(io_in_621); // @[Modules.scala 43:47:@42689.4]
  assign _T_90324 = _T_90323[4:0]; // @[Modules.scala 43:47:@42690.4]
  assign _T_90325 = $signed(_T_90324); // @[Modules.scala 43:47:@42691.4]
  assign _T_90592 = $signed(_T_65599) + $signed(io_in_723); // @[Modules.scala 43:47:@42980.4]
  assign _T_90593 = _T_90592[4:0]; // @[Modules.scala 43:47:@42981.4]
  assign _T_90594 = $signed(_T_90593); // @[Modules.scala 43:47:@42982.4]
  assign _T_90793 = $signed(buffer_0_8) + $signed(buffer_1_9); // @[Modules.scala 50:57:@43192.4]
  assign _T_90794 = _T_90793[10:0]; // @[Modules.scala 50:57:@43193.4]
  assign buffer_11_396 = $signed(_T_90794); // @[Modules.scala 50:57:@43194.4]
  assign _T_90796 = $signed(buffer_7_10) + $signed(buffer_4_11); // @[Modules.scala 50:57:@43196.4]
  assign _T_90797 = _T_90796[10:0]; // @[Modules.scala 50:57:@43197.4]
  assign buffer_11_397 = $signed(_T_90797); // @[Modules.scala 50:57:@43198.4]
  assign _T_90802 = $signed(buffer_3_14) + $signed(buffer_1_15); // @[Modules.scala 50:57:@43204.4]
  assign _T_90803 = _T_90802[10:0]; // @[Modules.scala 50:57:@43205.4]
  assign buffer_11_399 = $signed(_T_90803); // @[Modules.scala 50:57:@43206.4]
  assign buffer_11_19 = {{6{_T_88752[4]}},_T_88752}; // @[Modules.scala 32:22:@8.4]
  assign _T_90808 = $signed(buffer_0_18) + $signed(buffer_11_19); // @[Modules.scala 50:57:@43212.4]
  assign _T_90809 = _T_90808[10:0]; // @[Modules.scala 50:57:@43213.4]
  assign buffer_11_401 = $signed(_T_90809); // @[Modules.scala 50:57:@43214.4]
  assign buffer_11_22 = {{6{_T_88761[4]}},_T_88761}; // @[Modules.scala 32:22:@8.4]
  assign buffer_11_23 = {{6{_T_88768[4]}},_T_88768}; // @[Modules.scala 32:22:@8.4]
  assign _T_90814 = $signed(buffer_11_22) + $signed(buffer_11_23); // @[Modules.scala 50:57:@43220.4]
  assign _T_90815 = _T_90814[10:0]; // @[Modules.scala 50:57:@43221.4]
  assign buffer_11_403 = $signed(_T_90815); // @[Modules.scala 50:57:@43222.4]
  assign _T_90820 = $signed(buffer_3_26) + $signed(buffer_1_27); // @[Modules.scala 50:57:@43228.4]
  assign _T_90821 = _T_90820[10:0]; // @[Modules.scala 50:57:@43229.4]
  assign buffer_11_405 = $signed(_T_90821); // @[Modules.scala 50:57:@43230.4]
  assign _T_90823 = $signed(buffer_3_28) + $signed(buffer_2_29); // @[Modules.scala 50:57:@43232.4]
  assign _T_90824 = _T_90823[10:0]; // @[Modules.scala 50:57:@43233.4]
  assign buffer_11_406 = $signed(_T_90824); // @[Modules.scala 50:57:@43234.4]
  assign _T_90832 = $signed(buffer_0_34) + $signed(buffer_1_35); // @[Modules.scala 50:57:@43244.4]
  assign _T_90833 = _T_90832[10:0]; // @[Modules.scala 50:57:@43245.4]
  assign buffer_11_409 = $signed(_T_90833); // @[Modules.scala 50:57:@43246.4]
  assign buffer_11_43 = {{6{_T_88880[4]}},_T_88880}; // @[Modules.scala 32:22:@8.4]
  assign _T_90844 = $signed(buffer_2_42) + $signed(buffer_11_43); // @[Modules.scala 50:57:@43260.4]
  assign _T_90845 = _T_90844[10:0]; // @[Modules.scala 50:57:@43261.4]
  assign buffer_11_413 = $signed(_T_90845); // @[Modules.scala 50:57:@43262.4]
  assign _T_90847 = $signed(buffer_2_44) + $signed(buffer_3_45); // @[Modules.scala 50:57:@43264.4]
  assign _T_90848 = _T_90847[10:0]; // @[Modules.scala 50:57:@43265.4]
  assign buffer_11_414 = $signed(_T_90848); // @[Modules.scala 50:57:@43266.4]
  assign _T_90883 = $signed(buffer_0_68) + $signed(buffer_3_69); // @[Modules.scala 50:57:@43312.4]
  assign _T_90884 = _T_90883[10:0]; // @[Modules.scala 50:57:@43313.4]
  assign buffer_11_426 = $signed(_T_90884); // @[Modules.scala 50:57:@43314.4]
  assign _T_90886 = $signed(buffer_0_70) + $signed(buffer_2_71); // @[Modules.scala 50:57:@43316.4]
  assign _T_90887 = _T_90886[10:0]; // @[Modules.scala 50:57:@43317.4]
  assign buffer_11_427 = $signed(_T_90887); // @[Modules.scala 50:57:@43318.4]
  assign _T_90904 = $signed(buffer_5_82) + $signed(buffer_1_83); // @[Modules.scala 50:57:@43340.4]
  assign _T_90905 = _T_90904[10:0]; // @[Modules.scala 50:57:@43341.4]
  assign buffer_11_433 = $signed(_T_90905); // @[Modules.scala 50:57:@43342.4]
  assign buffer_11_90 = {{6{_T_89149[4]}},_T_89149}; // @[Modules.scala 32:22:@8.4]
  assign _T_90916 = $signed(buffer_11_90) + $signed(buffer_1_91); // @[Modules.scala 50:57:@43356.4]
  assign _T_90917 = _T_90916[10:0]; // @[Modules.scala 50:57:@43357.4]
  assign buffer_11_437 = $signed(_T_90917); // @[Modules.scala 50:57:@43358.4]
  assign _T_90919 = $signed(buffer_3_92) + $signed(buffer_0_93); // @[Modules.scala 50:57:@43360.4]
  assign _T_90920 = _T_90919[10:0]; // @[Modules.scala 50:57:@43361.4]
  assign buffer_11_438 = $signed(_T_90920); // @[Modules.scala 50:57:@43362.4]
  assign _T_90922 = $signed(buffer_1_94) + $signed(buffer_2_95); // @[Modules.scala 50:57:@43364.4]
  assign _T_90923 = _T_90922[10:0]; // @[Modules.scala 50:57:@43365.4]
  assign buffer_11_439 = $signed(_T_90923); // @[Modules.scala 50:57:@43366.4]
  assign _T_90928 = $signed(buffer_6_98) + $signed(buffer_2_99); // @[Modules.scala 50:57:@43372.4]
  assign _T_90929 = _T_90928[10:0]; // @[Modules.scala 50:57:@43373.4]
  assign buffer_11_441 = $signed(_T_90929); // @[Modules.scala 50:57:@43374.4]
  assign buffer_11_105 = {{6{_T_89222[4]}},_T_89222}; // @[Modules.scala 32:22:@8.4]
  assign _T_90937 = $signed(buffer_0_104) + $signed(buffer_11_105); // @[Modules.scala 50:57:@43384.4]
  assign _T_90938 = _T_90937[10:0]; // @[Modules.scala 50:57:@43385.4]
  assign buffer_11_444 = $signed(_T_90938); // @[Modules.scala 50:57:@43386.4]
  assign _T_90940 = $signed(buffer_4_106) + $signed(buffer_6_107); // @[Modules.scala 50:57:@43388.4]
  assign _T_90941 = _T_90940[10:0]; // @[Modules.scala 50:57:@43389.4]
  assign buffer_11_445 = $signed(_T_90941); // @[Modules.scala 50:57:@43390.4]
  assign buffer_11_112 = {{6{_T_89247[4]}},_T_89247}; // @[Modules.scala 32:22:@8.4]
  assign _T_90949 = $signed(buffer_11_112) + $signed(buffer_0_113); // @[Modules.scala 50:57:@43400.4]
  assign _T_90950 = _T_90949[10:0]; // @[Modules.scala 50:57:@43401.4]
  assign buffer_11_448 = $signed(_T_90950); // @[Modules.scala 50:57:@43402.4]
  assign _T_90955 = $signed(buffer_0_116) + $signed(buffer_7_117); // @[Modules.scala 50:57:@43408.4]
  assign _T_90956 = _T_90955[10:0]; // @[Modules.scala 50:57:@43409.4]
  assign buffer_11_450 = $signed(_T_90956); // @[Modules.scala 50:57:@43410.4]
  assign buffer_11_119 = {{6{_T_89288[4]}},_T_89288}; // @[Modules.scala 32:22:@8.4]
  assign _T_90958 = $signed(buffer_3_118) + $signed(buffer_11_119); // @[Modules.scala 50:57:@43412.4]
  assign _T_90959 = _T_90958[10:0]; // @[Modules.scala 50:57:@43413.4]
  assign buffer_11_451 = $signed(_T_90959); // @[Modules.scala 50:57:@43414.4]
  assign _T_90961 = $signed(buffer_6_120) + $signed(buffer_4_121); // @[Modules.scala 50:57:@43416.4]
  assign _T_90962 = _T_90961[10:0]; // @[Modules.scala 50:57:@43417.4]
  assign buffer_11_452 = $signed(_T_90962); // @[Modules.scala 50:57:@43418.4]
  assign _T_90964 = $signed(buffer_9_122) + $signed(buffer_3_123); // @[Modules.scala 50:57:@43420.4]
  assign _T_90965 = _T_90964[10:0]; // @[Modules.scala 50:57:@43421.4]
  assign buffer_11_453 = $signed(_T_90965); // @[Modules.scala 50:57:@43422.4]
  assign _T_90973 = $signed(buffer_0_128) + $signed(buffer_4_129); // @[Modules.scala 50:57:@43432.4]
  assign _T_90974 = _T_90973[10:0]; // @[Modules.scala 50:57:@43433.4]
  assign buffer_11_456 = $signed(_T_90974); // @[Modules.scala 50:57:@43434.4]
  assign _T_90979 = $signed(buffer_5_132) + $signed(buffer_0_133); // @[Modules.scala 50:57:@43440.4]
  assign _T_90980 = _T_90979[10:0]; // @[Modules.scala 50:57:@43441.4]
  assign buffer_11_458 = $signed(_T_90980); // @[Modules.scala 50:57:@43442.4]
  assign buffer_11_135 = {{6{_T_89368[4]}},_T_89368}; // @[Modules.scala 32:22:@8.4]
  assign _T_90982 = $signed(buffer_0_134) + $signed(buffer_11_135); // @[Modules.scala 50:57:@43444.4]
  assign _T_90983 = _T_90982[10:0]; // @[Modules.scala 50:57:@43445.4]
  assign buffer_11_459 = $signed(_T_90983); // @[Modules.scala 50:57:@43446.4]
  assign _T_90991 = $signed(buffer_3_140) + $signed(buffer_0_141); // @[Modules.scala 50:57:@43456.4]
  assign _T_90992 = _T_90991[10:0]; // @[Modules.scala 50:57:@43457.4]
  assign buffer_11_462 = $signed(_T_90992); // @[Modules.scala 50:57:@43458.4]
  assign _T_90994 = $signed(buffer_0_142) + $signed(buffer_7_143); // @[Modules.scala 50:57:@43460.4]
  assign _T_90995 = _T_90994[10:0]; // @[Modules.scala 50:57:@43461.4]
  assign buffer_11_463 = $signed(_T_90995); // @[Modules.scala 50:57:@43462.4]
  assign _T_91015 = $signed(buffer_6_156) + $signed(buffer_2_157); // @[Modules.scala 50:57:@43488.4]
  assign _T_91016 = _T_91015[10:0]; // @[Modules.scala 50:57:@43489.4]
  assign buffer_11_470 = $signed(_T_91016); // @[Modules.scala 50:57:@43490.4]
  assign _T_91021 = $signed(buffer_1_160) + $signed(buffer_5_161); // @[Modules.scala 50:57:@43496.4]
  assign _T_91022 = _T_91021[10:0]; // @[Modules.scala 50:57:@43497.4]
  assign buffer_11_472 = $signed(_T_91022); // @[Modules.scala 50:57:@43498.4]
  assign _T_91051 = $signed(buffer_1_180) + $signed(buffer_8_181); // @[Modules.scala 50:57:@43536.4]
  assign _T_91052 = _T_91051[10:0]; // @[Modules.scala 50:57:@43537.4]
  assign buffer_11_482 = $signed(_T_91052); // @[Modules.scala 50:57:@43538.4]
  assign buffer_11_185 = {{6{_T_89606[4]}},_T_89606}; // @[Modules.scala 32:22:@8.4]
  assign _T_91057 = $signed(buffer_3_184) + $signed(buffer_11_185); // @[Modules.scala 50:57:@43544.4]
  assign _T_91058 = _T_91057[10:0]; // @[Modules.scala 50:57:@43545.4]
  assign buffer_11_484 = $signed(_T_91058); // @[Modules.scala 50:57:@43546.4]
  assign buffer_11_186 = {{6{_T_89613[4]}},_T_89613}; // @[Modules.scala 32:22:@8.4]
  assign _T_91060 = $signed(buffer_11_186) + $signed(buffer_5_187); // @[Modules.scala 50:57:@43548.4]
  assign _T_91061 = _T_91060[10:0]; // @[Modules.scala 50:57:@43549.4]
  assign buffer_11_485 = $signed(_T_91061); // @[Modules.scala 50:57:@43550.4]
  assign _T_91072 = $signed(buffer_5_194) + $signed(buffer_4_195); // @[Modules.scala 50:57:@43564.4]
  assign _T_91073 = _T_91072[10:0]; // @[Modules.scala 50:57:@43565.4]
  assign buffer_11_489 = $signed(_T_91073); // @[Modules.scala 50:57:@43566.4]
  assign _T_91081 = $signed(buffer_5_200) + $signed(buffer_3_201); // @[Modules.scala 50:57:@43576.4]
  assign _T_91082 = _T_91081[10:0]; // @[Modules.scala 50:57:@43577.4]
  assign buffer_11_492 = $signed(_T_91082); // @[Modules.scala 50:57:@43578.4]
  assign _T_91087 = $signed(buffer_3_204) + $signed(buffer_1_205); // @[Modules.scala 50:57:@43584.4]
  assign _T_91088 = _T_91087[10:0]; // @[Modules.scala 50:57:@43585.4]
  assign buffer_11_494 = $signed(_T_91088); // @[Modules.scala 50:57:@43586.4]
  assign _T_91096 = $signed(buffer_3_210) + $signed(buffer_1_211); // @[Modules.scala 50:57:@43596.4]
  assign _T_91097 = _T_91096[10:0]; // @[Modules.scala 50:57:@43597.4]
  assign buffer_11_497 = $signed(_T_91097); // @[Modules.scala 50:57:@43598.4]
  assign buffer_11_214 = {{6{_T_89769[4]}},_T_89769}; // @[Modules.scala 32:22:@8.4]
  assign _T_91102 = $signed(buffer_11_214) + $signed(buffer_2_215); // @[Modules.scala 50:57:@43604.4]
  assign _T_91103 = _T_91102[10:0]; // @[Modules.scala 50:57:@43605.4]
  assign buffer_11_499 = $signed(_T_91103); // @[Modules.scala 50:57:@43606.4]
  assign buffer_11_217 = {{6{_T_89782[4]}},_T_89782}; // @[Modules.scala 32:22:@8.4]
  assign _T_91105 = $signed(buffer_0_216) + $signed(buffer_11_217); // @[Modules.scala 50:57:@43608.4]
  assign _T_91106 = _T_91105[10:0]; // @[Modules.scala 50:57:@43609.4]
  assign buffer_11_500 = $signed(_T_91106); // @[Modules.scala 50:57:@43610.4]
  assign buffer_11_225 = {{6{_T_89834[4]}},_T_89834}; // @[Modules.scala 32:22:@8.4]
  assign _T_91117 = $signed(buffer_1_224) + $signed(buffer_11_225); // @[Modules.scala 50:57:@43624.4]
  assign _T_91118 = _T_91117[10:0]; // @[Modules.scala 50:57:@43625.4]
  assign buffer_11_504 = $signed(_T_91118); // @[Modules.scala 50:57:@43626.4]
  assign _T_91123 = $signed(buffer_1_228) + $signed(buffer_2_229); // @[Modules.scala 50:57:@43632.4]
  assign _T_91124 = _T_91123[10:0]; // @[Modules.scala 50:57:@43633.4]
  assign buffer_11_506 = $signed(_T_91124); // @[Modules.scala 50:57:@43634.4]
  assign buffer_11_235 = {{6{_T_89896[4]}},_T_89896}; // @[Modules.scala 32:22:@8.4]
  assign _T_91132 = $signed(buffer_2_234) + $signed(buffer_11_235); // @[Modules.scala 50:57:@43644.4]
  assign _T_91133 = _T_91132[10:0]; // @[Modules.scala 50:57:@43645.4]
  assign buffer_11_509 = $signed(_T_91133); // @[Modules.scala 50:57:@43646.4]
  assign _T_91138 = $signed(buffer_1_238) + $signed(buffer_7_239); // @[Modules.scala 50:57:@43652.4]
  assign _T_91139 = _T_91138[10:0]; // @[Modules.scala 50:57:@43653.4]
  assign buffer_11_511 = $signed(_T_91139); // @[Modules.scala 50:57:@43654.4]
  assign buffer_11_240 = {{6{_T_89931[4]}},_T_89931}; // @[Modules.scala 32:22:@8.4]
  assign _T_91141 = $signed(buffer_11_240) + $signed(buffer_3_241); // @[Modules.scala 50:57:@43656.4]
  assign _T_91142 = _T_91141[10:0]; // @[Modules.scala 50:57:@43657.4]
  assign buffer_11_512 = $signed(_T_91142); // @[Modules.scala 50:57:@43658.4]
  assign buffer_11_249 = {{6{_T_89982[4]}},_T_89982}; // @[Modules.scala 32:22:@8.4]
  assign _T_91153 = $signed(buffer_0_248) + $signed(buffer_11_249); // @[Modules.scala 50:57:@43672.4]
  assign _T_91154 = _T_91153[10:0]; // @[Modules.scala 50:57:@43673.4]
  assign buffer_11_516 = $signed(_T_91154); // @[Modules.scala 50:57:@43674.4]
  assign _T_91165 = $signed(buffer_0_256) + $signed(buffer_4_257); // @[Modules.scala 50:57:@43688.4]
  assign _T_91166 = _T_91165[10:0]; // @[Modules.scala 50:57:@43689.4]
  assign buffer_11_520 = $signed(_T_91166); // @[Modules.scala 50:57:@43690.4]
  assign buffer_11_258 = {{6{_T_90033[4]}},_T_90033}; // @[Modules.scala 32:22:@8.4]
  assign _T_91168 = $signed(buffer_11_258) + $signed(buffer_1_259); // @[Modules.scala 50:57:@43692.4]
  assign _T_91169 = _T_91168[10:0]; // @[Modules.scala 50:57:@43693.4]
  assign buffer_11_521 = $signed(_T_91169); // @[Modules.scala 50:57:@43694.4]
  assign _T_91174 = $signed(buffer_7_262) + $signed(buffer_1_263); // @[Modules.scala 50:57:@43700.4]
  assign _T_91175 = _T_91174[10:0]; // @[Modules.scala 50:57:@43701.4]
  assign buffer_11_523 = $signed(_T_91175); // @[Modules.scala 50:57:@43702.4]
  assign _T_91186 = $signed(buffer_1_270) + $signed(buffer_0_271); // @[Modules.scala 50:57:@43716.4]
  assign _T_91187 = _T_91186[10:0]; // @[Modules.scala 50:57:@43717.4]
  assign buffer_11_527 = $signed(_T_91187); // @[Modules.scala 50:57:@43718.4]
  assign _T_91189 = $signed(buffer_1_272) + $signed(buffer_0_273); // @[Modules.scala 50:57:@43720.4]
  assign _T_91190 = _T_91189[10:0]; // @[Modules.scala 50:57:@43721.4]
  assign buffer_11_528 = $signed(_T_91190); // @[Modules.scala 50:57:@43722.4]
  assign _T_91195 = $signed(buffer_6_276) + $signed(buffer_3_277); // @[Modules.scala 50:57:@43728.4]
  assign _T_91196 = _T_91195[10:0]; // @[Modules.scala 50:57:@43729.4]
  assign buffer_11_530 = $signed(_T_91196); // @[Modules.scala 50:57:@43730.4]
  assign buffer_11_281 = {{6{_T_90170[4]}},_T_90170}; // @[Modules.scala 32:22:@8.4]
  assign _T_91201 = $signed(buffer_0_280) + $signed(buffer_11_281); // @[Modules.scala 50:57:@43736.4]
  assign _T_91202 = _T_91201[10:0]; // @[Modules.scala 50:57:@43737.4]
  assign buffer_11_532 = $signed(_T_91202); // @[Modules.scala 50:57:@43738.4]
  assign _T_91210 = $signed(buffer_3_286) + $signed(buffer_5_287); // @[Modules.scala 50:57:@43748.4]
  assign _T_91211 = _T_91210[10:0]; // @[Modules.scala 50:57:@43749.4]
  assign buffer_11_535 = $signed(_T_91211); // @[Modules.scala 50:57:@43750.4]
  assign _T_91216 = $signed(buffer_2_290) + $signed(buffer_3_291); // @[Modules.scala 50:57:@43756.4]
  assign _T_91217 = _T_91216[10:0]; // @[Modules.scala 50:57:@43757.4]
  assign buffer_11_537 = $signed(_T_91217); // @[Modules.scala 50:57:@43758.4]
  assign _T_91225 = $signed(buffer_0_296) + $signed(buffer_3_297); // @[Modules.scala 50:57:@43768.4]
  assign _T_91226 = _T_91225[10:0]; // @[Modules.scala 50:57:@43769.4]
  assign buffer_11_540 = $signed(_T_91226); // @[Modules.scala 50:57:@43770.4]
  assign _T_91234 = $signed(buffer_0_302) + $signed(buffer_8_303); // @[Modules.scala 50:57:@43780.4]
  assign _T_91235 = _T_91234[10:0]; // @[Modules.scala 50:57:@43781.4]
  assign buffer_11_543 = $signed(_T_91235); // @[Modules.scala 50:57:@43782.4]
  assign _T_91240 = $signed(buffer_1_306) + $signed(buffer_7_307); // @[Modules.scala 50:57:@43788.4]
  assign _T_91241 = _T_91240[10:0]; // @[Modules.scala 50:57:@43789.4]
  assign buffer_11_545 = $signed(_T_91241); // @[Modules.scala 50:57:@43790.4]
  assign buffer_11_310 = {{6{_T_90325[4]}},_T_90325}; // @[Modules.scala 32:22:@8.4]
  assign _T_91246 = $signed(buffer_11_310) + $signed(buffer_7_311); // @[Modules.scala 50:57:@43796.4]
  assign _T_91247 = _T_91246[10:0]; // @[Modules.scala 50:57:@43797.4]
  assign buffer_11_547 = $signed(_T_91247); // @[Modules.scala 50:57:@43798.4]
  assign _T_91249 = $signed(buffer_0_312) + $signed(buffer_3_313); // @[Modules.scala 50:57:@43800.4]
  assign _T_91250 = _T_91249[10:0]; // @[Modules.scala 50:57:@43801.4]
  assign buffer_11_548 = $signed(_T_91250); // @[Modules.scala 50:57:@43802.4]
  assign _T_91261 = $signed(buffer_1_320) + $signed(buffer_3_321); // @[Modules.scala 50:57:@43816.4]
  assign _T_91262 = _T_91261[10:0]; // @[Modules.scala 50:57:@43817.4]
  assign buffer_11_552 = $signed(_T_91262); // @[Modules.scala 50:57:@43818.4]
  assign _T_91270 = $signed(buffer_0_326) + $signed(buffer_8_327); // @[Modules.scala 50:57:@43828.4]
  assign _T_91271 = _T_91270[10:0]; // @[Modules.scala 50:57:@43829.4]
  assign buffer_11_555 = $signed(_T_91271); // @[Modules.scala 50:57:@43830.4]
  assign _T_91285 = $signed(buffer_1_336) + $signed(buffer_6_337); // @[Modules.scala 50:57:@43848.4]
  assign _T_91286 = _T_91285[10:0]; // @[Modules.scala 50:57:@43849.4]
  assign buffer_11_560 = $signed(_T_91286); // @[Modules.scala 50:57:@43850.4]
  assign _T_91300 = $signed(buffer_0_346) + $signed(buffer_3_347); // @[Modules.scala 50:57:@43868.4]
  assign _T_91301 = _T_91300[10:0]; // @[Modules.scala 50:57:@43869.4]
  assign buffer_11_565 = $signed(_T_91301); // @[Modules.scala 50:57:@43870.4]
  assign _T_91303 = $signed(buffer_2_348) + $signed(buffer_1_349); // @[Modules.scala 50:57:@43872.4]
  assign _T_91304 = _T_91303[10:0]; // @[Modules.scala 50:57:@43873.4]
  assign buffer_11_566 = $signed(_T_91304); // @[Modules.scala 50:57:@43874.4]
  assign _T_91306 = $signed(buffer_5_350) + $signed(buffer_1_351); // @[Modules.scala 50:57:@43876.4]
  assign _T_91307 = _T_91306[10:0]; // @[Modules.scala 50:57:@43877.4]
  assign buffer_11_567 = $signed(_T_91307); // @[Modules.scala 50:57:@43878.4]
  assign buffer_11_361 = {{6{_T_90594[4]}},_T_90594}; // @[Modules.scala 32:22:@8.4]
  assign _T_91321 = $signed(buffer_1_360) + $signed(buffer_11_361); // @[Modules.scala 50:57:@43896.4]
  assign _T_91322 = _T_91321[10:0]; // @[Modules.scala 50:57:@43897.4]
  assign buffer_11_572 = $signed(_T_91322); // @[Modules.scala 50:57:@43898.4]
  assign _T_91348 = $signed(buffer_2_378) + $signed(buffer_9_379); // @[Modules.scala 50:57:@43932.4]
  assign _T_91349 = _T_91348[10:0]; // @[Modules.scala 50:57:@43933.4]
  assign buffer_11_581 = $signed(_T_91349); // @[Modules.scala 50:57:@43934.4]
  assign _T_91369 = $signed(buffer_3_392) + $signed(buffer_6_393); // @[Modules.scala 53:83:@43960.4]
  assign _T_91370 = _T_91369[10:0]; // @[Modules.scala 53:83:@43961.4]
  assign buffer_11_588 = $signed(_T_91370); // @[Modules.scala 53:83:@43962.4]
  assign _T_91372 = $signed(buffer_10_394) + $signed(buffer_1_395); // @[Modules.scala 53:83:@43964.4]
  assign _T_91373 = _T_91372[10:0]; // @[Modules.scala 53:83:@43965.4]
  assign buffer_11_589 = $signed(_T_91373); // @[Modules.scala 53:83:@43966.4]
  assign _T_91375 = $signed(buffer_11_396) + $signed(buffer_11_397); // @[Modules.scala 53:83:@43968.4]
  assign _T_91376 = _T_91375[10:0]; // @[Modules.scala 53:83:@43969.4]
  assign buffer_11_590 = $signed(_T_91376); // @[Modules.scala 53:83:@43970.4]
  assign _T_91378 = $signed(buffer_0_398) + $signed(buffer_11_399); // @[Modules.scala 53:83:@43972.4]
  assign _T_91379 = _T_91378[10:0]; // @[Modules.scala 53:83:@43973.4]
  assign buffer_11_591 = $signed(_T_91379); // @[Modules.scala 53:83:@43974.4]
  assign _T_91381 = $signed(buffer_1_400) + $signed(buffer_11_401); // @[Modules.scala 53:83:@43976.4]
  assign _T_91382 = _T_91381[10:0]; // @[Modules.scala 53:83:@43977.4]
  assign buffer_11_592 = $signed(_T_91382); // @[Modules.scala 53:83:@43978.4]
  assign _T_91384 = $signed(buffer_2_402) + $signed(buffer_11_403); // @[Modules.scala 53:83:@43980.4]
  assign _T_91385 = _T_91384[10:0]; // @[Modules.scala 53:83:@43981.4]
  assign buffer_11_593 = $signed(_T_91385); // @[Modules.scala 53:83:@43982.4]
  assign _T_91387 = $signed(buffer_1_404) + $signed(buffer_11_405); // @[Modules.scala 53:83:@43984.4]
  assign _T_91388 = _T_91387[10:0]; // @[Modules.scala 53:83:@43985.4]
  assign buffer_11_594 = $signed(_T_91388); // @[Modules.scala 53:83:@43986.4]
  assign _T_91390 = $signed(buffer_11_406) + $signed(buffer_1_407); // @[Modules.scala 53:83:@43988.4]
  assign _T_91391 = _T_91390[10:0]; // @[Modules.scala 53:83:@43989.4]
  assign buffer_11_595 = $signed(_T_91391); // @[Modules.scala 53:83:@43990.4]
  assign _T_91393 = $signed(buffer_3_408) + $signed(buffer_11_409); // @[Modules.scala 53:83:@43992.4]
  assign _T_91394 = _T_91393[10:0]; // @[Modules.scala 53:83:@43993.4]
  assign buffer_11_596 = $signed(_T_91394); // @[Modules.scala 53:83:@43994.4]
  assign _T_91399 = $signed(buffer_0_412) + $signed(buffer_11_413); // @[Modules.scala 53:83:@44000.4]
  assign _T_91400 = _T_91399[10:0]; // @[Modules.scala 53:83:@44001.4]
  assign buffer_11_598 = $signed(_T_91400); // @[Modules.scala 53:83:@44002.4]
  assign _T_91402 = $signed(buffer_11_414) + $signed(buffer_6_415); // @[Modules.scala 53:83:@44004.4]
  assign _T_91403 = _T_91402[10:0]; // @[Modules.scala 53:83:@44005.4]
  assign buffer_11_599 = $signed(_T_91403); // @[Modules.scala 53:83:@44006.4]
  assign _T_91414 = $signed(buffer_0_422) + $signed(buffer_7_423); // @[Modules.scala 53:83:@44020.4]
  assign _T_91415 = _T_91414[10:0]; // @[Modules.scala 53:83:@44021.4]
  assign buffer_11_603 = $signed(_T_91415); // @[Modules.scala 53:83:@44022.4]
  assign _T_91417 = $signed(buffer_6_424) + $signed(buffer_7_425); // @[Modules.scala 53:83:@44024.4]
  assign _T_91418 = _T_91417[10:0]; // @[Modules.scala 53:83:@44025.4]
  assign buffer_11_604 = $signed(_T_91418); // @[Modules.scala 53:83:@44026.4]
  assign _T_91420 = $signed(buffer_11_426) + $signed(buffer_11_427); // @[Modules.scala 53:83:@44028.4]
  assign _T_91421 = _T_91420[10:0]; // @[Modules.scala 53:83:@44029.4]
  assign buffer_11_605 = $signed(_T_91421); // @[Modules.scala 53:83:@44030.4]
  assign _T_91426 = $signed(buffer_10_430) + $signed(buffer_4_431); // @[Modules.scala 53:83:@44036.4]
  assign _T_91427 = _T_91426[10:0]; // @[Modules.scala 53:83:@44037.4]
  assign buffer_11_607 = $signed(_T_91427); // @[Modules.scala 53:83:@44038.4]
  assign _T_91429 = $signed(buffer_2_432) + $signed(buffer_11_433); // @[Modules.scala 53:83:@44040.4]
  assign _T_91430 = _T_91429[10:0]; // @[Modules.scala 53:83:@44041.4]
  assign buffer_11_608 = $signed(_T_91430); // @[Modules.scala 53:83:@44042.4]
  assign _T_91432 = $signed(buffer_4_434) + $signed(buffer_2_435); // @[Modules.scala 53:83:@44044.4]
  assign _T_91433 = _T_91432[10:0]; // @[Modules.scala 53:83:@44045.4]
  assign buffer_11_609 = $signed(_T_91433); // @[Modules.scala 53:83:@44046.4]
  assign _T_91435 = $signed(buffer_0_436) + $signed(buffer_11_437); // @[Modules.scala 53:83:@44048.4]
  assign _T_91436 = _T_91435[10:0]; // @[Modules.scala 53:83:@44049.4]
  assign buffer_11_610 = $signed(_T_91436); // @[Modules.scala 53:83:@44050.4]
  assign _T_91438 = $signed(buffer_11_438) + $signed(buffer_11_439); // @[Modules.scala 53:83:@44052.4]
  assign _T_91439 = _T_91438[10:0]; // @[Modules.scala 53:83:@44053.4]
  assign buffer_11_611 = $signed(_T_91439); // @[Modules.scala 53:83:@44054.4]
  assign _T_91441 = $signed(buffer_2_440) + $signed(buffer_11_441); // @[Modules.scala 53:83:@44056.4]
  assign _T_91442 = _T_91441[10:0]; // @[Modules.scala 53:83:@44057.4]
  assign buffer_11_612 = $signed(_T_91442); // @[Modules.scala 53:83:@44058.4]
  assign _T_91444 = $signed(buffer_0_442) + $signed(buffer_1_443); // @[Modules.scala 53:83:@44060.4]
  assign _T_91445 = _T_91444[10:0]; // @[Modules.scala 53:83:@44061.4]
  assign buffer_11_613 = $signed(_T_91445); // @[Modules.scala 53:83:@44062.4]
  assign _T_91447 = $signed(buffer_11_444) + $signed(buffer_11_445); // @[Modules.scala 53:83:@44064.4]
  assign _T_91448 = _T_91447[10:0]; // @[Modules.scala 53:83:@44065.4]
  assign buffer_11_614 = $signed(_T_91448); // @[Modules.scala 53:83:@44066.4]
  assign _T_91453 = $signed(buffer_11_448) + $signed(buffer_0_449); // @[Modules.scala 53:83:@44072.4]
  assign _T_91454 = _T_91453[10:0]; // @[Modules.scala 53:83:@44073.4]
  assign buffer_11_616 = $signed(_T_91454); // @[Modules.scala 53:83:@44074.4]
  assign _T_91456 = $signed(buffer_11_450) + $signed(buffer_11_451); // @[Modules.scala 53:83:@44076.4]
  assign _T_91457 = _T_91456[10:0]; // @[Modules.scala 53:83:@44077.4]
  assign buffer_11_617 = $signed(_T_91457); // @[Modules.scala 53:83:@44078.4]
  assign _T_91459 = $signed(buffer_11_452) + $signed(buffer_11_453); // @[Modules.scala 53:83:@44080.4]
  assign _T_91460 = _T_91459[10:0]; // @[Modules.scala 53:83:@44081.4]
  assign buffer_11_618 = $signed(_T_91460); // @[Modules.scala 53:83:@44082.4]
  assign _T_91462 = $signed(buffer_1_454) + $signed(buffer_8_455); // @[Modules.scala 53:83:@44084.4]
  assign _T_91463 = _T_91462[10:0]; // @[Modules.scala 53:83:@44085.4]
  assign buffer_11_619 = $signed(_T_91463); // @[Modules.scala 53:83:@44086.4]
  assign _T_91465 = $signed(buffer_11_456) + $signed(buffer_6_457); // @[Modules.scala 53:83:@44088.4]
  assign _T_91466 = _T_91465[10:0]; // @[Modules.scala 53:83:@44089.4]
  assign buffer_11_620 = $signed(_T_91466); // @[Modules.scala 53:83:@44090.4]
  assign _T_91468 = $signed(buffer_11_458) + $signed(buffer_11_459); // @[Modules.scala 53:83:@44092.4]
  assign _T_91469 = _T_91468[10:0]; // @[Modules.scala 53:83:@44093.4]
  assign buffer_11_621 = $signed(_T_91469); // @[Modules.scala 53:83:@44094.4]
  assign _T_91474 = $signed(buffer_11_462) + $signed(buffer_11_463); // @[Modules.scala 53:83:@44100.4]
  assign _T_91475 = _T_91474[10:0]; // @[Modules.scala 53:83:@44101.4]
  assign buffer_11_623 = $signed(_T_91475); // @[Modules.scala 53:83:@44102.4]
  assign _T_91477 = $signed(buffer_2_464) + $signed(buffer_1_465); // @[Modules.scala 53:83:@44104.4]
  assign _T_91478 = _T_91477[10:0]; // @[Modules.scala 53:83:@44105.4]
  assign buffer_11_624 = $signed(_T_91478); // @[Modules.scala 53:83:@44106.4]
  assign _T_91486 = $signed(buffer_11_470) + $signed(buffer_0_471); // @[Modules.scala 53:83:@44116.4]
  assign _T_91487 = _T_91486[10:0]; // @[Modules.scala 53:83:@44117.4]
  assign buffer_11_627 = $signed(_T_91487); // @[Modules.scala 53:83:@44118.4]
  assign _T_91489 = $signed(buffer_11_472) + $signed(buffer_1_473); // @[Modules.scala 53:83:@44120.4]
  assign _T_91490 = _T_91489[10:0]; // @[Modules.scala 53:83:@44121.4]
  assign buffer_11_628 = $signed(_T_91490); // @[Modules.scala 53:83:@44122.4]
  assign _T_91501 = $signed(buffer_8_480) + $signed(buffer_1_481); // @[Modules.scala 53:83:@44136.4]
  assign _T_91502 = _T_91501[10:0]; // @[Modules.scala 53:83:@44137.4]
  assign buffer_11_632 = $signed(_T_91502); // @[Modules.scala 53:83:@44138.4]
  assign _T_91504 = $signed(buffer_11_482) + $signed(buffer_4_483); // @[Modules.scala 53:83:@44140.4]
  assign _T_91505 = _T_91504[10:0]; // @[Modules.scala 53:83:@44141.4]
  assign buffer_11_633 = $signed(_T_91505); // @[Modules.scala 53:83:@44142.4]
  assign _T_91507 = $signed(buffer_11_484) + $signed(buffer_11_485); // @[Modules.scala 53:83:@44144.4]
  assign _T_91508 = _T_91507[10:0]; // @[Modules.scala 53:83:@44145.4]
  assign buffer_11_634 = $signed(_T_91508); // @[Modules.scala 53:83:@44146.4]
  assign _T_91510 = $signed(buffer_5_486) + $signed(buffer_7_487); // @[Modules.scala 53:83:@44148.4]
  assign _T_91511 = _T_91510[10:0]; // @[Modules.scala 53:83:@44149.4]
  assign buffer_11_635 = $signed(_T_91511); // @[Modules.scala 53:83:@44150.4]
  assign _T_91513 = $signed(buffer_8_488) + $signed(buffer_11_489); // @[Modules.scala 53:83:@44152.4]
  assign _T_91514 = _T_91513[10:0]; // @[Modules.scala 53:83:@44153.4]
  assign buffer_11_636 = $signed(_T_91514); // @[Modules.scala 53:83:@44154.4]
  assign _T_91519 = $signed(buffer_11_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@44160.4]
  assign _T_91520 = _T_91519[10:0]; // @[Modules.scala 53:83:@44161.4]
  assign buffer_11_638 = $signed(_T_91520); // @[Modules.scala 53:83:@44162.4]
  assign _T_91522 = $signed(buffer_11_494) + $signed(buffer_3_495); // @[Modules.scala 53:83:@44164.4]
  assign _T_91523 = _T_91522[10:0]; // @[Modules.scala 53:83:@44165.4]
  assign buffer_11_639 = $signed(_T_91523); // @[Modules.scala 53:83:@44166.4]
  assign _T_91525 = $signed(buffer_2_496) + $signed(buffer_11_497); // @[Modules.scala 53:83:@44168.4]
  assign _T_91526 = _T_91525[10:0]; // @[Modules.scala 53:83:@44169.4]
  assign buffer_11_640 = $signed(_T_91526); // @[Modules.scala 53:83:@44170.4]
  assign _T_91528 = $signed(buffer_9_498) + $signed(buffer_11_499); // @[Modules.scala 53:83:@44172.4]
  assign _T_91529 = _T_91528[10:0]; // @[Modules.scala 53:83:@44173.4]
  assign buffer_11_641 = $signed(_T_91529); // @[Modules.scala 53:83:@44174.4]
  assign _T_91531 = $signed(buffer_11_500) + $signed(buffer_2_501); // @[Modules.scala 53:83:@44176.4]
  assign _T_91532 = _T_91531[10:0]; // @[Modules.scala 53:83:@44177.4]
  assign buffer_11_642 = $signed(_T_91532); // @[Modules.scala 53:83:@44178.4]
  assign _T_91534 = $signed(buffer_5_502) + $signed(buffer_0_503); // @[Modules.scala 53:83:@44180.4]
  assign _T_91535 = _T_91534[10:0]; // @[Modules.scala 53:83:@44181.4]
  assign buffer_11_643 = $signed(_T_91535); // @[Modules.scala 53:83:@44182.4]
  assign _T_91537 = $signed(buffer_11_504) + $signed(buffer_1_505); // @[Modules.scala 53:83:@44184.4]
  assign _T_91538 = _T_91537[10:0]; // @[Modules.scala 53:83:@44185.4]
  assign buffer_11_644 = $signed(_T_91538); // @[Modules.scala 53:83:@44186.4]
  assign _T_91540 = $signed(buffer_11_506) + $signed(buffer_5_507); // @[Modules.scala 53:83:@44188.4]
  assign _T_91541 = _T_91540[10:0]; // @[Modules.scala 53:83:@44189.4]
  assign buffer_11_645 = $signed(_T_91541); // @[Modules.scala 53:83:@44190.4]
  assign _T_91543 = $signed(buffer_9_508) + $signed(buffer_11_509); // @[Modules.scala 53:83:@44192.4]
  assign _T_91544 = _T_91543[10:0]; // @[Modules.scala 53:83:@44193.4]
  assign buffer_11_646 = $signed(_T_91544); // @[Modules.scala 53:83:@44194.4]
  assign _T_91546 = $signed(buffer_0_510) + $signed(buffer_11_511); // @[Modules.scala 53:83:@44196.4]
  assign _T_91547 = _T_91546[10:0]; // @[Modules.scala 53:83:@44197.4]
  assign buffer_11_647 = $signed(_T_91547); // @[Modules.scala 53:83:@44198.4]
  assign _T_91549 = $signed(buffer_11_512) + $signed(buffer_1_513); // @[Modules.scala 53:83:@44200.4]
  assign _T_91550 = _T_91549[10:0]; // @[Modules.scala 53:83:@44201.4]
  assign buffer_11_648 = $signed(_T_91550); // @[Modules.scala 53:83:@44202.4]
  assign _T_91552 = $signed(buffer_9_514) + $signed(buffer_5_515); // @[Modules.scala 53:83:@44204.4]
  assign _T_91553 = _T_91552[10:0]; // @[Modules.scala 53:83:@44205.4]
  assign buffer_11_649 = $signed(_T_91553); // @[Modules.scala 53:83:@44206.4]
  assign _T_91555 = $signed(buffer_11_516) + $signed(buffer_0_517); // @[Modules.scala 53:83:@44208.4]
  assign _T_91556 = _T_91555[10:0]; // @[Modules.scala 53:83:@44209.4]
  assign buffer_11_650 = $signed(_T_91556); // @[Modules.scala 53:83:@44210.4]
  assign _T_91558 = $signed(buffer_2_518) + $signed(buffer_8_519); // @[Modules.scala 53:83:@44212.4]
  assign _T_91559 = _T_91558[10:0]; // @[Modules.scala 53:83:@44213.4]
  assign buffer_11_651 = $signed(_T_91559); // @[Modules.scala 53:83:@44214.4]
  assign _T_91561 = $signed(buffer_11_520) + $signed(buffer_11_521); // @[Modules.scala 53:83:@44216.4]
  assign _T_91562 = _T_91561[10:0]; // @[Modules.scala 53:83:@44217.4]
  assign buffer_11_652 = $signed(_T_91562); // @[Modules.scala 53:83:@44218.4]
  assign _T_91564 = $signed(buffer_6_522) + $signed(buffer_11_523); // @[Modules.scala 53:83:@44220.4]
  assign _T_91565 = _T_91564[10:0]; // @[Modules.scala 53:83:@44221.4]
  assign buffer_11_653 = $signed(_T_91565); // @[Modules.scala 53:83:@44222.4]
  assign _T_91570 = $signed(buffer_0_526) + $signed(buffer_11_527); // @[Modules.scala 53:83:@44228.4]
  assign _T_91571 = _T_91570[10:0]; // @[Modules.scala 53:83:@44229.4]
  assign buffer_11_655 = $signed(_T_91571); // @[Modules.scala 53:83:@44230.4]
  assign _T_91573 = $signed(buffer_11_528) + $signed(buffer_3_529); // @[Modules.scala 53:83:@44232.4]
  assign _T_91574 = _T_91573[10:0]; // @[Modules.scala 53:83:@44233.4]
  assign buffer_11_656 = $signed(_T_91574); // @[Modules.scala 53:83:@44234.4]
  assign _T_91576 = $signed(buffer_11_530) + $signed(buffer_2_531); // @[Modules.scala 53:83:@44236.4]
  assign _T_91577 = _T_91576[10:0]; // @[Modules.scala 53:83:@44237.4]
  assign buffer_11_657 = $signed(_T_91577); // @[Modules.scala 53:83:@44238.4]
  assign _T_91579 = $signed(buffer_11_532) + $signed(buffer_7_533); // @[Modules.scala 53:83:@44240.4]
  assign _T_91580 = _T_91579[10:0]; // @[Modules.scala 53:83:@44241.4]
  assign buffer_11_658 = $signed(_T_91580); // @[Modules.scala 53:83:@44242.4]
  assign _T_91582 = $signed(buffer_1_534) + $signed(buffer_11_535); // @[Modules.scala 53:83:@44244.4]
  assign _T_91583 = _T_91582[10:0]; // @[Modules.scala 53:83:@44245.4]
  assign buffer_11_659 = $signed(_T_91583); // @[Modules.scala 53:83:@44246.4]
  assign _T_91585 = $signed(buffer_6_536) + $signed(buffer_11_537); // @[Modules.scala 53:83:@44248.4]
  assign _T_91586 = _T_91585[10:0]; // @[Modules.scala 53:83:@44249.4]
  assign buffer_11_660 = $signed(_T_91586); // @[Modules.scala 53:83:@44250.4]
  assign _T_91588 = $signed(buffer_1_538) + $signed(buffer_7_539); // @[Modules.scala 53:83:@44252.4]
  assign _T_91589 = _T_91588[10:0]; // @[Modules.scala 53:83:@44253.4]
  assign buffer_11_661 = $signed(_T_91589); // @[Modules.scala 53:83:@44254.4]
  assign _T_91591 = $signed(buffer_11_540) + $signed(buffer_4_541); // @[Modules.scala 53:83:@44256.4]
  assign _T_91592 = _T_91591[10:0]; // @[Modules.scala 53:83:@44257.4]
  assign buffer_11_662 = $signed(_T_91592); // @[Modules.scala 53:83:@44258.4]
  assign _T_91594 = $signed(buffer_2_542) + $signed(buffer_11_543); // @[Modules.scala 53:83:@44260.4]
  assign _T_91595 = _T_91594[10:0]; // @[Modules.scala 53:83:@44261.4]
  assign buffer_11_663 = $signed(_T_91595); // @[Modules.scala 53:83:@44262.4]
  assign _T_91597 = $signed(buffer_2_544) + $signed(buffer_11_545); // @[Modules.scala 53:83:@44264.4]
  assign _T_91598 = _T_91597[10:0]; // @[Modules.scala 53:83:@44265.4]
  assign buffer_11_664 = $signed(_T_91598); // @[Modules.scala 53:83:@44266.4]
  assign _T_91600 = $signed(buffer_7_546) + $signed(buffer_11_547); // @[Modules.scala 53:83:@44268.4]
  assign _T_91601 = _T_91600[10:0]; // @[Modules.scala 53:83:@44269.4]
  assign buffer_11_665 = $signed(_T_91601); // @[Modules.scala 53:83:@44270.4]
  assign _T_91603 = $signed(buffer_11_548) + $signed(buffer_1_549); // @[Modules.scala 53:83:@44272.4]
  assign _T_91604 = _T_91603[10:0]; // @[Modules.scala 53:83:@44273.4]
  assign buffer_11_666 = $signed(_T_91604); // @[Modules.scala 53:83:@44274.4]
  assign _T_91609 = $signed(buffer_11_552) + $signed(buffer_7_553); // @[Modules.scala 53:83:@44280.4]
  assign _T_91610 = _T_91609[10:0]; // @[Modules.scala 53:83:@44281.4]
  assign buffer_11_668 = $signed(_T_91610); // @[Modules.scala 53:83:@44282.4]
  assign _T_91612 = $signed(buffer_0_554) + $signed(buffer_11_555); // @[Modules.scala 53:83:@44284.4]
  assign _T_91613 = _T_91612[10:0]; // @[Modules.scala 53:83:@44285.4]
  assign buffer_11_669 = $signed(_T_91613); // @[Modules.scala 53:83:@44286.4]
  assign _T_91615 = $signed(buffer_1_556) + $signed(buffer_2_557); // @[Modules.scala 53:83:@44288.4]
  assign _T_91616 = _T_91615[10:0]; // @[Modules.scala 53:83:@44289.4]
  assign buffer_11_670 = $signed(_T_91616); // @[Modules.scala 53:83:@44290.4]
  assign _T_91618 = $signed(buffer_4_558) + $signed(buffer_2_559); // @[Modules.scala 53:83:@44292.4]
  assign _T_91619 = _T_91618[10:0]; // @[Modules.scala 53:83:@44293.4]
  assign buffer_11_671 = $signed(_T_91619); // @[Modules.scala 53:83:@44294.4]
  assign _T_91621 = $signed(buffer_11_560) + $signed(buffer_2_561); // @[Modules.scala 53:83:@44296.4]
  assign _T_91622 = _T_91621[10:0]; // @[Modules.scala 53:83:@44297.4]
  assign buffer_11_672 = $signed(_T_91622); // @[Modules.scala 53:83:@44298.4]
  assign _T_91627 = $signed(buffer_0_564) + $signed(buffer_11_565); // @[Modules.scala 53:83:@44304.4]
  assign _T_91628 = _T_91627[10:0]; // @[Modules.scala 53:83:@44305.4]
  assign buffer_11_674 = $signed(_T_91628); // @[Modules.scala 53:83:@44306.4]
  assign _T_91630 = $signed(buffer_11_566) + $signed(buffer_11_567); // @[Modules.scala 53:83:@44308.4]
  assign _T_91631 = _T_91630[10:0]; // @[Modules.scala 53:83:@44309.4]
  assign buffer_11_675 = $signed(_T_91631); // @[Modules.scala 53:83:@44310.4]
  assign _T_91639 = $signed(buffer_11_572) + $signed(buffer_0_573); // @[Modules.scala 53:83:@44320.4]
  assign _T_91640 = _T_91639[10:0]; // @[Modules.scala 53:83:@44321.4]
  assign buffer_11_678 = $signed(_T_91640); // @[Modules.scala 53:83:@44322.4]
  assign _T_91651 = $signed(buffer_9_580) + $signed(buffer_11_581); // @[Modules.scala 53:83:@44336.4]
  assign _T_91652 = _T_91651[10:0]; // @[Modules.scala 53:83:@44337.4]
  assign buffer_11_682 = $signed(_T_91652); // @[Modules.scala 53:83:@44338.4]
  assign _T_91663 = $signed(buffer_11_588) + $signed(buffer_11_589); // @[Modules.scala 56:109:@44352.4]
  assign _T_91664 = _T_91663[10:0]; // @[Modules.scala 56:109:@44353.4]
  assign buffer_11_686 = $signed(_T_91664); // @[Modules.scala 56:109:@44354.4]
  assign _T_91666 = $signed(buffer_11_590) + $signed(buffer_11_591); // @[Modules.scala 56:109:@44356.4]
  assign _T_91667 = _T_91666[10:0]; // @[Modules.scala 56:109:@44357.4]
  assign buffer_11_687 = $signed(_T_91667); // @[Modules.scala 56:109:@44358.4]
  assign _T_91669 = $signed(buffer_11_592) + $signed(buffer_11_593); // @[Modules.scala 56:109:@44360.4]
  assign _T_91670 = _T_91669[10:0]; // @[Modules.scala 56:109:@44361.4]
  assign buffer_11_688 = $signed(_T_91670); // @[Modules.scala 56:109:@44362.4]
  assign _T_91672 = $signed(buffer_11_594) + $signed(buffer_11_595); // @[Modules.scala 56:109:@44364.4]
  assign _T_91673 = _T_91672[10:0]; // @[Modules.scala 56:109:@44365.4]
  assign buffer_11_689 = $signed(_T_91673); // @[Modules.scala 56:109:@44366.4]
  assign _T_91675 = $signed(buffer_11_596) + $signed(buffer_3_597); // @[Modules.scala 56:109:@44368.4]
  assign _T_91676 = _T_91675[10:0]; // @[Modules.scala 56:109:@44369.4]
  assign buffer_11_690 = $signed(_T_91676); // @[Modules.scala 56:109:@44370.4]
  assign _T_91678 = $signed(buffer_11_598) + $signed(buffer_11_599); // @[Modules.scala 56:109:@44372.4]
  assign _T_91679 = _T_91678[10:0]; // @[Modules.scala 56:109:@44373.4]
  assign buffer_11_691 = $signed(_T_91679); // @[Modules.scala 56:109:@44374.4]
  assign _T_91684 = $signed(buffer_6_602) + $signed(buffer_11_603); // @[Modules.scala 56:109:@44380.4]
  assign _T_91685 = _T_91684[10:0]; // @[Modules.scala 56:109:@44381.4]
  assign buffer_11_693 = $signed(_T_91685); // @[Modules.scala 56:109:@44382.4]
  assign _T_91687 = $signed(buffer_11_604) + $signed(buffer_11_605); // @[Modules.scala 56:109:@44384.4]
  assign _T_91688 = _T_91687[10:0]; // @[Modules.scala 56:109:@44385.4]
  assign buffer_11_694 = $signed(_T_91688); // @[Modules.scala 56:109:@44386.4]
  assign _T_91690 = $signed(buffer_2_606) + $signed(buffer_11_607); // @[Modules.scala 56:109:@44388.4]
  assign _T_91691 = _T_91690[10:0]; // @[Modules.scala 56:109:@44389.4]
  assign buffer_11_695 = $signed(_T_91691); // @[Modules.scala 56:109:@44390.4]
  assign _T_91693 = $signed(buffer_11_608) + $signed(buffer_11_609); // @[Modules.scala 56:109:@44392.4]
  assign _T_91694 = _T_91693[10:0]; // @[Modules.scala 56:109:@44393.4]
  assign buffer_11_696 = $signed(_T_91694); // @[Modules.scala 56:109:@44394.4]
  assign _T_91696 = $signed(buffer_11_610) + $signed(buffer_11_611); // @[Modules.scala 56:109:@44396.4]
  assign _T_91697 = _T_91696[10:0]; // @[Modules.scala 56:109:@44397.4]
  assign buffer_11_697 = $signed(_T_91697); // @[Modules.scala 56:109:@44398.4]
  assign _T_91699 = $signed(buffer_11_612) + $signed(buffer_11_613); // @[Modules.scala 56:109:@44400.4]
  assign _T_91700 = _T_91699[10:0]; // @[Modules.scala 56:109:@44401.4]
  assign buffer_11_698 = $signed(_T_91700); // @[Modules.scala 56:109:@44402.4]
  assign _T_91702 = $signed(buffer_11_614) + $signed(buffer_7_615); // @[Modules.scala 56:109:@44404.4]
  assign _T_91703 = _T_91702[10:0]; // @[Modules.scala 56:109:@44405.4]
  assign buffer_11_699 = $signed(_T_91703); // @[Modules.scala 56:109:@44406.4]
  assign _T_91705 = $signed(buffer_11_616) + $signed(buffer_11_617); // @[Modules.scala 56:109:@44408.4]
  assign _T_91706 = _T_91705[10:0]; // @[Modules.scala 56:109:@44409.4]
  assign buffer_11_700 = $signed(_T_91706); // @[Modules.scala 56:109:@44410.4]
  assign _T_91708 = $signed(buffer_11_618) + $signed(buffer_11_619); // @[Modules.scala 56:109:@44412.4]
  assign _T_91709 = _T_91708[10:0]; // @[Modules.scala 56:109:@44413.4]
  assign buffer_11_701 = $signed(_T_91709); // @[Modules.scala 56:109:@44414.4]
  assign _T_91711 = $signed(buffer_11_620) + $signed(buffer_11_621); // @[Modules.scala 56:109:@44416.4]
  assign _T_91712 = _T_91711[10:0]; // @[Modules.scala 56:109:@44417.4]
  assign buffer_11_702 = $signed(_T_91712); // @[Modules.scala 56:109:@44418.4]
  assign _T_91714 = $signed(buffer_7_622) + $signed(buffer_11_623); // @[Modules.scala 56:109:@44420.4]
  assign _T_91715 = _T_91714[10:0]; // @[Modules.scala 56:109:@44421.4]
  assign buffer_11_703 = $signed(_T_91715); // @[Modules.scala 56:109:@44422.4]
  assign _T_91717 = $signed(buffer_11_624) + $signed(buffer_9_625); // @[Modules.scala 56:109:@44424.4]
  assign _T_91718 = _T_91717[10:0]; // @[Modules.scala 56:109:@44425.4]
  assign buffer_11_704 = $signed(_T_91718); // @[Modules.scala 56:109:@44426.4]
  assign _T_91720 = $signed(buffer_1_626) + $signed(buffer_11_627); // @[Modules.scala 56:109:@44428.4]
  assign _T_91721 = _T_91720[10:0]; // @[Modules.scala 56:109:@44429.4]
  assign buffer_11_705 = $signed(_T_91721); // @[Modules.scala 56:109:@44430.4]
  assign _T_91723 = $signed(buffer_11_628) + $signed(buffer_1_629); // @[Modules.scala 56:109:@44432.4]
  assign _T_91724 = _T_91723[10:0]; // @[Modules.scala 56:109:@44433.4]
  assign buffer_11_706 = $signed(_T_91724); // @[Modules.scala 56:109:@44434.4]
  assign _T_91729 = $signed(buffer_11_632) + $signed(buffer_11_633); // @[Modules.scala 56:109:@44440.4]
  assign _T_91730 = _T_91729[10:0]; // @[Modules.scala 56:109:@44441.4]
  assign buffer_11_708 = $signed(_T_91730); // @[Modules.scala 56:109:@44442.4]
  assign _T_91732 = $signed(buffer_11_634) + $signed(buffer_11_635); // @[Modules.scala 56:109:@44444.4]
  assign _T_91733 = _T_91732[10:0]; // @[Modules.scala 56:109:@44445.4]
  assign buffer_11_709 = $signed(_T_91733); // @[Modules.scala 56:109:@44446.4]
  assign _T_91735 = $signed(buffer_11_636) + $signed(buffer_3_637); // @[Modules.scala 56:109:@44448.4]
  assign _T_91736 = _T_91735[10:0]; // @[Modules.scala 56:109:@44449.4]
  assign buffer_11_710 = $signed(_T_91736); // @[Modules.scala 56:109:@44450.4]
  assign _T_91738 = $signed(buffer_11_638) + $signed(buffer_11_639); // @[Modules.scala 56:109:@44452.4]
  assign _T_91739 = _T_91738[10:0]; // @[Modules.scala 56:109:@44453.4]
  assign buffer_11_711 = $signed(_T_91739); // @[Modules.scala 56:109:@44454.4]
  assign _T_91741 = $signed(buffer_11_640) + $signed(buffer_11_641); // @[Modules.scala 56:109:@44456.4]
  assign _T_91742 = _T_91741[10:0]; // @[Modules.scala 56:109:@44457.4]
  assign buffer_11_712 = $signed(_T_91742); // @[Modules.scala 56:109:@44458.4]
  assign _T_91744 = $signed(buffer_11_642) + $signed(buffer_11_643); // @[Modules.scala 56:109:@44460.4]
  assign _T_91745 = _T_91744[10:0]; // @[Modules.scala 56:109:@44461.4]
  assign buffer_11_713 = $signed(_T_91745); // @[Modules.scala 56:109:@44462.4]
  assign _T_91747 = $signed(buffer_11_644) + $signed(buffer_11_645); // @[Modules.scala 56:109:@44464.4]
  assign _T_91748 = _T_91747[10:0]; // @[Modules.scala 56:109:@44465.4]
  assign buffer_11_714 = $signed(_T_91748); // @[Modules.scala 56:109:@44466.4]
  assign _T_91750 = $signed(buffer_11_646) + $signed(buffer_11_647); // @[Modules.scala 56:109:@44468.4]
  assign _T_91751 = _T_91750[10:0]; // @[Modules.scala 56:109:@44469.4]
  assign buffer_11_715 = $signed(_T_91751); // @[Modules.scala 56:109:@44470.4]
  assign _T_91753 = $signed(buffer_11_648) + $signed(buffer_11_649); // @[Modules.scala 56:109:@44472.4]
  assign _T_91754 = _T_91753[10:0]; // @[Modules.scala 56:109:@44473.4]
  assign buffer_11_716 = $signed(_T_91754); // @[Modules.scala 56:109:@44474.4]
  assign _T_91756 = $signed(buffer_11_650) + $signed(buffer_11_651); // @[Modules.scala 56:109:@44476.4]
  assign _T_91757 = _T_91756[10:0]; // @[Modules.scala 56:109:@44477.4]
  assign buffer_11_717 = $signed(_T_91757); // @[Modules.scala 56:109:@44478.4]
  assign _T_91759 = $signed(buffer_11_652) + $signed(buffer_11_653); // @[Modules.scala 56:109:@44480.4]
  assign _T_91760 = _T_91759[10:0]; // @[Modules.scala 56:109:@44481.4]
  assign buffer_11_718 = $signed(_T_91760); // @[Modules.scala 56:109:@44482.4]
  assign _T_91762 = $signed(buffer_2_654) + $signed(buffer_11_655); // @[Modules.scala 56:109:@44484.4]
  assign _T_91763 = _T_91762[10:0]; // @[Modules.scala 56:109:@44485.4]
  assign buffer_11_719 = $signed(_T_91763); // @[Modules.scala 56:109:@44486.4]
  assign _T_91765 = $signed(buffer_11_656) + $signed(buffer_11_657); // @[Modules.scala 56:109:@44488.4]
  assign _T_91766 = _T_91765[10:0]; // @[Modules.scala 56:109:@44489.4]
  assign buffer_11_720 = $signed(_T_91766); // @[Modules.scala 56:109:@44490.4]
  assign _T_91768 = $signed(buffer_11_658) + $signed(buffer_11_659); // @[Modules.scala 56:109:@44492.4]
  assign _T_91769 = _T_91768[10:0]; // @[Modules.scala 56:109:@44493.4]
  assign buffer_11_721 = $signed(_T_91769); // @[Modules.scala 56:109:@44494.4]
  assign _T_91771 = $signed(buffer_11_660) + $signed(buffer_11_661); // @[Modules.scala 56:109:@44496.4]
  assign _T_91772 = _T_91771[10:0]; // @[Modules.scala 56:109:@44497.4]
  assign buffer_11_722 = $signed(_T_91772); // @[Modules.scala 56:109:@44498.4]
  assign _T_91774 = $signed(buffer_11_662) + $signed(buffer_11_663); // @[Modules.scala 56:109:@44500.4]
  assign _T_91775 = _T_91774[10:0]; // @[Modules.scala 56:109:@44501.4]
  assign buffer_11_723 = $signed(_T_91775); // @[Modules.scala 56:109:@44502.4]
  assign _T_91777 = $signed(buffer_11_664) + $signed(buffer_11_665); // @[Modules.scala 56:109:@44504.4]
  assign _T_91778 = _T_91777[10:0]; // @[Modules.scala 56:109:@44505.4]
  assign buffer_11_724 = $signed(_T_91778); // @[Modules.scala 56:109:@44506.4]
  assign _T_91780 = $signed(buffer_11_666) + $signed(buffer_2_667); // @[Modules.scala 56:109:@44508.4]
  assign _T_91781 = _T_91780[10:0]; // @[Modules.scala 56:109:@44509.4]
  assign buffer_11_725 = $signed(_T_91781); // @[Modules.scala 56:109:@44510.4]
  assign _T_91783 = $signed(buffer_11_668) + $signed(buffer_11_669); // @[Modules.scala 56:109:@44512.4]
  assign _T_91784 = _T_91783[10:0]; // @[Modules.scala 56:109:@44513.4]
  assign buffer_11_726 = $signed(_T_91784); // @[Modules.scala 56:109:@44514.4]
  assign _T_91786 = $signed(buffer_11_670) + $signed(buffer_11_671); // @[Modules.scala 56:109:@44516.4]
  assign _T_91787 = _T_91786[10:0]; // @[Modules.scala 56:109:@44517.4]
  assign buffer_11_727 = $signed(_T_91787); // @[Modules.scala 56:109:@44518.4]
  assign _T_91789 = $signed(buffer_11_672) + $signed(buffer_7_673); // @[Modules.scala 56:109:@44520.4]
  assign _T_91790 = _T_91789[10:0]; // @[Modules.scala 56:109:@44521.4]
  assign buffer_11_728 = $signed(_T_91790); // @[Modules.scala 56:109:@44522.4]
  assign _T_91792 = $signed(buffer_11_674) + $signed(buffer_11_675); // @[Modules.scala 56:109:@44524.4]
  assign _T_91793 = _T_91792[10:0]; // @[Modules.scala 56:109:@44525.4]
  assign buffer_11_729 = $signed(_T_91793); // @[Modules.scala 56:109:@44526.4]
  assign _T_91798 = $signed(buffer_11_678) + $signed(buffer_10_679); // @[Modules.scala 56:109:@44532.4]
  assign _T_91799 = _T_91798[10:0]; // @[Modules.scala 56:109:@44533.4]
  assign buffer_11_731 = $signed(_T_91799); // @[Modules.scala 56:109:@44534.4]
  assign _T_91804 = $signed(buffer_11_682) + $signed(buffer_6_683); // @[Modules.scala 56:109:@44540.4]
  assign _T_91805 = _T_91804[10:0]; // @[Modules.scala 56:109:@44541.4]
  assign buffer_11_733 = $signed(_T_91805); // @[Modules.scala 56:109:@44542.4]
  assign _T_91810 = $signed(buffer_11_686) + $signed(buffer_11_687); // @[Modules.scala 63:156:@44549.4]
  assign _T_91811 = _T_91810[10:0]; // @[Modules.scala 63:156:@44550.4]
  assign buffer_11_736 = $signed(_T_91811); // @[Modules.scala 63:156:@44551.4]
  assign _T_91813 = $signed(buffer_11_736) + $signed(buffer_11_688); // @[Modules.scala 63:156:@44553.4]
  assign _T_91814 = _T_91813[10:0]; // @[Modules.scala 63:156:@44554.4]
  assign buffer_11_737 = $signed(_T_91814); // @[Modules.scala 63:156:@44555.4]
  assign _T_91816 = $signed(buffer_11_737) + $signed(buffer_11_689); // @[Modules.scala 63:156:@44557.4]
  assign _T_91817 = _T_91816[10:0]; // @[Modules.scala 63:156:@44558.4]
  assign buffer_11_738 = $signed(_T_91817); // @[Modules.scala 63:156:@44559.4]
  assign _T_91819 = $signed(buffer_11_738) + $signed(buffer_11_690); // @[Modules.scala 63:156:@44561.4]
  assign _T_91820 = _T_91819[10:0]; // @[Modules.scala 63:156:@44562.4]
  assign buffer_11_739 = $signed(_T_91820); // @[Modules.scala 63:156:@44563.4]
  assign _T_91822 = $signed(buffer_11_739) + $signed(buffer_11_691); // @[Modules.scala 63:156:@44565.4]
  assign _T_91823 = _T_91822[10:0]; // @[Modules.scala 63:156:@44566.4]
  assign buffer_11_740 = $signed(_T_91823); // @[Modules.scala 63:156:@44567.4]
  assign _T_91825 = $signed(buffer_11_740) + $signed(buffer_8_692); // @[Modules.scala 63:156:@44569.4]
  assign _T_91826 = _T_91825[10:0]; // @[Modules.scala 63:156:@44570.4]
  assign buffer_11_741 = $signed(_T_91826); // @[Modules.scala 63:156:@44571.4]
  assign _T_91828 = $signed(buffer_11_741) + $signed(buffer_11_693); // @[Modules.scala 63:156:@44573.4]
  assign _T_91829 = _T_91828[10:0]; // @[Modules.scala 63:156:@44574.4]
  assign buffer_11_742 = $signed(_T_91829); // @[Modules.scala 63:156:@44575.4]
  assign _T_91831 = $signed(buffer_11_742) + $signed(buffer_11_694); // @[Modules.scala 63:156:@44577.4]
  assign _T_91832 = _T_91831[10:0]; // @[Modules.scala 63:156:@44578.4]
  assign buffer_11_743 = $signed(_T_91832); // @[Modules.scala 63:156:@44579.4]
  assign _T_91834 = $signed(buffer_11_743) + $signed(buffer_11_695); // @[Modules.scala 63:156:@44581.4]
  assign _T_91835 = _T_91834[10:0]; // @[Modules.scala 63:156:@44582.4]
  assign buffer_11_744 = $signed(_T_91835); // @[Modules.scala 63:156:@44583.4]
  assign _T_91837 = $signed(buffer_11_744) + $signed(buffer_11_696); // @[Modules.scala 63:156:@44585.4]
  assign _T_91838 = _T_91837[10:0]; // @[Modules.scala 63:156:@44586.4]
  assign buffer_11_745 = $signed(_T_91838); // @[Modules.scala 63:156:@44587.4]
  assign _T_91840 = $signed(buffer_11_745) + $signed(buffer_11_697); // @[Modules.scala 63:156:@44589.4]
  assign _T_91841 = _T_91840[10:0]; // @[Modules.scala 63:156:@44590.4]
  assign buffer_11_746 = $signed(_T_91841); // @[Modules.scala 63:156:@44591.4]
  assign _T_91843 = $signed(buffer_11_746) + $signed(buffer_11_698); // @[Modules.scala 63:156:@44593.4]
  assign _T_91844 = _T_91843[10:0]; // @[Modules.scala 63:156:@44594.4]
  assign buffer_11_747 = $signed(_T_91844); // @[Modules.scala 63:156:@44595.4]
  assign _T_91846 = $signed(buffer_11_747) + $signed(buffer_11_699); // @[Modules.scala 63:156:@44597.4]
  assign _T_91847 = _T_91846[10:0]; // @[Modules.scala 63:156:@44598.4]
  assign buffer_11_748 = $signed(_T_91847); // @[Modules.scala 63:156:@44599.4]
  assign _T_91849 = $signed(buffer_11_748) + $signed(buffer_11_700); // @[Modules.scala 63:156:@44601.4]
  assign _T_91850 = _T_91849[10:0]; // @[Modules.scala 63:156:@44602.4]
  assign buffer_11_749 = $signed(_T_91850); // @[Modules.scala 63:156:@44603.4]
  assign _T_91852 = $signed(buffer_11_749) + $signed(buffer_11_701); // @[Modules.scala 63:156:@44605.4]
  assign _T_91853 = _T_91852[10:0]; // @[Modules.scala 63:156:@44606.4]
  assign buffer_11_750 = $signed(_T_91853); // @[Modules.scala 63:156:@44607.4]
  assign _T_91855 = $signed(buffer_11_750) + $signed(buffer_11_702); // @[Modules.scala 63:156:@44609.4]
  assign _T_91856 = _T_91855[10:0]; // @[Modules.scala 63:156:@44610.4]
  assign buffer_11_751 = $signed(_T_91856); // @[Modules.scala 63:156:@44611.4]
  assign _T_91858 = $signed(buffer_11_751) + $signed(buffer_11_703); // @[Modules.scala 63:156:@44613.4]
  assign _T_91859 = _T_91858[10:0]; // @[Modules.scala 63:156:@44614.4]
  assign buffer_11_752 = $signed(_T_91859); // @[Modules.scala 63:156:@44615.4]
  assign _T_91861 = $signed(buffer_11_752) + $signed(buffer_11_704); // @[Modules.scala 63:156:@44617.4]
  assign _T_91862 = _T_91861[10:0]; // @[Modules.scala 63:156:@44618.4]
  assign buffer_11_753 = $signed(_T_91862); // @[Modules.scala 63:156:@44619.4]
  assign _T_91864 = $signed(buffer_11_753) + $signed(buffer_11_705); // @[Modules.scala 63:156:@44621.4]
  assign _T_91865 = _T_91864[10:0]; // @[Modules.scala 63:156:@44622.4]
  assign buffer_11_754 = $signed(_T_91865); // @[Modules.scala 63:156:@44623.4]
  assign _T_91867 = $signed(buffer_11_754) + $signed(buffer_11_706); // @[Modules.scala 63:156:@44625.4]
  assign _T_91868 = _T_91867[10:0]; // @[Modules.scala 63:156:@44626.4]
  assign buffer_11_755 = $signed(_T_91868); // @[Modules.scala 63:156:@44627.4]
  assign _T_91870 = $signed(buffer_11_755) + $signed(buffer_0_707); // @[Modules.scala 63:156:@44629.4]
  assign _T_91871 = _T_91870[10:0]; // @[Modules.scala 63:156:@44630.4]
  assign buffer_11_756 = $signed(_T_91871); // @[Modules.scala 63:156:@44631.4]
  assign _T_91873 = $signed(buffer_11_756) + $signed(buffer_11_708); // @[Modules.scala 63:156:@44633.4]
  assign _T_91874 = _T_91873[10:0]; // @[Modules.scala 63:156:@44634.4]
  assign buffer_11_757 = $signed(_T_91874); // @[Modules.scala 63:156:@44635.4]
  assign _T_91876 = $signed(buffer_11_757) + $signed(buffer_11_709); // @[Modules.scala 63:156:@44637.4]
  assign _T_91877 = _T_91876[10:0]; // @[Modules.scala 63:156:@44638.4]
  assign buffer_11_758 = $signed(_T_91877); // @[Modules.scala 63:156:@44639.4]
  assign _T_91879 = $signed(buffer_11_758) + $signed(buffer_11_710); // @[Modules.scala 63:156:@44641.4]
  assign _T_91880 = _T_91879[10:0]; // @[Modules.scala 63:156:@44642.4]
  assign buffer_11_759 = $signed(_T_91880); // @[Modules.scala 63:156:@44643.4]
  assign _T_91882 = $signed(buffer_11_759) + $signed(buffer_11_711); // @[Modules.scala 63:156:@44645.4]
  assign _T_91883 = _T_91882[10:0]; // @[Modules.scala 63:156:@44646.4]
  assign buffer_11_760 = $signed(_T_91883); // @[Modules.scala 63:156:@44647.4]
  assign _T_91885 = $signed(buffer_11_760) + $signed(buffer_11_712); // @[Modules.scala 63:156:@44649.4]
  assign _T_91886 = _T_91885[10:0]; // @[Modules.scala 63:156:@44650.4]
  assign buffer_11_761 = $signed(_T_91886); // @[Modules.scala 63:156:@44651.4]
  assign _T_91888 = $signed(buffer_11_761) + $signed(buffer_11_713); // @[Modules.scala 63:156:@44653.4]
  assign _T_91889 = _T_91888[10:0]; // @[Modules.scala 63:156:@44654.4]
  assign buffer_11_762 = $signed(_T_91889); // @[Modules.scala 63:156:@44655.4]
  assign _T_91891 = $signed(buffer_11_762) + $signed(buffer_11_714); // @[Modules.scala 63:156:@44657.4]
  assign _T_91892 = _T_91891[10:0]; // @[Modules.scala 63:156:@44658.4]
  assign buffer_11_763 = $signed(_T_91892); // @[Modules.scala 63:156:@44659.4]
  assign _T_91894 = $signed(buffer_11_763) + $signed(buffer_11_715); // @[Modules.scala 63:156:@44661.4]
  assign _T_91895 = _T_91894[10:0]; // @[Modules.scala 63:156:@44662.4]
  assign buffer_11_764 = $signed(_T_91895); // @[Modules.scala 63:156:@44663.4]
  assign _T_91897 = $signed(buffer_11_764) + $signed(buffer_11_716); // @[Modules.scala 63:156:@44665.4]
  assign _T_91898 = _T_91897[10:0]; // @[Modules.scala 63:156:@44666.4]
  assign buffer_11_765 = $signed(_T_91898); // @[Modules.scala 63:156:@44667.4]
  assign _T_91900 = $signed(buffer_11_765) + $signed(buffer_11_717); // @[Modules.scala 63:156:@44669.4]
  assign _T_91901 = _T_91900[10:0]; // @[Modules.scala 63:156:@44670.4]
  assign buffer_11_766 = $signed(_T_91901); // @[Modules.scala 63:156:@44671.4]
  assign _T_91903 = $signed(buffer_11_766) + $signed(buffer_11_718); // @[Modules.scala 63:156:@44673.4]
  assign _T_91904 = _T_91903[10:0]; // @[Modules.scala 63:156:@44674.4]
  assign buffer_11_767 = $signed(_T_91904); // @[Modules.scala 63:156:@44675.4]
  assign _T_91906 = $signed(buffer_11_767) + $signed(buffer_11_719); // @[Modules.scala 63:156:@44677.4]
  assign _T_91907 = _T_91906[10:0]; // @[Modules.scala 63:156:@44678.4]
  assign buffer_11_768 = $signed(_T_91907); // @[Modules.scala 63:156:@44679.4]
  assign _T_91909 = $signed(buffer_11_768) + $signed(buffer_11_720); // @[Modules.scala 63:156:@44681.4]
  assign _T_91910 = _T_91909[10:0]; // @[Modules.scala 63:156:@44682.4]
  assign buffer_11_769 = $signed(_T_91910); // @[Modules.scala 63:156:@44683.4]
  assign _T_91912 = $signed(buffer_11_769) + $signed(buffer_11_721); // @[Modules.scala 63:156:@44685.4]
  assign _T_91913 = _T_91912[10:0]; // @[Modules.scala 63:156:@44686.4]
  assign buffer_11_770 = $signed(_T_91913); // @[Modules.scala 63:156:@44687.4]
  assign _T_91915 = $signed(buffer_11_770) + $signed(buffer_11_722); // @[Modules.scala 63:156:@44689.4]
  assign _T_91916 = _T_91915[10:0]; // @[Modules.scala 63:156:@44690.4]
  assign buffer_11_771 = $signed(_T_91916); // @[Modules.scala 63:156:@44691.4]
  assign _T_91918 = $signed(buffer_11_771) + $signed(buffer_11_723); // @[Modules.scala 63:156:@44693.4]
  assign _T_91919 = _T_91918[10:0]; // @[Modules.scala 63:156:@44694.4]
  assign buffer_11_772 = $signed(_T_91919); // @[Modules.scala 63:156:@44695.4]
  assign _T_91921 = $signed(buffer_11_772) + $signed(buffer_11_724); // @[Modules.scala 63:156:@44697.4]
  assign _T_91922 = _T_91921[10:0]; // @[Modules.scala 63:156:@44698.4]
  assign buffer_11_773 = $signed(_T_91922); // @[Modules.scala 63:156:@44699.4]
  assign _T_91924 = $signed(buffer_11_773) + $signed(buffer_11_725); // @[Modules.scala 63:156:@44701.4]
  assign _T_91925 = _T_91924[10:0]; // @[Modules.scala 63:156:@44702.4]
  assign buffer_11_774 = $signed(_T_91925); // @[Modules.scala 63:156:@44703.4]
  assign _T_91927 = $signed(buffer_11_774) + $signed(buffer_11_726); // @[Modules.scala 63:156:@44705.4]
  assign _T_91928 = _T_91927[10:0]; // @[Modules.scala 63:156:@44706.4]
  assign buffer_11_775 = $signed(_T_91928); // @[Modules.scala 63:156:@44707.4]
  assign _T_91930 = $signed(buffer_11_775) + $signed(buffer_11_727); // @[Modules.scala 63:156:@44709.4]
  assign _T_91931 = _T_91930[10:0]; // @[Modules.scala 63:156:@44710.4]
  assign buffer_11_776 = $signed(_T_91931); // @[Modules.scala 63:156:@44711.4]
  assign _T_91933 = $signed(buffer_11_776) + $signed(buffer_11_728); // @[Modules.scala 63:156:@44713.4]
  assign _T_91934 = _T_91933[10:0]; // @[Modules.scala 63:156:@44714.4]
  assign buffer_11_777 = $signed(_T_91934); // @[Modules.scala 63:156:@44715.4]
  assign _T_91936 = $signed(buffer_11_777) + $signed(buffer_11_729); // @[Modules.scala 63:156:@44717.4]
  assign _T_91937 = _T_91936[10:0]; // @[Modules.scala 63:156:@44718.4]
  assign buffer_11_778 = $signed(_T_91937); // @[Modules.scala 63:156:@44719.4]
  assign _T_91939 = $signed(buffer_11_778) + $signed(buffer_2_730); // @[Modules.scala 63:156:@44721.4]
  assign _T_91940 = _T_91939[10:0]; // @[Modules.scala 63:156:@44722.4]
  assign buffer_11_779 = $signed(_T_91940); // @[Modules.scala 63:156:@44723.4]
  assign _T_91942 = $signed(buffer_11_779) + $signed(buffer_11_731); // @[Modules.scala 63:156:@44725.4]
  assign _T_91943 = _T_91942[10:0]; // @[Modules.scala 63:156:@44726.4]
  assign buffer_11_780 = $signed(_T_91943); // @[Modules.scala 63:156:@44727.4]
  assign _T_91945 = $signed(buffer_11_780) + $signed(buffer_4_732); // @[Modules.scala 63:156:@44729.4]
  assign _T_91946 = _T_91945[10:0]; // @[Modules.scala 63:156:@44730.4]
  assign buffer_11_781 = $signed(_T_91946); // @[Modules.scala 63:156:@44731.4]
  assign _T_91948 = $signed(buffer_11_781) + $signed(buffer_11_733); // @[Modules.scala 63:156:@44733.4]
  assign _T_91949 = _T_91948[10:0]; // @[Modules.scala 63:156:@44734.4]
  assign buffer_11_782 = $signed(_T_91949); // @[Modules.scala 63:156:@44735.4]
  assign _T_91951 = $signed(buffer_11_782) + $signed(buffer_2_734); // @[Modules.scala 63:156:@44737.4]
  assign _T_91952 = _T_91951[10:0]; // @[Modules.scala 63:156:@44738.4]
  assign buffer_11_783 = $signed(_T_91952); // @[Modules.scala 63:156:@44739.4]
  assign _T_91991 = $signed(io_in_14) - $signed(io_in_15); // @[Modules.scala 40:46:@44782.4]
  assign _T_91992 = _T_91991[4:0]; // @[Modules.scala 40:46:@44783.4]
  assign _T_91993 = $signed(_T_91992); // @[Modules.scala 40:46:@44784.4]
  assign _T_92493 = $signed(io_in_226) - $signed(io_in_227); // @[Modules.scala 40:46:@45344.4]
  assign _T_92494 = _T_92493[4:0]; // @[Modules.scala 40:46:@45345.4]
  assign _T_92495 = $signed(_T_92494); // @[Modules.scala 40:46:@45346.4]
  assign _T_92715 = $signed(io_in_310) - $signed(io_in_311); // @[Modules.scala 40:46:@45584.4]
  assign _T_92716 = _T_92715[4:0]; // @[Modules.scala 40:46:@45585.4]
  assign _T_92717 = $signed(_T_92716); // @[Modules.scala 40:46:@45586.4]
  assign _T_92771 = $signed(_T_55242) + $signed(io_in_327); // @[Modules.scala 43:47:@45640.4]
  assign _T_92772 = _T_92771[4:0]; // @[Modules.scala 43:47:@45641.4]
  assign _T_92773 = $signed(_T_92772); // @[Modules.scala 43:47:@45642.4]
  assign _T_92778 = $signed(_T_58354) + $signed(io_in_329); // @[Modules.scala 43:47:@45647.4]
  assign _T_92779 = _T_92778[4:0]; // @[Modules.scala 43:47:@45648.4]
  assign _T_92780 = $signed(_T_92779); // @[Modules.scala 43:47:@45649.4]
  assign _T_92784 = $signed(io_in_332) - $signed(io_in_333); // @[Modules.scala 40:46:@45655.4]
  assign _T_92785 = _T_92784[4:0]; // @[Modules.scala 40:46:@45656.4]
  assign _T_92786 = $signed(_T_92785); // @[Modules.scala 40:46:@45657.4]
  assign _T_93012 = $signed(_T_64898) + $signed(io_in_413); // @[Modules.scala 43:47:@45896.4]
  assign _T_93013 = _T_93012[4:0]; // @[Modules.scala 43:47:@45897.4]
  assign _T_93014 = $signed(_T_93013); // @[Modules.scala 43:47:@45898.4]
  assign _T_93144 = $signed(io_in_476) - $signed(io_in_477); // @[Modules.scala 40:46:@46051.4]
  assign _T_93145 = _T_93144[4:0]; // @[Modules.scala 40:46:@46052.4]
  assign _T_93146 = $signed(_T_93145); // @[Modules.scala 40:46:@46053.4]
  assign _T_93166 = $signed(io_in_488) - $signed(io_in_489); // @[Modules.scala 40:46:@46078.4]
  assign _T_93167 = _T_93166[4:0]; // @[Modules.scala 40:46:@46079.4]
  assign _T_93168 = $signed(_T_93167); // @[Modules.scala 40:46:@46080.4]
  assign _T_93173 = $signed(_T_58777) + $signed(io_in_491); // @[Modules.scala 43:47:@46085.4]
  assign _T_93174 = _T_93173[4:0]; // @[Modules.scala 43:47:@46086.4]
  assign _T_93175 = $signed(_T_93174); // @[Modules.scala 43:47:@46087.4]
  assign _T_93314 = $signed(io_in_560) + $signed(io_in_561); // @[Modules.scala 37:46:@46252.4]
  assign _T_93315 = _T_93314[4:0]; // @[Modules.scala 37:46:@46253.4]
  assign _T_93316 = $signed(_T_93315); // @[Modules.scala 37:46:@46254.4]
  assign _T_93346 = $signed(_T_71330) + $signed(io_in_577); // @[Modules.scala 43:47:@46290.4]
  assign _T_93347 = _T_93346[4:0]; // @[Modules.scala 43:47:@46291.4]
  assign _T_93348 = $signed(_T_93347); // @[Modules.scala 43:47:@46292.4]
  assign _T_93374 = $signed(_T_55889) + $signed(io_in_593); // @[Modules.scala 43:47:@46325.4]
  assign _T_93375 = _T_93374[4:0]; // @[Modules.scala 43:47:@46326.4]
  assign _T_93376 = $signed(_T_93375); // @[Modules.scala 43:47:@46327.4]
  assign _T_93425 = $signed(_T_62298) + $signed(io_in_619); // @[Modules.scala 43:47:@46386.4]
  assign _T_93426 = _T_93425[4:0]; // @[Modules.scala 43:47:@46387.4]
  assign _T_93427 = $signed(_T_93426); // @[Modules.scala 43:47:@46388.4]
  assign _T_93858 = $signed(io_in_776) - $signed(io_in_777); // @[Modules.scala 40:46:@46849.4]
  assign _T_93859 = _T_93858[4:0]; // @[Modules.scala 40:46:@46850.4]
  assign _T_93860 = $signed(_T_93859); // @[Modules.scala 40:46:@46851.4]
  assign _T_93878 = $signed(buffer_7_0) + $signed(buffer_4_1); // @[Modules.scala 50:57:@46871.4]
  assign _T_93879 = _T_93878[10:0]; // @[Modules.scala 50:57:@46872.4]
  assign buffer_12_392 = $signed(_T_93879); // @[Modules.scala 50:57:@46873.4]
  assign _T_93881 = $signed(buffer_9_2) + $signed(buffer_2_3); // @[Modules.scala 50:57:@46875.4]
  assign _T_93882 = _T_93881[10:0]; // @[Modules.scala 50:57:@46876.4]
  assign buffer_12_393 = $signed(_T_93882); // @[Modules.scala 50:57:@46877.4]
  assign buffer_12_7 = {{6{_T_91993[4]}},_T_91993}; // @[Modules.scala 32:22:@8.4]
  assign _T_93887 = $signed(buffer_1_6) + $signed(buffer_12_7); // @[Modules.scala 50:57:@46883.4]
  assign _T_93888 = _T_93887[10:0]; // @[Modules.scala 50:57:@46884.4]
  assign buffer_12_395 = $signed(_T_93888); // @[Modules.scala 50:57:@46885.4]
  assign _T_93890 = $signed(buffer_7_8) + $signed(buffer_1_9); // @[Modules.scala 50:57:@46887.4]
  assign _T_93891 = _T_93890[10:0]; // @[Modules.scala 50:57:@46888.4]
  assign buffer_12_396 = $signed(_T_93891); // @[Modules.scala 50:57:@46889.4]
  assign _T_93893 = $signed(buffer_7_10) + $signed(buffer_1_11); // @[Modules.scala 50:57:@46891.4]
  assign _T_93894 = _T_93893[10:0]; // @[Modules.scala 50:57:@46892.4]
  assign buffer_12_397 = $signed(_T_93894); // @[Modules.scala 50:57:@46893.4]
  assign _T_93896 = $signed(buffer_0_12) + $signed(buffer_1_13); // @[Modules.scala 50:57:@46895.4]
  assign _T_93897 = _T_93896[10:0]; // @[Modules.scala 50:57:@46896.4]
  assign buffer_12_398 = $signed(_T_93897); // @[Modules.scala 50:57:@46897.4]
  assign _T_93899 = $signed(buffer_1_14) + $signed(buffer_2_15); // @[Modules.scala 50:57:@46899.4]
  assign _T_93900 = _T_93899[10:0]; // @[Modules.scala 50:57:@46900.4]
  assign buffer_12_399 = $signed(_T_93900); // @[Modules.scala 50:57:@46901.4]
  assign _T_93959 = $signed(buffer_1_54) + $signed(buffer_3_55); // @[Modules.scala 50:57:@46979.4]
  assign _T_93960 = _T_93959[10:0]; // @[Modules.scala 50:57:@46980.4]
  assign buffer_12_419 = $signed(_T_93960); // @[Modules.scala 50:57:@46981.4]
  assign _T_93965 = $signed(buffer_2_58) + $signed(buffer_4_59); // @[Modules.scala 50:57:@46987.4]
  assign _T_93966 = _T_93965[10:0]; // @[Modules.scala 50:57:@46988.4]
  assign buffer_12_421 = $signed(_T_93966); // @[Modules.scala 50:57:@46989.4]
  assign _T_93971 = $signed(buffer_8_62) + $signed(buffer_0_63); // @[Modules.scala 50:57:@46995.4]
  assign _T_93972 = _T_93971[10:0]; // @[Modules.scala 50:57:@46996.4]
  assign buffer_12_423 = $signed(_T_93972); // @[Modules.scala 50:57:@46997.4]
  assign _T_93977 = $signed(buffer_5_66) + $signed(buffer_3_67); // @[Modules.scala 50:57:@47003.4]
  assign _T_93978 = _T_93977[10:0]; // @[Modules.scala 50:57:@47004.4]
  assign buffer_12_425 = $signed(_T_93978); // @[Modules.scala 50:57:@47005.4]
  assign _T_93980 = $signed(buffer_8_68) + $signed(buffer_1_69); // @[Modules.scala 50:57:@47007.4]
  assign _T_93981 = _T_93980[10:0]; // @[Modules.scala 50:57:@47008.4]
  assign buffer_12_426 = $signed(_T_93981); // @[Modules.scala 50:57:@47009.4]
  assign _T_93986 = $signed(buffer_0_72) + $signed(buffer_1_73); // @[Modules.scala 50:57:@47015.4]
  assign _T_93987 = _T_93986[10:0]; // @[Modules.scala 50:57:@47016.4]
  assign buffer_12_428 = $signed(_T_93987); // @[Modules.scala 50:57:@47017.4]
  assign _T_93989 = $signed(buffer_0_74) + $signed(buffer_1_75); // @[Modules.scala 50:57:@47019.4]
  assign _T_93990 = _T_93989[10:0]; // @[Modules.scala 50:57:@47020.4]
  assign buffer_12_429 = $signed(_T_93990); // @[Modules.scala 50:57:@47021.4]
  assign _T_93995 = $signed(buffer_9_78) + $signed(buffer_3_79); // @[Modules.scala 50:57:@47027.4]
  assign _T_93996 = _T_93995[10:0]; // @[Modules.scala 50:57:@47028.4]
  assign buffer_12_431 = $signed(_T_93996); // @[Modules.scala 50:57:@47029.4]
  assign _T_94001 = $signed(buffer_1_82) + $signed(buffer_0_83); // @[Modules.scala 50:57:@47035.4]
  assign _T_94002 = _T_94001[10:0]; // @[Modules.scala 50:57:@47036.4]
  assign buffer_12_433 = $signed(_T_94002); // @[Modules.scala 50:57:@47037.4]
  assign _T_94016 = $signed(buffer_4_92) + $signed(buffer_3_93); // @[Modules.scala 50:57:@47055.4]
  assign _T_94017 = _T_94016[10:0]; // @[Modules.scala 50:57:@47056.4]
  assign buffer_12_438 = $signed(_T_94017); // @[Modules.scala 50:57:@47057.4]
  assign _T_94028 = $signed(buffer_0_100) + $signed(buffer_5_101); // @[Modules.scala 50:57:@47071.4]
  assign _T_94029 = _T_94028[10:0]; // @[Modules.scala 50:57:@47072.4]
  assign buffer_12_442 = $signed(_T_94029); // @[Modules.scala 50:57:@47073.4]
  assign _T_94031 = $signed(buffer_1_102) + $signed(buffer_0_103); // @[Modules.scala 50:57:@47075.4]
  assign _T_94032 = _T_94031[10:0]; // @[Modules.scala 50:57:@47076.4]
  assign buffer_12_443 = $signed(_T_94032); // @[Modules.scala 50:57:@47077.4]
  assign _T_94037 = $signed(buffer_1_106) + $signed(buffer_2_107); // @[Modules.scala 50:57:@47083.4]
  assign _T_94038 = _T_94037[10:0]; // @[Modules.scala 50:57:@47084.4]
  assign buffer_12_445 = $signed(_T_94038); // @[Modules.scala 50:57:@47085.4]
  assign buffer_12_113 = {{6{_T_92495[4]}},_T_92495}; // @[Modules.scala 32:22:@8.4]
  assign _T_94046 = $signed(buffer_1_112) + $signed(buffer_12_113); // @[Modules.scala 50:57:@47095.4]
  assign _T_94047 = _T_94046[10:0]; // @[Modules.scala 50:57:@47096.4]
  assign buffer_12_448 = $signed(_T_94047); // @[Modules.scala 50:57:@47097.4]
  assign _T_94052 = $signed(buffer_7_116) + $signed(buffer_3_117); // @[Modules.scala 50:57:@47103.4]
  assign _T_94053 = _T_94052[10:0]; // @[Modules.scala 50:57:@47104.4]
  assign buffer_12_450 = $signed(_T_94053); // @[Modules.scala 50:57:@47105.4]
  assign _T_94055 = $signed(buffer_1_118) + $signed(buffer_3_119); // @[Modules.scala 50:57:@47107.4]
  assign _T_94056 = _T_94055[10:0]; // @[Modules.scala 50:57:@47108.4]
  assign buffer_12_451 = $signed(_T_94056); // @[Modules.scala 50:57:@47109.4]
  assign _T_94067 = $signed(buffer_3_126) + $signed(buffer_8_127); // @[Modules.scala 50:57:@47123.4]
  assign _T_94068 = _T_94067[10:0]; // @[Modules.scala 50:57:@47124.4]
  assign buffer_12_455 = $signed(_T_94068); // @[Modules.scala 50:57:@47125.4]
  assign _T_94070 = $signed(buffer_4_128) + $signed(buffer_0_129); // @[Modules.scala 50:57:@47127.4]
  assign _T_94071 = _T_94070[10:0]; // @[Modules.scala 50:57:@47128.4]
  assign buffer_12_456 = $signed(_T_94071); // @[Modules.scala 50:57:@47129.4]
  assign _T_94073 = $signed(buffer_1_130) + $signed(buffer_0_131); // @[Modules.scala 50:57:@47131.4]
  assign _T_94074 = _T_94073[10:0]; // @[Modules.scala 50:57:@47132.4]
  assign buffer_12_457 = $signed(_T_94074); // @[Modules.scala 50:57:@47133.4]
  assign _T_94076 = $signed(buffer_3_132) + $signed(buffer_9_133); // @[Modules.scala 50:57:@47135.4]
  assign _T_94077 = _T_94076[10:0]; // @[Modules.scala 50:57:@47136.4]
  assign buffer_12_458 = $signed(_T_94077); // @[Modules.scala 50:57:@47137.4]
  assign _T_94079 = $signed(buffer_3_134) + $signed(buffer_11_135); // @[Modules.scala 50:57:@47139.4]
  assign _T_94080 = _T_94079[10:0]; // @[Modules.scala 50:57:@47140.4]
  assign buffer_12_459 = $signed(_T_94080); // @[Modules.scala 50:57:@47141.4]
  assign _T_94088 = $signed(buffer_3_140) + $signed(buffer_8_141); // @[Modules.scala 50:57:@47151.4]
  assign _T_94089 = _T_94088[10:0]; // @[Modules.scala 50:57:@47152.4]
  assign buffer_12_462 = $signed(_T_94089); // @[Modules.scala 50:57:@47153.4]
  assign _T_94100 = $signed(buffer_0_148) + $signed(buffer_3_149); // @[Modules.scala 50:57:@47167.4]
  assign _T_94101 = _T_94100[10:0]; // @[Modules.scala 50:57:@47168.4]
  assign buffer_12_466 = $signed(_T_94101); // @[Modules.scala 50:57:@47169.4]
  assign _T_94103 = $signed(buffer_6_150) + $signed(buffer_5_151); // @[Modules.scala 50:57:@47171.4]
  assign _T_94104 = _T_94103[10:0]; // @[Modules.scala 50:57:@47172.4]
  assign buffer_12_467 = $signed(_T_94104); // @[Modules.scala 50:57:@47173.4]
  assign buffer_12_155 = {{6{_T_92717[4]}},_T_92717}; // @[Modules.scala 32:22:@8.4]
  assign _T_94109 = $signed(buffer_10_154) + $signed(buffer_12_155); // @[Modules.scala 50:57:@47179.4]
  assign _T_94110 = _T_94109[10:0]; // @[Modules.scala 50:57:@47180.4]
  assign buffer_12_469 = $signed(_T_94110); // @[Modules.scala 50:57:@47181.4]
  assign buffer_12_163 = {{6{_T_92773[4]}},_T_92773}; // @[Modules.scala 32:22:@8.4]
  assign _T_94121 = $signed(buffer_1_162) + $signed(buffer_12_163); // @[Modules.scala 50:57:@47195.4]
  assign _T_94122 = _T_94121[10:0]; // @[Modules.scala 50:57:@47196.4]
  assign buffer_12_473 = $signed(_T_94122); // @[Modules.scala 50:57:@47197.4]
  assign buffer_12_164 = {{6{_T_92780[4]}},_T_92780}; // @[Modules.scala 32:22:@8.4]
  assign _T_94124 = $signed(buffer_12_164) + $signed(buffer_5_165); // @[Modules.scala 50:57:@47199.4]
  assign _T_94125 = _T_94124[10:0]; // @[Modules.scala 50:57:@47200.4]
  assign buffer_12_474 = $signed(_T_94125); // @[Modules.scala 50:57:@47201.4]
  assign buffer_12_166 = {{6{_T_92786[4]}},_T_92786}; // @[Modules.scala 32:22:@8.4]
  assign _T_94127 = $signed(buffer_12_166) + $signed(buffer_6_167); // @[Modules.scala 50:57:@47203.4]
  assign _T_94128 = _T_94127[10:0]; // @[Modules.scala 50:57:@47204.4]
  assign buffer_12_475 = $signed(_T_94128); // @[Modules.scala 50:57:@47205.4]
  assign _T_94130 = $signed(buffer_5_168) + $signed(buffer_3_169); // @[Modules.scala 50:57:@47207.4]
  assign _T_94131 = _T_94130[10:0]; // @[Modules.scala 50:57:@47208.4]
  assign buffer_12_476 = $signed(_T_94131); // @[Modules.scala 50:57:@47209.4]
  assign _T_94172 = $signed(buffer_0_196) + $signed(buffer_3_197); // @[Modules.scala 50:57:@47263.4]
  assign _T_94173 = _T_94172[10:0]; // @[Modules.scala 50:57:@47264.4]
  assign buffer_12_490 = $signed(_T_94173); // @[Modules.scala 50:57:@47265.4]
  assign _T_94175 = $signed(buffer_3_198) + $signed(buffer_4_199); // @[Modules.scala 50:57:@47267.4]
  assign _T_94176 = _T_94175[10:0]; // @[Modules.scala 50:57:@47268.4]
  assign buffer_12_491 = $signed(_T_94176); // @[Modules.scala 50:57:@47269.4]
  assign buffer_12_206 = {{6{_T_93014[4]}},_T_93014}; // @[Modules.scala 32:22:@8.4]
  assign _T_94187 = $signed(buffer_12_206) + $signed(buffer_0_207); // @[Modules.scala 50:57:@47283.4]
  assign _T_94188 = _T_94187[10:0]; // @[Modules.scala 50:57:@47284.4]
  assign buffer_12_495 = $signed(_T_94188); // @[Modules.scala 50:57:@47285.4]
  assign _T_94193 = $signed(buffer_3_210) + $signed(buffer_0_211); // @[Modules.scala 50:57:@47291.4]
  assign _T_94194 = _T_94193[10:0]; // @[Modules.scala 50:57:@47292.4]
  assign buffer_12_497 = $signed(_T_94194); // @[Modules.scala 50:57:@47293.4]
  assign _T_94208 = $signed(buffer_0_220) + $signed(buffer_1_221); // @[Modules.scala 50:57:@47311.4]
  assign _T_94209 = _T_94208[10:0]; // @[Modules.scala 50:57:@47312.4]
  assign buffer_12_502 = $signed(_T_94209); // @[Modules.scala 50:57:@47313.4]
  assign _T_94223 = $signed(buffer_0_230) + $signed(buffer_1_231); // @[Modules.scala 50:57:@47331.4]
  assign _T_94224 = _T_94223[10:0]; // @[Modules.scala 50:57:@47332.4]
  assign buffer_12_507 = $signed(_T_94224); // @[Modules.scala 50:57:@47333.4]
  assign _T_94229 = $signed(buffer_1_234) + $signed(buffer_0_235); // @[Modules.scala 50:57:@47339.4]
  assign _T_94230 = _T_94229[10:0]; // @[Modules.scala 50:57:@47340.4]
  assign buffer_12_509 = $signed(_T_94230); // @[Modules.scala 50:57:@47341.4]
  assign buffer_12_238 = {{6{_T_93146[4]}},_T_93146}; // @[Modules.scala 32:22:@8.4]
  assign _T_94235 = $signed(buffer_12_238) + $signed(buffer_7_239); // @[Modules.scala 50:57:@47347.4]
  assign _T_94236 = _T_94235[10:0]; // @[Modules.scala 50:57:@47348.4]
  assign buffer_12_511 = $signed(_T_94236); // @[Modules.scala 50:57:@47349.4]
  assign buffer_12_244 = {{6{_T_93168[4]}},_T_93168}; // @[Modules.scala 32:22:@8.4]
  assign buffer_12_245 = {{6{_T_93175[4]}},_T_93175}; // @[Modules.scala 32:22:@8.4]
  assign _T_94244 = $signed(buffer_12_244) + $signed(buffer_12_245); // @[Modules.scala 50:57:@47359.4]
  assign _T_94245 = _T_94244[10:0]; // @[Modules.scala 50:57:@47360.4]
  assign buffer_12_514 = $signed(_T_94245); // @[Modules.scala 50:57:@47361.4]
  assign _T_94256 = $signed(buffer_3_252) + $signed(buffer_2_253); // @[Modules.scala 50:57:@47375.4]
  assign _T_94257 = _T_94256[10:0]; // @[Modules.scala 50:57:@47376.4]
  assign buffer_12_518 = $signed(_T_94257); // @[Modules.scala 50:57:@47377.4]
  assign _T_94259 = $signed(buffer_8_254) + $signed(buffer_10_255); // @[Modules.scala 50:57:@47379.4]
  assign _T_94260 = _T_94259[10:0]; // @[Modules.scala 50:57:@47380.4]
  assign buffer_12_519 = $signed(_T_94260); // @[Modules.scala 50:57:@47381.4]
  assign _T_94265 = $signed(buffer_2_258) + $signed(buffer_4_259); // @[Modules.scala 50:57:@47387.4]
  assign _T_94266 = _T_94265[10:0]; // @[Modules.scala 50:57:@47388.4]
  assign buffer_12_521 = $signed(_T_94266); // @[Modules.scala 50:57:@47389.4]
  assign _T_94271 = $signed(buffer_7_262) + $signed(buffer_0_263); // @[Modules.scala 50:57:@47395.4]
  assign _T_94272 = _T_94271[10:0]; // @[Modules.scala 50:57:@47396.4]
  assign buffer_12_523 = $signed(_T_94272); // @[Modules.scala 50:57:@47397.4]
  assign _T_94277 = $signed(buffer_1_266) + $signed(buffer_2_267); // @[Modules.scala 50:57:@47403.4]
  assign _T_94278 = _T_94277[10:0]; // @[Modules.scala 50:57:@47404.4]
  assign buffer_12_525 = $signed(_T_94278); // @[Modules.scala 50:57:@47405.4]
  assign _T_94289 = $signed(buffer_0_274) + $signed(buffer_2_275); // @[Modules.scala 50:57:@47419.4]
  assign _T_94290 = _T_94289[10:0]; // @[Modules.scala 50:57:@47420.4]
  assign buffer_12_529 = $signed(_T_94290); // @[Modules.scala 50:57:@47421.4]
  assign buffer_12_280 = {{6{_T_93316[4]}},_T_93316}; // @[Modules.scala 32:22:@8.4]
  assign _T_94298 = $signed(buffer_12_280) + $signed(buffer_0_281); // @[Modules.scala 50:57:@47431.4]
  assign _T_94299 = _T_94298[10:0]; // @[Modules.scala 50:57:@47432.4]
  assign buffer_12_532 = $signed(_T_94299); // @[Modules.scala 50:57:@47433.4]
  assign buffer_12_288 = {{6{_T_93348[4]}},_T_93348}; // @[Modules.scala 32:22:@8.4]
  assign _T_94310 = $signed(buffer_12_288) + $signed(buffer_1_289); // @[Modules.scala 50:57:@47447.4]
  assign _T_94311 = _T_94310[10:0]; // @[Modules.scala 50:57:@47448.4]
  assign buffer_12_536 = $signed(_T_94311); // @[Modules.scala 50:57:@47449.4]
  assign _T_94319 = $signed(buffer_2_294) + $signed(buffer_1_295); // @[Modules.scala 50:57:@47459.4]
  assign _T_94320 = _T_94319[10:0]; // @[Modules.scala 50:57:@47460.4]
  assign buffer_12_539 = $signed(_T_94320); // @[Modules.scala 50:57:@47461.4]
  assign buffer_12_296 = {{6{_T_93376[4]}},_T_93376}; // @[Modules.scala 32:22:@8.4]
  assign _T_94322 = $signed(buffer_12_296) + $signed(buffer_2_297); // @[Modules.scala 50:57:@47463.4]
  assign _T_94323 = _T_94322[10:0]; // @[Modules.scala 50:57:@47464.4]
  assign buffer_12_540 = $signed(_T_94323); // @[Modules.scala 50:57:@47465.4]
  assign _T_94325 = $signed(buffer_8_298) + $signed(buffer_1_299); // @[Modules.scala 50:57:@47467.4]
  assign _T_94326 = _T_94325[10:0]; // @[Modules.scala 50:57:@47468.4]
  assign buffer_12_541 = $signed(_T_94326); // @[Modules.scala 50:57:@47469.4]
  assign buffer_12_309 = {{6{_T_93427[4]}},_T_93427}; // @[Modules.scala 32:22:@8.4]
  assign _T_94340 = $signed(buffer_2_308) + $signed(buffer_12_309); // @[Modules.scala 50:57:@47487.4]
  assign _T_94341 = _T_94340[10:0]; // @[Modules.scala 50:57:@47488.4]
  assign buffer_12_546 = $signed(_T_94341); // @[Modules.scala 50:57:@47489.4]
  assign _T_94361 = $signed(buffer_10_322) + $signed(buffer_6_323); // @[Modules.scala 50:57:@47515.4]
  assign _T_94362 = _T_94361[10:0]; // @[Modules.scala 50:57:@47516.4]
  assign buffer_12_553 = $signed(_T_94362); // @[Modules.scala 50:57:@47517.4]
  assign _T_94379 = $signed(buffer_0_334) + $signed(buffer_4_335); // @[Modules.scala 50:57:@47539.4]
  assign _T_94380 = _T_94379[10:0]; // @[Modules.scala 50:57:@47540.4]
  assign buffer_12_559 = $signed(_T_94380); // @[Modules.scala 50:57:@47541.4]
  assign _T_94388 = $signed(buffer_1_340) + $signed(buffer_2_341); // @[Modules.scala 50:57:@47551.4]
  assign _T_94389 = _T_94388[10:0]; // @[Modules.scala 50:57:@47552.4]
  assign buffer_12_562 = $signed(_T_94389); // @[Modules.scala 50:57:@47553.4]
  assign _T_94391 = $signed(buffer_1_342) + $signed(buffer_0_343); // @[Modules.scala 50:57:@47555.4]
  assign _T_94392 = _T_94391[10:0]; // @[Modules.scala 50:57:@47556.4]
  assign buffer_12_563 = $signed(_T_94392); // @[Modules.scala 50:57:@47557.4]
  assign _T_94400 = $signed(buffer_0_348) + $signed(buffer_4_349); // @[Modules.scala 50:57:@47567.4]
  assign _T_94401 = _T_94400[10:0]; // @[Modules.scala 50:57:@47568.4]
  assign buffer_12_566 = $signed(_T_94401); // @[Modules.scala 50:57:@47569.4]
  assign _T_94403 = $signed(buffer_0_350) + $signed(buffer_5_351); // @[Modules.scala 50:57:@47571.4]
  assign _T_94404 = _T_94403[10:0]; // @[Modules.scala 50:57:@47572.4]
  assign buffer_12_567 = $signed(_T_94404); // @[Modules.scala 50:57:@47573.4]
  assign _T_94424 = $signed(buffer_0_364) + $signed(buffer_3_365); // @[Modules.scala 50:57:@47599.4]
  assign _T_94425 = _T_94424[10:0]; // @[Modules.scala 50:57:@47600.4]
  assign buffer_12_574 = $signed(_T_94425); // @[Modules.scala 50:57:@47601.4]
  assign _T_94442 = $signed(buffer_8_376) + $signed(buffer_0_377); // @[Modules.scala 50:57:@47623.4]
  assign _T_94443 = _T_94442[10:0]; // @[Modules.scala 50:57:@47624.4]
  assign buffer_12_580 = $signed(_T_94443); // @[Modules.scala 50:57:@47625.4]
  assign _T_94445 = $signed(buffer_3_378) + $signed(buffer_8_379); // @[Modules.scala 50:57:@47627.4]
  assign _T_94446 = _T_94445[10:0]; // @[Modules.scala 50:57:@47628.4]
  assign buffer_12_581 = $signed(_T_94446); // @[Modules.scala 50:57:@47629.4]
  assign _T_94451 = $signed(buffer_8_382) + $signed(buffer_4_383); // @[Modules.scala 50:57:@47635.4]
  assign _T_94452 = _T_94451[10:0]; // @[Modules.scala 50:57:@47636.4]
  assign buffer_12_583 = $signed(_T_94452); // @[Modules.scala 50:57:@47637.4]
  assign buffer_12_388 = {{6{_T_93860[4]}},_T_93860}; // @[Modules.scala 32:22:@8.4]
  assign _T_94460 = $signed(buffer_12_388) + $signed(buffer_0_389); // @[Modules.scala 50:57:@47647.4]
  assign _T_94461 = _T_94460[10:0]; // @[Modules.scala 50:57:@47648.4]
  assign buffer_12_586 = $signed(_T_94461); // @[Modules.scala 50:57:@47649.4]
  assign _T_94466 = $signed(buffer_12_392) + $signed(buffer_12_393); // @[Modules.scala 53:83:@47655.4]
  assign _T_94467 = _T_94466[10:0]; // @[Modules.scala 53:83:@47656.4]
  assign buffer_12_588 = $signed(_T_94467); // @[Modules.scala 53:83:@47657.4]
  assign _T_94469 = $signed(buffer_1_394) + $signed(buffer_12_395); // @[Modules.scala 53:83:@47659.4]
  assign _T_94470 = _T_94469[10:0]; // @[Modules.scala 53:83:@47660.4]
  assign buffer_12_589 = $signed(_T_94470); // @[Modules.scala 53:83:@47661.4]
  assign _T_94472 = $signed(buffer_12_396) + $signed(buffer_12_397); // @[Modules.scala 53:83:@47663.4]
  assign _T_94473 = _T_94472[10:0]; // @[Modules.scala 53:83:@47664.4]
  assign buffer_12_590 = $signed(_T_94473); // @[Modules.scala 53:83:@47665.4]
  assign _T_94475 = $signed(buffer_12_398) + $signed(buffer_12_399); // @[Modules.scala 53:83:@47667.4]
  assign _T_94476 = _T_94475[10:0]; // @[Modules.scala 53:83:@47668.4]
  assign buffer_12_591 = $signed(_T_94476); // @[Modules.scala 53:83:@47669.4]
  assign _T_94487 = $signed(buffer_1_406) + $signed(buffer_7_407); // @[Modules.scala 53:83:@47683.4]
  assign _T_94488 = _T_94487[10:0]; // @[Modules.scala 53:83:@47684.4]
  assign buffer_12_595 = $signed(_T_94488); // @[Modules.scala 53:83:@47685.4]
  assign _T_94496 = $signed(buffer_1_412) + $signed(buffer_4_413); // @[Modules.scala 53:83:@47695.4]
  assign _T_94497 = _T_94496[10:0]; // @[Modules.scala 53:83:@47696.4]
  assign buffer_12_598 = $signed(_T_94497); // @[Modules.scala 53:83:@47697.4]
  assign _T_94505 = $signed(buffer_0_418) + $signed(buffer_12_419); // @[Modules.scala 53:83:@47707.4]
  assign _T_94506 = _T_94505[10:0]; // @[Modules.scala 53:83:@47708.4]
  assign buffer_12_601 = $signed(_T_94506); // @[Modules.scala 53:83:@47709.4]
  assign _T_94508 = $signed(buffer_4_420) + $signed(buffer_12_421); // @[Modules.scala 53:83:@47711.4]
  assign _T_94509 = _T_94508[10:0]; // @[Modules.scala 53:83:@47712.4]
  assign buffer_12_602 = $signed(_T_94509); // @[Modules.scala 53:83:@47713.4]
  assign _T_94511 = $signed(buffer_4_422) + $signed(buffer_12_423); // @[Modules.scala 53:83:@47715.4]
  assign _T_94512 = _T_94511[10:0]; // @[Modules.scala 53:83:@47716.4]
  assign buffer_12_603 = $signed(_T_94512); // @[Modules.scala 53:83:@47717.4]
  assign _T_94514 = $signed(buffer_6_424) + $signed(buffer_12_425); // @[Modules.scala 53:83:@47719.4]
  assign _T_94515 = _T_94514[10:0]; // @[Modules.scala 53:83:@47720.4]
  assign buffer_12_604 = $signed(_T_94515); // @[Modules.scala 53:83:@47721.4]
  assign _T_94517 = $signed(buffer_12_426) + $signed(buffer_0_427); // @[Modules.scala 53:83:@47723.4]
  assign _T_94518 = _T_94517[10:0]; // @[Modules.scala 53:83:@47724.4]
  assign buffer_12_605 = $signed(_T_94518); // @[Modules.scala 53:83:@47725.4]
  assign _T_94520 = $signed(buffer_12_428) + $signed(buffer_12_429); // @[Modules.scala 53:83:@47727.4]
  assign _T_94521 = _T_94520[10:0]; // @[Modules.scala 53:83:@47728.4]
  assign buffer_12_606 = $signed(_T_94521); // @[Modules.scala 53:83:@47729.4]
  assign _T_94523 = $signed(buffer_4_430) + $signed(buffer_12_431); // @[Modules.scala 53:83:@47731.4]
  assign _T_94524 = _T_94523[10:0]; // @[Modules.scala 53:83:@47732.4]
  assign buffer_12_607 = $signed(_T_94524); // @[Modules.scala 53:83:@47733.4]
  assign _T_94526 = $signed(buffer_5_432) + $signed(buffer_12_433); // @[Modules.scala 53:83:@47735.4]
  assign _T_94527 = _T_94526[10:0]; // @[Modules.scala 53:83:@47736.4]
  assign buffer_12_608 = $signed(_T_94527); // @[Modules.scala 53:83:@47737.4]
  assign _T_94532 = $signed(buffer_0_436) + $signed(buffer_5_437); // @[Modules.scala 53:83:@47743.4]
  assign _T_94533 = _T_94532[10:0]; // @[Modules.scala 53:83:@47744.4]
  assign buffer_12_610 = $signed(_T_94533); // @[Modules.scala 53:83:@47745.4]
  assign _T_94535 = $signed(buffer_12_438) + $signed(buffer_9_439); // @[Modules.scala 53:83:@47747.4]
  assign _T_94536 = _T_94535[10:0]; // @[Modules.scala 53:83:@47748.4]
  assign buffer_12_611 = $signed(_T_94536); // @[Modules.scala 53:83:@47749.4]
  assign _T_94541 = $signed(buffer_12_442) + $signed(buffer_12_443); // @[Modules.scala 53:83:@47755.4]
  assign _T_94542 = _T_94541[10:0]; // @[Modules.scala 53:83:@47756.4]
  assign buffer_12_613 = $signed(_T_94542); // @[Modules.scala 53:83:@47757.4]
  assign _T_94544 = $signed(buffer_1_444) + $signed(buffer_12_445); // @[Modules.scala 53:83:@47759.4]
  assign _T_94545 = _T_94544[10:0]; // @[Modules.scala 53:83:@47760.4]
  assign buffer_12_614 = $signed(_T_94545); // @[Modules.scala 53:83:@47761.4]
  assign _T_94550 = $signed(buffer_12_448) + $signed(buffer_7_449); // @[Modules.scala 53:83:@47767.4]
  assign _T_94551 = _T_94550[10:0]; // @[Modules.scala 53:83:@47768.4]
  assign buffer_12_616 = $signed(_T_94551); // @[Modules.scala 53:83:@47769.4]
  assign _T_94553 = $signed(buffer_12_450) + $signed(buffer_12_451); // @[Modules.scala 53:83:@47771.4]
  assign _T_94554 = _T_94553[10:0]; // @[Modules.scala 53:83:@47772.4]
  assign buffer_12_617 = $signed(_T_94554); // @[Modules.scala 53:83:@47773.4]
  assign _T_94556 = $signed(buffer_1_452) + $signed(buffer_9_453); // @[Modules.scala 53:83:@47775.4]
  assign _T_94557 = _T_94556[10:0]; // @[Modules.scala 53:83:@47776.4]
  assign buffer_12_618 = $signed(_T_94557); // @[Modules.scala 53:83:@47777.4]
  assign _T_94559 = $signed(buffer_0_454) + $signed(buffer_12_455); // @[Modules.scala 53:83:@47779.4]
  assign _T_94560 = _T_94559[10:0]; // @[Modules.scala 53:83:@47780.4]
  assign buffer_12_619 = $signed(_T_94560); // @[Modules.scala 53:83:@47781.4]
  assign _T_94562 = $signed(buffer_12_456) + $signed(buffer_12_457); // @[Modules.scala 53:83:@47783.4]
  assign _T_94563 = _T_94562[10:0]; // @[Modules.scala 53:83:@47784.4]
  assign buffer_12_620 = $signed(_T_94563); // @[Modules.scala 53:83:@47785.4]
  assign _T_94565 = $signed(buffer_12_458) + $signed(buffer_12_459); // @[Modules.scala 53:83:@47787.4]
  assign _T_94566 = _T_94565[10:0]; // @[Modules.scala 53:83:@47788.4]
  assign buffer_12_621 = $signed(_T_94566); // @[Modules.scala 53:83:@47789.4]
  assign _T_94571 = $signed(buffer_12_462) + $signed(buffer_0_463); // @[Modules.scala 53:83:@47795.4]
  assign _T_94572 = _T_94571[10:0]; // @[Modules.scala 53:83:@47796.4]
  assign buffer_12_623 = $signed(_T_94572); // @[Modules.scala 53:83:@47797.4]
  assign _T_94574 = $signed(buffer_3_464) + $signed(buffer_7_465); // @[Modules.scala 53:83:@47799.4]
  assign _T_94575 = _T_94574[10:0]; // @[Modules.scala 53:83:@47800.4]
  assign buffer_12_624 = $signed(_T_94575); // @[Modules.scala 53:83:@47801.4]
  assign _T_94577 = $signed(buffer_12_466) + $signed(buffer_12_467); // @[Modules.scala 53:83:@47803.4]
  assign _T_94578 = _T_94577[10:0]; // @[Modules.scala 53:83:@47804.4]
  assign buffer_12_625 = $signed(_T_94578); // @[Modules.scala 53:83:@47805.4]
  assign _T_94580 = $signed(buffer_0_468) + $signed(buffer_12_469); // @[Modules.scala 53:83:@47807.4]
  assign _T_94581 = _T_94580[10:0]; // @[Modules.scala 53:83:@47808.4]
  assign buffer_12_626 = $signed(_T_94581); // @[Modules.scala 53:83:@47809.4]
  assign _T_94586 = $signed(buffer_0_472) + $signed(buffer_12_473); // @[Modules.scala 53:83:@47815.4]
  assign _T_94587 = _T_94586[10:0]; // @[Modules.scala 53:83:@47816.4]
  assign buffer_12_628 = $signed(_T_94587); // @[Modules.scala 53:83:@47817.4]
  assign _T_94589 = $signed(buffer_12_474) + $signed(buffer_12_475); // @[Modules.scala 53:83:@47819.4]
  assign _T_94590 = _T_94589[10:0]; // @[Modules.scala 53:83:@47820.4]
  assign buffer_12_629 = $signed(_T_94590); // @[Modules.scala 53:83:@47821.4]
  assign _T_94592 = $signed(buffer_12_476) + $signed(buffer_3_477); // @[Modules.scala 53:83:@47823.4]
  assign _T_94593 = _T_94592[10:0]; // @[Modules.scala 53:83:@47824.4]
  assign buffer_12_630 = $signed(_T_94593); // @[Modules.scala 53:83:@47825.4]
  assign _T_94598 = $signed(buffer_1_480) + $signed(buffer_0_481); // @[Modules.scala 53:83:@47831.4]
  assign _T_94599 = _T_94598[10:0]; // @[Modules.scala 53:83:@47832.4]
  assign buffer_12_632 = $signed(_T_94599); // @[Modules.scala 53:83:@47833.4]
  assign _T_94601 = $signed(buffer_11_482) + $signed(buffer_3_483); // @[Modules.scala 53:83:@47835.4]
  assign _T_94602 = _T_94601[10:0]; // @[Modules.scala 53:83:@47836.4]
  assign buffer_12_633 = $signed(_T_94602); // @[Modules.scala 53:83:@47837.4]
  assign _T_94607 = $signed(buffer_3_486) + $signed(buffer_1_487); // @[Modules.scala 53:83:@47843.4]
  assign _T_94608 = _T_94607[10:0]; // @[Modules.scala 53:83:@47844.4]
  assign buffer_12_635 = $signed(_T_94608); // @[Modules.scala 53:83:@47845.4]
  assign _T_94610 = $signed(buffer_0_488) + $signed(buffer_9_489); // @[Modules.scala 53:83:@47847.4]
  assign _T_94611 = _T_94610[10:0]; // @[Modules.scala 53:83:@47848.4]
  assign buffer_12_636 = $signed(_T_94611); // @[Modules.scala 53:83:@47849.4]
  assign _T_94613 = $signed(buffer_12_490) + $signed(buffer_12_491); // @[Modules.scala 53:83:@47851.4]
  assign _T_94614 = _T_94613[10:0]; // @[Modules.scala 53:83:@47852.4]
  assign buffer_12_637 = $signed(_T_94614); // @[Modules.scala 53:83:@47853.4]
  assign _T_94616 = $signed(buffer_4_492) + $signed(buffer_3_493); // @[Modules.scala 53:83:@47855.4]
  assign _T_94617 = _T_94616[10:0]; // @[Modules.scala 53:83:@47856.4]
  assign buffer_12_638 = $signed(_T_94617); // @[Modules.scala 53:83:@47857.4]
  assign _T_94619 = $signed(buffer_1_494) + $signed(buffer_12_495); // @[Modules.scala 53:83:@47859.4]
  assign _T_94620 = _T_94619[10:0]; // @[Modules.scala 53:83:@47860.4]
  assign buffer_12_639 = $signed(_T_94620); // @[Modules.scala 53:83:@47861.4]
  assign _T_94622 = $signed(buffer_10_496) + $signed(buffer_12_497); // @[Modules.scala 53:83:@47863.4]
  assign _T_94623 = _T_94622[10:0]; // @[Modules.scala 53:83:@47864.4]
  assign buffer_12_640 = $signed(_T_94623); // @[Modules.scala 53:83:@47865.4]
  assign _T_94631 = $signed(buffer_12_502) + $signed(buffer_3_503); // @[Modules.scala 53:83:@47875.4]
  assign _T_94632 = _T_94631[10:0]; // @[Modules.scala 53:83:@47876.4]
  assign buffer_12_643 = $signed(_T_94632); // @[Modules.scala 53:83:@47877.4]
  assign _T_94637 = $signed(buffer_0_506) + $signed(buffer_12_507); // @[Modules.scala 53:83:@47883.4]
  assign _T_94638 = _T_94637[10:0]; // @[Modules.scala 53:83:@47884.4]
  assign buffer_12_645 = $signed(_T_94638); // @[Modules.scala 53:83:@47885.4]
  assign _T_94640 = $signed(buffer_0_508) + $signed(buffer_12_509); // @[Modules.scala 53:83:@47887.4]
  assign _T_94641 = _T_94640[10:0]; // @[Modules.scala 53:83:@47888.4]
  assign buffer_12_646 = $signed(_T_94641); // @[Modules.scala 53:83:@47889.4]
  assign _T_94643 = $signed(buffer_3_510) + $signed(buffer_12_511); // @[Modules.scala 53:83:@47891.4]
  assign _T_94644 = _T_94643[10:0]; // @[Modules.scala 53:83:@47892.4]
  assign buffer_12_647 = $signed(_T_94644); // @[Modules.scala 53:83:@47893.4]
  assign _T_94646 = $signed(buffer_4_512) + $signed(buffer_0_513); // @[Modules.scala 53:83:@47895.4]
  assign _T_94647 = _T_94646[10:0]; // @[Modules.scala 53:83:@47896.4]
  assign buffer_12_648 = $signed(_T_94647); // @[Modules.scala 53:83:@47897.4]
  assign _T_94649 = $signed(buffer_12_514) + $signed(buffer_8_515); // @[Modules.scala 53:83:@47899.4]
  assign _T_94650 = _T_94649[10:0]; // @[Modules.scala 53:83:@47900.4]
  assign buffer_12_649 = $signed(_T_94650); // @[Modules.scala 53:83:@47901.4]
  assign _T_94655 = $signed(buffer_12_518) + $signed(buffer_12_519); // @[Modules.scala 53:83:@47907.4]
  assign _T_94656 = _T_94655[10:0]; // @[Modules.scala 53:83:@47908.4]
  assign buffer_12_651 = $signed(_T_94656); // @[Modules.scala 53:83:@47909.4]
  assign _T_94658 = $signed(buffer_0_520) + $signed(buffer_12_521); // @[Modules.scala 53:83:@47911.4]
  assign _T_94659 = _T_94658[10:0]; // @[Modules.scala 53:83:@47912.4]
  assign buffer_12_652 = $signed(_T_94659); // @[Modules.scala 53:83:@47913.4]
  assign _T_94661 = $signed(buffer_4_522) + $signed(buffer_12_523); // @[Modules.scala 53:83:@47915.4]
  assign _T_94662 = _T_94661[10:0]; // @[Modules.scala 53:83:@47916.4]
  assign buffer_12_653 = $signed(_T_94662); // @[Modules.scala 53:83:@47917.4]
  assign _T_94664 = $signed(buffer_3_524) + $signed(buffer_12_525); // @[Modules.scala 53:83:@47919.4]
  assign _T_94665 = _T_94664[10:0]; // @[Modules.scala 53:83:@47920.4]
  assign buffer_12_654 = $signed(_T_94665); // @[Modules.scala 53:83:@47921.4]
  assign _T_94670 = $signed(buffer_7_528) + $signed(buffer_12_529); // @[Modules.scala 53:83:@47927.4]
  assign _T_94671 = _T_94670[10:0]; // @[Modules.scala 53:83:@47928.4]
  assign buffer_12_656 = $signed(_T_94671); // @[Modules.scala 53:83:@47929.4]
  assign _T_94676 = $signed(buffer_12_532) + $signed(buffer_3_533); // @[Modules.scala 53:83:@47935.4]
  assign _T_94677 = _T_94676[10:0]; // @[Modules.scala 53:83:@47936.4]
  assign buffer_12_658 = $signed(_T_94677); // @[Modules.scala 53:83:@47937.4]
  assign _T_94682 = $signed(buffer_12_536) + $signed(buffer_4_537); // @[Modules.scala 53:83:@47943.4]
  assign _T_94683 = _T_94682[10:0]; // @[Modules.scala 53:83:@47944.4]
  assign buffer_12_660 = $signed(_T_94683); // @[Modules.scala 53:83:@47945.4]
  assign _T_94685 = $signed(buffer_3_538) + $signed(buffer_12_539); // @[Modules.scala 53:83:@47947.4]
  assign _T_94686 = _T_94685[10:0]; // @[Modules.scala 53:83:@47948.4]
  assign buffer_12_661 = $signed(_T_94686); // @[Modules.scala 53:83:@47949.4]
  assign _T_94688 = $signed(buffer_12_540) + $signed(buffer_12_541); // @[Modules.scala 53:83:@47951.4]
  assign _T_94689 = _T_94688[10:0]; // @[Modules.scala 53:83:@47952.4]
  assign buffer_12_662 = $signed(_T_94689); // @[Modules.scala 53:83:@47953.4]
  assign _T_94694 = $signed(buffer_4_544) + $signed(buffer_10_545); // @[Modules.scala 53:83:@47959.4]
  assign _T_94695 = _T_94694[10:0]; // @[Modules.scala 53:83:@47960.4]
  assign buffer_12_664 = $signed(_T_94695); // @[Modules.scala 53:83:@47961.4]
  assign _T_94697 = $signed(buffer_12_546) + $signed(buffer_3_547); // @[Modules.scala 53:83:@47963.4]
  assign _T_94698 = _T_94697[10:0]; // @[Modules.scala 53:83:@47964.4]
  assign buffer_12_665 = $signed(_T_94698); // @[Modules.scala 53:83:@47965.4]
  assign _T_94700 = $signed(buffer_8_548) + $signed(buffer_6_549); // @[Modules.scala 53:83:@47967.4]
  assign _T_94701 = _T_94700[10:0]; // @[Modules.scala 53:83:@47968.4]
  assign buffer_12_666 = $signed(_T_94701); // @[Modules.scala 53:83:@47969.4]
  assign _T_94703 = $signed(buffer_2_550) + $signed(buffer_3_551); // @[Modules.scala 53:83:@47971.4]
  assign _T_94704 = _T_94703[10:0]; // @[Modules.scala 53:83:@47972.4]
  assign buffer_12_667 = $signed(_T_94704); // @[Modules.scala 53:83:@47973.4]
  assign _T_94706 = $signed(buffer_0_552) + $signed(buffer_12_553); // @[Modules.scala 53:83:@47975.4]
  assign _T_94707 = _T_94706[10:0]; // @[Modules.scala 53:83:@47976.4]
  assign buffer_12_668 = $signed(_T_94707); // @[Modules.scala 53:83:@47977.4]
  assign _T_94709 = $signed(buffer_1_554) + $signed(buffer_8_555); // @[Modules.scala 53:83:@47979.4]
  assign _T_94710 = _T_94709[10:0]; // @[Modules.scala 53:83:@47980.4]
  assign buffer_12_669 = $signed(_T_94710); // @[Modules.scala 53:83:@47981.4]
  assign _T_94715 = $signed(buffer_5_558) + $signed(buffer_12_559); // @[Modules.scala 53:83:@47987.4]
  assign _T_94716 = _T_94715[10:0]; // @[Modules.scala 53:83:@47988.4]
  assign buffer_12_671 = $signed(_T_94716); // @[Modules.scala 53:83:@47989.4]
  assign _T_94721 = $signed(buffer_12_562) + $signed(buffer_12_563); // @[Modules.scala 53:83:@47995.4]
  assign _T_94722 = _T_94721[10:0]; // @[Modules.scala 53:83:@47996.4]
  assign buffer_12_673 = $signed(_T_94722); // @[Modules.scala 53:83:@47997.4]
  assign _T_94727 = $signed(buffer_12_566) + $signed(buffer_12_567); // @[Modules.scala 53:83:@48003.4]
  assign _T_94728 = _T_94727[10:0]; // @[Modules.scala 53:83:@48004.4]
  assign buffer_12_675 = $signed(_T_94728); // @[Modules.scala 53:83:@48005.4]
  assign _T_94739 = $signed(buffer_12_574) + $signed(buffer_1_575); // @[Modules.scala 53:83:@48019.4]
  assign _T_94740 = _T_94739[10:0]; // @[Modules.scala 53:83:@48020.4]
  assign buffer_12_679 = $signed(_T_94740); // @[Modules.scala 53:83:@48021.4]
  assign _T_94748 = $signed(buffer_12_580) + $signed(buffer_12_581); // @[Modules.scala 53:83:@48031.4]
  assign _T_94749 = _T_94748[10:0]; // @[Modules.scala 53:83:@48032.4]
  assign buffer_12_682 = $signed(_T_94749); // @[Modules.scala 53:83:@48033.4]
  assign _T_94751 = $signed(buffer_1_582) + $signed(buffer_12_583); // @[Modules.scala 53:83:@48035.4]
  assign _T_94752 = _T_94751[10:0]; // @[Modules.scala 53:83:@48036.4]
  assign buffer_12_683 = $signed(_T_94752); // @[Modules.scala 53:83:@48037.4]
  assign _T_94757 = $signed(buffer_12_586) + $signed(buffer_0_587); // @[Modules.scala 53:83:@48043.4]
  assign _T_94758 = _T_94757[10:0]; // @[Modules.scala 53:83:@48044.4]
  assign buffer_12_685 = $signed(_T_94758); // @[Modules.scala 53:83:@48045.4]
  assign _T_94760 = $signed(buffer_12_588) + $signed(buffer_12_589); // @[Modules.scala 56:109:@48047.4]
  assign _T_94761 = _T_94760[10:0]; // @[Modules.scala 56:109:@48048.4]
  assign buffer_12_686 = $signed(_T_94761); // @[Modules.scala 56:109:@48049.4]
  assign _T_94763 = $signed(buffer_12_590) + $signed(buffer_12_591); // @[Modules.scala 56:109:@48051.4]
  assign _T_94764 = _T_94763[10:0]; // @[Modules.scala 56:109:@48052.4]
  assign buffer_12_687 = $signed(_T_94764); // @[Modules.scala 56:109:@48053.4]
  assign _T_94766 = $signed(buffer_1_592) + $signed(buffer_9_593); // @[Modules.scala 56:109:@48055.4]
  assign _T_94767 = _T_94766[10:0]; // @[Modules.scala 56:109:@48056.4]
  assign buffer_12_688 = $signed(_T_94767); // @[Modules.scala 56:109:@48057.4]
  assign _T_94769 = $signed(buffer_2_594) + $signed(buffer_12_595); // @[Modules.scala 56:109:@48059.4]
  assign _T_94770 = _T_94769[10:0]; // @[Modules.scala 56:109:@48060.4]
  assign buffer_12_689 = $signed(_T_94770); // @[Modules.scala 56:109:@48061.4]
  assign _T_94775 = $signed(buffer_12_598) + $signed(buffer_1_599); // @[Modules.scala 56:109:@48067.4]
  assign _T_94776 = _T_94775[10:0]; // @[Modules.scala 56:109:@48068.4]
  assign buffer_12_691 = $signed(_T_94776); // @[Modules.scala 56:109:@48069.4]
  assign _T_94778 = $signed(buffer_1_600) + $signed(buffer_12_601); // @[Modules.scala 56:109:@48071.4]
  assign _T_94779 = _T_94778[10:0]; // @[Modules.scala 56:109:@48072.4]
  assign buffer_12_692 = $signed(_T_94779); // @[Modules.scala 56:109:@48073.4]
  assign _T_94781 = $signed(buffer_12_602) + $signed(buffer_12_603); // @[Modules.scala 56:109:@48075.4]
  assign _T_94782 = _T_94781[10:0]; // @[Modules.scala 56:109:@48076.4]
  assign buffer_12_693 = $signed(_T_94782); // @[Modules.scala 56:109:@48077.4]
  assign _T_94784 = $signed(buffer_12_604) + $signed(buffer_12_605); // @[Modules.scala 56:109:@48079.4]
  assign _T_94785 = _T_94784[10:0]; // @[Modules.scala 56:109:@48080.4]
  assign buffer_12_694 = $signed(_T_94785); // @[Modules.scala 56:109:@48081.4]
  assign _T_94787 = $signed(buffer_12_606) + $signed(buffer_12_607); // @[Modules.scala 56:109:@48083.4]
  assign _T_94788 = _T_94787[10:0]; // @[Modules.scala 56:109:@48084.4]
  assign buffer_12_695 = $signed(_T_94788); // @[Modules.scala 56:109:@48085.4]
  assign _T_94790 = $signed(buffer_12_608) + $signed(buffer_0_609); // @[Modules.scala 56:109:@48087.4]
  assign _T_94791 = _T_94790[10:0]; // @[Modules.scala 56:109:@48088.4]
  assign buffer_12_696 = $signed(_T_94791); // @[Modules.scala 56:109:@48089.4]
  assign _T_94793 = $signed(buffer_12_610) + $signed(buffer_12_611); // @[Modules.scala 56:109:@48091.4]
  assign _T_94794 = _T_94793[10:0]; // @[Modules.scala 56:109:@48092.4]
  assign buffer_12_697 = $signed(_T_94794); // @[Modules.scala 56:109:@48093.4]
  assign _T_94796 = $signed(buffer_0_612) + $signed(buffer_12_613); // @[Modules.scala 56:109:@48095.4]
  assign _T_94797 = _T_94796[10:0]; // @[Modules.scala 56:109:@48096.4]
  assign buffer_12_698 = $signed(_T_94797); // @[Modules.scala 56:109:@48097.4]
  assign _T_94799 = $signed(buffer_12_614) + $signed(buffer_0_615); // @[Modules.scala 56:109:@48099.4]
  assign _T_94800 = _T_94799[10:0]; // @[Modules.scala 56:109:@48100.4]
  assign buffer_12_699 = $signed(_T_94800); // @[Modules.scala 56:109:@48101.4]
  assign _T_94802 = $signed(buffer_12_616) + $signed(buffer_12_617); // @[Modules.scala 56:109:@48103.4]
  assign _T_94803 = _T_94802[10:0]; // @[Modules.scala 56:109:@48104.4]
  assign buffer_12_700 = $signed(_T_94803); // @[Modules.scala 56:109:@48105.4]
  assign _T_94805 = $signed(buffer_12_618) + $signed(buffer_12_619); // @[Modules.scala 56:109:@48107.4]
  assign _T_94806 = _T_94805[10:0]; // @[Modules.scala 56:109:@48108.4]
  assign buffer_12_701 = $signed(_T_94806); // @[Modules.scala 56:109:@48109.4]
  assign _T_94808 = $signed(buffer_12_620) + $signed(buffer_12_621); // @[Modules.scala 56:109:@48111.4]
  assign _T_94809 = _T_94808[10:0]; // @[Modules.scala 56:109:@48112.4]
  assign buffer_12_702 = $signed(_T_94809); // @[Modules.scala 56:109:@48113.4]
  assign _T_94811 = $signed(buffer_6_622) + $signed(buffer_12_623); // @[Modules.scala 56:109:@48115.4]
  assign _T_94812 = _T_94811[10:0]; // @[Modules.scala 56:109:@48116.4]
  assign buffer_12_703 = $signed(_T_94812); // @[Modules.scala 56:109:@48117.4]
  assign _T_94814 = $signed(buffer_12_624) + $signed(buffer_12_625); // @[Modules.scala 56:109:@48119.4]
  assign _T_94815 = _T_94814[10:0]; // @[Modules.scala 56:109:@48120.4]
  assign buffer_12_704 = $signed(_T_94815); // @[Modules.scala 56:109:@48121.4]
  assign _T_94817 = $signed(buffer_12_626) + $signed(buffer_3_627); // @[Modules.scala 56:109:@48123.4]
  assign _T_94818 = _T_94817[10:0]; // @[Modules.scala 56:109:@48124.4]
  assign buffer_12_705 = $signed(_T_94818); // @[Modules.scala 56:109:@48125.4]
  assign _T_94820 = $signed(buffer_12_628) + $signed(buffer_12_629); // @[Modules.scala 56:109:@48127.4]
  assign _T_94821 = _T_94820[10:0]; // @[Modules.scala 56:109:@48128.4]
  assign buffer_12_706 = $signed(_T_94821); // @[Modules.scala 56:109:@48129.4]
  assign _T_94823 = $signed(buffer_12_630) + $signed(buffer_3_631); // @[Modules.scala 56:109:@48131.4]
  assign _T_94824 = _T_94823[10:0]; // @[Modules.scala 56:109:@48132.4]
  assign buffer_12_707 = $signed(_T_94824); // @[Modules.scala 56:109:@48133.4]
  assign _T_94826 = $signed(buffer_12_632) + $signed(buffer_12_633); // @[Modules.scala 56:109:@48135.4]
  assign _T_94827 = _T_94826[10:0]; // @[Modules.scala 56:109:@48136.4]
  assign buffer_12_708 = $signed(_T_94827); // @[Modules.scala 56:109:@48137.4]
  assign _T_94829 = $signed(buffer_9_634) + $signed(buffer_12_635); // @[Modules.scala 56:109:@48139.4]
  assign _T_94830 = _T_94829[10:0]; // @[Modules.scala 56:109:@48140.4]
  assign buffer_12_709 = $signed(_T_94830); // @[Modules.scala 56:109:@48141.4]
  assign _T_94832 = $signed(buffer_12_636) + $signed(buffer_12_637); // @[Modules.scala 56:109:@48143.4]
  assign _T_94833 = _T_94832[10:0]; // @[Modules.scala 56:109:@48144.4]
  assign buffer_12_710 = $signed(_T_94833); // @[Modules.scala 56:109:@48145.4]
  assign _T_94835 = $signed(buffer_12_638) + $signed(buffer_12_639); // @[Modules.scala 56:109:@48147.4]
  assign _T_94836 = _T_94835[10:0]; // @[Modules.scala 56:109:@48148.4]
  assign buffer_12_711 = $signed(_T_94836); // @[Modules.scala 56:109:@48149.4]
  assign _T_94838 = $signed(buffer_12_640) + $signed(buffer_0_641); // @[Modules.scala 56:109:@48151.4]
  assign _T_94839 = _T_94838[10:0]; // @[Modules.scala 56:109:@48152.4]
  assign buffer_12_712 = $signed(_T_94839); // @[Modules.scala 56:109:@48153.4]
  assign _T_94841 = $signed(buffer_1_642) + $signed(buffer_12_643); // @[Modules.scala 56:109:@48155.4]
  assign _T_94842 = _T_94841[10:0]; // @[Modules.scala 56:109:@48156.4]
  assign buffer_12_713 = $signed(_T_94842); // @[Modules.scala 56:109:@48157.4]
  assign _T_94844 = $signed(buffer_6_644) + $signed(buffer_12_645); // @[Modules.scala 56:109:@48159.4]
  assign _T_94845 = _T_94844[10:0]; // @[Modules.scala 56:109:@48160.4]
  assign buffer_12_714 = $signed(_T_94845); // @[Modules.scala 56:109:@48161.4]
  assign _T_94847 = $signed(buffer_12_646) + $signed(buffer_12_647); // @[Modules.scala 56:109:@48163.4]
  assign _T_94848 = _T_94847[10:0]; // @[Modules.scala 56:109:@48164.4]
  assign buffer_12_715 = $signed(_T_94848); // @[Modules.scala 56:109:@48165.4]
  assign _T_94850 = $signed(buffer_12_648) + $signed(buffer_12_649); // @[Modules.scala 56:109:@48167.4]
  assign _T_94851 = _T_94850[10:0]; // @[Modules.scala 56:109:@48168.4]
  assign buffer_12_716 = $signed(_T_94851); // @[Modules.scala 56:109:@48169.4]
  assign _T_94853 = $signed(buffer_3_650) + $signed(buffer_12_651); // @[Modules.scala 56:109:@48171.4]
  assign _T_94854 = _T_94853[10:0]; // @[Modules.scala 56:109:@48172.4]
  assign buffer_12_717 = $signed(_T_94854); // @[Modules.scala 56:109:@48173.4]
  assign _T_94856 = $signed(buffer_12_652) + $signed(buffer_12_653); // @[Modules.scala 56:109:@48175.4]
  assign _T_94857 = _T_94856[10:0]; // @[Modules.scala 56:109:@48176.4]
  assign buffer_12_718 = $signed(_T_94857); // @[Modules.scala 56:109:@48177.4]
  assign _T_94859 = $signed(buffer_12_654) + $signed(buffer_9_655); // @[Modules.scala 56:109:@48179.4]
  assign _T_94860 = _T_94859[10:0]; // @[Modules.scala 56:109:@48180.4]
  assign buffer_12_719 = $signed(_T_94860); // @[Modules.scala 56:109:@48181.4]
  assign _T_94862 = $signed(buffer_12_656) + $signed(buffer_3_657); // @[Modules.scala 56:109:@48183.4]
  assign _T_94863 = _T_94862[10:0]; // @[Modules.scala 56:109:@48184.4]
  assign buffer_12_720 = $signed(_T_94863); // @[Modules.scala 56:109:@48185.4]
  assign _T_94865 = $signed(buffer_12_658) + $signed(buffer_1_659); // @[Modules.scala 56:109:@48187.4]
  assign _T_94866 = _T_94865[10:0]; // @[Modules.scala 56:109:@48188.4]
  assign buffer_12_721 = $signed(_T_94866); // @[Modules.scala 56:109:@48189.4]
  assign _T_94868 = $signed(buffer_12_660) + $signed(buffer_12_661); // @[Modules.scala 56:109:@48191.4]
  assign _T_94869 = _T_94868[10:0]; // @[Modules.scala 56:109:@48192.4]
  assign buffer_12_722 = $signed(_T_94869); // @[Modules.scala 56:109:@48193.4]
  assign _T_94871 = $signed(buffer_12_662) + $signed(buffer_0_663); // @[Modules.scala 56:109:@48195.4]
  assign _T_94872 = _T_94871[10:0]; // @[Modules.scala 56:109:@48196.4]
  assign buffer_12_723 = $signed(_T_94872); // @[Modules.scala 56:109:@48197.4]
  assign _T_94874 = $signed(buffer_12_664) + $signed(buffer_12_665); // @[Modules.scala 56:109:@48199.4]
  assign _T_94875 = _T_94874[10:0]; // @[Modules.scala 56:109:@48200.4]
  assign buffer_12_724 = $signed(_T_94875); // @[Modules.scala 56:109:@48201.4]
  assign _T_94877 = $signed(buffer_12_666) + $signed(buffer_12_667); // @[Modules.scala 56:109:@48203.4]
  assign _T_94878 = _T_94877[10:0]; // @[Modules.scala 56:109:@48204.4]
  assign buffer_12_725 = $signed(_T_94878); // @[Modules.scala 56:109:@48205.4]
  assign _T_94880 = $signed(buffer_12_668) + $signed(buffer_12_669); // @[Modules.scala 56:109:@48207.4]
  assign _T_94881 = _T_94880[10:0]; // @[Modules.scala 56:109:@48208.4]
  assign buffer_12_726 = $signed(_T_94881); // @[Modules.scala 56:109:@48209.4]
  assign _T_94883 = $signed(buffer_6_670) + $signed(buffer_12_671); // @[Modules.scala 56:109:@48211.4]
  assign _T_94884 = _T_94883[10:0]; // @[Modules.scala 56:109:@48212.4]
  assign buffer_12_727 = $signed(_T_94884); // @[Modules.scala 56:109:@48213.4]
  assign _T_94886 = $signed(buffer_2_672) + $signed(buffer_12_673); // @[Modules.scala 56:109:@48215.4]
  assign _T_94887 = _T_94886[10:0]; // @[Modules.scala 56:109:@48216.4]
  assign buffer_12_728 = $signed(_T_94887); // @[Modules.scala 56:109:@48217.4]
  assign _T_94889 = $signed(buffer_3_674) + $signed(buffer_12_675); // @[Modules.scala 56:109:@48219.4]
  assign _T_94890 = _T_94889[10:0]; // @[Modules.scala 56:109:@48220.4]
  assign buffer_12_729 = $signed(_T_94890); // @[Modules.scala 56:109:@48221.4]
  assign _T_94895 = $signed(buffer_9_678) + $signed(buffer_12_679); // @[Modules.scala 56:109:@48227.4]
  assign _T_94896 = _T_94895[10:0]; // @[Modules.scala 56:109:@48228.4]
  assign buffer_12_731 = $signed(_T_94896); // @[Modules.scala 56:109:@48229.4]
  assign _T_94901 = $signed(buffer_12_682) + $signed(buffer_12_683); // @[Modules.scala 56:109:@48235.4]
  assign _T_94902 = _T_94901[10:0]; // @[Modules.scala 56:109:@48236.4]
  assign buffer_12_733 = $signed(_T_94902); // @[Modules.scala 56:109:@48237.4]
  assign _T_94904 = $signed(buffer_3_684) + $signed(buffer_12_685); // @[Modules.scala 56:109:@48239.4]
  assign _T_94905 = _T_94904[10:0]; // @[Modules.scala 56:109:@48240.4]
  assign buffer_12_734 = $signed(_T_94905); // @[Modules.scala 56:109:@48241.4]
  assign _T_94907 = $signed(buffer_12_686) + $signed(buffer_12_687); // @[Modules.scala 63:156:@48244.4]
  assign _T_94908 = _T_94907[10:0]; // @[Modules.scala 63:156:@48245.4]
  assign buffer_12_736 = $signed(_T_94908); // @[Modules.scala 63:156:@48246.4]
  assign _T_94910 = $signed(buffer_12_736) + $signed(buffer_12_688); // @[Modules.scala 63:156:@48248.4]
  assign _T_94911 = _T_94910[10:0]; // @[Modules.scala 63:156:@48249.4]
  assign buffer_12_737 = $signed(_T_94911); // @[Modules.scala 63:156:@48250.4]
  assign _T_94913 = $signed(buffer_12_737) + $signed(buffer_12_689); // @[Modules.scala 63:156:@48252.4]
  assign _T_94914 = _T_94913[10:0]; // @[Modules.scala 63:156:@48253.4]
  assign buffer_12_738 = $signed(_T_94914); // @[Modules.scala 63:156:@48254.4]
  assign _T_94916 = $signed(buffer_12_738) + $signed(buffer_1_690); // @[Modules.scala 63:156:@48256.4]
  assign _T_94917 = _T_94916[10:0]; // @[Modules.scala 63:156:@48257.4]
  assign buffer_12_739 = $signed(_T_94917); // @[Modules.scala 63:156:@48258.4]
  assign _T_94919 = $signed(buffer_12_739) + $signed(buffer_12_691); // @[Modules.scala 63:156:@48260.4]
  assign _T_94920 = _T_94919[10:0]; // @[Modules.scala 63:156:@48261.4]
  assign buffer_12_740 = $signed(_T_94920); // @[Modules.scala 63:156:@48262.4]
  assign _T_94922 = $signed(buffer_12_740) + $signed(buffer_12_692); // @[Modules.scala 63:156:@48264.4]
  assign _T_94923 = _T_94922[10:0]; // @[Modules.scala 63:156:@48265.4]
  assign buffer_12_741 = $signed(_T_94923); // @[Modules.scala 63:156:@48266.4]
  assign _T_94925 = $signed(buffer_12_741) + $signed(buffer_12_693); // @[Modules.scala 63:156:@48268.4]
  assign _T_94926 = _T_94925[10:0]; // @[Modules.scala 63:156:@48269.4]
  assign buffer_12_742 = $signed(_T_94926); // @[Modules.scala 63:156:@48270.4]
  assign _T_94928 = $signed(buffer_12_742) + $signed(buffer_12_694); // @[Modules.scala 63:156:@48272.4]
  assign _T_94929 = _T_94928[10:0]; // @[Modules.scala 63:156:@48273.4]
  assign buffer_12_743 = $signed(_T_94929); // @[Modules.scala 63:156:@48274.4]
  assign _T_94931 = $signed(buffer_12_743) + $signed(buffer_12_695); // @[Modules.scala 63:156:@48276.4]
  assign _T_94932 = _T_94931[10:0]; // @[Modules.scala 63:156:@48277.4]
  assign buffer_12_744 = $signed(_T_94932); // @[Modules.scala 63:156:@48278.4]
  assign _T_94934 = $signed(buffer_12_744) + $signed(buffer_12_696); // @[Modules.scala 63:156:@48280.4]
  assign _T_94935 = _T_94934[10:0]; // @[Modules.scala 63:156:@48281.4]
  assign buffer_12_745 = $signed(_T_94935); // @[Modules.scala 63:156:@48282.4]
  assign _T_94937 = $signed(buffer_12_745) + $signed(buffer_12_697); // @[Modules.scala 63:156:@48284.4]
  assign _T_94938 = _T_94937[10:0]; // @[Modules.scala 63:156:@48285.4]
  assign buffer_12_746 = $signed(_T_94938); // @[Modules.scala 63:156:@48286.4]
  assign _T_94940 = $signed(buffer_12_746) + $signed(buffer_12_698); // @[Modules.scala 63:156:@48288.4]
  assign _T_94941 = _T_94940[10:0]; // @[Modules.scala 63:156:@48289.4]
  assign buffer_12_747 = $signed(_T_94941); // @[Modules.scala 63:156:@48290.4]
  assign _T_94943 = $signed(buffer_12_747) + $signed(buffer_12_699); // @[Modules.scala 63:156:@48292.4]
  assign _T_94944 = _T_94943[10:0]; // @[Modules.scala 63:156:@48293.4]
  assign buffer_12_748 = $signed(_T_94944); // @[Modules.scala 63:156:@48294.4]
  assign _T_94946 = $signed(buffer_12_748) + $signed(buffer_12_700); // @[Modules.scala 63:156:@48296.4]
  assign _T_94947 = _T_94946[10:0]; // @[Modules.scala 63:156:@48297.4]
  assign buffer_12_749 = $signed(_T_94947); // @[Modules.scala 63:156:@48298.4]
  assign _T_94949 = $signed(buffer_12_749) + $signed(buffer_12_701); // @[Modules.scala 63:156:@48300.4]
  assign _T_94950 = _T_94949[10:0]; // @[Modules.scala 63:156:@48301.4]
  assign buffer_12_750 = $signed(_T_94950); // @[Modules.scala 63:156:@48302.4]
  assign _T_94952 = $signed(buffer_12_750) + $signed(buffer_12_702); // @[Modules.scala 63:156:@48304.4]
  assign _T_94953 = _T_94952[10:0]; // @[Modules.scala 63:156:@48305.4]
  assign buffer_12_751 = $signed(_T_94953); // @[Modules.scala 63:156:@48306.4]
  assign _T_94955 = $signed(buffer_12_751) + $signed(buffer_12_703); // @[Modules.scala 63:156:@48308.4]
  assign _T_94956 = _T_94955[10:0]; // @[Modules.scala 63:156:@48309.4]
  assign buffer_12_752 = $signed(_T_94956); // @[Modules.scala 63:156:@48310.4]
  assign _T_94958 = $signed(buffer_12_752) + $signed(buffer_12_704); // @[Modules.scala 63:156:@48312.4]
  assign _T_94959 = _T_94958[10:0]; // @[Modules.scala 63:156:@48313.4]
  assign buffer_12_753 = $signed(_T_94959); // @[Modules.scala 63:156:@48314.4]
  assign _T_94961 = $signed(buffer_12_753) + $signed(buffer_12_705); // @[Modules.scala 63:156:@48316.4]
  assign _T_94962 = _T_94961[10:0]; // @[Modules.scala 63:156:@48317.4]
  assign buffer_12_754 = $signed(_T_94962); // @[Modules.scala 63:156:@48318.4]
  assign _T_94964 = $signed(buffer_12_754) + $signed(buffer_12_706); // @[Modules.scala 63:156:@48320.4]
  assign _T_94965 = _T_94964[10:0]; // @[Modules.scala 63:156:@48321.4]
  assign buffer_12_755 = $signed(_T_94965); // @[Modules.scala 63:156:@48322.4]
  assign _T_94967 = $signed(buffer_12_755) + $signed(buffer_12_707); // @[Modules.scala 63:156:@48324.4]
  assign _T_94968 = _T_94967[10:0]; // @[Modules.scala 63:156:@48325.4]
  assign buffer_12_756 = $signed(_T_94968); // @[Modules.scala 63:156:@48326.4]
  assign _T_94970 = $signed(buffer_12_756) + $signed(buffer_12_708); // @[Modules.scala 63:156:@48328.4]
  assign _T_94971 = _T_94970[10:0]; // @[Modules.scala 63:156:@48329.4]
  assign buffer_12_757 = $signed(_T_94971); // @[Modules.scala 63:156:@48330.4]
  assign _T_94973 = $signed(buffer_12_757) + $signed(buffer_12_709); // @[Modules.scala 63:156:@48332.4]
  assign _T_94974 = _T_94973[10:0]; // @[Modules.scala 63:156:@48333.4]
  assign buffer_12_758 = $signed(_T_94974); // @[Modules.scala 63:156:@48334.4]
  assign _T_94976 = $signed(buffer_12_758) + $signed(buffer_12_710); // @[Modules.scala 63:156:@48336.4]
  assign _T_94977 = _T_94976[10:0]; // @[Modules.scala 63:156:@48337.4]
  assign buffer_12_759 = $signed(_T_94977); // @[Modules.scala 63:156:@48338.4]
  assign _T_94979 = $signed(buffer_12_759) + $signed(buffer_12_711); // @[Modules.scala 63:156:@48340.4]
  assign _T_94980 = _T_94979[10:0]; // @[Modules.scala 63:156:@48341.4]
  assign buffer_12_760 = $signed(_T_94980); // @[Modules.scala 63:156:@48342.4]
  assign _T_94982 = $signed(buffer_12_760) + $signed(buffer_12_712); // @[Modules.scala 63:156:@48344.4]
  assign _T_94983 = _T_94982[10:0]; // @[Modules.scala 63:156:@48345.4]
  assign buffer_12_761 = $signed(_T_94983); // @[Modules.scala 63:156:@48346.4]
  assign _T_94985 = $signed(buffer_12_761) + $signed(buffer_12_713); // @[Modules.scala 63:156:@48348.4]
  assign _T_94986 = _T_94985[10:0]; // @[Modules.scala 63:156:@48349.4]
  assign buffer_12_762 = $signed(_T_94986); // @[Modules.scala 63:156:@48350.4]
  assign _T_94988 = $signed(buffer_12_762) + $signed(buffer_12_714); // @[Modules.scala 63:156:@48352.4]
  assign _T_94989 = _T_94988[10:0]; // @[Modules.scala 63:156:@48353.4]
  assign buffer_12_763 = $signed(_T_94989); // @[Modules.scala 63:156:@48354.4]
  assign _T_94991 = $signed(buffer_12_763) + $signed(buffer_12_715); // @[Modules.scala 63:156:@48356.4]
  assign _T_94992 = _T_94991[10:0]; // @[Modules.scala 63:156:@48357.4]
  assign buffer_12_764 = $signed(_T_94992); // @[Modules.scala 63:156:@48358.4]
  assign _T_94994 = $signed(buffer_12_764) + $signed(buffer_12_716); // @[Modules.scala 63:156:@48360.4]
  assign _T_94995 = _T_94994[10:0]; // @[Modules.scala 63:156:@48361.4]
  assign buffer_12_765 = $signed(_T_94995); // @[Modules.scala 63:156:@48362.4]
  assign _T_94997 = $signed(buffer_12_765) + $signed(buffer_12_717); // @[Modules.scala 63:156:@48364.4]
  assign _T_94998 = _T_94997[10:0]; // @[Modules.scala 63:156:@48365.4]
  assign buffer_12_766 = $signed(_T_94998); // @[Modules.scala 63:156:@48366.4]
  assign _T_95000 = $signed(buffer_12_766) + $signed(buffer_12_718); // @[Modules.scala 63:156:@48368.4]
  assign _T_95001 = _T_95000[10:0]; // @[Modules.scala 63:156:@48369.4]
  assign buffer_12_767 = $signed(_T_95001); // @[Modules.scala 63:156:@48370.4]
  assign _T_95003 = $signed(buffer_12_767) + $signed(buffer_12_719); // @[Modules.scala 63:156:@48372.4]
  assign _T_95004 = _T_95003[10:0]; // @[Modules.scala 63:156:@48373.4]
  assign buffer_12_768 = $signed(_T_95004); // @[Modules.scala 63:156:@48374.4]
  assign _T_95006 = $signed(buffer_12_768) + $signed(buffer_12_720); // @[Modules.scala 63:156:@48376.4]
  assign _T_95007 = _T_95006[10:0]; // @[Modules.scala 63:156:@48377.4]
  assign buffer_12_769 = $signed(_T_95007); // @[Modules.scala 63:156:@48378.4]
  assign _T_95009 = $signed(buffer_12_769) + $signed(buffer_12_721); // @[Modules.scala 63:156:@48380.4]
  assign _T_95010 = _T_95009[10:0]; // @[Modules.scala 63:156:@48381.4]
  assign buffer_12_770 = $signed(_T_95010); // @[Modules.scala 63:156:@48382.4]
  assign _T_95012 = $signed(buffer_12_770) + $signed(buffer_12_722); // @[Modules.scala 63:156:@48384.4]
  assign _T_95013 = _T_95012[10:0]; // @[Modules.scala 63:156:@48385.4]
  assign buffer_12_771 = $signed(_T_95013); // @[Modules.scala 63:156:@48386.4]
  assign _T_95015 = $signed(buffer_12_771) + $signed(buffer_12_723); // @[Modules.scala 63:156:@48388.4]
  assign _T_95016 = _T_95015[10:0]; // @[Modules.scala 63:156:@48389.4]
  assign buffer_12_772 = $signed(_T_95016); // @[Modules.scala 63:156:@48390.4]
  assign _T_95018 = $signed(buffer_12_772) + $signed(buffer_12_724); // @[Modules.scala 63:156:@48392.4]
  assign _T_95019 = _T_95018[10:0]; // @[Modules.scala 63:156:@48393.4]
  assign buffer_12_773 = $signed(_T_95019); // @[Modules.scala 63:156:@48394.4]
  assign _T_95021 = $signed(buffer_12_773) + $signed(buffer_12_725); // @[Modules.scala 63:156:@48396.4]
  assign _T_95022 = _T_95021[10:0]; // @[Modules.scala 63:156:@48397.4]
  assign buffer_12_774 = $signed(_T_95022); // @[Modules.scala 63:156:@48398.4]
  assign _T_95024 = $signed(buffer_12_774) + $signed(buffer_12_726); // @[Modules.scala 63:156:@48400.4]
  assign _T_95025 = _T_95024[10:0]; // @[Modules.scala 63:156:@48401.4]
  assign buffer_12_775 = $signed(_T_95025); // @[Modules.scala 63:156:@48402.4]
  assign _T_95027 = $signed(buffer_12_775) + $signed(buffer_12_727); // @[Modules.scala 63:156:@48404.4]
  assign _T_95028 = _T_95027[10:0]; // @[Modules.scala 63:156:@48405.4]
  assign buffer_12_776 = $signed(_T_95028); // @[Modules.scala 63:156:@48406.4]
  assign _T_95030 = $signed(buffer_12_776) + $signed(buffer_12_728); // @[Modules.scala 63:156:@48408.4]
  assign _T_95031 = _T_95030[10:0]; // @[Modules.scala 63:156:@48409.4]
  assign buffer_12_777 = $signed(_T_95031); // @[Modules.scala 63:156:@48410.4]
  assign _T_95033 = $signed(buffer_12_777) + $signed(buffer_12_729); // @[Modules.scala 63:156:@48412.4]
  assign _T_95034 = _T_95033[10:0]; // @[Modules.scala 63:156:@48413.4]
  assign buffer_12_778 = $signed(_T_95034); // @[Modules.scala 63:156:@48414.4]
  assign _T_95036 = $signed(buffer_12_778) + $signed(buffer_2_730); // @[Modules.scala 63:156:@48416.4]
  assign _T_95037 = _T_95036[10:0]; // @[Modules.scala 63:156:@48417.4]
  assign buffer_12_779 = $signed(_T_95037); // @[Modules.scala 63:156:@48418.4]
  assign _T_95039 = $signed(buffer_12_779) + $signed(buffer_12_731); // @[Modules.scala 63:156:@48420.4]
  assign _T_95040 = _T_95039[10:0]; // @[Modules.scala 63:156:@48421.4]
  assign buffer_12_780 = $signed(_T_95040); // @[Modules.scala 63:156:@48422.4]
  assign _T_95042 = $signed(buffer_12_780) + $signed(buffer_4_732); // @[Modules.scala 63:156:@48424.4]
  assign _T_95043 = _T_95042[10:0]; // @[Modules.scala 63:156:@48425.4]
  assign buffer_12_781 = $signed(_T_95043); // @[Modules.scala 63:156:@48426.4]
  assign _T_95045 = $signed(buffer_12_781) + $signed(buffer_12_733); // @[Modules.scala 63:156:@48428.4]
  assign _T_95046 = _T_95045[10:0]; // @[Modules.scala 63:156:@48429.4]
  assign buffer_12_782 = $signed(_T_95046); // @[Modules.scala 63:156:@48430.4]
  assign _T_95048 = $signed(buffer_12_782) + $signed(buffer_12_734); // @[Modules.scala 63:156:@48432.4]
  assign _T_95049 = _T_95048[10:0]; // @[Modules.scala 63:156:@48433.4]
  assign buffer_12_783 = $signed(_T_95049); // @[Modules.scala 63:156:@48434.4]
  assign _T_95085 = $signed(io_in_12) - $signed(io_in_13); // @[Modules.scala 40:46:@48473.4]
  assign _T_95086 = _T_95085[4:0]; // @[Modules.scala 40:46:@48474.4]
  assign _T_95087 = $signed(_T_95086); // @[Modules.scala 40:46:@48475.4]
  assign _T_95149 = $signed(io_in_36) - $signed(io_in_37); // @[Modules.scala 40:46:@48542.4]
  assign _T_95150 = _T_95149[4:0]; // @[Modules.scala 40:46:@48543.4]
  assign _T_95151 = $signed(_T_95150); // @[Modules.scala 40:46:@48544.4]
  assign _T_95236 = $signed(io_in_70) - $signed(io_in_71); // @[Modules.scala 40:46:@48637.4]
  assign _T_95237 = _T_95236[4:0]; // @[Modules.scala 40:46:@48638.4]
  assign _T_95238 = $signed(_T_95237); // @[Modules.scala 40:46:@48639.4]
  assign _T_95255 = $signed(io_in_80) - $signed(io_in_81); // @[Modules.scala 40:46:@48660.4]
  assign _T_95256 = _T_95255[4:0]; // @[Modules.scala 40:46:@48661.4]
  assign _T_95257 = $signed(_T_95256); // @[Modules.scala 40:46:@48662.4]
  assign _T_95448 = $signed(io_in_158) - $signed(io_in_159); // @[Modules.scala 40:46:@48873.4]
  assign _T_95449 = _T_95448[4:0]; // @[Modules.scala 40:46:@48874.4]
  assign _T_95450 = $signed(_T_95449); // @[Modules.scala 40:46:@48875.4]
  assign _T_95482 = $signed(io_in_170) - $signed(io_in_171); // @[Modules.scala 40:46:@48909.4]
  assign _T_95483 = _T_95482[4:0]; // @[Modules.scala 40:46:@48910.4]
  assign _T_95484 = $signed(_T_95483); // @[Modules.scala 40:46:@48911.4]
  assign _T_95513 = $signed(io_in_180) - $signed(io_in_181); // @[Modules.scala 40:46:@48941.4]
  assign _T_95514 = _T_95513[4:0]; // @[Modules.scala 40:46:@48942.4]
  assign _T_95515 = $signed(_T_95514); // @[Modules.scala 40:46:@48943.4]
  assign _T_95530 = $signed(_T_61118) + $signed(io_in_187); // @[Modules.scala 43:47:@48959.4]
  assign _T_95531 = _T_95530[4:0]; // @[Modules.scala 43:47:@48960.4]
  assign _T_95532 = $signed(_T_95531); // @[Modules.scala 43:47:@48961.4]
  assign _T_95671 = $signed(io_in_240) - $signed(io_in_241); // @[Modules.scala 40:46:@49112.4]
  assign _T_95672 = _T_95671[4:0]; // @[Modules.scala 40:46:@49113.4]
  assign _T_95673 = $signed(_T_95672); // @[Modules.scala 40:46:@49114.4]
  assign _T_95747 = $signed(io_in_264) - $signed(io_in_265); // @[Modules.scala 40:46:@49190.4]
  assign _T_95748 = _T_95747[4:0]; // @[Modules.scala 40:46:@49191.4]
  assign _T_95749 = $signed(_T_95748); // @[Modules.scala 40:46:@49192.4]
  assign _T_95822 = $signed(_T_55124) + $signed(io_in_291); // @[Modules.scala 43:47:@49269.4]
  assign _T_95823 = _T_95822[4:0]; // @[Modules.scala 43:47:@49270.4]
  assign _T_95824 = $signed(_T_95823); // @[Modules.scala 43:47:@49271.4]
  assign _T_95889 = $signed(io_in_316) - $signed(io_in_317); // @[Modules.scala 40:46:@49342.4]
  assign _T_95890 = _T_95889[4:0]; // @[Modules.scala 40:46:@49343.4]
  assign _T_95891 = $signed(_T_95890); // @[Modules.scala 40:46:@49344.4]
  assign _T_95952 = $signed(io_in_342) - $signed(io_in_343); // @[Modules.scala 40:46:@49412.4]
  assign _T_95953 = _T_95952[4:0]; // @[Modules.scala 40:46:@49413.4]
  assign _T_95954 = $signed(_T_95953); // @[Modules.scala 40:46:@49414.4]
  assign _T_95959 = $signed(_T_64688) + $signed(io_in_345); // @[Modules.scala 43:47:@49419.4]
  assign _T_95960 = _T_95959[4:0]; // @[Modules.scala 43:47:@49420.4]
  assign _T_95961 = $signed(_T_95960); // @[Modules.scala 43:47:@49421.4]
  assign _T_95969 = $signed(io_in_348) - $signed(io_in_349); // @[Modules.scala 40:46:@49430.4]
  assign _T_95970 = _T_95969[4:0]; // @[Modules.scala 40:46:@49431.4]
  assign _T_95971 = $signed(_T_95970); // @[Modules.scala 40:46:@49432.4]
  assign _T_95983 = $signed(_T_58410) + $signed(io_in_353); // @[Modules.scala 43:47:@49444.4]
  assign _T_95984 = _T_95983[4:0]; // @[Modules.scala 43:47:@49445.4]
  assign _T_95985 = $signed(_T_95984); // @[Modules.scala 43:47:@49446.4]
  assign _T_96303 = $signed(io_in_496) - $signed(io_in_497); // @[Modules.scala 40:46:@49810.4]
  assign _T_96304 = _T_96303[4:0]; // @[Modules.scala 40:46:@49811.4]
  assign _T_96305 = $signed(_T_96304); // @[Modules.scala 40:46:@49812.4]
  assign _T_96378 = $signed(io_in_530) - $signed(io_in_531); // @[Modules.scala 40:46:@49896.4]
  assign _T_96379 = _T_96378[4:0]; // @[Modules.scala 40:46:@49897.4]
  assign _T_96380 = $signed(_T_96379); // @[Modules.scala 40:46:@49898.4]
  assign _T_96461 = $signed(_T_55807) + $signed(io_in_565); // @[Modules.scala 43:47:@49988.4]
  assign _T_96462 = _T_96461[4:0]; // @[Modules.scala 43:47:@49989.4]
  assign _T_96463 = $signed(_T_96462); // @[Modules.scala 43:47:@49990.4]
  assign _T_96602 = $signed(io_in_618) - $signed(io_in_619); // @[Modules.scala 40:46:@50141.4]
  assign _T_96603 = _T_96602[4:0]; // @[Modules.scala 40:46:@50142.4]
  assign _T_96604 = $signed(_T_96603); // @[Modules.scala 40:46:@50143.4]
  assign _T_96654 = $signed(_T_56036) - $signed(io_in_643); // @[Modules.scala 46:47:@50201.4]
  assign _T_96655 = _T_96654[4:0]; // @[Modules.scala 46:47:@50202.4]
  assign _T_96656 = $signed(_T_96655); // @[Modules.scala 46:47:@50203.4]
  assign _T_96706 = $signed(_T_56088) + $signed(io_in_659); // @[Modules.scala 43:47:@50254.4]
  assign _T_96707 = _T_96706[4:0]; // @[Modules.scala 43:47:@50255.4]
  assign _T_96708 = $signed(_T_96707); // @[Modules.scala 43:47:@50256.4]
  assign _T_97076 = $signed(io_in_782) - $signed(io_in_783); // @[Modules.scala 40:46:@50640.4]
  assign _T_97077 = _T_97076[4:0]; // @[Modules.scala 40:46:@50641.4]
  assign _T_97078 = $signed(_T_97077); // @[Modules.scala 40:46:@50642.4]
  assign _T_97079 = $signed(buffer_7_0) + $signed(buffer_3_1); // @[Modules.scala 50:57:@50644.4]
  assign _T_97080 = _T_97079[10:0]; // @[Modules.scala 50:57:@50645.4]
  assign buffer_13_392 = $signed(_T_97080); // @[Modules.scala 50:57:@50646.4]
  assign buffer_13_6 = {{6{_T_95087[4]}},_T_95087}; // @[Modules.scala 32:22:@8.4]
  assign _T_97088 = $signed(buffer_13_6) + $signed(buffer_0_7); // @[Modules.scala 50:57:@50656.4]
  assign _T_97089 = _T_97088[10:0]; // @[Modules.scala 50:57:@50657.4]
  assign buffer_13_395 = $signed(_T_97089); // @[Modules.scala 50:57:@50658.4]
  assign _T_97097 = $signed(buffer_2_12) + $signed(buffer_1_13); // @[Modules.scala 50:57:@50668.4]
  assign _T_97098 = _T_97097[10:0]; // @[Modules.scala 50:57:@50669.4]
  assign buffer_13_398 = $signed(_T_97098); // @[Modules.scala 50:57:@50670.4]
  assign _T_97100 = $signed(buffer_4_14) + $signed(buffer_0_15); // @[Modules.scala 50:57:@50672.4]
  assign _T_97101 = _T_97100[10:0]; // @[Modules.scala 50:57:@50673.4]
  assign buffer_13_399 = $signed(_T_97101); // @[Modules.scala 50:57:@50674.4]
  assign buffer_13_18 = {{6{_T_95151[4]}},_T_95151}; // @[Modules.scala 32:22:@8.4]
  assign _T_97106 = $signed(buffer_13_18) + $signed(buffer_0_19); // @[Modules.scala 50:57:@50680.4]
  assign _T_97107 = _T_97106[10:0]; // @[Modules.scala 50:57:@50681.4]
  assign buffer_13_401 = $signed(_T_97107); // @[Modules.scala 50:57:@50682.4]
  assign _T_97118 = $signed(buffer_1_26) + $signed(buffer_3_27); // @[Modules.scala 50:57:@50696.4]
  assign _T_97119 = _T_97118[10:0]; // @[Modules.scala 50:57:@50697.4]
  assign buffer_13_405 = $signed(_T_97119); // @[Modules.scala 50:57:@50698.4]
  assign buffer_13_35 = {{6{_T_95238[4]}},_T_95238}; // @[Modules.scala 32:22:@8.4]
  assign _T_97130 = $signed(buffer_1_34) + $signed(buffer_13_35); // @[Modules.scala 50:57:@50712.4]
  assign _T_97131 = _T_97130[10:0]; // @[Modules.scala 50:57:@50713.4]
  assign buffer_13_409 = $signed(_T_97131); // @[Modules.scala 50:57:@50714.4]
  assign _T_97133 = $signed(buffer_5_36) + $signed(buffer_1_37); // @[Modules.scala 50:57:@50716.4]
  assign _T_97134 = _T_97133[10:0]; // @[Modules.scala 50:57:@50717.4]
  assign buffer_13_410 = $signed(_T_97134); // @[Modules.scala 50:57:@50718.4]
  assign buffer_13_40 = {{6{_T_95257[4]}},_T_95257}; // @[Modules.scala 32:22:@8.4]
  assign _T_97139 = $signed(buffer_13_40) + $signed(buffer_0_41); // @[Modules.scala 50:57:@50724.4]
  assign _T_97140 = _T_97139[10:0]; // @[Modules.scala 50:57:@50725.4]
  assign buffer_13_412 = $signed(_T_97140); // @[Modules.scala 50:57:@50726.4]
  assign _T_97151 = $signed(buffer_1_48) + $signed(buffer_2_49); // @[Modules.scala 50:57:@50740.4]
  assign _T_97152 = _T_97151[10:0]; // @[Modules.scala 50:57:@50741.4]
  assign buffer_13_416 = $signed(_T_97152); // @[Modules.scala 50:57:@50742.4]
  assign _T_97169 = $signed(buffer_8_60) + $signed(buffer_4_61); // @[Modules.scala 50:57:@50764.4]
  assign _T_97170 = _T_97169[10:0]; // @[Modules.scala 50:57:@50765.4]
  assign buffer_13_422 = $signed(_T_97170); // @[Modules.scala 50:57:@50766.4]
  assign buffer_13_79 = {{6{_T_95450[4]}},_T_95450}; // @[Modules.scala 32:22:@8.4]
  assign _T_97196 = $signed(buffer_4_78) + $signed(buffer_13_79); // @[Modules.scala 50:57:@50800.4]
  assign _T_97197 = _T_97196[10:0]; // @[Modules.scala 50:57:@50801.4]
  assign buffer_13_431 = $signed(_T_97197); // @[Modules.scala 50:57:@50802.4]
  assign _T_97199 = $signed(buffer_4_80) + $signed(buffer_5_81); // @[Modules.scala 50:57:@50804.4]
  assign _T_97200 = _T_97199[10:0]; // @[Modules.scala 50:57:@50805.4]
  assign buffer_13_432 = $signed(_T_97200); // @[Modules.scala 50:57:@50806.4]
  assign buffer_13_85 = {{6{_T_95484[4]}},_T_95484}; // @[Modules.scala 32:22:@8.4]
  assign _T_97205 = $signed(buffer_0_84) + $signed(buffer_13_85); // @[Modules.scala 50:57:@50812.4]
  assign _T_97206 = _T_97205[10:0]; // @[Modules.scala 50:57:@50813.4]
  assign buffer_13_434 = $signed(_T_97206); // @[Modules.scala 50:57:@50814.4]
  assign buffer_13_90 = {{6{_T_95515[4]}},_T_95515}; // @[Modules.scala 32:22:@8.4]
  assign _T_97214 = $signed(buffer_13_90) + $signed(buffer_9_91); // @[Modules.scala 50:57:@50824.4]
  assign _T_97215 = _T_97214[10:0]; // @[Modules.scala 50:57:@50825.4]
  assign buffer_13_437 = $signed(_T_97215); // @[Modules.scala 50:57:@50826.4]
  assign buffer_13_93 = {{6{_T_95532[4]}},_T_95532}; // @[Modules.scala 32:22:@8.4]
  assign _T_97217 = $signed(buffer_5_92) + $signed(buffer_13_93); // @[Modules.scala 50:57:@50828.4]
  assign _T_97218 = _T_97217[10:0]; // @[Modules.scala 50:57:@50829.4]
  assign buffer_13_438 = $signed(_T_97218); // @[Modules.scala 50:57:@50830.4]
  assign _T_97220 = $signed(buffer_4_94) + $signed(buffer_0_95); // @[Modules.scala 50:57:@50832.4]
  assign _T_97221 = _T_97220[10:0]; // @[Modules.scala 50:57:@50833.4]
  assign buffer_13_439 = $signed(_T_97221); // @[Modules.scala 50:57:@50834.4]
  assign _T_97226 = $signed(buffer_6_98) + $signed(buffer_0_99); // @[Modules.scala 50:57:@50840.4]
  assign _T_97227 = _T_97226[10:0]; // @[Modules.scala 50:57:@50841.4]
  assign buffer_13_441 = $signed(_T_97227); // @[Modules.scala 50:57:@50842.4]
  assign _T_97229 = $signed(buffer_10_100) + $signed(buffer_0_101); // @[Modules.scala 50:57:@50844.4]
  assign _T_97230 = _T_97229[10:0]; // @[Modules.scala 50:57:@50845.4]
  assign buffer_13_442 = $signed(_T_97230); // @[Modules.scala 50:57:@50846.4]
  assign _T_97235 = $signed(buffer_2_104) + $signed(buffer_11_105); // @[Modules.scala 50:57:@50852.4]
  assign _T_97236 = _T_97235[10:0]; // @[Modules.scala 50:57:@50853.4]
  assign buffer_13_444 = $signed(_T_97236); // @[Modules.scala 50:57:@50854.4]
  assign _T_97247 = $signed(buffer_0_112) + $signed(buffer_12_113); // @[Modules.scala 50:57:@50868.4]
  assign _T_97248 = _T_97247[10:0]; // @[Modules.scala 50:57:@50869.4]
  assign buffer_13_448 = $signed(_T_97248); // @[Modules.scala 50:57:@50870.4]
  assign _T_97250 = $signed(buffer_0_114) + $signed(buffer_5_115); // @[Modules.scala 50:57:@50872.4]
  assign _T_97251 = _T_97250[10:0]; // @[Modules.scala 50:57:@50873.4]
  assign buffer_13_449 = $signed(_T_97251); // @[Modules.scala 50:57:@50874.4]
  assign buffer_13_120 = {{6{_T_95673[4]}},_T_95673}; // @[Modules.scala 32:22:@8.4]
  assign _T_97259 = $signed(buffer_13_120) + $signed(buffer_4_121); // @[Modules.scala 50:57:@50884.4]
  assign _T_97260 = _T_97259[10:0]; // @[Modules.scala 50:57:@50885.4]
  assign buffer_13_452 = $signed(_T_97260); // @[Modules.scala 50:57:@50886.4]
  assign _T_97274 = $signed(buffer_2_130) + $signed(buffer_0_131); // @[Modules.scala 50:57:@50904.4]
  assign _T_97275 = _T_97274[10:0]; // @[Modules.scala 50:57:@50905.4]
  assign buffer_13_457 = $signed(_T_97275); // @[Modules.scala 50:57:@50906.4]
  assign buffer_13_132 = {{6{_T_95749[4]}},_T_95749}; // @[Modules.scala 32:22:@8.4]
  assign _T_97277 = $signed(buffer_13_132) + $signed(buffer_0_133); // @[Modules.scala 50:57:@50908.4]
  assign _T_97278 = _T_97277[10:0]; // @[Modules.scala 50:57:@50909.4]
  assign buffer_13_458 = $signed(_T_97278); // @[Modules.scala 50:57:@50910.4]
  assign _T_97283 = $signed(buffer_0_136) + $signed(buffer_3_137); // @[Modules.scala 50:57:@50916.4]
  assign _T_97284 = _T_97283[10:0]; // @[Modules.scala 50:57:@50917.4]
  assign buffer_13_460 = $signed(_T_97284); // @[Modules.scala 50:57:@50918.4]
  assign buffer_13_145 = {{6{_T_95824[4]}},_T_95824}; // @[Modules.scala 32:22:@8.4]
  assign _T_97295 = $signed(buffer_2_144) + $signed(buffer_13_145); // @[Modules.scala 50:57:@50932.4]
  assign _T_97296 = _T_97295[10:0]; // @[Modules.scala 50:57:@50933.4]
  assign buffer_13_464 = $signed(_T_97296); // @[Modules.scala 50:57:@50934.4]
  assign _T_97301 = $signed(buffer_4_148) + $signed(buffer_3_149); // @[Modules.scala 50:57:@50940.4]
  assign _T_97302 = _T_97301[10:0]; // @[Modules.scala 50:57:@50941.4]
  assign buffer_13_466 = $signed(_T_97302); // @[Modules.scala 50:57:@50942.4]
  assign _T_97304 = $signed(buffer_5_150) + $signed(buffer_4_151); // @[Modules.scala 50:57:@50944.4]
  assign _T_97305 = _T_97304[10:0]; // @[Modules.scala 50:57:@50945.4]
  assign buffer_13_467 = $signed(_T_97305); // @[Modules.scala 50:57:@50946.4]
  assign _T_97313 = $signed(buffer_6_156) + $signed(buffer_1_157); // @[Modules.scala 50:57:@50956.4]
  assign _T_97314 = _T_97313[10:0]; // @[Modules.scala 50:57:@50957.4]
  assign buffer_13_470 = $signed(_T_97314); // @[Modules.scala 50:57:@50958.4]
  assign buffer_13_158 = {{6{_T_95891[4]}},_T_95891}; // @[Modules.scala 32:22:@8.4]
  assign _T_97316 = $signed(buffer_13_158) + $signed(buffer_0_159); // @[Modules.scala 50:57:@50960.4]
  assign _T_97317 = _T_97316[10:0]; // @[Modules.scala 50:57:@50961.4]
  assign buffer_13_471 = $signed(_T_97317); // @[Modules.scala 50:57:@50962.4]
  assign _T_97322 = $signed(buffer_1_162) + $signed(buffer_5_163); // @[Modules.scala 50:57:@50968.4]
  assign _T_97323 = _T_97322[10:0]; // @[Modules.scala 50:57:@50969.4]
  assign buffer_13_473 = $signed(_T_97323); // @[Modules.scala 50:57:@50970.4]
  assign _T_97331 = $signed(buffer_3_168) + $signed(buffer_0_169); // @[Modules.scala 50:57:@50980.4]
  assign _T_97332 = _T_97331[10:0]; // @[Modules.scala 50:57:@50981.4]
  assign buffer_13_476 = $signed(_T_97332); // @[Modules.scala 50:57:@50982.4]
  assign buffer_13_171 = {{6{_T_95954[4]}},_T_95954}; // @[Modules.scala 32:22:@8.4]
  assign _T_97334 = $signed(buffer_0_170) + $signed(buffer_13_171); // @[Modules.scala 50:57:@50984.4]
  assign _T_97335 = _T_97334[10:0]; // @[Modules.scala 50:57:@50985.4]
  assign buffer_13_477 = $signed(_T_97335); // @[Modules.scala 50:57:@50986.4]
  assign buffer_13_172 = {{6{_T_95961[4]}},_T_95961}; // @[Modules.scala 32:22:@8.4]
  assign _T_97337 = $signed(buffer_13_172) + $signed(buffer_3_173); // @[Modules.scala 50:57:@50988.4]
  assign _T_97338 = _T_97337[10:0]; // @[Modules.scala 50:57:@50989.4]
  assign buffer_13_478 = $signed(_T_97338); // @[Modules.scala 50:57:@50990.4]
  assign buffer_13_174 = {{6{_T_95971[4]}},_T_95971}; // @[Modules.scala 32:22:@8.4]
  assign _T_97340 = $signed(buffer_13_174) + $signed(buffer_1_175); // @[Modules.scala 50:57:@50992.4]
  assign _T_97341 = _T_97340[10:0]; // @[Modules.scala 50:57:@50993.4]
  assign buffer_13_479 = $signed(_T_97341); // @[Modules.scala 50:57:@50994.4]
  assign buffer_13_176 = {{6{_T_95985[4]}},_T_95985}; // @[Modules.scala 32:22:@8.4]
  assign _T_97343 = $signed(buffer_13_176) + $signed(buffer_5_177); // @[Modules.scala 50:57:@50996.4]
  assign _T_97344 = _T_97343[10:0]; // @[Modules.scala 50:57:@50997.4]
  assign buffer_13_480 = $signed(_T_97344); // @[Modules.scala 50:57:@50998.4]
  assign _T_97352 = $signed(buffer_7_182) + $signed(buffer_0_183); // @[Modules.scala 50:57:@51008.4]
  assign _T_97353 = _T_97352[10:0]; // @[Modules.scala 50:57:@51009.4]
  assign buffer_13_483 = $signed(_T_97353); // @[Modules.scala 50:57:@51010.4]
  assign _T_97358 = $signed(buffer_3_186) + $signed(buffer_0_187); // @[Modules.scala 50:57:@51016.4]
  assign _T_97359 = _T_97358[10:0]; // @[Modules.scala 50:57:@51017.4]
  assign buffer_13_485 = $signed(_T_97359); // @[Modules.scala 50:57:@51018.4]
  assign _T_97364 = $signed(buffer_4_190) + $signed(buffer_0_191); // @[Modules.scala 50:57:@51024.4]
  assign _T_97365 = _T_97364[10:0]; // @[Modules.scala 50:57:@51025.4]
  assign buffer_13_487 = $signed(_T_97365); // @[Modules.scala 50:57:@51026.4]
  assign _T_97367 = $signed(buffer_2_192) + $signed(buffer_0_193); // @[Modules.scala 50:57:@51028.4]
  assign _T_97368 = _T_97367[10:0]; // @[Modules.scala 50:57:@51029.4]
  assign buffer_13_488 = $signed(_T_97368); // @[Modules.scala 50:57:@51030.4]
  assign _T_97382 = $signed(buffer_1_202) + $signed(buffer_0_203); // @[Modules.scala 50:57:@51048.4]
  assign _T_97383 = _T_97382[10:0]; // @[Modules.scala 50:57:@51049.4]
  assign buffer_13_493 = $signed(_T_97383); // @[Modules.scala 50:57:@51050.4]
  assign _T_97385 = $signed(buffer_8_204) + $signed(buffer_1_205); // @[Modules.scala 50:57:@51052.4]
  assign _T_97386 = _T_97385[10:0]; // @[Modules.scala 50:57:@51053.4]
  assign buffer_13_494 = $signed(_T_97386); // @[Modules.scala 50:57:@51054.4]
  assign _T_97394 = $signed(buffer_5_210) + $signed(buffer_0_211); // @[Modules.scala 50:57:@51064.4]
  assign _T_97395 = _T_97394[10:0]; // @[Modules.scala 50:57:@51065.4]
  assign buffer_13_497 = $signed(_T_97395); // @[Modules.scala 50:57:@51066.4]
  assign _T_97415 = $signed(buffer_7_224) + $signed(buffer_0_225); // @[Modules.scala 50:57:@51092.4]
  assign _T_97416 = _T_97415[10:0]; // @[Modules.scala 50:57:@51093.4]
  assign buffer_13_504 = $signed(_T_97416); // @[Modules.scala 50:57:@51094.4]
  assign _T_97424 = $signed(buffer_2_230) + $signed(buffer_1_231); // @[Modules.scala 50:57:@51104.4]
  assign _T_97425 = _T_97424[10:0]; // @[Modules.scala 50:57:@51105.4]
  assign buffer_13_507 = $signed(_T_97425); // @[Modules.scala 50:57:@51106.4]
  assign _T_97427 = $signed(buffer_5_232) + $signed(buffer_1_233); // @[Modules.scala 50:57:@51108.4]
  assign _T_97428 = _T_97427[10:0]; // @[Modules.scala 50:57:@51109.4]
  assign buffer_13_508 = $signed(_T_97428); // @[Modules.scala 50:57:@51110.4]
  assign _T_97430 = $signed(buffer_0_234) + $signed(buffer_11_235); // @[Modules.scala 50:57:@51112.4]
  assign _T_97431 = _T_97430[10:0]; // @[Modules.scala 50:57:@51113.4]
  assign buffer_13_509 = $signed(_T_97431); // @[Modules.scala 50:57:@51114.4]
  assign _T_97439 = $signed(buffer_11_240) + $signed(buffer_0_241); // @[Modules.scala 50:57:@51124.4]
  assign _T_97440 = _T_97439[10:0]; // @[Modules.scala 50:57:@51125.4]
  assign buffer_13_512 = $signed(_T_97440); // @[Modules.scala 50:57:@51126.4]
  assign _T_97448 = $signed(buffer_1_246) + $signed(buffer_0_247); // @[Modules.scala 50:57:@51136.4]
  assign _T_97449 = _T_97448[10:0]; // @[Modules.scala 50:57:@51137.4]
  assign buffer_13_515 = $signed(_T_97449); // @[Modules.scala 50:57:@51138.4]
  assign buffer_13_248 = {{6{_T_96305[4]}},_T_96305}; // @[Modules.scala 32:22:@8.4]
  assign _T_97451 = $signed(buffer_13_248) + $signed(buffer_11_249); // @[Modules.scala 50:57:@51140.4]
  assign _T_97452 = _T_97451[10:0]; // @[Modules.scala 50:57:@51141.4]
  assign buffer_13_516 = $signed(_T_97452); // @[Modules.scala 50:57:@51142.4]
  assign _T_97469 = $signed(buffer_4_260) + $signed(buffer_0_261); // @[Modules.scala 50:57:@51164.4]
  assign _T_97470 = _T_97469[10:0]; // @[Modules.scala 50:57:@51165.4]
  assign buffer_13_522 = $signed(_T_97470); // @[Modules.scala 50:57:@51166.4]
  assign _T_97472 = $signed(buffer_2_262) + $signed(buffer_0_263); // @[Modules.scala 50:57:@51168.4]
  assign _T_97473 = _T_97472[10:0]; // @[Modules.scala 50:57:@51169.4]
  assign buffer_13_523 = $signed(_T_97473); // @[Modules.scala 50:57:@51170.4]
  assign buffer_13_265 = {{6{_T_96380[4]}},_T_96380}; // @[Modules.scala 32:22:@8.4]
  assign _T_97475 = $signed(buffer_0_264) + $signed(buffer_13_265); // @[Modules.scala 50:57:@51172.4]
  assign _T_97476 = _T_97475[10:0]; // @[Modules.scala 50:57:@51173.4]
  assign buffer_13_524 = $signed(_T_97476); // @[Modules.scala 50:57:@51174.4]
  assign _T_97481 = $signed(buffer_0_268) + $signed(buffer_5_269); // @[Modules.scala 50:57:@51180.4]
  assign _T_97482 = _T_97481[10:0]; // @[Modules.scala 50:57:@51181.4]
  assign buffer_13_526 = $signed(_T_97482); // @[Modules.scala 50:57:@51182.4]
  assign _T_97487 = $signed(buffer_4_272) + $signed(buffer_1_273); // @[Modules.scala 50:57:@51188.4]
  assign _T_97488 = _T_97487[10:0]; // @[Modules.scala 50:57:@51189.4]
  assign buffer_13_528 = $signed(_T_97488); // @[Modules.scala 50:57:@51190.4]
  assign _T_97499 = $signed(buffer_1_280) + $signed(buffer_0_281); // @[Modules.scala 50:57:@51204.4]
  assign _T_97500 = _T_97499[10:0]; // @[Modules.scala 50:57:@51205.4]
  assign buffer_13_532 = $signed(_T_97500); // @[Modules.scala 50:57:@51206.4]
  assign buffer_13_282 = {{6{_T_96463[4]}},_T_96463}; // @[Modules.scala 32:22:@8.4]
  assign _T_97502 = $signed(buffer_13_282) + $signed(buffer_9_283); // @[Modules.scala 50:57:@51208.4]
  assign _T_97503 = _T_97502[10:0]; // @[Modules.scala 50:57:@51209.4]
  assign buffer_13_533 = $signed(_T_97503); // @[Modules.scala 50:57:@51210.4]
  assign _T_97514 = $signed(buffer_5_290) + $signed(buffer_3_291); // @[Modules.scala 50:57:@51224.4]
  assign _T_97515 = _T_97514[10:0]; // @[Modules.scala 50:57:@51225.4]
  assign buffer_13_537 = $signed(_T_97515); // @[Modules.scala 50:57:@51226.4]
  assign _T_97517 = $signed(buffer_0_292) + $signed(buffer_4_293); // @[Modules.scala 50:57:@51228.4]
  assign _T_97518 = _T_97517[10:0]; // @[Modules.scala 50:57:@51229.4]
  assign buffer_13_538 = $signed(_T_97518); // @[Modules.scala 50:57:@51230.4]
  assign _T_97523 = $signed(buffer_12_296) + $signed(buffer_0_297); // @[Modules.scala 50:57:@51236.4]
  assign _T_97524 = _T_97523[10:0]; // @[Modules.scala 50:57:@51237.4]
  assign buffer_13_540 = $signed(_T_97524); // @[Modules.scala 50:57:@51238.4]
  assign buffer_13_309 = {{6{_T_96604[4]}},_T_96604}; // @[Modules.scala 32:22:@8.4]
  assign _T_97541 = $signed(buffer_2_308) + $signed(buffer_13_309); // @[Modules.scala 50:57:@51260.4]
  assign _T_97542 = _T_97541[10:0]; // @[Modules.scala 50:57:@51261.4]
  assign buffer_13_546 = $signed(_T_97542); // @[Modules.scala 50:57:@51262.4]
  assign _T_97544 = $signed(buffer_0_310) + $signed(buffer_4_311); // @[Modules.scala 50:57:@51264.4]
  assign _T_97545 = _T_97544[10:0]; // @[Modules.scala 50:57:@51265.4]
  assign buffer_13_547 = $signed(_T_97545); // @[Modules.scala 50:57:@51266.4]
  assign _T_97547 = $signed(buffer_2_312) + $signed(buffer_3_313); // @[Modules.scala 50:57:@51268.4]
  assign _T_97548 = _T_97547[10:0]; // @[Modules.scala 50:57:@51269.4]
  assign buffer_13_548 = $signed(_T_97548); // @[Modules.scala 50:57:@51270.4]
  assign _T_97550 = $signed(buffer_1_314) + $signed(buffer_0_315); // @[Modules.scala 50:57:@51272.4]
  assign _T_97551 = _T_97550[10:0]; // @[Modules.scala 50:57:@51273.4]
  assign buffer_13_549 = $signed(_T_97551); // @[Modules.scala 50:57:@51274.4]
  assign _T_97553 = $signed(buffer_3_316) + $signed(buffer_1_317); // @[Modules.scala 50:57:@51276.4]
  assign _T_97554 = _T_97553[10:0]; // @[Modules.scala 50:57:@51277.4]
  assign buffer_13_550 = $signed(_T_97554); // @[Modules.scala 50:57:@51278.4]
  assign buffer_13_321 = {{6{_T_96656[4]}},_T_96656}; // @[Modules.scala 32:22:@8.4]
  assign _T_97559 = $signed(buffer_0_320) + $signed(buffer_13_321); // @[Modules.scala 50:57:@51284.4]
  assign _T_97560 = _T_97559[10:0]; // @[Modules.scala 50:57:@51285.4]
  assign buffer_13_552 = $signed(_T_97560); // @[Modules.scala 50:57:@51286.4]
  assign buffer_13_329 = {{6{_T_96708[4]}},_T_96708}; // @[Modules.scala 32:22:@8.4]
  assign _T_97571 = $signed(buffer_1_328) + $signed(buffer_13_329); // @[Modules.scala 50:57:@51300.4]
  assign _T_97572 = _T_97571[10:0]; // @[Modules.scala 50:57:@51301.4]
  assign buffer_13_556 = $signed(_T_97572); // @[Modules.scala 50:57:@51302.4]
  assign _T_97583 = $signed(buffer_3_336) + $signed(buffer_6_337); // @[Modules.scala 50:57:@51316.4]
  assign _T_97584 = _T_97583[10:0]; // @[Modules.scala 50:57:@51317.4]
  assign buffer_13_560 = $signed(_T_97584); // @[Modules.scala 50:57:@51318.4]
  assign _T_97592 = $signed(buffer_0_342) + $signed(buffer_3_343); // @[Modules.scala 50:57:@51328.4]
  assign _T_97593 = _T_97592[10:0]; // @[Modules.scala 50:57:@51329.4]
  assign buffer_13_563 = $signed(_T_97593); // @[Modules.scala 50:57:@51330.4]
  assign _T_97604 = $signed(buffer_1_350) + $signed(buffer_0_351); // @[Modules.scala 50:57:@51344.4]
  assign _T_97605 = _T_97604[10:0]; // @[Modules.scala 50:57:@51345.4]
  assign buffer_13_567 = $signed(_T_97605); // @[Modules.scala 50:57:@51346.4]
  assign _T_97625 = $signed(buffer_1_364) + $signed(buffer_2_365); // @[Modules.scala 50:57:@51372.4]
  assign _T_97626 = _T_97625[10:0]; // @[Modules.scala 50:57:@51373.4]
  assign buffer_13_574 = $signed(_T_97626); // @[Modules.scala 50:57:@51374.4]
  assign _T_97646 = $signed(buffer_2_378) + $signed(buffer_8_379); // @[Modules.scala 50:57:@51400.4]
  assign _T_97647 = _T_97646[10:0]; // @[Modules.scala 50:57:@51401.4]
  assign buffer_13_581 = $signed(_T_97647); // @[Modules.scala 50:57:@51402.4]
  assign buffer_13_391 = {{6{_T_97078[4]}},_T_97078}; // @[Modules.scala 32:22:@8.4]
  assign _T_97664 = $signed(buffer_4_390) + $signed(buffer_13_391); // @[Modules.scala 50:57:@51424.4]
  assign _T_97665 = _T_97664[10:0]; // @[Modules.scala 50:57:@51425.4]
  assign buffer_13_587 = $signed(_T_97665); // @[Modules.scala 50:57:@51426.4]
  assign _T_97667 = $signed(buffer_13_392) + $signed(buffer_0_393); // @[Modules.scala 53:83:@51428.4]
  assign _T_97668 = _T_97667[10:0]; // @[Modules.scala 53:83:@51429.4]
  assign buffer_13_588 = $signed(_T_97668); // @[Modules.scala 53:83:@51430.4]
  assign _T_97670 = $signed(buffer_4_394) + $signed(buffer_13_395); // @[Modules.scala 53:83:@51432.4]
  assign _T_97671 = _T_97670[10:0]; // @[Modules.scala 53:83:@51433.4]
  assign buffer_13_589 = $signed(_T_97671); // @[Modules.scala 53:83:@51434.4]
  assign _T_97673 = $signed(buffer_2_396) + $signed(buffer_3_397); // @[Modules.scala 53:83:@51436.4]
  assign _T_97674 = _T_97673[10:0]; // @[Modules.scala 53:83:@51437.4]
  assign buffer_13_590 = $signed(_T_97674); // @[Modules.scala 53:83:@51438.4]
  assign _T_97676 = $signed(buffer_13_398) + $signed(buffer_13_399); // @[Modules.scala 53:83:@51440.4]
  assign _T_97677 = _T_97676[10:0]; // @[Modules.scala 53:83:@51441.4]
  assign buffer_13_591 = $signed(_T_97677); // @[Modules.scala 53:83:@51442.4]
  assign _T_97679 = $signed(buffer_1_400) + $signed(buffer_13_401); // @[Modules.scala 53:83:@51444.4]
  assign _T_97680 = _T_97679[10:0]; // @[Modules.scala 53:83:@51445.4]
  assign buffer_13_592 = $signed(_T_97680); // @[Modules.scala 53:83:@51446.4]
  assign _T_97682 = $signed(buffer_4_402) + $signed(buffer_3_403); // @[Modules.scala 53:83:@51448.4]
  assign _T_97683 = _T_97682[10:0]; // @[Modules.scala 53:83:@51449.4]
  assign buffer_13_593 = $signed(_T_97683); // @[Modules.scala 53:83:@51450.4]
  assign _T_97685 = $signed(buffer_0_404) + $signed(buffer_13_405); // @[Modules.scala 53:83:@51452.4]
  assign _T_97686 = _T_97685[10:0]; // @[Modules.scala 53:83:@51453.4]
  assign buffer_13_594 = $signed(_T_97686); // @[Modules.scala 53:83:@51454.4]
  assign _T_97688 = $signed(buffer_1_406) + $signed(buffer_10_407); // @[Modules.scala 53:83:@51456.4]
  assign _T_97689 = _T_97688[10:0]; // @[Modules.scala 53:83:@51457.4]
  assign buffer_13_595 = $signed(_T_97689); // @[Modules.scala 53:83:@51458.4]
  assign _T_97691 = $signed(buffer_1_408) + $signed(buffer_13_409); // @[Modules.scala 53:83:@51460.4]
  assign _T_97692 = _T_97691[10:0]; // @[Modules.scala 53:83:@51461.4]
  assign buffer_13_596 = $signed(_T_97692); // @[Modules.scala 53:83:@51462.4]
  assign _T_97694 = $signed(buffer_13_410) + $signed(buffer_1_411); // @[Modules.scala 53:83:@51464.4]
  assign _T_97695 = _T_97694[10:0]; // @[Modules.scala 53:83:@51465.4]
  assign buffer_13_597 = $signed(_T_97695); // @[Modules.scala 53:83:@51466.4]
  assign _T_97697 = $signed(buffer_13_412) + $signed(buffer_5_413); // @[Modules.scala 53:83:@51468.4]
  assign _T_97698 = _T_97697[10:0]; // @[Modules.scala 53:83:@51469.4]
  assign buffer_13_598 = $signed(_T_97698); // @[Modules.scala 53:83:@51470.4]
  assign _T_97703 = $signed(buffer_13_416) + $signed(buffer_0_417); // @[Modules.scala 53:83:@51476.4]
  assign _T_97704 = _T_97703[10:0]; // @[Modules.scala 53:83:@51477.4]
  assign buffer_13_600 = $signed(_T_97704); // @[Modules.scala 53:83:@51478.4]
  assign _T_97709 = $signed(buffer_0_420) + $signed(buffer_4_421); // @[Modules.scala 53:83:@51484.4]
  assign _T_97710 = _T_97709[10:0]; // @[Modules.scala 53:83:@51485.4]
  assign buffer_13_602 = $signed(_T_97710); // @[Modules.scala 53:83:@51486.4]
  assign _T_97712 = $signed(buffer_13_422) + $signed(buffer_12_423); // @[Modules.scala 53:83:@51488.4]
  assign _T_97713 = _T_97712[10:0]; // @[Modules.scala 53:83:@51489.4]
  assign buffer_13_603 = $signed(_T_97713); // @[Modules.scala 53:83:@51490.4]
  assign _T_97718 = $signed(buffer_10_426) + $signed(buffer_4_427); // @[Modules.scala 53:83:@51496.4]
  assign _T_97719 = _T_97718[10:0]; // @[Modules.scala 53:83:@51497.4]
  assign buffer_13_605 = $signed(_T_97719); // @[Modules.scala 53:83:@51498.4]
  assign _T_97721 = $signed(buffer_7_428) + $signed(buffer_3_429); // @[Modules.scala 53:83:@51500.4]
  assign _T_97722 = _T_97721[10:0]; // @[Modules.scala 53:83:@51501.4]
  assign buffer_13_606 = $signed(_T_97722); // @[Modules.scala 53:83:@51502.4]
  assign _T_97724 = $signed(buffer_4_430) + $signed(buffer_13_431); // @[Modules.scala 53:83:@51504.4]
  assign _T_97725 = _T_97724[10:0]; // @[Modules.scala 53:83:@51505.4]
  assign buffer_13_607 = $signed(_T_97725); // @[Modules.scala 53:83:@51506.4]
  assign _T_97727 = $signed(buffer_13_432) + $signed(buffer_12_433); // @[Modules.scala 53:83:@51508.4]
  assign _T_97728 = _T_97727[10:0]; // @[Modules.scala 53:83:@51509.4]
  assign buffer_13_608 = $signed(_T_97728); // @[Modules.scala 53:83:@51510.4]
  assign _T_97730 = $signed(buffer_13_434) + $signed(buffer_2_435); // @[Modules.scala 53:83:@51512.4]
  assign _T_97731 = _T_97730[10:0]; // @[Modules.scala 53:83:@51513.4]
  assign buffer_13_609 = $signed(_T_97731); // @[Modules.scala 53:83:@51514.4]
  assign _T_97733 = $signed(buffer_0_436) + $signed(buffer_13_437); // @[Modules.scala 53:83:@51516.4]
  assign _T_97734 = _T_97733[10:0]; // @[Modules.scala 53:83:@51517.4]
  assign buffer_13_610 = $signed(_T_97734); // @[Modules.scala 53:83:@51518.4]
  assign _T_97736 = $signed(buffer_13_438) + $signed(buffer_13_439); // @[Modules.scala 53:83:@51520.4]
  assign _T_97737 = _T_97736[10:0]; // @[Modules.scala 53:83:@51521.4]
  assign buffer_13_611 = $signed(_T_97737); // @[Modules.scala 53:83:@51522.4]
  assign _T_97739 = $signed(buffer_0_440) + $signed(buffer_13_441); // @[Modules.scala 53:83:@51524.4]
  assign _T_97740 = _T_97739[10:0]; // @[Modules.scala 53:83:@51525.4]
  assign buffer_13_612 = $signed(_T_97740); // @[Modules.scala 53:83:@51526.4]
  assign _T_97742 = $signed(buffer_13_442) + $signed(buffer_9_443); // @[Modules.scala 53:83:@51528.4]
  assign _T_97743 = _T_97742[10:0]; // @[Modules.scala 53:83:@51529.4]
  assign buffer_13_613 = $signed(_T_97743); // @[Modules.scala 53:83:@51530.4]
  assign _T_97745 = $signed(buffer_13_444) + $signed(buffer_11_445); // @[Modules.scala 53:83:@51532.4]
  assign _T_97746 = _T_97745[10:0]; // @[Modules.scala 53:83:@51533.4]
  assign buffer_13_614 = $signed(_T_97746); // @[Modules.scala 53:83:@51534.4]
  assign _T_97748 = $signed(buffer_3_446) + $signed(buffer_0_447); // @[Modules.scala 53:83:@51536.4]
  assign _T_97749 = _T_97748[10:0]; // @[Modules.scala 53:83:@51537.4]
  assign buffer_13_615 = $signed(_T_97749); // @[Modules.scala 53:83:@51538.4]
  assign _T_97751 = $signed(buffer_13_448) + $signed(buffer_13_449); // @[Modules.scala 53:83:@51540.4]
  assign _T_97752 = _T_97751[10:0]; // @[Modules.scala 53:83:@51541.4]
  assign buffer_13_616 = $signed(_T_97752); // @[Modules.scala 53:83:@51542.4]
  assign _T_97754 = $signed(buffer_4_450) + $signed(buffer_0_451); // @[Modules.scala 53:83:@51544.4]
  assign _T_97755 = _T_97754[10:0]; // @[Modules.scala 53:83:@51545.4]
  assign buffer_13_617 = $signed(_T_97755); // @[Modules.scala 53:83:@51546.4]
  assign _T_97757 = $signed(buffer_13_452) + $signed(buffer_0_453); // @[Modules.scala 53:83:@51548.4]
  assign _T_97758 = _T_97757[10:0]; // @[Modules.scala 53:83:@51549.4]
  assign buffer_13_618 = $signed(_T_97758); // @[Modules.scala 53:83:@51550.4]
  assign _T_97763 = $signed(buffer_0_456) + $signed(buffer_13_457); // @[Modules.scala 53:83:@51556.4]
  assign _T_97764 = _T_97763[10:0]; // @[Modules.scala 53:83:@51557.4]
  assign buffer_13_620 = $signed(_T_97764); // @[Modules.scala 53:83:@51558.4]
  assign _T_97766 = $signed(buffer_13_458) + $signed(buffer_7_459); // @[Modules.scala 53:83:@51560.4]
  assign _T_97767 = _T_97766[10:0]; // @[Modules.scala 53:83:@51561.4]
  assign buffer_13_621 = $signed(_T_97767); // @[Modules.scala 53:83:@51562.4]
  assign _T_97769 = $signed(buffer_13_460) + $signed(buffer_0_461); // @[Modules.scala 53:83:@51564.4]
  assign _T_97770 = _T_97769[10:0]; // @[Modules.scala 53:83:@51565.4]
  assign buffer_13_622 = $signed(_T_97770); // @[Modules.scala 53:83:@51566.4]
  assign _T_97772 = $signed(buffer_0_462) + $signed(buffer_11_463); // @[Modules.scala 53:83:@51568.4]
  assign _T_97773 = _T_97772[10:0]; // @[Modules.scala 53:83:@51569.4]
  assign buffer_13_623 = $signed(_T_97773); // @[Modules.scala 53:83:@51570.4]
  assign _T_97775 = $signed(buffer_13_464) + $signed(buffer_7_465); // @[Modules.scala 53:83:@51572.4]
  assign _T_97776 = _T_97775[10:0]; // @[Modules.scala 53:83:@51573.4]
  assign buffer_13_624 = $signed(_T_97776); // @[Modules.scala 53:83:@51574.4]
  assign _T_97778 = $signed(buffer_13_466) + $signed(buffer_13_467); // @[Modules.scala 53:83:@51576.4]
  assign _T_97779 = _T_97778[10:0]; // @[Modules.scala 53:83:@51577.4]
  assign buffer_13_625 = $signed(_T_97779); // @[Modules.scala 53:83:@51578.4]
  assign _T_97784 = $signed(buffer_13_470) + $signed(buffer_13_471); // @[Modules.scala 53:83:@51584.4]
  assign _T_97785 = _T_97784[10:0]; // @[Modules.scala 53:83:@51585.4]
  assign buffer_13_627 = $signed(_T_97785); // @[Modules.scala 53:83:@51586.4]
  assign _T_97787 = $signed(buffer_4_472) + $signed(buffer_13_473); // @[Modules.scala 53:83:@51588.4]
  assign _T_97788 = _T_97787[10:0]; // @[Modules.scala 53:83:@51589.4]
  assign buffer_13_628 = $signed(_T_97788); // @[Modules.scala 53:83:@51590.4]
  assign _T_97790 = $signed(buffer_5_474) + $signed(buffer_12_475); // @[Modules.scala 53:83:@51592.4]
  assign _T_97791 = _T_97790[10:0]; // @[Modules.scala 53:83:@51593.4]
  assign buffer_13_629 = $signed(_T_97791); // @[Modules.scala 53:83:@51594.4]
  assign _T_97793 = $signed(buffer_13_476) + $signed(buffer_13_477); // @[Modules.scala 53:83:@51596.4]
  assign _T_97794 = _T_97793[10:0]; // @[Modules.scala 53:83:@51597.4]
  assign buffer_13_630 = $signed(_T_97794); // @[Modules.scala 53:83:@51598.4]
  assign _T_97796 = $signed(buffer_13_478) + $signed(buffer_13_479); // @[Modules.scala 53:83:@51600.4]
  assign _T_97797 = _T_97796[10:0]; // @[Modules.scala 53:83:@51601.4]
  assign buffer_13_631 = $signed(_T_97797); // @[Modules.scala 53:83:@51602.4]
  assign _T_97799 = $signed(buffer_13_480) + $signed(buffer_0_481); // @[Modules.scala 53:83:@51604.4]
  assign _T_97800 = _T_97799[10:0]; // @[Modules.scala 53:83:@51605.4]
  assign buffer_13_632 = $signed(_T_97800); // @[Modules.scala 53:83:@51606.4]
  assign _T_97802 = $signed(buffer_4_482) + $signed(buffer_13_483); // @[Modules.scala 53:83:@51608.4]
  assign _T_97803 = _T_97802[10:0]; // @[Modules.scala 53:83:@51609.4]
  assign buffer_13_633 = $signed(_T_97803); // @[Modules.scala 53:83:@51610.4]
  assign _T_97805 = $signed(buffer_11_484) + $signed(buffer_13_485); // @[Modules.scala 53:83:@51612.4]
  assign _T_97806 = _T_97805[10:0]; // @[Modules.scala 53:83:@51613.4]
  assign buffer_13_634 = $signed(_T_97806); // @[Modules.scala 53:83:@51614.4]
  assign _T_97808 = $signed(buffer_3_486) + $signed(buffer_13_487); // @[Modules.scala 53:83:@51616.4]
  assign _T_97809 = _T_97808[10:0]; // @[Modules.scala 53:83:@51617.4]
  assign buffer_13_635 = $signed(_T_97809); // @[Modules.scala 53:83:@51618.4]
  assign _T_97811 = $signed(buffer_13_488) + $signed(buffer_9_489); // @[Modules.scala 53:83:@51620.4]
  assign _T_97812 = _T_97811[10:0]; // @[Modules.scala 53:83:@51621.4]
  assign buffer_13_636 = $signed(_T_97812); // @[Modules.scala 53:83:@51622.4]
  assign _T_97814 = $signed(buffer_12_490) + $signed(buffer_1_491); // @[Modules.scala 53:83:@51624.4]
  assign _T_97815 = _T_97814[10:0]; // @[Modules.scala 53:83:@51625.4]
  assign buffer_13_637 = $signed(_T_97815); // @[Modules.scala 53:83:@51626.4]
  assign _T_97817 = $signed(buffer_0_492) + $signed(buffer_13_493); // @[Modules.scala 53:83:@51628.4]
  assign _T_97818 = _T_97817[10:0]; // @[Modules.scala 53:83:@51629.4]
  assign buffer_13_638 = $signed(_T_97818); // @[Modules.scala 53:83:@51630.4]
  assign _T_97820 = $signed(buffer_13_494) + $signed(buffer_0_495); // @[Modules.scala 53:83:@51632.4]
  assign _T_97821 = _T_97820[10:0]; // @[Modules.scala 53:83:@51633.4]
  assign buffer_13_639 = $signed(_T_97821); // @[Modules.scala 53:83:@51634.4]
  assign _T_97823 = $signed(buffer_10_496) + $signed(buffer_13_497); // @[Modules.scala 53:83:@51636.4]
  assign _T_97824 = _T_97823[10:0]; // @[Modules.scala 53:83:@51637.4]
  assign buffer_13_640 = $signed(_T_97824); // @[Modules.scala 53:83:@51638.4]
  assign _T_97826 = $signed(buffer_7_498) + $signed(buffer_0_499); // @[Modules.scala 53:83:@51640.4]
  assign _T_97827 = _T_97826[10:0]; // @[Modules.scala 53:83:@51641.4]
  assign buffer_13_641 = $signed(_T_97827); // @[Modules.scala 53:83:@51642.4]
  assign _T_97829 = $signed(buffer_11_500) + $signed(buffer_5_501); // @[Modules.scala 53:83:@51644.4]
  assign _T_97830 = _T_97829[10:0]; // @[Modules.scala 53:83:@51645.4]
  assign buffer_13_642 = $signed(_T_97830); // @[Modules.scala 53:83:@51646.4]
  assign _T_97832 = $signed(buffer_2_502) + $signed(buffer_3_503); // @[Modules.scala 53:83:@51648.4]
  assign _T_97833 = _T_97832[10:0]; // @[Modules.scala 53:83:@51649.4]
  assign buffer_13_643 = $signed(_T_97833); // @[Modules.scala 53:83:@51650.4]
  assign _T_97835 = $signed(buffer_13_504) + $signed(buffer_0_505); // @[Modules.scala 53:83:@51652.4]
  assign _T_97836 = _T_97835[10:0]; // @[Modules.scala 53:83:@51653.4]
  assign buffer_13_644 = $signed(_T_97836); // @[Modules.scala 53:83:@51654.4]
  assign _T_97838 = $signed(buffer_0_506) + $signed(buffer_13_507); // @[Modules.scala 53:83:@51656.4]
  assign _T_97839 = _T_97838[10:0]; // @[Modules.scala 53:83:@51657.4]
  assign buffer_13_645 = $signed(_T_97839); // @[Modules.scala 53:83:@51658.4]
  assign _T_97841 = $signed(buffer_13_508) + $signed(buffer_13_509); // @[Modules.scala 53:83:@51660.4]
  assign _T_97842 = _T_97841[10:0]; // @[Modules.scala 53:83:@51661.4]
  assign buffer_13_646 = $signed(_T_97842); // @[Modules.scala 53:83:@51662.4]
  assign _T_97847 = $signed(buffer_13_512) + $signed(buffer_0_513); // @[Modules.scala 53:83:@51668.4]
  assign _T_97848 = _T_97847[10:0]; // @[Modules.scala 53:83:@51669.4]
  assign buffer_13_648 = $signed(_T_97848); // @[Modules.scala 53:83:@51670.4]
  assign _T_97850 = $signed(buffer_2_514) + $signed(buffer_13_515); // @[Modules.scala 53:83:@51672.4]
  assign _T_97851 = _T_97850[10:0]; // @[Modules.scala 53:83:@51673.4]
  assign buffer_13_649 = $signed(_T_97851); // @[Modules.scala 53:83:@51674.4]
  assign _T_97853 = $signed(buffer_13_516) + $signed(buffer_3_517); // @[Modules.scala 53:83:@51676.4]
  assign _T_97854 = _T_97853[10:0]; // @[Modules.scala 53:83:@51677.4]
  assign buffer_13_650 = $signed(_T_97854); // @[Modules.scala 53:83:@51678.4]
  assign _T_97862 = $signed(buffer_13_522) + $signed(buffer_13_523); // @[Modules.scala 53:83:@51688.4]
  assign _T_97863 = _T_97862[10:0]; // @[Modules.scala 53:83:@51689.4]
  assign buffer_13_653 = $signed(_T_97863); // @[Modules.scala 53:83:@51690.4]
  assign _T_97865 = $signed(buffer_13_524) + $signed(buffer_2_525); // @[Modules.scala 53:83:@51692.4]
  assign _T_97866 = _T_97865[10:0]; // @[Modules.scala 53:83:@51693.4]
  assign buffer_13_654 = $signed(_T_97866); // @[Modules.scala 53:83:@51694.4]
  assign _T_97868 = $signed(buffer_13_526) + $signed(buffer_1_527); // @[Modules.scala 53:83:@51696.4]
  assign _T_97869 = _T_97868[10:0]; // @[Modules.scala 53:83:@51697.4]
  assign buffer_13_655 = $signed(_T_97869); // @[Modules.scala 53:83:@51698.4]
  assign _T_97871 = $signed(buffer_13_528) + $signed(buffer_7_529); // @[Modules.scala 53:83:@51700.4]
  assign _T_97872 = _T_97871[10:0]; // @[Modules.scala 53:83:@51701.4]
  assign buffer_13_656 = $signed(_T_97872); // @[Modules.scala 53:83:@51702.4]
  assign _T_97877 = $signed(buffer_13_532) + $signed(buffer_13_533); // @[Modules.scala 53:83:@51708.4]
  assign _T_97878 = _T_97877[10:0]; // @[Modules.scala 53:83:@51709.4]
  assign buffer_13_658 = $signed(_T_97878); // @[Modules.scala 53:83:@51710.4]
  assign _T_97883 = $signed(buffer_5_536) + $signed(buffer_13_537); // @[Modules.scala 53:83:@51716.4]
  assign _T_97884 = _T_97883[10:0]; // @[Modules.scala 53:83:@51717.4]
  assign buffer_13_660 = $signed(_T_97884); // @[Modules.scala 53:83:@51718.4]
  assign _T_97886 = $signed(buffer_13_538) + $signed(buffer_6_539); // @[Modules.scala 53:83:@51720.4]
  assign _T_97887 = _T_97886[10:0]; // @[Modules.scala 53:83:@51721.4]
  assign buffer_13_661 = $signed(_T_97887); // @[Modules.scala 53:83:@51722.4]
  assign _T_97889 = $signed(buffer_13_540) + $signed(buffer_0_541); // @[Modules.scala 53:83:@51724.4]
  assign _T_97890 = _T_97889[10:0]; // @[Modules.scala 53:83:@51725.4]
  assign buffer_13_662 = $signed(_T_97890); // @[Modules.scala 53:83:@51726.4]
  assign _T_97898 = $signed(buffer_13_546) + $signed(buffer_13_547); // @[Modules.scala 53:83:@51736.4]
  assign _T_97899 = _T_97898[10:0]; // @[Modules.scala 53:83:@51737.4]
  assign buffer_13_665 = $signed(_T_97899); // @[Modules.scala 53:83:@51738.4]
  assign _T_97901 = $signed(buffer_13_548) + $signed(buffer_13_549); // @[Modules.scala 53:83:@51740.4]
  assign _T_97902 = _T_97901[10:0]; // @[Modules.scala 53:83:@51741.4]
  assign buffer_13_666 = $signed(_T_97902); // @[Modules.scala 53:83:@51742.4]
  assign _T_97904 = $signed(buffer_13_550) + $signed(buffer_3_551); // @[Modules.scala 53:83:@51744.4]
  assign _T_97905 = _T_97904[10:0]; // @[Modules.scala 53:83:@51745.4]
  assign buffer_13_667 = $signed(_T_97905); // @[Modules.scala 53:83:@51746.4]
  assign _T_97907 = $signed(buffer_13_552) + $signed(buffer_6_553); // @[Modules.scala 53:83:@51748.4]
  assign _T_97908 = _T_97907[10:0]; // @[Modules.scala 53:83:@51749.4]
  assign buffer_13_668 = $signed(_T_97908); // @[Modules.scala 53:83:@51750.4]
  assign _T_97913 = $signed(buffer_13_556) + $signed(buffer_1_557); // @[Modules.scala 53:83:@51756.4]
  assign _T_97914 = _T_97913[10:0]; // @[Modules.scala 53:83:@51757.4]
  assign buffer_13_670 = $signed(_T_97914); // @[Modules.scala 53:83:@51758.4]
  assign _T_97919 = $signed(buffer_13_560) + $signed(buffer_2_561); // @[Modules.scala 53:83:@51764.4]
  assign _T_97920 = _T_97919[10:0]; // @[Modules.scala 53:83:@51765.4]
  assign buffer_13_672 = $signed(_T_97920); // @[Modules.scala 53:83:@51766.4]
  assign _T_97922 = $signed(buffer_2_562) + $signed(buffer_13_563); // @[Modules.scala 53:83:@51768.4]
  assign _T_97923 = _T_97922[10:0]; // @[Modules.scala 53:83:@51769.4]
  assign buffer_13_673 = $signed(_T_97923); // @[Modules.scala 53:83:@51770.4]
  assign _T_97928 = $signed(buffer_0_566) + $signed(buffer_13_567); // @[Modules.scala 53:83:@51776.4]
  assign _T_97929 = _T_97928[10:0]; // @[Modules.scala 53:83:@51777.4]
  assign buffer_13_675 = $signed(_T_97929); // @[Modules.scala 53:83:@51778.4]
  assign _T_97937 = $signed(buffer_3_572) + $signed(buffer_6_573); // @[Modules.scala 53:83:@51788.4]
  assign _T_97938 = _T_97937[10:0]; // @[Modules.scala 53:83:@51789.4]
  assign buffer_13_678 = $signed(_T_97938); // @[Modules.scala 53:83:@51790.4]
  assign _T_97940 = $signed(buffer_13_574) + $signed(buffer_1_575); // @[Modules.scala 53:83:@51792.4]
  assign _T_97941 = _T_97940[10:0]; // @[Modules.scala 53:83:@51793.4]
  assign buffer_13_679 = $signed(_T_97941); // @[Modules.scala 53:83:@51794.4]
  assign _T_97949 = $signed(buffer_7_580) + $signed(buffer_13_581); // @[Modules.scala 53:83:@51804.4]
  assign _T_97950 = _T_97949[10:0]; // @[Modules.scala 53:83:@51805.4]
  assign buffer_13_682 = $signed(_T_97950); // @[Modules.scala 53:83:@51806.4]
  assign _T_97958 = $signed(buffer_1_586) + $signed(buffer_13_587); // @[Modules.scala 53:83:@51816.4]
  assign _T_97959 = _T_97958[10:0]; // @[Modules.scala 53:83:@51817.4]
  assign buffer_13_685 = $signed(_T_97959); // @[Modules.scala 53:83:@51818.4]
  assign _T_97961 = $signed(buffer_13_588) + $signed(buffer_13_589); // @[Modules.scala 56:109:@51820.4]
  assign _T_97962 = _T_97961[10:0]; // @[Modules.scala 56:109:@51821.4]
  assign buffer_13_686 = $signed(_T_97962); // @[Modules.scala 56:109:@51822.4]
  assign _T_97964 = $signed(buffer_13_590) + $signed(buffer_13_591); // @[Modules.scala 56:109:@51824.4]
  assign _T_97965 = _T_97964[10:0]; // @[Modules.scala 56:109:@51825.4]
  assign buffer_13_687 = $signed(_T_97965); // @[Modules.scala 56:109:@51826.4]
  assign _T_97967 = $signed(buffer_13_592) + $signed(buffer_13_593); // @[Modules.scala 56:109:@51828.4]
  assign _T_97968 = _T_97967[10:0]; // @[Modules.scala 56:109:@51829.4]
  assign buffer_13_688 = $signed(_T_97968); // @[Modules.scala 56:109:@51830.4]
  assign _T_97970 = $signed(buffer_13_594) + $signed(buffer_13_595); // @[Modules.scala 56:109:@51832.4]
  assign _T_97971 = _T_97970[10:0]; // @[Modules.scala 56:109:@51833.4]
  assign buffer_13_689 = $signed(_T_97971); // @[Modules.scala 56:109:@51834.4]
  assign _T_97973 = $signed(buffer_13_596) + $signed(buffer_13_597); // @[Modules.scala 56:109:@51836.4]
  assign _T_97974 = _T_97973[10:0]; // @[Modules.scala 56:109:@51837.4]
  assign buffer_13_690 = $signed(_T_97974); // @[Modules.scala 56:109:@51838.4]
  assign _T_97976 = $signed(buffer_13_598) + $signed(buffer_0_599); // @[Modules.scala 56:109:@51840.4]
  assign _T_97977 = _T_97976[10:0]; // @[Modules.scala 56:109:@51841.4]
  assign buffer_13_691 = $signed(_T_97977); // @[Modules.scala 56:109:@51842.4]
  assign _T_97979 = $signed(buffer_13_600) + $signed(buffer_1_601); // @[Modules.scala 56:109:@51844.4]
  assign _T_97980 = _T_97979[10:0]; // @[Modules.scala 56:109:@51845.4]
  assign buffer_13_692 = $signed(_T_97980); // @[Modules.scala 56:109:@51846.4]
  assign _T_97982 = $signed(buffer_13_602) + $signed(buffer_13_603); // @[Modules.scala 56:109:@51848.4]
  assign _T_97983 = _T_97982[10:0]; // @[Modules.scala 56:109:@51849.4]
  assign buffer_13_693 = $signed(_T_97983); // @[Modules.scala 56:109:@51850.4]
  assign _T_97985 = $signed(buffer_8_604) + $signed(buffer_13_605); // @[Modules.scala 56:109:@51852.4]
  assign _T_97986 = _T_97985[10:0]; // @[Modules.scala 56:109:@51853.4]
  assign buffer_13_694 = $signed(_T_97986); // @[Modules.scala 56:109:@51854.4]
  assign _T_97988 = $signed(buffer_13_606) + $signed(buffer_13_607); // @[Modules.scala 56:109:@51856.4]
  assign _T_97989 = _T_97988[10:0]; // @[Modules.scala 56:109:@51857.4]
  assign buffer_13_695 = $signed(_T_97989); // @[Modules.scala 56:109:@51858.4]
  assign _T_97991 = $signed(buffer_13_608) + $signed(buffer_13_609); // @[Modules.scala 56:109:@51860.4]
  assign _T_97992 = _T_97991[10:0]; // @[Modules.scala 56:109:@51861.4]
  assign buffer_13_696 = $signed(_T_97992); // @[Modules.scala 56:109:@51862.4]
  assign _T_97994 = $signed(buffer_13_610) + $signed(buffer_13_611); // @[Modules.scala 56:109:@51864.4]
  assign _T_97995 = _T_97994[10:0]; // @[Modules.scala 56:109:@51865.4]
  assign buffer_13_697 = $signed(_T_97995); // @[Modules.scala 56:109:@51866.4]
  assign _T_97997 = $signed(buffer_13_612) + $signed(buffer_13_613); // @[Modules.scala 56:109:@51868.4]
  assign _T_97998 = _T_97997[10:0]; // @[Modules.scala 56:109:@51869.4]
  assign buffer_13_698 = $signed(_T_97998); // @[Modules.scala 56:109:@51870.4]
  assign _T_98000 = $signed(buffer_13_614) + $signed(buffer_13_615); // @[Modules.scala 56:109:@51872.4]
  assign _T_98001 = _T_98000[10:0]; // @[Modules.scala 56:109:@51873.4]
  assign buffer_13_699 = $signed(_T_98001); // @[Modules.scala 56:109:@51874.4]
  assign _T_98003 = $signed(buffer_13_616) + $signed(buffer_13_617); // @[Modules.scala 56:109:@51876.4]
  assign _T_98004 = _T_98003[10:0]; // @[Modules.scala 56:109:@51877.4]
  assign buffer_13_700 = $signed(_T_98004); // @[Modules.scala 56:109:@51878.4]
  assign _T_98006 = $signed(buffer_13_618) + $signed(buffer_0_619); // @[Modules.scala 56:109:@51880.4]
  assign _T_98007 = _T_98006[10:0]; // @[Modules.scala 56:109:@51881.4]
  assign buffer_13_701 = $signed(_T_98007); // @[Modules.scala 56:109:@51882.4]
  assign _T_98009 = $signed(buffer_13_620) + $signed(buffer_13_621); // @[Modules.scala 56:109:@51884.4]
  assign _T_98010 = _T_98009[10:0]; // @[Modules.scala 56:109:@51885.4]
  assign buffer_13_702 = $signed(_T_98010); // @[Modules.scala 56:109:@51886.4]
  assign _T_98012 = $signed(buffer_13_622) + $signed(buffer_13_623); // @[Modules.scala 56:109:@51888.4]
  assign _T_98013 = _T_98012[10:0]; // @[Modules.scala 56:109:@51889.4]
  assign buffer_13_703 = $signed(_T_98013); // @[Modules.scala 56:109:@51890.4]
  assign _T_98015 = $signed(buffer_13_624) + $signed(buffer_13_625); // @[Modules.scala 56:109:@51892.4]
  assign _T_98016 = _T_98015[10:0]; // @[Modules.scala 56:109:@51893.4]
  assign buffer_13_704 = $signed(_T_98016); // @[Modules.scala 56:109:@51894.4]
  assign _T_98018 = $signed(buffer_0_626) + $signed(buffer_13_627); // @[Modules.scala 56:109:@51896.4]
  assign _T_98019 = _T_98018[10:0]; // @[Modules.scala 56:109:@51897.4]
  assign buffer_13_705 = $signed(_T_98019); // @[Modules.scala 56:109:@51898.4]
  assign _T_98021 = $signed(buffer_13_628) + $signed(buffer_13_629); // @[Modules.scala 56:109:@51900.4]
  assign _T_98022 = _T_98021[10:0]; // @[Modules.scala 56:109:@51901.4]
  assign buffer_13_706 = $signed(_T_98022); // @[Modules.scala 56:109:@51902.4]
  assign _T_98024 = $signed(buffer_13_630) + $signed(buffer_13_631); // @[Modules.scala 56:109:@51904.4]
  assign _T_98025 = _T_98024[10:0]; // @[Modules.scala 56:109:@51905.4]
  assign buffer_13_707 = $signed(_T_98025); // @[Modules.scala 56:109:@51906.4]
  assign _T_98027 = $signed(buffer_13_632) + $signed(buffer_13_633); // @[Modules.scala 56:109:@51908.4]
  assign _T_98028 = _T_98027[10:0]; // @[Modules.scala 56:109:@51909.4]
  assign buffer_13_708 = $signed(_T_98028); // @[Modules.scala 56:109:@51910.4]
  assign _T_98030 = $signed(buffer_13_634) + $signed(buffer_13_635); // @[Modules.scala 56:109:@51912.4]
  assign _T_98031 = _T_98030[10:0]; // @[Modules.scala 56:109:@51913.4]
  assign buffer_13_709 = $signed(_T_98031); // @[Modules.scala 56:109:@51914.4]
  assign _T_98033 = $signed(buffer_13_636) + $signed(buffer_13_637); // @[Modules.scala 56:109:@51916.4]
  assign _T_98034 = _T_98033[10:0]; // @[Modules.scala 56:109:@51917.4]
  assign buffer_13_710 = $signed(_T_98034); // @[Modules.scala 56:109:@51918.4]
  assign _T_98036 = $signed(buffer_13_638) + $signed(buffer_13_639); // @[Modules.scala 56:109:@51920.4]
  assign _T_98037 = _T_98036[10:0]; // @[Modules.scala 56:109:@51921.4]
  assign buffer_13_711 = $signed(_T_98037); // @[Modules.scala 56:109:@51922.4]
  assign _T_98039 = $signed(buffer_13_640) + $signed(buffer_13_641); // @[Modules.scala 56:109:@51924.4]
  assign _T_98040 = _T_98039[10:0]; // @[Modules.scala 56:109:@51925.4]
  assign buffer_13_712 = $signed(_T_98040); // @[Modules.scala 56:109:@51926.4]
  assign _T_98042 = $signed(buffer_13_642) + $signed(buffer_13_643); // @[Modules.scala 56:109:@51928.4]
  assign _T_98043 = _T_98042[10:0]; // @[Modules.scala 56:109:@51929.4]
  assign buffer_13_713 = $signed(_T_98043); // @[Modules.scala 56:109:@51930.4]
  assign _T_98045 = $signed(buffer_13_644) + $signed(buffer_13_645); // @[Modules.scala 56:109:@51932.4]
  assign _T_98046 = _T_98045[10:0]; // @[Modules.scala 56:109:@51933.4]
  assign buffer_13_714 = $signed(_T_98046); // @[Modules.scala 56:109:@51934.4]
  assign _T_98048 = $signed(buffer_13_646) + $signed(buffer_7_647); // @[Modules.scala 56:109:@51936.4]
  assign _T_98049 = _T_98048[10:0]; // @[Modules.scala 56:109:@51937.4]
  assign buffer_13_715 = $signed(_T_98049); // @[Modules.scala 56:109:@51938.4]
  assign _T_98051 = $signed(buffer_13_648) + $signed(buffer_13_649); // @[Modules.scala 56:109:@51940.4]
  assign _T_98052 = _T_98051[10:0]; // @[Modules.scala 56:109:@51941.4]
  assign buffer_13_716 = $signed(_T_98052); // @[Modules.scala 56:109:@51942.4]
  assign _T_98054 = $signed(buffer_13_650) + $signed(buffer_11_651); // @[Modules.scala 56:109:@51944.4]
  assign _T_98055 = _T_98054[10:0]; // @[Modules.scala 56:109:@51945.4]
  assign buffer_13_717 = $signed(_T_98055); // @[Modules.scala 56:109:@51946.4]
  assign _T_98057 = $signed(buffer_7_652) + $signed(buffer_13_653); // @[Modules.scala 56:109:@51948.4]
  assign _T_98058 = _T_98057[10:0]; // @[Modules.scala 56:109:@51949.4]
  assign buffer_13_718 = $signed(_T_98058); // @[Modules.scala 56:109:@51950.4]
  assign _T_98060 = $signed(buffer_13_654) + $signed(buffer_13_655); // @[Modules.scala 56:109:@51952.4]
  assign _T_98061 = _T_98060[10:0]; // @[Modules.scala 56:109:@51953.4]
  assign buffer_13_719 = $signed(_T_98061); // @[Modules.scala 56:109:@51954.4]
  assign _T_98063 = $signed(buffer_13_656) + $signed(buffer_3_657); // @[Modules.scala 56:109:@51956.4]
  assign _T_98064 = _T_98063[10:0]; // @[Modules.scala 56:109:@51957.4]
  assign buffer_13_720 = $signed(_T_98064); // @[Modules.scala 56:109:@51958.4]
  assign _T_98066 = $signed(buffer_13_658) + $signed(buffer_9_659); // @[Modules.scala 56:109:@51960.4]
  assign _T_98067 = _T_98066[10:0]; // @[Modules.scala 56:109:@51961.4]
  assign buffer_13_721 = $signed(_T_98067); // @[Modules.scala 56:109:@51962.4]
  assign _T_98069 = $signed(buffer_13_660) + $signed(buffer_13_661); // @[Modules.scala 56:109:@51964.4]
  assign _T_98070 = _T_98069[10:0]; // @[Modules.scala 56:109:@51965.4]
  assign buffer_13_722 = $signed(_T_98070); // @[Modules.scala 56:109:@51966.4]
  assign _T_98072 = $signed(buffer_13_662) + $signed(buffer_7_663); // @[Modules.scala 56:109:@51968.4]
  assign _T_98073 = _T_98072[10:0]; // @[Modules.scala 56:109:@51969.4]
  assign buffer_13_723 = $signed(_T_98073); // @[Modules.scala 56:109:@51970.4]
  assign _T_98075 = $signed(buffer_3_664) + $signed(buffer_13_665); // @[Modules.scala 56:109:@51972.4]
  assign _T_98076 = _T_98075[10:0]; // @[Modules.scala 56:109:@51973.4]
  assign buffer_13_724 = $signed(_T_98076); // @[Modules.scala 56:109:@51974.4]
  assign _T_98078 = $signed(buffer_13_666) + $signed(buffer_13_667); // @[Modules.scala 56:109:@51976.4]
  assign _T_98079 = _T_98078[10:0]; // @[Modules.scala 56:109:@51977.4]
  assign buffer_13_725 = $signed(_T_98079); // @[Modules.scala 56:109:@51978.4]
  assign _T_98081 = $signed(buffer_13_668) + $signed(buffer_0_669); // @[Modules.scala 56:109:@51980.4]
  assign _T_98082 = _T_98081[10:0]; // @[Modules.scala 56:109:@51981.4]
  assign buffer_13_726 = $signed(_T_98082); // @[Modules.scala 56:109:@51982.4]
  assign _T_98084 = $signed(buffer_13_670) + $signed(buffer_0_671); // @[Modules.scala 56:109:@51984.4]
  assign _T_98085 = _T_98084[10:0]; // @[Modules.scala 56:109:@51985.4]
  assign buffer_13_727 = $signed(_T_98085); // @[Modules.scala 56:109:@51986.4]
  assign _T_98087 = $signed(buffer_13_672) + $signed(buffer_13_673); // @[Modules.scala 56:109:@51988.4]
  assign _T_98088 = _T_98087[10:0]; // @[Modules.scala 56:109:@51989.4]
  assign buffer_13_728 = $signed(_T_98088); // @[Modules.scala 56:109:@51990.4]
  assign _T_98090 = $signed(buffer_0_674) + $signed(buffer_13_675); // @[Modules.scala 56:109:@51992.4]
  assign _T_98091 = _T_98090[10:0]; // @[Modules.scala 56:109:@51993.4]
  assign buffer_13_729 = $signed(_T_98091); // @[Modules.scala 56:109:@51994.4]
  assign _T_98096 = $signed(buffer_13_678) + $signed(buffer_13_679); // @[Modules.scala 56:109:@52000.4]
  assign _T_98097 = _T_98096[10:0]; // @[Modules.scala 56:109:@52001.4]
  assign buffer_13_731 = $signed(_T_98097); // @[Modules.scala 56:109:@52002.4]
  assign _T_98102 = $signed(buffer_13_682) + $signed(buffer_6_683); // @[Modules.scala 56:109:@52008.4]
  assign _T_98103 = _T_98102[10:0]; // @[Modules.scala 56:109:@52009.4]
  assign buffer_13_733 = $signed(_T_98103); // @[Modules.scala 56:109:@52010.4]
  assign _T_98105 = $signed(buffer_1_684) + $signed(buffer_13_685); // @[Modules.scala 56:109:@52012.4]
  assign _T_98106 = _T_98105[10:0]; // @[Modules.scala 56:109:@52013.4]
  assign buffer_13_734 = $signed(_T_98106); // @[Modules.scala 56:109:@52014.4]
  assign _T_98108 = $signed(buffer_13_686) + $signed(buffer_13_687); // @[Modules.scala 63:156:@52017.4]
  assign _T_98109 = _T_98108[10:0]; // @[Modules.scala 63:156:@52018.4]
  assign buffer_13_736 = $signed(_T_98109); // @[Modules.scala 63:156:@52019.4]
  assign _T_98111 = $signed(buffer_13_736) + $signed(buffer_13_688); // @[Modules.scala 63:156:@52021.4]
  assign _T_98112 = _T_98111[10:0]; // @[Modules.scala 63:156:@52022.4]
  assign buffer_13_737 = $signed(_T_98112); // @[Modules.scala 63:156:@52023.4]
  assign _T_98114 = $signed(buffer_13_737) + $signed(buffer_13_689); // @[Modules.scala 63:156:@52025.4]
  assign _T_98115 = _T_98114[10:0]; // @[Modules.scala 63:156:@52026.4]
  assign buffer_13_738 = $signed(_T_98115); // @[Modules.scala 63:156:@52027.4]
  assign _T_98117 = $signed(buffer_13_738) + $signed(buffer_13_690); // @[Modules.scala 63:156:@52029.4]
  assign _T_98118 = _T_98117[10:0]; // @[Modules.scala 63:156:@52030.4]
  assign buffer_13_739 = $signed(_T_98118); // @[Modules.scala 63:156:@52031.4]
  assign _T_98120 = $signed(buffer_13_739) + $signed(buffer_13_691); // @[Modules.scala 63:156:@52033.4]
  assign _T_98121 = _T_98120[10:0]; // @[Modules.scala 63:156:@52034.4]
  assign buffer_13_740 = $signed(_T_98121); // @[Modules.scala 63:156:@52035.4]
  assign _T_98123 = $signed(buffer_13_740) + $signed(buffer_13_692); // @[Modules.scala 63:156:@52037.4]
  assign _T_98124 = _T_98123[10:0]; // @[Modules.scala 63:156:@52038.4]
  assign buffer_13_741 = $signed(_T_98124); // @[Modules.scala 63:156:@52039.4]
  assign _T_98126 = $signed(buffer_13_741) + $signed(buffer_13_693); // @[Modules.scala 63:156:@52041.4]
  assign _T_98127 = _T_98126[10:0]; // @[Modules.scala 63:156:@52042.4]
  assign buffer_13_742 = $signed(_T_98127); // @[Modules.scala 63:156:@52043.4]
  assign _T_98129 = $signed(buffer_13_742) + $signed(buffer_13_694); // @[Modules.scala 63:156:@52045.4]
  assign _T_98130 = _T_98129[10:0]; // @[Modules.scala 63:156:@52046.4]
  assign buffer_13_743 = $signed(_T_98130); // @[Modules.scala 63:156:@52047.4]
  assign _T_98132 = $signed(buffer_13_743) + $signed(buffer_13_695); // @[Modules.scala 63:156:@52049.4]
  assign _T_98133 = _T_98132[10:0]; // @[Modules.scala 63:156:@52050.4]
  assign buffer_13_744 = $signed(_T_98133); // @[Modules.scala 63:156:@52051.4]
  assign _T_98135 = $signed(buffer_13_744) + $signed(buffer_13_696); // @[Modules.scala 63:156:@52053.4]
  assign _T_98136 = _T_98135[10:0]; // @[Modules.scala 63:156:@52054.4]
  assign buffer_13_745 = $signed(_T_98136); // @[Modules.scala 63:156:@52055.4]
  assign _T_98138 = $signed(buffer_13_745) + $signed(buffer_13_697); // @[Modules.scala 63:156:@52057.4]
  assign _T_98139 = _T_98138[10:0]; // @[Modules.scala 63:156:@52058.4]
  assign buffer_13_746 = $signed(_T_98139); // @[Modules.scala 63:156:@52059.4]
  assign _T_98141 = $signed(buffer_13_746) + $signed(buffer_13_698); // @[Modules.scala 63:156:@52061.4]
  assign _T_98142 = _T_98141[10:0]; // @[Modules.scala 63:156:@52062.4]
  assign buffer_13_747 = $signed(_T_98142); // @[Modules.scala 63:156:@52063.4]
  assign _T_98144 = $signed(buffer_13_747) + $signed(buffer_13_699); // @[Modules.scala 63:156:@52065.4]
  assign _T_98145 = _T_98144[10:0]; // @[Modules.scala 63:156:@52066.4]
  assign buffer_13_748 = $signed(_T_98145); // @[Modules.scala 63:156:@52067.4]
  assign _T_98147 = $signed(buffer_13_748) + $signed(buffer_13_700); // @[Modules.scala 63:156:@52069.4]
  assign _T_98148 = _T_98147[10:0]; // @[Modules.scala 63:156:@52070.4]
  assign buffer_13_749 = $signed(_T_98148); // @[Modules.scala 63:156:@52071.4]
  assign _T_98150 = $signed(buffer_13_749) + $signed(buffer_13_701); // @[Modules.scala 63:156:@52073.4]
  assign _T_98151 = _T_98150[10:0]; // @[Modules.scala 63:156:@52074.4]
  assign buffer_13_750 = $signed(_T_98151); // @[Modules.scala 63:156:@52075.4]
  assign _T_98153 = $signed(buffer_13_750) + $signed(buffer_13_702); // @[Modules.scala 63:156:@52077.4]
  assign _T_98154 = _T_98153[10:0]; // @[Modules.scala 63:156:@52078.4]
  assign buffer_13_751 = $signed(_T_98154); // @[Modules.scala 63:156:@52079.4]
  assign _T_98156 = $signed(buffer_13_751) + $signed(buffer_13_703); // @[Modules.scala 63:156:@52081.4]
  assign _T_98157 = _T_98156[10:0]; // @[Modules.scala 63:156:@52082.4]
  assign buffer_13_752 = $signed(_T_98157); // @[Modules.scala 63:156:@52083.4]
  assign _T_98159 = $signed(buffer_13_752) + $signed(buffer_13_704); // @[Modules.scala 63:156:@52085.4]
  assign _T_98160 = _T_98159[10:0]; // @[Modules.scala 63:156:@52086.4]
  assign buffer_13_753 = $signed(_T_98160); // @[Modules.scala 63:156:@52087.4]
  assign _T_98162 = $signed(buffer_13_753) + $signed(buffer_13_705); // @[Modules.scala 63:156:@52089.4]
  assign _T_98163 = _T_98162[10:0]; // @[Modules.scala 63:156:@52090.4]
  assign buffer_13_754 = $signed(_T_98163); // @[Modules.scala 63:156:@52091.4]
  assign _T_98165 = $signed(buffer_13_754) + $signed(buffer_13_706); // @[Modules.scala 63:156:@52093.4]
  assign _T_98166 = _T_98165[10:0]; // @[Modules.scala 63:156:@52094.4]
  assign buffer_13_755 = $signed(_T_98166); // @[Modules.scala 63:156:@52095.4]
  assign _T_98168 = $signed(buffer_13_755) + $signed(buffer_13_707); // @[Modules.scala 63:156:@52097.4]
  assign _T_98169 = _T_98168[10:0]; // @[Modules.scala 63:156:@52098.4]
  assign buffer_13_756 = $signed(_T_98169); // @[Modules.scala 63:156:@52099.4]
  assign _T_98171 = $signed(buffer_13_756) + $signed(buffer_13_708); // @[Modules.scala 63:156:@52101.4]
  assign _T_98172 = _T_98171[10:0]; // @[Modules.scala 63:156:@52102.4]
  assign buffer_13_757 = $signed(_T_98172); // @[Modules.scala 63:156:@52103.4]
  assign _T_98174 = $signed(buffer_13_757) + $signed(buffer_13_709); // @[Modules.scala 63:156:@52105.4]
  assign _T_98175 = _T_98174[10:0]; // @[Modules.scala 63:156:@52106.4]
  assign buffer_13_758 = $signed(_T_98175); // @[Modules.scala 63:156:@52107.4]
  assign _T_98177 = $signed(buffer_13_758) + $signed(buffer_13_710); // @[Modules.scala 63:156:@52109.4]
  assign _T_98178 = _T_98177[10:0]; // @[Modules.scala 63:156:@52110.4]
  assign buffer_13_759 = $signed(_T_98178); // @[Modules.scala 63:156:@52111.4]
  assign _T_98180 = $signed(buffer_13_759) + $signed(buffer_13_711); // @[Modules.scala 63:156:@52113.4]
  assign _T_98181 = _T_98180[10:0]; // @[Modules.scala 63:156:@52114.4]
  assign buffer_13_760 = $signed(_T_98181); // @[Modules.scala 63:156:@52115.4]
  assign _T_98183 = $signed(buffer_13_760) + $signed(buffer_13_712); // @[Modules.scala 63:156:@52117.4]
  assign _T_98184 = _T_98183[10:0]; // @[Modules.scala 63:156:@52118.4]
  assign buffer_13_761 = $signed(_T_98184); // @[Modules.scala 63:156:@52119.4]
  assign _T_98186 = $signed(buffer_13_761) + $signed(buffer_13_713); // @[Modules.scala 63:156:@52121.4]
  assign _T_98187 = _T_98186[10:0]; // @[Modules.scala 63:156:@52122.4]
  assign buffer_13_762 = $signed(_T_98187); // @[Modules.scala 63:156:@52123.4]
  assign _T_98189 = $signed(buffer_13_762) + $signed(buffer_13_714); // @[Modules.scala 63:156:@52125.4]
  assign _T_98190 = _T_98189[10:0]; // @[Modules.scala 63:156:@52126.4]
  assign buffer_13_763 = $signed(_T_98190); // @[Modules.scala 63:156:@52127.4]
  assign _T_98192 = $signed(buffer_13_763) + $signed(buffer_13_715); // @[Modules.scala 63:156:@52129.4]
  assign _T_98193 = _T_98192[10:0]; // @[Modules.scala 63:156:@52130.4]
  assign buffer_13_764 = $signed(_T_98193); // @[Modules.scala 63:156:@52131.4]
  assign _T_98195 = $signed(buffer_13_764) + $signed(buffer_13_716); // @[Modules.scala 63:156:@52133.4]
  assign _T_98196 = _T_98195[10:0]; // @[Modules.scala 63:156:@52134.4]
  assign buffer_13_765 = $signed(_T_98196); // @[Modules.scala 63:156:@52135.4]
  assign _T_98198 = $signed(buffer_13_765) + $signed(buffer_13_717); // @[Modules.scala 63:156:@52137.4]
  assign _T_98199 = _T_98198[10:0]; // @[Modules.scala 63:156:@52138.4]
  assign buffer_13_766 = $signed(_T_98199); // @[Modules.scala 63:156:@52139.4]
  assign _T_98201 = $signed(buffer_13_766) + $signed(buffer_13_718); // @[Modules.scala 63:156:@52141.4]
  assign _T_98202 = _T_98201[10:0]; // @[Modules.scala 63:156:@52142.4]
  assign buffer_13_767 = $signed(_T_98202); // @[Modules.scala 63:156:@52143.4]
  assign _T_98204 = $signed(buffer_13_767) + $signed(buffer_13_719); // @[Modules.scala 63:156:@52145.4]
  assign _T_98205 = _T_98204[10:0]; // @[Modules.scala 63:156:@52146.4]
  assign buffer_13_768 = $signed(_T_98205); // @[Modules.scala 63:156:@52147.4]
  assign _T_98207 = $signed(buffer_13_768) + $signed(buffer_13_720); // @[Modules.scala 63:156:@52149.4]
  assign _T_98208 = _T_98207[10:0]; // @[Modules.scala 63:156:@52150.4]
  assign buffer_13_769 = $signed(_T_98208); // @[Modules.scala 63:156:@52151.4]
  assign _T_98210 = $signed(buffer_13_769) + $signed(buffer_13_721); // @[Modules.scala 63:156:@52153.4]
  assign _T_98211 = _T_98210[10:0]; // @[Modules.scala 63:156:@52154.4]
  assign buffer_13_770 = $signed(_T_98211); // @[Modules.scala 63:156:@52155.4]
  assign _T_98213 = $signed(buffer_13_770) + $signed(buffer_13_722); // @[Modules.scala 63:156:@52157.4]
  assign _T_98214 = _T_98213[10:0]; // @[Modules.scala 63:156:@52158.4]
  assign buffer_13_771 = $signed(_T_98214); // @[Modules.scala 63:156:@52159.4]
  assign _T_98216 = $signed(buffer_13_771) + $signed(buffer_13_723); // @[Modules.scala 63:156:@52161.4]
  assign _T_98217 = _T_98216[10:0]; // @[Modules.scala 63:156:@52162.4]
  assign buffer_13_772 = $signed(_T_98217); // @[Modules.scala 63:156:@52163.4]
  assign _T_98219 = $signed(buffer_13_772) + $signed(buffer_13_724); // @[Modules.scala 63:156:@52165.4]
  assign _T_98220 = _T_98219[10:0]; // @[Modules.scala 63:156:@52166.4]
  assign buffer_13_773 = $signed(_T_98220); // @[Modules.scala 63:156:@52167.4]
  assign _T_98222 = $signed(buffer_13_773) + $signed(buffer_13_725); // @[Modules.scala 63:156:@52169.4]
  assign _T_98223 = _T_98222[10:0]; // @[Modules.scala 63:156:@52170.4]
  assign buffer_13_774 = $signed(_T_98223); // @[Modules.scala 63:156:@52171.4]
  assign _T_98225 = $signed(buffer_13_774) + $signed(buffer_13_726); // @[Modules.scala 63:156:@52173.4]
  assign _T_98226 = _T_98225[10:0]; // @[Modules.scala 63:156:@52174.4]
  assign buffer_13_775 = $signed(_T_98226); // @[Modules.scala 63:156:@52175.4]
  assign _T_98228 = $signed(buffer_13_775) + $signed(buffer_13_727); // @[Modules.scala 63:156:@52177.4]
  assign _T_98229 = _T_98228[10:0]; // @[Modules.scala 63:156:@52178.4]
  assign buffer_13_776 = $signed(_T_98229); // @[Modules.scala 63:156:@52179.4]
  assign _T_98231 = $signed(buffer_13_776) + $signed(buffer_13_728); // @[Modules.scala 63:156:@52181.4]
  assign _T_98232 = _T_98231[10:0]; // @[Modules.scala 63:156:@52182.4]
  assign buffer_13_777 = $signed(_T_98232); // @[Modules.scala 63:156:@52183.4]
  assign _T_98234 = $signed(buffer_13_777) + $signed(buffer_13_729); // @[Modules.scala 63:156:@52185.4]
  assign _T_98235 = _T_98234[10:0]; // @[Modules.scala 63:156:@52186.4]
  assign buffer_13_778 = $signed(_T_98235); // @[Modules.scala 63:156:@52187.4]
  assign _T_98237 = $signed(buffer_13_778) + $signed(buffer_2_730); // @[Modules.scala 63:156:@52189.4]
  assign _T_98238 = _T_98237[10:0]; // @[Modules.scala 63:156:@52190.4]
  assign buffer_13_779 = $signed(_T_98238); // @[Modules.scala 63:156:@52191.4]
  assign _T_98240 = $signed(buffer_13_779) + $signed(buffer_13_731); // @[Modules.scala 63:156:@52193.4]
  assign _T_98241 = _T_98240[10:0]; // @[Modules.scala 63:156:@52194.4]
  assign buffer_13_780 = $signed(_T_98241); // @[Modules.scala 63:156:@52195.4]
  assign _T_98243 = $signed(buffer_13_780) + $signed(buffer_4_732); // @[Modules.scala 63:156:@52197.4]
  assign _T_98244 = _T_98243[10:0]; // @[Modules.scala 63:156:@52198.4]
  assign buffer_13_781 = $signed(_T_98244); // @[Modules.scala 63:156:@52199.4]
  assign _T_98246 = $signed(buffer_13_781) + $signed(buffer_13_733); // @[Modules.scala 63:156:@52201.4]
  assign _T_98247 = _T_98246[10:0]; // @[Modules.scala 63:156:@52202.4]
  assign buffer_13_782 = $signed(_T_98247); // @[Modules.scala 63:156:@52203.4]
  assign _T_98249 = $signed(buffer_13_782) + $signed(buffer_13_734); // @[Modules.scala 63:156:@52205.4]
  assign _T_98250 = _T_98249[10:0]; // @[Modules.scala 63:156:@52206.4]
  assign buffer_13_783 = $signed(_T_98250); // @[Modules.scala 63:156:@52207.4]
  assign _T_98414 = $signed(io_in_60) - $signed(io_in_61); // @[Modules.scala 40:46:@52384.4]
  assign _T_98415 = _T_98414[4:0]; // @[Modules.scala 40:46:@52385.4]
  assign _T_98416 = $signed(_T_98415); // @[Modules.scala 40:46:@52386.4]
  assign _T_98499 = $signed(_T_64143) + $signed(io_in_91); // @[Modules.scala 43:47:@52474.4]
  assign _T_98500 = _T_98499[4:0]; // @[Modules.scala 43:47:@52475.4]
  assign _T_98501 = $signed(_T_98500); // @[Modules.scala 43:47:@52476.4]
  assign _T_98508 = $signed(io_in_96) - $signed(io_in_97); // @[Modules.scala 40:46:@52486.4]
  assign _T_98509 = _T_98508[4:0]; // @[Modules.scala 40:46:@52487.4]
  assign _T_98510 = $signed(_T_98509); // @[Modules.scala 40:46:@52488.4]
  assign _T_98630 = $signed(_T_60981) - $signed(io_in_141); // @[Modules.scala 46:47:@52616.4]
  assign _T_98631 = _T_98630[4:0]; // @[Modules.scala 46:47:@52617.4]
  assign _T_98632 = $signed(_T_98631); // @[Modules.scala 46:47:@52618.4]
  assign _T_98712 = $signed(_T_54753) + $signed(io_in_177); // @[Modules.scala 43:47:@52709.4]
  assign _T_98713 = _T_98712[4:0]; // @[Modules.scala 43:47:@52710.4]
  assign _T_98714 = $signed(_T_98713); // @[Modules.scala 43:47:@52711.4]
  assign _T_98934 = $signed(_T_55047) + $signed(io_in_269); // @[Modules.scala 43:47:@52956.4]
  assign _T_98935 = _T_98934[4:0]; // @[Modules.scala 43:47:@52957.4]
  assign _T_98936 = $signed(_T_98935); // @[Modules.scala 43:47:@52958.4]
  assign _T_99080 = $signed(io_in_328) - $signed(io_in_329); // @[Modules.scala 40:46:@53118.4]
  assign _T_99081 = _T_99080[4:0]; // @[Modules.scala 40:46:@53119.4]
  assign _T_99082 = $signed(_T_99081); // @[Modules.scala 40:46:@53120.4]
  assign _T_99127 = $signed(io_in_346) - $signed(io_in_347); // @[Modules.scala 40:46:@53169.4]
  assign _T_99128 = _T_99127[4:0]; // @[Modules.scala 40:46:@53170.4]
  assign _T_99129 = $signed(_T_99128); // @[Modules.scala 40:46:@53171.4]
  assign _T_99156 = $signed(io_in_360) - $signed(io_in_361); // @[Modules.scala 40:46:@53203.4]
  assign _T_99157 = _T_99156[4:0]; // @[Modules.scala 40:46:@53204.4]
  assign _T_99158 = $signed(_T_99157); // @[Modules.scala 40:46:@53205.4]
  assign _T_99349 = $signed(io_in_430) - $signed(io_in_431); // @[Modules.scala 40:46:@53409.4]
  assign _T_99350 = _T_99349[4:0]; // @[Modules.scala 40:46:@53410.4]
  assign _T_99351 = $signed(_T_99350); // @[Modules.scala 40:46:@53411.4]
  assign _T_99356 = $signed(_T_58614) + $signed(io_in_433); // @[Modules.scala 43:47:@53416.4]
  assign _T_99357 = _T_99356[4:0]; // @[Modules.scala 43:47:@53417.4]
  assign _T_99358 = $signed(_T_99357); // @[Modules.scala 43:47:@53418.4]
  assign _T_99640 = $signed(io_in_568) - $signed(io_in_569); // @[Modules.scala 40:46:@53748.4]
  assign _T_99641 = _T_99640[4:0]; // @[Modules.scala 40:46:@53749.4]
  assign _T_99642 = $signed(_T_99641); // @[Modules.scala 40:46:@53750.4]
  assign _T_99942 = $signed(_T_59244) + $signed(io_in_709); // @[Modules.scala 43:47:@54097.4]
  assign _T_99943 = _T_99942[4:0]; // @[Modules.scala 43:47:@54098.4]
  assign _T_99944 = $signed(_T_99943); // @[Modules.scala 43:47:@54099.4]
  assign _T_99973 = $signed(_T_56226) + $signed(io_in_727); // @[Modules.scala 43:47:@54136.4]
  assign _T_99974 = _T_99973[4:0]; // @[Modules.scala 43:47:@54137.4]
  assign _T_99975 = $signed(_T_99974); // @[Modules.scala 43:47:@54138.4]
  assign _T_99997 = $signed(_T_59319) + $signed(io_in_735); // @[Modules.scala 43:47:@54161.4]
  assign _T_99998 = _T_99997[4:0]; // @[Modules.scala 43:47:@54162.4]
  assign _T_99999 = $signed(_T_99998); // @[Modules.scala 43:47:@54163.4]
  assign _T_100000 = $signed(io_in_736) - $signed(io_in_737); // @[Modules.scala 40:46:@54165.4]
  assign _T_100001 = _T_100000[4:0]; // @[Modules.scala 40:46:@54166.4]
  assign _T_100002 = $signed(_T_100001); // @[Modules.scala 40:46:@54167.4]
  assign _T_100003 = $signed(io_in_738) - $signed(io_in_739); // @[Modules.scala 40:46:@54169.4]
  assign _T_100004 = _T_100003[4:0]; // @[Modules.scala 40:46:@54170.4]
  assign _T_100005 = $signed(_T_100004); // @[Modules.scala 40:46:@54171.4]
  assign _T_100116 = $signed(buffer_0_0) + $signed(buffer_3_1); // @[Modules.scala 50:57:@54294.4]
  assign _T_100117 = _T_100116[10:0]; // @[Modules.scala 50:57:@54295.4]
  assign buffer_14_392 = $signed(_T_100117); // @[Modules.scala 50:57:@54296.4]
  assign _T_100122 = $signed(buffer_0_4) + $signed(buffer_4_5); // @[Modules.scala 50:57:@54302.4]
  assign _T_100123 = _T_100122[10:0]; // @[Modules.scala 50:57:@54303.4]
  assign buffer_14_394 = $signed(_T_100123); // @[Modules.scala 50:57:@54304.4]
  assign _T_100137 = $signed(buffer_3_14) + $signed(buffer_2_15); // @[Modules.scala 50:57:@54322.4]
  assign _T_100138 = _T_100137[10:0]; // @[Modules.scala 50:57:@54323.4]
  assign buffer_14_399 = $signed(_T_100138); // @[Modules.scala 50:57:@54324.4]
  assign _T_100146 = $signed(buffer_0_20) + $signed(buffer_1_21); // @[Modules.scala 50:57:@54334.4]
  assign _T_100147 = _T_100146[10:0]; // @[Modules.scala 50:57:@54335.4]
  assign buffer_14_402 = $signed(_T_100147); // @[Modules.scala 50:57:@54336.4]
  assign _T_100155 = $signed(buffer_1_26) + $signed(buffer_7_27); // @[Modules.scala 50:57:@54346.4]
  assign _T_100156 = _T_100155[10:0]; // @[Modules.scala 50:57:@54347.4]
  assign buffer_14_405 = $signed(_T_100156); // @[Modules.scala 50:57:@54348.4]
  assign buffer_14_30 = {{6{_T_98416[4]}},_T_98416}; // @[Modules.scala 32:22:@8.4]
  assign _T_100161 = $signed(buffer_14_30) + $signed(buffer_1_31); // @[Modules.scala 50:57:@54354.4]
  assign _T_100162 = _T_100161[10:0]; // @[Modules.scala 50:57:@54355.4]
  assign buffer_14_407 = $signed(_T_100162); // @[Modules.scala 50:57:@54356.4]
  assign _T_100179 = $signed(buffer_5_42) + $signed(buffer_1_43); // @[Modules.scala 50:57:@54378.4]
  assign _T_100180 = _T_100179[10:0]; // @[Modules.scala 50:57:@54379.4]
  assign buffer_14_413 = $signed(_T_100180); // @[Modules.scala 50:57:@54380.4]
  assign buffer_14_45 = {{6{_T_98501[4]}},_T_98501}; // @[Modules.scala 32:22:@8.4]
  assign _T_100182 = $signed(buffer_2_44) + $signed(buffer_14_45); // @[Modules.scala 50:57:@54382.4]
  assign _T_100183 = _T_100182[10:0]; // @[Modules.scala 50:57:@54383.4]
  assign buffer_14_414 = $signed(_T_100183); // @[Modules.scala 50:57:@54384.4]
  assign buffer_14_48 = {{6{_T_98510[4]}},_T_98510}; // @[Modules.scala 32:22:@8.4]
  assign _T_100188 = $signed(buffer_14_48) + $signed(buffer_2_49); // @[Modules.scala 50:57:@54390.4]
  assign _T_100189 = _T_100188[10:0]; // @[Modules.scala 50:57:@54391.4]
  assign buffer_14_416 = $signed(_T_100189); // @[Modules.scala 50:57:@54392.4]
  assign _T_100200 = $signed(buffer_3_56) + $signed(buffer_0_57); // @[Modules.scala 50:57:@54406.4]
  assign _T_100201 = _T_100200[10:0]; // @[Modules.scala 50:57:@54407.4]
  assign buffer_14_420 = $signed(_T_100201); // @[Modules.scala 50:57:@54408.4]
  assign _T_100209 = $signed(buffer_3_62) + $signed(buffer_0_63); // @[Modules.scala 50:57:@54418.4]
  assign _T_100210 = _T_100209[10:0]; // @[Modules.scala 50:57:@54419.4]
  assign buffer_14_423 = $signed(_T_100210); // @[Modules.scala 50:57:@54420.4]
  assign buffer_14_70 = {{6{_T_98632[4]}},_T_98632}; // @[Modules.scala 32:22:@8.4]
  assign _T_100221 = $signed(buffer_14_70) + $signed(buffer_5_71); // @[Modules.scala 50:57:@54434.4]
  assign _T_100222 = _T_100221[10:0]; // @[Modules.scala 50:57:@54435.4]
  assign buffer_14_427 = $signed(_T_100222); // @[Modules.scala 50:57:@54436.4]
  assign buffer_14_88 = {{6{_T_98714[4]}},_T_98714}; // @[Modules.scala 32:22:@8.4]
  assign _T_100248 = $signed(buffer_14_88) + $signed(buffer_0_89); // @[Modules.scala 50:57:@54470.4]
  assign _T_100249 = _T_100248[10:0]; // @[Modules.scala 50:57:@54471.4]
  assign buffer_14_436 = $signed(_T_100249); // @[Modules.scala 50:57:@54472.4]
  assign _T_100254 = $signed(buffer_5_92) + $signed(buffer_0_93); // @[Modules.scala 50:57:@54478.4]
  assign _T_100255 = _T_100254[10:0]; // @[Modules.scala 50:57:@54479.4]
  assign buffer_14_438 = $signed(_T_100255); // @[Modules.scala 50:57:@54480.4]
  assign _T_100257 = $signed(buffer_4_94) + $signed(buffer_5_95); // @[Modules.scala 50:57:@54482.4]
  assign _T_100258 = _T_100257[10:0]; // @[Modules.scala 50:57:@54483.4]
  assign buffer_14_439 = $signed(_T_100258); // @[Modules.scala 50:57:@54484.4]
  assign _T_100296 = $signed(buffer_1_120) + $signed(buffer_6_121); // @[Modules.scala 50:57:@54534.4]
  assign _T_100297 = _T_100296[10:0]; // @[Modules.scala 50:57:@54535.4]
  assign buffer_14_452 = $signed(_T_100297); // @[Modules.scala 50:57:@54536.4]
  assign buffer_14_134 = {{6{_T_98936[4]}},_T_98936}; // @[Modules.scala 32:22:@8.4]
  assign _T_100317 = $signed(buffer_14_134) + $signed(buffer_3_135); // @[Modules.scala 50:57:@54562.4]
  assign _T_100318 = _T_100317[10:0]; // @[Modules.scala 50:57:@54563.4]
  assign buffer_14_459 = $signed(_T_100318); // @[Modules.scala 50:57:@54564.4]
  assign _T_100320 = $signed(buffer_5_136) + $signed(buffer_1_137); // @[Modules.scala 50:57:@54566.4]
  assign _T_100321 = _T_100320[10:0]; // @[Modules.scala 50:57:@54567.4]
  assign buffer_14_460 = $signed(_T_100321); // @[Modules.scala 50:57:@54568.4]
  assign _T_100323 = $signed(buffer_1_138) + $signed(buffer_5_139); // @[Modules.scala 50:57:@54570.4]
  assign _T_100324 = _T_100323[10:0]; // @[Modules.scala 50:57:@54571.4]
  assign buffer_14_461 = $signed(_T_100324); // @[Modules.scala 50:57:@54572.4]
  assign buffer_14_164 = {{6{_T_99082[4]}},_T_99082}; // @[Modules.scala 32:22:@8.4]
  assign _T_100362 = $signed(buffer_14_164) + $signed(buffer_5_165); // @[Modules.scala 50:57:@54622.4]
  assign _T_100363 = _T_100362[10:0]; // @[Modules.scala 50:57:@54623.4]
  assign buffer_14_474 = $signed(_T_100363); // @[Modules.scala 50:57:@54624.4]
  assign _T_100371 = $signed(buffer_0_170) + $signed(buffer_3_171); // @[Modules.scala 50:57:@54634.4]
  assign _T_100372 = _T_100371[10:0]; // @[Modules.scala 50:57:@54635.4]
  assign buffer_14_477 = $signed(_T_100372); // @[Modules.scala 50:57:@54636.4]
  assign buffer_14_173 = {{6{_T_99129[4]}},_T_99129}; // @[Modules.scala 32:22:@8.4]
  assign _T_100374 = $signed(buffer_3_172) + $signed(buffer_14_173); // @[Modules.scala 50:57:@54638.4]
  assign _T_100375 = _T_100374[10:0]; // @[Modules.scala 50:57:@54639.4]
  assign buffer_14_478 = $signed(_T_100375); // @[Modules.scala 50:57:@54640.4]
  assign buffer_14_180 = {{6{_T_99158[4]}},_T_99158}; // @[Modules.scala 32:22:@8.4]
  assign _T_100386 = $signed(buffer_14_180) + $signed(buffer_2_181); // @[Modules.scala 50:57:@54654.4]
  assign _T_100387 = _T_100386[10:0]; // @[Modules.scala 50:57:@54655.4]
  assign buffer_14_482 = $signed(_T_100387); // @[Modules.scala 50:57:@54656.4]
  assign _T_100392 = $signed(buffer_1_184) + $signed(buffer_11_185); // @[Modules.scala 50:57:@54662.4]
  assign _T_100393 = _T_100392[10:0]; // @[Modules.scala 50:57:@54663.4]
  assign buffer_14_484 = $signed(_T_100393); // @[Modules.scala 50:57:@54664.4]
  assign _T_100395 = $signed(buffer_11_186) + $signed(buffer_3_187); // @[Modules.scala 50:57:@54666.4]
  assign _T_100396 = _T_100395[10:0]; // @[Modules.scala 50:57:@54667.4]
  assign buffer_14_485 = $signed(_T_100396); // @[Modules.scala 50:57:@54668.4]
  assign _T_100404 = $signed(buffer_0_192) + $signed(buffer_2_193); // @[Modules.scala 50:57:@54678.4]
  assign _T_100405 = _T_100404[10:0]; // @[Modules.scala 50:57:@54679.4]
  assign buffer_14_488 = $signed(_T_100405); // @[Modules.scala 50:57:@54680.4]
  assign _T_100428 = $signed(buffer_2_208) + $signed(buffer_4_209); // @[Modules.scala 50:57:@54710.4]
  assign _T_100429 = _T_100428[10:0]; // @[Modules.scala 50:57:@54711.4]
  assign buffer_14_496 = $signed(_T_100429); // @[Modules.scala 50:57:@54712.4]
  assign buffer_14_215 = {{6{_T_99351[4]}},_T_99351}; // @[Modules.scala 32:22:@8.4]
  assign _T_100437 = $signed(buffer_0_214) + $signed(buffer_14_215); // @[Modules.scala 50:57:@54722.4]
  assign _T_100438 = _T_100437[10:0]; // @[Modules.scala 50:57:@54723.4]
  assign buffer_14_499 = $signed(_T_100438); // @[Modules.scala 50:57:@54724.4]
  assign buffer_14_216 = {{6{_T_99358[4]}},_T_99358}; // @[Modules.scala 32:22:@8.4]
  assign _T_100440 = $signed(buffer_14_216) + $signed(buffer_1_217); // @[Modules.scala 50:57:@54726.4]
  assign _T_100441 = _T_100440[10:0]; // @[Modules.scala 50:57:@54727.4]
  assign buffer_14_500 = $signed(_T_100441); // @[Modules.scala 50:57:@54728.4]
  assign _T_100443 = $signed(buffer_4_218) + $signed(buffer_2_219); // @[Modules.scala 50:57:@54730.4]
  assign _T_100444 = _T_100443[10:0]; // @[Modules.scala 50:57:@54731.4]
  assign buffer_14_501 = $signed(_T_100444); // @[Modules.scala 50:57:@54732.4]
  assign _T_100464 = $signed(buffer_1_232) + $signed(buffer_6_233); // @[Modules.scala 50:57:@54758.4]
  assign _T_100465 = _T_100464[10:0]; // @[Modules.scala 50:57:@54759.4]
  assign buffer_14_508 = $signed(_T_100465); // @[Modules.scala 50:57:@54760.4]
  assign _T_100467 = $signed(buffer_2_234) + $signed(buffer_6_235); // @[Modules.scala 50:57:@54762.4]
  assign _T_100468 = _T_100467[10:0]; // @[Modules.scala 50:57:@54763.4]
  assign buffer_14_509 = $signed(_T_100468); // @[Modules.scala 50:57:@54764.4]
  assign _T_100470 = $signed(buffer_0_236) + $signed(buffer_3_237); // @[Modules.scala 50:57:@54766.4]
  assign _T_100471 = _T_100470[10:0]; // @[Modules.scala 50:57:@54767.4]
  assign buffer_14_510 = $signed(_T_100471); // @[Modules.scala 50:57:@54768.4]
  assign _T_100473 = $signed(buffer_12_238) + $signed(buffer_1_239); // @[Modules.scala 50:57:@54770.4]
  assign _T_100474 = _T_100473[10:0]; // @[Modules.scala 50:57:@54771.4]
  assign buffer_14_511 = $signed(_T_100474); // @[Modules.scala 50:57:@54772.4]
  assign _T_100482 = $signed(buffer_12_244) + $signed(buffer_1_245); // @[Modules.scala 50:57:@54782.4]
  assign _T_100483 = _T_100482[10:0]; // @[Modules.scala 50:57:@54783.4]
  assign buffer_14_514 = $signed(_T_100483); // @[Modules.scala 50:57:@54784.4]
  assign _T_100488 = $signed(buffer_13_248) + $signed(buffer_0_249); // @[Modules.scala 50:57:@54790.4]
  assign _T_100489 = _T_100488[10:0]; // @[Modules.scala 50:57:@54791.4]
  assign buffer_14_516 = $signed(_T_100489); // @[Modules.scala 50:57:@54792.4]
  assign _T_100494 = $signed(buffer_3_252) + $signed(buffer_0_253); // @[Modules.scala 50:57:@54798.4]
  assign _T_100495 = _T_100494[10:0]; // @[Modules.scala 50:57:@54799.4]
  assign buffer_14_518 = $signed(_T_100495); // @[Modules.scala 50:57:@54800.4]
  assign _T_100503 = $signed(buffer_1_258) + $signed(buffer_4_259); // @[Modules.scala 50:57:@54810.4]
  assign _T_100504 = _T_100503[10:0]; // @[Modules.scala 50:57:@54811.4]
  assign buffer_14_521 = $signed(_T_100504); // @[Modules.scala 50:57:@54812.4]
  assign _T_100515 = $signed(buffer_0_266) + $signed(buffer_1_267); // @[Modules.scala 50:57:@54826.4]
  assign _T_100516 = _T_100515[10:0]; // @[Modules.scala 50:57:@54827.4]
  assign buffer_14_525 = $signed(_T_100516); // @[Modules.scala 50:57:@54828.4]
  assign _T_100521 = $signed(buffer_1_270) + $signed(buffer_3_271); // @[Modules.scala 50:57:@54834.4]
  assign _T_100522 = _T_100521[10:0]; // @[Modules.scala 50:57:@54835.4]
  assign buffer_14_527 = $signed(_T_100522); // @[Modules.scala 50:57:@54836.4]
  assign _T_100536 = $signed(buffer_12_280) + $signed(buffer_1_281); // @[Modules.scala 50:57:@54854.4]
  assign _T_100537 = _T_100536[10:0]; // @[Modules.scala 50:57:@54855.4]
  assign buffer_14_532 = $signed(_T_100537); // @[Modules.scala 50:57:@54856.4]
  assign buffer_14_284 = {{6{_T_99642[4]}},_T_99642}; // @[Modules.scala 32:22:@8.4]
  assign _T_100542 = $signed(buffer_14_284) + $signed(buffer_5_285); // @[Modules.scala 50:57:@54862.4]
  assign _T_100543 = _T_100542[10:0]; // @[Modules.scala 50:57:@54863.4]
  assign buffer_14_534 = $signed(_T_100543); // @[Modules.scala 50:57:@54864.4]
  assign _T_100548 = $signed(buffer_12_288) + $signed(buffer_5_289); // @[Modules.scala 50:57:@54870.4]
  assign _T_100549 = _T_100548[10:0]; // @[Modules.scala 50:57:@54871.4]
  assign buffer_14_536 = $signed(_T_100549); // @[Modules.scala 50:57:@54872.4]
  assign _T_100557 = $signed(buffer_6_294) + $signed(buffer_1_295); // @[Modules.scala 50:57:@54882.4]
  assign _T_100558 = _T_100557[10:0]; // @[Modules.scala 50:57:@54883.4]
  assign buffer_14_539 = $signed(_T_100558); // @[Modules.scala 50:57:@54884.4]
  assign _T_100569 = $signed(buffer_6_302) + $signed(buffer_0_303); // @[Modules.scala 50:57:@54898.4]
  assign _T_100570 = _T_100569[10:0]; // @[Modules.scala 50:57:@54899.4]
  assign buffer_14_543 = $signed(_T_100570); // @[Modules.scala 50:57:@54900.4]
  assign _T_100578 = $signed(buffer_2_308) + $signed(buffer_0_309); // @[Modules.scala 50:57:@54910.4]
  assign _T_100579 = _T_100578[10:0]; // @[Modules.scala 50:57:@54911.4]
  assign buffer_14_546 = $signed(_T_100579); // @[Modules.scala 50:57:@54912.4]
  assign _T_100581 = $signed(buffer_1_310) + $signed(buffer_4_311); // @[Modules.scala 50:57:@54914.4]
  assign _T_100582 = _T_100581[10:0]; // @[Modules.scala 50:57:@54915.4]
  assign buffer_14_547 = $signed(_T_100582); // @[Modules.scala 50:57:@54916.4]
  assign _T_100596 = $signed(buffer_5_320) + $signed(buffer_13_321); // @[Modules.scala 50:57:@54934.4]
  assign _T_100597 = _T_100596[10:0]; // @[Modules.scala 50:57:@54935.4]
  assign buffer_14_552 = $signed(_T_100597); // @[Modules.scala 50:57:@54936.4]
  assign _T_100605 = $signed(buffer_0_326) + $signed(buffer_1_327); // @[Modules.scala 50:57:@54946.4]
  assign _T_100606 = _T_100605[10:0]; // @[Modules.scala 50:57:@54947.4]
  assign buffer_14_555 = $signed(_T_100606); // @[Modules.scala 50:57:@54948.4]
  assign _T_100638 = $signed(buffer_1_348) + $signed(buffer_0_349); // @[Modules.scala 50:57:@54990.4]
  assign _T_100639 = _T_100638[10:0]; // @[Modules.scala 50:57:@54991.4]
  assign buffer_14_566 = $signed(_T_100639); // @[Modules.scala 50:57:@54992.4]
  assign _T_100644 = $signed(buffer_5_352) + $signed(buffer_10_353); // @[Modules.scala 50:57:@54998.4]
  assign _T_100645 = _T_100644[10:0]; // @[Modules.scala 50:57:@54999.4]
  assign buffer_14_568 = $signed(_T_100645); // @[Modules.scala 50:57:@55000.4]
  assign buffer_14_354 = {{6{_T_99944[4]}},_T_99944}; // @[Modules.scala 32:22:@8.4]
  assign _T_100647 = $signed(buffer_14_354) + $signed(buffer_0_355); // @[Modules.scala 50:57:@55002.4]
  assign _T_100648 = _T_100647[10:0]; // @[Modules.scala 50:57:@55003.4]
  assign buffer_14_569 = $signed(_T_100648); // @[Modules.scala 50:57:@55004.4]
  assign _T_100650 = $signed(buffer_9_356) + $signed(buffer_0_357); // @[Modules.scala 50:57:@55006.4]
  assign _T_100651 = _T_100650[10:0]; // @[Modules.scala 50:57:@55007.4]
  assign buffer_14_570 = $signed(_T_100651); // @[Modules.scala 50:57:@55008.4]
  assign buffer_14_363 = {{6{_T_99975[4]}},_T_99975}; // @[Modules.scala 32:22:@8.4]
  assign _T_100659 = $signed(buffer_1_362) + $signed(buffer_14_363); // @[Modules.scala 50:57:@55018.4]
  assign _T_100660 = _T_100659[10:0]; // @[Modules.scala 50:57:@55019.4]
  assign buffer_14_573 = $signed(_T_100660); // @[Modules.scala 50:57:@55020.4]
  assign _T_100662 = $signed(buffer_9_364) + $signed(buffer_0_365); // @[Modules.scala 50:57:@55022.4]
  assign _T_100663 = _T_100662[10:0]; // @[Modules.scala 50:57:@55023.4]
  assign buffer_14_574 = $signed(_T_100663); // @[Modules.scala 50:57:@55024.4]
  assign buffer_14_367 = {{6{_T_99999[4]}},_T_99999}; // @[Modules.scala 32:22:@8.4]
  assign _T_100665 = $signed(buffer_0_366) + $signed(buffer_14_367); // @[Modules.scala 50:57:@55026.4]
  assign _T_100666 = _T_100665[10:0]; // @[Modules.scala 50:57:@55027.4]
  assign buffer_14_575 = $signed(_T_100666); // @[Modules.scala 50:57:@55028.4]
  assign buffer_14_368 = {{6{_T_100002[4]}},_T_100002}; // @[Modules.scala 32:22:@8.4]
  assign buffer_14_369 = {{6{_T_100005[4]}},_T_100005}; // @[Modules.scala 32:22:@8.4]
  assign _T_100668 = $signed(buffer_14_368) + $signed(buffer_14_369); // @[Modules.scala 50:57:@55030.4]
  assign _T_100669 = _T_100668[10:0]; // @[Modules.scala 50:57:@55031.4]
  assign buffer_14_576 = $signed(_T_100669); // @[Modules.scala 50:57:@55032.4]
  assign _T_100671 = $signed(buffer_0_370) + $signed(buffer_5_371); // @[Modules.scala 50:57:@55034.4]
  assign _T_100672 = _T_100671[10:0]; // @[Modules.scala 50:57:@55035.4]
  assign buffer_14_577 = $signed(_T_100672); // @[Modules.scala 50:57:@55036.4]
  assign _T_100701 = $signed(buffer_0_390) + $signed(buffer_1_391); // @[Modules.scala 50:57:@55074.4]
  assign _T_100702 = _T_100701[10:0]; // @[Modules.scala 50:57:@55075.4]
  assign buffer_14_587 = $signed(_T_100702); // @[Modules.scala 50:57:@55076.4]
  assign _T_100704 = $signed(buffer_14_392) + $signed(buffer_7_393); // @[Modules.scala 53:83:@55078.4]
  assign _T_100705 = _T_100704[10:0]; // @[Modules.scala 53:83:@55079.4]
  assign buffer_14_588 = $signed(_T_100705); // @[Modules.scala 53:83:@55080.4]
  assign _T_100707 = $signed(buffer_14_394) + $signed(buffer_0_395); // @[Modules.scala 53:83:@55082.4]
  assign _T_100708 = _T_100707[10:0]; // @[Modules.scala 53:83:@55083.4]
  assign buffer_14_589 = $signed(_T_100708); // @[Modules.scala 53:83:@55084.4]
  assign _T_100710 = $signed(buffer_2_396) + $signed(buffer_7_397); // @[Modules.scala 53:83:@55086.4]
  assign _T_100711 = _T_100710[10:0]; // @[Modules.scala 53:83:@55087.4]
  assign buffer_14_590 = $signed(_T_100711); // @[Modules.scala 53:83:@55088.4]
  assign _T_100713 = $signed(buffer_3_398) + $signed(buffer_14_399); // @[Modules.scala 53:83:@55090.4]
  assign _T_100714 = _T_100713[10:0]; // @[Modules.scala 53:83:@55091.4]
  assign buffer_14_591 = $signed(_T_100714); // @[Modules.scala 53:83:@55092.4]
  assign _T_100716 = $signed(buffer_2_400) + $signed(buffer_0_401); // @[Modules.scala 53:83:@55094.4]
  assign _T_100717 = _T_100716[10:0]; // @[Modules.scala 53:83:@55095.4]
  assign buffer_14_592 = $signed(_T_100717); // @[Modules.scala 53:83:@55096.4]
  assign _T_100719 = $signed(buffer_14_402) + $signed(buffer_4_403); // @[Modules.scala 53:83:@55098.4]
  assign _T_100720 = _T_100719[10:0]; // @[Modules.scala 53:83:@55099.4]
  assign buffer_14_593 = $signed(_T_100720); // @[Modules.scala 53:83:@55100.4]
  assign _T_100722 = $signed(buffer_0_404) + $signed(buffer_14_405); // @[Modules.scala 53:83:@55102.4]
  assign _T_100723 = _T_100722[10:0]; // @[Modules.scala 53:83:@55103.4]
  assign buffer_14_594 = $signed(_T_100723); // @[Modules.scala 53:83:@55104.4]
  assign _T_100725 = $signed(buffer_11_406) + $signed(buffer_14_407); // @[Modules.scala 53:83:@55106.4]
  assign _T_100726 = _T_100725[10:0]; // @[Modules.scala 53:83:@55107.4]
  assign buffer_14_595 = $signed(_T_100726); // @[Modules.scala 53:83:@55108.4]
  assign _T_100734 = $signed(buffer_3_412) + $signed(buffer_14_413); // @[Modules.scala 53:83:@55118.4]
  assign _T_100735 = _T_100734[10:0]; // @[Modules.scala 53:83:@55119.4]
  assign buffer_14_598 = $signed(_T_100735); // @[Modules.scala 53:83:@55120.4]
  assign _T_100737 = $signed(buffer_14_414) + $signed(buffer_1_415); // @[Modules.scala 53:83:@55122.4]
  assign _T_100738 = _T_100737[10:0]; // @[Modules.scala 53:83:@55123.4]
  assign buffer_14_599 = $signed(_T_100738); // @[Modules.scala 53:83:@55124.4]
  assign _T_100740 = $signed(buffer_14_416) + $signed(buffer_6_417); // @[Modules.scala 53:83:@55126.4]
  assign _T_100741 = _T_100740[10:0]; // @[Modules.scala 53:83:@55127.4]
  assign buffer_14_600 = $signed(_T_100741); // @[Modules.scala 53:83:@55128.4]
  assign _T_100743 = $signed(buffer_3_418) + $signed(buffer_6_419); // @[Modules.scala 53:83:@55130.4]
  assign _T_100744 = _T_100743[10:0]; // @[Modules.scala 53:83:@55131.4]
  assign buffer_14_601 = $signed(_T_100744); // @[Modules.scala 53:83:@55132.4]
  assign _T_100746 = $signed(buffer_14_420) + $signed(buffer_5_421); // @[Modules.scala 53:83:@55134.4]
  assign _T_100747 = _T_100746[10:0]; // @[Modules.scala 53:83:@55135.4]
  assign buffer_14_602 = $signed(_T_100747); // @[Modules.scala 53:83:@55136.4]
  assign _T_100749 = $signed(buffer_3_422) + $signed(buffer_14_423); // @[Modules.scala 53:83:@55138.4]
  assign _T_100750 = _T_100749[10:0]; // @[Modules.scala 53:83:@55139.4]
  assign buffer_14_603 = $signed(_T_100750); // @[Modules.scala 53:83:@55140.4]
  assign _T_100752 = $signed(buffer_2_424) + $signed(buffer_4_425); // @[Modules.scala 53:83:@55142.4]
  assign _T_100753 = _T_100752[10:0]; // @[Modules.scala 53:83:@55143.4]
  assign buffer_14_604 = $signed(_T_100753); // @[Modules.scala 53:83:@55144.4]
  assign _T_100755 = $signed(buffer_10_426) + $signed(buffer_14_427); // @[Modules.scala 53:83:@55146.4]
  assign _T_100756 = _T_100755[10:0]; // @[Modules.scala 53:83:@55147.4]
  assign buffer_14_605 = $signed(_T_100756); // @[Modules.scala 53:83:@55148.4]
  assign _T_100758 = $signed(buffer_0_428) + $signed(buffer_3_429); // @[Modules.scala 53:83:@55150.4]
  assign _T_100759 = _T_100758[10:0]; // @[Modules.scala 53:83:@55151.4]
  assign buffer_14_606 = $signed(_T_100759); // @[Modules.scala 53:83:@55152.4]
  assign _T_100764 = $signed(buffer_9_432) + $signed(buffer_5_433); // @[Modules.scala 53:83:@55158.4]
  assign _T_100765 = _T_100764[10:0]; // @[Modules.scala 53:83:@55159.4]
  assign buffer_14_608 = $signed(_T_100765); // @[Modules.scala 53:83:@55160.4]
  assign _T_100767 = $signed(buffer_1_434) + $signed(buffer_2_435); // @[Modules.scala 53:83:@55162.4]
  assign _T_100768 = _T_100767[10:0]; // @[Modules.scala 53:83:@55163.4]
  assign buffer_14_609 = $signed(_T_100768); // @[Modules.scala 53:83:@55164.4]
  assign _T_100770 = $signed(buffer_14_436) + $signed(buffer_5_437); // @[Modules.scala 53:83:@55166.4]
  assign _T_100771 = _T_100770[10:0]; // @[Modules.scala 53:83:@55167.4]
  assign buffer_14_610 = $signed(_T_100771); // @[Modules.scala 53:83:@55168.4]
  assign _T_100773 = $signed(buffer_14_438) + $signed(buffer_14_439); // @[Modules.scala 53:83:@55170.4]
  assign _T_100774 = _T_100773[10:0]; // @[Modules.scala 53:83:@55171.4]
  assign buffer_14_611 = $signed(_T_100774); // @[Modules.scala 53:83:@55172.4]
  assign _T_100779 = $signed(buffer_0_442) + $signed(buffer_5_443); // @[Modules.scala 53:83:@55178.4]
  assign _T_100780 = _T_100779[10:0]; // @[Modules.scala 53:83:@55179.4]
  assign buffer_14_613 = $signed(_T_100780); // @[Modules.scala 53:83:@55180.4]
  assign _T_100782 = $signed(buffer_5_444) + $signed(buffer_3_445); // @[Modules.scala 53:83:@55182.4]
  assign _T_100783 = _T_100782[10:0]; // @[Modules.scala 53:83:@55183.4]
  assign buffer_14_614 = $signed(_T_100783); // @[Modules.scala 53:83:@55184.4]
  assign _T_100785 = $signed(buffer_1_446) + $signed(buffer_2_447); // @[Modules.scala 53:83:@55186.4]
  assign _T_100786 = _T_100785[10:0]; // @[Modules.scala 53:83:@55187.4]
  assign buffer_14_615 = $signed(_T_100786); // @[Modules.scala 53:83:@55188.4]
  assign _T_100791 = $signed(buffer_0_450) + $signed(buffer_3_451); // @[Modules.scala 53:83:@55194.4]
  assign _T_100792 = _T_100791[10:0]; // @[Modules.scala 53:83:@55195.4]
  assign buffer_14_617 = $signed(_T_100792); // @[Modules.scala 53:83:@55196.4]
  assign _T_100794 = $signed(buffer_14_452) + $signed(buffer_4_453); // @[Modules.scala 53:83:@55198.4]
  assign _T_100795 = _T_100794[10:0]; // @[Modules.scala 53:83:@55199.4]
  assign buffer_14_618 = $signed(_T_100795); // @[Modules.scala 53:83:@55200.4]
  assign _T_100803 = $signed(buffer_11_458) + $signed(buffer_14_459); // @[Modules.scala 53:83:@55210.4]
  assign _T_100804 = _T_100803[10:0]; // @[Modules.scala 53:83:@55211.4]
  assign buffer_14_621 = $signed(_T_100804); // @[Modules.scala 53:83:@55212.4]
  assign _T_100806 = $signed(buffer_14_460) + $signed(buffer_14_461); // @[Modules.scala 53:83:@55214.4]
  assign _T_100807 = _T_100806[10:0]; // @[Modules.scala 53:83:@55215.4]
  assign buffer_14_622 = $signed(_T_100807); // @[Modules.scala 53:83:@55216.4]
  assign _T_100812 = $signed(buffer_2_464) + $signed(buffer_7_465); // @[Modules.scala 53:83:@55222.4]
  assign _T_100813 = _T_100812[10:0]; // @[Modules.scala 53:83:@55223.4]
  assign buffer_14_624 = $signed(_T_100813); // @[Modules.scala 53:83:@55224.4]
  assign _T_100815 = $signed(buffer_12_466) + $signed(buffer_9_467); // @[Modules.scala 53:83:@55226.4]
  assign _T_100816 = _T_100815[10:0]; // @[Modules.scala 53:83:@55227.4]
  assign buffer_14_625 = $signed(_T_100816); // @[Modules.scala 53:83:@55228.4]
  assign _T_100824 = $signed(buffer_4_472) + $signed(buffer_12_473); // @[Modules.scala 53:83:@55238.4]
  assign _T_100825 = _T_100824[10:0]; // @[Modules.scala 53:83:@55239.4]
  assign buffer_14_628 = $signed(_T_100825); // @[Modules.scala 53:83:@55240.4]
  assign _T_100827 = $signed(buffer_14_474) + $signed(buffer_1_475); // @[Modules.scala 53:83:@55242.4]
  assign _T_100828 = _T_100827[10:0]; // @[Modules.scala 53:83:@55243.4]
  assign buffer_14_629 = $signed(_T_100828); // @[Modules.scala 53:83:@55244.4]
  assign _T_100830 = $signed(buffer_7_476) + $signed(buffer_14_477); // @[Modules.scala 53:83:@55246.4]
  assign _T_100831 = _T_100830[10:0]; // @[Modules.scala 53:83:@55247.4]
  assign buffer_14_630 = $signed(_T_100831); // @[Modules.scala 53:83:@55248.4]
  assign _T_100833 = $signed(buffer_14_478) + $signed(buffer_0_479); // @[Modules.scala 53:83:@55250.4]
  assign _T_100834 = _T_100833[10:0]; // @[Modules.scala 53:83:@55251.4]
  assign buffer_14_631 = $signed(_T_100834); // @[Modules.scala 53:83:@55252.4]
  assign _T_100839 = $signed(buffer_14_482) + $signed(buffer_4_483); // @[Modules.scala 53:83:@55258.4]
  assign _T_100840 = _T_100839[10:0]; // @[Modules.scala 53:83:@55259.4]
  assign buffer_14_633 = $signed(_T_100840); // @[Modules.scala 53:83:@55260.4]
  assign _T_100842 = $signed(buffer_14_484) + $signed(buffer_14_485); // @[Modules.scala 53:83:@55262.4]
  assign _T_100843 = _T_100842[10:0]; // @[Modules.scala 53:83:@55263.4]
  assign buffer_14_634 = $signed(_T_100843); // @[Modules.scala 53:83:@55264.4]
  assign _T_100845 = $signed(buffer_8_486) + $signed(buffer_4_487); // @[Modules.scala 53:83:@55266.4]
  assign _T_100846 = _T_100845[10:0]; // @[Modules.scala 53:83:@55267.4]
  assign buffer_14_635 = $signed(_T_100846); // @[Modules.scala 53:83:@55268.4]
  assign _T_100848 = $signed(buffer_14_488) + $signed(buffer_3_489); // @[Modules.scala 53:83:@55270.4]
  assign _T_100849 = _T_100848[10:0]; // @[Modules.scala 53:83:@55271.4]
  assign buffer_14_636 = $signed(_T_100849); // @[Modules.scala 53:83:@55272.4]
  assign _T_100851 = $signed(buffer_0_490) + $signed(buffer_3_491); // @[Modules.scala 53:83:@55274.4]
  assign _T_100852 = _T_100851[10:0]; // @[Modules.scala 53:83:@55275.4]
  assign buffer_14_637 = $signed(_T_100852); // @[Modules.scala 53:83:@55276.4]
  assign _T_100854 = $signed(buffer_4_492) + $signed(buffer_0_493); // @[Modules.scala 53:83:@55278.4]
  assign _T_100855 = _T_100854[10:0]; // @[Modules.scala 53:83:@55279.4]
  assign buffer_14_638 = $signed(_T_100855); // @[Modules.scala 53:83:@55280.4]
  assign _T_100857 = $signed(buffer_13_494) + $signed(buffer_3_495); // @[Modules.scala 53:83:@55282.4]
  assign _T_100858 = _T_100857[10:0]; // @[Modules.scala 53:83:@55283.4]
  assign buffer_14_639 = $signed(_T_100858); // @[Modules.scala 53:83:@55284.4]
  assign _T_100860 = $signed(buffer_14_496) + $signed(buffer_13_497); // @[Modules.scala 53:83:@55286.4]
  assign _T_100861 = _T_100860[10:0]; // @[Modules.scala 53:83:@55287.4]
  assign buffer_14_640 = $signed(_T_100861); // @[Modules.scala 53:83:@55288.4]
  assign _T_100863 = $signed(buffer_3_498) + $signed(buffer_14_499); // @[Modules.scala 53:83:@55290.4]
  assign _T_100864 = _T_100863[10:0]; // @[Modules.scala 53:83:@55291.4]
  assign buffer_14_641 = $signed(_T_100864); // @[Modules.scala 53:83:@55292.4]
  assign _T_100866 = $signed(buffer_14_500) + $signed(buffer_14_501); // @[Modules.scala 53:83:@55294.4]
  assign _T_100867 = _T_100866[10:0]; // @[Modules.scala 53:83:@55295.4]
  assign buffer_14_642 = $signed(_T_100867); // @[Modules.scala 53:83:@55296.4]
  assign _T_100869 = $signed(buffer_5_502) + $signed(buffer_8_503); // @[Modules.scala 53:83:@55298.4]
  assign _T_100870 = _T_100869[10:0]; // @[Modules.scala 53:83:@55299.4]
  assign buffer_14_643 = $signed(_T_100870); // @[Modules.scala 53:83:@55300.4]
  assign _T_100872 = $signed(buffer_1_504) + $signed(buffer_5_505); // @[Modules.scala 53:83:@55302.4]
  assign _T_100873 = _T_100872[10:0]; // @[Modules.scala 53:83:@55303.4]
  assign buffer_14_644 = $signed(_T_100873); // @[Modules.scala 53:83:@55304.4]
  assign _T_100878 = $signed(buffer_14_508) + $signed(buffer_14_509); // @[Modules.scala 53:83:@55310.4]
  assign _T_100879 = _T_100878[10:0]; // @[Modules.scala 53:83:@55311.4]
  assign buffer_14_646 = $signed(_T_100879); // @[Modules.scala 53:83:@55312.4]
  assign _T_100881 = $signed(buffer_14_510) + $signed(buffer_14_511); // @[Modules.scala 53:83:@55314.4]
  assign _T_100882 = _T_100881[10:0]; // @[Modules.scala 53:83:@55315.4]
  assign buffer_14_647 = $signed(_T_100882); // @[Modules.scala 53:83:@55316.4]
  assign _T_100887 = $signed(buffer_14_514) + $signed(buffer_10_515); // @[Modules.scala 53:83:@55322.4]
  assign _T_100888 = _T_100887[10:0]; // @[Modules.scala 53:83:@55323.4]
  assign buffer_14_649 = $signed(_T_100888); // @[Modules.scala 53:83:@55324.4]
  assign _T_100890 = $signed(buffer_14_516) + $signed(buffer_3_517); // @[Modules.scala 53:83:@55326.4]
  assign _T_100891 = _T_100890[10:0]; // @[Modules.scala 53:83:@55327.4]
  assign buffer_14_650 = $signed(_T_100891); // @[Modules.scala 53:83:@55328.4]
  assign _T_100893 = $signed(buffer_14_518) + $signed(buffer_3_519); // @[Modules.scala 53:83:@55330.4]
  assign _T_100894 = _T_100893[10:0]; // @[Modules.scala 53:83:@55331.4]
  assign buffer_14_651 = $signed(_T_100894); // @[Modules.scala 53:83:@55332.4]
  assign _T_100896 = $signed(buffer_10_520) + $signed(buffer_14_521); // @[Modules.scala 53:83:@55334.4]
  assign _T_100897 = _T_100896[10:0]; // @[Modules.scala 53:83:@55335.4]
  assign buffer_14_652 = $signed(_T_100897); // @[Modules.scala 53:83:@55336.4]
  assign _T_100899 = $signed(buffer_7_522) + $signed(buffer_4_523); // @[Modules.scala 53:83:@55338.4]
  assign _T_100900 = _T_100899[10:0]; // @[Modules.scala 53:83:@55339.4]
  assign buffer_14_653 = $signed(_T_100900); // @[Modules.scala 53:83:@55340.4]
  assign _T_100902 = $signed(buffer_13_524) + $signed(buffer_14_525); // @[Modules.scala 53:83:@55342.4]
  assign _T_100903 = _T_100902[10:0]; // @[Modules.scala 53:83:@55343.4]
  assign buffer_14_654 = $signed(_T_100903); // @[Modules.scala 53:83:@55344.4]
  assign _T_100905 = $signed(buffer_1_526) + $signed(buffer_14_527); // @[Modules.scala 53:83:@55346.4]
  assign _T_100906 = _T_100905[10:0]; // @[Modules.scala 53:83:@55347.4]
  assign buffer_14_655 = $signed(_T_100906); // @[Modules.scala 53:83:@55348.4]
  assign _T_100908 = $signed(buffer_0_528) + $signed(buffer_1_529); // @[Modules.scala 53:83:@55350.4]
  assign _T_100909 = _T_100908[10:0]; // @[Modules.scala 53:83:@55351.4]
  assign buffer_14_656 = $signed(_T_100909); // @[Modules.scala 53:83:@55352.4]
  assign _T_100914 = $signed(buffer_14_532) + $signed(buffer_3_533); // @[Modules.scala 53:83:@55358.4]
  assign _T_100915 = _T_100914[10:0]; // @[Modules.scala 53:83:@55359.4]
  assign buffer_14_658 = $signed(_T_100915); // @[Modules.scala 53:83:@55360.4]
  assign _T_100917 = $signed(buffer_14_534) + $signed(buffer_5_535); // @[Modules.scala 53:83:@55362.4]
  assign _T_100918 = _T_100917[10:0]; // @[Modules.scala 53:83:@55363.4]
  assign buffer_14_659 = $signed(_T_100918); // @[Modules.scala 53:83:@55364.4]
  assign _T_100920 = $signed(buffer_14_536) + $signed(buffer_4_537); // @[Modules.scala 53:83:@55366.4]
  assign _T_100921 = _T_100920[10:0]; // @[Modules.scala 53:83:@55367.4]
  assign buffer_14_660 = $signed(_T_100921); // @[Modules.scala 53:83:@55368.4]
  assign _T_100923 = $signed(buffer_13_538) + $signed(buffer_14_539); // @[Modules.scala 53:83:@55370.4]
  assign _T_100924 = _T_100923[10:0]; // @[Modules.scala 53:83:@55371.4]
  assign buffer_14_661 = $signed(_T_100924); // @[Modules.scala 53:83:@55372.4]
  assign _T_100926 = $signed(buffer_3_540) + $signed(buffer_5_541); // @[Modules.scala 53:83:@55374.4]
  assign _T_100927 = _T_100926[10:0]; // @[Modules.scala 53:83:@55375.4]
  assign buffer_14_662 = $signed(_T_100927); // @[Modules.scala 53:83:@55376.4]
  assign _T_100929 = $signed(buffer_5_542) + $signed(buffer_14_543); // @[Modules.scala 53:83:@55378.4]
  assign _T_100930 = _T_100929[10:0]; // @[Modules.scala 53:83:@55379.4]
  assign buffer_14_663 = $signed(_T_100930); // @[Modules.scala 53:83:@55380.4]
  assign _T_100935 = $signed(buffer_14_546) + $signed(buffer_14_547); // @[Modules.scala 53:83:@55386.4]
  assign _T_100936 = _T_100935[10:0]; // @[Modules.scala 53:83:@55387.4]
  assign buffer_14_665 = $signed(_T_100936); // @[Modules.scala 53:83:@55388.4]
  assign _T_100944 = $signed(buffer_14_552) + $signed(buffer_1_553); // @[Modules.scala 53:83:@55398.4]
  assign _T_100945 = _T_100944[10:0]; // @[Modules.scala 53:83:@55399.4]
  assign buffer_14_668 = $signed(_T_100945); // @[Modules.scala 53:83:@55400.4]
  assign _T_100947 = $signed(buffer_4_554) + $signed(buffer_14_555); // @[Modules.scala 53:83:@55402.4]
  assign _T_100948 = _T_100947[10:0]; // @[Modules.scala 53:83:@55403.4]
  assign buffer_14_669 = $signed(_T_100948); // @[Modules.scala 53:83:@55404.4]
  assign _T_100956 = $signed(buffer_1_560) + $signed(buffer_8_561); // @[Modules.scala 53:83:@55414.4]
  assign _T_100957 = _T_100956[10:0]; // @[Modules.scala 53:83:@55415.4]
  assign buffer_14_672 = $signed(_T_100957); // @[Modules.scala 53:83:@55416.4]
  assign _T_100959 = $signed(buffer_5_562) + $signed(buffer_4_563); // @[Modules.scala 53:83:@55418.4]
  assign _T_100960 = _T_100959[10:0]; // @[Modules.scala 53:83:@55419.4]
  assign buffer_14_673 = $signed(_T_100960); // @[Modules.scala 53:83:@55420.4]
  assign _T_100965 = $signed(buffer_14_566) + $signed(buffer_2_567); // @[Modules.scala 53:83:@55426.4]
  assign _T_100966 = _T_100965[10:0]; // @[Modules.scala 53:83:@55427.4]
  assign buffer_14_675 = $signed(_T_100966); // @[Modules.scala 53:83:@55428.4]
  assign _T_100968 = $signed(buffer_14_568) + $signed(buffer_14_569); // @[Modules.scala 53:83:@55430.4]
  assign _T_100969 = _T_100968[10:0]; // @[Modules.scala 53:83:@55431.4]
  assign buffer_14_676 = $signed(_T_100969); // @[Modules.scala 53:83:@55432.4]
  assign _T_100971 = $signed(buffer_14_570) + $signed(buffer_0_571); // @[Modules.scala 53:83:@55434.4]
  assign _T_100972 = _T_100971[10:0]; // @[Modules.scala 53:83:@55435.4]
  assign buffer_14_677 = $signed(_T_100972); // @[Modules.scala 53:83:@55436.4]
  assign _T_100974 = $signed(buffer_0_572) + $signed(buffer_14_573); // @[Modules.scala 53:83:@55438.4]
  assign _T_100975 = _T_100974[10:0]; // @[Modules.scala 53:83:@55439.4]
  assign buffer_14_678 = $signed(_T_100975); // @[Modules.scala 53:83:@55440.4]
  assign _T_100977 = $signed(buffer_14_574) + $signed(buffer_14_575); // @[Modules.scala 53:83:@55442.4]
  assign _T_100978 = _T_100977[10:0]; // @[Modules.scala 53:83:@55443.4]
  assign buffer_14_679 = $signed(_T_100978); // @[Modules.scala 53:83:@55444.4]
  assign _T_100980 = $signed(buffer_14_576) + $signed(buffer_14_577); // @[Modules.scala 53:83:@55446.4]
  assign _T_100981 = _T_100980[10:0]; // @[Modules.scala 53:83:@55447.4]
  assign buffer_14_680 = $signed(_T_100981); // @[Modules.scala 53:83:@55448.4]
  assign _T_100983 = $signed(buffer_3_578) + $signed(buffer_9_579); // @[Modules.scala 53:83:@55450.4]
  assign _T_100984 = _T_100983[10:0]; // @[Modules.scala 53:83:@55451.4]
  assign buffer_14_681 = $signed(_T_100984); // @[Modules.scala 53:83:@55452.4]
  assign _T_100986 = $signed(buffer_12_580) + $signed(buffer_10_581); // @[Modules.scala 53:83:@55454.4]
  assign _T_100987 = _T_100986[10:0]; // @[Modules.scala 53:83:@55455.4]
  assign buffer_14_682 = $signed(_T_100987); // @[Modules.scala 53:83:@55456.4]
  assign _T_100989 = $signed(buffer_1_582) + $signed(buffer_5_583); // @[Modules.scala 53:83:@55458.4]
  assign _T_100990 = _T_100989[10:0]; // @[Modules.scala 53:83:@55459.4]
  assign buffer_14_683 = $signed(_T_100990); // @[Modules.scala 53:83:@55460.4]
  assign _T_100995 = $signed(buffer_1_586) + $signed(buffer_14_587); // @[Modules.scala 53:83:@55466.4]
  assign _T_100996 = _T_100995[10:0]; // @[Modules.scala 53:83:@55467.4]
  assign buffer_14_685 = $signed(_T_100996); // @[Modules.scala 53:83:@55468.4]
  assign _T_100998 = $signed(buffer_14_588) + $signed(buffer_14_589); // @[Modules.scala 56:109:@55470.4]
  assign _T_100999 = _T_100998[10:0]; // @[Modules.scala 56:109:@55471.4]
  assign buffer_14_686 = $signed(_T_100999); // @[Modules.scala 56:109:@55472.4]
  assign _T_101001 = $signed(buffer_14_590) + $signed(buffer_14_591); // @[Modules.scala 56:109:@55474.4]
  assign _T_101002 = _T_101001[10:0]; // @[Modules.scala 56:109:@55475.4]
  assign buffer_14_687 = $signed(_T_101002); // @[Modules.scala 56:109:@55476.4]
  assign _T_101004 = $signed(buffer_14_592) + $signed(buffer_14_593); // @[Modules.scala 56:109:@55478.4]
  assign _T_101005 = _T_101004[10:0]; // @[Modules.scala 56:109:@55479.4]
  assign buffer_14_688 = $signed(_T_101005); // @[Modules.scala 56:109:@55480.4]
  assign _T_101007 = $signed(buffer_14_594) + $signed(buffer_14_595); // @[Modules.scala 56:109:@55482.4]
  assign _T_101008 = _T_101007[10:0]; // @[Modules.scala 56:109:@55483.4]
  assign buffer_14_689 = $signed(_T_101008); // @[Modules.scala 56:109:@55484.4]
  assign _T_101013 = $signed(buffer_14_598) + $signed(buffer_14_599); // @[Modules.scala 56:109:@55490.4]
  assign _T_101014 = _T_101013[10:0]; // @[Modules.scala 56:109:@55491.4]
  assign buffer_14_691 = $signed(_T_101014); // @[Modules.scala 56:109:@55492.4]
  assign _T_101016 = $signed(buffer_14_600) + $signed(buffer_14_601); // @[Modules.scala 56:109:@55494.4]
  assign _T_101017 = _T_101016[10:0]; // @[Modules.scala 56:109:@55495.4]
  assign buffer_14_692 = $signed(_T_101017); // @[Modules.scala 56:109:@55496.4]
  assign _T_101019 = $signed(buffer_14_602) + $signed(buffer_14_603); // @[Modules.scala 56:109:@55498.4]
  assign _T_101020 = _T_101019[10:0]; // @[Modules.scala 56:109:@55499.4]
  assign buffer_14_693 = $signed(_T_101020); // @[Modules.scala 56:109:@55500.4]
  assign _T_101022 = $signed(buffer_14_604) + $signed(buffer_14_605); // @[Modules.scala 56:109:@55502.4]
  assign _T_101023 = _T_101022[10:0]; // @[Modules.scala 56:109:@55503.4]
  assign buffer_14_694 = $signed(_T_101023); // @[Modules.scala 56:109:@55504.4]
  assign _T_101025 = $signed(buffer_14_606) + $signed(buffer_4_607); // @[Modules.scala 56:109:@55506.4]
  assign _T_101026 = _T_101025[10:0]; // @[Modules.scala 56:109:@55507.4]
  assign buffer_14_695 = $signed(_T_101026); // @[Modules.scala 56:109:@55508.4]
  assign _T_101028 = $signed(buffer_14_608) + $signed(buffer_14_609); // @[Modules.scala 56:109:@55510.4]
  assign _T_101029 = _T_101028[10:0]; // @[Modules.scala 56:109:@55511.4]
  assign buffer_14_696 = $signed(_T_101029); // @[Modules.scala 56:109:@55512.4]
  assign _T_101031 = $signed(buffer_14_610) + $signed(buffer_14_611); // @[Modules.scala 56:109:@55514.4]
  assign _T_101032 = _T_101031[10:0]; // @[Modules.scala 56:109:@55515.4]
  assign buffer_14_697 = $signed(_T_101032); // @[Modules.scala 56:109:@55516.4]
  assign _T_101034 = $signed(buffer_4_612) + $signed(buffer_14_613); // @[Modules.scala 56:109:@55518.4]
  assign _T_101035 = _T_101034[10:0]; // @[Modules.scala 56:109:@55519.4]
  assign buffer_14_698 = $signed(_T_101035); // @[Modules.scala 56:109:@55520.4]
  assign _T_101037 = $signed(buffer_14_614) + $signed(buffer_14_615); // @[Modules.scala 56:109:@55522.4]
  assign _T_101038 = _T_101037[10:0]; // @[Modules.scala 56:109:@55523.4]
  assign buffer_14_699 = $signed(_T_101038); // @[Modules.scala 56:109:@55524.4]
  assign _T_101040 = $signed(buffer_11_616) + $signed(buffer_14_617); // @[Modules.scala 56:109:@55526.4]
  assign _T_101041 = _T_101040[10:0]; // @[Modules.scala 56:109:@55527.4]
  assign buffer_14_700 = $signed(_T_101041); // @[Modules.scala 56:109:@55528.4]
  assign _T_101043 = $signed(buffer_14_618) + $signed(buffer_2_619); // @[Modules.scala 56:109:@55530.4]
  assign _T_101044 = _T_101043[10:0]; // @[Modules.scala 56:109:@55531.4]
  assign buffer_14_701 = $signed(_T_101044); // @[Modules.scala 56:109:@55532.4]
  assign _T_101046 = $signed(buffer_0_620) + $signed(buffer_14_621); // @[Modules.scala 56:109:@55534.4]
  assign _T_101047 = _T_101046[10:0]; // @[Modules.scala 56:109:@55535.4]
  assign buffer_14_702 = $signed(_T_101047); // @[Modules.scala 56:109:@55536.4]
  assign _T_101049 = $signed(buffer_14_622) + $signed(buffer_0_623); // @[Modules.scala 56:109:@55538.4]
  assign _T_101050 = _T_101049[10:0]; // @[Modules.scala 56:109:@55539.4]
  assign buffer_14_703 = $signed(_T_101050); // @[Modules.scala 56:109:@55540.4]
  assign _T_101052 = $signed(buffer_14_624) + $signed(buffer_14_625); // @[Modules.scala 56:109:@55542.4]
  assign _T_101053 = _T_101052[10:0]; // @[Modules.scala 56:109:@55543.4]
  assign buffer_14_704 = $signed(_T_101053); // @[Modules.scala 56:109:@55544.4]
  assign _T_101055 = $signed(buffer_1_626) + $signed(buffer_2_627); // @[Modules.scala 56:109:@55546.4]
  assign _T_101056 = _T_101055[10:0]; // @[Modules.scala 56:109:@55547.4]
  assign buffer_14_705 = $signed(_T_101056); // @[Modules.scala 56:109:@55548.4]
  assign _T_101058 = $signed(buffer_14_628) + $signed(buffer_14_629); // @[Modules.scala 56:109:@55550.4]
  assign _T_101059 = _T_101058[10:0]; // @[Modules.scala 56:109:@55551.4]
  assign buffer_14_706 = $signed(_T_101059); // @[Modules.scala 56:109:@55552.4]
  assign _T_101061 = $signed(buffer_14_630) + $signed(buffer_14_631); // @[Modules.scala 56:109:@55554.4]
  assign _T_101062 = _T_101061[10:0]; // @[Modules.scala 56:109:@55555.4]
  assign buffer_14_707 = $signed(_T_101062); // @[Modules.scala 56:109:@55556.4]
  assign _T_101064 = $signed(buffer_13_632) + $signed(buffer_14_633); // @[Modules.scala 56:109:@55558.4]
  assign _T_101065 = _T_101064[10:0]; // @[Modules.scala 56:109:@55559.4]
  assign buffer_14_708 = $signed(_T_101065); // @[Modules.scala 56:109:@55560.4]
  assign _T_101067 = $signed(buffer_14_634) + $signed(buffer_14_635); // @[Modules.scala 56:109:@55562.4]
  assign _T_101068 = _T_101067[10:0]; // @[Modules.scala 56:109:@55563.4]
  assign buffer_14_709 = $signed(_T_101068); // @[Modules.scala 56:109:@55564.4]
  assign _T_101070 = $signed(buffer_14_636) + $signed(buffer_14_637); // @[Modules.scala 56:109:@55566.4]
  assign _T_101071 = _T_101070[10:0]; // @[Modules.scala 56:109:@55567.4]
  assign buffer_14_710 = $signed(_T_101071); // @[Modules.scala 56:109:@55568.4]
  assign _T_101073 = $signed(buffer_14_638) + $signed(buffer_14_639); // @[Modules.scala 56:109:@55570.4]
  assign _T_101074 = _T_101073[10:0]; // @[Modules.scala 56:109:@55571.4]
  assign buffer_14_711 = $signed(_T_101074); // @[Modules.scala 56:109:@55572.4]
  assign _T_101076 = $signed(buffer_14_640) + $signed(buffer_14_641); // @[Modules.scala 56:109:@55574.4]
  assign _T_101077 = _T_101076[10:0]; // @[Modules.scala 56:109:@55575.4]
  assign buffer_14_712 = $signed(_T_101077); // @[Modules.scala 56:109:@55576.4]
  assign _T_101079 = $signed(buffer_14_642) + $signed(buffer_14_643); // @[Modules.scala 56:109:@55578.4]
  assign _T_101080 = _T_101079[10:0]; // @[Modules.scala 56:109:@55579.4]
  assign buffer_14_713 = $signed(_T_101080); // @[Modules.scala 56:109:@55580.4]
  assign _T_101082 = $signed(buffer_14_644) + $signed(buffer_12_645); // @[Modules.scala 56:109:@55582.4]
  assign _T_101083 = _T_101082[10:0]; // @[Modules.scala 56:109:@55583.4]
  assign buffer_14_714 = $signed(_T_101083); // @[Modules.scala 56:109:@55584.4]
  assign _T_101085 = $signed(buffer_14_646) + $signed(buffer_14_647); // @[Modules.scala 56:109:@55586.4]
  assign _T_101086 = _T_101085[10:0]; // @[Modules.scala 56:109:@55587.4]
  assign buffer_14_715 = $signed(_T_101086); // @[Modules.scala 56:109:@55588.4]
  assign _T_101088 = $signed(buffer_8_648) + $signed(buffer_14_649); // @[Modules.scala 56:109:@55590.4]
  assign _T_101089 = _T_101088[10:0]; // @[Modules.scala 56:109:@55591.4]
  assign buffer_14_716 = $signed(_T_101089); // @[Modules.scala 56:109:@55592.4]
  assign _T_101091 = $signed(buffer_14_650) + $signed(buffer_14_651); // @[Modules.scala 56:109:@55594.4]
  assign _T_101092 = _T_101091[10:0]; // @[Modules.scala 56:109:@55595.4]
  assign buffer_14_717 = $signed(_T_101092); // @[Modules.scala 56:109:@55596.4]
  assign _T_101094 = $signed(buffer_14_652) + $signed(buffer_14_653); // @[Modules.scala 56:109:@55598.4]
  assign _T_101095 = _T_101094[10:0]; // @[Modules.scala 56:109:@55599.4]
  assign buffer_14_718 = $signed(_T_101095); // @[Modules.scala 56:109:@55600.4]
  assign _T_101097 = $signed(buffer_14_654) + $signed(buffer_14_655); // @[Modules.scala 56:109:@55602.4]
  assign _T_101098 = _T_101097[10:0]; // @[Modules.scala 56:109:@55603.4]
  assign buffer_14_719 = $signed(_T_101098); // @[Modules.scala 56:109:@55604.4]
  assign _T_101100 = $signed(buffer_14_656) + $signed(buffer_3_657); // @[Modules.scala 56:109:@55606.4]
  assign _T_101101 = _T_101100[10:0]; // @[Modules.scala 56:109:@55607.4]
  assign buffer_14_720 = $signed(_T_101101); // @[Modules.scala 56:109:@55608.4]
  assign _T_101103 = $signed(buffer_14_658) + $signed(buffer_14_659); // @[Modules.scala 56:109:@55610.4]
  assign _T_101104 = _T_101103[10:0]; // @[Modules.scala 56:109:@55611.4]
  assign buffer_14_721 = $signed(_T_101104); // @[Modules.scala 56:109:@55612.4]
  assign _T_101106 = $signed(buffer_14_660) + $signed(buffer_14_661); // @[Modules.scala 56:109:@55614.4]
  assign _T_101107 = _T_101106[10:0]; // @[Modules.scala 56:109:@55615.4]
  assign buffer_14_722 = $signed(_T_101107); // @[Modules.scala 56:109:@55616.4]
  assign _T_101109 = $signed(buffer_14_662) + $signed(buffer_14_663); // @[Modules.scala 56:109:@55618.4]
  assign _T_101110 = _T_101109[10:0]; // @[Modules.scala 56:109:@55619.4]
  assign buffer_14_723 = $signed(_T_101110); // @[Modules.scala 56:109:@55620.4]
  assign _T_101112 = $signed(buffer_12_664) + $signed(buffer_14_665); // @[Modules.scala 56:109:@55622.4]
  assign _T_101113 = _T_101112[10:0]; // @[Modules.scala 56:109:@55623.4]
  assign buffer_14_724 = $signed(_T_101113); // @[Modules.scala 56:109:@55624.4]
  assign _T_101115 = $signed(buffer_1_666) + $signed(buffer_4_667); // @[Modules.scala 56:109:@55626.4]
  assign _T_101116 = _T_101115[10:0]; // @[Modules.scala 56:109:@55627.4]
  assign buffer_14_725 = $signed(_T_101116); // @[Modules.scala 56:109:@55628.4]
  assign _T_101118 = $signed(buffer_14_668) + $signed(buffer_14_669); // @[Modules.scala 56:109:@55630.4]
  assign _T_101119 = _T_101118[10:0]; // @[Modules.scala 56:109:@55631.4]
  assign buffer_14_726 = $signed(_T_101119); // @[Modules.scala 56:109:@55632.4]
  assign _T_101121 = $signed(buffer_11_670) + $signed(buffer_0_671); // @[Modules.scala 56:109:@55634.4]
  assign _T_101122 = _T_101121[10:0]; // @[Modules.scala 56:109:@55635.4]
  assign buffer_14_727 = $signed(_T_101122); // @[Modules.scala 56:109:@55636.4]
  assign _T_101124 = $signed(buffer_14_672) + $signed(buffer_14_673); // @[Modules.scala 56:109:@55638.4]
  assign _T_101125 = _T_101124[10:0]; // @[Modules.scala 56:109:@55639.4]
  assign buffer_14_728 = $signed(_T_101125); // @[Modules.scala 56:109:@55640.4]
  assign _T_101127 = $signed(buffer_0_674) + $signed(buffer_14_675); // @[Modules.scala 56:109:@55642.4]
  assign _T_101128 = _T_101127[10:0]; // @[Modules.scala 56:109:@55643.4]
  assign buffer_14_729 = $signed(_T_101128); // @[Modules.scala 56:109:@55644.4]
  assign _T_101130 = $signed(buffer_14_676) + $signed(buffer_14_677); // @[Modules.scala 56:109:@55646.4]
  assign _T_101131 = _T_101130[10:0]; // @[Modules.scala 56:109:@55647.4]
  assign buffer_14_730 = $signed(_T_101131); // @[Modules.scala 56:109:@55648.4]
  assign _T_101133 = $signed(buffer_14_678) + $signed(buffer_14_679); // @[Modules.scala 56:109:@55650.4]
  assign _T_101134 = _T_101133[10:0]; // @[Modules.scala 56:109:@55651.4]
  assign buffer_14_731 = $signed(_T_101134); // @[Modules.scala 56:109:@55652.4]
  assign _T_101136 = $signed(buffer_14_680) + $signed(buffer_14_681); // @[Modules.scala 56:109:@55654.4]
  assign _T_101137 = _T_101136[10:0]; // @[Modules.scala 56:109:@55655.4]
  assign buffer_14_732 = $signed(_T_101137); // @[Modules.scala 56:109:@55656.4]
  assign _T_101139 = $signed(buffer_14_682) + $signed(buffer_14_683); // @[Modules.scala 56:109:@55658.4]
  assign _T_101140 = _T_101139[10:0]; // @[Modules.scala 56:109:@55659.4]
  assign buffer_14_733 = $signed(_T_101140); // @[Modules.scala 56:109:@55660.4]
  assign _T_101142 = $signed(buffer_1_684) + $signed(buffer_14_685); // @[Modules.scala 56:109:@55662.4]
  assign _T_101143 = _T_101142[10:0]; // @[Modules.scala 56:109:@55663.4]
  assign buffer_14_734 = $signed(_T_101143); // @[Modules.scala 56:109:@55664.4]
  assign _T_101145 = $signed(buffer_14_686) + $signed(buffer_14_687); // @[Modules.scala 63:156:@55667.4]
  assign _T_101146 = _T_101145[10:0]; // @[Modules.scala 63:156:@55668.4]
  assign buffer_14_736 = $signed(_T_101146); // @[Modules.scala 63:156:@55669.4]
  assign _T_101148 = $signed(buffer_14_736) + $signed(buffer_14_688); // @[Modules.scala 63:156:@55671.4]
  assign _T_101149 = _T_101148[10:0]; // @[Modules.scala 63:156:@55672.4]
  assign buffer_14_737 = $signed(_T_101149); // @[Modules.scala 63:156:@55673.4]
  assign _T_101151 = $signed(buffer_14_737) + $signed(buffer_14_689); // @[Modules.scala 63:156:@55675.4]
  assign _T_101152 = _T_101151[10:0]; // @[Modules.scala 63:156:@55676.4]
  assign buffer_14_738 = $signed(_T_101152); // @[Modules.scala 63:156:@55677.4]
  assign _T_101154 = $signed(buffer_14_738) + $signed(buffer_3_690); // @[Modules.scala 63:156:@55679.4]
  assign _T_101155 = _T_101154[10:0]; // @[Modules.scala 63:156:@55680.4]
  assign buffer_14_739 = $signed(_T_101155); // @[Modules.scala 63:156:@55681.4]
  assign _T_101157 = $signed(buffer_14_739) + $signed(buffer_14_691); // @[Modules.scala 63:156:@55683.4]
  assign _T_101158 = _T_101157[10:0]; // @[Modules.scala 63:156:@55684.4]
  assign buffer_14_740 = $signed(_T_101158); // @[Modules.scala 63:156:@55685.4]
  assign _T_101160 = $signed(buffer_14_740) + $signed(buffer_14_692); // @[Modules.scala 63:156:@55687.4]
  assign _T_101161 = _T_101160[10:0]; // @[Modules.scala 63:156:@55688.4]
  assign buffer_14_741 = $signed(_T_101161); // @[Modules.scala 63:156:@55689.4]
  assign _T_101163 = $signed(buffer_14_741) + $signed(buffer_14_693); // @[Modules.scala 63:156:@55691.4]
  assign _T_101164 = _T_101163[10:0]; // @[Modules.scala 63:156:@55692.4]
  assign buffer_14_742 = $signed(_T_101164); // @[Modules.scala 63:156:@55693.4]
  assign _T_101166 = $signed(buffer_14_742) + $signed(buffer_14_694); // @[Modules.scala 63:156:@55695.4]
  assign _T_101167 = _T_101166[10:0]; // @[Modules.scala 63:156:@55696.4]
  assign buffer_14_743 = $signed(_T_101167); // @[Modules.scala 63:156:@55697.4]
  assign _T_101169 = $signed(buffer_14_743) + $signed(buffer_14_695); // @[Modules.scala 63:156:@55699.4]
  assign _T_101170 = _T_101169[10:0]; // @[Modules.scala 63:156:@55700.4]
  assign buffer_14_744 = $signed(_T_101170); // @[Modules.scala 63:156:@55701.4]
  assign _T_101172 = $signed(buffer_14_744) + $signed(buffer_14_696); // @[Modules.scala 63:156:@55703.4]
  assign _T_101173 = _T_101172[10:0]; // @[Modules.scala 63:156:@55704.4]
  assign buffer_14_745 = $signed(_T_101173); // @[Modules.scala 63:156:@55705.4]
  assign _T_101175 = $signed(buffer_14_745) + $signed(buffer_14_697); // @[Modules.scala 63:156:@55707.4]
  assign _T_101176 = _T_101175[10:0]; // @[Modules.scala 63:156:@55708.4]
  assign buffer_14_746 = $signed(_T_101176); // @[Modules.scala 63:156:@55709.4]
  assign _T_101178 = $signed(buffer_14_746) + $signed(buffer_14_698); // @[Modules.scala 63:156:@55711.4]
  assign _T_101179 = _T_101178[10:0]; // @[Modules.scala 63:156:@55712.4]
  assign buffer_14_747 = $signed(_T_101179); // @[Modules.scala 63:156:@55713.4]
  assign _T_101181 = $signed(buffer_14_747) + $signed(buffer_14_699); // @[Modules.scala 63:156:@55715.4]
  assign _T_101182 = _T_101181[10:0]; // @[Modules.scala 63:156:@55716.4]
  assign buffer_14_748 = $signed(_T_101182); // @[Modules.scala 63:156:@55717.4]
  assign _T_101184 = $signed(buffer_14_748) + $signed(buffer_14_700); // @[Modules.scala 63:156:@55719.4]
  assign _T_101185 = _T_101184[10:0]; // @[Modules.scala 63:156:@55720.4]
  assign buffer_14_749 = $signed(_T_101185); // @[Modules.scala 63:156:@55721.4]
  assign _T_101187 = $signed(buffer_14_749) + $signed(buffer_14_701); // @[Modules.scala 63:156:@55723.4]
  assign _T_101188 = _T_101187[10:0]; // @[Modules.scala 63:156:@55724.4]
  assign buffer_14_750 = $signed(_T_101188); // @[Modules.scala 63:156:@55725.4]
  assign _T_101190 = $signed(buffer_14_750) + $signed(buffer_14_702); // @[Modules.scala 63:156:@55727.4]
  assign _T_101191 = _T_101190[10:0]; // @[Modules.scala 63:156:@55728.4]
  assign buffer_14_751 = $signed(_T_101191); // @[Modules.scala 63:156:@55729.4]
  assign _T_101193 = $signed(buffer_14_751) + $signed(buffer_14_703); // @[Modules.scala 63:156:@55731.4]
  assign _T_101194 = _T_101193[10:0]; // @[Modules.scala 63:156:@55732.4]
  assign buffer_14_752 = $signed(_T_101194); // @[Modules.scala 63:156:@55733.4]
  assign _T_101196 = $signed(buffer_14_752) + $signed(buffer_14_704); // @[Modules.scala 63:156:@55735.4]
  assign _T_101197 = _T_101196[10:0]; // @[Modules.scala 63:156:@55736.4]
  assign buffer_14_753 = $signed(_T_101197); // @[Modules.scala 63:156:@55737.4]
  assign _T_101199 = $signed(buffer_14_753) + $signed(buffer_14_705); // @[Modules.scala 63:156:@55739.4]
  assign _T_101200 = _T_101199[10:0]; // @[Modules.scala 63:156:@55740.4]
  assign buffer_14_754 = $signed(_T_101200); // @[Modules.scala 63:156:@55741.4]
  assign _T_101202 = $signed(buffer_14_754) + $signed(buffer_14_706); // @[Modules.scala 63:156:@55743.4]
  assign _T_101203 = _T_101202[10:0]; // @[Modules.scala 63:156:@55744.4]
  assign buffer_14_755 = $signed(_T_101203); // @[Modules.scala 63:156:@55745.4]
  assign _T_101205 = $signed(buffer_14_755) + $signed(buffer_14_707); // @[Modules.scala 63:156:@55747.4]
  assign _T_101206 = _T_101205[10:0]; // @[Modules.scala 63:156:@55748.4]
  assign buffer_14_756 = $signed(_T_101206); // @[Modules.scala 63:156:@55749.4]
  assign _T_101208 = $signed(buffer_14_756) + $signed(buffer_14_708); // @[Modules.scala 63:156:@55751.4]
  assign _T_101209 = _T_101208[10:0]; // @[Modules.scala 63:156:@55752.4]
  assign buffer_14_757 = $signed(_T_101209); // @[Modules.scala 63:156:@55753.4]
  assign _T_101211 = $signed(buffer_14_757) + $signed(buffer_14_709); // @[Modules.scala 63:156:@55755.4]
  assign _T_101212 = _T_101211[10:0]; // @[Modules.scala 63:156:@55756.4]
  assign buffer_14_758 = $signed(_T_101212); // @[Modules.scala 63:156:@55757.4]
  assign _T_101214 = $signed(buffer_14_758) + $signed(buffer_14_710); // @[Modules.scala 63:156:@55759.4]
  assign _T_101215 = _T_101214[10:0]; // @[Modules.scala 63:156:@55760.4]
  assign buffer_14_759 = $signed(_T_101215); // @[Modules.scala 63:156:@55761.4]
  assign _T_101217 = $signed(buffer_14_759) + $signed(buffer_14_711); // @[Modules.scala 63:156:@55763.4]
  assign _T_101218 = _T_101217[10:0]; // @[Modules.scala 63:156:@55764.4]
  assign buffer_14_760 = $signed(_T_101218); // @[Modules.scala 63:156:@55765.4]
  assign _T_101220 = $signed(buffer_14_760) + $signed(buffer_14_712); // @[Modules.scala 63:156:@55767.4]
  assign _T_101221 = _T_101220[10:0]; // @[Modules.scala 63:156:@55768.4]
  assign buffer_14_761 = $signed(_T_101221); // @[Modules.scala 63:156:@55769.4]
  assign _T_101223 = $signed(buffer_14_761) + $signed(buffer_14_713); // @[Modules.scala 63:156:@55771.4]
  assign _T_101224 = _T_101223[10:0]; // @[Modules.scala 63:156:@55772.4]
  assign buffer_14_762 = $signed(_T_101224); // @[Modules.scala 63:156:@55773.4]
  assign _T_101226 = $signed(buffer_14_762) + $signed(buffer_14_714); // @[Modules.scala 63:156:@55775.4]
  assign _T_101227 = _T_101226[10:0]; // @[Modules.scala 63:156:@55776.4]
  assign buffer_14_763 = $signed(_T_101227); // @[Modules.scala 63:156:@55777.4]
  assign _T_101229 = $signed(buffer_14_763) + $signed(buffer_14_715); // @[Modules.scala 63:156:@55779.4]
  assign _T_101230 = _T_101229[10:0]; // @[Modules.scala 63:156:@55780.4]
  assign buffer_14_764 = $signed(_T_101230); // @[Modules.scala 63:156:@55781.4]
  assign _T_101232 = $signed(buffer_14_764) + $signed(buffer_14_716); // @[Modules.scala 63:156:@55783.4]
  assign _T_101233 = _T_101232[10:0]; // @[Modules.scala 63:156:@55784.4]
  assign buffer_14_765 = $signed(_T_101233); // @[Modules.scala 63:156:@55785.4]
  assign _T_101235 = $signed(buffer_14_765) + $signed(buffer_14_717); // @[Modules.scala 63:156:@55787.4]
  assign _T_101236 = _T_101235[10:0]; // @[Modules.scala 63:156:@55788.4]
  assign buffer_14_766 = $signed(_T_101236); // @[Modules.scala 63:156:@55789.4]
  assign _T_101238 = $signed(buffer_14_766) + $signed(buffer_14_718); // @[Modules.scala 63:156:@55791.4]
  assign _T_101239 = _T_101238[10:0]; // @[Modules.scala 63:156:@55792.4]
  assign buffer_14_767 = $signed(_T_101239); // @[Modules.scala 63:156:@55793.4]
  assign _T_101241 = $signed(buffer_14_767) + $signed(buffer_14_719); // @[Modules.scala 63:156:@55795.4]
  assign _T_101242 = _T_101241[10:0]; // @[Modules.scala 63:156:@55796.4]
  assign buffer_14_768 = $signed(_T_101242); // @[Modules.scala 63:156:@55797.4]
  assign _T_101244 = $signed(buffer_14_768) + $signed(buffer_14_720); // @[Modules.scala 63:156:@55799.4]
  assign _T_101245 = _T_101244[10:0]; // @[Modules.scala 63:156:@55800.4]
  assign buffer_14_769 = $signed(_T_101245); // @[Modules.scala 63:156:@55801.4]
  assign _T_101247 = $signed(buffer_14_769) + $signed(buffer_14_721); // @[Modules.scala 63:156:@55803.4]
  assign _T_101248 = _T_101247[10:0]; // @[Modules.scala 63:156:@55804.4]
  assign buffer_14_770 = $signed(_T_101248); // @[Modules.scala 63:156:@55805.4]
  assign _T_101250 = $signed(buffer_14_770) + $signed(buffer_14_722); // @[Modules.scala 63:156:@55807.4]
  assign _T_101251 = _T_101250[10:0]; // @[Modules.scala 63:156:@55808.4]
  assign buffer_14_771 = $signed(_T_101251); // @[Modules.scala 63:156:@55809.4]
  assign _T_101253 = $signed(buffer_14_771) + $signed(buffer_14_723); // @[Modules.scala 63:156:@55811.4]
  assign _T_101254 = _T_101253[10:0]; // @[Modules.scala 63:156:@55812.4]
  assign buffer_14_772 = $signed(_T_101254); // @[Modules.scala 63:156:@55813.4]
  assign _T_101256 = $signed(buffer_14_772) + $signed(buffer_14_724); // @[Modules.scala 63:156:@55815.4]
  assign _T_101257 = _T_101256[10:0]; // @[Modules.scala 63:156:@55816.4]
  assign buffer_14_773 = $signed(_T_101257); // @[Modules.scala 63:156:@55817.4]
  assign _T_101259 = $signed(buffer_14_773) + $signed(buffer_14_725); // @[Modules.scala 63:156:@55819.4]
  assign _T_101260 = _T_101259[10:0]; // @[Modules.scala 63:156:@55820.4]
  assign buffer_14_774 = $signed(_T_101260); // @[Modules.scala 63:156:@55821.4]
  assign _T_101262 = $signed(buffer_14_774) + $signed(buffer_14_726); // @[Modules.scala 63:156:@55823.4]
  assign _T_101263 = _T_101262[10:0]; // @[Modules.scala 63:156:@55824.4]
  assign buffer_14_775 = $signed(_T_101263); // @[Modules.scala 63:156:@55825.4]
  assign _T_101265 = $signed(buffer_14_775) + $signed(buffer_14_727); // @[Modules.scala 63:156:@55827.4]
  assign _T_101266 = _T_101265[10:0]; // @[Modules.scala 63:156:@55828.4]
  assign buffer_14_776 = $signed(_T_101266); // @[Modules.scala 63:156:@55829.4]
  assign _T_101268 = $signed(buffer_14_776) + $signed(buffer_14_728); // @[Modules.scala 63:156:@55831.4]
  assign _T_101269 = _T_101268[10:0]; // @[Modules.scala 63:156:@55832.4]
  assign buffer_14_777 = $signed(_T_101269); // @[Modules.scala 63:156:@55833.4]
  assign _T_101271 = $signed(buffer_14_777) + $signed(buffer_14_729); // @[Modules.scala 63:156:@55835.4]
  assign _T_101272 = _T_101271[10:0]; // @[Modules.scala 63:156:@55836.4]
  assign buffer_14_778 = $signed(_T_101272); // @[Modules.scala 63:156:@55837.4]
  assign _T_101274 = $signed(buffer_14_778) + $signed(buffer_14_730); // @[Modules.scala 63:156:@55839.4]
  assign _T_101275 = _T_101274[10:0]; // @[Modules.scala 63:156:@55840.4]
  assign buffer_14_779 = $signed(_T_101275); // @[Modules.scala 63:156:@55841.4]
  assign _T_101277 = $signed(buffer_14_779) + $signed(buffer_14_731); // @[Modules.scala 63:156:@55843.4]
  assign _T_101278 = _T_101277[10:0]; // @[Modules.scala 63:156:@55844.4]
  assign buffer_14_780 = $signed(_T_101278); // @[Modules.scala 63:156:@55845.4]
  assign _T_101280 = $signed(buffer_14_780) + $signed(buffer_14_732); // @[Modules.scala 63:156:@55847.4]
  assign _T_101281 = _T_101280[10:0]; // @[Modules.scala 63:156:@55848.4]
  assign buffer_14_781 = $signed(_T_101281); // @[Modules.scala 63:156:@55849.4]
  assign _T_101283 = $signed(buffer_14_781) + $signed(buffer_14_733); // @[Modules.scala 63:156:@55851.4]
  assign _T_101284 = _T_101283[10:0]; // @[Modules.scala 63:156:@55852.4]
  assign buffer_14_782 = $signed(_T_101284); // @[Modules.scala 63:156:@55853.4]
  assign _T_101286 = $signed(buffer_14_782) + $signed(buffer_14_734); // @[Modules.scala 63:156:@55855.4]
  assign _T_101287 = _T_101286[10:0]; // @[Modules.scala 63:156:@55856.4]
  assign buffer_14_783 = $signed(_T_101287); // @[Modules.scala 63:156:@55857.4]
  assign _T_101401 = $signed(io_in_48) - $signed(io_in_49); // @[Modules.scala 40:46:@55986.4]
  assign _T_101402 = _T_101401[4:0]; // @[Modules.scala 40:46:@55987.4]
  assign _T_101403 = $signed(_T_101402); // @[Modules.scala 40:46:@55988.4]
  assign _T_101459 = $signed(_T_64110) + $signed(io_in_77); // @[Modules.scala 43:47:@56054.4]
  assign _T_101460 = _T_101459[4:0]; // @[Modules.scala 43:47:@56055.4]
  assign _T_101461 = $signed(_T_101460); // @[Modules.scala 43:47:@56056.4]
  assign _T_101932 = $signed(_T_55016) + $signed(io_in_259); // @[Modules.scala 43:47:@56568.4]
  assign _T_101933 = _T_101932[4:0]; // @[Modules.scala 43:47:@56569.4]
  assign _T_101934 = $signed(_T_101933); // @[Modules.scala 43:47:@56570.4]
  assign _T_102198 = $signed(io_in_366) + $signed(io_in_367); // @[Modules.scala 37:46:@56862.4]
  assign _T_102199 = _T_102198[4:0]; // @[Modules.scala 37:46:@56863.4]
  assign _T_102200 = $signed(_T_102199); // @[Modules.scala 37:46:@56864.4]
  assign _T_102496 = $signed(io_in_498) - $signed(io_in_499); // @[Modules.scala 40:46:@57201.4]
  assign _T_102497 = _T_102496[4:0]; // @[Modules.scala 40:46:@57202.4]
  assign _T_102498 = $signed(_T_102497); // @[Modules.scala 40:46:@57203.4]
  assign _T_102670 = $signed(io_in_574) - $signed(io_in_575); // @[Modules.scala 40:46:@57398.4]
  assign _T_102671 = _T_102670[4:0]; // @[Modules.scala 40:46:@57399.4]
  assign _T_102672 = $signed(_T_102671); // @[Modules.scala 40:46:@57400.4]
  assign _T_102769 = $signed(io_in_616) - $signed(io_in_617); // @[Modules.scala 40:46:@57509.4]
  assign _T_102770 = _T_102769[4:0]; // @[Modules.scala 40:46:@57510.4]
  assign _T_102771 = $signed(_T_102770); // @[Modules.scala 40:46:@57511.4]
  assign _T_102935 = $signed(_T_62429) + $signed(io_in_677); // @[Modules.scala 43:47:@57686.4]
  assign _T_102936 = _T_102935[4:0]; // @[Modules.scala 43:47:@57687.4]
  assign _T_102937 = $signed(_T_102936); // @[Modules.scala 43:47:@57688.4]
  assign _T_103033 = $signed(_T_59258) + $signed(io_in_713); // @[Modules.scala 43:47:@57791.4]
  assign _T_103034 = _T_103033[4:0]; // @[Modules.scala 43:47:@57792.4]
  assign _T_103035 = $signed(_T_103034); // @[Modules.scala 43:47:@57793.4]
  assign _T_103087 = $signed(_T_59312) + $signed(io_in_733); // @[Modules.scala 43:47:@57849.4]
  assign _T_103088 = _T_103087[4:0]; // @[Modules.scala 43:47:@57850.4]
  assign _T_103089 = $signed(_T_103088); // @[Modules.scala 43:47:@57851.4]
  assign _T_103176 = $signed(io_in_778) - $signed(io_in_779); // @[Modules.scala 40:46:@57956.4]
  assign _T_103177 = _T_103176[4:0]; // @[Modules.scala 40:46:@57957.4]
  assign _T_103178 = $signed(_T_103177); // @[Modules.scala 40:46:@57958.4]
  assign _T_103198 = $signed(buffer_1_6) + $signed(buffer_0_7); // @[Modules.scala 50:57:@57983.4]
  assign _T_103199 = _T_103198[10:0]; // @[Modules.scala 50:57:@57984.4]
  assign buffer_15_395 = $signed(_T_103199); // @[Modules.scala 50:57:@57985.4]
  assign _T_103201 = $signed(buffer_0_8) + $signed(buffer_9_9); // @[Modules.scala 50:57:@57987.4]
  assign _T_103202 = _T_103201[10:0]; // @[Modules.scala 50:57:@57988.4]
  assign buffer_15_396 = $signed(_T_103202); // @[Modules.scala 50:57:@57989.4]
  assign _T_103204 = $signed(buffer_5_10) + $signed(buffer_1_11); // @[Modules.scala 50:57:@57991.4]
  assign _T_103205 = _T_103204[10:0]; // @[Modules.scala 50:57:@57992.4]
  assign buffer_15_397 = $signed(_T_103205); // @[Modules.scala 50:57:@57993.4]
  assign _T_103207 = $signed(buffer_0_12) + $signed(buffer_4_13); // @[Modules.scala 50:57:@57995.4]
  assign _T_103208 = _T_103207[10:0]; // @[Modules.scala 50:57:@57996.4]
  assign buffer_15_398 = $signed(_T_103208); // @[Modules.scala 50:57:@57997.4]
  assign _T_103216 = $signed(buffer_0_18) + $signed(buffer_1_19); // @[Modules.scala 50:57:@58007.4]
  assign _T_103217 = _T_103216[10:0]; // @[Modules.scala 50:57:@58008.4]
  assign buffer_15_401 = $signed(_T_103217); // @[Modules.scala 50:57:@58009.4]
  assign _T_103222 = $signed(buffer_4_22) + $signed(buffer_11_23); // @[Modules.scala 50:57:@58015.4]
  assign _T_103223 = _T_103222[10:0]; // @[Modules.scala 50:57:@58016.4]
  assign buffer_15_403 = $signed(_T_103223); // @[Modules.scala 50:57:@58017.4]
  assign buffer_15_24 = {{6{_T_101403[4]}},_T_101403}; // @[Modules.scala 32:22:@8.4]
  assign _T_103225 = $signed(buffer_15_24) + $signed(buffer_1_25); // @[Modules.scala 50:57:@58019.4]
  assign _T_103226 = _T_103225[10:0]; // @[Modules.scala 50:57:@58020.4]
  assign buffer_15_404 = $signed(_T_103226); // @[Modules.scala 50:57:@58021.4]
  assign _T_103228 = $signed(buffer_2_26) + $signed(buffer_3_27); // @[Modules.scala 50:57:@58023.4]
  assign _T_103229 = _T_103228[10:0]; // @[Modules.scala 50:57:@58024.4]
  assign buffer_15_405 = $signed(_T_103229); // @[Modules.scala 50:57:@58025.4]
  assign buffer_15_38 = {{6{_T_101461[4]}},_T_101461}; // @[Modules.scala 32:22:@8.4]
  assign _T_103246 = $signed(buffer_15_38) + $signed(buffer_0_39); // @[Modules.scala 50:57:@58047.4]
  assign _T_103247 = _T_103246[10:0]; // @[Modules.scala 50:57:@58048.4]
  assign buffer_15_411 = $signed(_T_103247); // @[Modules.scala 50:57:@58049.4]
  assign _T_103252 = $signed(buffer_1_42) + $signed(buffer_11_43); // @[Modules.scala 50:57:@58055.4]
  assign _T_103253 = _T_103252[10:0]; // @[Modules.scala 50:57:@58056.4]
  assign buffer_15_413 = $signed(_T_103253); // @[Modules.scala 50:57:@58057.4]
  assign _T_103255 = $signed(buffer_3_44) + $signed(buffer_14_45); // @[Modules.scala 50:57:@58059.4]
  assign _T_103256 = _T_103255[10:0]; // @[Modules.scala 50:57:@58060.4]
  assign buffer_15_414 = $signed(_T_103256); // @[Modules.scala 50:57:@58061.4]
  assign _T_103279 = $signed(buffer_8_60) + $signed(buffer_0_61); // @[Modules.scala 50:57:@58091.4]
  assign _T_103280 = _T_103279[10:0]; // @[Modules.scala 50:57:@58092.4]
  assign buffer_15_422 = $signed(_T_103280); // @[Modules.scala 50:57:@58093.4]
  assign _T_103285 = $signed(buffer_1_64) + $signed(buffer_0_65); // @[Modules.scala 50:57:@58099.4]
  assign _T_103286 = _T_103285[10:0]; // @[Modules.scala 50:57:@58100.4]
  assign buffer_15_424 = $signed(_T_103286); // @[Modules.scala 50:57:@58101.4]
  assign _T_103294 = $signed(buffer_14_70) + $signed(buffer_1_71); // @[Modules.scala 50:57:@58111.4]
  assign _T_103295 = _T_103294[10:0]; // @[Modules.scala 50:57:@58112.4]
  assign buffer_15_427 = $signed(_T_103295); // @[Modules.scala 50:57:@58113.4]
  assign _T_103303 = $signed(buffer_3_76) + $signed(buffer_10_77); // @[Modules.scala 50:57:@58123.4]
  assign _T_103304 = _T_103303[10:0]; // @[Modules.scala 50:57:@58124.4]
  assign buffer_15_430 = $signed(_T_103304); // @[Modules.scala 50:57:@58125.4]
  assign _T_103306 = $signed(buffer_0_78) + $signed(buffer_3_79); // @[Modules.scala 50:57:@58127.4]
  assign _T_103307 = _T_103306[10:0]; // @[Modules.scala 50:57:@58128.4]
  assign buffer_15_431 = $signed(_T_103307); // @[Modules.scala 50:57:@58129.4]
  assign _T_103312 = $signed(buffer_1_82) + $signed(buffer_6_83); // @[Modules.scala 50:57:@58135.4]
  assign _T_103313 = _T_103312[10:0]; // @[Modules.scala 50:57:@58136.4]
  assign buffer_15_433 = $signed(_T_103313); // @[Modules.scala 50:57:@58137.4]
  assign _T_103315 = $signed(buffer_0_84) + $signed(buffer_9_85); // @[Modules.scala 50:57:@58139.4]
  assign _T_103316 = _T_103315[10:0]; // @[Modules.scala 50:57:@58140.4]
  assign buffer_15_434 = $signed(_T_103316); // @[Modules.scala 50:57:@58141.4]
  assign _T_103318 = $signed(buffer_2_86) + $signed(buffer_1_87); // @[Modules.scala 50:57:@58143.4]
  assign _T_103319 = _T_103318[10:0]; // @[Modules.scala 50:57:@58144.4]
  assign buffer_15_435 = $signed(_T_103319); // @[Modules.scala 50:57:@58145.4]
  assign _T_103321 = $signed(buffer_10_88) + $signed(buffer_1_89); // @[Modules.scala 50:57:@58147.4]
  assign _T_103322 = _T_103321[10:0]; // @[Modules.scala 50:57:@58148.4]
  assign buffer_15_436 = $signed(_T_103322); // @[Modules.scala 50:57:@58149.4]
  assign _T_103336 = $signed(buffer_0_98) + $signed(buffer_3_99); // @[Modules.scala 50:57:@58167.4]
  assign _T_103337 = _T_103336[10:0]; // @[Modules.scala 50:57:@58168.4]
  assign buffer_15_441 = $signed(_T_103337); // @[Modules.scala 50:57:@58169.4]
  assign _T_103339 = $signed(buffer_0_100) + $signed(buffer_1_101); // @[Modules.scala 50:57:@58171.4]
  assign _T_103340 = _T_103339[10:0]; // @[Modules.scala 50:57:@58172.4]
  assign buffer_15_442 = $signed(_T_103340); // @[Modules.scala 50:57:@58173.4]
  assign _T_103348 = $signed(buffer_4_106) + $signed(buffer_2_107); // @[Modules.scala 50:57:@58183.4]
  assign _T_103349 = _T_103348[10:0]; // @[Modules.scala 50:57:@58184.4]
  assign buffer_15_445 = $signed(_T_103349); // @[Modules.scala 50:57:@58185.4]
  assign _T_103363 = $signed(buffer_0_116) + $signed(buffer_3_117); // @[Modules.scala 50:57:@58203.4]
  assign _T_103364 = _T_103363[10:0]; // @[Modules.scala 50:57:@58204.4]
  assign buffer_15_450 = $signed(_T_103364); // @[Modules.scala 50:57:@58205.4]
  assign buffer_15_129 = {{6{_T_101934[4]}},_T_101934}; // @[Modules.scala 32:22:@8.4]
  assign _T_103381 = $signed(buffer_3_128) + $signed(buffer_15_129); // @[Modules.scala 50:57:@58227.4]
  assign _T_103382 = _T_103381[10:0]; // @[Modules.scala 50:57:@58228.4]
  assign buffer_15_456 = $signed(_T_103382); // @[Modules.scala 50:57:@58229.4]
  assign _T_103402 = $signed(buffer_7_142) + $signed(buffer_2_143); // @[Modules.scala 50:57:@58255.4]
  assign _T_103403 = _T_103402[10:0]; // @[Modules.scala 50:57:@58256.4]
  assign buffer_15_463 = $signed(_T_103403); // @[Modules.scala 50:57:@58257.4]
  assign _T_103414 = $signed(buffer_5_150) + $signed(buffer_0_151); // @[Modules.scala 50:57:@58271.4]
  assign _T_103415 = _T_103414[10:0]; // @[Modules.scala 50:57:@58272.4]
  assign buffer_15_467 = $signed(_T_103415); // @[Modules.scala 50:57:@58273.4]
  assign _T_103423 = $signed(buffer_9_156) + $signed(buffer_2_157); // @[Modules.scala 50:57:@58283.4]
  assign _T_103424 = _T_103423[10:0]; // @[Modules.scala 50:57:@58284.4]
  assign buffer_15_470 = $signed(_T_103424); // @[Modules.scala 50:57:@58285.4]
  assign _T_103426 = $signed(buffer_13_158) + $signed(buffer_3_159); // @[Modules.scala 50:57:@58287.4]
  assign _T_103427 = _T_103426[10:0]; // @[Modules.scala 50:57:@58288.4]
  assign buffer_15_471 = $signed(_T_103427); // @[Modules.scala 50:57:@58289.4]
  assign _T_103432 = $signed(buffer_0_162) + $signed(buffer_5_163); // @[Modules.scala 50:57:@58295.4]
  assign _T_103433 = _T_103432[10:0]; // @[Modules.scala 50:57:@58296.4]
  assign buffer_15_473 = $signed(_T_103433); // @[Modules.scala 50:57:@58297.4]
  assign _T_103441 = $signed(buffer_5_168) + $signed(buffer_6_169); // @[Modules.scala 50:57:@58307.4]
  assign _T_103442 = _T_103441[10:0]; // @[Modules.scala 50:57:@58308.4]
  assign buffer_15_476 = $signed(_T_103442); // @[Modules.scala 50:57:@58309.4]
  assign _T_103459 = $signed(buffer_14_180) + $signed(buffer_0_181); // @[Modules.scala 50:57:@58331.4]
  assign _T_103460 = _T_103459[10:0]; // @[Modules.scala 50:57:@58332.4]
  assign buffer_15_482 = $signed(_T_103460); // @[Modules.scala 50:57:@58333.4]
  assign buffer_15_183 = {{6{_T_102200[4]}},_T_102200}; // @[Modules.scala 32:22:@8.4]
  assign _T_103462 = $signed(buffer_3_182) + $signed(buffer_15_183); // @[Modules.scala 50:57:@58335.4]
  assign _T_103463 = _T_103462[10:0]; // @[Modules.scala 50:57:@58336.4]
  assign buffer_15_483 = $signed(_T_103463); // @[Modules.scala 50:57:@58337.4]
  assign _T_103465 = $signed(buffer_0_184) + $signed(buffer_3_185); // @[Modules.scala 50:57:@58339.4]
  assign _T_103466 = _T_103465[10:0]; // @[Modules.scala 50:57:@58340.4]
  assign buffer_15_484 = $signed(_T_103466); // @[Modules.scala 50:57:@58341.4]
  assign _T_103495 = $signed(buffer_3_204) + $signed(buffer_2_205); // @[Modules.scala 50:57:@58379.4]
  assign _T_103496 = _T_103495[10:0]; // @[Modules.scala 50:57:@58380.4]
  assign buffer_15_494 = $signed(_T_103496); // @[Modules.scala 50:57:@58381.4]
  assign _T_103516 = $signed(buffer_1_218) + $signed(buffer_6_219); // @[Modules.scala 50:57:@58407.4]
  assign _T_103517 = _T_103516[10:0]; // @[Modules.scala 50:57:@58408.4]
  assign buffer_15_501 = $signed(_T_103517); // @[Modules.scala 50:57:@58409.4]
  assign _T_103531 = $signed(buffer_0_228) + $signed(buffer_1_229); // @[Modules.scala 50:57:@58427.4]
  assign _T_103532 = _T_103531[10:0]; // @[Modules.scala 50:57:@58428.4]
  assign buffer_15_506 = $signed(_T_103532); // @[Modules.scala 50:57:@58429.4]
  assign _T_103534 = $signed(buffer_1_230) + $signed(buffer_4_231); // @[Modules.scala 50:57:@58431.4]
  assign _T_103535 = _T_103534[10:0]; // @[Modules.scala 50:57:@58432.4]
  assign buffer_15_507 = $signed(_T_103535); // @[Modules.scala 50:57:@58433.4]
  assign _T_103558 = $signed(buffer_0_246) + $signed(buffer_1_247); // @[Modules.scala 50:57:@58463.4]
  assign _T_103559 = _T_103558[10:0]; // @[Modules.scala 50:57:@58464.4]
  assign buffer_15_515 = $signed(_T_103559); // @[Modules.scala 50:57:@58465.4]
  assign buffer_15_249 = {{6{_T_102498[4]}},_T_102498}; // @[Modules.scala 32:22:@8.4]
  assign _T_103561 = $signed(buffer_13_248) + $signed(buffer_15_249); // @[Modules.scala 50:57:@58467.4]
  assign _T_103562 = _T_103561[10:0]; // @[Modules.scala 50:57:@58468.4]
  assign buffer_15_516 = $signed(_T_103562); // @[Modules.scala 50:57:@58469.4]
  assign _T_103582 = $signed(buffer_2_262) + $signed(buffer_7_263); // @[Modules.scala 50:57:@58495.4]
  assign _T_103583 = _T_103582[10:0]; // @[Modules.scala 50:57:@58496.4]
  assign buffer_15_523 = $signed(_T_103583); // @[Modules.scala 50:57:@58497.4]
  assign _T_103597 = $signed(buffer_1_272) + $signed(buffer_3_273); // @[Modules.scala 50:57:@58515.4]
  assign _T_103598 = _T_103597[10:0]; // @[Modules.scala 50:57:@58516.4]
  assign buffer_15_528 = $signed(_T_103598); // @[Modules.scala 50:57:@58517.4]
  assign _T_103600 = $signed(buffer_2_274) + $signed(buffer_0_275); // @[Modules.scala 50:57:@58519.4]
  assign _T_103601 = _T_103600[10:0]; // @[Modules.scala 50:57:@58520.4]
  assign buffer_15_529 = $signed(_T_103601); // @[Modules.scala 50:57:@58521.4]
  assign _T_103615 = $signed(buffer_0_284) + $signed(buffer_1_285); // @[Modules.scala 50:57:@58539.4]
  assign _T_103616 = _T_103615[10:0]; // @[Modules.scala 50:57:@58540.4]
  assign buffer_15_534 = $signed(_T_103616); // @[Modules.scala 50:57:@58541.4]
  assign buffer_15_287 = {{6{_T_102672[4]}},_T_102672}; // @[Modules.scala 32:22:@8.4]
  assign _T_103618 = $signed(buffer_1_286) + $signed(buffer_15_287); // @[Modules.scala 50:57:@58543.4]
  assign _T_103619 = _T_103618[10:0]; // @[Modules.scala 50:57:@58544.4]
  assign buffer_15_535 = $signed(_T_103619); // @[Modules.scala 50:57:@58545.4]
  assign _T_103621 = $signed(buffer_0_288) + $signed(buffer_5_289); // @[Modules.scala 50:57:@58547.4]
  assign _T_103622 = _T_103621[10:0]; // @[Modules.scala 50:57:@58548.4]
  assign buffer_15_536 = $signed(_T_103622); // @[Modules.scala 50:57:@58549.4]
  assign _T_103630 = $signed(buffer_2_294) + $signed(buffer_0_295); // @[Modules.scala 50:57:@58559.4]
  assign _T_103631 = _T_103630[10:0]; // @[Modules.scala 50:57:@58560.4]
  assign buffer_15_539 = $signed(_T_103631); // @[Modules.scala 50:57:@58561.4]
  assign _T_103636 = $signed(buffer_0_298) + $signed(buffer_7_299); // @[Modules.scala 50:57:@58567.4]
  assign _T_103637 = _T_103636[10:0]; // @[Modules.scala 50:57:@58568.4]
  assign buffer_15_541 = $signed(_T_103637); // @[Modules.scala 50:57:@58569.4]
  assign _T_103639 = $signed(buffer_2_300) + $signed(buffer_0_301); // @[Modules.scala 50:57:@58571.4]
  assign _T_103640 = _T_103639[10:0]; // @[Modules.scala 50:57:@58572.4]
  assign buffer_15_542 = $signed(_T_103640); // @[Modules.scala 50:57:@58573.4]
  assign _T_103642 = $signed(buffer_5_302) + $signed(buffer_8_303); // @[Modules.scala 50:57:@58575.4]
  assign _T_103643 = _T_103642[10:0]; // @[Modules.scala 50:57:@58576.4]
  assign buffer_15_543 = $signed(_T_103643); // @[Modules.scala 50:57:@58577.4]
  assign _T_103645 = $signed(buffer_0_304) + $signed(buffer_3_305); // @[Modules.scala 50:57:@58579.4]
  assign _T_103646 = _T_103645[10:0]; // @[Modules.scala 50:57:@58580.4]
  assign buffer_15_544 = $signed(_T_103646); // @[Modules.scala 50:57:@58581.4]
  assign buffer_15_308 = {{6{_T_102771[4]}},_T_102771}; // @[Modules.scala 32:22:@8.4]
  assign _T_103651 = $signed(buffer_15_308) + $signed(buffer_2_309); // @[Modules.scala 50:57:@58587.4]
  assign _T_103652 = _T_103651[10:0]; // @[Modules.scala 50:57:@58588.4]
  assign buffer_15_546 = $signed(_T_103652); // @[Modules.scala 50:57:@58589.4]
  assign _T_103654 = $signed(buffer_11_310) + $signed(buffer_0_311); // @[Modules.scala 50:57:@58591.4]
  assign _T_103655 = _T_103654[10:0]; // @[Modules.scala 50:57:@58592.4]
  assign buffer_15_547 = $signed(_T_103655); // @[Modules.scala 50:57:@58593.4]
  assign _T_103660 = $signed(buffer_0_314) + $signed(buffer_1_315); // @[Modules.scala 50:57:@58599.4]
  assign _T_103661 = _T_103660[10:0]; // @[Modules.scala 50:57:@58600.4]
  assign buffer_15_549 = $signed(_T_103661); // @[Modules.scala 50:57:@58601.4]
  assign _T_103669 = $signed(buffer_0_320) + $signed(buffer_1_321); // @[Modules.scala 50:57:@58611.4]
  assign _T_103670 = _T_103669[10:0]; // @[Modules.scala 50:57:@58612.4]
  assign buffer_15_552 = $signed(_T_103670); // @[Modules.scala 50:57:@58613.4]
  assign _T_103672 = $signed(buffer_0_322) + $signed(buffer_6_323); // @[Modules.scala 50:57:@58615.4]
  assign _T_103673 = _T_103672[10:0]; // @[Modules.scala 50:57:@58616.4]
  assign buffer_15_553 = $signed(_T_103673); // @[Modules.scala 50:57:@58617.4]
  assign _T_103675 = $signed(buffer_0_324) + $signed(buffer_3_325); // @[Modules.scala 50:57:@58619.4]
  assign _T_103676 = _T_103675[10:0]; // @[Modules.scala 50:57:@58620.4]
  assign buffer_15_554 = $signed(_T_103676); // @[Modules.scala 50:57:@58621.4]
  assign buffer_15_338 = {{6{_T_102937[4]}},_T_102937}; // @[Modules.scala 32:22:@8.4]
  assign _T_103696 = $signed(buffer_15_338) + $signed(buffer_2_339); // @[Modules.scala 50:57:@58647.4]
  assign _T_103697 = _T_103696[10:0]; // @[Modules.scala 50:57:@58648.4]
  assign buffer_15_561 = $signed(_T_103697); // @[Modules.scala 50:57:@58649.4]
  assign _T_103699 = $signed(buffer_2_340) + $signed(buffer_1_341); // @[Modules.scala 50:57:@58651.4]
  assign _T_103700 = _T_103699[10:0]; // @[Modules.scala 50:57:@58652.4]
  assign buffer_15_562 = $signed(_T_103700); // @[Modules.scala 50:57:@58653.4]
  assign _T_103714 = $signed(buffer_1_350) + $signed(buffer_5_351); // @[Modules.scala 50:57:@58671.4]
  assign _T_103715 = _T_103714[10:0]; // @[Modules.scala 50:57:@58672.4]
  assign buffer_15_567 = $signed(_T_103715); // @[Modules.scala 50:57:@58673.4]
  assign _T_103717 = $signed(buffer_0_352) + $signed(buffer_2_353); // @[Modules.scala 50:57:@58675.4]
  assign _T_103718 = _T_103717[10:0]; // @[Modules.scala 50:57:@58676.4]
  assign buffer_15_568 = $signed(_T_103718); // @[Modules.scala 50:57:@58677.4]
  assign buffer_15_356 = {{6{_T_103035[4]}},_T_103035}; // @[Modules.scala 32:22:@8.4]
  assign _T_103723 = $signed(buffer_15_356) + $signed(buffer_2_357); // @[Modules.scala 50:57:@58683.4]
  assign _T_103724 = _T_103723[10:0]; // @[Modules.scala 50:57:@58684.4]
  assign buffer_15_570 = $signed(_T_103724); // @[Modules.scala 50:57:@58685.4]
  assign buffer_15_366 = {{6{_T_103089[4]}},_T_103089}; // @[Modules.scala 32:22:@8.4]
  assign _T_103738 = $signed(buffer_15_366) + $signed(buffer_0_367); // @[Modules.scala 50:57:@58703.4]
  assign _T_103739 = _T_103738[10:0]; // @[Modules.scala 50:57:@58704.4]
  assign buffer_15_575 = $signed(_T_103739); // @[Modules.scala 50:57:@58705.4]
  assign buffer_15_389 = {{6{_T_103178[4]}},_T_103178}; // @[Modules.scala 32:22:@8.4]
  assign _T_103771 = $signed(buffer_0_388) + $signed(buffer_15_389); // @[Modules.scala 50:57:@58747.4]
  assign _T_103772 = _T_103771[10:0]; // @[Modules.scala 50:57:@58748.4]
  assign buffer_15_586 = $signed(_T_103772); // @[Modules.scala 50:57:@58749.4]
  assign _T_103777 = $signed(buffer_14_392) + $signed(buffer_0_393); // @[Modules.scala 53:83:@58755.4]
  assign _T_103778 = _T_103777[10:0]; // @[Modules.scala 53:83:@58756.4]
  assign buffer_15_588 = $signed(_T_103778); // @[Modules.scala 53:83:@58757.4]
  assign _T_103780 = $signed(buffer_8_394) + $signed(buffer_15_395); // @[Modules.scala 53:83:@58759.4]
  assign _T_103781 = _T_103780[10:0]; // @[Modules.scala 53:83:@58760.4]
  assign buffer_15_589 = $signed(_T_103781); // @[Modules.scala 53:83:@58761.4]
  assign _T_103783 = $signed(buffer_15_396) + $signed(buffer_15_397); // @[Modules.scala 53:83:@58763.4]
  assign _T_103784 = _T_103783[10:0]; // @[Modules.scala 53:83:@58764.4]
  assign buffer_15_590 = $signed(_T_103784); // @[Modules.scala 53:83:@58765.4]
  assign _T_103786 = $signed(buffer_15_398) + $signed(buffer_12_399); // @[Modules.scala 53:83:@58767.4]
  assign _T_103787 = _T_103786[10:0]; // @[Modules.scala 53:83:@58768.4]
  assign buffer_15_591 = $signed(_T_103787); // @[Modules.scala 53:83:@58769.4]
  assign _T_103789 = $signed(buffer_2_400) + $signed(buffer_15_401); // @[Modules.scala 53:83:@58771.4]
  assign _T_103790 = _T_103789[10:0]; // @[Modules.scala 53:83:@58772.4]
  assign buffer_15_592 = $signed(_T_103790); // @[Modules.scala 53:83:@58773.4]
  assign _T_103792 = $signed(buffer_1_402) + $signed(buffer_15_403); // @[Modules.scala 53:83:@58775.4]
  assign _T_103793 = _T_103792[10:0]; // @[Modules.scala 53:83:@58776.4]
  assign buffer_15_593 = $signed(_T_103793); // @[Modules.scala 53:83:@58777.4]
  assign _T_103795 = $signed(buffer_15_404) + $signed(buffer_15_405); // @[Modules.scala 53:83:@58779.4]
  assign _T_103796 = _T_103795[10:0]; // @[Modules.scala 53:83:@58780.4]
  assign buffer_15_594 = $signed(_T_103796); // @[Modules.scala 53:83:@58781.4]
  assign _T_103798 = $signed(buffer_5_406) + $signed(buffer_1_407); // @[Modules.scala 53:83:@58783.4]
  assign _T_103799 = _T_103798[10:0]; // @[Modules.scala 53:83:@58784.4]
  assign buffer_15_595 = $signed(_T_103799); // @[Modules.scala 53:83:@58785.4]
  assign _T_103804 = $signed(buffer_1_410) + $signed(buffer_15_411); // @[Modules.scala 53:83:@58791.4]
  assign _T_103805 = _T_103804[10:0]; // @[Modules.scala 53:83:@58792.4]
  assign buffer_15_597 = $signed(_T_103805); // @[Modules.scala 53:83:@58793.4]
  assign _T_103807 = $signed(buffer_3_412) + $signed(buffer_15_413); // @[Modules.scala 53:83:@58795.4]
  assign _T_103808 = _T_103807[10:0]; // @[Modules.scala 53:83:@58796.4]
  assign buffer_15_598 = $signed(_T_103808); // @[Modules.scala 53:83:@58797.4]
  assign _T_103810 = $signed(buffer_15_414) + $signed(buffer_1_415); // @[Modules.scala 53:83:@58799.4]
  assign _T_103811 = _T_103810[10:0]; // @[Modules.scala 53:83:@58800.4]
  assign buffer_15_599 = $signed(_T_103811); // @[Modules.scala 53:83:@58801.4]
  assign _T_103819 = $signed(buffer_0_420) + $signed(buffer_12_421); // @[Modules.scala 53:83:@58811.4]
  assign _T_103820 = _T_103819[10:0]; // @[Modules.scala 53:83:@58812.4]
  assign buffer_15_602 = $signed(_T_103820); // @[Modules.scala 53:83:@58813.4]
  assign _T_103822 = $signed(buffer_15_422) + $signed(buffer_14_423); // @[Modules.scala 53:83:@58815.4]
  assign _T_103823 = _T_103822[10:0]; // @[Modules.scala 53:83:@58816.4]
  assign buffer_15_603 = $signed(_T_103823); // @[Modules.scala 53:83:@58817.4]
  assign _T_103825 = $signed(buffer_15_424) + $signed(buffer_0_425); // @[Modules.scala 53:83:@58819.4]
  assign _T_103826 = _T_103825[10:0]; // @[Modules.scala 53:83:@58820.4]
  assign buffer_15_604 = $signed(_T_103826); // @[Modules.scala 53:83:@58821.4]
  assign _T_103828 = $signed(buffer_12_426) + $signed(buffer_15_427); // @[Modules.scala 53:83:@58823.4]
  assign _T_103829 = _T_103828[10:0]; // @[Modules.scala 53:83:@58824.4]
  assign buffer_15_605 = $signed(_T_103829); // @[Modules.scala 53:83:@58825.4]
  assign _T_103831 = $signed(buffer_1_428) + $signed(buffer_0_429); // @[Modules.scala 53:83:@58827.4]
  assign _T_103832 = _T_103831[10:0]; // @[Modules.scala 53:83:@58828.4]
  assign buffer_15_606 = $signed(_T_103832); // @[Modules.scala 53:83:@58829.4]
  assign _T_103834 = $signed(buffer_15_430) + $signed(buffer_15_431); // @[Modules.scala 53:83:@58831.4]
  assign _T_103835 = _T_103834[10:0]; // @[Modules.scala 53:83:@58832.4]
  assign buffer_15_607 = $signed(_T_103835); // @[Modules.scala 53:83:@58833.4]
  assign _T_103837 = $signed(buffer_5_432) + $signed(buffer_15_433); // @[Modules.scala 53:83:@58835.4]
  assign _T_103838 = _T_103837[10:0]; // @[Modules.scala 53:83:@58836.4]
  assign buffer_15_608 = $signed(_T_103838); // @[Modules.scala 53:83:@58837.4]
  assign _T_103840 = $signed(buffer_15_434) + $signed(buffer_15_435); // @[Modules.scala 53:83:@58839.4]
  assign _T_103841 = _T_103840[10:0]; // @[Modules.scala 53:83:@58840.4]
  assign buffer_15_609 = $signed(_T_103841); // @[Modules.scala 53:83:@58841.4]
  assign _T_103843 = $signed(buffer_15_436) + $signed(buffer_1_437); // @[Modules.scala 53:83:@58843.4]
  assign _T_103844 = _T_103843[10:0]; // @[Modules.scala 53:83:@58844.4]
  assign buffer_15_610 = $signed(_T_103844); // @[Modules.scala 53:83:@58845.4]
  assign _T_103846 = $signed(buffer_4_438) + $signed(buffer_6_439); // @[Modules.scala 53:83:@58847.4]
  assign _T_103847 = _T_103846[10:0]; // @[Modules.scala 53:83:@58848.4]
  assign buffer_15_611 = $signed(_T_103847); // @[Modules.scala 53:83:@58849.4]
  assign _T_103849 = $signed(buffer_0_440) + $signed(buffer_15_441); // @[Modules.scala 53:83:@58851.4]
  assign _T_103850 = _T_103849[10:0]; // @[Modules.scala 53:83:@58852.4]
  assign buffer_15_612 = $signed(_T_103850); // @[Modules.scala 53:83:@58853.4]
  assign _T_103852 = $signed(buffer_15_442) + $signed(buffer_1_443); // @[Modules.scala 53:83:@58855.4]
  assign _T_103853 = _T_103852[10:0]; // @[Modules.scala 53:83:@58856.4]
  assign buffer_15_613 = $signed(_T_103853); // @[Modules.scala 53:83:@58857.4]
  assign _T_103855 = $signed(buffer_6_444) + $signed(buffer_15_445); // @[Modules.scala 53:83:@58859.4]
  assign _T_103856 = _T_103855[10:0]; // @[Modules.scala 53:83:@58860.4]
  assign buffer_15_614 = $signed(_T_103856); // @[Modules.scala 53:83:@58861.4]
  assign _T_103858 = $signed(buffer_9_446) + $signed(buffer_0_447); // @[Modules.scala 53:83:@58863.4]
  assign _T_103859 = _T_103858[10:0]; // @[Modules.scala 53:83:@58864.4]
  assign buffer_15_615 = $signed(_T_103859); // @[Modules.scala 53:83:@58865.4]
  assign _T_103861 = $signed(buffer_3_448) + $signed(buffer_13_449); // @[Modules.scala 53:83:@58867.4]
  assign _T_103862 = _T_103861[10:0]; // @[Modules.scala 53:83:@58868.4]
  assign buffer_15_616 = $signed(_T_103862); // @[Modules.scala 53:83:@58869.4]
  assign _T_103864 = $signed(buffer_15_450) + $signed(buffer_12_451); // @[Modules.scala 53:83:@58871.4]
  assign _T_103865 = _T_103864[10:0]; // @[Modules.scala 53:83:@58872.4]
  assign buffer_15_617 = $signed(_T_103865); // @[Modules.scala 53:83:@58873.4]
  assign _T_103867 = $signed(buffer_6_452) + $signed(buffer_9_453); // @[Modules.scala 53:83:@58875.4]
  assign _T_103868 = _T_103867[10:0]; // @[Modules.scala 53:83:@58876.4]
  assign buffer_15_618 = $signed(_T_103868); // @[Modules.scala 53:83:@58877.4]
  assign _T_103873 = $signed(buffer_15_456) + $signed(buffer_12_457); // @[Modules.scala 53:83:@58883.4]
  assign _T_103874 = _T_103873[10:0]; // @[Modules.scala 53:83:@58884.4]
  assign buffer_15_620 = $signed(_T_103874); // @[Modules.scala 53:83:@58885.4]
  assign _T_103876 = $signed(buffer_5_458) + $signed(buffer_3_459); // @[Modules.scala 53:83:@58887.4]
  assign _T_103877 = _T_103876[10:0]; // @[Modules.scala 53:83:@58888.4]
  assign buffer_15_621 = $signed(_T_103877); // @[Modules.scala 53:83:@58889.4]
  assign _T_103882 = $signed(buffer_3_462) + $signed(buffer_15_463); // @[Modules.scala 53:83:@58895.4]
  assign _T_103883 = _T_103882[10:0]; // @[Modules.scala 53:83:@58896.4]
  assign buffer_15_623 = $signed(_T_103883); // @[Modules.scala 53:83:@58897.4]
  assign _T_103888 = $signed(buffer_3_466) + $signed(buffer_15_467); // @[Modules.scala 53:83:@58903.4]
  assign _T_103889 = _T_103888[10:0]; // @[Modules.scala 53:83:@58904.4]
  assign buffer_15_625 = $signed(_T_103889); // @[Modules.scala 53:83:@58905.4]
  assign _T_103891 = $signed(buffer_0_468) + $signed(buffer_10_469); // @[Modules.scala 53:83:@58907.4]
  assign _T_103892 = _T_103891[10:0]; // @[Modules.scala 53:83:@58908.4]
  assign buffer_15_626 = $signed(_T_103892); // @[Modules.scala 53:83:@58909.4]
  assign _T_103894 = $signed(buffer_15_470) + $signed(buffer_15_471); // @[Modules.scala 53:83:@58911.4]
  assign _T_103895 = _T_103894[10:0]; // @[Modules.scala 53:83:@58912.4]
  assign buffer_15_627 = $signed(_T_103895); // @[Modules.scala 53:83:@58913.4]
  assign _T_103897 = $signed(buffer_0_472) + $signed(buffer_15_473); // @[Modules.scala 53:83:@58915.4]
  assign _T_103898 = _T_103897[10:0]; // @[Modules.scala 53:83:@58916.4]
  assign buffer_15_628 = $signed(_T_103898); // @[Modules.scala 53:83:@58917.4]
  assign _T_103900 = $signed(buffer_5_474) + $signed(buffer_6_475); // @[Modules.scala 53:83:@58919.4]
  assign _T_103901 = _T_103900[10:0]; // @[Modules.scala 53:83:@58920.4]
  assign buffer_15_629 = $signed(_T_103901); // @[Modules.scala 53:83:@58921.4]
  assign _T_103903 = $signed(buffer_15_476) + $signed(buffer_6_477); // @[Modules.scala 53:83:@58923.4]
  assign _T_103904 = _T_103903[10:0]; // @[Modules.scala 53:83:@58924.4]
  assign buffer_15_630 = $signed(_T_103904); // @[Modules.scala 53:83:@58925.4]
  assign _T_103909 = $signed(buffer_9_480) + $signed(buffer_0_481); // @[Modules.scala 53:83:@58931.4]
  assign _T_103910 = _T_103909[10:0]; // @[Modules.scala 53:83:@58932.4]
  assign buffer_15_632 = $signed(_T_103910); // @[Modules.scala 53:83:@58933.4]
  assign _T_103912 = $signed(buffer_15_482) + $signed(buffer_15_483); // @[Modules.scala 53:83:@58935.4]
  assign _T_103913 = _T_103912[10:0]; // @[Modules.scala 53:83:@58936.4]
  assign buffer_15_633 = $signed(_T_103913); // @[Modules.scala 53:83:@58937.4]
  assign _T_103915 = $signed(buffer_15_484) + $signed(buffer_9_485); // @[Modules.scala 53:83:@58939.4]
  assign _T_103916 = _T_103915[10:0]; // @[Modules.scala 53:83:@58940.4]
  assign buffer_15_634 = $signed(_T_103916); // @[Modules.scala 53:83:@58941.4]
  assign _T_103921 = $signed(buffer_4_488) + $signed(buffer_9_489); // @[Modules.scala 53:83:@58947.4]
  assign _T_103922 = _T_103921[10:0]; // @[Modules.scala 53:83:@58948.4]
  assign buffer_15_636 = $signed(_T_103922); // @[Modules.scala 53:83:@58949.4]
  assign _T_103927 = $signed(buffer_5_492) + $signed(buffer_3_493); // @[Modules.scala 53:83:@58955.4]
  assign _T_103928 = _T_103927[10:0]; // @[Modules.scala 53:83:@58956.4]
  assign buffer_15_638 = $signed(_T_103928); // @[Modules.scala 53:83:@58957.4]
  assign _T_103930 = $signed(buffer_15_494) + $signed(buffer_0_495); // @[Modules.scala 53:83:@58959.4]
  assign _T_103931 = _T_103930[10:0]; // @[Modules.scala 53:83:@58960.4]
  assign buffer_15_639 = $signed(_T_103931); // @[Modules.scala 53:83:@58961.4]
  assign _T_103933 = $signed(buffer_10_496) + $signed(buffer_7_497); // @[Modules.scala 53:83:@58963.4]
  assign _T_103934 = _T_103933[10:0]; // @[Modules.scala 53:83:@58964.4]
  assign buffer_15_640 = $signed(_T_103934); // @[Modules.scala 53:83:@58965.4]
  assign _T_103939 = $signed(buffer_1_500) + $signed(buffer_15_501); // @[Modules.scala 53:83:@58971.4]
  assign _T_103940 = _T_103939[10:0]; // @[Modules.scala 53:83:@58972.4]
  assign buffer_15_642 = $signed(_T_103940); // @[Modules.scala 53:83:@58973.4]
  assign _T_103942 = $signed(buffer_1_502) + $signed(buffer_3_503); // @[Modules.scala 53:83:@58975.4]
  assign _T_103943 = _T_103942[10:0]; // @[Modules.scala 53:83:@58976.4]
  assign buffer_15_643 = $signed(_T_103943); // @[Modules.scala 53:83:@58977.4]
  assign _T_103948 = $signed(buffer_15_506) + $signed(buffer_15_507); // @[Modules.scala 53:83:@58983.4]
  assign _T_103949 = _T_103948[10:0]; // @[Modules.scala 53:83:@58984.4]
  assign buffer_15_645 = $signed(_T_103949); // @[Modules.scala 53:83:@58985.4]
  assign _T_103951 = $signed(buffer_0_508) + $signed(buffer_10_509); // @[Modules.scala 53:83:@58987.4]
  assign _T_103952 = _T_103951[10:0]; // @[Modules.scala 53:83:@58988.4]
  assign buffer_15_646 = $signed(_T_103952); // @[Modules.scala 53:83:@58989.4]
  assign _T_103960 = $signed(buffer_2_514) + $signed(buffer_15_515); // @[Modules.scala 53:83:@58999.4]
  assign _T_103961 = _T_103960[10:0]; // @[Modules.scala 53:83:@59000.4]
  assign buffer_15_649 = $signed(_T_103961); // @[Modules.scala 53:83:@59001.4]
  assign _T_103963 = $signed(buffer_15_516) + $signed(buffer_3_517); // @[Modules.scala 53:83:@59003.4]
  assign _T_103964 = _T_103963[10:0]; // @[Modules.scala 53:83:@59004.4]
  assign buffer_15_650 = $signed(_T_103964); // @[Modules.scala 53:83:@59005.4]
  assign _T_103966 = $signed(buffer_12_518) + $signed(buffer_8_519); // @[Modules.scala 53:83:@59007.4]
  assign _T_103967 = _T_103966[10:0]; // @[Modules.scala 53:83:@59008.4]
  assign buffer_15_651 = $signed(_T_103967); // @[Modules.scala 53:83:@59009.4]
  assign _T_103969 = $signed(buffer_0_520) + $signed(buffer_2_521); // @[Modules.scala 53:83:@59011.4]
  assign _T_103970 = _T_103969[10:0]; // @[Modules.scala 53:83:@59012.4]
  assign buffer_15_652 = $signed(_T_103970); // @[Modules.scala 53:83:@59013.4]
  assign _T_103972 = $signed(buffer_5_522) + $signed(buffer_15_523); // @[Modules.scala 53:83:@59015.4]
  assign _T_103973 = _T_103972[10:0]; // @[Modules.scala 53:83:@59016.4]
  assign buffer_15_653 = $signed(_T_103973); // @[Modules.scala 53:83:@59017.4]
  assign _T_103978 = $signed(buffer_0_526) + $signed(buffer_1_527); // @[Modules.scala 53:83:@59023.4]
  assign _T_103979 = _T_103978[10:0]; // @[Modules.scala 53:83:@59024.4]
  assign buffer_15_655 = $signed(_T_103979); // @[Modules.scala 53:83:@59025.4]
  assign _T_103981 = $signed(buffer_15_528) + $signed(buffer_15_529); // @[Modules.scala 53:83:@59027.4]
  assign _T_103982 = _T_103981[10:0]; // @[Modules.scala 53:83:@59028.4]
  assign buffer_15_656 = $signed(_T_103982); // @[Modules.scala 53:83:@59029.4]
  assign _T_103990 = $signed(buffer_15_534) + $signed(buffer_15_535); // @[Modules.scala 53:83:@59039.4]
  assign _T_103991 = _T_103990[10:0]; // @[Modules.scala 53:83:@59040.4]
  assign buffer_15_659 = $signed(_T_103991); // @[Modules.scala 53:83:@59041.4]
  assign _T_103993 = $signed(buffer_15_536) + $signed(buffer_10_537); // @[Modules.scala 53:83:@59043.4]
  assign _T_103994 = _T_103993[10:0]; // @[Modules.scala 53:83:@59044.4]
  assign buffer_15_660 = $signed(_T_103994); // @[Modules.scala 53:83:@59045.4]
  assign _T_103996 = $signed(buffer_8_538) + $signed(buffer_15_539); // @[Modules.scala 53:83:@59047.4]
  assign _T_103997 = _T_103996[10:0]; // @[Modules.scala 53:83:@59048.4]
  assign buffer_15_661 = $signed(_T_103997); // @[Modules.scala 53:83:@59049.4]
  assign _T_103999 = $signed(buffer_11_540) + $signed(buffer_15_541); // @[Modules.scala 53:83:@59051.4]
  assign _T_104000 = _T_103999[10:0]; // @[Modules.scala 53:83:@59052.4]
  assign buffer_15_662 = $signed(_T_104000); // @[Modules.scala 53:83:@59053.4]
  assign _T_104002 = $signed(buffer_15_542) + $signed(buffer_15_543); // @[Modules.scala 53:83:@59055.4]
  assign _T_104003 = _T_104002[10:0]; // @[Modules.scala 53:83:@59056.4]
  assign buffer_15_663 = $signed(_T_104003); // @[Modules.scala 53:83:@59057.4]
  assign _T_104005 = $signed(buffer_15_544) + $signed(buffer_10_545); // @[Modules.scala 53:83:@59059.4]
  assign _T_104006 = _T_104005[10:0]; // @[Modules.scala 53:83:@59060.4]
  assign buffer_15_664 = $signed(_T_104006); // @[Modules.scala 53:83:@59061.4]
  assign _T_104008 = $signed(buffer_15_546) + $signed(buffer_15_547); // @[Modules.scala 53:83:@59063.4]
  assign _T_104009 = _T_104008[10:0]; // @[Modules.scala 53:83:@59064.4]
  assign buffer_15_665 = $signed(_T_104009); // @[Modules.scala 53:83:@59065.4]
  assign _T_104011 = $signed(buffer_8_548) + $signed(buffer_15_549); // @[Modules.scala 53:83:@59067.4]
  assign _T_104012 = _T_104011[10:0]; // @[Modules.scala 53:83:@59068.4]
  assign buffer_15_666 = $signed(_T_104012); // @[Modules.scala 53:83:@59069.4]
  assign _T_104017 = $signed(buffer_15_552) + $signed(buffer_15_553); // @[Modules.scala 53:83:@59075.4]
  assign _T_104018 = _T_104017[10:0]; // @[Modules.scala 53:83:@59076.4]
  assign buffer_15_668 = $signed(_T_104018); // @[Modules.scala 53:83:@59077.4]
  assign _T_104020 = $signed(buffer_15_554) + $signed(buffer_8_555); // @[Modules.scala 53:83:@59079.4]
  assign _T_104021 = _T_104020[10:0]; // @[Modules.scala 53:83:@59080.4]
  assign buffer_15_669 = $signed(_T_104021); // @[Modules.scala 53:83:@59081.4]
  assign _T_104026 = $signed(buffer_5_558) + $signed(buffer_3_559); // @[Modules.scala 53:83:@59087.4]
  assign _T_104027 = _T_104026[10:0]; // @[Modules.scala 53:83:@59088.4]
  assign buffer_15_671 = $signed(_T_104027); // @[Modules.scala 53:83:@59089.4]
  assign _T_104029 = $signed(buffer_6_560) + $signed(buffer_15_561); // @[Modules.scala 53:83:@59091.4]
  assign _T_104030 = _T_104029[10:0]; // @[Modules.scala 53:83:@59092.4]
  assign buffer_15_672 = $signed(_T_104030); // @[Modules.scala 53:83:@59093.4]
  assign _T_104032 = $signed(buffer_15_562) + $signed(buffer_3_563); // @[Modules.scala 53:83:@59095.4]
  assign _T_104033 = _T_104032[10:0]; // @[Modules.scala 53:83:@59096.4]
  assign buffer_15_673 = $signed(_T_104033); // @[Modules.scala 53:83:@59097.4]
  assign _T_104038 = $signed(buffer_12_566) + $signed(buffer_15_567); // @[Modules.scala 53:83:@59103.4]
  assign _T_104039 = _T_104038[10:0]; // @[Modules.scala 53:83:@59104.4]
  assign buffer_15_675 = $signed(_T_104039); // @[Modules.scala 53:83:@59105.4]
  assign _T_104041 = $signed(buffer_15_568) + $signed(buffer_6_569); // @[Modules.scala 53:83:@59107.4]
  assign _T_104042 = _T_104041[10:0]; // @[Modules.scala 53:83:@59108.4]
  assign buffer_15_676 = $signed(_T_104042); // @[Modules.scala 53:83:@59109.4]
  assign _T_104044 = $signed(buffer_15_570) + $signed(buffer_1_571); // @[Modules.scala 53:83:@59111.4]
  assign _T_104045 = _T_104044[10:0]; // @[Modules.scala 53:83:@59112.4]
  assign buffer_15_677 = $signed(_T_104045); // @[Modules.scala 53:83:@59113.4]
  assign _T_104050 = $signed(buffer_3_574) + $signed(buffer_15_575); // @[Modules.scala 53:83:@59119.4]
  assign _T_104051 = _T_104050[10:0]; // @[Modules.scala 53:83:@59120.4]
  assign buffer_15_679 = $signed(_T_104051); // @[Modules.scala 53:83:@59121.4]
  assign _T_104068 = $signed(buffer_15_586) + $signed(buffer_13_587); // @[Modules.scala 53:83:@59143.4]
  assign _T_104069 = _T_104068[10:0]; // @[Modules.scala 53:83:@59144.4]
  assign buffer_15_685 = $signed(_T_104069); // @[Modules.scala 53:83:@59145.4]
  assign _T_104071 = $signed(buffer_15_588) + $signed(buffer_15_589); // @[Modules.scala 56:109:@59147.4]
  assign _T_104072 = _T_104071[10:0]; // @[Modules.scala 56:109:@59148.4]
  assign buffer_15_686 = $signed(_T_104072); // @[Modules.scala 56:109:@59149.4]
  assign _T_104074 = $signed(buffer_15_590) + $signed(buffer_15_591); // @[Modules.scala 56:109:@59151.4]
  assign _T_104075 = _T_104074[10:0]; // @[Modules.scala 56:109:@59152.4]
  assign buffer_15_687 = $signed(_T_104075); // @[Modules.scala 56:109:@59153.4]
  assign _T_104077 = $signed(buffer_15_592) + $signed(buffer_15_593); // @[Modules.scala 56:109:@59155.4]
  assign _T_104078 = _T_104077[10:0]; // @[Modules.scala 56:109:@59156.4]
  assign buffer_15_688 = $signed(_T_104078); // @[Modules.scala 56:109:@59157.4]
  assign _T_104080 = $signed(buffer_15_594) + $signed(buffer_15_595); // @[Modules.scala 56:109:@59159.4]
  assign _T_104081 = _T_104080[10:0]; // @[Modules.scala 56:109:@59160.4]
  assign buffer_15_689 = $signed(_T_104081); // @[Modules.scala 56:109:@59161.4]
  assign _T_104083 = $signed(buffer_1_596) + $signed(buffer_15_597); // @[Modules.scala 56:109:@59163.4]
  assign _T_104084 = _T_104083[10:0]; // @[Modules.scala 56:109:@59164.4]
  assign buffer_15_690 = $signed(_T_104084); // @[Modules.scala 56:109:@59165.4]
  assign _T_104086 = $signed(buffer_15_598) + $signed(buffer_15_599); // @[Modules.scala 56:109:@59167.4]
  assign _T_104087 = _T_104086[10:0]; // @[Modules.scala 56:109:@59168.4]
  assign buffer_15_691 = $signed(_T_104087); // @[Modules.scala 56:109:@59169.4]
  assign _T_104092 = $signed(buffer_15_602) + $signed(buffer_15_603); // @[Modules.scala 56:109:@59175.4]
  assign _T_104093 = _T_104092[10:0]; // @[Modules.scala 56:109:@59176.4]
  assign buffer_15_693 = $signed(_T_104093); // @[Modules.scala 56:109:@59177.4]
  assign _T_104095 = $signed(buffer_15_604) + $signed(buffer_15_605); // @[Modules.scala 56:109:@59179.4]
  assign _T_104096 = _T_104095[10:0]; // @[Modules.scala 56:109:@59180.4]
  assign buffer_15_694 = $signed(_T_104096); // @[Modules.scala 56:109:@59181.4]
  assign _T_104098 = $signed(buffer_15_606) + $signed(buffer_15_607); // @[Modules.scala 56:109:@59183.4]
  assign _T_104099 = _T_104098[10:0]; // @[Modules.scala 56:109:@59184.4]
  assign buffer_15_695 = $signed(_T_104099); // @[Modules.scala 56:109:@59185.4]
  assign _T_104101 = $signed(buffer_15_608) + $signed(buffer_15_609); // @[Modules.scala 56:109:@59187.4]
  assign _T_104102 = _T_104101[10:0]; // @[Modules.scala 56:109:@59188.4]
  assign buffer_15_696 = $signed(_T_104102); // @[Modules.scala 56:109:@59189.4]
  assign _T_104104 = $signed(buffer_15_610) + $signed(buffer_15_611); // @[Modules.scala 56:109:@59191.4]
  assign _T_104105 = _T_104104[10:0]; // @[Modules.scala 56:109:@59192.4]
  assign buffer_15_697 = $signed(_T_104105); // @[Modules.scala 56:109:@59193.4]
  assign _T_104107 = $signed(buffer_15_612) + $signed(buffer_15_613); // @[Modules.scala 56:109:@59195.4]
  assign _T_104108 = _T_104107[10:0]; // @[Modules.scala 56:109:@59196.4]
  assign buffer_15_698 = $signed(_T_104108); // @[Modules.scala 56:109:@59197.4]
  assign _T_104110 = $signed(buffer_15_614) + $signed(buffer_15_615); // @[Modules.scala 56:109:@59199.4]
  assign _T_104111 = _T_104110[10:0]; // @[Modules.scala 56:109:@59200.4]
  assign buffer_15_699 = $signed(_T_104111); // @[Modules.scala 56:109:@59201.4]
  assign _T_104113 = $signed(buffer_15_616) + $signed(buffer_15_617); // @[Modules.scala 56:109:@59203.4]
  assign _T_104114 = _T_104113[10:0]; // @[Modules.scala 56:109:@59204.4]
  assign buffer_15_700 = $signed(_T_104114); // @[Modules.scala 56:109:@59205.4]
  assign _T_104116 = $signed(buffer_15_618) + $signed(buffer_10_619); // @[Modules.scala 56:109:@59207.4]
  assign _T_104117 = _T_104116[10:0]; // @[Modules.scala 56:109:@59208.4]
  assign buffer_15_701 = $signed(_T_104117); // @[Modules.scala 56:109:@59209.4]
  assign _T_104119 = $signed(buffer_15_620) + $signed(buffer_15_621); // @[Modules.scala 56:109:@59211.4]
  assign _T_104120 = _T_104119[10:0]; // @[Modules.scala 56:109:@59212.4]
  assign buffer_15_702 = $signed(_T_104120); // @[Modules.scala 56:109:@59213.4]
  assign _T_104122 = $signed(buffer_0_622) + $signed(buffer_15_623); // @[Modules.scala 56:109:@59215.4]
  assign _T_104123 = _T_104122[10:0]; // @[Modules.scala 56:109:@59216.4]
  assign buffer_15_703 = $signed(_T_104123); // @[Modules.scala 56:109:@59217.4]
  assign _T_104125 = $signed(buffer_5_624) + $signed(buffer_15_625); // @[Modules.scala 56:109:@59219.4]
  assign _T_104126 = _T_104125[10:0]; // @[Modules.scala 56:109:@59220.4]
  assign buffer_15_704 = $signed(_T_104126); // @[Modules.scala 56:109:@59221.4]
  assign _T_104128 = $signed(buffer_15_626) + $signed(buffer_15_627); // @[Modules.scala 56:109:@59223.4]
  assign _T_104129 = _T_104128[10:0]; // @[Modules.scala 56:109:@59224.4]
  assign buffer_15_705 = $signed(_T_104129); // @[Modules.scala 56:109:@59225.4]
  assign _T_104131 = $signed(buffer_15_628) + $signed(buffer_15_629); // @[Modules.scala 56:109:@59227.4]
  assign _T_104132 = _T_104131[10:0]; // @[Modules.scala 56:109:@59228.4]
  assign buffer_15_706 = $signed(_T_104132); // @[Modules.scala 56:109:@59229.4]
  assign _T_104134 = $signed(buffer_15_630) + $signed(buffer_3_631); // @[Modules.scala 56:109:@59231.4]
  assign _T_104135 = _T_104134[10:0]; // @[Modules.scala 56:109:@59232.4]
  assign buffer_15_707 = $signed(_T_104135); // @[Modules.scala 56:109:@59233.4]
  assign _T_104137 = $signed(buffer_15_632) + $signed(buffer_15_633); // @[Modules.scala 56:109:@59235.4]
  assign _T_104138 = _T_104137[10:0]; // @[Modules.scala 56:109:@59236.4]
  assign buffer_15_708 = $signed(_T_104138); // @[Modules.scala 56:109:@59237.4]
  assign _T_104140 = $signed(buffer_15_634) + $signed(buffer_12_635); // @[Modules.scala 56:109:@59239.4]
  assign _T_104141 = _T_104140[10:0]; // @[Modules.scala 56:109:@59240.4]
  assign buffer_15_709 = $signed(_T_104141); // @[Modules.scala 56:109:@59241.4]
  assign _T_104143 = $signed(buffer_15_636) + $signed(buffer_8_637); // @[Modules.scala 56:109:@59243.4]
  assign _T_104144 = _T_104143[10:0]; // @[Modules.scala 56:109:@59244.4]
  assign buffer_15_710 = $signed(_T_104144); // @[Modules.scala 56:109:@59245.4]
  assign _T_104146 = $signed(buffer_15_638) + $signed(buffer_15_639); // @[Modules.scala 56:109:@59247.4]
  assign _T_104147 = _T_104146[10:0]; // @[Modules.scala 56:109:@59248.4]
  assign buffer_15_711 = $signed(_T_104147); // @[Modules.scala 56:109:@59249.4]
  assign _T_104149 = $signed(buffer_15_640) + $signed(buffer_8_641); // @[Modules.scala 56:109:@59251.4]
  assign _T_104150 = _T_104149[10:0]; // @[Modules.scala 56:109:@59252.4]
  assign buffer_15_712 = $signed(_T_104150); // @[Modules.scala 56:109:@59253.4]
  assign _T_104152 = $signed(buffer_15_642) + $signed(buffer_15_643); // @[Modules.scala 56:109:@59255.4]
  assign _T_104153 = _T_104152[10:0]; // @[Modules.scala 56:109:@59256.4]
  assign buffer_15_713 = $signed(_T_104153); // @[Modules.scala 56:109:@59257.4]
  assign _T_104155 = $signed(buffer_8_644) + $signed(buffer_15_645); // @[Modules.scala 56:109:@59259.4]
  assign _T_104156 = _T_104155[10:0]; // @[Modules.scala 56:109:@59260.4]
  assign buffer_15_714 = $signed(_T_104156); // @[Modules.scala 56:109:@59261.4]
  assign _T_104158 = $signed(buffer_15_646) + $signed(buffer_7_647); // @[Modules.scala 56:109:@59263.4]
  assign _T_104159 = _T_104158[10:0]; // @[Modules.scala 56:109:@59264.4]
  assign buffer_15_715 = $signed(_T_104159); // @[Modules.scala 56:109:@59265.4]
  assign _T_104161 = $signed(buffer_12_648) + $signed(buffer_15_649); // @[Modules.scala 56:109:@59267.4]
  assign _T_104162 = _T_104161[10:0]; // @[Modules.scala 56:109:@59268.4]
  assign buffer_15_716 = $signed(_T_104162); // @[Modules.scala 56:109:@59269.4]
  assign _T_104164 = $signed(buffer_15_650) + $signed(buffer_15_651); // @[Modules.scala 56:109:@59271.4]
  assign _T_104165 = _T_104164[10:0]; // @[Modules.scala 56:109:@59272.4]
  assign buffer_15_717 = $signed(_T_104165); // @[Modules.scala 56:109:@59273.4]
  assign _T_104167 = $signed(buffer_15_652) + $signed(buffer_15_653); // @[Modules.scala 56:109:@59275.4]
  assign _T_104168 = _T_104167[10:0]; // @[Modules.scala 56:109:@59276.4]
  assign buffer_15_718 = $signed(_T_104168); // @[Modules.scala 56:109:@59277.4]
  assign _T_104170 = $signed(buffer_12_654) + $signed(buffer_15_655); // @[Modules.scala 56:109:@59279.4]
  assign _T_104171 = _T_104170[10:0]; // @[Modules.scala 56:109:@59280.4]
  assign buffer_15_719 = $signed(_T_104171); // @[Modules.scala 56:109:@59281.4]
  assign _T_104173 = $signed(buffer_15_656) + $signed(buffer_8_657); // @[Modules.scala 56:109:@59283.4]
  assign _T_104174 = _T_104173[10:0]; // @[Modules.scala 56:109:@59284.4]
  assign buffer_15_720 = $signed(_T_104174); // @[Modules.scala 56:109:@59285.4]
  assign _T_104176 = $signed(buffer_2_658) + $signed(buffer_15_659); // @[Modules.scala 56:109:@59287.4]
  assign _T_104177 = _T_104176[10:0]; // @[Modules.scala 56:109:@59288.4]
  assign buffer_15_721 = $signed(_T_104177); // @[Modules.scala 56:109:@59289.4]
  assign _T_104179 = $signed(buffer_15_660) + $signed(buffer_15_661); // @[Modules.scala 56:109:@59291.4]
  assign _T_104180 = _T_104179[10:0]; // @[Modules.scala 56:109:@59292.4]
  assign buffer_15_722 = $signed(_T_104180); // @[Modules.scala 56:109:@59293.4]
  assign _T_104182 = $signed(buffer_15_662) + $signed(buffer_15_663); // @[Modules.scala 56:109:@59295.4]
  assign _T_104183 = _T_104182[10:0]; // @[Modules.scala 56:109:@59296.4]
  assign buffer_15_723 = $signed(_T_104183); // @[Modules.scala 56:109:@59297.4]
  assign _T_104185 = $signed(buffer_15_664) + $signed(buffer_15_665); // @[Modules.scala 56:109:@59299.4]
  assign _T_104186 = _T_104185[10:0]; // @[Modules.scala 56:109:@59300.4]
  assign buffer_15_724 = $signed(_T_104186); // @[Modules.scala 56:109:@59301.4]
  assign _T_104188 = $signed(buffer_15_666) + $signed(buffer_3_667); // @[Modules.scala 56:109:@59303.4]
  assign _T_104189 = _T_104188[10:0]; // @[Modules.scala 56:109:@59304.4]
  assign buffer_15_725 = $signed(_T_104189); // @[Modules.scala 56:109:@59305.4]
  assign _T_104191 = $signed(buffer_15_668) + $signed(buffer_15_669); // @[Modules.scala 56:109:@59307.4]
  assign _T_104192 = _T_104191[10:0]; // @[Modules.scala 56:109:@59308.4]
  assign buffer_15_726 = $signed(_T_104192); // @[Modules.scala 56:109:@59309.4]
  assign _T_104194 = $signed(buffer_0_670) + $signed(buffer_15_671); // @[Modules.scala 56:109:@59311.4]
  assign _T_104195 = _T_104194[10:0]; // @[Modules.scala 56:109:@59312.4]
  assign buffer_15_727 = $signed(_T_104195); // @[Modules.scala 56:109:@59313.4]
  assign _T_104197 = $signed(buffer_15_672) + $signed(buffer_15_673); // @[Modules.scala 56:109:@59315.4]
  assign _T_104198 = _T_104197[10:0]; // @[Modules.scala 56:109:@59316.4]
  assign buffer_15_728 = $signed(_T_104198); // @[Modules.scala 56:109:@59317.4]
  assign _T_104200 = $signed(buffer_3_674) + $signed(buffer_15_675); // @[Modules.scala 56:109:@59319.4]
  assign _T_104201 = _T_104200[10:0]; // @[Modules.scala 56:109:@59320.4]
  assign buffer_15_729 = $signed(_T_104201); // @[Modules.scala 56:109:@59321.4]
  assign _T_104203 = $signed(buffer_15_676) + $signed(buffer_15_677); // @[Modules.scala 56:109:@59323.4]
  assign _T_104204 = _T_104203[10:0]; // @[Modules.scala 56:109:@59324.4]
  assign buffer_15_730 = $signed(_T_104204); // @[Modules.scala 56:109:@59325.4]
  assign _T_104206 = $signed(buffer_9_678) + $signed(buffer_15_679); // @[Modules.scala 56:109:@59327.4]
  assign _T_104207 = _T_104206[10:0]; // @[Modules.scala 56:109:@59328.4]
  assign buffer_15_731 = $signed(_T_104207); // @[Modules.scala 56:109:@59329.4]
  assign _T_104209 = $signed(buffer_5_680) + $signed(buffer_3_681); // @[Modules.scala 56:109:@59331.4]
  assign _T_104210 = _T_104209[10:0]; // @[Modules.scala 56:109:@59332.4]
  assign buffer_15_732 = $signed(_T_104210); // @[Modules.scala 56:109:@59333.4]
  assign _T_104212 = $signed(buffer_8_682) + $signed(buffer_10_683); // @[Modules.scala 56:109:@59335.4]
  assign _T_104213 = _T_104212[10:0]; // @[Modules.scala 56:109:@59336.4]
  assign buffer_15_733 = $signed(_T_104213); // @[Modules.scala 56:109:@59337.4]
  assign _T_104215 = $signed(buffer_3_684) + $signed(buffer_15_685); // @[Modules.scala 56:109:@59339.4]
  assign _T_104216 = _T_104215[10:0]; // @[Modules.scala 56:109:@59340.4]
  assign buffer_15_734 = $signed(_T_104216); // @[Modules.scala 56:109:@59341.4]
  assign _T_104218 = $signed(buffer_15_686) + $signed(buffer_15_687); // @[Modules.scala 63:156:@59344.4]
  assign _T_104219 = _T_104218[10:0]; // @[Modules.scala 63:156:@59345.4]
  assign buffer_15_736 = $signed(_T_104219); // @[Modules.scala 63:156:@59346.4]
  assign _T_104221 = $signed(buffer_15_736) + $signed(buffer_15_688); // @[Modules.scala 63:156:@59348.4]
  assign _T_104222 = _T_104221[10:0]; // @[Modules.scala 63:156:@59349.4]
  assign buffer_15_737 = $signed(_T_104222); // @[Modules.scala 63:156:@59350.4]
  assign _T_104224 = $signed(buffer_15_737) + $signed(buffer_15_689); // @[Modules.scala 63:156:@59352.4]
  assign _T_104225 = _T_104224[10:0]; // @[Modules.scala 63:156:@59353.4]
  assign buffer_15_738 = $signed(_T_104225); // @[Modules.scala 63:156:@59354.4]
  assign _T_104227 = $signed(buffer_15_738) + $signed(buffer_15_690); // @[Modules.scala 63:156:@59356.4]
  assign _T_104228 = _T_104227[10:0]; // @[Modules.scala 63:156:@59357.4]
  assign buffer_15_739 = $signed(_T_104228); // @[Modules.scala 63:156:@59358.4]
  assign _T_104230 = $signed(buffer_15_739) + $signed(buffer_15_691); // @[Modules.scala 63:156:@59360.4]
  assign _T_104231 = _T_104230[10:0]; // @[Modules.scala 63:156:@59361.4]
  assign buffer_15_740 = $signed(_T_104231); // @[Modules.scala 63:156:@59362.4]
  assign _T_104233 = $signed(buffer_15_740) + $signed(buffer_12_692); // @[Modules.scala 63:156:@59364.4]
  assign _T_104234 = _T_104233[10:0]; // @[Modules.scala 63:156:@59365.4]
  assign buffer_15_741 = $signed(_T_104234); // @[Modules.scala 63:156:@59366.4]
  assign _T_104236 = $signed(buffer_15_741) + $signed(buffer_15_693); // @[Modules.scala 63:156:@59368.4]
  assign _T_104237 = _T_104236[10:0]; // @[Modules.scala 63:156:@59369.4]
  assign buffer_15_742 = $signed(_T_104237); // @[Modules.scala 63:156:@59370.4]
  assign _T_104239 = $signed(buffer_15_742) + $signed(buffer_15_694); // @[Modules.scala 63:156:@59372.4]
  assign _T_104240 = _T_104239[10:0]; // @[Modules.scala 63:156:@59373.4]
  assign buffer_15_743 = $signed(_T_104240); // @[Modules.scala 63:156:@59374.4]
  assign _T_104242 = $signed(buffer_15_743) + $signed(buffer_15_695); // @[Modules.scala 63:156:@59376.4]
  assign _T_104243 = _T_104242[10:0]; // @[Modules.scala 63:156:@59377.4]
  assign buffer_15_744 = $signed(_T_104243); // @[Modules.scala 63:156:@59378.4]
  assign _T_104245 = $signed(buffer_15_744) + $signed(buffer_15_696); // @[Modules.scala 63:156:@59380.4]
  assign _T_104246 = _T_104245[10:0]; // @[Modules.scala 63:156:@59381.4]
  assign buffer_15_745 = $signed(_T_104246); // @[Modules.scala 63:156:@59382.4]
  assign _T_104248 = $signed(buffer_15_745) + $signed(buffer_15_697); // @[Modules.scala 63:156:@59384.4]
  assign _T_104249 = _T_104248[10:0]; // @[Modules.scala 63:156:@59385.4]
  assign buffer_15_746 = $signed(_T_104249); // @[Modules.scala 63:156:@59386.4]
  assign _T_104251 = $signed(buffer_15_746) + $signed(buffer_15_698); // @[Modules.scala 63:156:@59388.4]
  assign _T_104252 = _T_104251[10:0]; // @[Modules.scala 63:156:@59389.4]
  assign buffer_15_747 = $signed(_T_104252); // @[Modules.scala 63:156:@59390.4]
  assign _T_104254 = $signed(buffer_15_747) + $signed(buffer_15_699); // @[Modules.scala 63:156:@59392.4]
  assign _T_104255 = _T_104254[10:0]; // @[Modules.scala 63:156:@59393.4]
  assign buffer_15_748 = $signed(_T_104255); // @[Modules.scala 63:156:@59394.4]
  assign _T_104257 = $signed(buffer_15_748) + $signed(buffer_15_700); // @[Modules.scala 63:156:@59396.4]
  assign _T_104258 = _T_104257[10:0]; // @[Modules.scala 63:156:@59397.4]
  assign buffer_15_749 = $signed(_T_104258); // @[Modules.scala 63:156:@59398.4]
  assign _T_104260 = $signed(buffer_15_749) + $signed(buffer_15_701); // @[Modules.scala 63:156:@59400.4]
  assign _T_104261 = _T_104260[10:0]; // @[Modules.scala 63:156:@59401.4]
  assign buffer_15_750 = $signed(_T_104261); // @[Modules.scala 63:156:@59402.4]
  assign _T_104263 = $signed(buffer_15_750) + $signed(buffer_15_702); // @[Modules.scala 63:156:@59404.4]
  assign _T_104264 = _T_104263[10:0]; // @[Modules.scala 63:156:@59405.4]
  assign buffer_15_751 = $signed(_T_104264); // @[Modules.scala 63:156:@59406.4]
  assign _T_104266 = $signed(buffer_15_751) + $signed(buffer_15_703); // @[Modules.scala 63:156:@59408.4]
  assign _T_104267 = _T_104266[10:0]; // @[Modules.scala 63:156:@59409.4]
  assign buffer_15_752 = $signed(_T_104267); // @[Modules.scala 63:156:@59410.4]
  assign _T_104269 = $signed(buffer_15_752) + $signed(buffer_15_704); // @[Modules.scala 63:156:@59412.4]
  assign _T_104270 = _T_104269[10:0]; // @[Modules.scala 63:156:@59413.4]
  assign buffer_15_753 = $signed(_T_104270); // @[Modules.scala 63:156:@59414.4]
  assign _T_104272 = $signed(buffer_15_753) + $signed(buffer_15_705); // @[Modules.scala 63:156:@59416.4]
  assign _T_104273 = _T_104272[10:0]; // @[Modules.scala 63:156:@59417.4]
  assign buffer_15_754 = $signed(_T_104273); // @[Modules.scala 63:156:@59418.4]
  assign _T_104275 = $signed(buffer_15_754) + $signed(buffer_15_706); // @[Modules.scala 63:156:@59420.4]
  assign _T_104276 = _T_104275[10:0]; // @[Modules.scala 63:156:@59421.4]
  assign buffer_15_755 = $signed(_T_104276); // @[Modules.scala 63:156:@59422.4]
  assign _T_104278 = $signed(buffer_15_755) + $signed(buffer_15_707); // @[Modules.scala 63:156:@59424.4]
  assign _T_104279 = _T_104278[10:0]; // @[Modules.scala 63:156:@59425.4]
  assign buffer_15_756 = $signed(_T_104279); // @[Modules.scala 63:156:@59426.4]
  assign _T_104281 = $signed(buffer_15_756) + $signed(buffer_15_708); // @[Modules.scala 63:156:@59428.4]
  assign _T_104282 = _T_104281[10:0]; // @[Modules.scala 63:156:@59429.4]
  assign buffer_15_757 = $signed(_T_104282); // @[Modules.scala 63:156:@59430.4]
  assign _T_104284 = $signed(buffer_15_757) + $signed(buffer_15_709); // @[Modules.scala 63:156:@59432.4]
  assign _T_104285 = _T_104284[10:0]; // @[Modules.scala 63:156:@59433.4]
  assign buffer_15_758 = $signed(_T_104285); // @[Modules.scala 63:156:@59434.4]
  assign _T_104287 = $signed(buffer_15_758) + $signed(buffer_15_710); // @[Modules.scala 63:156:@59436.4]
  assign _T_104288 = _T_104287[10:0]; // @[Modules.scala 63:156:@59437.4]
  assign buffer_15_759 = $signed(_T_104288); // @[Modules.scala 63:156:@59438.4]
  assign _T_104290 = $signed(buffer_15_759) + $signed(buffer_15_711); // @[Modules.scala 63:156:@59440.4]
  assign _T_104291 = _T_104290[10:0]; // @[Modules.scala 63:156:@59441.4]
  assign buffer_15_760 = $signed(_T_104291); // @[Modules.scala 63:156:@59442.4]
  assign _T_104293 = $signed(buffer_15_760) + $signed(buffer_15_712); // @[Modules.scala 63:156:@59444.4]
  assign _T_104294 = _T_104293[10:0]; // @[Modules.scala 63:156:@59445.4]
  assign buffer_15_761 = $signed(_T_104294); // @[Modules.scala 63:156:@59446.4]
  assign _T_104296 = $signed(buffer_15_761) + $signed(buffer_15_713); // @[Modules.scala 63:156:@59448.4]
  assign _T_104297 = _T_104296[10:0]; // @[Modules.scala 63:156:@59449.4]
  assign buffer_15_762 = $signed(_T_104297); // @[Modules.scala 63:156:@59450.4]
  assign _T_104299 = $signed(buffer_15_762) + $signed(buffer_15_714); // @[Modules.scala 63:156:@59452.4]
  assign _T_104300 = _T_104299[10:0]; // @[Modules.scala 63:156:@59453.4]
  assign buffer_15_763 = $signed(_T_104300); // @[Modules.scala 63:156:@59454.4]
  assign _T_104302 = $signed(buffer_15_763) + $signed(buffer_15_715); // @[Modules.scala 63:156:@59456.4]
  assign _T_104303 = _T_104302[10:0]; // @[Modules.scala 63:156:@59457.4]
  assign buffer_15_764 = $signed(_T_104303); // @[Modules.scala 63:156:@59458.4]
  assign _T_104305 = $signed(buffer_15_764) + $signed(buffer_15_716); // @[Modules.scala 63:156:@59460.4]
  assign _T_104306 = _T_104305[10:0]; // @[Modules.scala 63:156:@59461.4]
  assign buffer_15_765 = $signed(_T_104306); // @[Modules.scala 63:156:@59462.4]
  assign _T_104308 = $signed(buffer_15_765) + $signed(buffer_15_717); // @[Modules.scala 63:156:@59464.4]
  assign _T_104309 = _T_104308[10:0]; // @[Modules.scala 63:156:@59465.4]
  assign buffer_15_766 = $signed(_T_104309); // @[Modules.scala 63:156:@59466.4]
  assign _T_104311 = $signed(buffer_15_766) + $signed(buffer_15_718); // @[Modules.scala 63:156:@59468.4]
  assign _T_104312 = _T_104311[10:0]; // @[Modules.scala 63:156:@59469.4]
  assign buffer_15_767 = $signed(_T_104312); // @[Modules.scala 63:156:@59470.4]
  assign _T_104314 = $signed(buffer_15_767) + $signed(buffer_15_719); // @[Modules.scala 63:156:@59472.4]
  assign _T_104315 = _T_104314[10:0]; // @[Modules.scala 63:156:@59473.4]
  assign buffer_15_768 = $signed(_T_104315); // @[Modules.scala 63:156:@59474.4]
  assign _T_104317 = $signed(buffer_15_768) + $signed(buffer_15_720); // @[Modules.scala 63:156:@59476.4]
  assign _T_104318 = _T_104317[10:0]; // @[Modules.scala 63:156:@59477.4]
  assign buffer_15_769 = $signed(_T_104318); // @[Modules.scala 63:156:@59478.4]
  assign _T_104320 = $signed(buffer_15_769) + $signed(buffer_15_721); // @[Modules.scala 63:156:@59480.4]
  assign _T_104321 = _T_104320[10:0]; // @[Modules.scala 63:156:@59481.4]
  assign buffer_15_770 = $signed(_T_104321); // @[Modules.scala 63:156:@59482.4]
  assign _T_104323 = $signed(buffer_15_770) + $signed(buffer_15_722); // @[Modules.scala 63:156:@59484.4]
  assign _T_104324 = _T_104323[10:0]; // @[Modules.scala 63:156:@59485.4]
  assign buffer_15_771 = $signed(_T_104324); // @[Modules.scala 63:156:@59486.4]
  assign _T_104326 = $signed(buffer_15_771) + $signed(buffer_15_723); // @[Modules.scala 63:156:@59488.4]
  assign _T_104327 = _T_104326[10:0]; // @[Modules.scala 63:156:@59489.4]
  assign buffer_15_772 = $signed(_T_104327); // @[Modules.scala 63:156:@59490.4]
  assign _T_104329 = $signed(buffer_15_772) + $signed(buffer_15_724); // @[Modules.scala 63:156:@59492.4]
  assign _T_104330 = _T_104329[10:0]; // @[Modules.scala 63:156:@59493.4]
  assign buffer_15_773 = $signed(_T_104330); // @[Modules.scala 63:156:@59494.4]
  assign _T_104332 = $signed(buffer_15_773) + $signed(buffer_15_725); // @[Modules.scala 63:156:@59496.4]
  assign _T_104333 = _T_104332[10:0]; // @[Modules.scala 63:156:@59497.4]
  assign buffer_15_774 = $signed(_T_104333); // @[Modules.scala 63:156:@59498.4]
  assign _T_104335 = $signed(buffer_15_774) + $signed(buffer_15_726); // @[Modules.scala 63:156:@59500.4]
  assign _T_104336 = _T_104335[10:0]; // @[Modules.scala 63:156:@59501.4]
  assign buffer_15_775 = $signed(_T_104336); // @[Modules.scala 63:156:@59502.4]
  assign _T_104338 = $signed(buffer_15_775) + $signed(buffer_15_727); // @[Modules.scala 63:156:@59504.4]
  assign _T_104339 = _T_104338[10:0]; // @[Modules.scala 63:156:@59505.4]
  assign buffer_15_776 = $signed(_T_104339); // @[Modules.scala 63:156:@59506.4]
  assign _T_104341 = $signed(buffer_15_776) + $signed(buffer_15_728); // @[Modules.scala 63:156:@59508.4]
  assign _T_104342 = _T_104341[10:0]; // @[Modules.scala 63:156:@59509.4]
  assign buffer_15_777 = $signed(_T_104342); // @[Modules.scala 63:156:@59510.4]
  assign _T_104344 = $signed(buffer_15_777) + $signed(buffer_15_729); // @[Modules.scala 63:156:@59512.4]
  assign _T_104345 = _T_104344[10:0]; // @[Modules.scala 63:156:@59513.4]
  assign buffer_15_778 = $signed(_T_104345); // @[Modules.scala 63:156:@59514.4]
  assign _T_104347 = $signed(buffer_15_778) + $signed(buffer_15_730); // @[Modules.scala 63:156:@59516.4]
  assign _T_104348 = _T_104347[10:0]; // @[Modules.scala 63:156:@59517.4]
  assign buffer_15_779 = $signed(_T_104348); // @[Modules.scala 63:156:@59518.4]
  assign _T_104350 = $signed(buffer_15_779) + $signed(buffer_15_731); // @[Modules.scala 63:156:@59520.4]
  assign _T_104351 = _T_104350[10:0]; // @[Modules.scala 63:156:@59521.4]
  assign buffer_15_780 = $signed(_T_104351); // @[Modules.scala 63:156:@59522.4]
  assign _T_104353 = $signed(buffer_15_780) + $signed(buffer_15_732); // @[Modules.scala 63:156:@59524.4]
  assign _T_104354 = _T_104353[10:0]; // @[Modules.scala 63:156:@59525.4]
  assign buffer_15_781 = $signed(_T_104354); // @[Modules.scala 63:156:@59526.4]
  assign _T_104356 = $signed(buffer_15_781) + $signed(buffer_15_733); // @[Modules.scala 63:156:@59528.4]
  assign _T_104357 = _T_104356[10:0]; // @[Modules.scala 63:156:@59529.4]
  assign buffer_15_782 = $signed(_T_104357); // @[Modules.scala 63:156:@59530.4]
  assign _T_104359 = $signed(buffer_15_782) + $signed(buffer_15_734); // @[Modules.scala 63:156:@59532.4]
  assign _T_104360 = _T_104359[10:0]; // @[Modules.scala 63:156:@59533.4]
  assign buffer_15_783 = $signed(_T_104360); // @[Modules.scala 63:156:@59534.4]
  assign io_out_0 = buffer_0_783;
  assign io_out_1 = buffer_1_783;
  assign io_out_2 = buffer_2_783;
  assign io_out_3 = buffer_3_783;
  assign io_out_4 = buffer_4_783;
  assign io_out_5 = buffer_5_783;
  assign io_out_6 = buffer_6_783;
  assign io_out_7 = buffer_7_783;
  assign io_out_8 = buffer_8_783;
  assign io_out_9 = buffer_9_783;
  assign io_out_10 = buffer_10_783;
  assign io_out_11 = buffer_11_783;
  assign io_out_12 = buffer_12_783;
  assign io_out_13 = buffer_13_783;
  assign io_out_14 = buffer_14_783;
  assign io_out_15 = buffer_15_783;
endmodule
