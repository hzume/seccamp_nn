`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Ex( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [3:0] io_in_0, // @[:@6.4]
  input  [3:0] io_in_1, // @[:@6.4]
  input  [3:0] io_in_2, // @[:@6.4]
  input  [3:0] io_in_3, // @[:@6.4]
  input  [3:0] io_in_4, // @[:@6.4]
  input  [3:0] io_in_5, // @[:@6.4]
  input  [3:0] io_in_6, // @[:@6.4]
  input  [3:0] io_in_7, // @[:@6.4]
  input  [3:0] io_in_8, // @[:@6.4]
  input  [3:0] io_in_9, // @[:@6.4]
  input  [3:0] io_in_10, // @[:@6.4]
  input  [3:0] io_in_11, // @[:@6.4]
  input  [3:0] io_in_12, // @[:@6.4]
  input  [3:0] io_in_13, // @[:@6.4]
  input  [3:0] io_in_14, // @[:@6.4]
  input  [3:0] io_in_15, // @[:@6.4]
  input  [3:0] io_in_16, // @[:@6.4]
  input  [3:0] io_in_17, // @[:@6.4]
  input  [3:0] io_in_18, // @[:@6.4]
  input  [3:0] io_in_19, // @[:@6.4]
  input  [3:0] io_in_20, // @[:@6.4]
  input  [3:0] io_in_21, // @[:@6.4]
  input  [3:0] io_in_22, // @[:@6.4]
  input  [3:0] io_in_23, // @[:@6.4]
  input  [3:0] io_in_24, // @[:@6.4]
  input  [3:0] io_in_25, // @[:@6.4]
  input  [3:0] io_in_26, // @[:@6.4]
  input  [3:0] io_in_27, // @[:@6.4]
  input  [3:0] io_in_28, // @[:@6.4]
  input  [3:0] io_in_29, // @[:@6.4]
  input  [3:0] io_in_30, // @[:@6.4]
  input  [3:0] io_in_31, // @[:@6.4]
  input  [3:0] io_in_32, // @[:@6.4]
  input  [3:0] io_in_33, // @[:@6.4]
  input  [3:0] io_in_34, // @[:@6.4]
  input  [3:0] io_in_35, // @[:@6.4]
  input  [3:0] io_in_36, // @[:@6.4]
  input  [3:0] io_in_37, // @[:@6.4]
  input  [3:0] io_in_38, // @[:@6.4]
  input  [3:0] io_in_39, // @[:@6.4]
  input  [3:0] io_in_40, // @[:@6.4]
  input  [3:0] io_in_41, // @[:@6.4]
  input  [3:0] io_in_42, // @[:@6.4]
  input  [3:0] io_in_43, // @[:@6.4]
  input  [3:0] io_in_44, // @[:@6.4]
  input  [3:0] io_in_45, // @[:@6.4]
  input  [3:0] io_in_46, // @[:@6.4]
  input  [3:0] io_in_47, // @[:@6.4]
  input  [3:0] io_in_48, // @[:@6.4]
  input  [3:0] io_in_49, // @[:@6.4]
  input  [3:0] io_in_50, // @[:@6.4]
  input  [3:0] io_in_51, // @[:@6.4]
  input  [3:0] io_in_52, // @[:@6.4]
  input  [3:0] io_in_53, // @[:@6.4]
  input  [3:0] io_in_54, // @[:@6.4]
  input  [3:0] io_in_55, // @[:@6.4]
  input  [3:0] io_in_56, // @[:@6.4]
  input  [3:0] io_in_57, // @[:@6.4]
  input  [3:0] io_in_58, // @[:@6.4]
  input  [3:0] io_in_59, // @[:@6.4]
  input  [3:0] io_in_60, // @[:@6.4]
  input  [3:0] io_in_61, // @[:@6.4]
  input  [3:0] io_in_62, // @[:@6.4]
  input  [3:0] io_in_63, // @[:@6.4]
  input  [3:0] io_in_64, // @[:@6.4]
  input  [3:0] io_in_65, // @[:@6.4]
  input  [3:0] io_in_66, // @[:@6.4]
  input  [3:0] io_in_67, // @[:@6.4]
  input  [3:0] io_in_68, // @[:@6.4]
  input  [3:0] io_in_69, // @[:@6.4]
  input  [3:0] io_in_70, // @[:@6.4]
  input  [3:0] io_in_71, // @[:@6.4]
  input  [3:0] io_in_72, // @[:@6.4]
  input  [3:0] io_in_73, // @[:@6.4]
  input  [3:0] io_in_74, // @[:@6.4]
  input  [3:0] io_in_75, // @[:@6.4]
  input  [3:0] io_in_76, // @[:@6.4]
  input  [3:0] io_in_77, // @[:@6.4]
  input  [3:0] io_in_78, // @[:@6.4]
  input  [3:0] io_in_79, // @[:@6.4]
  input  [3:0] io_in_80, // @[:@6.4]
  input  [3:0] io_in_81, // @[:@6.4]
  input  [3:0] io_in_82, // @[:@6.4]
  input  [3:0] io_in_83, // @[:@6.4]
  input  [3:0] io_in_84, // @[:@6.4]
  input  [3:0] io_in_85, // @[:@6.4]
  input  [3:0] io_in_86, // @[:@6.4]
  input  [3:0] io_in_87, // @[:@6.4]
  input  [3:0] io_in_88, // @[:@6.4]
  input  [3:0] io_in_89, // @[:@6.4]
  input  [3:0] io_in_90, // @[:@6.4]
  input  [3:0] io_in_91, // @[:@6.4]
  input  [3:0] io_in_92, // @[:@6.4]
  input  [3:0] io_in_93, // @[:@6.4]
  input  [3:0] io_in_94, // @[:@6.4]
  input  [3:0] io_in_95, // @[:@6.4]
  input  [3:0] io_in_96, // @[:@6.4]
  input  [3:0] io_in_97, // @[:@6.4]
  input  [3:0] io_in_98, // @[:@6.4]
  input  [3:0] io_in_99, // @[:@6.4]
  input  [3:0] io_in_100, // @[:@6.4]
  input  [3:0] io_in_101, // @[:@6.4]
  input  [3:0] io_in_102, // @[:@6.4]
  input  [3:0] io_in_103, // @[:@6.4]
  input  [3:0] io_in_104, // @[:@6.4]
  input  [3:0] io_in_105, // @[:@6.4]
  input  [3:0] io_in_106, // @[:@6.4]
  input  [3:0] io_in_107, // @[:@6.4]
  input  [3:0] io_in_108, // @[:@6.4]
  input  [3:0] io_in_109, // @[:@6.4]
  input  [3:0] io_in_110, // @[:@6.4]
  input  [3:0] io_in_111, // @[:@6.4]
  input  [3:0] io_in_112, // @[:@6.4]
  input  [3:0] io_in_113, // @[:@6.4]
  input  [3:0] io_in_114, // @[:@6.4]
  input  [3:0] io_in_115, // @[:@6.4]
  input  [3:0] io_in_116, // @[:@6.4]
  input  [3:0] io_in_117, // @[:@6.4]
  input  [3:0] io_in_118, // @[:@6.4]
  input  [3:0] io_in_119, // @[:@6.4]
  input  [3:0] io_in_120, // @[:@6.4]
  input  [3:0] io_in_121, // @[:@6.4]
  input  [3:0] io_in_122, // @[:@6.4]
  input  [3:0] io_in_123, // @[:@6.4]
  input  [3:0] io_in_124, // @[:@6.4]
  input  [3:0] io_in_125, // @[:@6.4]
  input  [3:0] io_in_126, // @[:@6.4]
  input  [3:0] io_in_127, // @[:@6.4]
  input  [3:0] io_in_128, // @[:@6.4]
  input  [3:0] io_in_129, // @[:@6.4]
  input  [3:0] io_in_130, // @[:@6.4]
  input  [3:0] io_in_131, // @[:@6.4]
  input  [3:0] io_in_132, // @[:@6.4]
  input  [3:0] io_in_133, // @[:@6.4]
  input  [3:0] io_in_134, // @[:@6.4]
  input  [3:0] io_in_135, // @[:@6.4]
  input  [3:0] io_in_136, // @[:@6.4]
  input  [3:0] io_in_137, // @[:@6.4]
  input  [3:0] io_in_138, // @[:@6.4]
  input  [3:0] io_in_139, // @[:@6.4]
  input  [3:0] io_in_140, // @[:@6.4]
  input  [3:0] io_in_141, // @[:@6.4]
  input  [3:0] io_in_142, // @[:@6.4]
  input  [3:0] io_in_143, // @[:@6.4]
  input  [3:0] io_in_144, // @[:@6.4]
  input  [3:0] io_in_145, // @[:@6.4]
  input  [3:0] io_in_146, // @[:@6.4]
  input  [3:0] io_in_147, // @[:@6.4]
  input  [3:0] io_in_148, // @[:@6.4]
  input  [3:0] io_in_149, // @[:@6.4]
  input  [3:0] io_in_150, // @[:@6.4]
  input  [3:0] io_in_151, // @[:@6.4]
  input  [3:0] io_in_152, // @[:@6.4]
  input  [3:0] io_in_153, // @[:@6.4]
  input  [3:0] io_in_154, // @[:@6.4]
  input  [3:0] io_in_155, // @[:@6.4]
  input  [3:0] io_in_156, // @[:@6.4]
  input  [3:0] io_in_157, // @[:@6.4]
  input  [3:0] io_in_158, // @[:@6.4]
  input  [3:0] io_in_159, // @[:@6.4]
  input  [3:0] io_in_160, // @[:@6.4]
  input  [3:0] io_in_161, // @[:@6.4]
  input  [3:0] io_in_162, // @[:@6.4]
  input  [3:0] io_in_163, // @[:@6.4]
  input  [3:0] io_in_164, // @[:@6.4]
  input  [3:0] io_in_165, // @[:@6.4]
  input  [3:0] io_in_166, // @[:@6.4]
  input  [3:0] io_in_167, // @[:@6.4]
  input  [3:0] io_in_168, // @[:@6.4]
  input  [3:0] io_in_169, // @[:@6.4]
  input  [3:0] io_in_170, // @[:@6.4]
  input  [3:0] io_in_171, // @[:@6.4]
  input  [3:0] io_in_172, // @[:@6.4]
  input  [3:0] io_in_173, // @[:@6.4]
  input  [3:0] io_in_174, // @[:@6.4]
  input  [3:0] io_in_175, // @[:@6.4]
  input  [3:0] io_in_176, // @[:@6.4]
  input  [3:0] io_in_177, // @[:@6.4]
  input  [3:0] io_in_178, // @[:@6.4]
  input  [3:0] io_in_179, // @[:@6.4]
  input  [3:0] io_in_180, // @[:@6.4]
  input  [3:0] io_in_181, // @[:@6.4]
  input  [3:0] io_in_182, // @[:@6.4]
  input  [3:0] io_in_183, // @[:@6.4]
  input  [3:0] io_in_184, // @[:@6.4]
  input  [3:0] io_in_185, // @[:@6.4]
  input  [3:0] io_in_186, // @[:@6.4]
  input  [3:0] io_in_187, // @[:@6.4]
  input  [3:0] io_in_188, // @[:@6.4]
  input  [3:0] io_in_189, // @[:@6.4]
  input  [3:0] io_in_190, // @[:@6.4]
  input  [3:0] io_in_191, // @[:@6.4]
  input  [3:0] io_in_192, // @[:@6.4]
  input  [3:0] io_in_193, // @[:@6.4]
  input  [3:0] io_in_194, // @[:@6.4]
  input  [3:0] io_in_195, // @[:@6.4]
  input  [3:0] io_in_196, // @[:@6.4]
  input  [3:0] io_in_197, // @[:@6.4]
  input  [3:0] io_in_198, // @[:@6.4]
  input  [3:0] io_in_199, // @[:@6.4]
  input  [3:0] io_in_200, // @[:@6.4]
  input  [3:0] io_in_201, // @[:@6.4]
  input  [3:0] io_in_202, // @[:@6.4]
  input  [3:0] io_in_203, // @[:@6.4]
  input  [3:0] io_in_204, // @[:@6.4]
  input  [3:0] io_in_205, // @[:@6.4]
  input  [3:0] io_in_206, // @[:@6.4]
  input  [3:0] io_in_207, // @[:@6.4]
  input  [3:0] io_in_208, // @[:@6.4]
  input  [3:0] io_in_209, // @[:@6.4]
  input  [3:0] io_in_210, // @[:@6.4]
  input  [3:0] io_in_211, // @[:@6.4]
  input  [3:0] io_in_212, // @[:@6.4]
  input  [3:0] io_in_213, // @[:@6.4]
  input  [3:0] io_in_214, // @[:@6.4]
  input  [3:0] io_in_215, // @[:@6.4]
  input  [3:0] io_in_216, // @[:@6.4]
  input  [3:0] io_in_217, // @[:@6.4]
  input  [3:0] io_in_218, // @[:@6.4]
  input  [3:0] io_in_219, // @[:@6.4]
  input  [3:0] io_in_220, // @[:@6.4]
  input  [3:0] io_in_221, // @[:@6.4]
  input  [3:0] io_in_222, // @[:@6.4]
  input  [3:0] io_in_223, // @[:@6.4]
  input  [3:0] io_in_224, // @[:@6.4]
  input  [3:0] io_in_225, // @[:@6.4]
  input  [3:0] io_in_226, // @[:@6.4]
  input  [3:0] io_in_227, // @[:@6.4]
  input  [3:0] io_in_228, // @[:@6.4]
  input  [3:0] io_in_229, // @[:@6.4]
  input  [3:0] io_in_230, // @[:@6.4]
  input  [3:0] io_in_231, // @[:@6.4]
  input  [3:0] io_in_232, // @[:@6.4]
  input  [3:0] io_in_233, // @[:@6.4]
  input  [3:0] io_in_234, // @[:@6.4]
  input  [3:0] io_in_235, // @[:@6.4]
  input  [3:0] io_in_236, // @[:@6.4]
  input  [3:0] io_in_237, // @[:@6.4]
  input  [3:0] io_in_238, // @[:@6.4]
  input  [3:0] io_in_239, // @[:@6.4]
  input  [3:0] io_in_240, // @[:@6.4]
  input  [3:0] io_in_241, // @[:@6.4]
  input  [3:0] io_in_242, // @[:@6.4]
  input  [3:0] io_in_243, // @[:@6.4]
  input  [3:0] io_in_244, // @[:@6.4]
  input  [3:0] io_in_245, // @[:@6.4]
  input  [3:0] io_in_246, // @[:@6.4]
  input  [3:0] io_in_247, // @[:@6.4]
  input  [3:0] io_in_248, // @[:@6.4]
  input  [3:0] io_in_249, // @[:@6.4]
  input  [3:0] io_in_250, // @[:@6.4]
  input  [3:0] io_in_251, // @[:@6.4]
  input  [3:0] io_in_252, // @[:@6.4]
  input  [3:0] io_in_253, // @[:@6.4]
  input  [3:0] io_in_254, // @[:@6.4]
  input  [3:0] io_in_255, // @[:@6.4]
  input  [3:0] io_in_256, // @[:@6.4]
  input  [3:0] io_in_257, // @[:@6.4]
  input  [3:0] io_in_258, // @[:@6.4]
  input  [3:0] io_in_259, // @[:@6.4]
  input  [3:0] io_in_260, // @[:@6.4]
  input  [3:0] io_in_261, // @[:@6.4]
  input  [3:0] io_in_262, // @[:@6.4]
  input  [3:0] io_in_263, // @[:@6.4]
  input  [3:0] io_in_264, // @[:@6.4]
  input  [3:0] io_in_265, // @[:@6.4]
  input  [3:0] io_in_266, // @[:@6.4]
  input  [3:0] io_in_267, // @[:@6.4]
  input  [3:0] io_in_268, // @[:@6.4]
  input  [3:0] io_in_269, // @[:@6.4]
  input  [3:0] io_in_270, // @[:@6.4]
  input  [3:0] io_in_271, // @[:@6.4]
  input  [3:0] io_in_272, // @[:@6.4]
  input  [3:0] io_in_273, // @[:@6.4]
  input  [3:0] io_in_274, // @[:@6.4]
  input  [3:0] io_in_275, // @[:@6.4]
  input  [3:0] io_in_276, // @[:@6.4]
  input  [3:0] io_in_277, // @[:@6.4]
  input  [3:0] io_in_278, // @[:@6.4]
  input  [3:0] io_in_279, // @[:@6.4]
  input  [3:0] io_in_280, // @[:@6.4]
  input  [3:0] io_in_281, // @[:@6.4]
  input  [3:0] io_in_282, // @[:@6.4]
  input  [3:0] io_in_283, // @[:@6.4]
  input  [3:0] io_in_284, // @[:@6.4]
  input  [3:0] io_in_285, // @[:@6.4]
  input  [3:0] io_in_286, // @[:@6.4]
  input  [3:0] io_in_287, // @[:@6.4]
  input  [3:0] io_in_288, // @[:@6.4]
  input  [3:0] io_in_289, // @[:@6.4]
  input  [3:0] io_in_290, // @[:@6.4]
  input  [3:0] io_in_291, // @[:@6.4]
  input  [3:0] io_in_292, // @[:@6.4]
  input  [3:0] io_in_293, // @[:@6.4]
  input  [3:0] io_in_294, // @[:@6.4]
  input  [3:0] io_in_295, // @[:@6.4]
  input  [3:0] io_in_296, // @[:@6.4]
  input  [3:0] io_in_297, // @[:@6.4]
  input  [3:0] io_in_298, // @[:@6.4]
  input  [3:0] io_in_299, // @[:@6.4]
  input  [3:0] io_in_300, // @[:@6.4]
  input  [3:0] io_in_301, // @[:@6.4]
  input  [3:0] io_in_302, // @[:@6.4]
  input  [3:0] io_in_303, // @[:@6.4]
  input  [3:0] io_in_304, // @[:@6.4]
  input  [3:0] io_in_305, // @[:@6.4]
  input  [3:0] io_in_306, // @[:@6.4]
  input  [3:0] io_in_307, // @[:@6.4]
  input  [3:0] io_in_308, // @[:@6.4]
  input  [3:0] io_in_309, // @[:@6.4]
  input  [3:0] io_in_310, // @[:@6.4]
  input  [3:0] io_in_311, // @[:@6.4]
  input  [3:0] io_in_312, // @[:@6.4]
  input  [3:0] io_in_313, // @[:@6.4]
  input  [3:0] io_in_314, // @[:@6.4]
  input  [3:0] io_in_315, // @[:@6.4]
  input  [3:0] io_in_316, // @[:@6.4]
  input  [3:0] io_in_317, // @[:@6.4]
  input  [3:0] io_in_318, // @[:@6.4]
  input  [3:0] io_in_319, // @[:@6.4]
  input  [3:0] io_in_320, // @[:@6.4]
  input  [3:0] io_in_321, // @[:@6.4]
  input  [3:0] io_in_322, // @[:@6.4]
  input  [3:0] io_in_323, // @[:@6.4]
  input  [3:0] io_in_324, // @[:@6.4]
  input  [3:0] io_in_325, // @[:@6.4]
  input  [3:0] io_in_326, // @[:@6.4]
  input  [3:0] io_in_327, // @[:@6.4]
  input  [3:0] io_in_328, // @[:@6.4]
  input  [3:0] io_in_329, // @[:@6.4]
  input  [3:0] io_in_330, // @[:@6.4]
  input  [3:0] io_in_331, // @[:@6.4]
  input  [3:0] io_in_332, // @[:@6.4]
  input  [3:0] io_in_333, // @[:@6.4]
  input  [3:0] io_in_334, // @[:@6.4]
  input  [3:0] io_in_335, // @[:@6.4]
  input  [3:0] io_in_336, // @[:@6.4]
  input  [3:0] io_in_337, // @[:@6.4]
  input  [3:0] io_in_338, // @[:@6.4]
  input  [3:0] io_in_339, // @[:@6.4]
  input  [3:0] io_in_340, // @[:@6.4]
  input  [3:0] io_in_341, // @[:@6.4]
  input  [3:0] io_in_342, // @[:@6.4]
  input  [3:0] io_in_343, // @[:@6.4]
  input  [3:0] io_in_344, // @[:@6.4]
  input  [3:0] io_in_345, // @[:@6.4]
  input  [3:0] io_in_346, // @[:@6.4]
  input  [3:0] io_in_347, // @[:@6.4]
  input  [3:0] io_in_348, // @[:@6.4]
  input  [3:0] io_in_349, // @[:@6.4]
  input  [3:0] io_in_350, // @[:@6.4]
  input  [3:0] io_in_351, // @[:@6.4]
  input  [3:0] io_in_352, // @[:@6.4]
  input  [3:0] io_in_353, // @[:@6.4]
  input  [3:0] io_in_354, // @[:@6.4]
  input  [3:0] io_in_355, // @[:@6.4]
  input  [3:0] io_in_356, // @[:@6.4]
  input  [3:0] io_in_357, // @[:@6.4]
  input  [3:0] io_in_358, // @[:@6.4]
  input  [3:0] io_in_359, // @[:@6.4]
  input  [3:0] io_in_360, // @[:@6.4]
  input  [3:0] io_in_361, // @[:@6.4]
  input  [3:0] io_in_362, // @[:@6.4]
  input  [3:0] io_in_363, // @[:@6.4]
  input  [3:0] io_in_364, // @[:@6.4]
  input  [3:0] io_in_365, // @[:@6.4]
  input  [3:0] io_in_366, // @[:@6.4]
  input  [3:0] io_in_367, // @[:@6.4]
  input  [3:0] io_in_368, // @[:@6.4]
  input  [3:0] io_in_369, // @[:@6.4]
  input  [3:0] io_in_370, // @[:@6.4]
  input  [3:0] io_in_371, // @[:@6.4]
  input  [3:0] io_in_372, // @[:@6.4]
  input  [3:0] io_in_373, // @[:@6.4]
  input  [3:0] io_in_374, // @[:@6.4]
  input  [3:0] io_in_375, // @[:@6.4]
  input  [3:0] io_in_376, // @[:@6.4]
  input  [3:0] io_in_377, // @[:@6.4]
  input  [3:0] io_in_378, // @[:@6.4]
  input  [3:0] io_in_379, // @[:@6.4]
  input  [3:0] io_in_380, // @[:@6.4]
  input  [3:0] io_in_381, // @[:@6.4]
  input  [3:0] io_in_382, // @[:@6.4]
  input  [3:0] io_in_383, // @[:@6.4]
  input  [3:0] io_in_384, // @[:@6.4]
  input  [3:0] io_in_385, // @[:@6.4]
  input  [3:0] io_in_386, // @[:@6.4]
  input  [3:0] io_in_387, // @[:@6.4]
  input  [3:0] io_in_388, // @[:@6.4]
  input  [3:0] io_in_389, // @[:@6.4]
  input  [3:0] io_in_390, // @[:@6.4]
  input  [3:0] io_in_391, // @[:@6.4]
  input  [3:0] io_in_392, // @[:@6.4]
  input  [3:0] io_in_393, // @[:@6.4]
  input  [3:0] io_in_394, // @[:@6.4]
  input  [3:0] io_in_395, // @[:@6.4]
  input  [3:0] io_in_396, // @[:@6.4]
  input  [3:0] io_in_397, // @[:@6.4]
  input  [3:0] io_in_398, // @[:@6.4]
  input  [3:0] io_in_399, // @[:@6.4]
  input  [3:0] io_in_400, // @[:@6.4]
  input  [3:0] io_in_401, // @[:@6.4]
  input  [3:0] io_in_402, // @[:@6.4]
  input  [3:0] io_in_403, // @[:@6.4]
  input  [3:0] io_in_404, // @[:@6.4]
  input  [3:0] io_in_405, // @[:@6.4]
  input  [3:0] io_in_406, // @[:@6.4]
  input  [3:0] io_in_407, // @[:@6.4]
  input  [3:0] io_in_408, // @[:@6.4]
  input  [3:0] io_in_409, // @[:@6.4]
  input  [3:0] io_in_410, // @[:@6.4]
  input  [3:0] io_in_411, // @[:@6.4]
  input  [3:0] io_in_412, // @[:@6.4]
  input  [3:0] io_in_413, // @[:@6.4]
  input  [3:0] io_in_414, // @[:@6.4]
  input  [3:0] io_in_415, // @[:@6.4]
  input  [3:0] io_in_416, // @[:@6.4]
  input  [3:0] io_in_417, // @[:@6.4]
  input  [3:0] io_in_418, // @[:@6.4]
  input  [3:0] io_in_419, // @[:@6.4]
  input  [3:0] io_in_420, // @[:@6.4]
  input  [3:0] io_in_421, // @[:@6.4]
  input  [3:0] io_in_422, // @[:@6.4]
  input  [3:0] io_in_423, // @[:@6.4]
  input  [3:0] io_in_424, // @[:@6.4]
  input  [3:0] io_in_425, // @[:@6.4]
  input  [3:0] io_in_426, // @[:@6.4]
  input  [3:0] io_in_427, // @[:@6.4]
  input  [3:0] io_in_428, // @[:@6.4]
  input  [3:0] io_in_429, // @[:@6.4]
  input  [3:0] io_in_430, // @[:@6.4]
  input  [3:0] io_in_431, // @[:@6.4]
  input  [3:0] io_in_432, // @[:@6.4]
  input  [3:0] io_in_433, // @[:@6.4]
  input  [3:0] io_in_434, // @[:@6.4]
  input  [3:0] io_in_435, // @[:@6.4]
  input  [3:0] io_in_436, // @[:@6.4]
  input  [3:0] io_in_437, // @[:@6.4]
  input  [3:0] io_in_438, // @[:@6.4]
  input  [3:0] io_in_439, // @[:@6.4]
  input  [3:0] io_in_440, // @[:@6.4]
  input  [3:0] io_in_441, // @[:@6.4]
  input  [3:0] io_in_442, // @[:@6.4]
  input  [3:0] io_in_443, // @[:@6.4]
  input  [3:0] io_in_444, // @[:@6.4]
  input  [3:0] io_in_445, // @[:@6.4]
  input  [3:0] io_in_446, // @[:@6.4]
  input  [3:0] io_in_447, // @[:@6.4]
  input  [3:0] io_in_448, // @[:@6.4]
  input  [3:0] io_in_449, // @[:@6.4]
  input  [3:0] io_in_450, // @[:@6.4]
  input  [3:0] io_in_451, // @[:@6.4]
  input  [3:0] io_in_452, // @[:@6.4]
  input  [3:0] io_in_453, // @[:@6.4]
  input  [3:0] io_in_454, // @[:@6.4]
  input  [3:0] io_in_455, // @[:@6.4]
  input  [3:0] io_in_456, // @[:@6.4]
  input  [3:0] io_in_457, // @[:@6.4]
  input  [3:0] io_in_458, // @[:@6.4]
  input  [3:0] io_in_459, // @[:@6.4]
  input  [3:0] io_in_460, // @[:@6.4]
  input  [3:0] io_in_461, // @[:@6.4]
  input  [3:0] io_in_462, // @[:@6.4]
  input  [3:0] io_in_463, // @[:@6.4]
  input  [3:0] io_in_464, // @[:@6.4]
  input  [3:0] io_in_465, // @[:@6.4]
  input  [3:0] io_in_466, // @[:@6.4]
  input  [3:0] io_in_467, // @[:@6.4]
  input  [3:0] io_in_468, // @[:@6.4]
  input  [3:0] io_in_469, // @[:@6.4]
  input  [3:0] io_in_470, // @[:@6.4]
  input  [3:0] io_in_471, // @[:@6.4]
  input  [3:0] io_in_472, // @[:@6.4]
  input  [3:0] io_in_473, // @[:@6.4]
  input  [3:0] io_in_474, // @[:@6.4]
  input  [3:0] io_in_475, // @[:@6.4]
  input  [3:0] io_in_476, // @[:@6.4]
  input  [3:0] io_in_477, // @[:@6.4]
  input  [3:0] io_in_478, // @[:@6.4]
  input  [3:0] io_in_479, // @[:@6.4]
  input  [3:0] io_in_480, // @[:@6.4]
  input  [3:0] io_in_481, // @[:@6.4]
  input  [3:0] io_in_482, // @[:@6.4]
  input  [3:0] io_in_483, // @[:@6.4]
  input  [3:0] io_in_484, // @[:@6.4]
  input  [3:0] io_in_485, // @[:@6.4]
  input  [3:0] io_in_486, // @[:@6.4]
  input  [3:0] io_in_487, // @[:@6.4]
  input  [3:0] io_in_488, // @[:@6.4]
  input  [3:0] io_in_489, // @[:@6.4]
  input  [3:0] io_in_490, // @[:@6.4]
  input  [3:0] io_in_491, // @[:@6.4]
  input  [3:0] io_in_492, // @[:@6.4]
  input  [3:0] io_in_493, // @[:@6.4]
  input  [3:0] io_in_494, // @[:@6.4]
  input  [3:0] io_in_495, // @[:@6.4]
  input  [3:0] io_in_496, // @[:@6.4]
  input  [3:0] io_in_497, // @[:@6.4]
  input  [3:0] io_in_498, // @[:@6.4]
  input  [3:0] io_in_499, // @[:@6.4]
  input  [3:0] io_in_500, // @[:@6.4]
  input  [3:0] io_in_501, // @[:@6.4]
  input  [3:0] io_in_502, // @[:@6.4]
  input  [3:0] io_in_503, // @[:@6.4]
  input  [3:0] io_in_504, // @[:@6.4]
  input  [3:0] io_in_505, // @[:@6.4]
  input  [3:0] io_in_506, // @[:@6.4]
  input  [3:0] io_in_507, // @[:@6.4]
  input  [3:0] io_in_508, // @[:@6.4]
  input  [3:0] io_in_509, // @[:@6.4]
  input  [3:0] io_in_510, // @[:@6.4]
  input  [3:0] io_in_511, // @[:@6.4]
  input  [3:0] io_in_512, // @[:@6.4]
  input  [3:0] io_in_513, // @[:@6.4]
  input  [3:0] io_in_514, // @[:@6.4]
  input  [3:0] io_in_515, // @[:@6.4]
  input  [3:0] io_in_516, // @[:@6.4]
  input  [3:0] io_in_517, // @[:@6.4]
  input  [3:0] io_in_518, // @[:@6.4]
  input  [3:0] io_in_519, // @[:@6.4]
  input  [3:0] io_in_520, // @[:@6.4]
  input  [3:0] io_in_521, // @[:@6.4]
  input  [3:0] io_in_522, // @[:@6.4]
  input  [3:0] io_in_523, // @[:@6.4]
  input  [3:0] io_in_524, // @[:@6.4]
  input  [3:0] io_in_525, // @[:@6.4]
  input  [3:0] io_in_526, // @[:@6.4]
  input  [3:0] io_in_527, // @[:@6.4]
  input  [3:0] io_in_528, // @[:@6.4]
  input  [3:0] io_in_529, // @[:@6.4]
  input  [3:0] io_in_530, // @[:@6.4]
  input  [3:0] io_in_531, // @[:@6.4]
  input  [3:0] io_in_532, // @[:@6.4]
  input  [3:0] io_in_533, // @[:@6.4]
  input  [3:0] io_in_534, // @[:@6.4]
  input  [3:0] io_in_535, // @[:@6.4]
  input  [3:0] io_in_536, // @[:@6.4]
  input  [3:0] io_in_537, // @[:@6.4]
  input  [3:0] io_in_538, // @[:@6.4]
  input  [3:0] io_in_539, // @[:@6.4]
  input  [3:0] io_in_540, // @[:@6.4]
  input  [3:0] io_in_541, // @[:@6.4]
  input  [3:0] io_in_542, // @[:@6.4]
  input  [3:0] io_in_543, // @[:@6.4]
  input  [3:0] io_in_544, // @[:@6.4]
  input  [3:0] io_in_545, // @[:@6.4]
  input  [3:0] io_in_546, // @[:@6.4]
  input  [3:0] io_in_547, // @[:@6.4]
  input  [3:0] io_in_548, // @[:@6.4]
  input  [3:0] io_in_549, // @[:@6.4]
  input  [3:0] io_in_550, // @[:@6.4]
  input  [3:0] io_in_551, // @[:@6.4]
  input  [3:0] io_in_552, // @[:@6.4]
  input  [3:0] io_in_553, // @[:@6.4]
  input  [3:0] io_in_554, // @[:@6.4]
  input  [3:0] io_in_555, // @[:@6.4]
  input  [3:0] io_in_556, // @[:@6.4]
  input  [3:0] io_in_557, // @[:@6.4]
  input  [3:0] io_in_558, // @[:@6.4]
  input  [3:0] io_in_559, // @[:@6.4]
  input  [3:0] io_in_560, // @[:@6.4]
  input  [3:0] io_in_561, // @[:@6.4]
  input  [3:0] io_in_562, // @[:@6.4]
  input  [3:0] io_in_563, // @[:@6.4]
  input  [3:0] io_in_564, // @[:@6.4]
  input  [3:0] io_in_565, // @[:@6.4]
  input  [3:0] io_in_566, // @[:@6.4]
  input  [3:0] io_in_567, // @[:@6.4]
  input  [3:0] io_in_568, // @[:@6.4]
  input  [3:0] io_in_569, // @[:@6.4]
  input  [3:0] io_in_570, // @[:@6.4]
  input  [3:0] io_in_571, // @[:@6.4]
  input  [3:0] io_in_572, // @[:@6.4]
  input  [3:0] io_in_573, // @[:@6.4]
  input  [3:0] io_in_574, // @[:@6.4]
  input  [3:0] io_in_575, // @[:@6.4]
  input  [3:0] io_in_576, // @[:@6.4]
  input  [3:0] io_in_577, // @[:@6.4]
  input  [3:0] io_in_578, // @[:@6.4]
  input  [3:0] io_in_579, // @[:@6.4]
  input  [3:0] io_in_580, // @[:@6.4]
  input  [3:0] io_in_581, // @[:@6.4]
  input  [3:0] io_in_582, // @[:@6.4]
  input  [3:0] io_in_583, // @[:@6.4]
  input  [3:0] io_in_584, // @[:@6.4]
  input  [3:0] io_in_585, // @[:@6.4]
  input  [3:0] io_in_586, // @[:@6.4]
  input  [3:0] io_in_587, // @[:@6.4]
  input  [3:0] io_in_588, // @[:@6.4]
  input  [3:0] io_in_589, // @[:@6.4]
  input  [3:0] io_in_590, // @[:@6.4]
  input  [3:0] io_in_591, // @[:@6.4]
  input  [3:0] io_in_592, // @[:@6.4]
  input  [3:0] io_in_593, // @[:@6.4]
  input  [3:0] io_in_594, // @[:@6.4]
  input  [3:0] io_in_595, // @[:@6.4]
  input  [3:0] io_in_596, // @[:@6.4]
  input  [3:0] io_in_597, // @[:@6.4]
  input  [3:0] io_in_598, // @[:@6.4]
  input  [3:0] io_in_599, // @[:@6.4]
  input  [3:0] io_in_600, // @[:@6.4]
  input  [3:0] io_in_601, // @[:@6.4]
  input  [3:0] io_in_602, // @[:@6.4]
  input  [3:0] io_in_603, // @[:@6.4]
  input  [3:0] io_in_604, // @[:@6.4]
  input  [3:0] io_in_605, // @[:@6.4]
  input  [3:0] io_in_606, // @[:@6.4]
  input  [3:0] io_in_607, // @[:@6.4]
  input  [3:0] io_in_608, // @[:@6.4]
  input  [3:0] io_in_609, // @[:@6.4]
  input  [3:0] io_in_610, // @[:@6.4]
  input  [3:0] io_in_611, // @[:@6.4]
  input  [3:0] io_in_612, // @[:@6.4]
  input  [3:0] io_in_613, // @[:@6.4]
  input  [3:0] io_in_614, // @[:@6.4]
  input  [3:0] io_in_615, // @[:@6.4]
  input  [3:0] io_in_616, // @[:@6.4]
  input  [3:0] io_in_617, // @[:@6.4]
  input  [3:0] io_in_618, // @[:@6.4]
  input  [3:0] io_in_619, // @[:@6.4]
  input  [3:0] io_in_620, // @[:@6.4]
  input  [3:0] io_in_621, // @[:@6.4]
  input  [3:0] io_in_622, // @[:@6.4]
  input  [3:0] io_in_623, // @[:@6.4]
  input  [3:0] io_in_624, // @[:@6.4]
  input  [3:0] io_in_625, // @[:@6.4]
  input  [3:0] io_in_626, // @[:@6.4]
  input  [3:0] io_in_627, // @[:@6.4]
  input  [3:0] io_in_628, // @[:@6.4]
  input  [3:0] io_in_629, // @[:@6.4]
  input  [3:0] io_in_630, // @[:@6.4]
  input  [3:0] io_in_631, // @[:@6.4]
  input  [3:0] io_in_632, // @[:@6.4]
  input  [3:0] io_in_633, // @[:@6.4]
  input  [3:0] io_in_634, // @[:@6.4]
  input  [3:0] io_in_635, // @[:@6.4]
  input  [3:0] io_in_636, // @[:@6.4]
  input  [3:0] io_in_637, // @[:@6.4]
  input  [3:0] io_in_638, // @[:@6.4]
  input  [3:0] io_in_639, // @[:@6.4]
  input  [3:0] io_in_640, // @[:@6.4]
  input  [3:0] io_in_641, // @[:@6.4]
  input  [3:0] io_in_642, // @[:@6.4]
  input  [3:0] io_in_643, // @[:@6.4]
  input  [3:0] io_in_644, // @[:@6.4]
  input  [3:0] io_in_645, // @[:@6.4]
  input  [3:0] io_in_646, // @[:@6.4]
  input  [3:0] io_in_647, // @[:@6.4]
  input  [3:0] io_in_648, // @[:@6.4]
  input  [3:0] io_in_649, // @[:@6.4]
  input  [3:0] io_in_650, // @[:@6.4]
  input  [3:0] io_in_651, // @[:@6.4]
  input  [3:0] io_in_652, // @[:@6.4]
  input  [3:0] io_in_653, // @[:@6.4]
  input  [3:0] io_in_654, // @[:@6.4]
  input  [3:0] io_in_655, // @[:@6.4]
  input  [3:0] io_in_656, // @[:@6.4]
  input  [3:0] io_in_657, // @[:@6.4]
  input  [3:0] io_in_658, // @[:@6.4]
  input  [3:0] io_in_659, // @[:@6.4]
  input  [3:0] io_in_660, // @[:@6.4]
  input  [3:0] io_in_661, // @[:@6.4]
  input  [3:0] io_in_662, // @[:@6.4]
  input  [3:0] io_in_663, // @[:@6.4]
  input  [3:0] io_in_664, // @[:@6.4]
  input  [3:0] io_in_665, // @[:@6.4]
  input  [3:0] io_in_666, // @[:@6.4]
  input  [3:0] io_in_667, // @[:@6.4]
  input  [3:0] io_in_668, // @[:@6.4]
  input  [3:0] io_in_669, // @[:@6.4]
  input  [3:0] io_in_670, // @[:@6.4]
  input  [3:0] io_in_671, // @[:@6.4]
  input  [3:0] io_in_672, // @[:@6.4]
  input  [3:0] io_in_673, // @[:@6.4]
  input  [3:0] io_in_674, // @[:@6.4]
  input  [3:0] io_in_675, // @[:@6.4]
  input  [3:0] io_in_676, // @[:@6.4]
  input  [3:0] io_in_677, // @[:@6.4]
  input  [3:0] io_in_678, // @[:@6.4]
  input  [3:0] io_in_679, // @[:@6.4]
  input  [3:0] io_in_680, // @[:@6.4]
  input  [3:0] io_in_681, // @[:@6.4]
  input  [3:0] io_in_682, // @[:@6.4]
  input  [3:0] io_in_683, // @[:@6.4]
  input  [3:0] io_in_684, // @[:@6.4]
  input  [3:0] io_in_685, // @[:@6.4]
  input  [3:0] io_in_686, // @[:@6.4]
  input  [3:0] io_in_687, // @[:@6.4]
  input  [3:0] io_in_688, // @[:@6.4]
  input  [3:0] io_in_689, // @[:@6.4]
  input  [3:0] io_in_690, // @[:@6.4]
  input  [3:0] io_in_691, // @[:@6.4]
  input  [3:0] io_in_692, // @[:@6.4]
  input  [3:0] io_in_693, // @[:@6.4]
  input  [3:0] io_in_694, // @[:@6.4]
  input  [3:0] io_in_695, // @[:@6.4]
  input  [3:0] io_in_696, // @[:@6.4]
  input  [3:0] io_in_697, // @[:@6.4]
  input  [3:0] io_in_698, // @[:@6.4]
  input  [3:0] io_in_699, // @[:@6.4]
  input  [3:0] io_in_700, // @[:@6.4]
  input  [3:0] io_in_701, // @[:@6.4]
  input  [3:0] io_in_702, // @[:@6.4]
  input  [3:0] io_in_703, // @[:@6.4]
  input  [3:0] io_in_704, // @[:@6.4]
  input  [3:0] io_in_705, // @[:@6.4]
  input  [3:0] io_in_706, // @[:@6.4]
  input  [3:0] io_in_707, // @[:@6.4]
  input  [3:0] io_in_708, // @[:@6.4]
  input  [3:0] io_in_709, // @[:@6.4]
  input  [3:0] io_in_710, // @[:@6.4]
  input  [3:0] io_in_711, // @[:@6.4]
  input  [3:0] io_in_712, // @[:@6.4]
  input  [3:0] io_in_713, // @[:@6.4]
  input  [3:0] io_in_714, // @[:@6.4]
  input  [3:0] io_in_715, // @[:@6.4]
  input  [3:0] io_in_716, // @[:@6.4]
  input  [3:0] io_in_717, // @[:@6.4]
  input  [3:0] io_in_718, // @[:@6.4]
  input  [3:0] io_in_719, // @[:@6.4]
  input  [3:0] io_in_720, // @[:@6.4]
  input  [3:0] io_in_721, // @[:@6.4]
  input  [3:0] io_in_722, // @[:@6.4]
  input  [3:0] io_in_723, // @[:@6.4]
  input  [3:0] io_in_724, // @[:@6.4]
  input  [3:0] io_in_725, // @[:@6.4]
  input  [3:0] io_in_726, // @[:@6.4]
  input  [3:0] io_in_727, // @[:@6.4]
  input  [3:0] io_in_728, // @[:@6.4]
  input  [3:0] io_in_729, // @[:@6.4]
  input  [3:0] io_in_730, // @[:@6.4]
  input  [3:0] io_in_731, // @[:@6.4]
  input  [3:0] io_in_732, // @[:@6.4]
  input  [3:0] io_in_733, // @[:@6.4]
  input  [3:0] io_in_734, // @[:@6.4]
  input  [3:0] io_in_735, // @[:@6.4]
  input  [3:0] io_in_736, // @[:@6.4]
  input  [3:0] io_in_737, // @[:@6.4]
  input  [3:0] io_in_738, // @[:@6.4]
  input  [3:0] io_in_739, // @[:@6.4]
  input  [3:0] io_in_740, // @[:@6.4]
  input  [3:0] io_in_741, // @[:@6.4]
  input  [3:0] io_in_742, // @[:@6.4]
  input  [3:0] io_in_743, // @[:@6.4]
  input  [3:0] io_in_744, // @[:@6.4]
  input  [3:0] io_in_745, // @[:@6.4]
  input  [3:0] io_in_746, // @[:@6.4]
  input  [3:0] io_in_747, // @[:@6.4]
  input  [3:0] io_in_748, // @[:@6.4]
  input  [3:0] io_in_749, // @[:@6.4]
  input  [3:0] io_in_750, // @[:@6.4]
  input  [3:0] io_in_751, // @[:@6.4]
  input  [3:0] io_in_752, // @[:@6.4]
  input  [3:0] io_in_753, // @[:@6.4]
  input  [3:0] io_in_754, // @[:@6.4]
  input  [3:0] io_in_755, // @[:@6.4]
  input  [3:0] io_in_756, // @[:@6.4]
  input  [3:0] io_in_757, // @[:@6.4]
  input  [3:0] io_in_758, // @[:@6.4]
  input  [3:0] io_in_759, // @[:@6.4]
  input  [3:0] io_in_760, // @[:@6.4]
  input  [3:0] io_in_761, // @[:@6.4]
  input  [3:0] io_in_762, // @[:@6.4]
  input  [3:0] io_in_763, // @[:@6.4]
  input  [3:0] io_in_764, // @[:@6.4]
  input  [3:0] io_in_765, // @[:@6.4]
  input  [3:0] io_in_766, // @[:@6.4]
  input  [3:0] io_in_767, // @[:@6.4]
  input  [3:0] io_in_768, // @[:@6.4]
  input  [3:0] io_in_769, // @[:@6.4]
  input  [3:0] io_in_770, // @[:@6.4]
  input  [3:0] io_in_771, // @[:@6.4]
  input  [3:0] io_in_772, // @[:@6.4]
  input  [3:0] io_in_773, // @[:@6.4]
  input  [3:0] io_in_774, // @[:@6.4]
  input  [3:0] io_in_775, // @[:@6.4]
  input  [3:0] io_in_776, // @[:@6.4]
  input  [3:0] io_in_777, // @[:@6.4]
  input  [3:0] io_in_778, // @[:@6.4]
  input  [3:0] io_in_779, // @[:@6.4]
  input  [3:0] io_in_780, // @[:@6.4]
  input  [3:0] io_in_781, // @[:@6.4]
  input  [3:0] io_in_782, // @[:@6.4]
  input  [3:0] io_in_783, // @[:@6.4]
  output [3:0] io_out_0, // @[:@6.4]
  output [3:0] io_out_1, // @[:@6.4]
  output [3:0] io_out_2, // @[:@6.4]
  output [3:0] io_out_3, // @[:@6.4]
  output [3:0] io_out_4, // @[:@6.4]
  output [3:0] io_out_5, // @[:@6.4]
  output [3:0] io_out_6, // @[:@6.4]
  output [3:0] io_out_7, // @[:@6.4]
  output [3:0] io_out_8, // @[:@6.4]
  output [3:0] io_out_9, // @[:@6.4]
  output [3:0] io_out_10, // @[:@6.4]
  output [3:0] io_out_11, // @[:@6.4]
  output [3:0] io_out_12, // @[:@6.4]
  output [3:0] io_out_13, // @[:@6.4]
  output [3:0] io_out_14, // @[:@6.4]
  output [3:0] io_out_15, // @[:@6.4]
  output [3:0] io_out_16, // @[:@6.4]
  output [3:0] io_out_17, // @[:@6.4]
  output [3:0] io_out_18, // @[:@6.4]
  output [3:0] io_out_19, // @[:@6.4]
  output [3:0] io_out_20, // @[:@6.4]
  output [3:0] io_out_21, // @[:@6.4]
  output [3:0] io_out_22, // @[:@6.4]
  output [3:0] io_out_23, // @[:@6.4]
  output [3:0] io_out_24, // @[:@6.4]
  output [3:0] io_out_25, // @[:@6.4]
  output [3:0] io_out_26, // @[:@6.4]
  output [3:0] io_out_27, // @[:@6.4]
  output [3:0] io_out_28, // @[:@6.4]
  output [3:0] io_out_29, // @[:@6.4]
  output [3:0] io_out_30, // @[:@6.4]
  output [3:0] io_out_31, // @[:@6.4]
  output [3:0] io_out_32, // @[:@6.4]
  output [3:0] io_out_33, // @[:@6.4]
  output [3:0] io_out_34, // @[:@6.4]
  output [3:0] io_out_35, // @[:@6.4]
  output [3:0] io_out_36, // @[:@6.4]
  output [3:0] io_out_37, // @[:@6.4]
  output [3:0] io_out_38, // @[:@6.4]
  output [3:0] io_out_39, // @[:@6.4]
  output [3:0] io_out_40, // @[:@6.4]
  output [3:0] io_out_41, // @[:@6.4]
  output [3:0] io_out_42, // @[:@6.4]
  output [3:0] io_out_43, // @[:@6.4]
  output [3:0] io_out_44, // @[:@6.4]
  output [3:0] io_out_45, // @[:@6.4]
  output [3:0] io_out_46, // @[:@6.4]
  output [3:0] io_out_47, // @[:@6.4]
  output [3:0] io_out_48, // @[:@6.4]
  output [3:0] io_out_49, // @[:@6.4]
  output [3:0] io_out_50, // @[:@6.4]
  output [3:0] io_out_51, // @[:@6.4]
  output [3:0] io_out_52, // @[:@6.4]
  output [3:0] io_out_53, // @[:@6.4]
  output [3:0] io_out_54, // @[:@6.4]
  output [3:0] io_out_55, // @[:@6.4]
  output [3:0] io_out_56, // @[:@6.4]
  output [3:0] io_out_57, // @[:@6.4]
  output [3:0] io_out_58, // @[:@6.4]
  output [3:0] io_out_59, // @[:@6.4]
  output [3:0] io_out_60, // @[:@6.4]
  output [3:0] io_out_61, // @[:@6.4]
  output [3:0] io_out_62, // @[:@6.4]
  output [3:0] io_out_63, // @[:@6.4]
  output [3:0] io_out_64, // @[:@6.4]
  output [3:0] io_out_65, // @[:@6.4]
  output [3:0] io_out_66, // @[:@6.4]
  output [3:0] io_out_67, // @[:@6.4]
  output [3:0] io_out_68, // @[:@6.4]
  output [3:0] io_out_69, // @[:@6.4]
  output [3:0] io_out_70, // @[:@6.4]
  output [3:0] io_out_71, // @[:@6.4]
  output [3:0] io_out_72, // @[:@6.4]
  output [3:0] io_out_73, // @[:@6.4]
  output [3:0] io_out_74, // @[:@6.4]
  output [3:0] io_out_75, // @[:@6.4]
  output [3:0] io_out_76, // @[:@6.4]
  output [3:0] io_out_77, // @[:@6.4]
  output [3:0] io_out_78, // @[:@6.4]
  output [3:0] io_out_79, // @[:@6.4]
  output [3:0] io_out_80, // @[:@6.4]
  output [3:0] io_out_81, // @[:@6.4]
  output [3:0] io_out_82, // @[:@6.4]
  output [3:0] io_out_83, // @[:@6.4]
  output [3:0] io_out_84, // @[:@6.4]
  output [3:0] io_out_85, // @[:@6.4]
  output [3:0] io_out_86, // @[:@6.4]
  output [3:0] io_out_87, // @[:@6.4]
  output [3:0] io_out_88, // @[:@6.4]
  output [3:0] io_out_89, // @[:@6.4]
  output [3:0] io_out_90, // @[:@6.4]
  output [3:0] io_out_91, // @[:@6.4]
  output [3:0] io_out_92, // @[:@6.4]
  output [3:0] io_out_93, // @[:@6.4]
  output [3:0] io_out_94, // @[:@6.4]
  output [3:0] io_out_95, // @[:@6.4]
  output [3:0] io_out_96, // @[:@6.4]
  output [3:0] io_out_97, // @[:@6.4]
  output [3:0] io_out_98, // @[:@6.4]
  output [3:0] io_out_99, // @[:@6.4]
  output [3:0] io_out_100, // @[:@6.4]
  output [3:0] io_out_101, // @[:@6.4]
  output [3:0] io_out_102, // @[:@6.4]
  output [3:0] io_out_103, // @[:@6.4]
  output [3:0] io_out_104, // @[:@6.4]
  output [3:0] io_out_105, // @[:@6.4]
  output [3:0] io_out_106, // @[:@6.4]
  output [3:0] io_out_107, // @[:@6.4]
  output [3:0] io_out_108, // @[:@6.4]
  output [3:0] io_out_109, // @[:@6.4]
  output [3:0] io_out_110, // @[:@6.4]
  output [3:0] io_out_111, // @[:@6.4]
  output [3:0] io_out_112, // @[:@6.4]
  output [3:0] io_out_113, // @[:@6.4]
  output [3:0] io_out_114, // @[:@6.4]
  output [3:0] io_out_115, // @[:@6.4]
  output [3:0] io_out_116, // @[:@6.4]
  output [3:0] io_out_117, // @[:@6.4]
  output [3:0] io_out_118, // @[:@6.4]
  output [3:0] io_out_119, // @[:@6.4]
  output [3:0] io_out_120, // @[:@6.4]
  output [3:0] io_out_121, // @[:@6.4]
  output [3:0] io_out_122, // @[:@6.4]
  output [3:0] io_out_123, // @[:@6.4]
  output [3:0] io_out_124, // @[:@6.4]
  output [3:0] io_out_125, // @[:@6.4]
  output [3:0] io_out_126, // @[:@6.4]
  output [3:0] io_out_127, // @[:@6.4]
  output [3:0] io_out_128, // @[:@6.4]
  output [3:0] io_out_129, // @[:@6.4]
  output [3:0] io_out_130, // @[:@6.4]
  output [3:0] io_out_131, // @[:@6.4]
  output [3:0] io_out_132, // @[:@6.4]
  output [3:0] io_out_133, // @[:@6.4]
  output [3:0] io_out_134, // @[:@6.4]
  output [3:0] io_out_135, // @[:@6.4]
  output [3:0] io_out_136, // @[:@6.4]
  output [3:0] io_out_137, // @[:@6.4]
  output [3:0] io_out_138, // @[:@6.4]
  output [3:0] io_out_139, // @[:@6.4]
  output [3:0] io_out_140, // @[:@6.4]
  output [3:0] io_out_141, // @[:@6.4]
  output [3:0] io_out_142, // @[:@6.4]
  output [3:0] io_out_143, // @[:@6.4]
  output [3:0] io_out_144, // @[:@6.4]
  output [3:0] io_out_145, // @[:@6.4]
  output [3:0] io_out_146, // @[:@6.4]
  output [3:0] io_out_147, // @[:@6.4]
  output [3:0] io_out_148, // @[:@6.4]
  output [3:0] io_out_149, // @[:@6.4]
  output [3:0] io_out_150, // @[:@6.4]
  output [3:0] io_out_151, // @[:@6.4]
  output [3:0] io_out_152, // @[:@6.4]
  output [3:0] io_out_153, // @[:@6.4]
  output [3:0] io_out_154, // @[:@6.4]
  output [3:0] io_out_155, // @[:@6.4]
  output [3:0] io_out_156, // @[:@6.4]
  output [3:0] io_out_157, // @[:@6.4]
  output [3:0] io_out_158, // @[:@6.4]
  output [3:0] io_out_159, // @[:@6.4]
  output [3:0] io_out_160, // @[:@6.4]
  output [3:0] io_out_161, // @[:@6.4]
  output [3:0] io_out_162, // @[:@6.4]
  output [3:0] io_out_163, // @[:@6.4]
  output [3:0] io_out_164, // @[:@6.4]
  output [3:0] io_out_165, // @[:@6.4]
  output [3:0] io_out_166, // @[:@6.4]
  output [3:0] io_out_167, // @[:@6.4]
  output [3:0] io_out_168, // @[:@6.4]
  output [3:0] io_out_169, // @[:@6.4]
  output [3:0] io_out_170, // @[:@6.4]
  output [3:0] io_out_171, // @[:@6.4]
  output [3:0] io_out_172, // @[:@6.4]
  output [3:0] io_out_173, // @[:@6.4]
  output [3:0] io_out_174, // @[:@6.4]
  output [3:0] io_out_175, // @[:@6.4]
  output [3:0] io_out_176, // @[:@6.4]
  output [3:0] io_out_177, // @[:@6.4]
  output [3:0] io_out_178, // @[:@6.4]
  output [3:0] io_out_179, // @[:@6.4]
  output [3:0] io_out_180, // @[:@6.4]
  output [3:0] io_out_181, // @[:@6.4]
  output [3:0] io_out_182, // @[:@6.4]
  output [3:0] io_out_183, // @[:@6.4]
  output [3:0] io_out_184, // @[:@6.4]
  output [3:0] io_out_185, // @[:@6.4]
  output [3:0] io_out_186, // @[:@6.4]
  output [3:0] io_out_187, // @[:@6.4]
  output [3:0] io_out_188, // @[:@6.4]
  output [3:0] io_out_189, // @[:@6.4]
  output [3:0] io_out_190, // @[:@6.4]
  output [3:0] io_out_191, // @[:@6.4]
  output [3:0] io_out_192, // @[:@6.4]
  output [3:0] io_out_193, // @[:@6.4]
  output [3:0] io_out_194, // @[:@6.4]
  output [3:0] io_out_195, // @[:@6.4]
  output [3:0] io_out_196, // @[:@6.4]
  output [3:0] io_out_197, // @[:@6.4]
  output [3:0] io_out_198, // @[:@6.4]
  output [3:0] io_out_199, // @[:@6.4]
  output [3:0] io_out_200, // @[:@6.4]
  output [3:0] io_out_201, // @[:@6.4]
  output [3:0] io_out_202, // @[:@6.4]
  output [3:0] io_out_203, // @[:@6.4]
  output [3:0] io_out_204, // @[:@6.4]
  output [3:0] io_out_205, // @[:@6.4]
  output [3:0] io_out_206, // @[:@6.4]
  output [3:0] io_out_207, // @[:@6.4]
  output [3:0] io_out_208, // @[:@6.4]
  output [3:0] io_out_209, // @[:@6.4]
  output [3:0] io_out_210, // @[:@6.4]
  output [3:0] io_out_211, // @[:@6.4]
  output [3:0] io_out_212, // @[:@6.4]
  output [3:0] io_out_213, // @[:@6.4]
  output [3:0] io_out_214, // @[:@6.4]
  output [3:0] io_out_215, // @[:@6.4]
  output [3:0] io_out_216, // @[:@6.4]
  output [3:0] io_out_217, // @[:@6.4]
  output [3:0] io_out_218, // @[:@6.4]
  output [3:0] io_out_219, // @[:@6.4]
  output [3:0] io_out_220, // @[:@6.4]
  output [3:0] io_out_221, // @[:@6.4]
  output [3:0] io_out_222, // @[:@6.4]
  output [3:0] io_out_223, // @[:@6.4]
  output [3:0] io_out_224, // @[:@6.4]
  output [3:0] io_out_225, // @[:@6.4]
  output [3:0] io_out_226, // @[:@6.4]
  output [3:0] io_out_227, // @[:@6.4]
  output [3:0] io_out_228, // @[:@6.4]
  output [3:0] io_out_229, // @[:@6.4]
  output [3:0] io_out_230, // @[:@6.4]
  output [3:0] io_out_231, // @[:@6.4]
  output [3:0] io_out_232, // @[:@6.4]
  output [3:0] io_out_233, // @[:@6.4]
  output [3:0] io_out_234, // @[:@6.4]
  output [3:0] io_out_235, // @[:@6.4]
  output [3:0] io_out_236, // @[:@6.4]
  output [3:0] io_out_237, // @[:@6.4]
  output [3:0] io_out_238, // @[:@6.4]
  output [3:0] io_out_239, // @[:@6.4]
  output [3:0] io_out_240, // @[:@6.4]
  output [3:0] io_out_241, // @[:@6.4]
  output [3:0] io_out_242, // @[:@6.4]
  output [3:0] io_out_243, // @[:@6.4]
  output [3:0] io_out_244, // @[:@6.4]
  output [3:0] io_out_245, // @[:@6.4]
  output [3:0] io_out_246, // @[:@6.4]
  output [3:0] io_out_247, // @[:@6.4]
  output [3:0] io_out_248, // @[:@6.4]
  output [3:0] io_out_249, // @[:@6.4]
  output [3:0] io_out_250, // @[:@6.4]
  output [3:0] io_out_251, // @[:@6.4]
  output [3:0] io_out_252, // @[:@6.4]
  output [3:0] io_out_253, // @[:@6.4]
  output [3:0] io_out_254, // @[:@6.4]
  output [3:0] io_out_255, // @[:@6.4]
  output [3:0] io_out_256, // @[:@6.4]
  output [3:0] io_out_257, // @[:@6.4]
  output [3:0] io_out_258, // @[:@6.4]
  output [3:0] io_out_259, // @[:@6.4]
  output [3:0] io_out_260, // @[:@6.4]
  output [3:0] io_out_261, // @[:@6.4]
  output [3:0] io_out_262, // @[:@6.4]
  output [3:0] io_out_263, // @[:@6.4]
  output [3:0] io_out_264, // @[:@6.4]
  output [3:0] io_out_265, // @[:@6.4]
  output [3:0] io_out_266, // @[:@6.4]
  output [3:0] io_out_267, // @[:@6.4]
  output [3:0] io_out_268, // @[:@6.4]
  output [3:0] io_out_269, // @[:@6.4]
  output [3:0] io_out_270, // @[:@6.4]
  output [3:0] io_out_271, // @[:@6.4]
  output [3:0] io_out_272, // @[:@6.4]
  output [3:0] io_out_273, // @[:@6.4]
  output [3:0] io_out_274, // @[:@6.4]
  output [3:0] io_out_275, // @[:@6.4]
  output [3:0] io_out_276, // @[:@6.4]
  output [3:0] io_out_277, // @[:@6.4]
  output [3:0] io_out_278, // @[:@6.4]
  output [3:0] io_out_279, // @[:@6.4]
  output [3:0] io_out_280, // @[:@6.4]
  output [3:0] io_out_281, // @[:@6.4]
  output [3:0] io_out_282, // @[:@6.4]
  output [3:0] io_out_283, // @[:@6.4]
  output [3:0] io_out_284, // @[:@6.4]
  output [3:0] io_out_285, // @[:@6.4]
  output [3:0] io_out_286, // @[:@6.4]
  output [3:0] io_out_287, // @[:@6.4]
  output [3:0] io_out_288, // @[:@6.4]
  output [3:0] io_out_289, // @[:@6.4]
  output [3:0] io_out_290, // @[:@6.4]
  output [3:0] io_out_291, // @[:@6.4]
  output [3:0] io_out_292, // @[:@6.4]
  output [3:0] io_out_293, // @[:@6.4]
  output [3:0] io_out_294, // @[:@6.4]
  output [3:0] io_out_295, // @[:@6.4]
  output [3:0] io_out_296, // @[:@6.4]
  output [3:0] io_out_297, // @[:@6.4]
  output [3:0] io_out_298, // @[:@6.4]
  output [3:0] io_out_299, // @[:@6.4]
  output [3:0] io_out_300, // @[:@6.4]
  output [3:0] io_out_301, // @[:@6.4]
  output [3:0] io_out_302, // @[:@6.4]
  output [3:0] io_out_303, // @[:@6.4]
  output [3:0] io_out_304, // @[:@6.4]
  output [3:0] io_out_305, // @[:@6.4]
  output [3:0] io_out_306, // @[:@6.4]
  output [3:0] io_out_307, // @[:@6.4]
  output [3:0] io_out_308, // @[:@6.4]
  output [3:0] io_out_309, // @[:@6.4]
  output [3:0] io_out_310, // @[:@6.4]
  output [3:0] io_out_311, // @[:@6.4]
  output [3:0] io_out_312, // @[:@6.4]
  output [3:0] io_out_313, // @[:@6.4]
  output [3:0] io_out_314, // @[:@6.4]
  output [3:0] io_out_315, // @[:@6.4]
  output [3:0] io_out_316, // @[:@6.4]
  output [3:0] io_out_317, // @[:@6.4]
  output [3:0] io_out_318, // @[:@6.4]
  output [3:0] io_out_319, // @[:@6.4]
  output [3:0] io_out_320, // @[:@6.4]
  output [3:0] io_out_321, // @[:@6.4]
  output [3:0] io_out_322, // @[:@6.4]
  output [3:0] io_out_323, // @[:@6.4]
  output [3:0] io_out_324, // @[:@6.4]
  output [3:0] io_out_325, // @[:@6.4]
  output [3:0] io_out_326, // @[:@6.4]
  output [3:0] io_out_327, // @[:@6.4]
  output [3:0] io_out_328, // @[:@6.4]
  output [3:0] io_out_329, // @[:@6.4]
  output [3:0] io_out_330, // @[:@6.4]
  output [3:0] io_out_331, // @[:@6.4]
  output [3:0] io_out_332, // @[:@6.4]
  output [3:0] io_out_333, // @[:@6.4]
  output [3:0] io_out_334, // @[:@6.4]
  output [3:0] io_out_335, // @[:@6.4]
  output [3:0] io_out_336, // @[:@6.4]
  output [3:0] io_out_337, // @[:@6.4]
  output [3:0] io_out_338, // @[:@6.4]
  output [3:0] io_out_339, // @[:@6.4]
  output [3:0] io_out_340, // @[:@6.4]
  output [3:0] io_out_341, // @[:@6.4]
  output [3:0] io_out_342, // @[:@6.4]
  output [3:0] io_out_343, // @[:@6.4]
  output [3:0] io_out_344, // @[:@6.4]
  output [3:0] io_out_345, // @[:@6.4]
  output [3:0] io_out_346, // @[:@6.4]
  output [3:0] io_out_347, // @[:@6.4]
  output [3:0] io_out_348, // @[:@6.4]
  output [3:0] io_out_349, // @[:@6.4]
  output [3:0] io_out_350, // @[:@6.4]
  output [3:0] io_out_351, // @[:@6.4]
  output [3:0] io_out_352, // @[:@6.4]
  output [3:0] io_out_353, // @[:@6.4]
  output [3:0] io_out_354, // @[:@6.4]
  output [3:0] io_out_355, // @[:@6.4]
  output [3:0] io_out_356, // @[:@6.4]
  output [3:0] io_out_357, // @[:@6.4]
  output [3:0] io_out_358, // @[:@6.4]
  output [3:0] io_out_359, // @[:@6.4]
  output [3:0] io_out_360, // @[:@6.4]
  output [3:0] io_out_361, // @[:@6.4]
  output [3:0] io_out_362, // @[:@6.4]
  output [3:0] io_out_363, // @[:@6.4]
  output [3:0] io_out_364, // @[:@6.4]
  output [3:0] io_out_365, // @[:@6.4]
  output [3:0] io_out_366, // @[:@6.4]
  output [3:0] io_out_367, // @[:@6.4]
  output [3:0] io_out_368, // @[:@6.4]
  output [3:0] io_out_369, // @[:@6.4]
  output [3:0] io_out_370, // @[:@6.4]
  output [3:0] io_out_371, // @[:@6.4]
  output [3:0] io_out_372, // @[:@6.4]
  output [3:0] io_out_373, // @[:@6.4]
  output [3:0] io_out_374, // @[:@6.4]
  output [3:0] io_out_375, // @[:@6.4]
  output [3:0] io_out_376, // @[:@6.4]
  output [3:0] io_out_377, // @[:@6.4]
  output [3:0] io_out_378, // @[:@6.4]
  output [3:0] io_out_379, // @[:@6.4]
  output [3:0] io_out_380, // @[:@6.4]
  output [3:0] io_out_381, // @[:@6.4]
  output [3:0] io_out_382, // @[:@6.4]
  output [3:0] io_out_383, // @[:@6.4]
  output [3:0] io_out_384, // @[:@6.4]
  output [3:0] io_out_385, // @[:@6.4]
  output [3:0] io_out_386, // @[:@6.4]
  output [3:0] io_out_387, // @[:@6.4]
  output [3:0] io_out_388, // @[:@6.4]
  output [3:0] io_out_389, // @[:@6.4]
  output [3:0] io_out_390, // @[:@6.4]
  output [3:0] io_out_391, // @[:@6.4]
  output [3:0] io_out_392, // @[:@6.4]
  output [3:0] io_out_393, // @[:@6.4]
  output [3:0] io_out_394, // @[:@6.4]
  output [3:0] io_out_395, // @[:@6.4]
  output [3:0] io_out_396, // @[:@6.4]
  output [3:0] io_out_397, // @[:@6.4]
  output [3:0] io_out_398, // @[:@6.4]
  output [3:0] io_out_399, // @[:@6.4]
  output [3:0] io_out_400, // @[:@6.4]
  output [3:0] io_out_401, // @[:@6.4]
  output [3:0] io_out_402, // @[:@6.4]
  output [3:0] io_out_403, // @[:@6.4]
  output [3:0] io_out_404, // @[:@6.4]
  output [3:0] io_out_405, // @[:@6.4]
  output [3:0] io_out_406, // @[:@6.4]
  output [3:0] io_out_407, // @[:@6.4]
  output [3:0] io_out_408, // @[:@6.4]
  output [3:0] io_out_409, // @[:@6.4]
  output [3:0] io_out_410, // @[:@6.4]
  output [3:0] io_out_411, // @[:@6.4]
  output [3:0] io_out_412, // @[:@6.4]
  output [3:0] io_out_413, // @[:@6.4]
  output [3:0] io_out_414, // @[:@6.4]
  output [3:0] io_out_415, // @[:@6.4]
  output [3:0] io_out_416, // @[:@6.4]
  output [3:0] io_out_417, // @[:@6.4]
  output [3:0] io_out_418, // @[:@6.4]
  output [3:0] io_out_419, // @[:@6.4]
  output [3:0] io_out_420, // @[:@6.4]
  output [3:0] io_out_421, // @[:@6.4]
  output [3:0] io_out_422, // @[:@6.4]
  output [3:0] io_out_423, // @[:@6.4]
  output [3:0] io_out_424, // @[:@6.4]
  output [3:0] io_out_425, // @[:@6.4]
  output [3:0] io_out_426, // @[:@6.4]
  output [3:0] io_out_427, // @[:@6.4]
  output [3:0] io_out_428, // @[:@6.4]
  output [3:0] io_out_429, // @[:@6.4]
  output [3:0] io_out_430, // @[:@6.4]
  output [3:0] io_out_431, // @[:@6.4]
  output [3:0] io_out_432, // @[:@6.4]
  output [3:0] io_out_433, // @[:@6.4]
  output [3:0] io_out_434, // @[:@6.4]
  output [3:0] io_out_435, // @[:@6.4]
  output [3:0] io_out_436, // @[:@6.4]
  output [3:0] io_out_437, // @[:@6.4]
  output [3:0] io_out_438, // @[:@6.4]
  output [3:0] io_out_439, // @[:@6.4]
  output [3:0] io_out_440, // @[:@6.4]
  output [3:0] io_out_441, // @[:@6.4]
  output [3:0] io_out_442, // @[:@6.4]
  output [3:0] io_out_443, // @[:@6.4]
  output [3:0] io_out_444, // @[:@6.4]
  output [3:0] io_out_445, // @[:@6.4]
  output [3:0] io_out_446, // @[:@6.4]
  output [3:0] io_out_447, // @[:@6.4]
  output [3:0] io_out_448, // @[:@6.4]
  output [3:0] io_out_449, // @[:@6.4]
  output [3:0] io_out_450, // @[:@6.4]
  output [3:0] io_out_451, // @[:@6.4]
  output [3:0] io_out_452, // @[:@6.4]
  output [3:0] io_out_453, // @[:@6.4]
  output [3:0] io_out_454, // @[:@6.4]
  output [3:0] io_out_455, // @[:@6.4]
  output [3:0] io_out_456, // @[:@6.4]
  output [3:0] io_out_457, // @[:@6.4]
  output [3:0] io_out_458, // @[:@6.4]
  output [3:0] io_out_459, // @[:@6.4]
  output [3:0] io_out_460, // @[:@6.4]
  output [3:0] io_out_461, // @[:@6.4]
  output [3:0] io_out_462, // @[:@6.4]
  output [3:0] io_out_463, // @[:@6.4]
  output [3:0] io_out_464, // @[:@6.4]
  output [3:0] io_out_465, // @[:@6.4]
  output [3:0] io_out_466, // @[:@6.4]
  output [3:0] io_out_467, // @[:@6.4]
  output [3:0] io_out_468, // @[:@6.4]
  output [3:0] io_out_469, // @[:@6.4]
  output [3:0] io_out_470, // @[:@6.4]
  output [3:0] io_out_471, // @[:@6.4]
  output [3:0] io_out_472, // @[:@6.4]
  output [3:0] io_out_473, // @[:@6.4]
  output [3:0] io_out_474, // @[:@6.4]
  output [3:0] io_out_475, // @[:@6.4]
  output [3:0] io_out_476, // @[:@6.4]
  output [3:0] io_out_477, // @[:@6.4]
  output [3:0] io_out_478, // @[:@6.4]
  output [3:0] io_out_479, // @[:@6.4]
  output [3:0] io_out_480, // @[:@6.4]
  output [3:0] io_out_481, // @[:@6.4]
  output [3:0] io_out_482, // @[:@6.4]
  output [3:0] io_out_483, // @[:@6.4]
  output [3:0] io_out_484, // @[:@6.4]
  output [3:0] io_out_485, // @[:@6.4]
  output [3:0] io_out_486, // @[:@6.4]
  output [3:0] io_out_487, // @[:@6.4]
  output [3:0] io_out_488, // @[:@6.4]
  output [3:0] io_out_489, // @[:@6.4]
  output [3:0] io_out_490, // @[:@6.4]
  output [3:0] io_out_491, // @[:@6.4]
  output [3:0] io_out_492, // @[:@6.4]
  output [3:0] io_out_493, // @[:@6.4]
  output [3:0] io_out_494, // @[:@6.4]
  output [3:0] io_out_495, // @[:@6.4]
  output [3:0] io_out_496, // @[:@6.4]
  output [3:0] io_out_497, // @[:@6.4]
  output [3:0] io_out_498, // @[:@6.4]
  output [3:0] io_out_499, // @[:@6.4]
  output [3:0] io_out_500, // @[:@6.4]
  output [3:0] io_out_501, // @[:@6.4]
  output [3:0] io_out_502, // @[:@6.4]
  output [3:0] io_out_503, // @[:@6.4]
  output [3:0] io_out_504, // @[:@6.4]
  output [3:0] io_out_505, // @[:@6.4]
  output [3:0] io_out_506, // @[:@6.4]
  output [3:0] io_out_507, // @[:@6.4]
  output [3:0] io_out_508, // @[:@6.4]
  output [3:0] io_out_509, // @[:@6.4]
  output [3:0] io_out_510, // @[:@6.4]
  output [3:0] io_out_511, // @[:@6.4]
  output [3:0] io_out_512, // @[:@6.4]
  output [3:0] io_out_513, // @[:@6.4]
  output [3:0] io_out_514, // @[:@6.4]
  output [3:0] io_out_515, // @[:@6.4]
  output [3:0] io_out_516, // @[:@6.4]
  output [3:0] io_out_517, // @[:@6.4]
  output [3:0] io_out_518, // @[:@6.4]
  output [3:0] io_out_519, // @[:@6.4]
  output [3:0] io_out_520, // @[:@6.4]
  output [3:0] io_out_521, // @[:@6.4]
  output [3:0] io_out_522, // @[:@6.4]
  output [3:0] io_out_523, // @[:@6.4]
  output [3:0] io_out_524, // @[:@6.4]
  output [3:0] io_out_525, // @[:@6.4]
  output [3:0] io_out_526, // @[:@6.4]
  output [3:0] io_out_527, // @[:@6.4]
  output [3:0] io_out_528, // @[:@6.4]
  output [3:0] io_out_529, // @[:@6.4]
  output [3:0] io_out_530, // @[:@6.4]
  output [3:0] io_out_531, // @[:@6.4]
  output [3:0] io_out_532, // @[:@6.4]
  output [3:0] io_out_533, // @[:@6.4]
  output [3:0] io_out_534, // @[:@6.4]
  output [3:0] io_out_535, // @[:@6.4]
  output [3:0] io_out_536, // @[:@6.4]
  output [3:0] io_out_537, // @[:@6.4]
  output [3:0] io_out_538, // @[:@6.4]
  output [3:0] io_out_539, // @[:@6.4]
  output [3:0] io_out_540, // @[:@6.4]
  output [3:0] io_out_541, // @[:@6.4]
  output [3:0] io_out_542, // @[:@6.4]
  output [3:0] io_out_543, // @[:@6.4]
  output [3:0] io_out_544, // @[:@6.4]
  output [3:0] io_out_545, // @[:@6.4]
  output [3:0] io_out_546, // @[:@6.4]
  output [3:0] io_out_547, // @[:@6.4]
  output [3:0] io_out_548, // @[:@6.4]
  output [3:0] io_out_549, // @[:@6.4]
  output [3:0] io_out_550, // @[:@6.4]
  output [3:0] io_out_551, // @[:@6.4]
  output [3:0] io_out_552, // @[:@6.4]
  output [3:0] io_out_553, // @[:@6.4]
  output [3:0] io_out_554, // @[:@6.4]
  output [3:0] io_out_555, // @[:@6.4]
  output [3:0] io_out_556, // @[:@6.4]
  output [3:0] io_out_557, // @[:@6.4]
  output [3:0] io_out_558, // @[:@6.4]
  output [3:0] io_out_559, // @[:@6.4]
  output [3:0] io_out_560, // @[:@6.4]
  output [3:0] io_out_561, // @[:@6.4]
  output [3:0] io_out_562, // @[:@6.4]
  output [3:0] io_out_563, // @[:@6.4]
  output [3:0] io_out_564, // @[:@6.4]
  output [3:0] io_out_565, // @[:@6.4]
  output [3:0] io_out_566, // @[:@6.4]
  output [3:0] io_out_567, // @[:@6.4]
  output [3:0] io_out_568, // @[:@6.4]
  output [3:0] io_out_569, // @[:@6.4]
  output [3:0] io_out_570, // @[:@6.4]
  output [3:0] io_out_571, // @[:@6.4]
  output [3:0] io_out_572, // @[:@6.4]
  output [3:0] io_out_573, // @[:@6.4]
  output [3:0] io_out_574, // @[:@6.4]
  output [3:0] io_out_575, // @[:@6.4]
  output [3:0] io_out_576, // @[:@6.4]
  output [3:0] io_out_577, // @[:@6.4]
  output [3:0] io_out_578, // @[:@6.4]
  output [3:0] io_out_579, // @[:@6.4]
  output [3:0] io_out_580, // @[:@6.4]
  output [3:0] io_out_581, // @[:@6.4]
  output [3:0] io_out_582, // @[:@6.4]
  output [3:0] io_out_583, // @[:@6.4]
  output [3:0] io_out_584, // @[:@6.4]
  output [3:0] io_out_585, // @[:@6.4]
  output [3:0] io_out_586, // @[:@6.4]
  output [3:0] io_out_587, // @[:@6.4]
  output [3:0] io_out_588, // @[:@6.4]
  output [3:0] io_out_589, // @[:@6.4]
  output [3:0] io_out_590, // @[:@6.4]
  output [3:0] io_out_591, // @[:@6.4]
  output [3:0] io_out_592, // @[:@6.4]
  output [3:0] io_out_593, // @[:@6.4]
  output [3:0] io_out_594, // @[:@6.4]
  output [3:0] io_out_595, // @[:@6.4]
  output [3:0] io_out_596, // @[:@6.4]
  output [3:0] io_out_597, // @[:@6.4]
  output [3:0] io_out_598, // @[:@6.4]
  output [3:0] io_out_599, // @[:@6.4]
  output [3:0] io_out_600, // @[:@6.4]
  output [3:0] io_out_601, // @[:@6.4]
  output [3:0] io_out_602, // @[:@6.4]
  output [3:0] io_out_603, // @[:@6.4]
  output [3:0] io_out_604, // @[:@6.4]
  output [3:0] io_out_605, // @[:@6.4]
  output [3:0] io_out_606, // @[:@6.4]
  output [3:0] io_out_607, // @[:@6.4]
  output [3:0] io_out_608, // @[:@6.4]
  output [3:0] io_out_609, // @[:@6.4]
  output [3:0] io_out_610, // @[:@6.4]
  output [3:0] io_out_611, // @[:@6.4]
  output [3:0] io_out_612, // @[:@6.4]
  output [3:0] io_out_613, // @[:@6.4]
  output [3:0] io_out_614, // @[:@6.4]
  output [3:0] io_out_615, // @[:@6.4]
  output [3:0] io_out_616, // @[:@6.4]
  output [3:0] io_out_617, // @[:@6.4]
  output [3:0] io_out_618, // @[:@6.4]
  output [3:0] io_out_619, // @[:@6.4]
  output [3:0] io_out_620, // @[:@6.4]
  output [3:0] io_out_621, // @[:@6.4]
  output [3:0] io_out_622, // @[:@6.4]
  output [3:0] io_out_623, // @[:@6.4]
  output [3:0] io_out_624, // @[:@6.4]
  output [3:0] io_out_625, // @[:@6.4]
  output [3:0] io_out_626, // @[:@6.4]
  output [3:0] io_out_627, // @[:@6.4]
  output [3:0] io_out_628, // @[:@6.4]
  output [3:0] io_out_629, // @[:@6.4]
  output [3:0] io_out_630, // @[:@6.4]
  output [3:0] io_out_631, // @[:@6.4]
  output [3:0] io_out_632, // @[:@6.4]
  output [3:0] io_out_633, // @[:@6.4]
  output [3:0] io_out_634, // @[:@6.4]
  output [3:0] io_out_635, // @[:@6.4]
  output [3:0] io_out_636, // @[:@6.4]
  output [3:0] io_out_637, // @[:@6.4]
  output [3:0] io_out_638, // @[:@6.4]
  output [3:0] io_out_639, // @[:@6.4]
  output [3:0] io_out_640, // @[:@6.4]
  output [3:0] io_out_641, // @[:@6.4]
  output [3:0] io_out_642, // @[:@6.4]
  output [3:0] io_out_643, // @[:@6.4]
  output [3:0] io_out_644, // @[:@6.4]
  output [3:0] io_out_645, // @[:@6.4]
  output [3:0] io_out_646, // @[:@6.4]
  output [3:0] io_out_647, // @[:@6.4]
  output [3:0] io_out_648, // @[:@6.4]
  output [3:0] io_out_649, // @[:@6.4]
  output [3:0] io_out_650, // @[:@6.4]
  output [3:0] io_out_651, // @[:@6.4]
  output [3:0] io_out_652, // @[:@6.4]
  output [3:0] io_out_653, // @[:@6.4]
  output [3:0] io_out_654, // @[:@6.4]
  output [3:0] io_out_655, // @[:@6.4]
  output [3:0] io_out_656, // @[:@6.4]
  output [3:0] io_out_657, // @[:@6.4]
  output [3:0] io_out_658, // @[:@6.4]
  output [3:0] io_out_659, // @[:@6.4]
  output [3:0] io_out_660, // @[:@6.4]
  output [3:0] io_out_661, // @[:@6.4]
  output [3:0] io_out_662, // @[:@6.4]
  output [3:0] io_out_663, // @[:@6.4]
  output [3:0] io_out_664, // @[:@6.4]
  output [3:0] io_out_665, // @[:@6.4]
  output [3:0] io_out_666, // @[:@6.4]
  output [3:0] io_out_667, // @[:@6.4]
  output [3:0] io_out_668, // @[:@6.4]
  output [3:0] io_out_669, // @[:@6.4]
  output [3:0] io_out_670, // @[:@6.4]
  output [3:0] io_out_671, // @[:@6.4]
  output [3:0] io_out_672, // @[:@6.4]
  output [3:0] io_out_673, // @[:@6.4]
  output [3:0] io_out_674, // @[:@6.4]
  output [3:0] io_out_675, // @[:@6.4]
  output [3:0] io_out_676, // @[:@6.4]
  output [3:0] io_out_677, // @[:@6.4]
  output [3:0] io_out_678, // @[:@6.4]
  output [3:0] io_out_679, // @[:@6.4]
  output [3:0] io_out_680, // @[:@6.4]
  output [3:0] io_out_681, // @[:@6.4]
  output [3:0] io_out_682, // @[:@6.4]
  output [3:0] io_out_683, // @[:@6.4]
  output [3:0] io_out_684, // @[:@6.4]
  output [3:0] io_out_685, // @[:@6.4]
  output [3:0] io_out_686, // @[:@6.4]
  output [3:0] io_out_687, // @[:@6.4]
  output [3:0] io_out_688, // @[:@6.4]
  output [3:0] io_out_689, // @[:@6.4]
  output [3:0] io_out_690, // @[:@6.4]
  output [3:0] io_out_691, // @[:@6.4]
  output [3:0] io_out_692, // @[:@6.4]
  output [3:0] io_out_693, // @[:@6.4]
  output [3:0] io_out_694, // @[:@6.4]
  output [3:0] io_out_695, // @[:@6.4]
  output [3:0] io_out_696, // @[:@6.4]
  output [3:0] io_out_697, // @[:@6.4]
  output [3:0] io_out_698, // @[:@6.4]
  output [3:0] io_out_699, // @[:@6.4]
  output [3:0] io_out_700, // @[:@6.4]
  output [3:0] io_out_701, // @[:@6.4]
  output [3:0] io_out_702, // @[:@6.4]
  output [3:0] io_out_703, // @[:@6.4]
  output [3:0] io_out_704, // @[:@6.4]
  output [3:0] io_out_705, // @[:@6.4]
  output [3:0] io_out_706, // @[:@6.4]
  output [3:0] io_out_707, // @[:@6.4]
  output [3:0] io_out_708, // @[:@6.4]
  output [3:0] io_out_709, // @[:@6.4]
  output [3:0] io_out_710, // @[:@6.4]
  output [3:0] io_out_711, // @[:@6.4]
  output [3:0] io_out_712, // @[:@6.4]
  output [3:0] io_out_713, // @[:@6.4]
  output [3:0] io_out_714, // @[:@6.4]
  output [3:0] io_out_715, // @[:@6.4]
  output [3:0] io_out_716, // @[:@6.4]
  output [3:0] io_out_717, // @[:@6.4]
  output [3:0] io_out_718, // @[:@6.4]
  output [3:0] io_out_719, // @[:@6.4]
  output [3:0] io_out_720, // @[:@6.4]
  output [3:0] io_out_721, // @[:@6.4]
  output [3:0] io_out_722, // @[:@6.4]
  output [3:0] io_out_723, // @[:@6.4]
  output [3:0] io_out_724, // @[:@6.4]
  output [3:0] io_out_725, // @[:@6.4]
  output [3:0] io_out_726, // @[:@6.4]
  output [3:0] io_out_727, // @[:@6.4]
  output [3:0] io_out_728, // @[:@6.4]
  output [3:0] io_out_729, // @[:@6.4]
  output [3:0] io_out_730, // @[:@6.4]
  output [3:0] io_out_731, // @[:@6.4]
  output [3:0] io_out_732, // @[:@6.4]
  output [3:0] io_out_733, // @[:@6.4]
  output [3:0] io_out_734, // @[:@6.4]
  output [3:0] io_out_735, // @[:@6.4]
  output [3:0] io_out_736, // @[:@6.4]
  output [3:0] io_out_737, // @[:@6.4]
  output [3:0] io_out_738, // @[:@6.4]
  output [3:0] io_out_739, // @[:@6.4]
  output [3:0] io_out_740, // @[:@6.4]
  output [3:0] io_out_741, // @[:@6.4]
  output [3:0] io_out_742, // @[:@6.4]
  output [3:0] io_out_743, // @[:@6.4]
  output [3:0] io_out_744, // @[:@6.4]
  output [3:0] io_out_745, // @[:@6.4]
  output [3:0] io_out_746, // @[:@6.4]
  output [3:0] io_out_747, // @[:@6.4]
  output [3:0] io_out_748, // @[:@6.4]
  output [3:0] io_out_749, // @[:@6.4]
  output [3:0] io_out_750, // @[:@6.4]
  output [3:0] io_out_751, // @[:@6.4]
  output [3:0] io_out_752, // @[:@6.4]
  output [3:0] io_out_753, // @[:@6.4]
  output [3:0] io_out_754, // @[:@6.4]
  output [3:0] io_out_755, // @[:@6.4]
  output [3:0] io_out_756, // @[:@6.4]
  output [3:0] io_out_757, // @[:@6.4]
  output [3:0] io_out_758, // @[:@6.4]
  output [3:0] io_out_759, // @[:@6.4]
  output [3:0] io_out_760, // @[:@6.4]
  output [3:0] io_out_761, // @[:@6.4]
  output [3:0] io_out_762, // @[:@6.4]
  output [3:0] io_out_763, // @[:@6.4]
  output [3:0] io_out_764, // @[:@6.4]
  output [3:0] io_out_765, // @[:@6.4]
  output [3:0] io_out_766, // @[:@6.4]
  output [3:0] io_out_767, // @[:@6.4]
  output [3:0] io_out_768, // @[:@6.4]
  output [3:0] io_out_769, // @[:@6.4]
  output [3:0] io_out_770, // @[:@6.4]
  output [3:0] io_out_771, // @[:@6.4]
  output [3:0] io_out_772, // @[:@6.4]
  output [3:0] io_out_773, // @[:@6.4]
  output [3:0] io_out_774, // @[:@6.4]
  output [3:0] io_out_775, // @[:@6.4]
  output [3:0] io_out_776, // @[:@6.4]
  output [3:0] io_out_777, // @[:@6.4]
  output [3:0] io_out_778, // @[:@6.4]
  output [3:0] io_out_779, // @[:@6.4]
  output [3:0] io_out_780, // @[:@6.4]
  output [3:0] io_out_781, // @[:@6.4]
  output [3:0] io_out_782, // @[:@6.4]
  output [3:0] io_out_783, // @[:@6.4]
  output       io_addr // @[:@6.4]
);
  assign io_out_0 = io_in_0;
  assign io_out_1 = io_in_1;
  assign io_out_2 = io_in_2;
  assign io_out_3 = io_in_3;
  assign io_out_4 = io_in_4;
  assign io_out_5 = io_in_5;
  assign io_out_6 = io_in_6;
  assign io_out_7 = io_in_7;
  assign io_out_8 = io_in_8;
  assign io_out_9 = io_in_9;
  assign io_out_10 = io_in_10;
  assign io_out_11 = io_in_11;
  assign io_out_12 = io_in_12;
  assign io_out_13 = io_in_13;
  assign io_out_14 = io_in_14;
  assign io_out_15 = io_in_15;
  assign io_out_16 = io_in_16;
  assign io_out_17 = io_in_17;
  assign io_out_18 = io_in_18;
  assign io_out_19 = io_in_19;
  assign io_out_20 = io_in_20;
  assign io_out_21 = io_in_21;
  assign io_out_22 = io_in_22;
  assign io_out_23 = io_in_23;
  assign io_out_24 = io_in_24;
  assign io_out_25 = io_in_25;
  assign io_out_26 = io_in_26;
  assign io_out_27 = io_in_27;
  assign io_out_28 = io_in_28;
  assign io_out_29 = io_in_29;
  assign io_out_30 = io_in_30;
  assign io_out_31 = io_in_31;
  assign io_out_32 = io_in_32;
  assign io_out_33 = io_in_33;
  assign io_out_34 = io_in_34;
  assign io_out_35 = io_in_35;
  assign io_out_36 = io_in_36;
  assign io_out_37 = io_in_37;
  assign io_out_38 = io_in_38;
  assign io_out_39 = io_in_39;
  assign io_out_40 = io_in_40;
  assign io_out_41 = io_in_41;
  assign io_out_42 = io_in_42;
  assign io_out_43 = io_in_43;
  assign io_out_44 = io_in_44;
  assign io_out_45 = io_in_45;
  assign io_out_46 = io_in_46;
  assign io_out_47 = io_in_47;
  assign io_out_48 = io_in_48;
  assign io_out_49 = io_in_49;
  assign io_out_50 = io_in_50;
  assign io_out_51 = io_in_51;
  assign io_out_52 = io_in_52;
  assign io_out_53 = io_in_53;
  assign io_out_54 = io_in_54;
  assign io_out_55 = io_in_55;
  assign io_out_56 = io_in_56;
  assign io_out_57 = io_in_57;
  assign io_out_58 = io_in_58;
  assign io_out_59 = io_in_59;
  assign io_out_60 = io_in_60;
  assign io_out_61 = io_in_61;
  assign io_out_62 = io_in_62;
  assign io_out_63 = io_in_63;
  assign io_out_64 = io_in_64;
  assign io_out_65 = io_in_65;
  assign io_out_66 = io_in_66;
  assign io_out_67 = io_in_67;
  assign io_out_68 = io_in_68;
  assign io_out_69 = io_in_69;
  assign io_out_70 = io_in_70;
  assign io_out_71 = io_in_71;
  assign io_out_72 = io_in_72;
  assign io_out_73 = io_in_73;
  assign io_out_74 = io_in_74;
  assign io_out_75 = io_in_75;
  assign io_out_76 = io_in_76;
  assign io_out_77 = io_in_77;
  assign io_out_78 = io_in_78;
  assign io_out_79 = io_in_79;
  assign io_out_80 = io_in_80;
  assign io_out_81 = io_in_81;
  assign io_out_82 = io_in_82;
  assign io_out_83 = io_in_83;
  assign io_out_84 = io_in_84;
  assign io_out_85 = io_in_85;
  assign io_out_86 = io_in_86;
  assign io_out_87 = io_in_87;
  assign io_out_88 = io_in_88;
  assign io_out_89 = io_in_89;
  assign io_out_90 = io_in_90;
  assign io_out_91 = io_in_91;
  assign io_out_92 = io_in_92;
  assign io_out_93 = io_in_93;
  assign io_out_94 = io_in_94;
  assign io_out_95 = io_in_95;
  assign io_out_96 = io_in_96;
  assign io_out_97 = io_in_97;
  assign io_out_98 = io_in_98;
  assign io_out_99 = io_in_99;
  assign io_out_100 = io_in_100;
  assign io_out_101 = io_in_101;
  assign io_out_102 = io_in_102;
  assign io_out_103 = io_in_103;
  assign io_out_104 = io_in_104;
  assign io_out_105 = io_in_105;
  assign io_out_106 = io_in_106;
  assign io_out_107 = io_in_107;
  assign io_out_108 = io_in_108;
  assign io_out_109 = io_in_109;
  assign io_out_110 = io_in_110;
  assign io_out_111 = io_in_111;
  assign io_out_112 = io_in_112;
  assign io_out_113 = io_in_113;
  assign io_out_114 = io_in_114;
  assign io_out_115 = io_in_115;
  assign io_out_116 = io_in_116;
  assign io_out_117 = io_in_117;
  assign io_out_118 = io_in_118;
  assign io_out_119 = io_in_119;
  assign io_out_120 = io_in_120;
  assign io_out_121 = io_in_121;
  assign io_out_122 = io_in_122;
  assign io_out_123 = io_in_123;
  assign io_out_124 = io_in_124;
  assign io_out_125 = io_in_125;
  assign io_out_126 = io_in_126;
  assign io_out_127 = io_in_127;
  assign io_out_128 = io_in_128;
  assign io_out_129 = io_in_129;
  assign io_out_130 = io_in_130;
  assign io_out_131 = io_in_131;
  assign io_out_132 = io_in_132;
  assign io_out_133 = io_in_133;
  assign io_out_134 = io_in_134;
  assign io_out_135 = io_in_135;
  assign io_out_136 = io_in_136;
  assign io_out_137 = io_in_137;
  assign io_out_138 = io_in_138;
  assign io_out_139 = io_in_139;
  assign io_out_140 = io_in_140;
  assign io_out_141 = io_in_141;
  assign io_out_142 = io_in_142;
  assign io_out_143 = io_in_143;
  assign io_out_144 = io_in_144;
  assign io_out_145 = io_in_145;
  assign io_out_146 = io_in_146;
  assign io_out_147 = io_in_147;
  assign io_out_148 = io_in_148;
  assign io_out_149 = io_in_149;
  assign io_out_150 = io_in_150;
  assign io_out_151 = io_in_151;
  assign io_out_152 = io_in_152;
  assign io_out_153 = io_in_153;
  assign io_out_154 = io_in_154;
  assign io_out_155 = io_in_155;
  assign io_out_156 = io_in_156;
  assign io_out_157 = io_in_157;
  assign io_out_158 = io_in_158;
  assign io_out_159 = io_in_159;
  assign io_out_160 = io_in_160;
  assign io_out_161 = io_in_161;
  assign io_out_162 = io_in_162;
  assign io_out_163 = io_in_163;
  assign io_out_164 = io_in_164;
  assign io_out_165 = io_in_165;
  assign io_out_166 = io_in_166;
  assign io_out_167 = io_in_167;
  assign io_out_168 = io_in_168;
  assign io_out_169 = io_in_169;
  assign io_out_170 = io_in_170;
  assign io_out_171 = io_in_171;
  assign io_out_172 = io_in_172;
  assign io_out_173 = io_in_173;
  assign io_out_174 = io_in_174;
  assign io_out_175 = io_in_175;
  assign io_out_176 = io_in_176;
  assign io_out_177 = io_in_177;
  assign io_out_178 = io_in_178;
  assign io_out_179 = io_in_179;
  assign io_out_180 = io_in_180;
  assign io_out_181 = io_in_181;
  assign io_out_182 = io_in_182;
  assign io_out_183 = io_in_183;
  assign io_out_184 = io_in_184;
  assign io_out_185 = io_in_185;
  assign io_out_186 = io_in_186;
  assign io_out_187 = io_in_187;
  assign io_out_188 = io_in_188;
  assign io_out_189 = io_in_189;
  assign io_out_190 = io_in_190;
  assign io_out_191 = io_in_191;
  assign io_out_192 = io_in_192;
  assign io_out_193 = io_in_193;
  assign io_out_194 = io_in_194;
  assign io_out_195 = io_in_195;
  assign io_out_196 = io_in_196;
  assign io_out_197 = io_in_197;
  assign io_out_198 = io_in_198;
  assign io_out_199 = io_in_199;
  assign io_out_200 = io_in_200;
  assign io_out_201 = io_in_201;
  assign io_out_202 = io_in_202;
  assign io_out_203 = io_in_203;
  assign io_out_204 = io_in_204;
  assign io_out_205 = io_in_205;
  assign io_out_206 = io_in_206;
  assign io_out_207 = io_in_207;
  assign io_out_208 = io_in_208;
  assign io_out_209 = io_in_209;
  assign io_out_210 = io_in_210;
  assign io_out_211 = io_in_211;
  assign io_out_212 = io_in_212;
  assign io_out_213 = io_in_213;
  assign io_out_214 = io_in_214;
  assign io_out_215 = io_in_215;
  assign io_out_216 = io_in_216;
  assign io_out_217 = io_in_217;
  assign io_out_218 = io_in_218;
  assign io_out_219 = io_in_219;
  assign io_out_220 = io_in_220;
  assign io_out_221 = io_in_221;
  assign io_out_222 = io_in_222;
  assign io_out_223 = io_in_223;
  assign io_out_224 = io_in_224;
  assign io_out_225 = io_in_225;
  assign io_out_226 = io_in_226;
  assign io_out_227 = io_in_227;
  assign io_out_228 = io_in_228;
  assign io_out_229 = io_in_229;
  assign io_out_230 = io_in_230;
  assign io_out_231 = io_in_231;
  assign io_out_232 = io_in_232;
  assign io_out_233 = io_in_233;
  assign io_out_234 = io_in_234;
  assign io_out_235 = io_in_235;
  assign io_out_236 = io_in_236;
  assign io_out_237 = io_in_237;
  assign io_out_238 = io_in_238;
  assign io_out_239 = io_in_239;
  assign io_out_240 = io_in_240;
  assign io_out_241 = io_in_241;
  assign io_out_242 = io_in_242;
  assign io_out_243 = io_in_243;
  assign io_out_244 = io_in_244;
  assign io_out_245 = io_in_245;
  assign io_out_246 = io_in_246;
  assign io_out_247 = io_in_247;
  assign io_out_248 = io_in_248;
  assign io_out_249 = io_in_249;
  assign io_out_250 = io_in_250;
  assign io_out_251 = io_in_251;
  assign io_out_252 = io_in_252;
  assign io_out_253 = io_in_253;
  assign io_out_254 = io_in_254;
  assign io_out_255 = io_in_255;
  assign io_out_256 = io_in_256;
  assign io_out_257 = io_in_257;
  assign io_out_258 = io_in_258;
  assign io_out_259 = io_in_259;
  assign io_out_260 = io_in_260;
  assign io_out_261 = io_in_261;
  assign io_out_262 = io_in_262;
  assign io_out_263 = io_in_263;
  assign io_out_264 = io_in_264;
  assign io_out_265 = io_in_265;
  assign io_out_266 = io_in_266;
  assign io_out_267 = io_in_267;
  assign io_out_268 = io_in_268;
  assign io_out_269 = io_in_269;
  assign io_out_270 = io_in_270;
  assign io_out_271 = io_in_271;
  assign io_out_272 = io_in_272;
  assign io_out_273 = io_in_273;
  assign io_out_274 = io_in_274;
  assign io_out_275 = io_in_275;
  assign io_out_276 = io_in_276;
  assign io_out_277 = io_in_277;
  assign io_out_278 = io_in_278;
  assign io_out_279 = io_in_279;
  assign io_out_280 = io_in_280;
  assign io_out_281 = io_in_281;
  assign io_out_282 = io_in_282;
  assign io_out_283 = io_in_283;
  assign io_out_284 = io_in_284;
  assign io_out_285 = io_in_285;
  assign io_out_286 = io_in_286;
  assign io_out_287 = io_in_287;
  assign io_out_288 = io_in_288;
  assign io_out_289 = io_in_289;
  assign io_out_290 = io_in_290;
  assign io_out_291 = io_in_291;
  assign io_out_292 = io_in_292;
  assign io_out_293 = io_in_293;
  assign io_out_294 = io_in_294;
  assign io_out_295 = io_in_295;
  assign io_out_296 = io_in_296;
  assign io_out_297 = io_in_297;
  assign io_out_298 = io_in_298;
  assign io_out_299 = io_in_299;
  assign io_out_300 = io_in_300;
  assign io_out_301 = io_in_301;
  assign io_out_302 = io_in_302;
  assign io_out_303 = io_in_303;
  assign io_out_304 = io_in_304;
  assign io_out_305 = io_in_305;
  assign io_out_306 = io_in_306;
  assign io_out_307 = io_in_307;
  assign io_out_308 = io_in_308;
  assign io_out_309 = io_in_309;
  assign io_out_310 = io_in_310;
  assign io_out_311 = io_in_311;
  assign io_out_312 = io_in_312;
  assign io_out_313 = io_in_313;
  assign io_out_314 = io_in_314;
  assign io_out_315 = io_in_315;
  assign io_out_316 = io_in_316;
  assign io_out_317 = io_in_317;
  assign io_out_318 = io_in_318;
  assign io_out_319 = io_in_319;
  assign io_out_320 = io_in_320;
  assign io_out_321 = io_in_321;
  assign io_out_322 = io_in_322;
  assign io_out_323 = io_in_323;
  assign io_out_324 = io_in_324;
  assign io_out_325 = io_in_325;
  assign io_out_326 = io_in_326;
  assign io_out_327 = io_in_327;
  assign io_out_328 = io_in_328;
  assign io_out_329 = io_in_329;
  assign io_out_330 = io_in_330;
  assign io_out_331 = io_in_331;
  assign io_out_332 = io_in_332;
  assign io_out_333 = io_in_333;
  assign io_out_334 = io_in_334;
  assign io_out_335 = io_in_335;
  assign io_out_336 = io_in_336;
  assign io_out_337 = io_in_337;
  assign io_out_338 = io_in_338;
  assign io_out_339 = io_in_339;
  assign io_out_340 = io_in_340;
  assign io_out_341 = io_in_341;
  assign io_out_342 = io_in_342;
  assign io_out_343 = io_in_343;
  assign io_out_344 = io_in_344;
  assign io_out_345 = io_in_345;
  assign io_out_346 = io_in_346;
  assign io_out_347 = io_in_347;
  assign io_out_348 = io_in_348;
  assign io_out_349 = io_in_349;
  assign io_out_350 = io_in_350;
  assign io_out_351 = io_in_351;
  assign io_out_352 = io_in_352;
  assign io_out_353 = io_in_353;
  assign io_out_354 = io_in_354;
  assign io_out_355 = io_in_355;
  assign io_out_356 = io_in_356;
  assign io_out_357 = io_in_357;
  assign io_out_358 = io_in_358;
  assign io_out_359 = io_in_359;
  assign io_out_360 = io_in_360;
  assign io_out_361 = io_in_361;
  assign io_out_362 = io_in_362;
  assign io_out_363 = io_in_363;
  assign io_out_364 = io_in_364;
  assign io_out_365 = io_in_365;
  assign io_out_366 = io_in_366;
  assign io_out_367 = io_in_367;
  assign io_out_368 = io_in_368;
  assign io_out_369 = io_in_369;
  assign io_out_370 = io_in_370;
  assign io_out_371 = io_in_371;
  assign io_out_372 = io_in_372;
  assign io_out_373 = io_in_373;
  assign io_out_374 = io_in_374;
  assign io_out_375 = io_in_375;
  assign io_out_376 = io_in_376;
  assign io_out_377 = io_in_377;
  assign io_out_378 = io_in_378;
  assign io_out_379 = io_in_379;
  assign io_out_380 = io_in_380;
  assign io_out_381 = io_in_381;
  assign io_out_382 = io_in_382;
  assign io_out_383 = io_in_383;
  assign io_out_384 = io_in_384;
  assign io_out_385 = io_in_385;
  assign io_out_386 = io_in_386;
  assign io_out_387 = io_in_387;
  assign io_out_388 = io_in_388;
  assign io_out_389 = io_in_389;
  assign io_out_390 = io_in_390;
  assign io_out_391 = io_in_391;
  assign io_out_392 = io_in_392;
  assign io_out_393 = io_in_393;
  assign io_out_394 = io_in_394;
  assign io_out_395 = io_in_395;
  assign io_out_396 = io_in_396;
  assign io_out_397 = io_in_397;
  assign io_out_398 = io_in_398;
  assign io_out_399 = io_in_399;
  assign io_out_400 = io_in_400;
  assign io_out_401 = io_in_401;
  assign io_out_402 = io_in_402;
  assign io_out_403 = io_in_403;
  assign io_out_404 = io_in_404;
  assign io_out_405 = io_in_405;
  assign io_out_406 = io_in_406;
  assign io_out_407 = io_in_407;
  assign io_out_408 = io_in_408;
  assign io_out_409 = io_in_409;
  assign io_out_410 = io_in_410;
  assign io_out_411 = io_in_411;
  assign io_out_412 = io_in_412;
  assign io_out_413 = io_in_413;
  assign io_out_414 = io_in_414;
  assign io_out_415 = io_in_415;
  assign io_out_416 = io_in_416;
  assign io_out_417 = io_in_417;
  assign io_out_418 = io_in_418;
  assign io_out_419 = io_in_419;
  assign io_out_420 = io_in_420;
  assign io_out_421 = io_in_421;
  assign io_out_422 = io_in_422;
  assign io_out_423 = io_in_423;
  assign io_out_424 = io_in_424;
  assign io_out_425 = io_in_425;
  assign io_out_426 = io_in_426;
  assign io_out_427 = io_in_427;
  assign io_out_428 = io_in_428;
  assign io_out_429 = io_in_429;
  assign io_out_430 = io_in_430;
  assign io_out_431 = io_in_431;
  assign io_out_432 = io_in_432;
  assign io_out_433 = io_in_433;
  assign io_out_434 = io_in_434;
  assign io_out_435 = io_in_435;
  assign io_out_436 = io_in_436;
  assign io_out_437 = io_in_437;
  assign io_out_438 = io_in_438;
  assign io_out_439 = io_in_439;
  assign io_out_440 = io_in_440;
  assign io_out_441 = io_in_441;
  assign io_out_442 = io_in_442;
  assign io_out_443 = io_in_443;
  assign io_out_444 = io_in_444;
  assign io_out_445 = io_in_445;
  assign io_out_446 = io_in_446;
  assign io_out_447 = io_in_447;
  assign io_out_448 = io_in_448;
  assign io_out_449 = io_in_449;
  assign io_out_450 = io_in_450;
  assign io_out_451 = io_in_451;
  assign io_out_452 = io_in_452;
  assign io_out_453 = io_in_453;
  assign io_out_454 = io_in_454;
  assign io_out_455 = io_in_455;
  assign io_out_456 = io_in_456;
  assign io_out_457 = io_in_457;
  assign io_out_458 = io_in_458;
  assign io_out_459 = io_in_459;
  assign io_out_460 = io_in_460;
  assign io_out_461 = io_in_461;
  assign io_out_462 = io_in_462;
  assign io_out_463 = io_in_463;
  assign io_out_464 = io_in_464;
  assign io_out_465 = io_in_465;
  assign io_out_466 = io_in_466;
  assign io_out_467 = io_in_467;
  assign io_out_468 = io_in_468;
  assign io_out_469 = io_in_469;
  assign io_out_470 = io_in_470;
  assign io_out_471 = io_in_471;
  assign io_out_472 = io_in_472;
  assign io_out_473 = io_in_473;
  assign io_out_474 = io_in_474;
  assign io_out_475 = io_in_475;
  assign io_out_476 = io_in_476;
  assign io_out_477 = io_in_477;
  assign io_out_478 = io_in_478;
  assign io_out_479 = io_in_479;
  assign io_out_480 = io_in_480;
  assign io_out_481 = io_in_481;
  assign io_out_482 = io_in_482;
  assign io_out_483 = io_in_483;
  assign io_out_484 = io_in_484;
  assign io_out_485 = io_in_485;
  assign io_out_486 = io_in_486;
  assign io_out_487 = io_in_487;
  assign io_out_488 = io_in_488;
  assign io_out_489 = io_in_489;
  assign io_out_490 = io_in_490;
  assign io_out_491 = io_in_491;
  assign io_out_492 = io_in_492;
  assign io_out_493 = io_in_493;
  assign io_out_494 = io_in_494;
  assign io_out_495 = io_in_495;
  assign io_out_496 = io_in_496;
  assign io_out_497 = io_in_497;
  assign io_out_498 = io_in_498;
  assign io_out_499 = io_in_499;
  assign io_out_500 = io_in_500;
  assign io_out_501 = io_in_501;
  assign io_out_502 = io_in_502;
  assign io_out_503 = io_in_503;
  assign io_out_504 = io_in_504;
  assign io_out_505 = io_in_505;
  assign io_out_506 = io_in_506;
  assign io_out_507 = io_in_507;
  assign io_out_508 = io_in_508;
  assign io_out_509 = io_in_509;
  assign io_out_510 = io_in_510;
  assign io_out_511 = io_in_511;
  assign io_out_512 = io_in_512;
  assign io_out_513 = io_in_513;
  assign io_out_514 = io_in_514;
  assign io_out_515 = io_in_515;
  assign io_out_516 = io_in_516;
  assign io_out_517 = io_in_517;
  assign io_out_518 = io_in_518;
  assign io_out_519 = io_in_519;
  assign io_out_520 = io_in_520;
  assign io_out_521 = io_in_521;
  assign io_out_522 = io_in_522;
  assign io_out_523 = io_in_523;
  assign io_out_524 = io_in_524;
  assign io_out_525 = io_in_525;
  assign io_out_526 = io_in_526;
  assign io_out_527 = io_in_527;
  assign io_out_528 = io_in_528;
  assign io_out_529 = io_in_529;
  assign io_out_530 = io_in_530;
  assign io_out_531 = io_in_531;
  assign io_out_532 = io_in_532;
  assign io_out_533 = io_in_533;
  assign io_out_534 = io_in_534;
  assign io_out_535 = io_in_535;
  assign io_out_536 = io_in_536;
  assign io_out_537 = io_in_537;
  assign io_out_538 = io_in_538;
  assign io_out_539 = io_in_539;
  assign io_out_540 = io_in_540;
  assign io_out_541 = io_in_541;
  assign io_out_542 = io_in_542;
  assign io_out_543 = io_in_543;
  assign io_out_544 = io_in_544;
  assign io_out_545 = io_in_545;
  assign io_out_546 = io_in_546;
  assign io_out_547 = io_in_547;
  assign io_out_548 = io_in_548;
  assign io_out_549 = io_in_549;
  assign io_out_550 = io_in_550;
  assign io_out_551 = io_in_551;
  assign io_out_552 = io_in_552;
  assign io_out_553 = io_in_553;
  assign io_out_554 = io_in_554;
  assign io_out_555 = io_in_555;
  assign io_out_556 = io_in_556;
  assign io_out_557 = io_in_557;
  assign io_out_558 = io_in_558;
  assign io_out_559 = io_in_559;
  assign io_out_560 = io_in_560;
  assign io_out_561 = io_in_561;
  assign io_out_562 = io_in_562;
  assign io_out_563 = io_in_563;
  assign io_out_564 = io_in_564;
  assign io_out_565 = io_in_565;
  assign io_out_566 = io_in_566;
  assign io_out_567 = io_in_567;
  assign io_out_568 = io_in_568;
  assign io_out_569 = io_in_569;
  assign io_out_570 = io_in_570;
  assign io_out_571 = io_in_571;
  assign io_out_572 = io_in_572;
  assign io_out_573 = io_in_573;
  assign io_out_574 = io_in_574;
  assign io_out_575 = io_in_575;
  assign io_out_576 = io_in_576;
  assign io_out_577 = io_in_577;
  assign io_out_578 = io_in_578;
  assign io_out_579 = io_in_579;
  assign io_out_580 = io_in_580;
  assign io_out_581 = io_in_581;
  assign io_out_582 = io_in_582;
  assign io_out_583 = io_in_583;
  assign io_out_584 = io_in_584;
  assign io_out_585 = io_in_585;
  assign io_out_586 = io_in_586;
  assign io_out_587 = io_in_587;
  assign io_out_588 = io_in_588;
  assign io_out_589 = io_in_589;
  assign io_out_590 = io_in_590;
  assign io_out_591 = io_in_591;
  assign io_out_592 = io_in_592;
  assign io_out_593 = io_in_593;
  assign io_out_594 = io_in_594;
  assign io_out_595 = io_in_595;
  assign io_out_596 = io_in_596;
  assign io_out_597 = io_in_597;
  assign io_out_598 = io_in_598;
  assign io_out_599 = io_in_599;
  assign io_out_600 = io_in_600;
  assign io_out_601 = io_in_601;
  assign io_out_602 = io_in_602;
  assign io_out_603 = io_in_603;
  assign io_out_604 = io_in_604;
  assign io_out_605 = io_in_605;
  assign io_out_606 = io_in_606;
  assign io_out_607 = io_in_607;
  assign io_out_608 = io_in_608;
  assign io_out_609 = io_in_609;
  assign io_out_610 = io_in_610;
  assign io_out_611 = io_in_611;
  assign io_out_612 = io_in_612;
  assign io_out_613 = io_in_613;
  assign io_out_614 = io_in_614;
  assign io_out_615 = io_in_615;
  assign io_out_616 = io_in_616;
  assign io_out_617 = io_in_617;
  assign io_out_618 = io_in_618;
  assign io_out_619 = io_in_619;
  assign io_out_620 = io_in_620;
  assign io_out_621 = io_in_621;
  assign io_out_622 = io_in_622;
  assign io_out_623 = io_in_623;
  assign io_out_624 = io_in_624;
  assign io_out_625 = io_in_625;
  assign io_out_626 = io_in_626;
  assign io_out_627 = io_in_627;
  assign io_out_628 = io_in_628;
  assign io_out_629 = io_in_629;
  assign io_out_630 = io_in_630;
  assign io_out_631 = io_in_631;
  assign io_out_632 = io_in_632;
  assign io_out_633 = io_in_633;
  assign io_out_634 = io_in_634;
  assign io_out_635 = io_in_635;
  assign io_out_636 = io_in_636;
  assign io_out_637 = io_in_637;
  assign io_out_638 = io_in_638;
  assign io_out_639 = io_in_639;
  assign io_out_640 = io_in_640;
  assign io_out_641 = io_in_641;
  assign io_out_642 = io_in_642;
  assign io_out_643 = io_in_643;
  assign io_out_644 = io_in_644;
  assign io_out_645 = io_in_645;
  assign io_out_646 = io_in_646;
  assign io_out_647 = io_in_647;
  assign io_out_648 = io_in_648;
  assign io_out_649 = io_in_649;
  assign io_out_650 = io_in_650;
  assign io_out_651 = io_in_651;
  assign io_out_652 = io_in_652;
  assign io_out_653 = io_in_653;
  assign io_out_654 = io_in_654;
  assign io_out_655 = io_in_655;
  assign io_out_656 = io_in_656;
  assign io_out_657 = io_in_657;
  assign io_out_658 = io_in_658;
  assign io_out_659 = io_in_659;
  assign io_out_660 = io_in_660;
  assign io_out_661 = io_in_661;
  assign io_out_662 = io_in_662;
  assign io_out_663 = io_in_663;
  assign io_out_664 = io_in_664;
  assign io_out_665 = io_in_665;
  assign io_out_666 = io_in_666;
  assign io_out_667 = io_in_667;
  assign io_out_668 = io_in_668;
  assign io_out_669 = io_in_669;
  assign io_out_670 = io_in_670;
  assign io_out_671 = io_in_671;
  assign io_out_672 = io_in_672;
  assign io_out_673 = io_in_673;
  assign io_out_674 = io_in_674;
  assign io_out_675 = io_in_675;
  assign io_out_676 = io_in_676;
  assign io_out_677 = io_in_677;
  assign io_out_678 = io_in_678;
  assign io_out_679 = io_in_679;
  assign io_out_680 = io_in_680;
  assign io_out_681 = io_in_681;
  assign io_out_682 = io_in_682;
  assign io_out_683 = io_in_683;
  assign io_out_684 = io_in_684;
  assign io_out_685 = io_in_685;
  assign io_out_686 = io_in_686;
  assign io_out_687 = io_in_687;
  assign io_out_688 = io_in_688;
  assign io_out_689 = io_in_689;
  assign io_out_690 = io_in_690;
  assign io_out_691 = io_in_691;
  assign io_out_692 = io_in_692;
  assign io_out_693 = io_in_693;
  assign io_out_694 = io_in_694;
  assign io_out_695 = io_in_695;
  assign io_out_696 = io_in_696;
  assign io_out_697 = io_in_697;
  assign io_out_698 = io_in_698;
  assign io_out_699 = io_in_699;
  assign io_out_700 = io_in_700;
  assign io_out_701 = io_in_701;
  assign io_out_702 = io_in_702;
  assign io_out_703 = io_in_703;
  assign io_out_704 = io_in_704;
  assign io_out_705 = io_in_705;
  assign io_out_706 = io_in_706;
  assign io_out_707 = io_in_707;
  assign io_out_708 = io_in_708;
  assign io_out_709 = io_in_709;
  assign io_out_710 = io_in_710;
  assign io_out_711 = io_in_711;
  assign io_out_712 = io_in_712;
  assign io_out_713 = io_in_713;
  assign io_out_714 = io_in_714;
  assign io_out_715 = io_in_715;
  assign io_out_716 = io_in_716;
  assign io_out_717 = io_in_717;
  assign io_out_718 = io_in_718;
  assign io_out_719 = io_in_719;
  assign io_out_720 = io_in_720;
  assign io_out_721 = io_in_721;
  assign io_out_722 = io_in_722;
  assign io_out_723 = io_in_723;
  assign io_out_724 = io_in_724;
  assign io_out_725 = io_in_725;
  assign io_out_726 = io_in_726;
  assign io_out_727 = io_in_727;
  assign io_out_728 = io_in_728;
  assign io_out_729 = io_in_729;
  assign io_out_730 = io_in_730;
  assign io_out_731 = io_in_731;
  assign io_out_732 = io_in_732;
  assign io_out_733 = io_in_733;
  assign io_out_734 = io_in_734;
  assign io_out_735 = io_in_735;
  assign io_out_736 = io_in_736;
  assign io_out_737 = io_in_737;
  assign io_out_738 = io_in_738;
  assign io_out_739 = io_in_739;
  assign io_out_740 = io_in_740;
  assign io_out_741 = io_in_741;
  assign io_out_742 = io_in_742;
  assign io_out_743 = io_in_743;
  assign io_out_744 = io_in_744;
  assign io_out_745 = io_in_745;
  assign io_out_746 = io_in_746;
  assign io_out_747 = io_in_747;
  assign io_out_748 = io_in_748;
  assign io_out_749 = io_in_749;
  assign io_out_750 = io_in_750;
  assign io_out_751 = io_in_751;
  assign io_out_752 = io_in_752;
  assign io_out_753 = io_in_753;
  assign io_out_754 = io_in_754;
  assign io_out_755 = io_in_755;
  assign io_out_756 = io_in_756;
  assign io_out_757 = io_in_757;
  assign io_out_758 = io_in_758;
  assign io_out_759 = io_in_759;
  assign io_out_760 = io_in_760;
  assign io_out_761 = io_in_761;
  assign io_out_762 = io_in_762;
  assign io_out_763 = io_in_763;
  assign io_out_764 = io_in_764;
  assign io_out_765 = io_in_765;
  assign io_out_766 = io_in_766;
  assign io_out_767 = io_in_767;
  assign io_out_768 = io_in_768;
  assign io_out_769 = io_in_769;
  assign io_out_770 = io_in_770;
  assign io_out_771 = io_in_771;
  assign io_out_772 = io_in_772;
  assign io_out_773 = io_in_773;
  assign io_out_774 = io_in_774;
  assign io_out_775 = io_in_775;
  assign io_out_776 = io_in_776;
  assign io_out_777 = io_in_777;
  assign io_out_778 = io_in_778;
  assign io_out_779 = io_in_779;
  assign io_out_780 = io_in_780;
  assign io_out_781 = io_in_781;
  assign io_out_782 = io_in_782;
  assign io_out_783 = io_in_783;
  assign io_addr = 1'h0;
endmodule
