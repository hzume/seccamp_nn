`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Linear_p( // @[:@3.2]
  input  [4:0]  io_in_0, // @[:@6.4]
  input  [4:0]  io_in_1, // @[:@6.4]
  input  [4:0]  io_in_2, // @[:@6.4]
  input  [4:0]  io_in_3, // @[:@6.4]
  input  [4:0]  io_in_4, // @[:@6.4]
  input  [4:0]  io_in_5, // @[:@6.4]
  input  [4:0]  io_in_6, // @[:@6.4]
  input  [4:0]  io_in_7, // @[:@6.4]
  input  [4:0]  io_in_8, // @[:@6.4]
  input  [4:0]  io_in_9, // @[:@6.4]
  input  [4:0]  io_in_10, // @[:@6.4]
  input  [4:0]  io_in_11, // @[:@6.4]
  input  [4:0]  io_in_12, // @[:@6.4]
  input  [4:0]  io_in_13, // @[:@6.4]
  input  [4:0]  io_in_14, // @[:@6.4]
  input  [4:0]  io_in_15, // @[:@6.4]
  input  [4:0]  io_in_16, // @[:@6.4]
  input  [4:0]  io_in_17, // @[:@6.4]
  input  [4:0]  io_in_18, // @[:@6.4]
  input  [4:0]  io_in_19, // @[:@6.4]
  input  [4:0]  io_in_20, // @[:@6.4]
  input  [4:0]  io_in_21, // @[:@6.4]
  input  [4:0]  io_in_22, // @[:@6.4]
  input  [4:0]  io_in_23, // @[:@6.4]
  input  [4:0]  io_in_24, // @[:@6.4]
  input  [4:0]  io_in_25, // @[:@6.4]
  input  [4:0]  io_in_26, // @[:@6.4]
  input  [4:0]  io_in_27, // @[:@6.4]
  input  [4:0]  io_in_28, // @[:@6.4]
  input  [4:0]  io_in_29, // @[:@6.4]
  input  [4:0]  io_in_30, // @[:@6.4]
  input  [4:0]  io_in_31, // @[:@6.4]
  input  [4:0]  io_in_32, // @[:@6.4]
  input  [4:0]  io_in_33, // @[:@6.4]
  input  [4:0]  io_in_34, // @[:@6.4]
  input  [4:0]  io_in_35, // @[:@6.4]
  input  [4:0]  io_in_36, // @[:@6.4]
  input  [4:0]  io_in_37, // @[:@6.4]
  input  [4:0]  io_in_38, // @[:@6.4]
  input  [4:0]  io_in_39, // @[:@6.4]
  input  [4:0]  io_in_40, // @[:@6.4]
  input  [4:0]  io_in_41, // @[:@6.4]
  input  [4:0]  io_in_42, // @[:@6.4]
  input  [4:0]  io_in_43, // @[:@6.4]
  input  [4:0]  io_in_44, // @[:@6.4]
  input  [4:0]  io_in_45, // @[:@6.4]
  input  [4:0]  io_in_46, // @[:@6.4]
  input  [4:0]  io_in_47, // @[:@6.4]
  input  [4:0]  io_in_48, // @[:@6.4]
  input  [4:0]  io_in_49, // @[:@6.4]
  input  [4:0]  io_in_50, // @[:@6.4]
  input  [4:0]  io_in_51, // @[:@6.4]
  input  [4:0]  io_in_52, // @[:@6.4]
  input  [4:0]  io_in_53, // @[:@6.4]
  input  [4:0]  io_in_54, // @[:@6.4]
  input  [4:0]  io_in_55, // @[:@6.4]
  input  [4:0]  io_in_56, // @[:@6.4]
  input  [4:0]  io_in_57, // @[:@6.4]
  input  [4:0]  io_in_58, // @[:@6.4]
  input  [4:0]  io_in_59, // @[:@6.4]
  input  [4:0]  io_in_60, // @[:@6.4]
  input  [4:0]  io_in_61, // @[:@6.4]
  input  [4:0]  io_in_62, // @[:@6.4]
  input  [4:0]  io_in_63, // @[:@6.4]
  input  [4:0]  io_in_64, // @[:@6.4]
  input  [4:0]  io_in_65, // @[:@6.4]
  input  [4:0]  io_in_66, // @[:@6.4]
  input  [4:0]  io_in_67, // @[:@6.4]
  input  [4:0]  io_in_68, // @[:@6.4]
  input  [4:0]  io_in_69, // @[:@6.4]
  input  [4:0]  io_in_70, // @[:@6.4]
  input  [4:0]  io_in_71, // @[:@6.4]
  input  [4:0]  io_in_72, // @[:@6.4]
  input  [4:0]  io_in_73, // @[:@6.4]
  input  [4:0]  io_in_74, // @[:@6.4]
  input  [4:0]  io_in_75, // @[:@6.4]
  input  [4:0]  io_in_76, // @[:@6.4]
  input  [4:0]  io_in_77, // @[:@6.4]
  input  [4:0]  io_in_78, // @[:@6.4]
  input  [4:0]  io_in_79, // @[:@6.4]
  input  [4:0]  io_in_80, // @[:@6.4]
  input  [4:0]  io_in_81, // @[:@6.4]
  input  [4:0]  io_in_82, // @[:@6.4]
  input  [4:0]  io_in_83, // @[:@6.4]
  input  [4:0]  io_in_84, // @[:@6.4]
  input  [4:0]  io_in_85, // @[:@6.4]
  input  [4:0]  io_in_86, // @[:@6.4]
  input  [4:0]  io_in_87, // @[:@6.4]
  input  [4:0]  io_in_88, // @[:@6.4]
  input  [4:0]  io_in_89, // @[:@6.4]
  input  [4:0]  io_in_90, // @[:@6.4]
  input  [4:0]  io_in_91, // @[:@6.4]
  input  [4:0]  io_in_92, // @[:@6.4]
  input  [4:0]  io_in_93, // @[:@6.4]
  input  [4:0]  io_in_94, // @[:@6.4]
  input  [4:0]  io_in_95, // @[:@6.4]
  input  [4:0]  io_in_96, // @[:@6.4]
  input  [4:0]  io_in_97, // @[:@6.4]
  input  [4:0]  io_in_98, // @[:@6.4]
  input  [4:0]  io_in_99, // @[:@6.4]
  input  [4:0]  io_in_100, // @[:@6.4]
  input  [4:0]  io_in_101, // @[:@6.4]
  input  [4:0]  io_in_102, // @[:@6.4]
  input  [4:0]  io_in_103, // @[:@6.4]
  input  [4:0]  io_in_104, // @[:@6.4]
  input  [4:0]  io_in_105, // @[:@6.4]
  input  [4:0]  io_in_106, // @[:@6.4]
  input  [4:0]  io_in_107, // @[:@6.4]
  input  [4:0]  io_in_108, // @[:@6.4]
  input  [4:0]  io_in_109, // @[:@6.4]
  input  [4:0]  io_in_110, // @[:@6.4]
  input  [4:0]  io_in_111, // @[:@6.4]
  input  [4:0]  io_in_112, // @[:@6.4]
  input  [4:0]  io_in_113, // @[:@6.4]
  input  [4:0]  io_in_114, // @[:@6.4]
  input  [4:0]  io_in_115, // @[:@6.4]
  input  [4:0]  io_in_116, // @[:@6.4]
  input  [4:0]  io_in_117, // @[:@6.4]
  input  [4:0]  io_in_118, // @[:@6.4]
  input  [4:0]  io_in_119, // @[:@6.4]
  input  [4:0]  io_in_120, // @[:@6.4]
  input  [4:0]  io_in_121, // @[:@6.4]
  input  [4:0]  io_in_122, // @[:@6.4]
  input  [4:0]  io_in_123, // @[:@6.4]
  input  [4:0]  io_in_124, // @[:@6.4]
  input  [4:0]  io_in_125, // @[:@6.4]
  input  [4:0]  io_in_126, // @[:@6.4]
  input  [4:0]  io_in_127, // @[:@6.4]
  input  [4:0]  io_in_128, // @[:@6.4]
  input  [4:0]  io_in_129, // @[:@6.4]
  input  [4:0]  io_in_130, // @[:@6.4]
  input  [4:0]  io_in_131, // @[:@6.4]
  input  [4:0]  io_in_132, // @[:@6.4]
  input  [4:0]  io_in_133, // @[:@6.4]
  input  [4:0]  io_in_134, // @[:@6.4]
  input  [4:0]  io_in_135, // @[:@6.4]
  input  [4:0]  io_in_136, // @[:@6.4]
  input  [4:0]  io_in_137, // @[:@6.4]
  input  [4:0]  io_in_138, // @[:@6.4]
  input  [4:0]  io_in_139, // @[:@6.4]
  input  [4:0]  io_in_140, // @[:@6.4]
  input  [4:0]  io_in_141, // @[:@6.4]
  input  [4:0]  io_in_142, // @[:@6.4]
  input  [4:0]  io_in_143, // @[:@6.4]
  input  [4:0]  io_in_144, // @[:@6.4]
  input  [4:0]  io_in_145, // @[:@6.4]
  input  [4:0]  io_in_146, // @[:@6.4]
  input  [4:0]  io_in_147, // @[:@6.4]
  input  [4:0]  io_in_148, // @[:@6.4]
  input  [4:0]  io_in_149, // @[:@6.4]
  input  [4:0]  io_in_150, // @[:@6.4]
  input  [4:0]  io_in_151, // @[:@6.4]
  input  [4:0]  io_in_152, // @[:@6.4]
  input  [4:0]  io_in_153, // @[:@6.4]
  input  [4:0]  io_in_154, // @[:@6.4]
  input  [4:0]  io_in_155, // @[:@6.4]
  input  [4:0]  io_in_156, // @[:@6.4]
  input  [4:0]  io_in_157, // @[:@6.4]
  input  [4:0]  io_in_158, // @[:@6.4]
  input  [4:0]  io_in_159, // @[:@6.4]
  input  [4:0]  io_in_160, // @[:@6.4]
  input  [4:0]  io_in_161, // @[:@6.4]
  input  [4:0]  io_in_162, // @[:@6.4]
  input  [4:0]  io_in_163, // @[:@6.4]
  input  [4:0]  io_in_164, // @[:@6.4]
  input  [4:0]  io_in_165, // @[:@6.4]
  input  [4:0]  io_in_166, // @[:@6.4]
  input  [4:0]  io_in_167, // @[:@6.4]
  input  [4:0]  io_in_168, // @[:@6.4]
  input  [4:0]  io_in_169, // @[:@6.4]
  input  [4:0]  io_in_170, // @[:@6.4]
  input  [4:0]  io_in_171, // @[:@6.4]
  input  [4:0]  io_in_172, // @[:@6.4]
  input  [4:0]  io_in_173, // @[:@6.4]
  input  [4:0]  io_in_174, // @[:@6.4]
  input  [4:0]  io_in_175, // @[:@6.4]
  input  [4:0]  io_in_176, // @[:@6.4]
  input  [4:0]  io_in_177, // @[:@6.4]
  input  [4:0]  io_in_178, // @[:@6.4]
  input  [4:0]  io_in_179, // @[:@6.4]
  input  [4:0]  io_in_180, // @[:@6.4]
  input  [4:0]  io_in_181, // @[:@6.4]
  input  [4:0]  io_in_182, // @[:@6.4]
  input  [4:0]  io_in_183, // @[:@6.4]
  input  [4:0]  io_in_184, // @[:@6.4]
  input  [4:0]  io_in_185, // @[:@6.4]
  input  [4:0]  io_in_186, // @[:@6.4]
  input  [4:0]  io_in_187, // @[:@6.4]
  input  [4:0]  io_in_188, // @[:@6.4]
  input  [4:0]  io_in_189, // @[:@6.4]
  input  [4:0]  io_in_190, // @[:@6.4]
  input  [4:0]  io_in_191, // @[:@6.4]
  input  [4:0]  io_in_192, // @[:@6.4]
  input  [4:0]  io_in_193, // @[:@6.4]
  input  [4:0]  io_in_194, // @[:@6.4]
  input  [4:0]  io_in_195, // @[:@6.4]
  input  [4:0]  io_in_196, // @[:@6.4]
  input  [4:0]  io_in_197, // @[:@6.4]
  input  [4:0]  io_in_198, // @[:@6.4]
  input  [4:0]  io_in_199, // @[:@6.4]
  input  [4:0]  io_in_200, // @[:@6.4]
  input  [4:0]  io_in_201, // @[:@6.4]
  input  [4:0]  io_in_202, // @[:@6.4]
  input  [4:0]  io_in_203, // @[:@6.4]
  input  [4:0]  io_in_204, // @[:@6.4]
  input  [4:0]  io_in_205, // @[:@6.4]
  input  [4:0]  io_in_206, // @[:@6.4]
  input  [4:0]  io_in_207, // @[:@6.4]
  input  [4:0]  io_in_208, // @[:@6.4]
  input  [4:0]  io_in_209, // @[:@6.4]
  input  [4:0]  io_in_210, // @[:@6.4]
  input  [4:0]  io_in_211, // @[:@6.4]
  input  [4:0]  io_in_212, // @[:@6.4]
  input  [4:0]  io_in_213, // @[:@6.4]
  input  [4:0]  io_in_214, // @[:@6.4]
  input  [4:0]  io_in_215, // @[:@6.4]
  input  [4:0]  io_in_216, // @[:@6.4]
  input  [4:0]  io_in_217, // @[:@6.4]
  input  [4:0]  io_in_218, // @[:@6.4]
  input  [4:0]  io_in_219, // @[:@6.4]
  input  [4:0]  io_in_220, // @[:@6.4]
  input  [4:0]  io_in_221, // @[:@6.4]
  input  [4:0]  io_in_222, // @[:@6.4]
  input  [4:0]  io_in_223, // @[:@6.4]
  input  [4:0]  io_in_224, // @[:@6.4]
  input  [4:0]  io_in_225, // @[:@6.4]
  input  [4:0]  io_in_226, // @[:@6.4]
  input  [4:0]  io_in_227, // @[:@6.4]
  input  [4:0]  io_in_228, // @[:@6.4]
  input  [4:0]  io_in_229, // @[:@6.4]
  input  [4:0]  io_in_230, // @[:@6.4]
  input  [4:0]  io_in_231, // @[:@6.4]
  input  [4:0]  io_in_232, // @[:@6.4]
  input  [4:0]  io_in_233, // @[:@6.4]
  input  [4:0]  io_in_234, // @[:@6.4]
  input  [4:0]  io_in_235, // @[:@6.4]
  input  [4:0]  io_in_236, // @[:@6.4]
  input  [4:0]  io_in_237, // @[:@6.4]
  input  [4:0]  io_in_238, // @[:@6.4]
  input  [4:0]  io_in_239, // @[:@6.4]
  input  [4:0]  io_in_240, // @[:@6.4]
  input  [4:0]  io_in_241, // @[:@6.4]
  input  [4:0]  io_in_242, // @[:@6.4]
  input  [4:0]  io_in_243, // @[:@6.4]
  input  [4:0]  io_in_244, // @[:@6.4]
  input  [4:0]  io_in_245, // @[:@6.4]
  input  [4:0]  io_in_246, // @[:@6.4]
  input  [4:0]  io_in_247, // @[:@6.4]
  input  [4:0]  io_in_248, // @[:@6.4]
  input  [4:0]  io_in_249, // @[:@6.4]
  input  [4:0]  io_in_250, // @[:@6.4]
  input  [4:0]  io_in_251, // @[:@6.4]
  input  [4:0]  io_in_252, // @[:@6.4]
  input  [4:0]  io_in_253, // @[:@6.4]
  input  [4:0]  io_in_254, // @[:@6.4]
  input  [4:0]  io_in_255, // @[:@6.4]
  input  [4:0]  io_in_256, // @[:@6.4]
  input  [4:0]  io_in_257, // @[:@6.4]
  input  [4:0]  io_in_258, // @[:@6.4]
  input  [4:0]  io_in_259, // @[:@6.4]
  input  [4:0]  io_in_260, // @[:@6.4]
  input  [4:0]  io_in_261, // @[:@6.4]
  input  [4:0]  io_in_262, // @[:@6.4]
  input  [4:0]  io_in_263, // @[:@6.4]
  input  [4:0]  io_in_264, // @[:@6.4]
  input  [4:0]  io_in_265, // @[:@6.4]
  input  [4:0]  io_in_266, // @[:@6.4]
  input  [4:0]  io_in_267, // @[:@6.4]
  input  [4:0]  io_in_268, // @[:@6.4]
  input  [4:0]  io_in_269, // @[:@6.4]
  input  [4:0]  io_in_270, // @[:@6.4]
  input  [4:0]  io_in_271, // @[:@6.4]
  input  [4:0]  io_in_272, // @[:@6.4]
  input  [4:0]  io_in_273, // @[:@6.4]
  input  [4:0]  io_in_274, // @[:@6.4]
  input  [4:0]  io_in_275, // @[:@6.4]
  input  [4:0]  io_in_276, // @[:@6.4]
  input  [4:0]  io_in_277, // @[:@6.4]
  input  [4:0]  io_in_278, // @[:@6.4]
  input  [4:0]  io_in_279, // @[:@6.4]
  input  [4:0]  io_in_280, // @[:@6.4]
  input  [4:0]  io_in_281, // @[:@6.4]
  input  [4:0]  io_in_282, // @[:@6.4]
  input  [4:0]  io_in_283, // @[:@6.4]
  input  [4:0]  io_in_284, // @[:@6.4]
  input  [4:0]  io_in_285, // @[:@6.4]
  input  [4:0]  io_in_286, // @[:@6.4]
  input  [4:0]  io_in_287, // @[:@6.4]
  input  [4:0]  io_in_288, // @[:@6.4]
  input  [4:0]  io_in_289, // @[:@6.4]
  input  [4:0]  io_in_290, // @[:@6.4]
  input  [4:0]  io_in_291, // @[:@6.4]
  input  [4:0]  io_in_292, // @[:@6.4]
  input  [4:0]  io_in_293, // @[:@6.4]
  input  [4:0]  io_in_294, // @[:@6.4]
  input  [4:0]  io_in_295, // @[:@6.4]
  input  [4:0]  io_in_296, // @[:@6.4]
  input  [4:0]  io_in_297, // @[:@6.4]
  input  [4:0]  io_in_298, // @[:@6.4]
  input  [4:0]  io_in_299, // @[:@6.4]
  input  [4:0]  io_in_300, // @[:@6.4]
  input  [4:0]  io_in_301, // @[:@6.4]
  input  [4:0]  io_in_302, // @[:@6.4]
  input  [4:0]  io_in_303, // @[:@6.4]
  input  [4:0]  io_in_304, // @[:@6.4]
  input  [4:0]  io_in_305, // @[:@6.4]
  input  [4:0]  io_in_306, // @[:@6.4]
  input  [4:0]  io_in_307, // @[:@6.4]
  input  [4:0]  io_in_308, // @[:@6.4]
  input  [4:0]  io_in_309, // @[:@6.4]
  input  [4:0]  io_in_310, // @[:@6.4]
  input  [4:0]  io_in_311, // @[:@6.4]
  input  [4:0]  io_in_312, // @[:@6.4]
  input  [4:0]  io_in_313, // @[:@6.4]
  input  [4:0]  io_in_314, // @[:@6.4]
  input  [4:0]  io_in_315, // @[:@6.4]
  input  [4:0]  io_in_316, // @[:@6.4]
  input  [4:0]  io_in_317, // @[:@6.4]
  input  [4:0]  io_in_318, // @[:@6.4]
  input  [4:0]  io_in_319, // @[:@6.4]
  input  [4:0]  io_in_320, // @[:@6.4]
  input  [4:0]  io_in_321, // @[:@6.4]
  input  [4:0]  io_in_322, // @[:@6.4]
  input  [4:0]  io_in_323, // @[:@6.4]
  input  [4:0]  io_in_324, // @[:@6.4]
  input  [4:0]  io_in_325, // @[:@6.4]
  input  [4:0]  io_in_326, // @[:@6.4]
  input  [4:0]  io_in_327, // @[:@6.4]
  input  [4:0]  io_in_328, // @[:@6.4]
  input  [4:0]  io_in_329, // @[:@6.4]
  input  [4:0]  io_in_330, // @[:@6.4]
  input  [4:0]  io_in_331, // @[:@6.4]
  input  [4:0]  io_in_332, // @[:@6.4]
  input  [4:0]  io_in_333, // @[:@6.4]
  input  [4:0]  io_in_334, // @[:@6.4]
  input  [4:0]  io_in_335, // @[:@6.4]
  input  [4:0]  io_in_336, // @[:@6.4]
  input  [4:0]  io_in_337, // @[:@6.4]
  input  [4:0]  io_in_338, // @[:@6.4]
  input  [4:0]  io_in_339, // @[:@6.4]
  input  [4:0]  io_in_340, // @[:@6.4]
  input  [4:0]  io_in_341, // @[:@6.4]
  input  [4:0]  io_in_342, // @[:@6.4]
  input  [4:0]  io_in_343, // @[:@6.4]
  input  [4:0]  io_in_344, // @[:@6.4]
  input  [4:0]  io_in_345, // @[:@6.4]
  input  [4:0]  io_in_346, // @[:@6.4]
  input  [4:0]  io_in_347, // @[:@6.4]
  input  [4:0]  io_in_348, // @[:@6.4]
  input  [4:0]  io_in_349, // @[:@6.4]
  input  [4:0]  io_in_350, // @[:@6.4]
  input  [4:0]  io_in_351, // @[:@6.4]
  input  [4:0]  io_in_352, // @[:@6.4]
  input  [4:0]  io_in_353, // @[:@6.4]
  input  [4:0]  io_in_354, // @[:@6.4]
  input  [4:0]  io_in_355, // @[:@6.4]
  input  [4:0]  io_in_356, // @[:@6.4]
  input  [4:0]  io_in_357, // @[:@6.4]
  input  [4:0]  io_in_358, // @[:@6.4]
  input  [4:0]  io_in_359, // @[:@6.4]
  input  [4:0]  io_in_360, // @[:@6.4]
  input  [4:0]  io_in_361, // @[:@6.4]
  input  [4:0]  io_in_362, // @[:@6.4]
  input  [4:0]  io_in_363, // @[:@6.4]
  input  [4:0]  io_in_364, // @[:@6.4]
  input  [4:0]  io_in_365, // @[:@6.4]
  input  [4:0]  io_in_366, // @[:@6.4]
  input  [4:0]  io_in_367, // @[:@6.4]
  input  [4:0]  io_in_368, // @[:@6.4]
  input  [4:0]  io_in_369, // @[:@6.4]
  input  [4:0]  io_in_370, // @[:@6.4]
  input  [4:0]  io_in_371, // @[:@6.4]
  input  [4:0]  io_in_372, // @[:@6.4]
  input  [4:0]  io_in_373, // @[:@6.4]
  input  [4:0]  io_in_374, // @[:@6.4]
  input  [4:0]  io_in_375, // @[:@6.4]
  input  [4:0]  io_in_376, // @[:@6.4]
  input  [4:0]  io_in_377, // @[:@6.4]
  input  [4:0]  io_in_378, // @[:@6.4]
  input  [4:0]  io_in_379, // @[:@6.4]
  input  [4:0]  io_in_380, // @[:@6.4]
  input  [4:0]  io_in_381, // @[:@6.4]
  input  [4:0]  io_in_382, // @[:@6.4]
  input  [4:0]  io_in_383, // @[:@6.4]
  input  [4:0]  io_in_384, // @[:@6.4]
  input  [4:0]  io_in_385, // @[:@6.4]
  input  [4:0]  io_in_386, // @[:@6.4]
  input  [4:0]  io_in_387, // @[:@6.4]
  input  [4:0]  io_in_388, // @[:@6.4]
  input  [4:0]  io_in_389, // @[:@6.4]
  input  [4:0]  io_in_390, // @[:@6.4]
  input  [4:0]  io_in_391, // @[:@6.4]
  input  [4:0]  io_in_392, // @[:@6.4]
  input  [4:0]  io_in_393, // @[:@6.4]
  input  [4:0]  io_in_394, // @[:@6.4]
  input  [4:0]  io_in_395, // @[:@6.4]
  input  [4:0]  io_in_396, // @[:@6.4]
  input  [4:0]  io_in_397, // @[:@6.4]
  input  [4:0]  io_in_398, // @[:@6.4]
  input  [4:0]  io_in_399, // @[:@6.4]
  input  [4:0]  io_in_400, // @[:@6.4]
  input  [4:0]  io_in_401, // @[:@6.4]
  input  [4:0]  io_in_402, // @[:@6.4]
  input  [4:0]  io_in_403, // @[:@6.4]
  input  [4:0]  io_in_404, // @[:@6.4]
  input  [4:0]  io_in_405, // @[:@6.4]
  input  [4:0]  io_in_406, // @[:@6.4]
  input  [4:0]  io_in_407, // @[:@6.4]
  input  [4:0]  io_in_408, // @[:@6.4]
  input  [4:0]  io_in_409, // @[:@6.4]
  input  [4:0]  io_in_410, // @[:@6.4]
  input  [4:0]  io_in_411, // @[:@6.4]
  input  [4:0]  io_in_412, // @[:@6.4]
  input  [4:0]  io_in_413, // @[:@6.4]
  input  [4:0]  io_in_414, // @[:@6.4]
  input  [4:0]  io_in_415, // @[:@6.4]
  input  [4:0]  io_in_416, // @[:@6.4]
  input  [4:0]  io_in_417, // @[:@6.4]
  input  [4:0]  io_in_418, // @[:@6.4]
  input  [4:0]  io_in_419, // @[:@6.4]
  input  [4:0]  io_in_420, // @[:@6.4]
  input  [4:0]  io_in_421, // @[:@6.4]
  input  [4:0]  io_in_422, // @[:@6.4]
  input  [4:0]  io_in_423, // @[:@6.4]
  input  [4:0]  io_in_424, // @[:@6.4]
  input  [4:0]  io_in_425, // @[:@6.4]
  input  [4:0]  io_in_426, // @[:@6.4]
  input  [4:0]  io_in_427, // @[:@6.4]
  input  [4:0]  io_in_428, // @[:@6.4]
  input  [4:0]  io_in_429, // @[:@6.4]
  input  [4:0]  io_in_430, // @[:@6.4]
  input  [4:0]  io_in_431, // @[:@6.4]
  input  [4:0]  io_in_432, // @[:@6.4]
  input  [4:0]  io_in_433, // @[:@6.4]
  input  [4:0]  io_in_434, // @[:@6.4]
  input  [4:0]  io_in_435, // @[:@6.4]
  input  [4:0]  io_in_436, // @[:@6.4]
  input  [4:0]  io_in_437, // @[:@6.4]
  input  [4:0]  io_in_438, // @[:@6.4]
  input  [4:0]  io_in_439, // @[:@6.4]
  input  [4:0]  io_in_440, // @[:@6.4]
  input  [4:0]  io_in_441, // @[:@6.4]
  input  [4:0]  io_in_442, // @[:@6.4]
  input  [4:0]  io_in_443, // @[:@6.4]
  input  [4:0]  io_in_444, // @[:@6.4]
  input  [4:0]  io_in_445, // @[:@6.4]
  input  [4:0]  io_in_446, // @[:@6.4]
  input  [4:0]  io_in_447, // @[:@6.4]
  input  [4:0]  io_in_448, // @[:@6.4]
  input  [4:0]  io_in_449, // @[:@6.4]
  input  [4:0]  io_in_450, // @[:@6.4]
  input  [4:0]  io_in_451, // @[:@6.4]
  input  [4:0]  io_in_452, // @[:@6.4]
  input  [4:0]  io_in_453, // @[:@6.4]
  input  [4:0]  io_in_454, // @[:@6.4]
  input  [4:0]  io_in_455, // @[:@6.4]
  input  [4:0]  io_in_456, // @[:@6.4]
  input  [4:0]  io_in_457, // @[:@6.4]
  input  [4:0]  io_in_458, // @[:@6.4]
  input  [4:0]  io_in_459, // @[:@6.4]
  input  [4:0]  io_in_460, // @[:@6.4]
  input  [4:0]  io_in_461, // @[:@6.4]
  input  [4:0]  io_in_462, // @[:@6.4]
  input  [4:0]  io_in_463, // @[:@6.4]
  input  [4:0]  io_in_464, // @[:@6.4]
  input  [4:0]  io_in_465, // @[:@6.4]
  input  [4:0]  io_in_466, // @[:@6.4]
  input  [4:0]  io_in_467, // @[:@6.4]
  input  [4:0]  io_in_468, // @[:@6.4]
  input  [4:0]  io_in_469, // @[:@6.4]
  input  [4:0]  io_in_470, // @[:@6.4]
  input  [4:0]  io_in_471, // @[:@6.4]
  input  [4:0]  io_in_472, // @[:@6.4]
  input  [4:0]  io_in_473, // @[:@6.4]
  input  [4:0]  io_in_474, // @[:@6.4]
  input  [4:0]  io_in_475, // @[:@6.4]
  input  [4:0]  io_in_476, // @[:@6.4]
  input  [4:0]  io_in_477, // @[:@6.4]
  input  [4:0]  io_in_478, // @[:@6.4]
  input  [4:0]  io_in_479, // @[:@6.4]
  input  [4:0]  io_in_480, // @[:@6.4]
  input  [4:0]  io_in_481, // @[:@6.4]
  input  [4:0]  io_in_482, // @[:@6.4]
  input  [4:0]  io_in_483, // @[:@6.4]
  input  [4:0]  io_in_484, // @[:@6.4]
  input  [4:0]  io_in_485, // @[:@6.4]
  input  [4:0]  io_in_486, // @[:@6.4]
  input  [4:0]  io_in_487, // @[:@6.4]
  input  [4:0]  io_in_488, // @[:@6.4]
  input  [4:0]  io_in_489, // @[:@6.4]
  input  [4:0]  io_in_490, // @[:@6.4]
  input  [4:0]  io_in_491, // @[:@6.4]
  input  [4:0]  io_in_492, // @[:@6.4]
  input  [4:0]  io_in_493, // @[:@6.4]
  input  [4:0]  io_in_494, // @[:@6.4]
  input  [4:0]  io_in_495, // @[:@6.4]
  input  [4:0]  io_in_496, // @[:@6.4]
  input  [4:0]  io_in_497, // @[:@6.4]
  input  [4:0]  io_in_498, // @[:@6.4]
  input  [4:0]  io_in_499, // @[:@6.4]
  input  [4:0]  io_in_500, // @[:@6.4]
  input  [4:0]  io_in_501, // @[:@6.4]
  input  [4:0]  io_in_502, // @[:@6.4]
  input  [4:0]  io_in_503, // @[:@6.4]
  input  [4:0]  io_in_504, // @[:@6.4]
  input  [4:0]  io_in_505, // @[:@6.4]
  input  [4:0]  io_in_506, // @[:@6.4]
  input  [4:0]  io_in_507, // @[:@6.4]
  input  [4:0]  io_in_508, // @[:@6.4]
  input  [4:0]  io_in_509, // @[:@6.4]
  input  [4:0]  io_in_510, // @[:@6.4]
  input  [4:0]  io_in_511, // @[:@6.4]
  input  [4:0]  io_in_512, // @[:@6.4]
  input  [4:0]  io_in_513, // @[:@6.4]
  input  [4:0]  io_in_514, // @[:@6.4]
  input  [4:0]  io_in_515, // @[:@6.4]
  input  [4:0]  io_in_516, // @[:@6.4]
  input  [4:0]  io_in_517, // @[:@6.4]
  input  [4:0]  io_in_518, // @[:@6.4]
  input  [4:0]  io_in_519, // @[:@6.4]
  input  [4:0]  io_in_520, // @[:@6.4]
  input  [4:0]  io_in_521, // @[:@6.4]
  input  [4:0]  io_in_522, // @[:@6.4]
  input  [4:0]  io_in_523, // @[:@6.4]
  input  [4:0]  io_in_524, // @[:@6.4]
  input  [4:0]  io_in_525, // @[:@6.4]
  input  [4:0]  io_in_526, // @[:@6.4]
  input  [4:0]  io_in_527, // @[:@6.4]
  input  [4:0]  io_in_528, // @[:@6.4]
  input  [4:0]  io_in_529, // @[:@6.4]
  input  [4:0]  io_in_530, // @[:@6.4]
  input  [4:0]  io_in_531, // @[:@6.4]
  input  [4:0]  io_in_532, // @[:@6.4]
  input  [4:0]  io_in_533, // @[:@6.4]
  input  [4:0]  io_in_534, // @[:@6.4]
  input  [4:0]  io_in_535, // @[:@6.4]
  input  [4:0]  io_in_536, // @[:@6.4]
  input  [4:0]  io_in_537, // @[:@6.4]
  input  [4:0]  io_in_538, // @[:@6.4]
  input  [4:0]  io_in_539, // @[:@6.4]
  input  [4:0]  io_in_540, // @[:@6.4]
  input  [4:0]  io_in_541, // @[:@6.4]
  input  [4:0]  io_in_542, // @[:@6.4]
  input  [4:0]  io_in_543, // @[:@6.4]
  input  [4:0]  io_in_544, // @[:@6.4]
  input  [4:0]  io_in_545, // @[:@6.4]
  input  [4:0]  io_in_546, // @[:@6.4]
  input  [4:0]  io_in_547, // @[:@6.4]
  input  [4:0]  io_in_548, // @[:@6.4]
  input  [4:0]  io_in_549, // @[:@6.4]
  input  [4:0]  io_in_550, // @[:@6.4]
  input  [4:0]  io_in_551, // @[:@6.4]
  input  [4:0]  io_in_552, // @[:@6.4]
  input  [4:0]  io_in_553, // @[:@6.4]
  input  [4:0]  io_in_554, // @[:@6.4]
  input  [4:0]  io_in_555, // @[:@6.4]
  input  [4:0]  io_in_556, // @[:@6.4]
  input  [4:0]  io_in_557, // @[:@6.4]
  input  [4:0]  io_in_558, // @[:@6.4]
  input  [4:0]  io_in_559, // @[:@6.4]
  input  [4:0]  io_in_560, // @[:@6.4]
  input  [4:0]  io_in_561, // @[:@6.4]
  input  [4:0]  io_in_562, // @[:@6.4]
  input  [4:0]  io_in_563, // @[:@6.4]
  input  [4:0]  io_in_564, // @[:@6.4]
  input  [4:0]  io_in_565, // @[:@6.4]
  input  [4:0]  io_in_566, // @[:@6.4]
  input  [4:0]  io_in_567, // @[:@6.4]
  input  [4:0]  io_in_568, // @[:@6.4]
  input  [4:0]  io_in_569, // @[:@6.4]
  input  [4:0]  io_in_570, // @[:@6.4]
  input  [4:0]  io_in_571, // @[:@6.4]
  input  [4:0]  io_in_572, // @[:@6.4]
  input  [4:0]  io_in_573, // @[:@6.4]
  input  [4:0]  io_in_574, // @[:@6.4]
  input  [4:0]  io_in_575, // @[:@6.4]
  input  [4:0]  io_in_576, // @[:@6.4]
  input  [4:0]  io_in_577, // @[:@6.4]
  input  [4:0]  io_in_578, // @[:@6.4]
  input  [4:0]  io_in_579, // @[:@6.4]
  input  [4:0]  io_in_580, // @[:@6.4]
  input  [4:0]  io_in_581, // @[:@6.4]
  input  [4:0]  io_in_582, // @[:@6.4]
  input  [4:0]  io_in_583, // @[:@6.4]
  input  [4:0]  io_in_584, // @[:@6.4]
  input  [4:0]  io_in_585, // @[:@6.4]
  input  [4:0]  io_in_586, // @[:@6.4]
  input  [4:0]  io_in_587, // @[:@6.4]
  input  [4:0]  io_in_588, // @[:@6.4]
  input  [4:0]  io_in_589, // @[:@6.4]
  input  [4:0]  io_in_590, // @[:@6.4]
  input  [4:0]  io_in_591, // @[:@6.4]
  input  [4:0]  io_in_592, // @[:@6.4]
  input  [4:0]  io_in_593, // @[:@6.4]
  input  [4:0]  io_in_594, // @[:@6.4]
  input  [4:0]  io_in_595, // @[:@6.4]
  input  [4:0]  io_in_596, // @[:@6.4]
  input  [4:0]  io_in_597, // @[:@6.4]
  input  [4:0]  io_in_598, // @[:@6.4]
  input  [4:0]  io_in_599, // @[:@6.4]
  input  [4:0]  io_in_600, // @[:@6.4]
  input  [4:0]  io_in_601, // @[:@6.4]
  input  [4:0]  io_in_602, // @[:@6.4]
  input  [4:0]  io_in_603, // @[:@6.4]
  input  [4:0]  io_in_604, // @[:@6.4]
  input  [4:0]  io_in_605, // @[:@6.4]
  input  [4:0]  io_in_606, // @[:@6.4]
  input  [4:0]  io_in_607, // @[:@6.4]
  input  [4:0]  io_in_608, // @[:@6.4]
  input  [4:0]  io_in_609, // @[:@6.4]
  input  [4:0]  io_in_610, // @[:@6.4]
  input  [4:0]  io_in_611, // @[:@6.4]
  input  [4:0]  io_in_612, // @[:@6.4]
  input  [4:0]  io_in_613, // @[:@6.4]
  input  [4:0]  io_in_614, // @[:@6.4]
  input  [4:0]  io_in_615, // @[:@6.4]
  input  [4:0]  io_in_616, // @[:@6.4]
  input  [4:0]  io_in_617, // @[:@6.4]
  input  [4:0]  io_in_618, // @[:@6.4]
  input  [4:0]  io_in_619, // @[:@6.4]
  input  [4:0]  io_in_620, // @[:@6.4]
  input  [4:0]  io_in_621, // @[:@6.4]
  input  [4:0]  io_in_622, // @[:@6.4]
  input  [4:0]  io_in_623, // @[:@6.4]
  input  [4:0]  io_in_624, // @[:@6.4]
  input  [4:0]  io_in_625, // @[:@6.4]
  input  [4:0]  io_in_626, // @[:@6.4]
  input  [4:0]  io_in_627, // @[:@6.4]
  input  [4:0]  io_in_628, // @[:@6.4]
  input  [4:0]  io_in_629, // @[:@6.4]
  input  [4:0]  io_in_630, // @[:@6.4]
  input  [4:0]  io_in_631, // @[:@6.4]
  input  [4:0]  io_in_632, // @[:@6.4]
  input  [4:0]  io_in_633, // @[:@6.4]
  input  [4:0]  io_in_634, // @[:@6.4]
  input  [4:0]  io_in_635, // @[:@6.4]
  input  [4:0]  io_in_636, // @[:@6.4]
  input  [4:0]  io_in_637, // @[:@6.4]
  input  [4:0]  io_in_638, // @[:@6.4]
  input  [4:0]  io_in_639, // @[:@6.4]
  input  [4:0]  io_in_640, // @[:@6.4]
  input  [4:0]  io_in_641, // @[:@6.4]
  input  [4:0]  io_in_642, // @[:@6.4]
  input  [4:0]  io_in_643, // @[:@6.4]
  input  [4:0]  io_in_644, // @[:@6.4]
  input  [4:0]  io_in_645, // @[:@6.4]
  input  [4:0]  io_in_646, // @[:@6.4]
  input  [4:0]  io_in_647, // @[:@6.4]
  input  [4:0]  io_in_648, // @[:@6.4]
  input  [4:0]  io_in_649, // @[:@6.4]
  input  [4:0]  io_in_650, // @[:@6.4]
  input  [4:0]  io_in_651, // @[:@6.4]
  input  [4:0]  io_in_652, // @[:@6.4]
  input  [4:0]  io_in_653, // @[:@6.4]
  input  [4:0]  io_in_654, // @[:@6.4]
  input  [4:0]  io_in_655, // @[:@6.4]
  input  [4:0]  io_in_656, // @[:@6.4]
  input  [4:0]  io_in_657, // @[:@6.4]
  input  [4:0]  io_in_658, // @[:@6.4]
  input  [4:0]  io_in_659, // @[:@6.4]
  input  [4:0]  io_in_660, // @[:@6.4]
  input  [4:0]  io_in_661, // @[:@6.4]
  input  [4:0]  io_in_662, // @[:@6.4]
  input  [4:0]  io_in_663, // @[:@6.4]
  input  [4:0]  io_in_664, // @[:@6.4]
  input  [4:0]  io_in_665, // @[:@6.4]
  input  [4:0]  io_in_666, // @[:@6.4]
  input  [4:0]  io_in_667, // @[:@6.4]
  input  [4:0]  io_in_668, // @[:@6.4]
  input  [4:0]  io_in_669, // @[:@6.4]
  input  [4:0]  io_in_670, // @[:@6.4]
  input  [4:0]  io_in_671, // @[:@6.4]
  input  [4:0]  io_in_672, // @[:@6.4]
  input  [4:0]  io_in_673, // @[:@6.4]
  input  [4:0]  io_in_674, // @[:@6.4]
  input  [4:0]  io_in_675, // @[:@6.4]
  input  [4:0]  io_in_676, // @[:@6.4]
  input  [4:0]  io_in_677, // @[:@6.4]
  input  [4:0]  io_in_678, // @[:@6.4]
  input  [4:0]  io_in_679, // @[:@6.4]
  input  [4:0]  io_in_680, // @[:@6.4]
  input  [4:0]  io_in_681, // @[:@6.4]
  input  [4:0]  io_in_682, // @[:@6.4]
  input  [4:0]  io_in_683, // @[:@6.4]
  input  [4:0]  io_in_684, // @[:@6.4]
  input  [4:0]  io_in_685, // @[:@6.4]
  input  [4:0]  io_in_686, // @[:@6.4]
  input  [4:0]  io_in_687, // @[:@6.4]
  input  [4:0]  io_in_688, // @[:@6.4]
  input  [4:0]  io_in_689, // @[:@6.4]
  input  [4:0]  io_in_690, // @[:@6.4]
  input  [4:0]  io_in_691, // @[:@6.4]
  input  [4:0]  io_in_692, // @[:@6.4]
  input  [4:0]  io_in_693, // @[:@6.4]
  input  [4:0]  io_in_694, // @[:@6.4]
  input  [4:0]  io_in_695, // @[:@6.4]
  input  [4:0]  io_in_696, // @[:@6.4]
  input  [4:0]  io_in_697, // @[:@6.4]
  input  [4:0]  io_in_698, // @[:@6.4]
  input  [4:0]  io_in_699, // @[:@6.4]
  input  [4:0]  io_in_700, // @[:@6.4]
  input  [4:0]  io_in_701, // @[:@6.4]
  input  [4:0]  io_in_702, // @[:@6.4]
  input  [4:0]  io_in_703, // @[:@6.4]
  input  [4:0]  io_in_704, // @[:@6.4]
  input  [4:0]  io_in_705, // @[:@6.4]
  input  [4:0]  io_in_706, // @[:@6.4]
  input  [4:0]  io_in_707, // @[:@6.4]
  input  [4:0]  io_in_708, // @[:@6.4]
  input  [4:0]  io_in_709, // @[:@6.4]
  input  [4:0]  io_in_710, // @[:@6.4]
  input  [4:0]  io_in_711, // @[:@6.4]
  input  [4:0]  io_in_712, // @[:@6.4]
  input  [4:0]  io_in_713, // @[:@6.4]
  input  [4:0]  io_in_714, // @[:@6.4]
  input  [4:0]  io_in_715, // @[:@6.4]
  input  [4:0]  io_in_716, // @[:@6.4]
  input  [4:0]  io_in_717, // @[:@6.4]
  input  [4:0]  io_in_718, // @[:@6.4]
  input  [4:0]  io_in_719, // @[:@6.4]
  input  [4:0]  io_in_720, // @[:@6.4]
  input  [4:0]  io_in_721, // @[:@6.4]
  input  [4:0]  io_in_722, // @[:@6.4]
  input  [4:0]  io_in_723, // @[:@6.4]
  input  [4:0]  io_in_724, // @[:@6.4]
  input  [4:0]  io_in_725, // @[:@6.4]
  input  [4:0]  io_in_726, // @[:@6.4]
  input  [4:0]  io_in_727, // @[:@6.4]
  input  [4:0]  io_in_728, // @[:@6.4]
  input  [4:0]  io_in_729, // @[:@6.4]
  input  [4:0]  io_in_730, // @[:@6.4]
  input  [4:0]  io_in_731, // @[:@6.4]
  input  [4:0]  io_in_732, // @[:@6.4]
  input  [4:0]  io_in_733, // @[:@6.4]
  input  [4:0]  io_in_734, // @[:@6.4]
  input  [4:0]  io_in_735, // @[:@6.4]
  input  [4:0]  io_in_736, // @[:@6.4]
  input  [4:0]  io_in_737, // @[:@6.4]
  input  [4:0]  io_in_738, // @[:@6.4]
  input  [4:0]  io_in_739, // @[:@6.4]
  input  [4:0]  io_in_740, // @[:@6.4]
  input  [4:0]  io_in_741, // @[:@6.4]
  input  [4:0]  io_in_742, // @[:@6.4]
  input  [4:0]  io_in_743, // @[:@6.4]
  input  [4:0]  io_in_744, // @[:@6.4]
  input  [4:0]  io_in_745, // @[:@6.4]
  input  [4:0]  io_in_746, // @[:@6.4]
  input  [4:0]  io_in_747, // @[:@6.4]
  input  [4:0]  io_in_748, // @[:@6.4]
  input  [4:0]  io_in_749, // @[:@6.4]
  input  [4:0]  io_in_750, // @[:@6.4]
  input  [4:0]  io_in_751, // @[:@6.4]
  input  [4:0]  io_in_752, // @[:@6.4]
  input  [4:0]  io_in_753, // @[:@6.4]
  input  [4:0]  io_in_754, // @[:@6.4]
  input  [4:0]  io_in_755, // @[:@6.4]
  input  [4:0]  io_in_756, // @[:@6.4]
  input  [4:0]  io_in_757, // @[:@6.4]
  input  [4:0]  io_in_758, // @[:@6.4]
  input  [4:0]  io_in_759, // @[:@6.4]
  input  [4:0]  io_in_760, // @[:@6.4]
  input  [4:0]  io_in_761, // @[:@6.4]
  input  [4:0]  io_in_762, // @[:@6.4]
  input  [4:0]  io_in_763, // @[:@6.4]
  input  [4:0]  io_in_764, // @[:@6.4]
  input  [4:0]  io_in_765, // @[:@6.4]
  input  [4:0]  io_in_766, // @[:@6.4]
  input  [4:0]  io_in_767, // @[:@6.4]
  input  [4:0]  io_in_768, // @[:@6.4]
  input  [4:0]  io_in_769, // @[:@6.4]
  input  [4:0]  io_in_770, // @[:@6.4]
  input  [4:0]  io_in_771, // @[:@6.4]
  input  [4:0]  io_in_772, // @[:@6.4]
  input  [4:0]  io_in_773, // @[:@6.4]
  input  [4:0]  io_in_774, // @[:@6.4]
  input  [4:0]  io_in_775, // @[:@6.4]
  input  [4:0]  io_in_776, // @[:@6.4]
  input  [4:0]  io_in_777, // @[:@6.4]
  input  [4:0]  io_in_778, // @[:@6.4]
  input  [4:0]  io_in_779, // @[:@6.4]
  input  [4:0]  io_in_780, // @[:@6.4]
  input  [4:0]  io_in_781, // @[:@6.4]
  input  [4:0]  io_in_782, // @[:@6.4]
  input  [4:0]  io_in_783, // @[:@6.4]
  output [10:0] io_out_0, // @[:@6.4]
  output [10:0] io_out_1, // @[:@6.4]
  output [10:0] io_out_2, // @[:@6.4]
  output [10:0] io_out_3, // @[:@6.4]
  output [10:0] io_out_4, // @[:@6.4]
  output [10:0] io_out_5, // @[:@6.4]
  output [10:0] io_out_6, // @[:@6.4]
  output [10:0] io_out_7, // @[:@6.4]
  output [10:0] io_out_8, // @[:@6.4]
  output [10:0] io_out_9, // @[:@6.4]
  output [10:0] io_out_10, // @[:@6.4]
  output [10:0] io_out_11, // @[:@6.4]
  output [10:0] io_out_12, // @[:@6.4]
  output [10:0] io_out_13, // @[:@6.4]
  output [10:0] io_out_14, // @[:@6.4]
  output [10:0] io_out_15 // @[:@6.4]
);
  wire [5:0] _T_54270; // @[Modules.scala 37:46:@17.4]
  wire [4:0] _T_54271; // @[Modules.scala 37:46:@18.4]
  wire [4:0] _T_54272; // @[Modules.scala 37:46:@19.4]
  wire [5:0] _T_54274; // @[Modules.scala 37:46:@22.4]
  wire [4:0] _T_54275; // @[Modules.scala 37:46:@23.4]
  wire [4:0] _T_54276; // @[Modules.scala 37:46:@24.4]
  wire [5:0] _T_54278; // @[Modules.scala 37:46:@31.4]
  wire [4:0] _T_54279; // @[Modules.scala 37:46:@32.4]
  wire [4:0] _T_54280; // @[Modules.scala 37:46:@33.4]
  wire [5:0] _T_54290; // @[Modules.scala 37:46:@44.4]
  wire [4:0] _T_54291; // @[Modules.scala 37:46:@45.4]
  wire [4:0] _T_54292; // @[Modules.scala 37:46:@46.4]
  wire [5:0] _T_54300; // @[Modules.scala 37:46:@60.4]
  wire [4:0] _T_54301; // @[Modules.scala 37:46:@61.4]
  wire [4:0] _T_54302; // @[Modules.scala 37:46:@62.4]
  wire [5:0] _T_54305; // @[Modules.scala 37:46:@68.4]
  wire [4:0] _T_54306; // @[Modules.scala 37:46:@69.4]
  wire [4:0] _T_54307; // @[Modules.scala 37:46:@70.4]
  wire [5:0] _T_54308; // @[Modules.scala 37:46:@72.4]
  wire [4:0] _T_54309; // @[Modules.scala 37:46:@73.4]
  wire [4:0] _T_54310; // @[Modules.scala 37:46:@74.4]
  wire [5:0] _T_54311; // @[Modules.scala 37:46:@77.4]
  wire [4:0] _T_54312; // @[Modules.scala 37:46:@78.4]
  wire [4:0] _T_54313; // @[Modules.scala 37:46:@79.4]
  wire [5:0] _T_54314; // @[Modules.scala 37:46:@82.4]
  wire [4:0] _T_54315; // @[Modules.scala 37:46:@83.4]
  wire [4:0] _T_54316; // @[Modules.scala 37:46:@84.4]
  wire [5:0] _T_54317; // @[Modules.scala 37:46:@86.4]
  wire [4:0] _T_54318; // @[Modules.scala 37:46:@87.4]
  wire [4:0] _T_54319; // @[Modules.scala 37:46:@88.4]
  wire [5:0] _T_54320; // @[Modules.scala 37:46:@90.4]
  wire [4:0] _T_54321; // @[Modules.scala 37:46:@91.4]
  wire [4:0] _T_54322; // @[Modules.scala 37:46:@92.4]
  wire [5:0] _T_54323; // @[Modules.scala 37:46:@94.4]
  wire [4:0] _T_54324; // @[Modules.scala 37:46:@95.4]
  wire [4:0] _T_54325; // @[Modules.scala 37:46:@96.4]
  wire [5:0] _T_54326; // @[Modules.scala 37:46:@98.4]
  wire [4:0] _T_54327; // @[Modules.scala 37:46:@99.4]
  wire [4:0] _T_54328; // @[Modules.scala 37:46:@100.4]
  wire [5:0] _T_54329; // @[Modules.scala 37:46:@103.4]
  wire [4:0] _T_54330; // @[Modules.scala 37:46:@104.4]
  wire [4:0] _T_54331; // @[Modules.scala 37:46:@105.4]
  wire [5:0] _T_54333; // @[Modules.scala 37:46:@110.4]
  wire [4:0] _T_54334; // @[Modules.scala 37:46:@111.4]
  wire [4:0] _T_54335; // @[Modules.scala 37:46:@112.4]
  wire [5:0] _T_54340; // @[Modules.scala 37:46:@120.4]
  wire [4:0] _T_54341; // @[Modules.scala 37:46:@121.4]
  wire [4:0] _T_54342; // @[Modules.scala 37:46:@122.4]
  wire [5:0] _T_54343; // @[Modules.scala 37:46:@124.4]
  wire [4:0] _T_54344; // @[Modules.scala 37:46:@125.4]
  wire [4:0] _T_54345; // @[Modules.scala 37:46:@126.4]
  wire [5:0] _T_54347; // @[Modules.scala 37:46:@130.4]
  wire [4:0] _T_54348; // @[Modules.scala 37:46:@131.4]
  wire [4:0] _T_54349; // @[Modules.scala 37:46:@132.4]
  wire [5:0] _T_54351; // @[Modules.scala 37:46:@136.4]
  wire [4:0] _T_54352; // @[Modules.scala 37:46:@137.4]
  wire [4:0] _T_54353; // @[Modules.scala 37:46:@138.4]
  wire [5:0] _T_54354; // @[Modules.scala 37:46:@140.4]
  wire [4:0] _T_54355; // @[Modules.scala 37:46:@141.4]
  wire [4:0] _T_54356; // @[Modules.scala 37:46:@142.4]
  wire [5:0] _T_54363; // @[Modules.scala 37:46:@150.4]
  wire [4:0] _T_54364; // @[Modules.scala 37:46:@151.4]
  wire [4:0] _T_54365; // @[Modules.scala 37:46:@152.4]
  wire [5:0] _T_54374; // @[Modules.scala 37:46:@165.4]
  wire [4:0] _T_54375; // @[Modules.scala 37:46:@166.4]
  wire [4:0] _T_54376; // @[Modules.scala 37:46:@167.4]
  wire [5:0] _T_54383; // @[Modules.scala 37:46:@180.4]
  wire [4:0] _T_54384; // @[Modules.scala 37:46:@181.4]
  wire [4:0] _T_54385; // @[Modules.scala 37:46:@182.4]
  wire [5:0] _T_54433; // @[Modules.scala 37:46:@236.4]
  wire [4:0] _T_54434; // @[Modules.scala 37:46:@237.4]
  wire [4:0] _T_54435; // @[Modules.scala 37:46:@238.4]
  wire [5:0] _T_54436; // @[Modules.scala 37:46:@240.4]
  wire [4:0] _T_54437; // @[Modules.scala 37:46:@241.4]
  wire [4:0] _T_54438; // @[Modules.scala 37:46:@242.4]
  wire [5:0] _T_54442; // @[Modules.scala 37:46:@248.4]
  wire [4:0] _T_54443; // @[Modules.scala 37:46:@249.4]
  wire [4:0] _T_54444; // @[Modules.scala 37:46:@250.4]
  wire [5:0] _T_54448; // @[Modules.scala 37:46:@258.4]
  wire [4:0] _T_54449; // @[Modules.scala 37:46:@259.4]
  wire [4:0] _T_54450; // @[Modules.scala 37:46:@260.4]
  wire [5:0] _T_54451; // @[Modules.scala 37:46:@262.4]
  wire [4:0] _T_54452; // @[Modules.scala 37:46:@263.4]
  wire [4:0] _T_54453; // @[Modules.scala 37:46:@264.4]
  wire [5:0] _T_54454; // @[Modules.scala 37:46:@266.4]
  wire [4:0] _T_54455; // @[Modules.scala 37:46:@267.4]
  wire [4:0] _T_54456; // @[Modules.scala 37:46:@268.4]
  wire [5:0] _T_54457; // @[Modules.scala 37:46:@270.4]
  wire [4:0] _T_54458; // @[Modules.scala 37:46:@271.4]
  wire [4:0] _T_54459; // @[Modules.scala 37:46:@272.4]
  wire [5:0] _T_54460; // @[Modules.scala 37:46:@274.4]
  wire [4:0] _T_54461; // @[Modules.scala 37:46:@275.4]
  wire [4:0] _T_54462; // @[Modules.scala 37:46:@276.4]
  wire [5:0] _T_54463; // @[Modules.scala 37:46:@278.4]
  wire [4:0] _T_54464; // @[Modules.scala 37:46:@279.4]
  wire [4:0] _T_54465; // @[Modules.scala 37:46:@280.4]
  wire [5:0] _T_54466; // @[Modules.scala 37:46:@282.4]
  wire [4:0] _T_54467; // @[Modules.scala 37:46:@283.4]
  wire [4:0] _T_54468; // @[Modules.scala 37:46:@284.4]
  wire [5:0] _T_54469; // @[Modules.scala 37:46:@286.4]
  wire [4:0] _T_54470; // @[Modules.scala 37:46:@287.4]
  wire [4:0] _T_54471; // @[Modules.scala 37:46:@288.4]
  wire [5:0] _T_54472; // @[Modules.scala 37:46:@290.4]
  wire [4:0] _T_54473; // @[Modules.scala 37:46:@291.4]
  wire [4:0] _T_54474; // @[Modules.scala 37:46:@292.4]
  wire [5:0] _T_54478; // @[Modules.scala 37:46:@298.4]
  wire [4:0] _T_54479; // @[Modules.scala 37:46:@299.4]
  wire [4:0] _T_54480; // @[Modules.scala 37:46:@300.4]
  wire [5:0] _T_54481; // @[Modules.scala 37:46:@302.4]
  wire [4:0] _T_54482; // @[Modules.scala 37:46:@303.4]
  wire [4:0] _T_54483; // @[Modules.scala 37:46:@304.4]
  wire [5:0] _T_54484; // @[Modules.scala 37:46:@306.4]
  wire [4:0] _T_54485; // @[Modules.scala 37:46:@307.4]
  wire [4:0] _T_54486; // @[Modules.scala 37:46:@308.4]
  wire [5:0] _T_54487; // @[Modules.scala 37:46:@310.4]
  wire [4:0] _T_54488; // @[Modules.scala 37:46:@311.4]
  wire [4:0] _T_54489; // @[Modules.scala 37:46:@312.4]
  wire [5:0] _T_54490; // @[Modules.scala 37:46:@314.4]
  wire [4:0] _T_54491; // @[Modules.scala 37:46:@315.4]
  wire [4:0] _T_54492; // @[Modules.scala 37:46:@316.4]
  wire [5:0] _T_54493; // @[Modules.scala 37:46:@318.4]
  wire [4:0] _T_54494; // @[Modules.scala 37:46:@319.4]
  wire [4:0] _T_54495; // @[Modules.scala 37:46:@320.4]
  wire [5:0] _T_54496; // @[Modules.scala 37:46:@322.4]
  wire [4:0] _T_54497; // @[Modules.scala 37:46:@323.4]
  wire [4:0] _T_54498; // @[Modules.scala 37:46:@324.4]
  wire [5:0] _T_54499; // @[Modules.scala 37:46:@326.4]
  wire [4:0] _T_54500; // @[Modules.scala 37:46:@327.4]
  wire [4:0] _T_54501; // @[Modules.scala 37:46:@328.4]
  wire [5:0] _T_54502; // @[Modules.scala 37:46:@331.4]
  wire [4:0] _T_54503; // @[Modules.scala 37:46:@332.4]
  wire [4:0] _T_54504; // @[Modules.scala 37:46:@333.4]
  wire [5:0] _T_54507; // @[Modules.scala 37:46:@339.4]
  wire [4:0] _T_54508; // @[Modules.scala 37:46:@340.4]
  wire [4:0] _T_54509; // @[Modules.scala 37:46:@341.4]
  wire [5:0] _T_54510; // @[Modules.scala 37:46:@343.4]
  wire [4:0] _T_54511; // @[Modules.scala 37:46:@344.4]
  wire [4:0] _T_54512; // @[Modules.scala 37:46:@345.4]
  wire [5:0] _T_54513; // @[Modules.scala 37:46:@347.4]
  wire [4:0] _T_54514; // @[Modules.scala 37:46:@348.4]
  wire [4:0] _T_54515; // @[Modules.scala 37:46:@349.4]
  wire [5:0] _T_54516; // @[Modules.scala 37:46:@351.4]
  wire [4:0] _T_54517; // @[Modules.scala 37:46:@352.4]
  wire [4:0] _T_54518; // @[Modules.scala 37:46:@353.4]
  wire [5:0] _T_54519; // @[Modules.scala 37:46:@355.4]
  wire [4:0] _T_54520; // @[Modules.scala 37:46:@356.4]
  wire [4:0] _T_54521; // @[Modules.scala 37:46:@357.4]
  wire [5:0] _T_54522; // @[Modules.scala 37:46:@359.4]
  wire [4:0] _T_54523; // @[Modules.scala 37:46:@360.4]
  wire [4:0] _T_54524; // @[Modules.scala 37:46:@361.4]
  wire [5:0] _T_54525; // @[Modules.scala 37:46:@363.4]
  wire [4:0] _T_54526; // @[Modules.scala 37:46:@364.4]
  wire [4:0] _T_54527; // @[Modules.scala 37:46:@365.4]
  wire [5:0] _T_54528; // @[Modules.scala 37:46:@367.4]
  wire [4:0] _T_54529; // @[Modules.scala 37:46:@368.4]
  wire [4:0] _T_54530; // @[Modules.scala 37:46:@369.4]
  wire [5:0] _T_54531; // @[Modules.scala 37:46:@371.4]
  wire [4:0] _T_54532; // @[Modules.scala 37:46:@372.4]
  wire [4:0] _T_54533; // @[Modules.scala 37:46:@373.4]
  wire [5:0] _T_54534; // @[Modules.scala 37:46:@375.4]
  wire [4:0] _T_54535; // @[Modules.scala 37:46:@376.4]
  wire [4:0] _T_54536; // @[Modules.scala 37:46:@377.4]
  wire [5:0] _T_54538; // @[Modules.scala 37:46:@384.4]
  wire [4:0] _T_54539; // @[Modules.scala 37:46:@385.4]
  wire [4:0] _T_54540; // @[Modules.scala 37:46:@386.4]
  wire [5:0] _T_54541; // @[Modules.scala 37:46:@388.4]
  wire [4:0] _T_54542; // @[Modules.scala 37:46:@389.4]
  wire [4:0] _T_54543; // @[Modules.scala 37:46:@390.4]
  wire [5:0] _T_54544; // @[Modules.scala 37:46:@392.4]
  wire [4:0] _T_54545; // @[Modules.scala 37:46:@393.4]
  wire [4:0] _T_54546; // @[Modules.scala 37:46:@394.4]
  wire [5:0] _T_54547; // @[Modules.scala 37:46:@396.4]
  wire [4:0] _T_54548; // @[Modules.scala 37:46:@397.4]
  wire [4:0] _T_54549; // @[Modules.scala 37:46:@398.4]
  wire [5:0] _T_54550; // @[Modules.scala 37:46:@400.4]
  wire [4:0] _T_54551; // @[Modules.scala 37:46:@401.4]
  wire [4:0] _T_54552; // @[Modules.scala 37:46:@402.4]
  wire [5:0] _T_54553; // @[Modules.scala 37:46:@404.4]
  wire [4:0] _T_54554; // @[Modules.scala 37:46:@405.4]
  wire [4:0] _T_54555; // @[Modules.scala 37:46:@406.4]
  wire [5:0] _T_54558; // @[Modules.scala 37:46:@413.4]
  wire [4:0] _T_54559; // @[Modules.scala 37:46:@414.4]
  wire [4:0] _T_54560; // @[Modules.scala 37:46:@415.4]
  wire [5:0] _T_54562; // @[Modules.scala 37:46:@419.4]
  wire [4:0] _T_54563; // @[Modules.scala 37:46:@420.4]
  wire [4:0] _T_54564; // @[Modules.scala 37:46:@421.4]
  wire [5:0] _T_54565; // @[Modules.scala 37:46:@423.4]
  wire [4:0] _T_54566; // @[Modules.scala 37:46:@424.4]
  wire [4:0] _T_54567; // @[Modules.scala 37:46:@425.4]
  wire [5:0] _T_54568; // @[Modules.scala 37:46:@427.4]
  wire [4:0] _T_54569; // @[Modules.scala 37:46:@428.4]
  wire [4:0] _T_54570; // @[Modules.scala 37:46:@429.4]
  wire [5:0] _T_54571; // @[Modules.scala 37:46:@432.4]
  wire [4:0] _T_54572; // @[Modules.scala 37:46:@433.4]
  wire [4:0] _T_54573; // @[Modules.scala 37:46:@434.4]
  wire [5:0] _T_54574; // @[Modules.scala 37:46:@436.4]
  wire [4:0] _T_54575; // @[Modules.scala 37:46:@437.4]
  wire [4:0] _T_54576; // @[Modules.scala 37:46:@438.4]
  wire [5:0] _T_54577; // @[Modules.scala 37:46:@440.4]
  wire [4:0] _T_54578; // @[Modules.scala 37:46:@441.4]
  wire [4:0] _T_54579; // @[Modules.scala 37:46:@442.4]
  wire [5:0] _T_54585; // @[Modules.scala 37:46:@451.4]
  wire [4:0] _T_54586; // @[Modules.scala 37:46:@452.4]
  wire [4:0] _T_54587; // @[Modules.scala 37:46:@453.4]
  wire [5:0] _T_54588; // @[Modules.scala 37:46:@455.4]
  wire [4:0] _T_54589; // @[Modules.scala 37:46:@456.4]
  wire [4:0] _T_54590; // @[Modules.scala 37:46:@457.4]
  wire [5:0] _T_54591; // @[Modules.scala 37:46:@459.4]
  wire [4:0] _T_54592; // @[Modules.scala 37:46:@460.4]
  wire [4:0] _T_54593; // @[Modules.scala 37:46:@461.4]
  wire [5:0] _T_54594; // @[Modules.scala 37:46:@464.4]
  wire [4:0] _T_54595; // @[Modules.scala 37:46:@465.4]
  wire [4:0] _T_54596; // @[Modules.scala 37:46:@466.4]
  wire [5:0] _T_54598; // @[Modules.scala 37:46:@471.4]
  wire [4:0] _T_54599; // @[Modules.scala 37:46:@472.4]
  wire [4:0] _T_54600; // @[Modules.scala 37:46:@473.4]
  wire [5:0] _T_54606; // @[Modules.scala 37:46:@481.4]
  wire [4:0] _T_54607; // @[Modules.scala 37:46:@482.4]
  wire [4:0] _T_54608; // @[Modules.scala 37:46:@483.4]
  wire [5:0] _T_54609; // @[Modules.scala 37:46:@485.4]
  wire [4:0] _T_54610; // @[Modules.scala 37:46:@486.4]
  wire [4:0] _T_54611; // @[Modules.scala 37:46:@487.4]
  wire [5:0] _T_54612; // @[Modules.scala 37:46:@490.4]
  wire [4:0] _T_54613; // @[Modules.scala 37:46:@491.4]
  wire [4:0] _T_54614; // @[Modules.scala 37:46:@492.4]
  wire [5:0] _T_54615; // @[Modules.scala 37:46:@497.4]
  wire [4:0] _T_54616; // @[Modules.scala 37:46:@498.4]
  wire [4:0] _T_54617; // @[Modules.scala 37:46:@499.4]
  wire [5:0] _T_54618; // @[Modules.scala 37:46:@501.4]
  wire [4:0] _T_54619; // @[Modules.scala 37:46:@502.4]
  wire [4:0] _T_54620; // @[Modules.scala 37:46:@503.4]
  wire [5:0] _T_54634; // @[Modules.scala 37:46:@528.4]
  wire [4:0] _T_54635; // @[Modules.scala 37:46:@529.4]
  wire [4:0] _T_54636; // @[Modules.scala 37:46:@530.4]
  wire [5:0] _T_54638; // @[Modules.scala 37:46:@535.4]
  wire [4:0] _T_54639; // @[Modules.scala 37:46:@536.4]
  wire [4:0] _T_54640; // @[Modules.scala 37:46:@537.4]
  wire [5:0] _T_54646; // @[Modules.scala 37:46:@546.4]
  wire [4:0] _T_54647; // @[Modules.scala 37:46:@547.4]
  wire [4:0] _T_54648; // @[Modules.scala 37:46:@548.4]
  wire [5:0] _T_54649; // @[Modules.scala 37:46:@551.4]
  wire [4:0] _T_54650; // @[Modules.scala 37:46:@552.4]
  wire [4:0] _T_54651; // @[Modules.scala 37:46:@553.4]
  wire [5:0] _T_54652; // @[Modules.scala 37:46:@555.4]
  wire [4:0] _T_54653; // @[Modules.scala 37:46:@556.4]
  wire [4:0] _T_54654; // @[Modules.scala 37:46:@557.4]
  wire [5:0] _T_54657; // @[Modules.scala 37:46:@561.4]
  wire [4:0] _T_54658; // @[Modules.scala 37:46:@562.4]
  wire [4:0] _T_54659; // @[Modules.scala 37:46:@563.4]
  wire [5:0] _T_54660; // @[Modules.scala 37:46:@567.4]
  wire [4:0] _T_54661; // @[Modules.scala 37:46:@568.4]
  wire [4:0] _T_54662; // @[Modules.scala 37:46:@569.4]
  wire [5:0] _T_54672; // @[Modules.scala 37:46:@581.4]
  wire [4:0] _T_54673; // @[Modules.scala 37:46:@582.4]
  wire [4:0] _T_54674; // @[Modules.scala 37:46:@583.4]
  wire [5:0] _T_54675; // @[Modules.scala 37:46:@587.4]
  wire [4:0] _T_54676; // @[Modules.scala 37:46:@588.4]
  wire [4:0] _T_54677; // @[Modules.scala 37:46:@589.4]
  wire [5:0] _T_54685; // @[Modules.scala 37:46:@599.4]
  wire [4:0] _T_54686; // @[Modules.scala 37:46:@600.4]
  wire [4:0] _T_54687; // @[Modules.scala 37:46:@601.4]
  wire [5:0] _T_54688; // @[Modules.scala 37:46:@603.4]
  wire [4:0] _T_54689; // @[Modules.scala 37:46:@604.4]
  wire [4:0] _T_54690; // @[Modules.scala 37:46:@605.4]
  wire [5:0] _T_54691; // @[Modules.scala 37:46:@607.4]
  wire [4:0] _T_54692; // @[Modules.scala 37:46:@608.4]
  wire [4:0] _T_54693; // @[Modules.scala 37:46:@609.4]
  wire [5:0] _T_54695; // @[Modules.scala 37:46:@614.4]
  wire [4:0] _T_54696; // @[Modules.scala 37:46:@615.4]
  wire [4:0] _T_54697; // @[Modules.scala 37:46:@616.4]
  wire [5:0] _T_54698; // @[Modules.scala 37:46:@618.4]
  wire [4:0] _T_54699; // @[Modules.scala 37:46:@619.4]
  wire [4:0] _T_54700; // @[Modules.scala 37:46:@620.4]
  wire [5:0] _T_54701; // @[Modules.scala 37:46:@622.4]
  wire [4:0] _T_54702; // @[Modules.scala 37:46:@623.4]
  wire [4:0] _T_54703; // @[Modules.scala 37:46:@624.4]
  wire [5:0] _T_54706; // @[Modules.scala 37:46:@629.4]
  wire [4:0] _T_54707; // @[Modules.scala 37:46:@630.4]
  wire [4:0] _T_54708; // @[Modules.scala 37:46:@631.4]
  wire [5:0] _T_54709; // @[Modules.scala 37:46:@633.4]
  wire [4:0] _T_54710; // @[Modules.scala 37:46:@634.4]
  wire [4:0] _T_54711; // @[Modules.scala 37:46:@635.4]
  wire [5:0] _T_54712; // @[Modules.scala 37:46:@637.4]
  wire [4:0] _T_54713; // @[Modules.scala 37:46:@638.4]
  wire [4:0] _T_54714; // @[Modules.scala 37:46:@639.4]
  wire [5:0] _T_54715; // @[Modules.scala 37:46:@641.4]
  wire [4:0] _T_54716; // @[Modules.scala 37:46:@642.4]
  wire [4:0] _T_54717; // @[Modules.scala 37:46:@643.4]
  wire [5:0] _T_54718; // @[Modules.scala 37:46:@645.4]
  wire [4:0] _T_54719; // @[Modules.scala 37:46:@646.4]
  wire [4:0] _T_54720; // @[Modules.scala 37:46:@647.4]
  wire [5:0] _T_54721; // @[Modules.scala 37:46:@652.4]
  wire [4:0] _T_54722; // @[Modules.scala 37:46:@653.4]
  wire [4:0] _T_54723; // @[Modules.scala 37:46:@654.4]
  wire [5:0] _T_54724; // @[Modules.scala 37:46:@656.4]
  wire [4:0] _T_54725; // @[Modules.scala 37:46:@657.4]
  wire [4:0] _T_54726; // @[Modules.scala 37:46:@658.4]
  wire [5:0] _T_54727; // @[Modules.scala 37:46:@660.4]
  wire [4:0] _T_54728; // @[Modules.scala 37:46:@661.4]
  wire [4:0] _T_54729; // @[Modules.scala 37:46:@662.4]
  wire [5:0] _T_54730; // @[Modules.scala 37:46:@665.4]
  wire [4:0] _T_54731; // @[Modules.scala 37:46:@666.4]
  wire [4:0] _T_54732; // @[Modules.scala 37:46:@667.4]
  wire [5:0] _T_54733; // @[Modules.scala 37:46:@669.4]
  wire [4:0] _T_54734; // @[Modules.scala 37:46:@670.4]
  wire [4:0] _T_54735; // @[Modules.scala 37:46:@671.4]
  wire [5:0] _T_54736; // @[Modules.scala 37:46:@673.4]
  wire [4:0] _T_54737; // @[Modules.scala 37:46:@674.4]
  wire [4:0] _T_54738; // @[Modules.scala 37:46:@675.4]
  wire [5:0] _T_54739; // @[Modules.scala 37:46:@677.4]
  wire [4:0] _T_54740; // @[Modules.scala 37:46:@678.4]
  wire [4:0] _T_54741; // @[Modules.scala 37:46:@679.4]
  wire [5:0] _T_54742; // @[Modules.scala 37:46:@681.4]
  wire [4:0] _T_54743; // @[Modules.scala 37:46:@682.4]
  wire [4:0] _T_54744; // @[Modules.scala 37:46:@683.4]
  wire [5:0] _T_54745; // @[Modules.scala 37:46:@685.4]
  wire [4:0] _T_54746; // @[Modules.scala 37:46:@686.4]
  wire [4:0] _T_54747; // @[Modules.scala 37:46:@687.4]
  wire [5:0] _T_54749; // @[Modules.scala 37:46:@693.4]
  wire [4:0] _T_54750; // @[Modules.scala 37:46:@694.4]
  wire [4:0] _T_54751; // @[Modules.scala 37:46:@695.4]
  wire [5:0] _T_54752; // @[Modules.scala 37:46:@697.4]
  wire [4:0] _T_54753; // @[Modules.scala 37:46:@698.4]
  wire [4:0] _T_54754; // @[Modules.scala 37:46:@699.4]
  wire [5:0] _T_54759; // @[Modules.scala 37:46:@707.4]
  wire [4:0] _T_54760; // @[Modules.scala 37:46:@708.4]
  wire [4:0] _T_54761; // @[Modules.scala 37:46:@709.4]
  wire [5:0] _T_54762; // @[Modules.scala 37:46:@712.4]
  wire [4:0] _T_54763; // @[Modules.scala 37:46:@713.4]
  wire [4:0] _T_54764; // @[Modules.scala 37:46:@714.4]
  wire [5:0] _T_54765; // @[Modules.scala 37:46:@716.4]
  wire [4:0] _T_54766; // @[Modules.scala 37:46:@717.4]
  wire [4:0] _T_54767; // @[Modules.scala 37:46:@718.4]
  wire [5:0] _T_54774; // @[Modules.scala 37:46:@730.4]
  wire [4:0] _T_54775; // @[Modules.scala 37:46:@731.4]
  wire [4:0] _T_54776; // @[Modules.scala 37:46:@732.4]
  wire [5:0] _T_54778; // @[Modules.scala 37:46:@736.4]
  wire [4:0] _T_54779; // @[Modules.scala 37:46:@737.4]
  wire [4:0] _T_54780; // @[Modules.scala 37:46:@738.4]
  wire [10:0] buffer_0_0; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54781; // @[Modules.scala 65:57:@740.4]
  wire [10:0] _T_54782; // @[Modules.scala 65:57:@741.4]
  wire [10:0] buffer_0_392; // @[Modules.scala 65:57:@742.4]
  wire [10:0] buffer_0_2; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_3; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54784; // @[Modules.scala 65:57:@744.4]
  wire [10:0] _T_54785; // @[Modules.scala 65:57:@745.4]
  wire [10:0] buffer_0_393; // @[Modules.scala 65:57:@746.4]
  wire [10:0] buffer_0_4; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54787; // @[Modules.scala 65:57:@748.4]
  wire [10:0] _T_54788; // @[Modules.scala 65:57:@749.4]
  wire [10:0] buffer_0_394; // @[Modules.scala 65:57:@750.4]
  wire [11:0] _T_54790; // @[Modules.scala 65:57:@752.4]
  wire [10:0] _T_54791; // @[Modules.scala 65:57:@753.4]
  wire [10:0] buffer_0_395; // @[Modules.scala 65:57:@754.4]
  wire [10:0] buffer_0_8; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54793; // @[Modules.scala 65:57:@756.4]
  wire [10:0] _T_54794; // @[Modules.scala 65:57:@757.4]
  wire [10:0] buffer_0_396; // @[Modules.scala 65:57:@758.4]
  wire [10:0] buffer_0_10; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54796; // @[Modules.scala 65:57:@760.4]
  wire [10:0] _T_54797; // @[Modules.scala 65:57:@761.4]
  wire [10:0] buffer_0_397; // @[Modules.scala 65:57:@762.4]
  wire [10:0] buffer_0_12; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54799; // @[Modules.scala 65:57:@764.4]
  wire [10:0] _T_54800; // @[Modules.scala 65:57:@765.4]
  wire [10:0] buffer_0_398; // @[Modules.scala 65:57:@766.4]
  wire [10:0] buffer_0_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54802; // @[Modules.scala 65:57:@768.4]
  wire [10:0] _T_54803; // @[Modules.scala 65:57:@769.4]
  wire [10:0] buffer_0_399; // @[Modules.scala 65:57:@770.4]
  wire [10:0] buffer_0_16; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54805; // @[Modules.scala 65:57:@772.4]
  wire [10:0] _T_54806; // @[Modules.scala 65:57:@773.4]
  wire [10:0] buffer_0_400; // @[Modules.scala 65:57:@774.4]
  wire [10:0] buffer_0_26; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54820; // @[Modules.scala 65:57:@792.4]
  wire [10:0] _T_54821; // @[Modules.scala 65:57:@793.4]
  wire [10:0] buffer_0_405; // @[Modules.scala 65:57:@794.4]
  wire [10:0] buffer_0_28; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54823; // @[Modules.scala 65:57:@796.4]
  wire [10:0] _T_54824; // @[Modules.scala 65:57:@797.4]
  wire [10:0] buffer_0_406; // @[Modules.scala 65:57:@798.4]
  wire [10:0] buffer_0_32; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54829; // @[Modules.scala 65:57:@804.4]
  wire [10:0] _T_54830; // @[Modules.scala 65:57:@805.4]
  wire [10:0] buffer_0_408; // @[Modules.scala 65:57:@806.4]
  wire [10:0] buffer_0_37; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54835; // @[Modules.scala 65:57:@812.4]
  wire [10:0] _T_54836; // @[Modules.scala 65:57:@813.4]
  wire [10:0] buffer_0_410; // @[Modules.scala 65:57:@814.4]
  wire [10:0] buffer_0_38; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_39; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54838; // @[Modules.scala 65:57:@816.4]
  wire [10:0] _T_54839; // @[Modules.scala 65:57:@817.4]
  wire [10:0] buffer_0_411; // @[Modules.scala 65:57:@818.4]
  wire [10:0] buffer_0_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54841; // @[Modules.scala 65:57:@820.4]
  wire [10:0] _T_54842; // @[Modules.scala 65:57:@821.4]
  wire [10:0] buffer_0_412; // @[Modules.scala 65:57:@822.4]
  wire [10:0] buffer_0_42; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54844; // @[Modules.scala 65:57:@824.4]
  wire [10:0] _T_54845; // @[Modules.scala 65:57:@825.4]
  wire [10:0] buffer_0_413; // @[Modules.scala 65:57:@826.4]
  wire [10:0] buffer_0_44; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_45; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54847; // @[Modules.scala 65:57:@828.4]
  wire [10:0] _T_54848; // @[Modules.scala 65:57:@829.4]
  wire [10:0] buffer_0_414; // @[Modules.scala 65:57:@830.4]
  wire [10:0] buffer_0_46; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_47; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54850; // @[Modules.scala 65:57:@832.4]
  wire [10:0] _T_54851; // @[Modules.scala 65:57:@833.4]
  wire [10:0] buffer_0_415; // @[Modules.scala 65:57:@834.4]
  wire [10:0] buffer_0_48; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_49; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54853; // @[Modules.scala 65:57:@836.4]
  wire [10:0] _T_54854; // @[Modules.scala 65:57:@837.4]
  wire [10:0] buffer_0_416; // @[Modules.scala 65:57:@838.4]
  wire [10:0] buffer_0_50; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_51; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54856; // @[Modules.scala 65:57:@840.4]
  wire [10:0] _T_54857; // @[Modules.scala 65:57:@841.4]
  wire [10:0] buffer_0_417; // @[Modules.scala 65:57:@842.4]
  wire [10:0] buffer_0_52; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_53; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54859; // @[Modules.scala 65:57:@844.4]
  wire [10:0] _T_54860; // @[Modules.scala 65:57:@845.4]
  wire [10:0] buffer_0_418; // @[Modules.scala 65:57:@846.4]
  wire [10:0] buffer_0_54; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54862; // @[Modules.scala 65:57:@848.4]
  wire [10:0] _T_54863; // @[Modules.scala 65:57:@849.4]
  wire [10:0] buffer_0_419; // @[Modules.scala 65:57:@850.4]
  wire [10:0] buffer_0_56; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54865; // @[Modules.scala 65:57:@852.4]
  wire [10:0] _T_54866; // @[Modules.scala 65:57:@853.4]
  wire [10:0] buffer_0_420; // @[Modules.scala 65:57:@854.4]
  wire [10:0] buffer_0_58; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_59; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54868; // @[Modules.scala 65:57:@856.4]
  wire [10:0] _T_54869; // @[Modules.scala 65:57:@857.4]
  wire [10:0] buffer_0_421; // @[Modules.scala 65:57:@858.4]
  wire [10:0] buffer_0_64; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_65; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54877; // @[Modules.scala 65:57:@868.4]
  wire [10:0] _T_54878; // @[Modules.scala 65:57:@869.4]
  wire [10:0] buffer_0_424; // @[Modules.scala 65:57:@870.4]
  wire [10:0] buffer_0_66; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_67; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54880; // @[Modules.scala 65:57:@872.4]
  wire [10:0] _T_54881; // @[Modules.scala 65:57:@873.4]
  wire [10:0] buffer_0_425; // @[Modules.scala 65:57:@874.4]
  wire [10:0] buffer_0_68; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54883; // @[Modules.scala 65:57:@876.4]
  wire [10:0] _T_54884; // @[Modules.scala 65:57:@877.4]
  wire [10:0] buffer_0_426; // @[Modules.scala 65:57:@878.4]
  wire [10:0] buffer_0_70; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54886; // @[Modules.scala 65:57:@880.4]
  wire [10:0] _T_54887; // @[Modules.scala 65:57:@881.4]
  wire [10:0] buffer_0_427; // @[Modules.scala 65:57:@882.4]
  wire [10:0] buffer_0_72; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54889; // @[Modules.scala 65:57:@884.4]
  wire [10:0] _T_54890; // @[Modules.scala 65:57:@885.4]
  wire [10:0] buffer_0_428; // @[Modules.scala 65:57:@886.4]
  wire [10:0] buffer_0_74; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54892; // @[Modules.scala 65:57:@888.4]
  wire [10:0] _T_54893; // @[Modules.scala 65:57:@889.4]
  wire [10:0] buffer_0_429; // @[Modules.scala 65:57:@890.4]
  wire [10:0] buffer_0_81; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54901; // @[Modules.scala 65:57:@900.4]
  wire [10:0] _T_54902; // @[Modules.scala 65:57:@901.4]
  wire [10:0] buffer_0_432; // @[Modules.scala 65:57:@902.4]
  wire [10:0] buffer_0_82; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54904; // @[Modules.scala 65:57:@904.4]
  wire [10:0] _T_54905; // @[Modules.scala 65:57:@905.4]
  wire [10:0] buffer_0_433; // @[Modules.scala 65:57:@906.4]
  wire [10:0] buffer_0_86; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54910; // @[Modules.scala 65:57:@912.4]
  wire [10:0] _T_54911; // @[Modules.scala 65:57:@913.4]
  wire [10:0] buffer_0_435; // @[Modules.scala 65:57:@914.4]
  wire [10:0] buffer_0_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54919; // @[Modules.scala 65:57:@924.4]
  wire [10:0] _T_54920; // @[Modules.scala 65:57:@925.4]
  wire [10:0] buffer_0_438; // @[Modules.scala 65:57:@926.4]
  wire [10:0] buffer_0_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54922; // @[Modules.scala 65:57:@928.4]
  wire [10:0] _T_54923; // @[Modules.scala 65:57:@929.4]
  wire [10:0] buffer_0_439; // @[Modules.scala 65:57:@930.4]
  wire [10:0] buffer_0_98; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54928; // @[Modules.scala 65:57:@936.4]
  wire [10:0] _T_54929; // @[Modules.scala 65:57:@937.4]
  wire [10:0] buffer_0_441; // @[Modules.scala 65:57:@938.4]
  wire [10:0] buffer_0_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54934; // @[Modules.scala 65:57:@944.4]
  wire [10:0] _T_54935; // @[Modules.scala 65:57:@945.4]
  wire [10:0] buffer_0_443; // @[Modules.scala 65:57:@946.4]
  wire [10:0] buffer_0_104; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54937; // @[Modules.scala 65:57:@948.4]
  wire [10:0] _T_54938; // @[Modules.scala 65:57:@949.4]
  wire [10:0] buffer_0_444; // @[Modules.scala 65:57:@950.4]
  wire [10:0] buffer_0_106; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54940; // @[Modules.scala 65:57:@952.4]
  wire [10:0] _T_54941; // @[Modules.scala 65:57:@953.4]
  wire [10:0] buffer_0_445; // @[Modules.scala 65:57:@954.4]
  wire [10:0] buffer_0_118; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54958; // @[Modules.scala 65:57:@976.4]
  wire [10:0] _T_54959; // @[Modules.scala 65:57:@977.4]
  wire [10:0] buffer_0_451; // @[Modules.scala 65:57:@978.4]
  wire [10:0] buffer_0_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54976; // @[Modules.scala 65:57:@1000.4]
  wire [10:0] _T_54977; // @[Modules.scala 65:57:@1001.4]
  wire [10:0] buffer_0_457; // @[Modules.scala 65:57:@1002.4]
  wire [10:0] buffer_0_144; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_54997; // @[Modules.scala 65:57:@1028.4]
  wire [10:0] _T_54998; // @[Modules.scala 65:57:@1029.4]
  wire [10:0] buffer_0_464; // @[Modules.scala 65:57:@1030.4]
  wire [10:0] buffer_0_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55015; // @[Modules.scala 65:57:@1052.4]
  wire [10:0] _T_55016; // @[Modules.scala 65:57:@1053.4]
  wire [10:0] buffer_0_470; // @[Modules.scala 65:57:@1054.4]
  wire [10:0] buffer_0_158; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_159; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55018; // @[Modules.scala 65:57:@1056.4]
  wire [10:0] _T_55019; // @[Modules.scala 65:57:@1057.4]
  wire [10:0] buffer_0_471; // @[Modules.scala 65:57:@1058.4]
  wire [10:0] buffer_0_162; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55024; // @[Modules.scala 65:57:@1064.4]
  wire [10:0] _T_55025; // @[Modules.scala 65:57:@1065.4]
  wire [10:0] buffer_0_473; // @[Modules.scala 65:57:@1066.4]
  wire [10:0] buffer_0_164; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55027; // @[Modules.scala 65:57:@1068.4]
  wire [10:0] _T_55028; // @[Modules.scala 65:57:@1069.4]
  wire [10:0] buffer_0_474; // @[Modules.scala 65:57:@1070.4]
  wire [10:0] buffer_0_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55030; // @[Modules.scala 65:57:@1072.4]
  wire [10:0] _T_55031; // @[Modules.scala 65:57:@1073.4]
  wire [10:0] buffer_0_475; // @[Modules.scala 65:57:@1074.4]
  wire [10:0] buffer_0_168; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55033; // @[Modules.scala 65:57:@1076.4]
  wire [10:0] _T_55034; // @[Modules.scala 65:57:@1077.4]
  wire [10:0] buffer_0_476; // @[Modules.scala 65:57:@1078.4]
  wire [10:0] buffer_0_170; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55036; // @[Modules.scala 65:57:@1080.4]
  wire [10:0] _T_55037; // @[Modules.scala 65:57:@1081.4]
  wire [10:0] buffer_0_477; // @[Modules.scala 65:57:@1082.4]
  wire [10:0] buffer_0_172; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55039; // @[Modules.scala 65:57:@1084.4]
  wire [10:0] _T_55040; // @[Modules.scala 65:57:@1085.4]
  wire [10:0] buffer_0_478; // @[Modules.scala 65:57:@1086.4]
  wire [10:0] buffer_0_174; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_175; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55042; // @[Modules.scala 65:57:@1088.4]
  wire [10:0] _T_55043; // @[Modules.scala 65:57:@1089.4]
  wire [10:0] buffer_0_479; // @[Modules.scala 65:57:@1090.4]
  wire [10:0] buffer_0_176; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55045; // @[Modules.scala 65:57:@1092.4]
  wire [10:0] _T_55046; // @[Modules.scala 65:57:@1093.4]
  wire [10:0] buffer_0_480; // @[Modules.scala 65:57:@1094.4]
  wire [10:0] buffer_0_178; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55048; // @[Modules.scala 65:57:@1096.4]
  wire [10:0] _T_55049; // @[Modules.scala 65:57:@1097.4]
  wire [10:0] buffer_0_481; // @[Modules.scala 65:57:@1098.4]
  wire [10:0] buffer_0_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55051; // @[Modules.scala 65:57:@1100.4]
  wire [10:0] _T_55052; // @[Modules.scala 65:57:@1101.4]
  wire [10:0] buffer_0_482; // @[Modules.scala 65:57:@1102.4]
  wire [10:0] buffer_0_184; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55057; // @[Modules.scala 65:57:@1108.4]
  wire [10:0] _T_55058; // @[Modules.scala 65:57:@1109.4]
  wire [10:0] buffer_0_484; // @[Modules.scala 65:57:@1110.4]
  wire [10:0] buffer_0_186; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_187; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55060; // @[Modules.scala 65:57:@1112.4]
  wire [10:0] _T_55061; // @[Modules.scala 65:57:@1113.4]
  wire [10:0] buffer_0_485; // @[Modules.scala 65:57:@1114.4]
  wire [10:0] buffer_0_188; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55063; // @[Modules.scala 65:57:@1116.4]
  wire [10:0] _T_55064; // @[Modules.scala 65:57:@1117.4]
  wire [10:0] buffer_0_486; // @[Modules.scala 65:57:@1118.4]
  wire [10:0] buffer_0_190; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55066; // @[Modules.scala 65:57:@1120.4]
  wire [10:0] _T_55067; // @[Modules.scala 65:57:@1121.4]
  wire [10:0] buffer_0_487; // @[Modules.scala 65:57:@1122.4]
  wire [10:0] buffer_0_192; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_193; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55069; // @[Modules.scala 65:57:@1124.4]
  wire [10:0] _T_55070; // @[Modules.scala 65:57:@1125.4]
  wire [10:0] buffer_0_488; // @[Modules.scala 65:57:@1126.4]
  wire [10:0] buffer_0_194; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55072; // @[Modules.scala 65:57:@1128.4]
  wire [10:0] _T_55073; // @[Modules.scala 65:57:@1129.4]
  wire [10:0] buffer_0_489; // @[Modules.scala 65:57:@1130.4]
  wire [10:0] buffer_0_198; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55078; // @[Modules.scala 65:57:@1136.4]
  wire [10:0] _T_55079; // @[Modules.scala 65:57:@1137.4]
  wire [10:0] buffer_0_491; // @[Modules.scala 65:57:@1138.4]
  wire [10:0] buffer_0_200; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_201; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55081; // @[Modules.scala 65:57:@1140.4]
  wire [10:0] _T_55082; // @[Modules.scala 65:57:@1141.4]
  wire [10:0] buffer_0_492; // @[Modules.scala 65:57:@1142.4]
  wire [10:0] buffer_0_202; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55084; // @[Modules.scala 65:57:@1144.4]
  wire [10:0] _T_55085; // @[Modules.scala 65:57:@1145.4]
  wire [10:0] buffer_0_493; // @[Modules.scala 65:57:@1146.4]
  wire [10:0] buffer_0_204; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55087; // @[Modules.scala 65:57:@1148.4]
  wire [10:0] _T_55088; // @[Modules.scala 65:57:@1149.4]
  wire [10:0] buffer_0_494; // @[Modules.scala 65:57:@1150.4]
  wire [10:0] buffer_0_206; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_207; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55090; // @[Modules.scala 65:57:@1152.4]
  wire [10:0] _T_55091; // @[Modules.scala 65:57:@1153.4]
  wire [10:0] buffer_0_495; // @[Modules.scala 65:57:@1154.4]
  wire [10:0] buffer_0_208; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55093; // @[Modules.scala 65:57:@1156.4]
  wire [10:0] _T_55094; // @[Modules.scala 65:57:@1157.4]
  wire [10:0] buffer_0_496; // @[Modules.scala 65:57:@1158.4]
  wire [10:0] buffer_0_210; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55096; // @[Modules.scala 65:57:@1160.4]
  wire [10:0] _T_55097; // @[Modules.scala 65:57:@1161.4]
  wire [10:0] buffer_0_497; // @[Modules.scala 65:57:@1162.4]
  wire [10:0] buffer_0_212; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55099; // @[Modules.scala 65:57:@1164.4]
  wire [10:0] _T_55100; // @[Modules.scala 65:57:@1165.4]
  wire [10:0] buffer_0_498; // @[Modules.scala 65:57:@1166.4]
  wire [10:0] buffer_0_214; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55102; // @[Modules.scala 65:57:@1168.4]
  wire [10:0] _T_55103; // @[Modules.scala 65:57:@1169.4]
  wire [10:0] buffer_0_499; // @[Modules.scala 65:57:@1170.4]
  wire [10:0] buffer_0_216; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55105; // @[Modules.scala 65:57:@1172.4]
  wire [10:0] _T_55106; // @[Modules.scala 65:57:@1173.4]
  wire [10:0] buffer_0_500; // @[Modules.scala 65:57:@1174.4]
  wire [10:0] buffer_0_218; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55108; // @[Modules.scala 65:57:@1176.4]
  wire [10:0] _T_55109; // @[Modules.scala 65:57:@1177.4]
  wire [10:0] buffer_0_501; // @[Modules.scala 65:57:@1178.4]
  wire [10:0] buffer_0_220; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55111; // @[Modules.scala 65:57:@1180.4]
  wire [10:0] _T_55112; // @[Modules.scala 65:57:@1181.4]
  wire [10:0] buffer_0_502; // @[Modules.scala 65:57:@1182.4]
  wire [10:0] buffer_0_224; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55117; // @[Modules.scala 65:57:@1188.4]
  wire [10:0] _T_55118; // @[Modules.scala 65:57:@1189.4]
  wire [10:0] buffer_0_504; // @[Modules.scala 65:57:@1190.4]
  wire [10:0] buffer_0_226; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55120; // @[Modules.scala 65:57:@1192.4]
  wire [10:0] _T_55121; // @[Modules.scala 65:57:@1193.4]
  wire [10:0] buffer_0_505; // @[Modules.scala 65:57:@1194.4]
  wire [10:0] buffer_0_228; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55123; // @[Modules.scala 65:57:@1196.4]
  wire [10:0] _T_55124; // @[Modules.scala 65:57:@1197.4]
  wire [10:0] buffer_0_506; // @[Modules.scala 65:57:@1198.4]
  wire [10:0] buffer_0_230; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55126; // @[Modules.scala 65:57:@1200.4]
  wire [10:0] _T_55127; // @[Modules.scala 65:57:@1201.4]
  wire [10:0] buffer_0_507; // @[Modules.scala 65:57:@1202.4]
  wire [10:0] buffer_0_232; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55129; // @[Modules.scala 65:57:@1204.4]
  wire [10:0] _T_55130; // @[Modules.scala 65:57:@1205.4]
  wire [10:0] buffer_0_508; // @[Modules.scala 65:57:@1206.4]
  wire [10:0] buffer_0_234; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55132; // @[Modules.scala 65:57:@1208.4]
  wire [10:0] _T_55133; // @[Modules.scala 65:57:@1209.4]
  wire [10:0] buffer_0_509; // @[Modules.scala 65:57:@1210.4]
  wire [10:0] buffer_0_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55138; // @[Modules.scala 65:57:@1216.4]
  wire [10:0] _T_55139; // @[Modules.scala 65:57:@1217.4]
  wire [10:0] buffer_0_511; // @[Modules.scala 65:57:@1218.4]
  wire [10:0] buffer_0_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55141; // @[Modules.scala 65:57:@1220.4]
  wire [10:0] _T_55142; // @[Modules.scala 65:57:@1221.4]
  wire [10:0] buffer_0_512; // @[Modules.scala 65:57:@1222.4]
  wire [10:0] buffer_0_242; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_243; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55144; // @[Modules.scala 65:57:@1224.4]
  wire [10:0] _T_55145; // @[Modules.scala 65:57:@1225.4]
  wire [10:0] buffer_0_513; // @[Modules.scala 65:57:@1226.4]
  wire [10:0] buffer_0_244; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55147; // @[Modules.scala 65:57:@1228.4]
  wire [10:0] _T_55148; // @[Modules.scala 65:57:@1229.4]
  wire [10:0] buffer_0_514; // @[Modules.scala 65:57:@1230.4]
  wire [10:0] buffer_0_246; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55150; // @[Modules.scala 65:57:@1232.4]
  wire [10:0] _T_55151; // @[Modules.scala 65:57:@1233.4]
  wire [10:0] buffer_0_515; // @[Modules.scala 65:57:@1234.4]
  wire [10:0] buffer_0_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55153; // @[Modules.scala 65:57:@1236.4]
  wire [10:0] _T_55154; // @[Modules.scala 65:57:@1237.4]
  wire [10:0] buffer_0_516; // @[Modules.scala 65:57:@1238.4]
  wire [10:0] buffer_0_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55159; // @[Modules.scala 65:57:@1244.4]
  wire [10:0] _T_55160; // @[Modules.scala 65:57:@1245.4]
  wire [10:0] buffer_0_518; // @[Modules.scala 65:57:@1246.4]
  wire [10:0] buffer_0_256; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_257; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55165; // @[Modules.scala 65:57:@1252.4]
  wire [10:0] _T_55166; // @[Modules.scala 65:57:@1253.4]
  wire [10:0] buffer_0_520; // @[Modules.scala 65:57:@1254.4]
  wire [10:0] buffer_0_258; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55168; // @[Modules.scala 65:57:@1256.4]
  wire [10:0] _T_55169; // @[Modules.scala 65:57:@1257.4]
  wire [10:0] buffer_0_521; // @[Modules.scala 65:57:@1258.4]
  wire [10:0] buffer_0_260; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_261; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55171; // @[Modules.scala 65:57:@1260.4]
  wire [10:0] _T_55172; // @[Modules.scala 65:57:@1261.4]
  wire [10:0] buffer_0_522; // @[Modules.scala 65:57:@1262.4]
  wire [10:0] buffer_0_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55174; // @[Modules.scala 65:57:@1264.4]
  wire [10:0] _T_55175; // @[Modules.scala 65:57:@1265.4]
  wire [10:0] buffer_0_523; // @[Modules.scala 65:57:@1266.4]
  wire [10:0] buffer_0_264; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55177; // @[Modules.scala 65:57:@1268.4]
  wire [10:0] _T_55178; // @[Modules.scala 65:57:@1269.4]
  wire [10:0] buffer_0_524; // @[Modules.scala 65:57:@1270.4]
  wire [10:0] buffer_0_266; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_267; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55180; // @[Modules.scala 65:57:@1272.4]
  wire [10:0] _T_55181; // @[Modules.scala 65:57:@1273.4]
  wire [10:0] buffer_0_525; // @[Modules.scala 65:57:@1274.4]
  wire [10:0] buffer_0_271; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55186; // @[Modules.scala 65:57:@1280.4]
  wire [10:0] _T_55187; // @[Modules.scala 65:57:@1281.4]
  wire [10:0] buffer_0_527; // @[Modules.scala 65:57:@1282.4]
  wire [10:0] buffer_0_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55192; // @[Modules.scala 65:57:@1288.4]
  wire [10:0] _T_55193; // @[Modules.scala 65:57:@1289.4]
  wire [10:0] buffer_0_529; // @[Modules.scala 65:57:@1290.4]
  wire [10:0] buffer_0_276; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55195; // @[Modules.scala 65:57:@1292.4]
  wire [10:0] _T_55196; // @[Modules.scala 65:57:@1293.4]
  wire [10:0] buffer_0_530; // @[Modules.scala 65:57:@1294.4]
  wire [10:0] buffer_0_278; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55198; // @[Modules.scala 65:57:@1296.4]
  wire [10:0] _T_55199; // @[Modules.scala 65:57:@1297.4]
  wire [10:0] buffer_0_531; // @[Modules.scala 65:57:@1298.4]
  wire [10:0] buffer_0_285; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55207; // @[Modules.scala 65:57:@1308.4]
  wire [10:0] _T_55208; // @[Modules.scala 65:57:@1309.4]
  wire [10:0] buffer_0_534; // @[Modules.scala 65:57:@1310.4]
  wire [10:0] buffer_0_286; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55210; // @[Modules.scala 65:57:@1312.4]
  wire [10:0] _T_55211; // @[Modules.scala 65:57:@1313.4]
  wire [10:0] buffer_0_535; // @[Modules.scala 65:57:@1314.4]
  wire [10:0] buffer_0_288; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55213; // @[Modules.scala 65:57:@1316.4]
  wire [10:0] _T_55214; // @[Modules.scala 65:57:@1317.4]
  wire [10:0] buffer_0_536; // @[Modules.scala 65:57:@1318.4]
  wire [10:0] buffer_0_290; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55216; // @[Modules.scala 65:57:@1320.4]
  wire [10:0] _T_55217; // @[Modules.scala 65:57:@1321.4]
  wire [10:0] buffer_0_537; // @[Modules.scala 65:57:@1322.4]
  wire [10:0] buffer_0_292; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55219; // @[Modules.scala 65:57:@1324.4]
  wire [10:0] _T_55220; // @[Modules.scala 65:57:@1325.4]
  wire [10:0] buffer_0_538; // @[Modules.scala 65:57:@1326.4]
  wire [10:0] buffer_0_294; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55222; // @[Modules.scala 65:57:@1328.4]
  wire [10:0] _T_55223; // @[Modules.scala 65:57:@1329.4]
  wire [10:0] buffer_0_539; // @[Modules.scala 65:57:@1330.4]
  wire [10:0] buffer_0_300; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55231; // @[Modules.scala 65:57:@1340.4]
  wire [10:0] _T_55232; // @[Modules.scala 65:57:@1341.4]
  wire [10:0] buffer_0_542; // @[Modules.scala 65:57:@1342.4]
  wire [10:0] buffer_0_302; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_303; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55234; // @[Modules.scala 65:57:@1344.4]
  wire [10:0] _T_55235; // @[Modules.scala 65:57:@1345.4]
  wire [10:0] buffer_0_543; // @[Modules.scala 65:57:@1346.4]
  wire [10:0] buffer_0_306; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55240; // @[Modules.scala 65:57:@1352.4]
  wire [10:0] _T_55241; // @[Modules.scala 65:57:@1353.4]
  wire [10:0] buffer_0_545; // @[Modules.scala 65:57:@1354.4]
  wire [10:0] buffer_0_308; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55243; // @[Modules.scala 65:57:@1356.4]
  wire [10:0] _T_55244; // @[Modules.scala 65:57:@1357.4]
  wire [10:0] buffer_0_546; // @[Modules.scala 65:57:@1358.4]
  wire [10:0] buffer_0_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55258; // @[Modules.scala 65:57:@1376.4]
  wire [10:0] _T_55259; // @[Modules.scala 65:57:@1377.4]
  wire [10:0] buffer_0_551; // @[Modules.scala 65:57:@1378.4]
  wire [10:0] buffer_0_320; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55261; // @[Modules.scala 65:57:@1380.4]
  wire [10:0] _T_55262; // @[Modules.scala 65:57:@1381.4]
  wire [10:0] buffer_0_552; // @[Modules.scala 65:57:@1382.4]
  wire [10:0] buffer_0_322; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_323; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55264; // @[Modules.scala 65:57:@1384.4]
  wire [10:0] _T_55265; // @[Modules.scala 65:57:@1385.4]
  wire [10:0] buffer_0_553; // @[Modules.scala 65:57:@1386.4]
  wire [10:0] buffer_0_331; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55276; // @[Modules.scala 65:57:@1400.4]
  wire [10:0] _T_55277; // @[Modules.scala 65:57:@1401.4]
  wire [10:0] buffer_0_557; // @[Modules.scala 65:57:@1402.4]
  wire [10:0] buffer_0_332; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_333; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55279; // @[Modules.scala 65:57:@1404.4]
  wire [10:0] _T_55280; // @[Modules.scala 65:57:@1405.4]
  wire [10:0] buffer_0_558; // @[Modules.scala 65:57:@1406.4]
  wire [10:0] buffer_0_334; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55282; // @[Modules.scala 65:57:@1408.4]
  wire [10:0] _T_55283; // @[Modules.scala 65:57:@1409.4]
  wire [10:0] buffer_0_559; // @[Modules.scala 65:57:@1410.4]
  wire [10:0] buffer_0_336; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55285; // @[Modules.scala 65:57:@1412.4]
  wire [10:0] _T_55286; // @[Modules.scala 65:57:@1413.4]
  wire [10:0] buffer_0_560; // @[Modules.scala 65:57:@1414.4]
  wire [10:0] buffer_0_338; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55288; // @[Modules.scala 65:57:@1416.4]
  wire [10:0] _T_55289; // @[Modules.scala 65:57:@1417.4]
  wire [10:0] buffer_0_561; // @[Modules.scala 65:57:@1418.4]
  wire [10:0] buffer_0_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55291; // @[Modules.scala 65:57:@1420.4]
  wire [10:0] _T_55292; // @[Modules.scala 65:57:@1421.4]
  wire [10:0] buffer_0_562; // @[Modules.scala 65:57:@1422.4]
  wire [10:0] buffer_0_344; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55297; // @[Modules.scala 65:57:@1428.4]
  wire [10:0] _T_55298; // @[Modules.scala 65:57:@1429.4]
  wire [10:0] buffer_0_564; // @[Modules.scala 65:57:@1430.4]
  wire [10:0] buffer_0_346; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55300; // @[Modules.scala 65:57:@1432.4]
  wire [10:0] _T_55301; // @[Modules.scala 65:57:@1433.4]
  wire [10:0] buffer_0_565; // @[Modules.scala 65:57:@1434.4]
  wire [10:0] buffer_0_348; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55303; // @[Modules.scala 65:57:@1436.4]
  wire [10:0] _T_55304; // @[Modules.scala 65:57:@1437.4]
  wire [10:0] buffer_0_566; // @[Modules.scala 65:57:@1438.4]
  wire [10:0] buffer_0_350; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55306; // @[Modules.scala 65:57:@1440.4]
  wire [10:0] _T_55307; // @[Modules.scala 65:57:@1441.4]
  wire [10:0] buffer_0_567; // @[Modules.scala 65:57:@1442.4]
  wire [10:0] buffer_0_352; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_353; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55309; // @[Modules.scala 65:57:@1444.4]
  wire [10:0] _T_55310; // @[Modules.scala 65:57:@1445.4]
  wire [10:0] buffer_0_568; // @[Modules.scala 65:57:@1446.4]
  wire [10:0] buffer_0_354; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55312; // @[Modules.scala 65:57:@1448.4]
  wire [10:0] _T_55313; // @[Modules.scala 65:57:@1449.4]
  wire [10:0] buffer_0_569; // @[Modules.scala 65:57:@1450.4]
  wire [10:0] buffer_0_356; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55315; // @[Modules.scala 65:57:@1452.4]
  wire [10:0] _T_55316; // @[Modules.scala 65:57:@1453.4]
  wire [10:0] buffer_0_570; // @[Modules.scala 65:57:@1454.4]
  wire [10:0] buffer_0_358; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_359; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55318; // @[Modules.scala 65:57:@1456.4]
  wire [10:0] _T_55319; // @[Modules.scala 65:57:@1457.4]
  wire [10:0] buffer_0_571; // @[Modules.scala 65:57:@1458.4]
  wire [10:0] buffer_0_360; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55321; // @[Modules.scala 65:57:@1460.4]
  wire [10:0] _T_55322; // @[Modules.scala 65:57:@1461.4]
  wire [10:0] buffer_0_572; // @[Modules.scala 65:57:@1462.4]
  wire [10:0] buffer_0_362; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55324; // @[Modules.scala 65:57:@1464.4]
  wire [10:0] _T_55325; // @[Modules.scala 65:57:@1465.4]
  wire [10:0] buffer_0_573; // @[Modules.scala 65:57:@1466.4]
  wire [10:0] buffer_0_364; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55327; // @[Modules.scala 65:57:@1468.4]
  wire [10:0] _T_55328; // @[Modules.scala 65:57:@1469.4]
  wire [10:0] buffer_0_574; // @[Modules.scala 65:57:@1470.4]
  wire [10:0] buffer_0_366; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55330; // @[Modules.scala 65:57:@1472.4]
  wire [10:0] _T_55331; // @[Modules.scala 65:57:@1473.4]
  wire [10:0] buffer_0_575; // @[Modules.scala 65:57:@1474.4]
  wire [10:0] buffer_0_370; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55336; // @[Modules.scala 65:57:@1480.4]
  wire [10:0] _T_55337; // @[Modules.scala 65:57:@1481.4]
  wire [10:0] buffer_0_577; // @[Modules.scala 65:57:@1482.4]
  wire [10:0] buffer_0_374; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55342; // @[Modules.scala 65:57:@1488.4]
  wire [10:0] _T_55343; // @[Modules.scala 65:57:@1489.4]
  wire [10:0] buffer_0_579; // @[Modules.scala 65:57:@1490.4]
  wire [10:0] buffer_0_376; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55345; // @[Modules.scala 65:57:@1492.4]
  wire [10:0] _T_55346; // @[Modules.scala 65:57:@1493.4]
  wire [10:0] buffer_0_580; // @[Modules.scala 65:57:@1494.4]
  wire [10:0] buffer_0_378; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55348; // @[Modules.scala 65:57:@1496.4]
  wire [10:0] _T_55349; // @[Modules.scala 65:57:@1497.4]
  wire [10:0] buffer_0_581; // @[Modules.scala 65:57:@1498.4]
  wire [10:0] buffer_0_380; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55351; // @[Modules.scala 65:57:@1500.4]
  wire [10:0] _T_55352; // @[Modules.scala 65:57:@1501.4]
  wire [10:0] buffer_0_582; // @[Modules.scala 65:57:@1502.4]
  wire [10:0] buffer_0_384; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_385; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55357; // @[Modules.scala 65:57:@1508.4]
  wire [10:0] _T_55358; // @[Modules.scala 65:57:@1509.4]
  wire [10:0] buffer_0_584; // @[Modules.scala 65:57:@1510.4]
  wire [10:0] buffer_0_388; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55363; // @[Modules.scala 65:57:@1516.4]
  wire [10:0] _T_55364; // @[Modules.scala 65:57:@1517.4]
  wire [10:0] buffer_0_586; // @[Modules.scala 65:57:@1518.4]
  wire [10:0] buffer_0_390; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_0_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_55366; // @[Modules.scala 65:57:@1520.4]
  wire [10:0] _T_55367; // @[Modules.scala 65:57:@1521.4]
  wire [10:0] buffer_0_587; // @[Modules.scala 65:57:@1522.4]
  wire [11:0] _T_55369; // @[Modules.scala 68:83:@1524.4]
  wire [10:0] _T_55370; // @[Modules.scala 68:83:@1525.4]
  wire [10:0] buffer_0_588; // @[Modules.scala 68:83:@1526.4]
  wire [11:0] _T_55372; // @[Modules.scala 68:83:@1528.4]
  wire [10:0] _T_55373; // @[Modules.scala 68:83:@1529.4]
  wire [10:0] buffer_0_589; // @[Modules.scala 68:83:@1530.4]
  wire [11:0] _T_55375; // @[Modules.scala 68:83:@1532.4]
  wire [10:0] _T_55376; // @[Modules.scala 68:83:@1533.4]
  wire [10:0] buffer_0_590; // @[Modules.scala 68:83:@1534.4]
  wire [11:0] _T_55378; // @[Modules.scala 68:83:@1536.4]
  wire [10:0] _T_55379; // @[Modules.scala 68:83:@1537.4]
  wire [10:0] buffer_0_591; // @[Modules.scala 68:83:@1538.4]
  wire [11:0] _T_55381; // @[Modules.scala 68:83:@1540.4]
  wire [10:0] _T_55382; // @[Modules.scala 68:83:@1541.4]
  wire [10:0] buffer_0_592; // @[Modules.scala 68:83:@1542.4]
  wire [11:0] _T_55384; // @[Modules.scala 68:83:@1544.4]
  wire [10:0] _T_55385; // @[Modules.scala 68:83:@1545.4]
  wire [10:0] buffer_0_593; // @[Modules.scala 68:83:@1546.4]
  wire [11:0] _T_55387; // @[Modules.scala 68:83:@1548.4]
  wire [10:0] _T_55388; // @[Modules.scala 68:83:@1549.4]
  wire [10:0] buffer_0_594; // @[Modules.scala 68:83:@1550.4]
  wire [11:0] _T_55390; // @[Modules.scala 68:83:@1552.4]
  wire [10:0] _T_55391; // @[Modules.scala 68:83:@1553.4]
  wire [10:0] buffer_0_595; // @[Modules.scala 68:83:@1554.4]
  wire [11:0] _T_55393; // @[Modules.scala 68:83:@1556.4]
  wire [10:0] _T_55394; // @[Modules.scala 68:83:@1557.4]
  wire [10:0] buffer_0_596; // @[Modules.scala 68:83:@1558.4]
  wire [11:0] _T_55396; // @[Modules.scala 68:83:@1560.4]
  wire [10:0] _T_55397; // @[Modules.scala 68:83:@1561.4]
  wire [10:0] buffer_0_597; // @[Modules.scala 68:83:@1562.4]
  wire [11:0] _T_55399; // @[Modules.scala 68:83:@1564.4]
  wire [10:0] _T_55400; // @[Modules.scala 68:83:@1565.4]
  wire [10:0] buffer_0_598; // @[Modules.scala 68:83:@1566.4]
  wire [11:0] _T_55402; // @[Modules.scala 68:83:@1568.4]
  wire [10:0] _T_55403; // @[Modules.scala 68:83:@1569.4]
  wire [10:0] buffer_0_599; // @[Modules.scala 68:83:@1570.4]
  wire [11:0] _T_55405; // @[Modules.scala 68:83:@1572.4]
  wire [10:0] _T_55406; // @[Modules.scala 68:83:@1573.4]
  wire [10:0] buffer_0_600; // @[Modules.scala 68:83:@1574.4]
  wire [11:0] _T_55408; // @[Modules.scala 68:83:@1576.4]
  wire [10:0] _T_55409; // @[Modules.scala 68:83:@1577.4]
  wire [10:0] buffer_0_601; // @[Modules.scala 68:83:@1578.4]
  wire [11:0] _T_55411; // @[Modules.scala 68:83:@1580.4]
  wire [10:0] _T_55412; // @[Modules.scala 68:83:@1581.4]
  wire [10:0] buffer_0_602; // @[Modules.scala 68:83:@1582.4]
  wire [11:0] _T_55417; // @[Modules.scala 68:83:@1588.4]
  wire [10:0] _T_55418; // @[Modules.scala 68:83:@1589.4]
  wire [10:0] buffer_0_604; // @[Modules.scala 68:83:@1590.4]
  wire [11:0] _T_55420; // @[Modules.scala 68:83:@1592.4]
  wire [10:0] _T_55421; // @[Modules.scala 68:83:@1593.4]
  wire [10:0] buffer_0_605; // @[Modules.scala 68:83:@1594.4]
  wire [11:0] _T_55423; // @[Modules.scala 68:83:@1596.4]
  wire [10:0] _T_55424; // @[Modules.scala 68:83:@1597.4]
  wire [10:0] buffer_0_606; // @[Modules.scala 68:83:@1598.4]
  wire [11:0] _T_55429; // @[Modules.scala 68:83:@1604.4]
  wire [10:0] _T_55430; // @[Modules.scala 68:83:@1605.4]
  wire [10:0] buffer_0_608; // @[Modules.scala 68:83:@1606.4]
  wire [11:0] _T_55432; // @[Modules.scala 68:83:@1608.4]
  wire [10:0] _T_55433; // @[Modules.scala 68:83:@1609.4]
  wire [10:0] buffer_0_609; // @[Modules.scala 68:83:@1610.4]
  wire [11:0] _T_55438; // @[Modules.scala 68:83:@1616.4]
  wire [10:0] _T_55439; // @[Modules.scala 68:83:@1617.4]
  wire [10:0] buffer_0_611; // @[Modules.scala 68:83:@1618.4]
  wire [11:0] _T_55441; // @[Modules.scala 68:83:@1620.4]
  wire [10:0] _T_55442; // @[Modules.scala 68:83:@1621.4]
  wire [10:0] buffer_0_612; // @[Modules.scala 68:83:@1622.4]
  wire [11:0] _T_55444; // @[Modules.scala 68:83:@1624.4]
  wire [10:0] _T_55445; // @[Modules.scala 68:83:@1625.4]
  wire [10:0] buffer_0_613; // @[Modules.scala 68:83:@1626.4]
  wire [11:0] _T_55447; // @[Modules.scala 68:83:@1628.4]
  wire [10:0] _T_55448; // @[Modules.scala 68:83:@1629.4]
  wire [10:0] buffer_0_614; // @[Modules.scala 68:83:@1630.4]
  wire [11:0] _T_55456; // @[Modules.scala 68:83:@1640.4]
  wire [10:0] _T_55457; // @[Modules.scala 68:83:@1641.4]
  wire [10:0] buffer_0_617; // @[Modules.scala 68:83:@1642.4]
  wire [11:0] _T_55465; // @[Modules.scala 68:83:@1652.4]
  wire [10:0] _T_55466; // @[Modules.scala 68:83:@1653.4]
  wire [10:0] buffer_0_620; // @[Modules.scala 68:83:@1654.4]
  wire [11:0] _T_55477; // @[Modules.scala 68:83:@1668.4]
  wire [10:0] _T_55478; // @[Modules.scala 68:83:@1669.4]
  wire [10:0] buffer_0_624; // @[Modules.scala 68:83:@1670.4]
  wire [11:0] _T_55486; // @[Modules.scala 68:83:@1680.4]
  wire [10:0] _T_55487; // @[Modules.scala 68:83:@1681.4]
  wire [10:0] buffer_0_627; // @[Modules.scala 68:83:@1682.4]
  wire [11:0] _T_55489; // @[Modules.scala 68:83:@1684.4]
  wire [10:0] _T_55490; // @[Modules.scala 68:83:@1685.4]
  wire [10:0] buffer_0_628; // @[Modules.scala 68:83:@1686.4]
  wire [11:0] _T_55492; // @[Modules.scala 68:83:@1688.4]
  wire [10:0] _T_55493; // @[Modules.scala 68:83:@1689.4]
  wire [10:0] buffer_0_629; // @[Modules.scala 68:83:@1690.4]
  wire [11:0] _T_55495; // @[Modules.scala 68:83:@1692.4]
  wire [10:0] _T_55496; // @[Modules.scala 68:83:@1693.4]
  wire [10:0] buffer_0_630; // @[Modules.scala 68:83:@1694.4]
  wire [11:0] _T_55498; // @[Modules.scala 68:83:@1696.4]
  wire [10:0] _T_55499; // @[Modules.scala 68:83:@1697.4]
  wire [10:0] buffer_0_631; // @[Modules.scala 68:83:@1698.4]
  wire [11:0] _T_55501; // @[Modules.scala 68:83:@1700.4]
  wire [10:0] _T_55502; // @[Modules.scala 68:83:@1701.4]
  wire [10:0] buffer_0_632; // @[Modules.scala 68:83:@1702.4]
  wire [11:0] _T_55504; // @[Modules.scala 68:83:@1704.4]
  wire [10:0] _T_55505; // @[Modules.scala 68:83:@1705.4]
  wire [10:0] buffer_0_633; // @[Modules.scala 68:83:@1706.4]
  wire [11:0] _T_55507; // @[Modules.scala 68:83:@1708.4]
  wire [10:0] _T_55508; // @[Modules.scala 68:83:@1709.4]
  wire [10:0] buffer_0_634; // @[Modules.scala 68:83:@1710.4]
  wire [11:0] _T_55510; // @[Modules.scala 68:83:@1712.4]
  wire [10:0] _T_55511; // @[Modules.scala 68:83:@1713.4]
  wire [10:0] buffer_0_635; // @[Modules.scala 68:83:@1714.4]
  wire [11:0] _T_55513; // @[Modules.scala 68:83:@1716.4]
  wire [10:0] _T_55514; // @[Modules.scala 68:83:@1717.4]
  wire [10:0] buffer_0_636; // @[Modules.scala 68:83:@1718.4]
  wire [11:0] _T_55516; // @[Modules.scala 68:83:@1720.4]
  wire [10:0] _T_55517; // @[Modules.scala 68:83:@1721.4]
  wire [10:0] buffer_0_637; // @[Modules.scala 68:83:@1722.4]
  wire [11:0] _T_55519; // @[Modules.scala 68:83:@1724.4]
  wire [10:0] _T_55520; // @[Modules.scala 68:83:@1725.4]
  wire [10:0] buffer_0_638; // @[Modules.scala 68:83:@1726.4]
  wire [11:0] _T_55522; // @[Modules.scala 68:83:@1728.4]
  wire [10:0] _T_55523; // @[Modules.scala 68:83:@1729.4]
  wire [10:0] buffer_0_639; // @[Modules.scala 68:83:@1730.4]
  wire [11:0] _T_55525; // @[Modules.scala 68:83:@1732.4]
  wire [10:0] _T_55526; // @[Modules.scala 68:83:@1733.4]
  wire [10:0] buffer_0_640; // @[Modules.scala 68:83:@1734.4]
  wire [11:0] _T_55528; // @[Modules.scala 68:83:@1736.4]
  wire [10:0] _T_55529; // @[Modules.scala 68:83:@1737.4]
  wire [10:0] buffer_0_641; // @[Modules.scala 68:83:@1738.4]
  wire [11:0] _T_55531; // @[Modules.scala 68:83:@1740.4]
  wire [10:0] _T_55532; // @[Modules.scala 68:83:@1741.4]
  wire [10:0] buffer_0_642; // @[Modules.scala 68:83:@1742.4]
  wire [11:0] _T_55534; // @[Modules.scala 68:83:@1744.4]
  wire [10:0] _T_55535; // @[Modules.scala 68:83:@1745.4]
  wire [10:0] buffer_0_643; // @[Modules.scala 68:83:@1746.4]
  wire [11:0] _T_55537; // @[Modules.scala 68:83:@1748.4]
  wire [10:0] _T_55538; // @[Modules.scala 68:83:@1749.4]
  wire [10:0] buffer_0_644; // @[Modules.scala 68:83:@1750.4]
  wire [11:0] _T_55540; // @[Modules.scala 68:83:@1752.4]
  wire [10:0] _T_55541; // @[Modules.scala 68:83:@1753.4]
  wire [10:0] buffer_0_645; // @[Modules.scala 68:83:@1754.4]
  wire [11:0] _T_55543; // @[Modules.scala 68:83:@1756.4]
  wire [10:0] _T_55544; // @[Modules.scala 68:83:@1757.4]
  wire [10:0] buffer_0_646; // @[Modules.scala 68:83:@1758.4]
  wire [11:0] _T_55546; // @[Modules.scala 68:83:@1760.4]
  wire [10:0] _T_55547; // @[Modules.scala 68:83:@1761.4]
  wire [10:0] buffer_0_647; // @[Modules.scala 68:83:@1762.4]
  wire [11:0] _T_55549; // @[Modules.scala 68:83:@1764.4]
  wire [10:0] _T_55550; // @[Modules.scala 68:83:@1765.4]
  wire [10:0] buffer_0_648; // @[Modules.scala 68:83:@1766.4]
  wire [11:0] _T_55552; // @[Modules.scala 68:83:@1768.4]
  wire [10:0] _T_55553; // @[Modules.scala 68:83:@1769.4]
  wire [10:0] buffer_0_649; // @[Modules.scala 68:83:@1770.4]
  wire [11:0] _T_55555; // @[Modules.scala 68:83:@1772.4]
  wire [10:0] _T_55556; // @[Modules.scala 68:83:@1773.4]
  wire [10:0] buffer_0_650; // @[Modules.scala 68:83:@1774.4]
  wire [11:0] _T_55558; // @[Modules.scala 68:83:@1776.4]
  wire [10:0] _T_55559; // @[Modules.scala 68:83:@1777.4]
  wire [10:0] buffer_0_651; // @[Modules.scala 68:83:@1778.4]
  wire [11:0] _T_55561; // @[Modules.scala 68:83:@1780.4]
  wire [10:0] _T_55562; // @[Modules.scala 68:83:@1781.4]
  wire [10:0] buffer_0_652; // @[Modules.scala 68:83:@1782.4]
  wire [11:0] _T_55564; // @[Modules.scala 68:83:@1784.4]
  wire [10:0] _T_55565; // @[Modules.scala 68:83:@1785.4]
  wire [10:0] buffer_0_653; // @[Modules.scala 68:83:@1786.4]
  wire [11:0] _T_55567; // @[Modules.scala 68:83:@1788.4]
  wire [10:0] _T_55568; // @[Modules.scala 68:83:@1789.4]
  wire [10:0] buffer_0_654; // @[Modules.scala 68:83:@1790.4]
  wire [11:0] _T_55570; // @[Modules.scala 68:83:@1792.4]
  wire [10:0] _T_55571; // @[Modules.scala 68:83:@1793.4]
  wire [10:0] buffer_0_655; // @[Modules.scala 68:83:@1794.4]
  wire [11:0] _T_55573; // @[Modules.scala 68:83:@1796.4]
  wire [10:0] _T_55574; // @[Modules.scala 68:83:@1797.4]
  wire [10:0] buffer_0_656; // @[Modules.scala 68:83:@1798.4]
  wire [11:0] _T_55576; // @[Modules.scala 68:83:@1800.4]
  wire [10:0] _T_55577; // @[Modules.scala 68:83:@1801.4]
  wire [10:0] buffer_0_657; // @[Modules.scala 68:83:@1802.4]
  wire [11:0] _T_55582; // @[Modules.scala 68:83:@1808.4]
  wire [10:0] _T_55583; // @[Modules.scala 68:83:@1809.4]
  wire [10:0] buffer_0_659; // @[Modules.scala 68:83:@1810.4]
  wire [11:0] _T_55585; // @[Modules.scala 68:83:@1812.4]
  wire [10:0] _T_55586; // @[Modules.scala 68:83:@1813.4]
  wire [10:0] buffer_0_660; // @[Modules.scala 68:83:@1814.4]
  wire [11:0] _T_55588; // @[Modules.scala 68:83:@1816.4]
  wire [10:0] _T_55589; // @[Modules.scala 68:83:@1817.4]
  wire [10:0] buffer_0_661; // @[Modules.scala 68:83:@1818.4]
  wire [11:0] _T_55594; // @[Modules.scala 68:83:@1824.4]
  wire [10:0] _T_55595; // @[Modules.scala 68:83:@1825.4]
  wire [10:0] buffer_0_663; // @[Modules.scala 68:83:@1826.4]
  wire [11:0] _T_55597; // @[Modules.scala 68:83:@1828.4]
  wire [10:0] _T_55598; // @[Modules.scala 68:83:@1829.4]
  wire [10:0] buffer_0_664; // @[Modules.scala 68:83:@1830.4]
  wire [11:0] _T_55600; // @[Modules.scala 68:83:@1832.4]
  wire [10:0] _T_55601; // @[Modules.scala 68:83:@1833.4]
  wire [10:0] buffer_0_665; // @[Modules.scala 68:83:@1834.4]
  wire [11:0] _T_55606; // @[Modules.scala 68:83:@1840.4]
  wire [10:0] _T_55607; // @[Modules.scala 68:83:@1841.4]
  wire [10:0] buffer_0_667; // @[Modules.scala 68:83:@1842.4]
  wire [11:0] _T_55609; // @[Modules.scala 68:83:@1844.4]
  wire [10:0] _T_55610; // @[Modules.scala 68:83:@1845.4]
  wire [10:0] buffer_0_668; // @[Modules.scala 68:83:@1846.4]
  wire [11:0] _T_55615; // @[Modules.scala 68:83:@1852.4]
  wire [10:0] _T_55616; // @[Modules.scala 68:83:@1853.4]
  wire [10:0] buffer_0_670; // @[Modules.scala 68:83:@1854.4]
  wire [11:0] _T_55618; // @[Modules.scala 68:83:@1856.4]
  wire [10:0] _T_55619; // @[Modules.scala 68:83:@1857.4]
  wire [10:0] buffer_0_671; // @[Modules.scala 68:83:@1858.4]
  wire [11:0] _T_55621; // @[Modules.scala 68:83:@1860.4]
  wire [10:0] _T_55622; // @[Modules.scala 68:83:@1861.4]
  wire [10:0] buffer_0_672; // @[Modules.scala 68:83:@1862.4]
  wire [11:0] _T_55624; // @[Modules.scala 68:83:@1864.4]
  wire [10:0] _T_55625; // @[Modules.scala 68:83:@1865.4]
  wire [10:0] buffer_0_673; // @[Modules.scala 68:83:@1866.4]
  wire [11:0] _T_55627; // @[Modules.scala 68:83:@1868.4]
  wire [10:0] _T_55628; // @[Modules.scala 68:83:@1869.4]
  wire [10:0] buffer_0_674; // @[Modules.scala 68:83:@1870.4]
  wire [11:0] _T_55630; // @[Modules.scala 68:83:@1872.4]
  wire [10:0] _T_55631; // @[Modules.scala 68:83:@1873.4]
  wire [10:0] buffer_0_675; // @[Modules.scala 68:83:@1874.4]
  wire [11:0] _T_55633; // @[Modules.scala 68:83:@1876.4]
  wire [10:0] _T_55634; // @[Modules.scala 68:83:@1877.4]
  wire [10:0] buffer_0_676; // @[Modules.scala 68:83:@1878.4]
  wire [11:0] _T_55636; // @[Modules.scala 68:83:@1880.4]
  wire [10:0] _T_55637; // @[Modules.scala 68:83:@1881.4]
  wire [10:0] buffer_0_677; // @[Modules.scala 68:83:@1882.4]
  wire [11:0] _T_55639; // @[Modules.scala 68:83:@1884.4]
  wire [10:0] _T_55640; // @[Modules.scala 68:83:@1885.4]
  wire [10:0] buffer_0_678; // @[Modules.scala 68:83:@1886.4]
  wire [11:0] _T_55642; // @[Modules.scala 68:83:@1888.4]
  wire [10:0] _T_55643; // @[Modules.scala 68:83:@1889.4]
  wire [10:0] buffer_0_679; // @[Modules.scala 68:83:@1890.4]
  wire [11:0] _T_55645; // @[Modules.scala 68:83:@1892.4]
  wire [10:0] _T_55646; // @[Modules.scala 68:83:@1893.4]
  wire [10:0] buffer_0_680; // @[Modules.scala 68:83:@1894.4]
  wire [11:0] _T_55648; // @[Modules.scala 68:83:@1896.4]
  wire [10:0] _T_55649; // @[Modules.scala 68:83:@1897.4]
  wire [10:0] buffer_0_681; // @[Modules.scala 68:83:@1898.4]
  wire [11:0] _T_55651; // @[Modules.scala 68:83:@1900.4]
  wire [10:0] _T_55652; // @[Modules.scala 68:83:@1901.4]
  wire [10:0] buffer_0_682; // @[Modules.scala 68:83:@1902.4]
  wire [11:0] _T_55654; // @[Modules.scala 68:83:@1904.4]
  wire [10:0] _T_55655; // @[Modules.scala 68:83:@1905.4]
  wire [10:0] buffer_0_683; // @[Modules.scala 68:83:@1906.4]
  wire [11:0] _T_55657; // @[Modules.scala 68:83:@1908.4]
  wire [10:0] _T_55658; // @[Modules.scala 68:83:@1909.4]
  wire [10:0] buffer_0_684; // @[Modules.scala 68:83:@1910.4]
  wire [11:0] _T_55660; // @[Modules.scala 68:83:@1912.4]
  wire [10:0] _T_55661; // @[Modules.scala 68:83:@1913.4]
  wire [10:0] buffer_0_685; // @[Modules.scala 68:83:@1914.4]
  wire [11:0] _T_55663; // @[Modules.scala 71:109:@1916.4]
  wire [10:0] _T_55664; // @[Modules.scala 71:109:@1917.4]
  wire [10:0] buffer_0_686; // @[Modules.scala 71:109:@1918.4]
  wire [11:0] _T_55666; // @[Modules.scala 71:109:@1920.4]
  wire [10:0] _T_55667; // @[Modules.scala 71:109:@1921.4]
  wire [10:0] buffer_0_687; // @[Modules.scala 71:109:@1922.4]
  wire [11:0] _T_55669; // @[Modules.scala 71:109:@1924.4]
  wire [10:0] _T_55670; // @[Modules.scala 71:109:@1925.4]
  wire [10:0] buffer_0_688; // @[Modules.scala 71:109:@1926.4]
  wire [11:0] _T_55672; // @[Modules.scala 71:109:@1928.4]
  wire [10:0] _T_55673; // @[Modules.scala 71:109:@1929.4]
  wire [10:0] buffer_0_689; // @[Modules.scala 71:109:@1930.4]
  wire [11:0] _T_55675; // @[Modules.scala 71:109:@1932.4]
  wire [10:0] _T_55676; // @[Modules.scala 71:109:@1933.4]
  wire [10:0] buffer_0_690; // @[Modules.scala 71:109:@1934.4]
  wire [11:0] _T_55678; // @[Modules.scala 71:109:@1936.4]
  wire [10:0] _T_55679; // @[Modules.scala 71:109:@1937.4]
  wire [10:0] buffer_0_691; // @[Modules.scala 71:109:@1938.4]
  wire [11:0] _T_55681; // @[Modules.scala 71:109:@1940.4]
  wire [10:0] _T_55682; // @[Modules.scala 71:109:@1941.4]
  wire [10:0] buffer_0_692; // @[Modules.scala 71:109:@1942.4]
  wire [11:0] _T_55684; // @[Modules.scala 71:109:@1944.4]
  wire [10:0] _T_55685; // @[Modules.scala 71:109:@1945.4]
  wire [10:0] buffer_0_693; // @[Modules.scala 71:109:@1946.4]
  wire [11:0] _T_55687; // @[Modules.scala 71:109:@1948.4]
  wire [10:0] _T_55688; // @[Modules.scala 71:109:@1949.4]
  wire [10:0] buffer_0_694; // @[Modules.scala 71:109:@1950.4]
  wire [11:0] _T_55690; // @[Modules.scala 71:109:@1952.4]
  wire [10:0] _T_55691; // @[Modules.scala 71:109:@1953.4]
  wire [10:0] buffer_0_695; // @[Modules.scala 71:109:@1954.4]
  wire [11:0] _T_55693; // @[Modules.scala 71:109:@1956.4]
  wire [10:0] _T_55694; // @[Modules.scala 71:109:@1957.4]
  wire [10:0] buffer_0_696; // @[Modules.scala 71:109:@1958.4]
  wire [11:0] _T_55696; // @[Modules.scala 71:109:@1960.4]
  wire [10:0] _T_55697; // @[Modules.scala 71:109:@1961.4]
  wire [10:0] buffer_0_697; // @[Modules.scala 71:109:@1962.4]
  wire [11:0] _T_55699; // @[Modules.scala 71:109:@1964.4]
  wire [10:0] _T_55700; // @[Modules.scala 71:109:@1965.4]
  wire [10:0] buffer_0_698; // @[Modules.scala 71:109:@1966.4]
  wire [11:0] _T_55702; // @[Modules.scala 71:109:@1968.4]
  wire [10:0] _T_55703; // @[Modules.scala 71:109:@1969.4]
  wire [10:0] buffer_0_699; // @[Modules.scala 71:109:@1970.4]
  wire [11:0] _T_55705; // @[Modules.scala 71:109:@1972.4]
  wire [10:0] _T_55706; // @[Modules.scala 71:109:@1973.4]
  wire [10:0] buffer_0_700; // @[Modules.scala 71:109:@1974.4]
  wire [11:0] _T_55708; // @[Modules.scala 71:109:@1976.4]
  wire [10:0] _T_55709; // @[Modules.scala 71:109:@1977.4]
  wire [10:0] buffer_0_701; // @[Modules.scala 71:109:@1978.4]
  wire [11:0] _T_55711; // @[Modules.scala 71:109:@1980.4]
  wire [10:0] _T_55712; // @[Modules.scala 71:109:@1981.4]
  wire [10:0] buffer_0_702; // @[Modules.scala 71:109:@1982.4]
  wire [11:0] _T_55717; // @[Modules.scala 71:109:@1988.4]
  wire [10:0] _T_55718; // @[Modules.scala 71:109:@1989.4]
  wire [10:0] buffer_0_704; // @[Modules.scala 71:109:@1990.4]
  wire [11:0] _T_55720; // @[Modules.scala 71:109:@1992.4]
  wire [10:0] _T_55721; // @[Modules.scala 71:109:@1993.4]
  wire [10:0] buffer_0_705; // @[Modules.scala 71:109:@1994.4]
  wire [11:0] _T_55723; // @[Modules.scala 71:109:@1996.4]
  wire [10:0] _T_55724; // @[Modules.scala 71:109:@1997.4]
  wire [10:0] buffer_0_706; // @[Modules.scala 71:109:@1998.4]
  wire [11:0] _T_55726; // @[Modules.scala 71:109:@2000.4]
  wire [10:0] _T_55727; // @[Modules.scala 71:109:@2001.4]
  wire [10:0] buffer_0_707; // @[Modules.scala 71:109:@2002.4]
  wire [11:0] _T_55729; // @[Modules.scala 71:109:@2004.4]
  wire [10:0] _T_55730; // @[Modules.scala 71:109:@2005.4]
  wire [10:0] buffer_0_708; // @[Modules.scala 71:109:@2006.4]
  wire [11:0] _T_55732; // @[Modules.scala 71:109:@2008.4]
  wire [10:0] _T_55733; // @[Modules.scala 71:109:@2009.4]
  wire [10:0] buffer_0_709; // @[Modules.scala 71:109:@2010.4]
  wire [11:0] _T_55735; // @[Modules.scala 71:109:@2012.4]
  wire [10:0] _T_55736; // @[Modules.scala 71:109:@2013.4]
  wire [10:0] buffer_0_710; // @[Modules.scala 71:109:@2014.4]
  wire [11:0] _T_55738; // @[Modules.scala 71:109:@2016.4]
  wire [10:0] _T_55739; // @[Modules.scala 71:109:@2017.4]
  wire [10:0] buffer_0_711; // @[Modules.scala 71:109:@2018.4]
  wire [11:0] _T_55741; // @[Modules.scala 71:109:@2020.4]
  wire [10:0] _T_55742; // @[Modules.scala 71:109:@2021.4]
  wire [10:0] buffer_0_712; // @[Modules.scala 71:109:@2022.4]
  wire [11:0] _T_55744; // @[Modules.scala 71:109:@2024.4]
  wire [10:0] _T_55745; // @[Modules.scala 71:109:@2025.4]
  wire [10:0] buffer_0_713; // @[Modules.scala 71:109:@2026.4]
  wire [11:0] _T_55747; // @[Modules.scala 71:109:@2028.4]
  wire [10:0] _T_55748; // @[Modules.scala 71:109:@2029.4]
  wire [10:0] buffer_0_714; // @[Modules.scala 71:109:@2030.4]
  wire [11:0] _T_55750; // @[Modules.scala 71:109:@2032.4]
  wire [10:0] _T_55751; // @[Modules.scala 71:109:@2033.4]
  wire [10:0] buffer_0_715; // @[Modules.scala 71:109:@2034.4]
  wire [11:0] _T_55753; // @[Modules.scala 71:109:@2036.4]
  wire [10:0] _T_55754; // @[Modules.scala 71:109:@2037.4]
  wire [10:0] buffer_0_716; // @[Modules.scala 71:109:@2038.4]
  wire [11:0] _T_55756; // @[Modules.scala 71:109:@2040.4]
  wire [10:0] _T_55757; // @[Modules.scala 71:109:@2041.4]
  wire [10:0] buffer_0_717; // @[Modules.scala 71:109:@2042.4]
  wire [11:0] _T_55759; // @[Modules.scala 71:109:@2044.4]
  wire [10:0] _T_55760; // @[Modules.scala 71:109:@2045.4]
  wire [10:0] buffer_0_718; // @[Modules.scala 71:109:@2046.4]
  wire [11:0] _T_55762; // @[Modules.scala 71:109:@2048.4]
  wire [10:0] _T_55763; // @[Modules.scala 71:109:@2049.4]
  wire [10:0] buffer_0_719; // @[Modules.scala 71:109:@2050.4]
  wire [11:0] _T_55765; // @[Modules.scala 71:109:@2052.4]
  wire [10:0] _T_55766; // @[Modules.scala 71:109:@2053.4]
  wire [10:0] buffer_0_720; // @[Modules.scala 71:109:@2054.4]
  wire [11:0] _T_55768; // @[Modules.scala 71:109:@2056.4]
  wire [10:0] _T_55769; // @[Modules.scala 71:109:@2057.4]
  wire [10:0] buffer_0_721; // @[Modules.scala 71:109:@2058.4]
  wire [11:0] _T_55771; // @[Modules.scala 71:109:@2060.4]
  wire [10:0] _T_55772; // @[Modules.scala 71:109:@2061.4]
  wire [10:0] buffer_0_722; // @[Modules.scala 71:109:@2062.4]
  wire [11:0] _T_55774; // @[Modules.scala 71:109:@2064.4]
  wire [10:0] _T_55775; // @[Modules.scala 71:109:@2065.4]
  wire [10:0] buffer_0_723; // @[Modules.scala 71:109:@2066.4]
  wire [11:0] _T_55777; // @[Modules.scala 71:109:@2068.4]
  wire [10:0] _T_55778; // @[Modules.scala 71:109:@2069.4]
  wire [10:0] buffer_0_724; // @[Modules.scala 71:109:@2070.4]
  wire [11:0] _T_55780; // @[Modules.scala 71:109:@2072.4]
  wire [10:0] _T_55781; // @[Modules.scala 71:109:@2073.4]
  wire [10:0] buffer_0_725; // @[Modules.scala 71:109:@2074.4]
  wire [11:0] _T_55783; // @[Modules.scala 71:109:@2076.4]
  wire [10:0] _T_55784; // @[Modules.scala 71:109:@2077.4]
  wire [10:0] buffer_0_726; // @[Modules.scala 71:109:@2078.4]
  wire [11:0] _T_55786; // @[Modules.scala 71:109:@2080.4]
  wire [10:0] _T_55787; // @[Modules.scala 71:109:@2081.4]
  wire [10:0] buffer_0_727; // @[Modules.scala 71:109:@2082.4]
  wire [11:0] _T_55789; // @[Modules.scala 71:109:@2084.4]
  wire [10:0] _T_55790; // @[Modules.scala 71:109:@2085.4]
  wire [10:0] buffer_0_728; // @[Modules.scala 71:109:@2086.4]
  wire [11:0] _T_55792; // @[Modules.scala 71:109:@2088.4]
  wire [10:0] _T_55793; // @[Modules.scala 71:109:@2089.4]
  wire [10:0] buffer_0_729; // @[Modules.scala 71:109:@2090.4]
  wire [11:0] _T_55795; // @[Modules.scala 71:109:@2092.4]
  wire [10:0] _T_55796; // @[Modules.scala 71:109:@2093.4]
  wire [10:0] buffer_0_730; // @[Modules.scala 71:109:@2094.4]
  wire [11:0] _T_55798; // @[Modules.scala 71:109:@2096.4]
  wire [10:0] _T_55799; // @[Modules.scala 71:109:@2097.4]
  wire [10:0] buffer_0_731; // @[Modules.scala 71:109:@2098.4]
  wire [11:0] _T_55801; // @[Modules.scala 71:109:@2100.4]
  wire [10:0] _T_55802; // @[Modules.scala 71:109:@2101.4]
  wire [10:0] buffer_0_732; // @[Modules.scala 71:109:@2102.4]
  wire [11:0] _T_55804; // @[Modules.scala 71:109:@2104.4]
  wire [10:0] _T_55805; // @[Modules.scala 71:109:@2105.4]
  wire [10:0] buffer_0_733; // @[Modules.scala 71:109:@2106.4]
  wire [11:0] _T_55807; // @[Modules.scala 71:109:@2108.4]
  wire [10:0] _T_55808; // @[Modules.scala 71:109:@2109.4]
  wire [10:0] buffer_0_734; // @[Modules.scala 71:109:@2110.4]
  wire [11:0] _T_55810; // @[Modules.scala 78:156:@2113.4]
  wire [10:0] _T_55811; // @[Modules.scala 78:156:@2114.4]
  wire [10:0] buffer_0_736; // @[Modules.scala 78:156:@2115.4]
  wire [11:0] _T_55813; // @[Modules.scala 78:156:@2117.4]
  wire [10:0] _T_55814; // @[Modules.scala 78:156:@2118.4]
  wire [10:0] buffer_0_737; // @[Modules.scala 78:156:@2119.4]
  wire [11:0] _T_55816; // @[Modules.scala 78:156:@2121.4]
  wire [10:0] _T_55817; // @[Modules.scala 78:156:@2122.4]
  wire [10:0] buffer_0_738; // @[Modules.scala 78:156:@2123.4]
  wire [11:0] _T_55819; // @[Modules.scala 78:156:@2125.4]
  wire [10:0] _T_55820; // @[Modules.scala 78:156:@2126.4]
  wire [10:0] buffer_0_739; // @[Modules.scala 78:156:@2127.4]
  wire [11:0] _T_55822; // @[Modules.scala 78:156:@2129.4]
  wire [10:0] _T_55823; // @[Modules.scala 78:156:@2130.4]
  wire [10:0] buffer_0_740; // @[Modules.scala 78:156:@2131.4]
  wire [11:0] _T_55825; // @[Modules.scala 78:156:@2133.4]
  wire [10:0] _T_55826; // @[Modules.scala 78:156:@2134.4]
  wire [10:0] buffer_0_741; // @[Modules.scala 78:156:@2135.4]
  wire [11:0] _T_55828; // @[Modules.scala 78:156:@2137.4]
  wire [10:0] _T_55829; // @[Modules.scala 78:156:@2138.4]
  wire [10:0] buffer_0_742; // @[Modules.scala 78:156:@2139.4]
  wire [11:0] _T_55831; // @[Modules.scala 78:156:@2141.4]
  wire [10:0] _T_55832; // @[Modules.scala 78:156:@2142.4]
  wire [10:0] buffer_0_743; // @[Modules.scala 78:156:@2143.4]
  wire [11:0] _T_55834; // @[Modules.scala 78:156:@2145.4]
  wire [10:0] _T_55835; // @[Modules.scala 78:156:@2146.4]
  wire [10:0] buffer_0_744; // @[Modules.scala 78:156:@2147.4]
  wire [11:0] _T_55837; // @[Modules.scala 78:156:@2149.4]
  wire [10:0] _T_55838; // @[Modules.scala 78:156:@2150.4]
  wire [10:0] buffer_0_745; // @[Modules.scala 78:156:@2151.4]
  wire [11:0] _T_55840; // @[Modules.scala 78:156:@2153.4]
  wire [10:0] _T_55841; // @[Modules.scala 78:156:@2154.4]
  wire [10:0] buffer_0_746; // @[Modules.scala 78:156:@2155.4]
  wire [11:0] _T_55843; // @[Modules.scala 78:156:@2157.4]
  wire [10:0] _T_55844; // @[Modules.scala 78:156:@2158.4]
  wire [10:0] buffer_0_747; // @[Modules.scala 78:156:@2159.4]
  wire [11:0] _T_55846; // @[Modules.scala 78:156:@2161.4]
  wire [10:0] _T_55847; // @[Modules.scala 78:156:@2162.4]
  wire [10:0] buffer_0_748; // @[Modules.scala 78:156:@2163.4]
  wire [11:0] _T_55849; // @[Modules.scala 78:156:@2165.4]
  wire [10:0] _T_55850; // @[Modules.scala 78:156:@2166.4]
  wire [10:0] buffer_0_749; // @[Modules.scala 78:156:@2167.4]
  wire [11:0] _T_55852; // @[Modules.scala 78:156:@2169.4]
  wire [10:0] _T_55853; // @[Modules.scala 78:156:@2170.4]
  wire [10:0] buffer_0_750; // @[Modules.scala 78:156:@2171.4]
  wire [11:0] _T_55855; // @[Modules.scala 78:156:@2173.4]
  wire [10:0] _T_55856; // @[Modules.scala 78:156:@2174.4]
  wire [10:0] buffer_0_751; // @[Modules.scala 78:156:@2175.4]
  wire [11:0] _T_55858; // @[Modules.scala 78:156:@2177.4]
  wire [10:0] _T_55859; // @[Modules.scala 78:156:@2178.4]
  wire [10:0] buffer_0_752; // @[Modules.scala 78:156:@2179.4]
  wire [11:0] _T_55861; // @[Modules.scala 78:156:@2181.4]
  wire [10:0] _T_55862; // @[Modules.scala 78:156:@2182.4]
  wire [10:0] buffer_0_753; // @[Modules.scala 78:156:@2183.4]
  wire [11:0] _T_55864; // @[Modules.scala 78:156:@2185.4]
  wire [10:0] _T_55865; // @[Modules.scala 78:156:@2186.4]
  wire [10:0] buffer_0_754; // @[Modules.scala 78:156:@2187.4]
  wire [11:0] _T_55867; // @[Modules.scala 78:156:@2189.4]
  wire [10:0] _T_55868; // @[Modules.scala 78:156:@2190.4]
  wire [10:0] buffer_0_755; // @[Modules.scala 78:156:@2191.4]
  wire [11:0] _T_55870; // @[Modules.scala 78:156:@2193.4]
  wire [10:0] _T_55871; // @[Modules.scala 78:156:@2194.4]
  wire [10:0] buffer_0_756; // @[Modules.scala 78:156:@2195.4]
  wire [11:0] _T_55873; // @[Modules.scala 78:156:@2197.4]
  wire [10:0] _T_55874; // @[Modules.scala 78:156:@2198.4]
  wire [10:0] buffer_0_757; // @[Modules.scala 78:156:@2199.4]
  wire [11:0] _T_55876; // @[Modules.scala 78:156:@2201.4]
  wire [10:0] _T_55877; // @[Modules.scala 78:156:@2202.4]
  wire [10:0] buffer_0_758; // @[Modules.scala 78:156:@2203.4]
  wire [11:0] _T_55879; // @[Modules.scala 78:156:@2205.4]
  wire [10:0] _T_55880; // @[Modules.scala 78:156:@2206.4]
  wire [10:0] buffer_0_759; // @[Modules.scala 78:156:@2207.4]
  wire [11:0] _T_55882; // @[Modules.scala 78:156:@2209.4]
  wire [10:0] _T_55883; // @[Modules.scala 78:156:@2210.4]
  wire [10:0] buffer_0_760; // @[Modules.scala 78:156:@2211.4]
  wire [11:0] _T_55885; // @[Modules.scala 78:156:@2213.4]
  wire [10:0] _T_55886; // @[Modules.scala 78:156:@2214.4]
  wire [10:0] buffer_0_761; // @[Modules.scala 78:156:@2215.4]
  wire [11:0] _T_55888; // @[Modules.scala 78:156:@2217.4]
  wire [10:0] _T_55889; // @[Modules.scala 78:156:@2218.4]
  wire [10:0] buffer_0_762; // @[Modules.scala 78:156:@2219.4]
  wire [11:0] _T_55891; // @[Modules.scala 78:156:@2221.4]
  wire [10:0] _T_55892; // @[Modules.scala 78:156:@2222.4]
  wire [10:0] buffer_0_763; // @[Modules.scala 78:156:@2223.4]
  wire [11:0] _T_55894; // @[Modules.scala 78:156:@2225.4]
  wire [10:0] _T_55895; // @[Modules.scala 78:156:@2226.4]
  wire [10:0] buffer_0_764; // @[Modules.scala 78:156:@2227.4]
  wire [11:0] _T_55897; // @[Modules.scala 78:156:@2229.4]
  wire [10:0] _T_55898; // @[Modules.scala 78:156:@2230.4]
  wire [10:0] buffer_0_765; // @[Modules.scala 78:156:@2231.4]
  wire [11:0] _T_55900; // @[Modules.scala 78:156:@2233.4]
  wire [10:0] _T_55901; // @[Modules.scala 78:156:@2234.4]
  wire [10:0] buffer_0_766; // @[Modules.scala 78:156:@2235.4]
  wire [11:0] _T_55903; // @[Modules.scala 78:156:@2237.4]
  wire [10:0] _T_55904; // @[Modules.scala 78:156:@2238.4]
  wire [10:0] buffer_0_767; // @[Modules.scala 78:156:@2239.4]
  wire [11:0] _T_55906; // @[Modules.scala 78:156:@2241.4]
  wire [10:0] _T_55907; // @[Modules.scala 78:156:@2242.4]
  wire [10:0] buffer_0_768; // @[Modules.scala 78:156:@2243.4]
  wire [11:0] _T_55909; // @[Modules.scala 78:156:@2245.4]
  wire [10:0] _T_55910; // @[Modules.scala 78:156:@2246.4]
  wire [10:0] buffer_0_769; // @[Modules.scala 78:156:@2247.4]
  wire [11:0] _T_55912; // @[Modules.scala 78:156:@2249.4]
  wire [10:0] _T_55913; // @[Modules.scala 78:156:@2250.4]
  wire [10:0] buffer_0_770; // @[Modules.scala 78:156:@2251.4]
  wire [11:0] _T_55915; // @[Modules.scala 78:156:@2253.4]
  wire [10:0] _T_55916; // @[Modules.scala 78:156:@2254.4]
  wire [10:0] buffer_0_771; // @[Modules.scala 78:156:@2255.4]
  wire [11:0] _T_55918; // @[Modules.scala 78:156:@2257.4]
  wire [10:0] _T_55919; // @[Modules.scala 78:156:@2258.4]
  wire [10:0] buffer_0_772; // @[Modules.scala 78:156:@2259.4]
  wire [11:0] _T_55921; // @[Modules.scala 78:156:@2261.4]
  wire [10:0] _T_55922; // @[Modules.scala 78:156:@2262.4]
  wire [10:0] buffer_0_773; // @[Modules.scala 78:156:@2263.4]
  wire [11:0] _T_55924; // @[Modules.scala 78:156:@2265.4]
  wire [10:0] _T_55925; // @[Modules.scala 78:156:@2266.4]
  wire [10:0] buffer_0_774; // @[Modules.scala 78:156:@2267.4]
  wire [11:0] _T_55927; // @[Modules.scala 78:156:@2269.4]
  wire [10:0] _T_55928; // @[Modules.scala 78:156:@2270.4]
  wire [10:0] buffer_0_775; // @[Modules.scala 78:156:@2271.4]
  wire [11:0] _T_55930; // @[Modules.scala 78:156:@2273.4]
  wire [10:0] _T_55931; // @[Modules.scala 78:156:@2274.4]
  wire [10:0] buffer_0_776; // @[Modules.scala 78:156:@2275.4]
  wire [11:0] _T_55933; // @[Modules.scala 78:156:@2277.4]
  wire [10:0] _T_55934; // @[Modules.scala 78:156:@2278.4]
  wire [10:0] buffer_0_777; // @[Modules.scala 78:156:@2279.4]
  wire [11:0] _T_55936; // @[Modules.scala 78:156:@2281.4]
  wire [10:0] _T_55937; // @[Modules.scala 78:156:@2282.4]
  wire [10:0] buffer_0_778; // @[Modules.scala 78:156:@2283.4]
  wire [11:0] _T_55939; // @[Modules.scala 78:156:@2285.4]
  wire [10:0] _T_55940; // @[Modules.scala 78:156:@2286.4]
  wire [10:0] buffer_0_779; // @[Modules.scala 78:156:@2287.4]
  wire [11:0] _T_55942; // @[Modules.scala 78:156:@2289.4]
  wire [10:0] _T_55943; // @[Modules.scala 78:156:@2290.4]
  wire [10:0] buffer_0_780; // @[Modules.scala 78:156:@2291.4]
  wire [11:0] _T_55945; // @[Modules.scala 78:156:@2293.4]
  wire [10:0] _T_55946; // @[Modules.scala 78:156:@2294.4]
  wire [10:0] buffer_0_781; // @[Modules.scala 78:156:@2295.4]
  wire [11:0] _T_55948; // @[Modules.scala 78:156:@2297.4]
  wire [10:0] _T_55949; // @[Modules.scala 78:156:@2298.4]
  wire [10:0] buffer_0_782; // @[Modules.scala 78:156:@2299.4]
  wire [11:0] _T_55951; // @[Modules.scala 78:156:@2301.4]
  wire [10:0] _T_55952; // @[Modules.scala 78:156:@2302.4]
  wire [10:0] buffer_0_783; // @[Modules.scala 78:156:@2303.4]
  wire [5:0] _T_55956; // @[Modules.scala 37:46:@2308.4]
  wire [4:0] _T_55957; // @[Modules.scala 37:46:@2309.4]
  wire [4:0] _T_55958; // @[Modules.scala 37:46:@2310.4]
  wire [5:0] _T_55959; // @[Modules.scala 37:46:@2312.4]
  wire [4:0] _T_55960; // @[Modules.scala 37:46:@2313.4]
  wire [4:0] _T_55961; // @[Modules.scala 37:46:@2314.4]
  wire [5:0] _T_55962; // @[Modules.scala 37:46:@2316.4]
  wire [4:0] _T_55963; // @[Modules.scala 37:46:@2317.4]
  wire [4:0] _T_55964; // @[Modules.scala 37:46:@2318.4]
  wire [5:0] _T_55966; // @[Modules.scala 37:46:@2321.4]
  wire [4:0] _T_55967; // @[Modules.scala 37:46:@2322.4]
  wire [4:0] _T_55968; // @[Modules.scala 37:46:@2323.4]
  wire [5:0] _T_55969; // @[Modules.scala 37:46:@2325.4]
  wire [4:0] _T_55970; // @[Modules.scala 37:46:@2326.4]
  wire [4:0] _T_55971; // @[Modules.scala 37:46:@2327.4]
  wire [5:0] _T_55975; // @[Modules.scala 37:46:@2336.4]
  wire [4:0] _T_55976; // @[Modules.scala 37:46:@2337.4]
  wire [4:0] _T_55977; // @[Modules.scala 37:46:@2338.4]
  wire [5:0] _T_55979; // @[Modules.scala 37:46:@2342.4]
  wire [4:0] _T_55980; // @[Modules.scala 37:46:@2343.4]
  wire [4:0] _T_55981; // @[Modules.scala 37:46:@2344.4]
  wire [5:0] _T_55985; // @[Modules.scala 37:46:@2350.4]
  wire [4:0] _T_55986; // @[Modules.scala 37:46:@2351.4]
  wire [4:0] _T_55987; // @[Modules.scala 37:46:@2352.4]
  wire [5:0] _T_55988; // @[Modules.scala 37:46:@2354.4]
  wire [4:0] _T_55989; // @[Modules.scala 37:46:@2355.4]
  wire [4:0] _T_55990; // @[Modules.scala 37:46:@2356.4]
  wire [5:0] _T_55991; // @[Modules.scala 37:46:@2358.4]
  wire [4:0] _T_55992; // @[Modules.scala 37:46:@2359.4]
  wire [4:0] _T_55993; // @[Modules.scala 37:46:@2360.4]
  wire [5:0] _T_55994; // @[Modules.scala 37:46:@2362.4]
  wire [4:0] _T_55995; // @[Modules.scala 37:46:@2363.4]
  wire [4:0] _T_55996; // @[Modules.scala 37:46:@2364.4]
  wire [5:0] _T_55997; // @[Modules.scala 37:46:@2366.4]
  wire [4:0] _T_55998; // @[Modules.scala 37:46:@2367.4]
  wire [4:0] _T_55999; // @[Modules.scala 37:46:@2368.4]
  wire [5:0] _T_56000; // @[Modules.scala 37:46:@2371.4]
  wire [4:0] _T_56001; // @[Modules.scala 37:46:@2372.4]
  wire [4:0] _T_56002; // @[Modules.scala 37:46:@2373.4]
  wire [5:0] _T_56003; // @[Modules.scala 37:46:@2375.4]
  wire [4:0] _T_56004; // @[Modules.scala 37:46:@2376.4]
  wire [4:0] _T_56005; // @[Modules.scala 37:46:@2377.4]
  wire [5:0] _T_56006; // @[Modules.scala 37:46:@2379.4]
  wire [4:0] _T_56007; // @[Modules.scala 37:46:@2380.4]
  wire [4:0] _T_56008; // @[Modules.scala 37:46:@2381.4]
  wire [5:0] _T_56009; // @[Modules.scala 37:46:@2386.4]
  wire [4:0] _T_56010; // @[Modules.scala 37:46:@2387.4]
  wire [4:0] _T_56011; // @[Modules.scala 37:46:@2388.4]
  wire [5:0] _T_56012; // @[Modules.scala 37:46:@2390.4]
  wire [4:0] _T_56013; // @[Modules.scala 37:46:@2391.4]
  wire [4:0] _T_56014; // @[Modules.scala 37:46:@2392.4]
  wire [5:0] _T_56015; // @[Modules.scala 37:46:@2394.4]
  wire [4:0] _T_56016; // @[Modules.scala 37:46:@2395.4]
  wire [4:0] _T_56017; // @[Modules.scala 37:46:@2396.4]
  wire [5:0] _T_56018; // @[Modules.scala 37:46:@2398.4]
  wire [4:0] _T_56019; // @[Modules.scala 37:46:@2399.4]
  wire [4:0] _T_56020; // @[Modules.scala 37:46:@2400.4]
  wire [5:0] _T_56021; // @[Modules.scala 37:46:@2402.4]
  wire [4:0] _T_56022; // @[Modules.scala 37:46:@2403.4]
  wire [4:0] _T_56023; // @[Modules.scala 37:46:@2404.4]
  wire [5:0] _T_56024; // @[Modules.scala 37:46:@2406.4]
  wire [4:0] _T_56025; // @[Modules.scala 37:46:@2407.4]
  wire [4:0] _T_56026; // @[Modules.scala 37:46:@2408.4]
  wire [5:0] _T_56027; // @[Modules.scala 37:46:@2410.4]
  wire [4:0] _T_56028; // @[Modules.scala 37:46:@2411.4]
  wire [4:0] _T_56029; // @[Modules.scala 37:46:@2412.4]
  wire [5:0] _T_56030; // @[Modules.scala 37:46:@2414.4]
  wire [4:0] _T_56031; // @[Modules.scala 37:46:@2415.4]
  wire [4:0] _T_56032; // @[Modules.scala 37:46:@2416.4]
  wire [5:0] _T_56033; // @[Modules.scala 37:46:@2418.4]
  wire [4:0] _T_56034; // @[Modules.scala 37:46:@2419.4]
  wire [4:0] _T_56035; // @[Modules.scala 37:46:@2420.4]
  wire [5:0] _T_56036; // @[Modules.scala 37:46:@2422.4]
  wire [4:0] _T_56037; // @[Modules.scala 37:46:@2423.4]
  wire [4:0] _T_56038; // @[Modules.scala 37:46:@2424.4]
  wire [5:0] _T_56042; // @[Modules.scala 37:46:@2430.4]
  wire [4:0] _T_56043; // @[Modules.scala 37:46:@2431.4]
  wire [4:0] _T_56044; // @[Modules.scala 37:46:@2432.4]
  wire [5:0] _T_56052; // @[Modules.scala 37:46:@2445.4]
  wire [4:0] _T_56053; // @[Modules.scala 37:46:@2446.4]
  wire [4:0] _T_56054; // @[Modules.scala 37:46:@2447.4]
  wire [5:0] _T_56058; // @[Modules.scala 37:46:@2453.4]
  wire [4:0] _T_56059; // @[Modules.scala 37:46:@2454.4]
  wire [4:0] _T_56060; // @[Modules.scala 37:46:@2455.4]
  wire [5:0] _T_56076; // @[Modules.scala 37:46:@2477.4]
  wire [4:0] _T_56077; // @[Modules.scala 37:46:@2478.4]
  wire [4:0] _T_56078; // @[Modules.scala 37:46:@2479.4]
  wire [5:0] _T_56087; // @[Modules.scala 37:46:@2493.4]
  wire [4:0] _T_56088; // @[Modules.scala 37:46:@2494.4]
  wire [4:0] _T_56089; // @[Modules.scala 37:46:@2495.4]
  wire [5:0] _T_56090; // @[Modules.scala 37:46:@2497.4]
  wire [4:0] _T_56091; // @[Modules.scala 37:46:@2498.4]
  wire [4:0] _T_56092; // @[Modules.scala 37:46:@2499.4]
  wire [5:0] _T_56096; // @[Modules.scala 37:46:@2506.4]
  wire [4:0] _T_56097; // @[Modules.scala 37:46:@2507.4]
  wire [4:0] _T_56098; // @[Modules.scala 37:46:@2508.4]
  wire [5:0] _T_56106; // @[Modules.scala 37:46:@2524.4]
  wire [4:0] _T_56107; // @[Modules.scala 37:46:@2525.4]
  wire [4:0] _T_56108; // @[Modules.scala 37:46:@2526.4]
  wire [5:0] _T_56109; // @[Modules.scala 37:46:@2529.4]
  wire [4:0] _T_56110; // @[Modules.scala 37:46:@2530.4]
  wire [4:0] _T_56111; // @[Modules.scala 37:46:@2531.4]
  wire [5:0] _T_56112; // @[Modules.scala 37:46:@2534.4]
  wire [4:0] _T_56113; // @[Modules.scala 37:46:@2535.4]
  wire [4:0] _T_56114; // @[Modules.scala 37:46:@2536.4]
  wire [5:0] _T_56115; // @[Modules.scala 37:46:@2538.4]
  wire [4:0] _T_56116; // @[Modules.scala 37:46:@2539.4]
  wire [4:0] _T_56117; // @[Modules.scala 37:46:@2540.4]
  wire [5:0] _T_56123; // @[Modules.scala 37:46:@2554.4]
  wire [4:0] _T_56124; // @[Modules.scala 37:46:@2555.4]
  wire [4:0] _T_56125; // @[Modules.scala 37:46:@2556.4]
  wire [5:0] _T_56126; // @[Modules.scala 37:46:@2560.4]
  wire [4:0] _T_56127; // @[Modules.scala 37:46:@2561.4]
  wire [4:0] _T_56128; // @[Modules.scala 37:46:@2562.4]
  wire [5:0] _T_56132; // @[Modules.scala 37:46:@2575.4]
  wire [4:0] _T_56133; // @[Modules.scala 37:46:@2576.4]
  wire [4:0] _T_56134; // @[Modules.scala 37:46:@2577.4]
  wire [5:0] _T_56135; // @[Modules.scala 37:46:@2580.4]
  wire [4:0] _T_56136; // @[Modules.scala 37:46:@2581.4]
  wire [4:0] _T_56137; // @[Modules.scala 37:46:@2582.4]
  wire [5:0] _T_56145; // @[Modules.scala 37:46:@2591.4]
  wire [4:0] _T_56146; // @[Modules.scala 37:46:@2592.4]
  wire [4:0] _T_56147; // @[Modules.scala 37:46:@2593.4]
  wire [5:0] _T_56150; // @[Modules.scala 37:46:@2598.4]
  wire [4:0] _T_56151; // @[Modules.scala 37:46:@2599.4]
  wire [4:0] _T_56152; // @[Modules.scala 37:46:@2600.4]
  wire [5:0] _T_56153; // @[Modules.scala 37:46:@2602.4]
  wire [4:0] _T_56154; // @[Modules.scala 37:46:@2603.4]
  wire [4:0] _T_56155; // @[Modules.scala 37:46:@2604.4]
  wire [5:0] _T_56161; // @[Modules.scala 37:46:@2613.4]
  wire [4:0] _T_56162; // @[Modules.scala 37:46:@2614.4]
  wire [4:0] _T_56163; // @[Modules.scala 37:46:@2615.4]
  wire [5:0] _T_56167; // @[Modules.scala 37:46:@2621.4]
  wire [4:0] _T_56168; // @[Modules.scala 37:46:@2622.4]
  wire [4:0] _T_56169; // @[Modules.scala 37:46:@2623.4]
  wire [5:0] _T_56170; // @[Modules.scala 37:46:@2625.4]
  wire [4:0] _T_56171; // @[Modules.scala 37:46:@2626.4]
  wire [4:0] _T_56172; // @[Modules.scala 37:46:@2627.4]
  wire [5:0] _T_56176; // @[Modules.scala 37:46:@2635.4]
  wire [4:0] _T_56177; // @[Modules.scala 37:46:@2636.4]
  wire [4:0] _T_56178; // @[Modules.scala 37:46:@2637.4]
  wire [5:0] _T_56182; // @[Modules.scala 37:46:@2644.4]
  wire [4:0] _T_56183; // @[Modules.scala 37:46:@2645.4]
  wire [4:0] _T_56184; // @[Modules.scala 37:46:@2646.4]
  wire [5:0] _T_56185; // @[Modules.scala 37:46:@2648.4]
  wire [4:0] _T_56186; // @[Modules.scala 37:46:@2649.4]
  wire [4:0] _T_56187; // @[Modules.scala 37:46:@2650.4]
  wire [5:0] _T_56195; // @[Modules.scala 37:46:@2661.4]
  wire [4:0] _T_56196; // @[Modules.scala 37:46:@2662.4]
  wire [4:0] _T_56197; // @[Modules.scala 37:46:@2663.4]
  wire [5:0] _T_56201; // @[Modules.scala 37:46:@2670.4]
  wire [4:0] _T_56202; // @[Modules.scala 37:46:@2671.4]
  wire [4:0] _T_56203; // @[Modules.scala 37:46:@2672.4]
  wire [5:0] _T_56204; // @[Modules.scala 37:46:@2674.4]
  wire [4:0] _T_56205; // @[Modules.scala 37:46:@2675.4]
  wire [4:0] _T_56206; // @[Modules.scala 37:46:@2676.4]
  wire [5:0] _T_56224; // @[Modules.scala 37:46:@2702.4]
  wire [4:0] _T_56225; // @[Modules.scala 37:46:@2703.4]
  wire [4:0] _T_56226; // @[Modules.scala 37:46:@2704.4]
  wire [5:0] _T_56249; // @[Modules.scala 37:46:@2736.4]
  wire [4:0] _T_56250; // @[Modules.scala 37:46:@2737.4]
  wire [4:0] _T_56251; // @[Modules.scala 37:46:@2738.4]
  wire [5:0] _T_56281; // @[Modules.scala 37:46:@2784.4]
  wire [4:0] _T_56282; // @[Modules.scala 37:46:@2785.4]
  wire [4:0] _T_56283; // @[Modules.scala 37:46:@2786.4]
  wire [5:0] _T_56284; // @[Modules.scala 37:46:@2788.4]
  wire [4:0] _T_56285; // @[Modules.scala 37:46:@2789.4]
  wire [4:0] _T_56286; // @[Modules.scala 37:46:@2790.4]
  wire [5:0] _T_56288; // @[Modules.scala 37:46:@2795.4]
  wire [4:0] _T_56289; // @[Modules.scala 37:46:@2796.4]
  wire [4:0] _T_56290; // @[Modules.scala 37:46:@2797.4]
  wire [5:0] _T_56296; // @[Modules.scala 37:46:@2807.4]
  wire [4:0] _T_56297; // @[Modules.scala 37:46:@2808.4]
  wire [4:0] _T_56298; // @[Modules.scala 37:46:@2809.4]
  wire [5:0] _T_56299; // @[Modules.scala 37:46:@2811.4]
  wire [4:0] _T_56300; // @[Modules.scala 37:46:@2812.4]
  wire [4:0] _T_56301; // @[Modules.scala 37:46:@2813.4]
  wire [5:0] _T_56303; // @[Modules.scala 37:46:@2818.4]
  wire [4:0] _T_56304; // @[Modules.scala 37:46:@2819.4]
  wire [4:0] _T_56305; // @[Modules.scala 37:46:@2820.4]
  wire [5:0] _T_56315; // @[Modules.scala 37:46:@2832.4]
  wire [4:0] _T_56316; // @[Modules.scala 37:46:@2833.4]
  wire [4:0] _T_56317; // @[Modules.scala 37:46:@2834.4]
  wire [5:0] _T_56318; // @[Modules.scala 37:46:@2836.4]
  wire [4:0] _T_56319; // @[Modules.scala 37:46:@2837.4]
  wire [4:0] _T_56320; // @[Modules.scala 37:46:@2838.4]
  wire [5:0] _T_56326; // @[Modules.scala 37:46:@2847.4]
  wire [4:0] _T_56327; // @[Modules.scala 37:46:@2848.4]
  wire [4:0] _T_56328; // @[Modules.scala 37:46:@2849.4]
  wire [5:0] _T_56329; // @[Modules.scala 37:46:@2852.4]
  wire [4:0] _T_56330; // @[Modules.scala 37:46:@2853.4]
  wire [4:0] _T_56331; // @[Modules.scala 37:46:@2854.4]
  wire [5:0] _T_56338; // @[Modules.scala 37:46:@2863.4]
  wire [4:0] _T_56339; // @[Modules.scala 37:46:@2864.4]
  wire [4:0] _T_56340; // @[Modules.scala 37:46:@2865.4]
  wire [5:0] _T_56341; // @[Modules.scala 37:46:@2867.4]
  wire [4:0] _T_56342; // @[Modules.scala 37:46:@2868.4]
  wire [4:0] _T_56343; // @[Modules.scala 37:46:@2869.4]
  wire [5:0] _T_56344; // @[Modules.scala 37:46:@2871.4]
  wire [4:0] _T_56345; // @[Modules.scala 37:46:@2872.4]
  wire [4:0] _T_56346; // @[Modules.scala 37:46:@2873.4]
  wire [5:0] _T_56349; // @[Modules.scala 37:46:@2878.4]
  wire [4:0] _T_56350; // @[Modules.scala 37:46:@2879.4]
  wire [4:0] _T_56351; // @[Modules.scala 37:46:@2880.4]
  wire [5:0] _T_56352; // @[Modules.scala 37:46:@2882.4]
  wire [4:0] _T_56353; // @[Modules.scala 37:46:@2883.4]
  wire [4:0] _T_56354; // @[Modules.scala 37:46:@2884.4]
  wire [5:0] _T_56355; // @[Modules.scala 37:46:@2886.4]
  wire [4:0] _T_56356; // @[Modules.scala 37:46:@2887.4]
  wire [4:0] _T_56357; // @[Modules.scala 37:46:@2888.4]
  wire [5:0] _T_56358; // @[Modules.scala 37:46:@2890.4]
  wire [4:0] _T_56359; // @[Modules.scala 37:46:@2891.4]
  wire [4:0] _T_56360; // @[Modules.scala 37:46:@2892.4]
  wire [5:0] _T_56361; // @[Modules.scala 37:46:@2894.4]
  wire [4:0] _T_56362; // @[Modules.scala 37:46:@2895.4]
  wire [4:0] _T_56363; // @[Modules.scala 37:46:@2896.4]
  wire [5:0] _T_56364; // @[Modules.scala 37:46:@2898.4]
  wire [4:0] _T_56365; // @[Modules.scala 37:46:@2899.4]
  wire [4:0] _T_56366; // @[Modules.scala 37:46:@2900.4]
  wire [5:0] _T_56367; // @[Modules.scala 37:46:@2902.4]
  wire [4:0] _T_56368; // @[Modules.scala 37:46:@2903.4]
  wire [4:0] _T_56369; // @[Modules.scala 37:46:@2904.4]
  wire [5:0] _T_56370; // @[Modules.scala 37:46:@2907.4]
  wire [4:0] _T_56371; // @[Modules.scala 37:46:@2908.4]
  wire [4:0] _T_56372; // @[Modules.scala 37:46:@2909.4]
  wire [5:0] _T_56373; // @[Modules.scala 37:46:@2911.4]
  wire [4:0] _T_56374; // @[Modules.scala 37:46:@2912.4]
  wire [4:0] _T_56375; // @[Modules.scala 37:46:@2913.4]
  wire [5:0] _T_56378; // @[Modules.scala 37:46:@2920.4]
  wire [4:0] _T_56379; // @[Modules.scala 37:46:@2921.4]
  wire [4:0] _T_56380; // @[Modules.scala 37:46:@2922.4]
  wire [5:0] _T_56381; // @[Modules.scala 37:46:@2924.4]
  wire [4:0] _T_56382; // @[Modules.scala 37:46:@2925.4]
  wire [4:0] _T_56383; // @[Modules.scala 37:46:@2926.4]
  wire [5:0] _T_56384; // @[Modules.scala 37:46:@2929.4]
  wire [4:0] _T_56385; // @[Modules.scala 37:46:@2930.4]
  wire [4:0] _T_56386; // @[Modules.scala 37:46:@2931.4]
  wire [5:0] _T_56387; // @[Modules.scala 37:46:@2933.4]
  wire [4:0] _T_56388; // @[Modules.scala 37:46:@2934.4]
  wire [4:0] _T_56389; // @[Modules.scala 37:46:@2935.4]
  wire [5:0] _T_56390; // @[Modules.scala 37:46:@2937.4]
  wire [4:0] _T_56391; // @[Modules.scala 37:46:@2938.4]
  wire [4:0] _T_56392; // @[Modules.scala 37:46:@2939.4]
  wire [5:0] _T_56393; // @[Modules.scala 37:46:@2941.4]
  wire [4:0] _T_56394; // @[Modules.scala 37:46:@2942.4]
  wire [4:0] _T_56395; // @[Modules.scala 37:46:@2943.4]
  wire [5:0] _T_56396; // @[Modules.scala 37:46:@2946.4]
  wire [4:0] _T_56397; // @[Modules.scala 37:46:@2947.4]
  wire [4:0] _T_56398; // @[Modules.scala 37:46:@2948.4]
  wire [5:0] _T_56401; // @[Modules.scala 37:46:@2955.4]
  wire [4:0] _T_56402; // @[Modules.scala 37:46:@2956.4]
  wire [4:0] _T_56403; // @[Modules.scala 37:46:@2957.4]
  wire [5:0] _T_56404; // @[Modules.scala 37:46:@2959.4]
  wire [4:0] _T_56405; // @[Modules.scala 37:46:@2960.4]
  wire [4:0] _T_56406; // @[Modules.scala 37:46:@2961.4]
  wire [5:0] _T_56407; // @[Modules.scala 37:46:@2965.4]
  wire [4:0] _T_56408; // @[Modules.scala 37:46:@2966.4]
  wire [4:0] _T_56409; // @[Modules.scala 37:46:@2967.4]
  wire [5:0] _T_56413; // @[Modules.scala 37:46:@2973.4]
  wire [4:0] _T_56414; // @[Modules.scala 37:46:@2974.4]
  wire [4:0] _T_56415; // @[Modules.scala 37:46:@2975.4]
  wire [5:0] _T_56430; // @[Modules.scala 37:46:@2996.4]
  wire [4:0] _T_56431; // @[Modules.scala 37:46:@2997.4]
  wire [4:0] _T_56432; // @[Modules.scala 37:46:@2998.4]
  wire [5:0] _T_56433; // @[Modules.scala 37:46:@3000.4]
  wire [4:0] _T_56434; // @[Modules.scala 37:46:@3001.4]
  wire [4:0] _T_56435; // @[Modules.scala 37:46:@3002.4]
  wire [5:0] _T_56436; // @[Modules.scala 37:46:@3004.4]
  wire [4:0] _T_56437; // @[Modules.scala 37:46:@3005.4]
  wire [4:0] _T_56438; // @[Modules.scala 37:46:@3006.4]
  wire [5:0] _T_56439; // @[Modules.scala 37:46:@3008.4]
  wire [4:0] _T_56440; // @[Modules.scala 37:46:@3009.4]
  wire [4:0] _T_56441; // @[Modules.scala 37:46:@3010.4]
  wire [5:0] _T_56442; // @[Modules.scala 37:46:@3012.4]
  wire [4:0] _T_56443; // @[Modules.scala 37:46:@3013.4]
  wire [4:0] _T_56444; // @[Modules.scala 37:46:@3014.4]
  wire [5:0] _T_56445; // @[Modules.scala 37:46:@3017.4]
  wire [4:0] _T_56446; // @[Modules.scala 37:46:@3018.4]
  wire [4:0] _T_56447; // @[Modules.scala 37:46:@3019.4]
  wire [5:0] _T_56449; // @[Modules.scala 37:46:@3023.4]
  wire [4:0] _T_56450; // @[Modules.scala 37:46:@3024.4]
  wire [4:0] _T_56451; // @[Modules.scala 37:46:@3025.4]
  wire [5:0] _T_56456; // @[Modules.scala 37:46:@3032.4]
  wire [4:0] _T_56457; // @[Modules.scala 37:46:@3033.4]
  wire [4:0] _T_56458; // @[Modules.scala 37:46:@3034.4]
  wire [5:0] _T_56459; // @[Modules.scala 37:46:@3036.4]
  wire [4:0] _T_56460; // @[Modules.scala 37:46:@3037.4]
  wire [4:0] _T_56461; // @[Modules.scala 37:46:@3038.4]
  wire [5:0] _T_56462; // @[Modules.scala 37:46:@3040.4]
  wire [4:0] _T_56463; // @[Modules.scala 37:46:@3041.4]
  wire [4:0] _T_56464; // @[Modules.scala 37:46:@3042.4]
  wire [5:0] _T_56465; // @[Modules.scala 37:46:@3044.4]
  wire [4:0] _T_56466; // @[Modules.scala 37:46:@3045.4]
  wire [4:0] _T_56467; // @[Modules.scala 37:46:@3046.4]
  wire [5:0] _T_56468; // @[Modules.scala 37:46:@3048.4]
  wire [4:0] _T_56469; // @[Modules.scala 37:46:@3049.4]
  wire [4:0] _T_56470; // @[Modules.scala 37:46:@3050.4]
  wire [5:0] _T_56471; // @[Modules.scala 37:46:@3052.4]
  wire [4:0] _T_56472; // @[Modules.scala 37:46:@3053.4]
  wire [4:0] _T_56473; // @[Modules.scala 37:46:@3054.4]
  wire [5:0] _T_56475; // @[Modules.scala 37:46:@3057.4]
  wire [4:0] _T_56476; // @[Modules.scala 37:46:@3058.4]
  wire [4:0] _T_56477; // @[Modules.scala 37:46:@3059.4]
  wire [5:0] _T_56483; // @[Modules.scala 37:46:@3066.4]
  wire [4:0] _T_56484; // @[Modules.scala 37:46:@3067.4]
  wire [4:0] _T_56485; // @[Modules.scala 37:46:@3068.4]
  wire [5:0] _T_56492; // @[Modules.scala 37:46:@3079.4]
  wire [4:0] _T_56493; // @[Modules.scala 37:46:@3080.4]
  wire [4:0] _T_56494; // @[Modules.scala 37:46:@3081.4]
  wire [5:0] _T_56495; // @[Modules.scala 37:46:@3083.4]
  wire [4:0] _T_56496; // @[Modules.scala 37:46:@3084.4]
  wire [4:0] _T_56497; // @[Modules.scala 37:46:@3085.4]
  wire [5:0] _T_56500; // @[Modules.scala 37:46:@3094.4]
  wire [4:0] _T_56501; // @[Modules.scala 37:46:@3095.4]
  wire [4:0] _T_56502; // @[Modules.scala 37:46:@3096.4]
  wire [5:0] _T_56503; // @[Modules.scala 37:46:@3098.4]
  wire [4:0] _T_56504; // @[Modules.scala 37:46:@3099.4]
  wire [4:0] _T_56505; // @[Modules.scala 37:46:@3100.4]
  wire [5:0] _T_56519; // @[Modules.scala 37:46:@3121.4]
  wire [4:0] _T_56520; // @[Modules.scala 37:46:@3122.4]
  wire [4:0] _T_56521; // @[Modules.scala 37:46:@3123.4]
  wire [5:0] _T_56541; // @[Modules.scala 37:46:@3150.4]
  wire [4:0] _T_56542; // @[Modules.scala 37:46:@3151.4]
  wire [4:0] _T_56543; // @[Modules.scala 37:46:@3152.4]
  wire [5:0] _T_56544; // @[Modules.scala 37:46:@3154.4]
  wire [4:0] _T_56545; // @[Modules.scala 37:46:@3155.4]
  wire [4:0] _T_56546; // @[Modules.scala 37:46:@3156.4]
  wire [5:0] _T_56547; // @[Modules.scala 37:46:@3158.4]
  wire [4:0] _T_56548; // @[Modules.scala 37:46:@3159.4]
  wire [4:0] _T_56549; // @[Modules.scala 37:46:@3160.4]
  wire [5:0] _T_56551; // @[Modules.scala 37:46:@3163.4]
  wire [4:0] _T_56552; // @[Modules.scala 37:46:@3164.4]
  wire [4:0] _T_56553; // @[Modules.scala 37:46:@3165.4]
  wire [10:0] buffer_1_2; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_3; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56564; // @[Modules.scala 65:57:@3179.4]
  wire [10:0] _T_56565; // @[Modules.scala 65:57:@3180.4]
  wire [10:0] buffer_1_393; // @[Modules.scala 65:57:@3181.4]
  wire [10:0] buffer_1_4; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56567; // @[Modules.scala 65:57:@3183.4]
  wire [10:0] _T_56568; // @[Modules.scala 65:57:@3184.4]
  wire [10:0] buffer_1_394; // @[Modules.scala 65:57:@3185.4]
  wire [10:0] buffer_1_6; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_7; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56570; // @[Modules.scala 65:57:@3187.4]
  wire [10:0] _T_56571; // @[Modules.scala 65:57:@3188.4]
  wire [10:0] buffer_1_395; // @[Modules.scala 65:57:@3189.4]
  wire [10:0] buffer_1_8; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56573; // @[Modules.scala 65:57:@3191.4]
  wire [10:0] _T_56574; // @[Modules.scala 65:57:@3192.4]
  wire [10:0] buffer_1_396; // @[Modules.scala 65:57:@3193.4]
  wire [10:0] buffer_1_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56576; // @[Modules.scala 65:57:@3195.4]
  wire [10:0] _T_56577; // @[Modules.scala 65:57:@3196.4]
  wire [10:0] buffer_1_397; // @[Modules.scala 65:57:@3197.4]
  wire [10:0] buffer_1_12; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56579; // @[Modules.scala 65:57:@3199.4]
  wire [10:0] _T_56580; // @[Modules.scala 65:57:@3200.4]
  wire [10:0] buffer_1_398; // @[Modules.scala 65:57:@3201.4]
  wire [10:0] buffer_1_14; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56582; // @[Modules.scala 65:57:@3203.4]
  wire [10:0] _T_56583; // @[Modules.scala 65:57:@3204.4]
  wire [10:0] buffer_1_399; // @[Modules.scala 65:57:@3205.4]
  wire [10:0] buffer_1_17; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56585; // @[Modules.scala 65:57:@3207.4]
  wire [10:0] _T_56586; // @[Modules.scala 65:57:@3208.4]
  wire [10:0] buffer_1_400; // @[Modules.scala 65:57:@3209.4]
  wire [10:0] buffer_1_18; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_19; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56588; // @[Modules.scala 65:57:@3211.4]
  wire [10:0] _T_56589; // @[Modules.scala 65:57:@3212.4]
  wire [10:0] buffer_1_401; // @[Modules.scala 65:57:@3213.4]
  wire [10:0] buffer_1_20; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_21; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56591; // @[Modules.scala 65:57:@3215.4]
  wire [10:0] _T_56592; // @[Modules.scala 65:57:@3216.4]
  wire [10:0] buffer_1_402; // @[Modules.scala 65:57:@3217.4]
  wire [10:0] buffer_1_22; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_23; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56594; // @[Modules.scala 65:57:@3219.4]
  wire [10:0] _T_56595; // @[Modules.scala 65:57:@3220.4]
  wire [10:0] buffer_1_403; // @[Modules.scala 65:57:@3221.4]
  wire [10:0] buffer_1_24; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_25; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56597; // @[Modules.scala 65:57:@3223.4]
  wire [10:0] _T_56598; // @[Modules.scala 65:57:@3224.4]
  wire [10:0] buffer_1_404; // @[Modules.scala 65:57:@3225.4]
  wire [10:0] buffer_1_26; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56600; // @[Modules.scala 65:57:@3227.4]
  wire [10:0] _T_56601; // @[Modules.scala 65:57:@3228.4]
  wire [10:0] buffer_1_405; // @[Modules.scala 65:57:@3229.4]
  wire [10:0] buffer_1_28; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56603; // @[Modules.scala 65:57:@3231.4]
  wire [10:0] _T_56604; // @[Modules.scala 65:57:@3232.4]
  wire [10:0] buffer_1_406; // @[Modules.scala 65:57:@3233.4]
  wire [10:0] buffer_1_30; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_31; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56606; // @[Modules.scala 65:57:@3235.4]
  wire [10:0] _T_56607; // @[Modules.scala 65:57:@3236.4]
  wire [10:0] buffer_1_407; // @[Modules.scala 65:57:@3237.4]
  wire [10:0] buffer_1_32; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_33; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56609; // @[Modules.scala 65:57:@3239.4]
  wire [10:0] _T_56610; // @[Modules.scala 65:57:@3240.4]
  wire [10:0] buffer_1_408; // @[Modules.scala 65:57:@3241.4]
  wire [10:0] buffer_1_34; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56612; // @[Modules.scala 65:57:@3243.4]
  wire [10:0] _T_56613; // @[Modules.scala 65:57:@3244.4]
  wire [10:0] buffer_1_409; // @[Modules.scala 65:57:@3245.4]
  wire [10:0] buffer_1_36; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_37; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56615; // @[Modules.scala 65:57:@3247.4]
  wire [10:0] _T_56616; // @[Modules.scala 65:57:@3248.4]
  wire [10:0] buffer_1_410; // @[Modules.scala 65:57:@3249.4]
  wire [10:0] buffer_1_38; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56618; // @[Modules.scala 65:57:@3251.4]
  wire [10:0] _T_56619; // @[Modules.scala 65:57:@3252.4]
  wire [10:0] buffer_1_411; // @[Modules.scala 65:57:@3253.4]
  wire [10:0] buffer_1_40; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56621; // @[Modules.scala 65:57:@3255.4]
  wire [10:0] _T_56622; // @[Modules.scala 65:57:@3256.4]
  wire [10:0] buffer_1_412; // @[Modules.scala 65:57:@3257.4]
  wire [10:0] buffer_1_42; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56624; // @[Modules.scala 65:57:@3259.4]
  wire [10:0] _T_56625; // @[Modules.scala 65:57:@3260.4]
  wire [10:0] buffer_1_413; // @[Modules.scala 65:57:@3261.4]
  wire [10:0] buffer_1_46; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56630; // @[Modules.scala 65:57:@3267.4]
  wire [10:0] _T_56631; // @[Modules.scala 65:57:@3268.4]
  wire [10:0] buffer_1_415; // @[Modules.scala 65:57:@3269.4]
  wire [10:0] buffer_1_48; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56633; // @[Modules.scala 65:57:@3271.4]
  wire [10:0] _T_56634; // @[Modules.scala 65:57:@3272.4]
  wire [10:0] buffer_1_416; // @[Modules.scala 65:57:@3273.4]
  wire [10:0] buffer_1_54; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56642; // @[Modules.scala 65:57:@3283.4]
  wire [10:0] _T_56643; // @[Modules.scala 65:57:@3284.4]
  wire [10:0] buffer_1_419; // @[Modules.scala 65:57:@3285.4]
  wire [10:0] buffer_1_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56645; // @[Modules.scala 65:57:@3287.4]
  wire [10:0] _T_56646; // @[Modules.scala 65:57:@3288.4]
  wire [10:0] buffer_1_420; // @[Modules.scala 65:57:@3289.4]
  wire [11:0] _T_56648; // @[Modules.scala 65:57:@3291.4]
  wire [10:0] _T_56649; // @[Modules.scala 65:57:@3292.4]
  wire [10:0] buffer_1_421; // @[Modules.scala 65:57:@3293.4]
  wire [10:0] buffer_1_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56654; // @[Modules.scala 65:57:@3299.4]
  wire [10:0] _T_56655; // @[Modules.scala 65:57:@3300.4]
  wire [10:0] buffer_1_423; // @[Modules.scala 65:57:@3301.4]
  wire [10:0] buffer_1_64; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_65; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56657; // @[Modules.scala 65:57:@3303.4]
  wire [10:0] _T_56658; // @[Modules.scala 65:57:@3304.4]
  wire [10:0] buffer_1_424; // @[Modules.scala 65:57:@3305.4]
  wire [10:0] buffer_1_66; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56660; // @[Modules.scala 65:57:@3307.4]
  wire [10:0] _T_56661; // @[Modules.scala 65:57:@3308.4]
  wire [10:0] buffer_1_425; // @[Modules.scala 65:57:@3309.4]
  wire [10:0] buffer_1_68; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56663; // @[Modules.scala 65:57:@3311.4]
  wire [10:0] _T_56664; // @[Modules.scala 65:57:@3312.4]
  wire [10:0] buffer_1_426; // @[Modules.scala 65:57:@3313.4]
  wire [10:0] buffer_1_70; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56666; // @[Modules.scala 65:57:@3315.4]
  wire [10:0] _T_56667; // @[Modules.scala 65:57:@3316.4]
  wire [10:0] buffer_1_427; // @[Modules.scala 65:57:@3317.4]
  wire [10:0] buffer_1_74; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56672; // @[Modules.scala 65:57:@3323.4]
  wire [10:0] _T_56673; // @[Modules.scala 65:57:@3324.4]
  wire [10:0] buffer_1_429; // @[Modules.scala 65:57:@3325.4]
  wire [10:0] buffer_1_78; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56678; // @[Modules.scala 65:57:@3331.4]
  wire [10:0] _T_56679; // @[Modules.scala 65:57:@3332.4]
  wire [10:0] buffer_1_431; // @[Modules.scala 65:57:@3333.4]
  wire [10:0] buffer_1_81; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56681; // @[Modules.scala 65:57:@3335.4]
  wire [10:0] _T_56682; // @[Modules.scala 65:57:@3336.4]
  wire [10:0] buffer_1_432; // @[Modules.scala 65:57:@3337.4]
  wire [10:0] buffer_1_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56684; // @[Modules.scala 65:57:@3339.4]
  wire [10:0] _T_56685; // @[Modules.scala 65:57:@3340.4]
  wire [10:0] buffer_1_433; // @[Modules.scala 65:57:@3341.4]
  wire [10:0] buffer_1_84; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56687; // @[Modules.scala 65:57:@3343.4]
  wire [10:0] _T_56688; // @[Modules.scala 65:57:@3344.4]
  wire [10:0] buffer_1_434; // @[Modules.scala 65:57:@3345.4]
  wire [10:0] buffer_1_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56690; // @[Modules.scala 65:57:@3347.4]
  wire [10:0] _T_56691; // @[Modules.scala 65:57:@3348.4]
  wire [10:0] buffer_1_435; // @[Modules.scala 65:57:@3349.4]
  wire [10:0] buffer_1_88; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56693; // @[Modules.scala 65:57:@3351.4]
  wire [10:0] _T_56694; // @[Modules.scala 65:57:@3352.4]
  wire [10:0] buffer_1_436; // @[Modules.scala 65:57:@3353.4]
  wire [10:0] buffer_1_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56696; // @[Modules.scala 65:57:@3355.4]
  wire [10:0] _T_56697; // @[Modules.scala 65:57:@3356.4]
  wire [10:0] buffer_1_437; // @[Modules.scala 65:57:@3357.4]
  wire [10:0] buffer_1_94; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56702; // @[Modules.scala 65:57:@3363.4]
  wire [10:0] _T_56703; // @[Modules.scala 65:57:@3364.4]
  wire [10:0] buffer_1_439; // @[Modules.scala 65:57:@3365.4]
  wire [10:0] buffer_1_96; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56705; // @[Modules.scala 65:57:@3367.4]
  wire [10:0] _T_56706; // @[Modules.scala 65:57:@3368.4]
  wire [10:0] buffer_1_440; // @[Modules.scala 65:57:@3369.4]
  wire [10:0] buffer_1_98; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56708; // @[Modules.scala 65:57:@3371.4]
  wire [10:0] _T_56709; // @[Modules.scala 65:57:@3372.4]
  wire [10:0] buffer_1_441; // @[Modules.scala 65:57:@3373.4]
  wire [10:0] buffer_1_100; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56711; // @[Modules.scala 65:57:@3375.4]
  wire [10:0] _T_56712; // @[Modules.scala 65:57:@3376.4]
  wire [10:0] buffer_1_442; // @[Modules.scala 65:57:@3377.4]
  wire [10:0] buffer_1_102; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56714; // @[Modules.scala 65:57:@3379.4]
  wire [10:0] _T_56715; // @[Modules.scala 65:57:@3380.4]
  wire [10:0] buffer_1_443; // @[Modules.scala 65:57:@3381.4]
  wire [10:0] buffer_1_104; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56717; // @[Modules.scala 65:57:@3383.4]
  wire [10:0] _T_56718; // @[Modules.scala 65:57:@3384.4]
  wire [10:0] buffer_1_444; // @[Modules.scala 65:57:@3385.4]
  wire [10:0] buffer_1_106; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56720; // @[Modules.scala 65:57:@3387.4]
  wire [10:0] _T_56721; // @[Modules.scala 65:57:@3388.4]
  wire [10:0] buffer_1_445; // @[Modules.scala 65:57:@3389.4]
  wire [10:0] buffer_1_108; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56723; // @[Modules.scala 65:57:@3391.4]
  wire [10:0] _T_56724; // @[Modules.scala 65:57:@3392.4]
  wire [10:0] buffer_1_446; // @[Modules.scala 65:57:@3393.4]
  wire [10:0] buffer_1_110; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56726; // @[Modules.scala 65:57:@3395.4]
  wire [10:0] _T_56727; // @[Modules.scala 65:57:@3396.4]
  wire [10:0] buffer_1_447; // @[Modules.scala 65:57:@3397.4]
  wire [10:0] buffer_1_112; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56729; // @[Modules.scala 65:57:@3399.4]
  wire [10:0] _T_56730; // @[Modules.scala 65:57:@3400.4]
  wire [10:0] buffer_1_448; // @[Modules.scala 65:57:@3401.4]
  wire [10:0] buffer_1_120; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56741; // @[Modules.scala 65:57:@3415.4]
  wire [10:0] _T_56742; // @[Modules.scala 65:57:@3416.4]
  wire [10:0] buffer_1_452; // @[Modules.scala 65:57:@3417.4]
  wire [10:0] buffer_1_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56744; // @[Modules.scala 65:57:@3419.4]
  wire [10:0] _T_56745; // @[Modules.scala 65:57:@3420.4]
  wire [10:0] buffer_1_453; // @[Modules.scala 65:57:@3421.4]
  wire [10:0] buffer_1_124; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_125; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56747; // @[Modules.scala 65:57:@3423.4]
  wire [10:0] _T_56748; // @[Modules.scala 65:57:@3424.4]
  wire [10:0] buffer_1_454; // @[Modules.scala 65:57:@3425.4]
  wire [10:0] buffer_1_126; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56750; // @[Modules.scala 65:57:@3427.4]
  wire [10:0] _T_56751; // @[Modules.scala 65:57:@3428.4]
  wire [10:0] buffer_1_455; // @[Modules.scala 65:57:@3429.4]
  wire [10:0] buffer_1_130; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56756; // @[Modules.scala 65:57:@3435.4]
  wire [10:0] _T_56757; // @[Modules.scala 65:57:@3436.4]
  wire [10:0] buffer_1_457; // @[Modules.scala 65:57:@3437.4]
  wire [10:0] buffer_1_133; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56759; // @[Modules.scala 65:57:@3439.4]
  wire [10:0] _T_56760; // @[Modules.scala 65:57:@3440.4]
  wire [10:0] buffer_1_458; // @[Modules.scala 65:57:@3441.4]
  wire [10:0] buffer_1_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56765; // @[Modules.scala 65:57:@3447.4]
  wire [10:0] _T_56766; // @[Modules.scala 65:57:@3448.4]
  wire [10:0] buffer_1_460; // @[Modules.scala 65:57:@3449.4]
  wire [10:0] buffer_1_138; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_139; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56768; // @[Modules.scala 65:57:@3451.4]
  wire [10:0] _T_56769; // @[Modules.scala 65:57:@3452.4]
  wire [10:0] buffer_1_461; // @[Modules.scala 65:57:@3453.4]
  wire [10:0] buffer_1_140; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56771; // @[Modules.scala 65:57:@3455.4]
  wire [10:0] _T_56772; // @[Modules.scala 65:57:@3456.4]
  wire [10:0] buffer_1_462; // @[Modules.scala 65:57:@3457.4]
  wire [10:0] buffer_1_146; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56780; // @[Modules.scala 65:57:@3467.4]
  wire [10:0] _T_56781; // @[Modules.scala 65:57:@3468.4]
  wire [10:0] buffer_1_465; // @[Modules.scala 65:57:@3469.4]
  wire [10:0] buffer_1_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56786; // @[Modules.scala 65:57:@3475.4]
  wire [10:0] _T_56787; // @[Modules.scala 65:57:@3476.4]
  wire [10:0] buffer_1_467; // @[Modules.scala 65:57:@3477.4]
  wire [10:0] buffer_1_152; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_153; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56789; // @[Modules.scala 65:57:@3479.4]
  wire [10:0] _T_56790; // @[Modules.scala 65:57:@3480.4]
  wire [10:0] buffer_1_468; // @[Modules.scala 65:57:@3481.4]
  wire [10:0] buffer_1_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56795; // @[Modules.scala 65:57:@3487.4]
  wire [10:0] _T_56796; // @[Modules.scala 65:57:@3488.4]
  wire [10:0] buffer_1_470; // @[Modules.scala 65:57:@3489.4]
  wire [11:0] _T_56798; // @[Modules.scala 65:57:@3491.4]
  wire [10:0] _T_56799; // @[Modules.scala 65:57:@3492.4]
  wire [10:0] buffer_1_471; // @[Modules.scala 65:57:@3493.4]
  wire [10:0] buffer_1_160; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56801; // @[Modules.scala 65:57:@3495.4]
  wire [10:0] _T_56802; // @[Modules.scala 65:57:@3496.4]
  wire [10:0] buffer_1_472; // @[Modules.scala 65:57:@3497.4]
  wire [10:0] buffer_1_165; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56807; // @[Modules.scala 65:57:@3503.4]
  wire [10:0] _T_56808; // @[Modules.scala 65:57:@3504.4]
  wire [10:0] buffer_1_474; // @[Modules.scala 65:57:@3505.4]
  wire [10:0] buffer_1_166; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56810; // @[Modules.scala 65:57:@3507.4]
  wire [10:0] _T_56811; // @[Modules.scala 65:57:@3508.4]
  wire [10:0] buffer_1_475; // @[Modules.scala 65:57:@3509.4]
  wire [11:0] _T_56822; // @[Modules.scala 65:57:@3523.4]
  wire [10:0] _T_56823; // @[Modules.scala 65:57:@3524.4]
  wire [10:0] buffer_1_479; // @[Modules.scala 65:57:@3525.4]
  wire [10:0] buffer_1_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56828; // @[Modules.scala 65:57:@3531.4]
  wire [10:0] _T_56829; // @[Modules.scala 65:57:@3532.4]
  wire [10:0] buffer_1_481; // @[Modules.scala 65:57:@3533.4]
  wire [10:0] buffer_1_180; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56831; // @[Modules.scala 65:57:@3535.4]
  wire [10:0] _T_56832; // @[Modules.scala 65:57:@3536.4]
  wire [10:0] buffer_1_482; // @[Modules.scala 65:57:@3537.4]
  wire [10:0] buffer_1_184; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56837; // @[Modules.scala 65:57:@3543.4]
  wire [10:0] _T_56838; // @[Modules.scala 65:57:@3544.4]
  wire [10:0] buffer_1_484; // @[Modules.scala 65:57:@3545.4]
  wire [11:0] _T_56843; // @[Modules.scala 65:57:@3551.4]
  wire [10:0] _T_56844; // @[Modules.scala 65:57:@3552.4]
  wire [10:0] buffer_1_486; // @[Modules.scala 65:57:@3553.4]
  wire [11:0] _T_56852; // @[Modules.scala 65:57:@3563.4]
  wire [10:0] _T_56853; // @[Modules.scala 65:57:@3564.4]
  wire [10:0] buffer_1_489; // @[Modules.scala 65:57:@3565.4]
  wire [10:0] buffer_1_196; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56855; // @[Modules.scala 65:57:@3567.4]
  wire [10:0] _T_56856; // @[Modules.scala 65:57:@3568.4]
  wire [10:0] buffer_1_490; // @[Modules.scala 65:57:@3569.4]
  wire [10:0] buffer_1_198; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56858; // @[Modules.scala 65:57:@3571.4]
  wire [10:0] _T_56859; // @[Modules.scala 65:57:@3572.4]
  wire [10:0] buffer_1_491; // @[Modules.scala 65:57:@3573.4]
  wire [10:0] buffer_1_202; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56864; // @[Modules.scala 65:57:@3579.4]
  wire [10:0] _T_56865; // @[Modules.scala 65:57:@3580.4]
  wire [10:0] buffer_1_493; // @[Modules.scala 65:57:@3581.4]
  wire [10:0] buffer_1_204; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56867; // @[Modules.scala 65:57:@3583.4]
  wire [10:0] _T_56868; // @[Modules.scala 65:57:@3584.4]
  wire [10:0] buffer_1_494; // @[Modules.scala 65:57:@3585.4]
  wire [11:0] _T_56873; // @[Modules.scala 65:57:@3591.4]
  wire [10:0] _T_56874; // @[Modules.scala 65:57:@3592.4]
  wire [10:0] buffer_1_496; // @[Modules.scala 65:57:@3593.4]
  wire [10:0] buffer_1_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56876; // @[Modules.scala 65:57:@3595.4]
  wire [10:0] _T_56877; // @[Modules.scala 65:57:@3596.4]
  wire [10:0] buffer_1_497; // @[Modules.scala 65:57:@3597.4]
  wire [11:0] _T_56879; // @[Modules.scala 65:57:@3599.4]
  wire [10:0] _T_56880; // @[Modules.scala 65:57:@3600.4]
  wire [10:0] buffer_1_498; // @[Modules.scala 65:57:@3601.4]
  wire [10:0] buffer_1_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56888; // @[Modules.scala 65:57:@3611.4]
  wire [10:0] _T_56889; // @[Modules.scala 65:57:@3612.4]
  wire [10:0] buffer_1_501; // @[Modules.scala 65:57:@3613.4]
  wire [10:0] buffer_1_220; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56891; // @[Modules.scala 65:57:@3615.4]
  wire [10:0] _T_56892; // @[Modules.scala 65:57:@3616.4]
  wire [10:0] buffer_1_502; // @[Modules.scala 65:57:@3617.4]
  wire [10:0] buffer_1_222; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56894; // @[Modules.scala 65:57:@3619.4]
  wire [10:0] _T_56895; // @[Modules.scala 65:57:@3620.4]
  wire [10:0] buffer_1_503; // @[Modules.scala 65:57:@3621.4]
  wire [10:0] buffer_1_224; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56897; // @[Modules.scala 65:57:@3623.4]
  wire [10:0] _T_56898; // @[Modules.scala 65:57:@3624.4]
  wire [10:0] buffer_1_504; // @[Modules.scala 65:57:@3625.4]
  wire [10:0] buffer_1_228; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56903; // @[Modules.scala 65:57:@3631.4]
  wire [10:0] _T_56904; // @[Modules.scala 65:57:@3632.4]
  wire [10:0] buffer_1_506; // @[Modules.scala 65:57:@3633.4]
  wire [10:0] buffer_1_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56909; // @[Modules.scala 65:57:@3639.4]
  wire [10:0] _T_56910; // @[Modules.scala 65:57:@3640.4]
  wire [10:0] buffer_1_508; // @[Modules.scala 65:57:@3641.4]
  wire [10:0] buffer_1_234; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56912; // @[Modules.scala 65:57:@3643.4]
  wire [10:0] _T_56913; // @[Modules.scala 65:57:@3644.4]
  wire [10:0] buffer_1_509; // @[Modules.scala 65:57:@3645.4]
  wire [10:0] buffer_1_236; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56915; // @[Modules.scala 65:57:@3647.4]
  wire [10:0] _T_56916; // @[Modules.scala 65:57:@3648.4]
  wire [10:0] buffer_1_510; // @[Modules.scala 65:57:@3649.4]
  wire [10:0] buffer_1_238; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56918; // @[Modules.scala 65:57:@3651.4]
  wire [10:0] _T_56919; // @[Modules.scala 65:57:@3652.4]
  wire [10:0] buffer_1_511; // @[Modules.scala 65:57:@3653.4]
  wire [10:0] buffer_1_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56930; // @[Modules.scala 65:57:@3667.4]
  wire [10:0] _T_56931; // @[Modules.scala 65:57:@3668.4]
  wire [10:0] buffer_1_515; // @[Modules.scala 65:57:@3669.4]
  wire [10:0] buffer_1_248; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56933; // @[Modules.scala 65:57:@3671.4]
  wire [10:0] _T_56934; // @[Modules.scala 65:57:@3672.4]
  wire [10:0] buffer_1_516; // @[Modules.scala 65:57:@3673.4]
  wire [10:0] buffer_1_252; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56939; // @[Modules.scala 65:57:@3679.4]
  wire [10:0] _T_56940; // @[Modules.scala 65:57:@3680.4]
  wire [10:0] buffer_1_518; // @[Modules.scala 65:57:@3681.4]
  wire [10:0] buffer_1_254; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56942; // @[Modules.scala 65:57:@3683.4]
  wire [10:0] _T_56943; // @[Modules.scala 65:57:@3684.4]
  wire [10:0] buffer_1_519; // @[Modules.scala 65:57:@3685.4]
  wire [11:0] _T_56945; // @[Modules.scala 65:57:@3687.4]
  wire [10:0] _T_56946; // @[Modules.scala 65:57:@3688.4]
  wire [10:0] buffer_1_520; // @[Modules.scala 65:57:@3689.4]
  wire [10:0] buffer_1_260; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_261; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56951; // @[Modules.scala 65:57:@3695.4]
  wire [10:0] _T_56952; // @[Modules.scala 65:57:@3696.4]
  wire [10:0] buffer_1_522; // @[Modules.scala 65:57:@3697.4]
  wire [10:0] buffer_1_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56954; // @[Modules.scala 65:57:@3699.4]
  wire [10:0] _T_56955; // @[Modules.scala 65:57:@3700.4]
  wire [10:0] buffer_1_523; // @[Modules.scala 65:57:@3701.4]
  wire [10:0] buffer_1_266; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_267; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56960; // @[Modules.scala 65:57:@3707.4]
  wire [10:0] _T_56961; // @[Modules.scala 65:57:@3708.4]
  wire [10:0] buffer_1_525; // @[Modules.scala 65:57:@3709.4]
  wire [10:0] buffer_1_268; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56963; // @[Modules.scala 65:57:@3711.4]
  wire [10:0] _T_56964; // @[Modules.scala 65:57:@3712.4]
  wire [10:0] buffer_1_526; // @[Modules.scala 65:57:@3713.4]
  wire [10:0] buffer_1_270; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_271; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56966; // @[Modules.scala 65:57:@3715.4]
  wire [10:0] _T_56967; // @[Modules.scala 65:57:@3716.4]
  wire [10:0] buffer_1_527; // @[Modules.scala 65:57:@3717.4]
  wire [10:0] buffer_1_272; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56969; // @[Modules.scala 65:57:@3719.4]
  wire [10:0] _T_56970; // @[Modules.scala 65:57:@3720.4]
  wire [10:0] buffer_1_528; // @[Modules.scala 65:57:@3721.4]
  wire [10:0] buffer_1_274; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56972; // @[Modules.scala 65:57:@3723.4]
  wire [10:0] _T_56973; // @[Modules.scala 65:57:@3724.4]
  wire [10:0] buffer_1_529; // @[Modules.scala 65:57:@3725.4]
  wire [10:0] buffer_1_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56975; // @[Modules.scala 65:57:@3727.4]
  wire [10:0] _T_56976; // @[Modules.scala 65:57:@3728.4]
  wire [10:0] buffer_1_530; // @[Modules.scala 65:57:@3729.4]
  wire [10:0] buffer_1_280; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56981; // @[Modules.scala 65:57:@3735.4]
  wire [10:0] _T_56982; // @[Modules.scala 65:57:@3736.4]
  wire [10:0] buffer_1_532; // @[Modules.scala 65:57:@3737.4]
  wire [10:0] buffer_1_282; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56984; // @[Modules.scala 65:57:@3739.4]
  wire [10:0] _T_56985; // @[Modules.scala 65:57:@3740.4]
  wire [10:0] buffer_1_533; // @[Modules.scala 65:57:@3741.4]
  wire [10:0] buffer_1_284; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_285; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56987; // @[Modules.scala 65:57:@3743.4]
  wire [10:0] _T_56988; // @[Modules.scala 65:57:@3744.4]
  wire [10:0] buffer_1_534; // @[Modules.scala 65:57:@3745.4]
  wire [10:0] buffer_1_286; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56990; // @[Modules.scala 65:57:@3747.4]
  wire [10:0] _T_56991; // @[Modules.scala 65:57:@3748.4]
  wire [10:0] buffer_1_535; // @[Modules.scala 65:57:@3749.4]
  wire [10:0] buffer_1_288; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56993; // @[Modules.scala 65:57:@3751.4]
  wire [10:0] _T_56994; // @[Modules.scala 65:57:@3752.4]
  wire [10:0] buffer_1_536; // @[Modules.scala 65:57:@3753.4]
  wire [10:0] buffer_1_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_56996; // @[Modules.scala 65:57:@3755.4]
  wire [10:0] _T_56997; // @[Modules.scala 65:57:@3756.4]
  wire [10:0] buffer_1_537; // @[Modules.scala 65:57:@3757.4]
  wire [11:0] _T_56999; // @[Modules.scala 65:57:@3759.4]
  wire [10:0] _T_57000; // @[Modules.scala 65:57:@3760.4]
  wire [10:0] buffer_1_538; // @[Modules.scala 65:57:@3761.4]
  wire [10:0] buffer_1_295; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57002; // @[Modules.scala 65:57:@3763.4]
  wire [10:0] _T_57003; // @[Modules.scala 65:57:@3764.4]
  wire [10:0] buffer_1_539; // @[Modules.scala 65:57:@3765.4]
  wire [10:0] buffer_1_296; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57005; // @[Modules.scala 65:57:@3767.4]
  wire [10:0] _T_57006; // @[Modules.scala 65:57:@3768.4]
  wire [10:0] buffer_1_540; // @[Modules.scala 65:57:@3769.4]
  wire [10:0] buffer_1_298; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57008; // @[Modules.scala 65:57:@3771.4]
  wire [10:0] _T_57009; // @[Modules.scala 65:57:@3772.4]
  wire [10:0] buffer_1_541; // @[Modules.scala 65:57:@3773.4]
  wire [10:0] buffer_1_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57011; // @[Modules.scala 65:57:@3775.4]
  wire [10:0] _T_57012; // @[Modules.scala 65:57:@3776.4]
  wire [10:0] buffer_1_542; // @[Modules.scala 65:57:@3777.4]
  wire [11:0] _T_57020; // @[Modules.scala 65:57:@3787.4]
  wire [10:0] _T_57021; // @[Modules.scala 65:57:@3788.4]
  wire [10:0] buffer_1_545; // @[Modules.scala 65:57:@3789.4]
  wire [11:0] _T_57023; // @[Modules.scala 65:57:@3791.4]
  wire [10:0] _T_57024; // @[Modules.scala 65:57:@3792.4]
  wire [10:0] buffer_1_546; // @[Modules.scala 65:57:@3793.4]
  wire [10:0] buffer_1_310; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57026; // @[Modules.scala 65:57:@3795.4]
  wire [10:0] _T_57027; // @[Modules.scala 65:57:@3796.4]
  wire [10:0] buffer_1_547; // @[Modules.scala 65:57:@3797.4]
  wire [10:0] buffer_1_312; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57029; // @[Modules.scala 65:57:@3799.4]
  wire [10:0] _T_57030; // @[Modules.scala 65:57:@3800.4]
  wire [10:0] buffer_1_548; // @[Modules.scala 65:57:@3801.4]
  wire [10:0] buffer_1_314; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57032; // @[Modules.scala 65:57:@3803.4]
  wire [10:0] _T_57033; // @[Modules.scala 65:57:@3804.4]
  wire [10:0] buffer_1_549; // @[Modules.scala 65:57:@3805.4]
  wire [10:0] buffer_1_316; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57035; // @[Modules.scala 65:57:@3807.4]
  wire [10:0] _T_57036; // @[Modules.scala 65:57:@3808.4]
  wire [10:0] buffer_1_550; // @[Modules.scala 65:57:@3809.4]
  wire [10:0] buffer_1_318; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57038; // @[Modules.scala 65:57:@3811.4]
  wire [10:0] _T_57039; // @[Modules.scala 65:57:@3812.4]
  wire [10:0] buffer_1_551; // @[Modules.scala 65:57:@3813.4]
  wire [10:0] buffer_1_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57041; // @[Modules.scala 65:57:@3815.4]
  wire [10:0] _T_57042; // @[Modules.scala 65:57:@3816.4]
  wire [10:0] buffer_1_552; // @[Modules.scala 65:57:@3817.4]
  wire [11:0] _T_57044; // @[Modules.scala 65:57:@3819.4]
  wire [10:0] _T_57045; // @[Modules.scala 65:57:@3820.4]
  wire [10:0] buffer_1_553; // @[Modules.scala 65:57:@3821.4]
  wire [10:0] buffer_1_324; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57047; // @[Modules.scala 65:57:@3823.4]
  wire [10:0] _T_57048; // @[Modules.scala 65:57:@3824.4]
  wire [10:0] buffer_1_554; // @[Modules.scala 65:57:@3825.4]
  wire [10:0] buffer_1_326; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57050; // @[Modules.scala 65:57:@3827.4]
  wire [10:0] _T_57051; // @[Modules.scala 65:57:@3828.4]
  wire [10:0] buffer_1_555; // @[Modules.scala 65:57:@3829.4]
  wire [10:0] buffer_1_328; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57053; // @[Modules.scala 65:57:@3831.4]
  wire [10:0] _T_57054; // @[Modules.scala 65:57:@3832.4]
  wire [10:0] buffer_1_556; // @[Modules.scala 65:57:@3833.4]
  wire [10:0] buffer_1_331; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57056; // @[Modules.scala 65:57:@3835.4]
  wire [10:0] _T_57057; // @[Modules.scala 65:57:@3836.4]
  wire [10:0] buffer_1_557; // @[Modules.scala 65:57:@3837.4]
  wire [10:0] buffer_1_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57065; // @[Modules.scala 65:57:@3847.4]
  wire [10:0] _T_57066; // @[Modules.scala 65:57:@3848.4]
  wire [10:0] buffer_1_560; // @[Modules.scala 65:57:@3849.4]
  wire [10:0] buffer_1_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57071; // @[Modules.scala 65:57:@3855.4]
  wire [10:0] _T_57072; // @[Modules.scala 65:57:@3856.4]
  wire [10:0] buffer_1_562; // @[Modules.scala 65:57:@3857.4]
  wire [10:0] buffer_1_342; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57074; // @[Modules.scala 65:57:@3859.4]
  wire [10:0] _T_57075; // @[Modules.scala 65:57:@3860.4]
  wire [10:0] buffer_1_563; // @[Modules.scala 65:57:@3861.4]
  wire [10:0] buffer_1_344; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57077; // @[Modules.scala 65:57:@3863.4]
  wire [10:0] _T_57078; // @[Modules.scala 65:57:@3864.4]
  wire [10:0] buffer_1_564; // @[Modules.scala 65:57:@3865.4]
  wire [10:0] buffer_1_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57080; // @[Modules.scala 65:57:@3867.4]
  wire [10:0] _T_57081; // @[Modules.scala 65:57:@3868.4]
  wire [10:0] buffer_1_565; // @[Modules.scala 65:57:@3869.4]
  wire [10:0] buffer_1_348; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57083; // @[Modules.scala 65:57:@3871.4]
  wire [10:0] _T_57084; // @[Modules.scala 65:57:@3872.4]
  wire [10:0] buffer_1_566; // @[Modules.scala 65:57:@3873.4]
  wire [10:0] buffer_1_350; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57086; // @[Modules.scala 65:57:@3875.4]
  wire [10:0] _T_57087; // @[Modules.scala 65:57:@3876.4]
  wire [10:0] buffer_1_567; // @[Modules.scala 65:57:@3877.4]
  wire [10:0] buffer_1_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57092; // @[Modules.scala 65:57:@3883.4]
  wire [10:0] _T_57093; // @[Modules.scala 65:57:@3884.4]
  wire [10:0] buffer_1_569; // @[Modules.scala 65:57:@3885.4]
  wire [10:0] buffer_1_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57095; // @[Modules.scala 65:57:@3887.4]
  wire [10:0] _T_57096; // @[Modules.scala 65:57:@3888.4]
  wire [10:0] buffer_1_570; // @[Modules.scala 65:57:@3889.4]
  wire [10:0] buffer_1_358; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57098; // @[Modules.scala 65:57:@3891.4]
  wire [10:0] _T_57099; // @[Modules.scala 65:57:@3892.4]
  wire [10:0] buffer_1_571; // @[Modules.scala 65:57:@3893.4]
  wire [11:0] _T_57101; // @[Modules.scala 65:57:@3895.4]
  wire [10:0] _T_57102; // @[Modules.scala 65:57:@3896.4]
  wire [10:0] buffer_1_572; // @[Modules.scala 65:57:@3897.4]
  wire [10:0] buffer_1_362; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57104; // @[Modules.scala 65:57:@3899.4]
  wire [10:0] _T_57105; // @[Modules.scala 65:57:@3900.4]
  wire [10:0] buffer_1_573; // @[Modules.scala 65:57:@3901.4]
  wire [10:0] buffer_1_378; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57128; // @[Modules.scala 65:57:@3931.4]
  wire [10:0] _T_57129; // @[Modules.scala 65:57:@3932.4]
  wire [10:0] buffer_1_581; // @[Modules.scala 65:57:@3933.4]
  wire [10:0] buffer_1_380; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_1_381; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57131; // @[Modules.scala 65:57:@3935.4]
  wire [10:0] _T_57132; // @[Modules.scala 65:57:@3936.4]
  wire [10:0] buffer_1_582; // @[Modules.scala 65:57:@3937.4]
  wire [10:0] buffer_1_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57134; // @[Modules.scala 65:57:@3939.4]
  wire [10:0] _T_57135; // @[Modules.scala 65:57:@3940.4]
  wire [10:0] buffer_1_583; // @[Modules.scala 65:57:@3941.4]
  wire [10:0] buffer_1_390; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_57146; // @[Modules.scala 65:57:@3955.4]
  wire [10:0] _T_57147; // @[Modules.scala 65:57:@3956.4]
  wire [10:0] buffer_1_587; // @[Modules.scala 65:57:@3957.4]
  wire [11:0] _T_57149; // @[Modules.scala 68:83:@3959.4]
  wire [10:0] _T_57150; // @[Modules.scala 68:83:@3960.4]
  wire [10:0] buffer_1_588; // @[Modules.scala 68:83:@3961.4]
  wire [11:0] _T_57152; // @[Modules.scala 68:83:@3963.4]
  wire [10:0] _T_57153; // @[Modules.scala 68:83:@3964.4]
  wire [10:0] buffer_1_589; // @[Modules.scala 68:83:@3965.4]
  wire [11:0] _T_57155; // @[Modules.scala 68:83:@3967.4]
  wire [10:0] _T_57156; // @[Modules.scala 68:83:@3968.4]
  wire [10:0] buffer_1_590; // @[Modules.scala 68:83:@3969.4]
  wire [11:0] _T_57158; // @[Modules.scala 68:83:@3971.4]
  wire [10:0] _T_57159; // @[Modules.scala 68:83:@3972.4]
  wire [10:0] buffer_1_591; // @[Modules.scala 68:83:@3973.4]
  wire [11:0] _T_57161; // @[Modules.scala 68:83:@3975.4]
  wire [10:0] _T_57162; // @[Modules.scala 68:83:@3976.4]
  wire [10:0] buffer_1_592; // @[Modules.scala 68:83:@3977.4]
  wire [11:0] _T_57164; // @[Modules.scala 68:83:@3979.4]
  wire [10:0] _T_57165; // @[Modules.scala 68:83:@3980.4]
  wire [10:0] buffer_1_593; // @[Modules.scala 68:83:@3981.4]
  wire [11:0] _T_57167; // @[Modules.scala 68:83:@3983.4]
  wire [10:0] _T_57168; // @[Modules.scala 68:83:@3984.4]
  wire [10:0] buffer_1_594; // @[Modules.scala 68:83:@3985.4]
  wire [11:0] _T_57170; // @[Modules.scala 68:83:@3987.4]
  wire [10:0] _T_57171; // @[Modules.scala 68:83:@3988.4]
  wire [10:0] buffer_1_595; // @[Modules.scala 68:83:@3989.4]
  wire [11:0] _T_57173; // @[Modules.scala 68:83:@3991.4]
  wire [10:0] _T_57174; // @[Modules.scala 68:83:@3992.4]
  wire [10:0] buffer_1_596; // @[Modules.scala 68:83:@3993.4]
  wire [11:0] _T_57176; // @[Modules.scala 68:83:@3995.4]
  wire [10:0] _T_57177; // @[Modules.scala 68:83:@3996.4]
  wire [10:0] buffer_1_597; // @[Modules.scala 68:83:@3997.4]
  wire [11:0] _T_57179; // @[Modules.scala 68:83:@3999.4]
  wire [10:0] _T_57180; // @[Modules.scala 68:83:@4000.4]
  wire [10:0] buffer_1_598; // @[Modules.scala 68:83:@4001.4]
  wire [11:0] _T_57182; // @[Modules.scala 68:83:@4003.4]
  wire [10:0] _T_57183; // @[Modules.scala 68:83:@4004.4]
  wire [10:0] buffer_1_599; // @[Modules.scala 68:83:@4005.4]
  wire [11:0] _T_57185; // @[Modules.scala 68:83:@4007.4]
  wire [10:0] _T_57186; // @[Modules.scala 68:83:@4008.4]
  wire [10:0] buffer_1_600; // @[Modules.scala 68:83:@4009.4]
  wire [11:0] _T_57188; // @[Modules.scala 68:83:@4011.4]
  wire [10:0] _T_57189; // @[Modules.scala 68:83:@4012.4]
  wire [10:0] buffer_1_601; // @[Modules.scala 68:83:@4013.4]
  wire [11:0] _T_57191; // @[Modules.scala 68:83:@4015.4]
  wire [10:0] _T_57192; // @[Modules.scala 68:83:@4016.4]
  wire [10:0] buffer_1_602; // @[Modules.scala 68:83:@4017.4]
  wire [11:0] _T_57194; // @[Modules.scala 68:83:@4019.4]
  wire [10:0] _T_57195; // @[Modules.scala 68:83:@4020.4]
  wire [10:0] buffer_1_603; // @[Modules.scala 68:83:@4021.4]
  wire [11:0] _T_57197; // @[Modules.scala 68:83:@4023.4]
  wire [10:0] _T_57198; // @[Modules.scala 68:83:@4024.4]
  wire [10:0] buffer_1_604; // @[Modules.scala 68:83:@4025.4]
  wire [11:0] _T_57200; // @[Modules.scala 68:83:@4027.4]
  wire [10:0] _T_57201; // @[Modules.scala 68:83:@4028.4]
  wire [10:0] buffer_1_605; // @[Modules.scala 68:83:@4029.4]
  wire [11:0] _T_57203; // @[Modules.scala 68:83:@4031.4]
  wire [10:0] _T_57204; // @[Modules.scala 68:83:@4032.4]
  wire [10:0] buffer_1_606; // @[Modules.scala 68:83:@4033.4]
  wire [11:0] _T_57206; // @[Modules.scala 68:83:@4035.4]
  wire [10:0] _T_57207; // @[Modules.scala 68:83:@4036.4]
  wire [10:0] buffer_1_607; // @[Modules.scala 68:83:@4037.4]
  wire [11:0] _T_57209; // @[Modules.scala 68:83:@4039.4]
  wire [10:0] _T_57210; // @[Modules.scala 68:83:@4040.4]
  wire [10:0] buffer_1_608; // @[Modules.scala 68:83:@4041.4]
  wire [11:0] _T_57212; // @[Modules.scala 68:83:@4043.4]
  wire [10:0] _T_57213; // @[Modules.scala 68:83:@4044.4]
  wire [10:0] buffer_1_609; // @[Modules.scala 68:83:@4045.4]
  wire [11:0] _T_57215; // @[Modules.scala 68:83:@4047.4]
  wire [10:0] _T_57216; // @[Modules.scala 68:83:@4048.4]
  wire [10:0] buffer_1_610; // @[Modules.scala 68:83:@4049.4]
  wire [11:0] _T_57218; // @[Modules.scala 68:83:@4051.4]
  wire [10:0] _T_57219; // @[Modules.scala 68:83:@4052.4]
  wire [10:0] buffer_1_611; // @[Modules.scala 68:83:@4053.4]
  wire [11:0] _T_57221; // @[Modules.scala 68:83:@4055.4]
  wire [10:0] _T_57222; // @[Modules.scala 68:83:@4056.4]
  wire [10:0] buffer_1_612; // @[Modules.scala 68:83:@4057.4]
  wire [11:0] _T_57224; // @[Modules.scala 68:83:@4059.4]
  wire [10:0] _T_57225; // @[Modules.scala 68:83:@4060.4]
  wire [10:0] buffer_1_613; // @[Modules.scala 68:83:@4061.4]
  wire [11:0] _T_57227; // @[Modules.scala 68:83:@4063.4]
  wire [10:0] _T_57228; // @[Modules.scala 68:83:@4064.4]
  wire [10:0] buffer_1_614; // @[Modules.scala 68:83:@4065.4]
  wire [11:0] _T_57230; // @[Modules.scala 68:83:@4067.4]
  wire [10:0] _T_57231; // @[Modules.scala 68:83:@4068.4]
  wire [10:0] buffer_1_615; // @[Modules.scala 68:83:@4069.4]
  wire [11:0] _T_57233; // @[Modules.scala 68:83:@4071.4]
  wire [10:0] _T_57234; // @[Modules.scala 68:83:@4072.4]
  wire [10:0] buffer_1_616; // @[Modules.scala 68:83:@4073.4]
  wire [11:0] _T_57239; // @[Modules.scala 68:83:@4079.4]
  wire [10:0] _T_57240; // @[Modules.scala 68:83:@4080.4]
  wire [10:0] buffer_1_618; // @[Modules.scala 68:83:@4081.4]
  wire [11:0] _T_57242; // @[Modules.scala 68:83:@4083.4]
  wire [10:0] _T_57243; // @[Modules.scala 68:83:@4084.4]
  wire [10:0] buffer_1_619; // @[Modules.scala 68:83:@4085.4]
  wire [11:0] _T_57245; // @[Modules.scala 68:83:@4087.4]
  wire [10:0] _T_57246; // @[Modules.scala 68:83:@4088.4]
  wire [10:0] buffer_1_620; // @[Modules.scala 68:83:@4089.4]
  wire [11:0] _T_57248; // @[Modules.scala 68:83:@4091.4]
  wire [10:0] _T_57249; // @[Modules.scala 68:83:@4092.4]
  wire [10:0] buffer_1_621; // @[Modules.scala 68:83:@4093.4]
  wire [11:0] _T_57251; // @[Modules.scala 68:83:@4095.4]
  wire [10:0] _T_57252; // @[Modules.scala 68:83:@4096.4]
  wire [10:0] buffer_1_622; // @[Modules.scala 68:83:@4097.4]
  wire [11:0] _T_57254; // @[Modules.scala 68:83:@4099.4]
  wire [10:0] _T_57255; // @[Modules.scala 68:83:@4100.4]
  wire [10:0] buffer_1_623; // @[Modules.scala 68:83:@4101.4]
  wire [11:0] _T_57257; // @[Modules.scala 68:83:@4103.4]
  wire [10:0] _T_57258; // @[Modules.scala 68:83:@4104.4]
  wire [10:0] buffer_1_624; // @[Modules.scala 68:83:@4105.4]
  wire [11:0] _T_57260; // @[Modules.scala 68:83:@4107.4]
  wire [10:0] _T_57261; // @[Modules.scala 68:83:@4108.4]
  wire [10:0] buffer_1_625; // @[Modules.scala 68:83:@4109.4]
  wire [11:0] _T_57263; // @[Modules.scala 68:83:@4111.4]
  wire [10:0] _T_57264; // @[Modules.scala 68:83:@4112.4]
  wire [10:0] buffer_1_626; // @[Modules.scala 68:83:@4113.4]
  wire [11:0] _T_57266; // @[Modules.scala 68:83:@4115.4]
  wire [10:0] _T_57267; // @[Modules.scala 68:83:@4116.4]
  wire [10:0] buffer_1_627; // @[Modules.scala 68:83:@4117.4]
  wire [11:0] _T_57269; // @[Modules.scala 68:83:@4119.4]
  wire [10:0] _T_57270; // @[Modules.scala 68:83:@4120.4]
  wire [10:0] buffer_1_628; // @[Modules.scala 68:83:@4121.4]
  wire [11:0] _T_57272; // @[Modules.scala 68:83:@4123.4]
  wire [10:0] _T_57273; // @[Modules.scala 68:83:@4124.4]
  wire [10:0] buffer_1_629; // @[Modules.scala 68:83:@4125.4]
  wire [11:0] _T_57278; // @[Modules.scala 68:83:@4131.4]
  wire [10:0] _T_57279; // @[Modules.scala 68:83:@4132.4]
  wire [10:0] buffer_1_631; // @[Modules.scala 68:83:@4133.4]
  wire [11:0] _T_57281; // @[Modules.scala 68:83:@4135.4]
  wire [10:0] _T_57282; // @[Modules.scala 68:83:@4136.4]
  wire [10:0] buffer_1_632; // @[Modules.scala 68:83:@4137.4]
  wire [11:0] _T_57284; // @[Modules.scala 68:83:@4139.4]
  wire [10:0] _T_57285; // @[Modules.scala 68:83:@4140.4]
  wire [10:0] buffer_1_633; // @[Modules.scala 68:83:@4141.4]
  wire [11:0] _T_57287; // @[Modules.scala 68:83:@4143.4]
  wire [10:0] _T_57288; // @[Modules.scala 68:83:@4144.4]
  wire [10:0] buffer_1_634; // @[Modules.scala 68:83:@4145.4]
  wire [11:0] _T_57290; // @[Modules.scala 68:83:@4147.4]
  wire [10:0] _T_57291; // @[Modules.scala 68:83:@4148.4]
  wire [10:0] buffer_1_635; // @[Modules.scala 68:83:@4149.4]
  wire [11:0] _T_57293; // @[Modules.scala 68:83:@4151.4]
  wire [10:0] _T_57294; // @[Modules.scala 68:83:@4152.4]
  wire [10:0] buffer_1_636; // @[Modules.scala 68:83:@4153.4]
  wire [11:0] _T_57296; // @[Modules.scala 68:83:@4155.4]
  wire [10:0] _T_57297; // @[Modules.scala 68:83:@4156.4]
  wire [10:0] buffer_1_637; // @[Modules.scala 68:83:@4157.4]
  wire [11:0] _T_57299; // @[Modules.scala 68:83:@4159.4]
  wire [10:0] _T_57300; // @[Modules.scala 68:83:@4160.4]
  wire [10:0] buffer_1_638; // @[Modules.scala 68:83:@4161.4]
  wire [11:0] _T_57302; // @[Modules.scala 68:83:@4163.4]
  wire [10:0] _T_57303; // @[Modules.scala 68:83:@4164.4]
  wire [10:0] buffer_1_639; // @[Modules.scala 68:83:@4165.4]
  wire [11:0] _T_57305; // @[Modules.scala 68:83:@4167.4]
  wire [10:0] _T_57306; // @[Modules.scala 68:83:@4168.4]
  wire [10:0] buffer_1_640; // @[Modules.scala 68:83:@4169.4]
  wire [11:0] _T_57308; // @[Modules.scala 68:83:@4171.4]
  wire [10:0] _T_57309; // @[Modules.scala 68:83:@4172.4]
  wire [10:0] buffer_1_641; // @[Modules.scala 68:83:@4173.4]
  wire [11:0] _T_57311; // @[Modules.scala 68:83:@4175.4]
  wire [10:0] _T_57312; // @[Modules.scala 68:83:@4176.4]
  wire [10:0] buffer_1_642; // @[Modules.scala 68:83:@4177.4]
  wire [11:0] _T_57314; // @[Modules.scala 68:83:@4179.4]
  wire [10:0] _T_57315; // @[Modules.scala 68:83:@4180.4]
  wire [10:0] buffer_1_643; // @[Modules.scala 68:83:@4181.4]
  wire [11:0] _T_57317; // @[Modules.scala 68:83:@4183.4]
  wire [10:0] _T_57318; // @[Modules.scala 68:83:@4184.4]
  wire [10:0] buffer_1_644; // @[Modules.scala 68:83:@4185.4]
  wire [11:0] _T_57320; // @[Modules.scala 68:83:@4187.4]
  wire [10:0] _T_57321; // @[Modules.scala 68:83:@4188.4]
  wire [10:0] buffer_1_645; // @[Modules.scala 68:83:@4189.4]
  wire [11:0] _T_57323; // @[Modules.scala 68:83:@4191.4]
  wire [10:0] _T_57324; // @[Modules.scala 68:83:@4192.4]
  wire [10:0] buffer_1_646; // @[Modules.scala 68:83:@4193.4]
  wire [11:0] _T_57326; // @[Modules.scala 68:83:@4195.4]
  wire [10:0] _T_57327; // @[Modules.scala 68:83:@4196.4]
  wire [10:0] buffer_1_647; // @[Modules.scala 68:83:@4197.4]
  wire [11:0] _T_57329; // @[Modules.scala 68:83:@4199.4]
  wire [10:0] _T_57330; // @[Modules.scala 68:83:@4200.4]
  wire [10:0] buffer_1_648; // @[Modules.scala 68:83:@4201.4]
  wire [11:0] _T_57332; // @[Modules.scala 68:83:@4203.4]
  wire [10:0] _T_57333; // @[Modules.scala 68:83:@4204.4]
  wire [10:0] buffer_1_649; // @[Modules.scala 68:83:@4205.4]
  wire [11:0] _T_57335; // @[Modules.scala 68:83:@4207.4]
  wire [10:0] _T_57336; // @[Modules.scala 68:83:@4208.4]
  wire [10:0] buffer_1_650; // @[Modules.scala 68:83:@4209.4]
  wire [11:0] _T_57338; // @[Modules.scala 68:83:@4211.4]
  wire [10:0] _T_57339; // @[Modules.scala 68:83:@4212.4]
  wire [10:0] buffer_1_651; // @[Modules.scala 68:83:@4213.4]
  wire [11:0] _T_57341; // @[Modules.scala 68:83:@4215.4]
  wire [10:0] _T_57342; // @[Modules.scala 68:83:@4216.4]
  wire [10:0] buffer_1_652; // @[Modules.scala 68:83:@4217.4]
  wire [11:0] _T_57344; // @[Modules.scala 68:83:@4219.4]
  wire [10:0] _T_57345; // @[Modules.scala 68:83:@4220.4]
  wire [10:0] buffer_1_653; // @[Modules.scala 68:83:@4221.4]
  wire [11:0] _T_57347; // @[Modules.scala 68:83:@4223.4]
  wire [10:0] _T_57348; // @[Modules.scala 68:83:@4224.4]
  wire [10:0] buffer_1_654; // @[Modules.scala 68:83:@4225.4]
  wire [11:0] _T_57350; // @[Modules.scala 68:83:@4227.4]
  wire [10:0] _T_57351; // @[Modules.scala 68:83:@4228.4]
  wire [10:0] buffer_1_655; // @[Modules.scala 68:83:@4229.4]
  wire [11:0] _T_57353; // @[Modules.scala 68:83:@4231.4]
  wire [10:0] _T_57354; // @[Modules.scala 68:83:@4232.4]
  wire [10:0] buffer_1_656; // @[Modules.scala 68:83:@4233.4]
  wire [11:0] _T_57356; // @[Modules.scala 68:83:@4235.4]
  wire [10:0] _T_57357; // @[Modules.scala 68:83:@4236.4]
  wire [10:0] buffer_1_657; // @[Modules.scala 68:83:@4237.4]
  wire [11:0] _T_57359; // @[Modules.scala 68:83:@4239.4]
  wire [10:0] _T_57360; // @[Modules.scala 68:83:@4240.4]
  wire [10:0] buffer_1_658; // @[Modules.scala 68:83:@4241.4]
  wire [11:0] _T_57362; // @[Modules.scala 68:83:@4243.4]
  wire [10:0] _T_57363; // @[Modules.scala 68:83:@4244.4]
  wire [10:0] buffer_1_659; // @[Modules.scala 68:83:@4245.4]
  wire [11:0] _T_57365; // @[Modules.scala 68:83:@4247.4]
  wire [10:0] _T_57366; // @[Modules.scala 68:83:@4248.4]
  wire [10:0] buffer_1_660; // @[Modules.scala 68:83:@4249.4]
  wire [11:0] _T_57368; // @[Modules.scala 68:83:@4251.4]
  wire [10:0] _T_57369; // @[Modules.scala 68:83:@4252.4]
  wire [10:0] buffer_1_661; // @[Modules.scala 68:83:@4253.4]
  wire [11:0] _T_57371; // @[Modules.scala 68:83:@4255.4]
  wire [10:0] _T_57372; // @[Modules.scala 68:83:@4256.4]
  wire [10:0] buffer_1_662; // @[Modules.scala 68:83:@4257.4]
  wire [11:0] _T_57374; // @[Modules.scala 68:83:@4259.4]
  wire [10:0] _T_57375; // @[Modules.scala 68:83:@4260.4]
  wire [10:0] buffer_1_663; // @[Modules.scala 68:83:@4261.4]
  wire [11:0] _T_57377; // @[Modules.scala 68:83:@4263.4]
  wire [10:0] _T_57378; // @[Modules.scala 68:83:@4264.4]
  wire [10:0] buffer_1_664; // @[Modules.scala 68:83:@4265.4]
  wire [11:0] _T_57380; // @[Modules.scala 68:83:@4267.4]
  wire [10:0] _T_57381; // @[Modules.scala 68:83:@4268.4]
  wire [10:0] buffer_1_665; // @[Modules.scala 68:83:@4269.4]
  wire [11:0] _T_57383; // @[Modules.scala 68:83:@4271.4]
  wire [10:0] _T_57384; // @[Modules.scala 68:83:@4272.4]
  wire [10:0] buffer_1_666; // @[Modules.scala 68:83:@4273.4]
  wire [11:0] _T_57386; // @[Modules.scala 68:83:@4275.4]
  wire [10:0] _T_57387; // @[Modules.scala 68:83:@4276.4]
  wire [10:0] buffer_1_667; // @[Modules.scala 68:83:@4277.4]
  wire [11:0] _T_57389; // @[Modules.scala 68:83:@4279.4]
  wire [10:0] _T_57390; // @[Modules.scala 68:83:@4280.4]
  wire [10:0] buffer_1_668; // @[Modules.scala 68:83:@4281.4]
  wire [11:0] _T_57392; // @[Modules.scala 68:83:@4283.4]
  wire [10:0] _T_57393; // @[Modules.scala 68:83:@4284.4]
  wire [10:0] buffer_1_669; // @[Modules.scala 68:83:@4285.4]
  wire [11:0] _T_57395; // @[Modules.scala 68:83:@4287.4]
  wire [10:0] _T_57396; // @[Modules.scala 68:83:@4288.4]
  wire [10:0] buffer_1_670; // @[Modules.scala 68:83:@4289.4]
  wire [11:0] _T_57401; // @[Modules.scala 68:83:@4295.4]
  wire [10:0] _T_57402; // @[Modules.scala 68:83:@4296.4]
  wire [10:0] buffer_1_672; // @[Modules.scala 68:83:@4297.4]
  wire [11:0] _T_57404; // @[Modules.scala 68:83:@4299.4]
  wire [10:0] _T_57405; // @[Modules.scala 68:83:@4300.4]
  wire [10:0] buffer_1_673; // @[Modules.scala 68:83:@4301.4]
  wire [11:0] _T_57407; // @[Modules.scala 68:83:@4303.4]
  wire [10:0] _T_57408; // @[Modules.scala 68:83:@4304.4]
  wire [10:0] buffer_1_674; // @[Modules.scala 68:83:@4305.4]
  wire [11:0] _T_57410; // @[Modules.scala 68:83:@4307.4]
  wire [10:0] _T_57411; // @[Modules.scala 68:83:@4308.4]
  wire [10:0] buffer_1_675; // @[Modules.scala 68:83:@4309.4]
  wire [11:0] _T_57413; // @[Modules.scala 68:83:@4311.4]
  wire [10:0] _T_57414; // @[Modules.scala 68:83:@4312.4]
  wire [10:0] buffer_1_676; // @[Modules.scala 68:83:@4313.4]
  wire [11:0] _T_57416; // @[Modules.scala 68:83:@4315.4]
  wire [10:0] _T_57417; // @[Modules.scala 68:83:@4316.4]
  wire [10:0] buffer_1_677; // @[Modules.scala 68:83:@4317.4]
  wire [11:0] _T_57419; // @[Modules.scala 68:83:@4319.4]
  wire [10:0] _T_57420; // @[Modules.scala 68:83:@4320.4]
  wire [10:0] buffer_1_678; // @[Modules.scala 68:83:@4321.4]
  wire [11:0] _T_57431; // @[Modules.scala 68:83:@4335.4]
  wire [10:0] _T_57432; // @[Modules.scala 68:83:@4336.4]
  wire [10:0] buffer_1_682; // @[Modules.scala 68:83:@4337.4]
  wire [11:0] _T_57434; // @[Modules.scala 68:83:@4339.4]
  wire [10:0] _T_57435; // @[Modules.scala 68:83:@4340.4]
  wire [10:0] buffer_1_683; // @[Modules.scala 68:83:@4341.4]
  wire [11:0] _T_57440; // @[Modules.scala 68:83:@4347.4]
  wire [10:0] _T_57441; // @[Modules.scala 68:83:@4348.4]
  wire [10:0] buffer_1_685; // @[Modules.scala 68:83:@4349.4]
  wire [11:0] _T_57443; // @[Modules.scala 71:109:@4351.4]
  wire [10:0] _T_57444; // @[Modules.scala 71:109:@4352.4]
  wire [10:0] buffer_1_686; // @[Modules.scala 71:109:@4353.4]
  wire [11:0] _T_57446; // @[Modules.scala 71:109:@4355.4]
  wire [10:0] _T_57447; // @[Modules.scala 71:109:@4356.4]
  wire [10:0] buffer_1_687; // @[Modules.scala 71:109:@4357.4]
  wire [11:0] _T_57449; // @[Modules.scala 71:109:@4359.4]
  wire [10:0] _T_57450; // @[Modules.scala 71:109:@4360.4]
  wire [10:0] buffer_1_688; // @[Modules.scala 71:109:@4361.4]
  wire [11:0] _T_57452; // @[Modules.scala 71:109:@4363.4]
  wire [10:0] _T_57453; // @[Modules.scala 71:109:@4364.4]
  wire [10:0] buffer_1_689; // @[Modules.scala 71:109:@4365.4]
  wire [11:0] _T_57455; // @[Modules.scala 71:109:@4367.4]
  wire [10:0] _T_57456; // @[Modules.scala 71:109:@4368.4]
  wire [10:0] buffer_1_690; // @[Modules.scala 71:109:@4369.4]
  wire [11:0] _T_57458; // @[Modules.scala 71:109:@4371.4]
  wire [10:0] _T_57459; // @[Modules.scala 71:109:@4372.4]
  wire [10:0] buffer_1_691; // @[Modules.scala 71:109:@4373.4]
  wire [11:0] _T_57461; // @[Modules.scala 71:109:@4375.4]
  wire [10:0] _T_57462; // @[Modules.scala 71:109:@4376.4]
  wire [10:0] buffer_1_692; // @[Modules.scala 71:109:@4377.4]
  wire [11:0] _T_57464; // @[Modules.scala 71:109:@4379.4]
  wire [10:0] _T_57465; // @[Modules.scala 71:109:@4380.4]
  wire [10:0] buffer_1_693; // @[Modules.scala 71:109:@4381.4]
  wire [11:0] _T_57467; // @[Modules.scala 71:109:@4383.4]
  wire [10:0] _T_57468; // @[Modules.scala 71:109:@4384.4]
  wire [10:0] buffer_1_694; // @[Modules.scala 71:109:@4385.4]
  wire [11:0] _T_57470; // @[Modules.scala 71:109:@4387.4]
  wire [10:0] _T_57471; // @[Modules.scala 71:109:@4388.4]
  wire [10:0] buffer_1_695; // @[Modules.scala 71:109:@4389.4]
  wire [11:0] _T_57473; // @[Modules.scala 71:109:@4391.4]
  wire [10:0] _T_57474; // @[Modules.scala 71:109:@4392.4]
  wire [10:0] buffer_1_696; // @[Modules.scala 71:109:@4393.4]
  wire [11:0] _T_57476; // @[Modules.scala 71:109:@4395.4]
  wire [10:0] _T_57477; // @[Modules.scala 71:109:@4396.4]
  wire [10:0] buffer_1_697; // @[Modules.scala 71:109:@4397.4]
  wire [11:0] _T_57479; // @[Modules.scala 71:109:@4399.4]
  wire [10:0] _T_57480; // @[Modules.scala 71:109:@4400.4]
  wire [10:0] buffer_1_698; // @[Modules.scala 71:109:@4401.4]
  wire [11:0] _T_57482; // @[Modules.scala 71:109:@4403.4]
  wire [10:0] _T_57483; // @[Modules.scala 71:109:@4404.4]
  wire [10:0] buffer_1_699; // @[Modules.scala 71:109:@4405.4]
  wire [11:0] _T_57485; // @[Modules.scala 71:109:@4407.4]
  wire [10:0] _T_57486; // @[Modules.scala 71:109:@4408.4]
  wire [10:0] buffer_1_700; // @[Modules.scala 71:109:@4409.4]
  wire [11:0] _T_57488; // @[Modules.scala 71:109:@4411.4]
  wire [10:0] _T_57489; // @[Modules.scala 71:109:@4412.4]
  wire [10:0] buffer_1_701; // @[Modules.scala 71:109:@4413.4]
  wire [11:0] _T_57491; // @[Modules.scala 71:109:@4415.4]
  wire [10:0] _T_57492; // @[Modules.scala 71:109:@4416.4]
  wire [10:0] buffer_1_702; // @[Modules.scala 71:109:@4417.4]
  wire [11:0] _T_57494; // @[Modules.scala 71:109:@4419.4]
  wire [10:0] _T_57495; // @[Modules.scala 71:109:@4420.4]
  wire [10:0] buffer_1_703; // @[Modules.scala 71:109:@4421.4]
  wire [11:0] _T_57497; // @[Modules.scala 71:109:@4423.4]
  wire [10:0] _T_57498; // @[Modules.scala 71:109:@4424.4]
  wire [10:0] buffer_1_704; // @[Modules.scala 71:109:@4425.4]
  wire [11:0] _T_57500; // @[Modules.scala 71:109:@4427.4]
  wire [10:0] _T_57501; // @[Modules.scala 71:109:@4428.4]
  wire [10:0] buffer_1_705; // @[Modules.scala 71:109:@4429.4]
  wire [11:0] _T_57503; // @[Modules.scala 71:109:@4431.4]
  wire [10:0] _T_57504; // @[Modules.scala 71:109:@4432.4]
  wire [10:0] buffer_1_706; // @[Modules.scala 71:109:@4433.4]
  wire [11:0] _T_57506; // @[Modules.scala 71:109:@4435.4]
  wire [10:0] _T_57507; // @[Modules.scala 71:109:@4436.4]
  wire [10:0] buffer_1_707; // @[Modules.scala 71:109:@4437.4]
  wire [11:0] _T_57509; // @[Modules.scala 71:109:@4439.4]
  wire [10:0] _T_57510; // @[Modules.scala 71:109:@4440.4]
  wire [10:0] buffer_1_708; // @[Modules.scala 71:109:@4441.4]
  wire [11:0] _T_57512; // @[Modules.scala 71:109:@4443.4]
  wire [10:0] _T_57513; // @[Modules.scala 71:109:@4444.4]
  wire [10:0] buffer_1_709; // @[Modules.scala 71:109:@4445.4]
  wire [11:0] _T_57515; // @[Modules.scala 71:109:@4447.4]
  wire [10:0] _T_57516; // @[Modules.scala 71:109:@4448.4]
  wire [10:0] buffer_1_710; // @[Modules.scala 71:109:@4449.4]
  wire [11:0] _T_57518; // @[Modules.scala 71:109:@4451.4]
  wire [10:0] _T_57519; // @[Modules.scala 71:109:@4452.4]
  wire [10:0] buffer_1_711; // @[Modules.scala 71:109:@4453.4]
  wire [11:0] _T_57521; // @[Modules.scala 71:109:@4455.4]
  wire [10:0] _T_57522; // @[Modules.scala 71:109:@4456.4]
  wire [10:0] buffer_1_712; // @[Modules.scala 71:109:@4457.4]
  wire [11:0] _T_57524; // @[Modules.scala 71:109:@4459.4]
  wire [10:0] _T_57525; // @[Modules.scala 71:109:@4460.4]
  wire [10:0] buffer_1_713; // @[Modules.scala 71:109:@4461.4]
  wire [11:0] _T_57527; // @[Modules.scala 71:109:@4463.4]
  wire [10:0] _T_57528; // @[Modules.scala 71:109:@4464.4]
  wire [10:0] buffer_1_714; // @[Modules.scala 71:109:@4465.4]
  wire [11:0] _T_57530; // @[Modules.scala 71:109:@4467.4]
  wire [10:0] _T_57531; // @[Modules.scala 71:109:@4468.4]
  wire [10:0] buffer_1_715; // @[Modules.scala 71:109:@4469.4]
  wire [11:0] _T_57533; // @[Modules.scala 71:109:@4471.4]
  wire [10:0] _T_57534; // @[Modules.scala 71:109:@4472.4]
  wire [10:0] buffer_1_716; // @[Modules.scala 71:109:@4473.4]
  wire [11:0] _T_57536; // @[Modules.scala 71:109:@4475.4]
  wire [10:0] _T_57537; // @[Modules.scala 71:109:@4476.4]
  wire [10:0] buffer_1_717; // @[Modules.scala 71:109:@4477.4]
  wire [11:0] _T_57539; // @[Modules.scala 71:109:@4479.4]
  wire [10:0] _T_57540; // @[Modules.scala 71:109:@4480.4]
  wire [10:0] buffer_1_718; // @[Modules.scala 71:109:@4481.4]
  wire [11:0] _T_57542; // @[Modules.scala 71:109:@4483.4]
  wire [10:0] _T_57543; // @[Modules.scala 71:109:@4484.4]
  wire [10:0] buffer_1_719; // @[Modules.scala 71:109:@4485.4]
  wire [11:0] _T_57545; // @[Modules.scala 71:109:@4487.4]
  wire [10:0] _T_57546; // @[Modules.scala 71:109:@4488.4]
  wire [10:0] buffer_1_720; // @[Modules.scala 71:109:@4489.4]
  wire [11:0] _T_57548; // @[Modules.scala 71:109:@4491.4]
  wire [10:0] _T_57549; // @[Modules.scala 71:109:@4492.4]
  wire [10:0] buffer_1_721; // @[Modules.scala 71:109:@4493.4]
  wire [11:0] _T_57551; // @[Modules.scala 71:109:@4495.4]
  wire [10:0] _T_57552; // @[Modules.scala 71:109:@4496.4]
  wire [10:0] buffer_1_722; // @[Modules.scala 71:109:@4497.4]
  wire [11:0] _T_57554; // @[Modules.scala 71:109:@4499.4]
  wire [10:0] _T_57555; // @[Modules.scala 71:109:@4500.4]
  wire [10:0] buffer_1_723; // @[Modules.scala 71:109:@4501.4]
  wire [11:0] _T_57557; // @[Modules.scala 71:109:@4503.4]
  wire [10:0] _T_57558; // @[Modules.scala 71:109:@4504.4]
  wire [10:0] buffer_1_724; // @[Modules.scala 71:109:@4505.4]
  wire [11:0] _T_57560; // @[Modules.scala 71:109:@4507.4]
  wire [10:0] _T_57561; // @[Modules.scala 71:109:@4508.4]
  wire [10:0] buffer_1_725; // @[Modules.scala 71:109:@4509.4]
  wire [11:0] _T_57563; // @[Modules.scala 71:109:@4511.4]
  wire [10:0] _T_57564; // @[Modules.scala 71:109:@4512.4]
  wire [10:0] buffer_1_726; // @[Modules.scala 71:109:@4513.4]
  wire [11:0] _T_57566; // @[Modules.scala 71:109:@4515.4]
  wire [10:0] _T_57567; // @[Modules.scala 71:109:@4516.4]
  wire [10:0] buffer_1_727; // @[Modules.scala 71:109:@4517.4]
  wire [11:0] _T_57569; // @[Modules.scala 71:109:@4519.4]
  wire [10:0] _T_57570; // @[Modules.scala 71:109:@4520.4]
  wire [10:0] buffer_1_728; // @[Modules.scala 71:109:@4521.4]
  wire [11:0] _T_57572; // @[Modules.scala 71:109:@4523.4]
  wire [10:0] _T_57573; // @[Modules.scala 71:109:@4524.4]
  wire [10:0] buffer_1_729; // @[Modules.scala 71:109:@4525.4]
  wire [11:0] _T_57575; // @[Modules.scala 71:109:@4527.4]
  wire [10:0] _T_57576; // @[Modules.scala 71:109:@4528.4]
  wire [10:0] buffer_1_730; // @[Modules.scala 71:109:@4529.4]
  wire [11:0] _T_57578; // @[Modules.scala 71:109:@4531.4]
  wire [10:0] _T_57579; // @[Modules.scala 71:109:@4532.4]
  wire [10:0] buffer_1_731; // @[Modules.scala 71:109:@4533.4]
  wire [11:0] _T_57581; // @[Modules.scala 71:109:@4535.4]
  wire [10:0] _T_57582; // @[Modules.scala 71:109:@4536.4]
  wire [10:0] buffer_1_732; // @[Modules.scala 71:109:@4537.4]
  wire [11:0] _T_57584; // @[Modules.scala 71:109:@4539.4]
  wire [10:0] _T_57585; // @[Modules.scala 71:109:@4540.4]
  wire [10:0] buffer_1_733; // @[Modules.scala 71:109:@4541.4]
  wire [11:0] _T_57587; // @[Modules.scala 71:109:@4543.4]
  wire [10:0] _T_57588; // @[Modules.scala 71:109:@4544.4]
  wire [10:0] buffer_1_734; // @[Modules.scala 71:109:@4545.4]
  wire [11:0] _T_57590; // @[Modules.scala 78:156:@4548.4]
  wire [10:0] _T_57591; // @[Modules.scala 78:156:@4549.4]
  wire [10:0] buffer_1_736; // @[Modules.scala 78:156:@4550.4]
  wire [11:0] _T_57593; // @[Modules.scala 78:156:@4552.4]
  wire [10:0] _T_57594; // @[Modules.scala 78:156:@4553.4]
  wire [10:0] buffer_1_737; // @[Modules.scala 78:156:@4554.4]
  wire [11:0] _T_57596; // @[Modules.scala 78:156:@4556.4]
  wire [10:0] _T_57597; // @[Modules.scala 78:156:@4557.4]
  wire [10:0] buffer_1_738; // @[Modules.scala 78:156:@4558.4]
  wire [11:0] _T_57599; // @[Modules.scala 78:156:@4560.4]
  wire [10:0] _T_57600; // @[Modules.scala 78:156:@4561.4]
  wire [10:0] buffer_1_739; // @[Modules.scala 78:156:@4562.4]
  wire [11:0] _T_57602; // @[Modules.scala 78:156:@4564.4]
  wire [10:0] _T_57603; // @[Modules.scala 78:156:@4565.4]
  wire [10:0] buffer_1_740; // @[Modules.scala 78:156:@4566.4]
  wire [11:0] _T_57605; // @[Modules.scala 78:156:@4568.4]
  wire [10:0] _T_57606; // @[Modules.scala 78:156:@4569.4]
  wire [10:0] buffer_1_741; // @[Modules.scala 78:156:@4570.4]
  wire [11:0] _T_57608; // @[Modules.scala 78:156:@4572.4]
  wire [10:0] _T_57609; // @[Modules.scala 78:156:@4573.4]
  wire [10:0] buffer_1_742; // @[Modules.scala 78:156:@4574.4]
  wire [11:0] _T_57611; // @[Modules.scala 78:156:@4576.4]
  wire [10:0] _T_57612; // @[Modules.scala 78:156:@4577.4]
  wire [10:0] buffer_1_743; // @[Modules.scala 78:156:@4578.4]
  wire [11:0] _T_57614; // @[Modules.scala 78:156:@4580.4]
  wire [10:0] _T_57615; // @[Modules.scala 78:156:@4581.4]
  wire [10:0] buffer_1_744; // @[Modules.scala 78:156:@4582.4]
  wire [11:0] _T_57617; // @[Modules.scala 78:156:@4584.4]
  wire [10:0] _T_57618; // @[Modules.scala 78:156:@4585.4]
  wire [10:0] buffer_1_745; // @[Modules.scala 78:156:@4586.4]
  wire [11:0] _T_57620; // @[Modules.scala 78:156:@4588.4]
  wire [10:0] _T_57621; // @[Modules.scala 78:156:@4589.4]
  wire [10:0] buffer_1_746; // @[Modules.scala 78:156:@4590.4]
  wire [11:0] _T_57623; // @[Modules.scala 78:156:@4592.4]
  wire [10:0] _T_57624; // @[Modules.scala 78:156:@4593.4]
  wire [10:0] buffer_1_747; // @[Modules.scala 78:156:@4594.4]
  wire [11:0] _T_57626; // @[Modules.scala 78:156:@4596.4]
  wire [10:0] _T_57627; // @[Modules.scala 78:156:@4597.4]
  wire [10:0] buffer_1_748; // @[Modules.scala 78:156:@4598.4]
  wire [11:0] _T_57629; // @[Modules.scala 78:156:@4600.4]
  wire [10:0] _T_57630; // @[Modules.scala 78:156:@4601.4]
  wire [10:0] buffer_1_749; // @[Modules.scala 78:156:@4602.4]
  wire [11:0] _T_57632; // @[Modules.scala 78:156:@4604.4]
  wire [10:0] _T_57633; // @[Modules.scala 78:156:@4605.4]
  wire [10:0] buffer_1_750; // @[Modules.scala 78:156:@4606.4]
  wire [11:0] _T_57635; // @[Modules.scala 78:156:@4608.4]
  wire [10:0] _T_57636; // @[Modules.scala 78:156:@4609.4]
  wire [10:0] buffer_1_751; // @[Modules.scala 78:156:@4610.4]
  wire [11:0] _T_57638; // @[Modules.scala 78:156:@4612.4]
  wire [10:0] _T_57639; // @[Modules.scala 78:156:@4613.4]
  wire [10:0] buffer_1_752; // @[Modules.scala 78:156:@4614.4]
  wire [11:0] _T_57641; // @[Modules.scala 78:156:@4616.4]
  wire [10:0] _T_57642; // @[Modules.scala 78:156:@4617.4]
  wire [10:0] buffer_1_753; // @[Modules.scala 78:156:@4618.4]
  wire [11:0] _T_57644; // @[Modules.scala 78:156:@4620.4]
  wire [10:0] _T_57645; // @[Modules.scala 78:156:@4621.4]
  wire [10:0] buffer_1_754; // @[Modules.scala 78:156:@4622.4]
  wire [11:0] _T_57647; // @[Modules.scala 78:156:@4624.4]
  wire [10:0] _T_57648; // @[Modules.scala 78:156:@4625.4]
  wire [10:0] buffer_1_755; // @[Modules.scala 78:156:@4626.4]
  wire [11:0] _T_57650; // @[Modules.scala 78:156:@4628.4]
  wire [10:0] _T_57651; // @[Modules.scala 78:156:@4629.4]
  wire [10:0] buffer_1_756; // @[Modules.scala 78:156:@4630.4]
  wire [11:0] _T_57653; // @[Modules.scala 78:156:@4632.4]
  wire [10:0] _T_57654; // @[Modules.scala 78:156:@4633.4]
  wire [10:0] buffer_1_757; // @[Modules.scala 78:156:@4634.4]
  wire [11:0] _T_57656; // @[Modules.scala 78:156:@4636.4]
  wire [10:0] _T_57657; // @[Modules.scala 78:156:@4637.4]
  wire [10:0] buffer_1_758; // @[Modules.scala 78:156:@4638.4]
  wire [11:0] _T_57659; // @[Modules.scala 78:156:@4640.4]
  wire [10:0] _T_57660; // @[Modules.scala 78:156:@4641.4]
  wire [10:0] buffer_1_759; // @[Modules.scala 78:156:@4642.4]
  wire [11:0] _T_57662; // @[Modules.scala 78:156:@4644.4]
  wire [10:0] _T_57663; // @[Modules.scala 78:156:@4645.4]
  wire [10:0] buffer_1_760; // @[Modules.scala 78:156:@4646.4]
  wire [11:0] _T_57665; // @[Modules.scala 78:156:@4648.4]
  wire [10:0] _T_57666; // @[Modules.scala 78:156:@4649.4]
  wire [10:0] buffer_1_761; // @[Modules.scala 78:156:@4650.4]
  wire [11:0] _T_57668; // @[Modules.scala 78:156:@4652.4]
  wire [10:0] _T_57669; // @[Modules.scala 78:156:@4653.4]
  wire [10:0] buffer_1_762; // @[Modules.scala 78:156:@4654.4]
  wire [11:0] _T_57671; // @[Modules.scala 78:156:@4656.4]
  wire [10:0] _T_57672; // @[Modules.scala 78:156:@4657.4]
  wire [10:0] buffer_1_763; // @[Modules.scala 78:156:@4658.4]
  wire [11:0] _T_57674; // @[Modules.scala 78:156:@4660.4]
  wire [10:0] _T_57675; // @[Modules.scala 78:156:@4661.4]
  wire [10:0] buffer_1_764; // @[Modules.scala 78:156:@4662.4]
  wire [11:0] _T_57677; // @[Modules.scala 78:156:@4664.4]
  wire [10:0] _T_57678; // @[Modules.scala 78:156:@4665.4]
  wire [10:0] buffer_1_765; // @[Modules.scala 78:156:@4666.4]
  wire [11:0] _T_57680; // @[Modules.scala 78:156:@4668.4]
  wire [10:0] _T_57681; // @[Modules.scala 78:156:@4669.4]
  wire [10:0] buffer_1_766; // @[Modules.scala 78:156:@4670.4]
  wire [11:0] _T_57683; // @[Modules.scala 78:156:@4672.4]
  wire [10:0] _T_57684; // @[Modules.scala 78:156:@4673.4]
  wire [10:0] buffer_1_767; // @[Modules.scala 78:156:@4674.4]
  wire [11:0] _T_57686; // @[Modules.scala 78:156:@4676.4]
  wire [10:0] _T_57687; // @[Modules.scala 78:156:@4677.4]
  wire [10:0] buffer_1_768; // @[Modules.scala 78:156:@4678.4]
  wire [11:0] _T_57689; // @[Modules.scala 78:156:@4680.4]
  wire [10:0] _T_57690; // @[Modules.scala 78:156:@4681.4]
  wire [10:0] buffer_1_769; // @[Modules.scala 78:156:@4682.4]
  wire [11:0] _T_57692; // @[Modules.scala 78:156:@4684.4]
  wire [10:0] _T_57693; // @[Modules.scala 78:156:@4685.4]
  wire [10:0] buffer_1_770; // @[Modules.scala 78:156:@4686.4]
  wire [11:0] _T_57695; // @[Modules.scala 78:156:@4688.4]
  wire [10:0] _T_57696; // @[Modules.scala 78:156:@4689.4]
  wire [10:0] buffer_1_771; // @[Modules.scala 78:156:@4690.4]
  wire [11:0] _T_57698; // @[Modules.scala 78:156:@4692.4]
  wire [10:0] _T_57699; // @[Modules.scala 78:156:@4693.4]
  wire [10:0] buffer_1_772; // @[Modules.scala 78:156:@4694.4]
  wire [11:0] _T_57701; // @[Modules.scala 78:156:@4696.4]
  wire [10:0] _T_57702; // @[Modules.scala 78:156:@4697.4]
  wire [10:0] buffer_1_773; // @[Modules.scala 78:156:@4698.4]
  wire [11:0] _T_57704; // @[Modules.scala 78:156:@4700.4]
  wire [10:0] _T_57705; // @[Modules.scala 78:156:@4701.4]
  wire [10:0] buffer_1_774; // @[Modules.scala 78:156:@4702.4]
  wire [11:0] _T_57707; // @[Modules.scala 78:156:@4704.4]
  wire [10:0] _T_57708; // @[Modules.scala 78:156:@4705.4]
  wire [10:0] buffer_1_775; // @[Modules.scala 78:156:@4706.4]
  wire [11:0] _T_57710; // @[Modules.scala 78:156:@4708.4]
  wire [10:0] _T_57711; // @[Modules.scala 78:156:@4709.4]
  wire [10:0] buffer_1_776; // @[Modules.scala 78:156:@4710.4]
  wire [11:0] _T_57713; // @[Modules.scala 78:156:@4712.4]
  wire [10:0] _T_57714; // @[Modules.scala 78:156:@4713.4]
  wire [10:0] buffer_1_777; // @[Modules.scala 78:156:@4714.4]
  wire [11:0] _T_57716; // @[Modules.scala 78:156:@4716.4]
  wire [10:0] _T_57717; // @[Modules.scala 78:156:@4717.4]
  wire [10:0] buffer_1_778; // @[Modules.scala 78:156:@4718.4]
  wire [11:0] _T_57719; // @[Modules.scala 78:156:@4720.4]
  wire [10:0] _T_57720; // @[Modules.scala 78:156:@4721.4]
  wire [10:0] buffer_1_779; // @[Modules.scala 78:156:@4722.4]
  wire [11:0] _T_57722; // @[Modules.scala 78:156:@4724.4]
  wire [10:0] _T_57723; // @[Modules.scala 78:156:@4725.4]
  wire [10:0] buffer_1_780; // @[Modules.scala 78:156:@4726.4]
  wire [11:0] _T_57725; // @[Modules.scala 78:156:@4728.4]
  wire [10:0] _T_57726; // @[Modules.scala 78:156:@4729.4]
  wire [10:0] buffer_1_781; // @[Modules.scala 78:156:@4730.4]
  wire [11:0] _T_57728; // @[Modules.scala 78:156:@4732.4]
  wire [10:0] _T_57729; // @[Modules.scala 78:156:@4733.4]
  wire [10:0] buffer_1_782; // @[Modules.scala 78:156:@4734.4]
  wire [11:0] _T_57731; // @[Modules.scala 78:156:@4736.4]
  wire [10:0] _T_57732; // @[Modules.scala 78:156:@4737.4]
  wire [10:0] buffer_1_783; // @[Modules.scala 78:156:@4738.4]
  wire [5:0] _T_57736; // @[Modules.scala 37:46:@4746.4]
  wire [4:0] _T_57737; // @[Modules.scala 37:46:@4747.4]
  wire [4:0] _T_57738; // @[Modules.scala 37:46:@4748.4]
  wire [5:0] _T_57741; // @[Modules.scala 37:46:@4755.4]
  wire [4:0] _T_57742; // @[Modules.scala 37:46:@4756.4]
  wire [4:0] _T_57743; // @[Modules.scala 37:46:@4757.4]
  wire [5:0] _T_57770; // @[Modules.scala 37:46:@4796.4]
  wire [4:0] _T_57771; // @[Modules.scala 37:46:@4797.4]
  wire [4:0] _T_57772; // @[Modules.scala 37:46:@4798.4]
  wire [5:0] _T_57793; // @[Modules.scala 37:46:@4830.4]
  wire [4:0] _T_57794; // @[Modules.scala 37:46:@4831.4]
  wire [4:0] _T_57795; // @[Modules.scala 37:46:@4832.4]
  wire [5:0] _T_57836; // @[Modules.scala 37:46:@4890.4]
  wire [4:0] _T_57837; // @[Modules.scala 37:46:@4891.4]
  wire [4:0] _T_57838; // @[Modules.scala 37:46:@4892.4]
  wire [5:0] _T_57842; // @[Modules.scala 37:46:@4898.4]
  wire [4:0] _T_57843; // @[Modules.scala 37:46:@4899.4]
  wire [4:0] _T_57844; // @[Modules.scala 37:46:@4900.4]
  wire [5:0] _T_57858; // @[Modules.scala 37:46:@4917.4]
  wire [4:0] _T_57859; // @[Modules.scala 37:46:@4918.4]
  wire [4:0] _T_57860; // @[Modules.scala 37:46:@4919.4]
  wire [5:0] _T_57861; // @[Modules.scala 37:46:@4921.4]
  wire [4:0] _T_57862; // @[Modules.scala 37:46:@4922.4]
  wire [4:0] _T_57863; // @[Modules.scala 37:46:@4923.4]
  wire [5:0] _T_57864; // @[Modules.scala 37:46:@4925.4]
  wire [4:0] _T_57865; // @[Modules.scala 37:46:@4926.4]
  wire [4:0] _T_57866; // @[Modules.scala 37:46:@4927.4]
  wire [5:0] _T_57876; // @[Modules.scala 37:46:@4941.4]
  wire [4:0] _T_57877; // @[Modules.scala 37:46:@4942.4]
  wire [4:0] _T_57878; // @[Modules.scala 37:46:@4943.4]
  wire [5:0] _T_57879; // @[Modules.scala 37:46:@4946.4]
  wire [4:0] _T_57880; // @[Modules.scala 37:46:@4947.4]
  wire [4:0] _T_57881; // @[Modules.scala 37:46:@4948.4]
  wire [5:0] _T_57885; // @[Modules.scala 37:46:@4954.4]
  wire [4:0] _T_57886; // @[Modules.scala 37:46:@4955.4]
  wire [4:0] _T_57887; // @[Modules.scala 37:46:@4956.4]
  wire [5:0] _T_57923; // @[Modules.scala 37:46:@5002.4]
  wire [4:0] _T_57924; // @[Modules.scala 37:46:@5003.4]
  wire [4:0] _T_57925; // @[Modules.scala 37:46:@5004.4]
  wire [5:0] _T_57926; // @[Modules.scala 37:46:@5006.4]
  wire [4:0] _T_57927; // @[Modules.scala 37:46:@5007.4]
  wire [4:0] _T_57928; // @[Modules.scala 37:46:@5008.4]
  wire [5:0] _T_57941; // @[Modules.scala 37:46:@5024.4]
  wire [4:0] _T_57942; // @[Modules.scala 37:46:@5025.4]
  wire [4:0] _T_57943; // @[Modules.scala 37:46:@5026.4]
  wire [5:0] _T_57999; // @[Modules.scala 37:46:@5107.4]
  wire [4:0] _T_58000; // @[Modules.scala 37:46:@5108.4]
  wire [4:0] _T_58001; // @[Modules.scala 37:46:@5109.4]
  wire [5:0] _T_58038; // @[Modules.scala 37:46:@5159.4]
  wire [4:0] _T_58039; // @[Modules.scala 37:46:@5160.4]
  wire [4:0] _T_58040; // @[Modules.scala 37:46:@5161.4]
  wire [5:0] _T_58066; // @[Modules.scala 37:46:@5196.4]
  wire [4:0] _T_58067; // @[Modules.scala 37:46:@5197.4]
  wire [4:0] _T_58068; // @[Modules.scala 37:46:@5198.4]
  wire [5:0] _T_58081; // @[Modules.scala 37:46:@5216.4]
  wire [4:0] _T_58082; // @[Modules.scala 37:46:@5217.4]
  wire [4:0] _T_58083; // @[Modules.scala 37:46:@5218.4]
  wire [5:0] _T_58089; // @[Modules.scala 37:46:@5228.4]
  wire [4:0] _T_58090; // @[Modules.scala 37:46:@5229.4]
  wire [4:0] _T_58091; // @[Modules.scala 37:46:@5230.4]
  wire [5:0] _T_58113; // @[Modules.scala 37:46:@5257.4]
  wire [4:0] _T_58114; // @[Modules.scala 37:46:@5258.4]
  wire [4:0] _T_58115; // @[Modules.scala 37:46:@5259.4]
  wire [5:0] _T_58126; // @[Modules.scala 37:46:@5278.4]
  wire [4:0] _T_58127; // @[Modules.scala 37:46:@5279.4]
  wire [4:0] _T_58128; // @[Modules.scala 37:46:@5280.4]
  wire [5:0] _T_58149; // @[Modules.scala 37:46:@5312.4]
  wire [4:0] _T_58150; // @[Modules.scala 37:46:@5313.4]
  wire [4:0] _T_58151; // @[Modules.scala 37:46:@5314.4]
  wire [5:0] _T_58156; // @[Modules.scala 37:46:@5324.4]
  wire [4:0] _T_58157; // @[Modules.scala 37:46:@5325.4]
  wire [4:0] _T_58158; // @[Modules.scala 37:46:@5326.4]
  wire [5:0] _T_58160; // @[Modules.scala 37:46:@5331.4]
  wire [4:0] _T_58161; // @[Modules.scala 37:46:@5332.4]
  wire [4:0] _T_58162; // @[Modules.scala 37:46:@5333.4]
  wire [5:0] _T_58172; // @[Modules.scala 37:46:@5346.4]
  wire [4:0] _T_58173; // @[Modules.scala 37:46:@5347.4]
  wire [4:0] _T_58174; // @[Modules.scala 37:46:@5348.4]
  wire [5:0] _T_58189; // @[Modules.scala 37:46:@5374.4]
  wire [4:0] _T_58190; // @[Modules.scala 37:46:@5375.4]
  wire [4:0] _T_58191; // @[Modules.scala 37:46:@5376.4]
  wire [5:0] _T_58202; // @[Modules.scala 37:46:@5391.4]
  wire [4:0] _T_58203; // @[Modules.scala 37:46:@5392.4]
  wire [4:0] _T_58204; // @[Modules.scala 37:46:@5393.4]
  wire [5:0] _T_58237; // @[Modules.scala 37:46:@5438.4]
  wire [4:0] _T_58238; // @[Modules.scala 37:46:@5439.4]
  wire [4:0] _T_58239; // @[Modules.scala 37:46:@5440.4]
  wire [5:0] _T_58240; // @[Modules.scala 37:46:@5442.4]
  wire [4:0] _T_58241; // @[Modules.scala 37:46:@5443.4]
  wire [4:0] _T_58242; // @[Modules.scala 37:46:@5444.4]
  wire [10:0] buffer_2_2; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58269; // @[Modules.scala 65:57:@5482.4]
  wire [10:0] _T_58270; // @[Modules.scala 65:57:@5483.4]
  wire [10:0] buffer_2_393; // @[Modules.scala 65:57:@5484.4]
  wire [10:0] buffer_2_4; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58272; // @[Modules.scala 65:57:@5486.4]
  wire [10:0] _T_58273; // @[Modules.scala 65:57:@5487.4]
  wire [10:0] buffer_2_394; // @[Modules.scala 65:57:@5488.4]
  wire [10:0] buffer_2_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58278; // @[Modules.scala 65:57:@5494.4]
  wire [10:0] _T_58279; // @[Modules.scala 65:57:@5495.4]
  wire [10:0] buffer_2_396; // @[Modules.scala 65:57:@5496.4]
  wire [10:0] buffer_2_10; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_11; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58281; // @[Modules.scala 65:57:@5498.4]
  wire [10:0] _T_58282; // @[Modules.scala 65:57:@5499.4]
  wire [10:0] buffer_2_397; // @[Modules.scala 65:57:@5500.4]
  wire [11:0] _T_58284; // @[Modules.scala 65:57:@5502.4]
  wire [10:0] _T_58285; // @[Modules.scala 65:57:@5503.4]
  wire [10:0] buffer_2_398; // @[Modules.scala 65:57:@5504.4]
  wire [10:0] buffer_2_15; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58287; // @[Modules.scala 65:57:@5506.4]
  wire [10:0] _T_58288; // @[Modules.scala 65:57:@5507.4]
  wire [10:0] buffer_2_399; // @[Modules.scala 65:57:@5508.4]
  wire [11:0] _T_58290; // @[Modules.scala 65:57:@5510.4]
  wire [10:0] _T_58291; // @[Modules.scala 65:57:@5511.4]
  wire [10:0] buffer_2_400; // @[Modules.scala 65:57:@5512.4]
  wire [10:0] buffer_2_20; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58296; // @[Modules.scala 65:57:@5518.4]
  wire [10:0] _T_58297; // @[Modules.scala 65:57:@5519.4]
  wire [10:0] buffer_2_402; // @[Modules.scala 65:57:@5520.4]
  wire [11:0] _T_58299; // @[Modules.scala 65:57:@5522.4]
  wire [10:0] _T_58300; // @[Modules.scala 65:57:@5523.4]
  wire [10:0] buffer_2_403; // @[Modules.scala 65:57:@5524.4]
  wire [11:0] _T_58305; // @[Modules.scala 65:57:@5530.4]
  wire [10:0] _T_58306; // @[Modules.scala 65:57:@5531.4]
  wire [10:0] buffer_2_405; // @[Modules.scala 65:57:@5532.4]
  wire [10:0] buffer_2_28; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58308; // @[Modules.scala 65:57:@5534.4]
  wire [10:0] _T_58309; // @[Modules.scala 65:57:@5535.4]
  wire [10:0] buffer_2_406; // @[Modules.scala 65:57:@5536.4]
  wire [10:0] buffer_2_31; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58311; // @[Modules.scala 65:57:@5538.4]
  wire [10:0] _T_58312; // @[Modules.scala 65:57:@5539.4]
  wire [10:0] buffer_2_407; // @[Modules.scala 65:57:@5540.4]
  wire [10:0] buffer_2_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58317; // @[Modules.scala 65:57:@5546.4]
  wire [10:0] _T_58318; // @[Modules.scala 65:57:@5547.4]
  wire [10:0] buffer_2_409; // @[Modules.scala 65:57:@5548.4]
  wire [10:0] buffer_2_39; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58323; // @[Modules.scala 65:57:@5554.4]
  wire [10:0] _T_58324; // @[Modules.scala 65:57:@5555.4]
  wire [10:0] buffer_2_411; // @[Modules.scala 65:57:@5556.4]
  wire [10:0] buffer_2_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58326; // @[Modules.scala 65:57:@5558.4]
  wire [10:0] _T_58327; // @[Modules.scala 65:57:@5559.4]
  wire [10:0] buffer_2_412; // @[Modules.scala 65:57:@5560.4]
  wire [11:0] _T_58329; // @[Modules.scala 65:57:@5562.4]
  wire [10:0] _T_58330; // @[Modules.scala 65:57:@5563.4]
  wire [10:0] buffer_2_413; // @[Modules.scala 65:57:@5564.4]
  wire [10:0] buffer_2_44; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58332; // @[Modules.scala 65:57:@5566.4]
  wire [10:0] _T_58333; // @[Modules.scala 65:57:@5567.4]
  wire [10:0] buffer_2_414; // @[Modules.scala 65:57:@5568.4]
  wire [11:0] _T_58335; // @[Modules.scala 65:57:@5570.4]
  wire [10:0] _T_58336; // @[Modules.scala 65:57:@5571.4]
  wire [10:0] buffer_2_415; // @[Modules.scala 65:57:@5572.4]
  wire [10:0] buffer_2_50; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58341; // @[Modules.scala 65:57:@5578.4]
  wire [10:0] _T_58342; // @[Modules.scala 65:57:@5579.4]
  wire [10:0] buffer_2_417; // @[Modules.scala 65:57:@5580.4]
  wire [11:0] _T_58362; // @[Modules.scala 65:57:@5606.4]
  wire [10:0] _T_58363; // @[Modules.scala 65:57:@5607.4]
  wire [10:0] buffer_2_424; // @[Modules.scala 65:57:@5608.4]
  wire [10:0] buffer_2_70; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58371; // @[Modules.scala 65:57:@5618.4]
  wire [10:0] _T_58372; // @[Modules.scala 65:57:@5619.4]
  wire [10:0] buffer_2_427; // @[Modules.scala 65:57:@5620.4]
  wire [10:0] buffer_2_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58383; // @[Modules.scala 65:57:@5634.4]
  wire [10:0] _T_58384; // @[Modules.scala 65:57:@5635.4]
  wire [10:0] buffer_2_431; // @[Modules.scala 65:57:@5636.4]
  wire [10:0] buffer_2_80; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58386; // @[Modules.scala 65:57:@5638.4]
  wire [10:0] _T_58387; // @[Modules.scala 65:57:@5639.4]
  wire [10:0] buffer_2_432; // @[Modules.scala 65:57:@5640.4]
  wire [10:0] buffer_2_82; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58389; // @[Modules.scala 65:57:@5642.4]
  wire [10:0] _T_58390; // @[Modules.scala 65:57:@5643.4]
  wire [10:0] buffer_2_433; // @[Modules.scala 65:57:@5644.4]
  wire [10:0] buffer_2_84; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58392; // @[Modules.scala 65:57:@5646.4]
  wire [10:0] _T_58393; // @[Modules.scala 65:57:@5647.4]
  wire [10:0] buffer_2_434; // @[Modules.scala 65:57:@5648.4]
  wire [10:0] buffer_2_95; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58407; // @[Modules.scala 65:57:@5666.4]
  wire [10:0] _T_58408; // @[Modules.scala 65:57:@5667.4]
  wire [10:0] buffer_2_439; // @[Modules.scala 65:57:@5668.4]
  wire [10:0] buffer_2_96; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58410; // @[Modules.scala 65:57:@5670.4]
  wire [10:0] _T_58411; // @[Modules.scala 65:57:@5671.4]
  wire [10:0] buffer_2_440; // @[Modules.scala 65:57:@5672.4]
  wire [11:0] _T_58413; // @[Modules.scala 65:57:@5674.4]
  wire [10:0] _T_58414; // @[Modules.scala 65:57:@5675.4]
  wire [10:0] buffer_2_441; // @[Modules.scala 65:57:@5676.4]
  wire [11:0] _T_58422; // @[Modules.scala 65:57:@5686.4]
  wire [10:0] _T_58423; // @[Modules.scala 65:57:@5687.4]
  wire [10:0] buffer_2_444; // @[Modules.scala 65:57:@5688.4]
  wire [10:0] buffer_2_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58425; // @[Modules.scala 65:57:@5690.4]
  wire [10:0] _T_58426; // @[Modules.scala 65:57:@5691.4]
  wire [10:0] buffer_2_445; // @[Modules.scala 65:57:@5692.4]
  wire [10:0] buffer_2_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58428; // @[Modules.scala 65:57:@5694.4]
  wire [10:0] _T_58429; // @[Modules.scala 65:57:@5695.4]
  wire [10:0] buffer_2_446; // @[Modules.scala 65:57:@5696.4]
  wire [10:0] buffer_2_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58431; // @[Modules.scala 65:57:@5698.4]
  wire [10:0] _T_58432; // @[Modules.scala 65:57:@5699.4]
  wire [10:0] buffer_2_447; // @[Modules.scala 65:57:@5700.4]
  wire [10:0] buffer_2_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58440; // @[Modules.scala 65:57:@5710.4]
  wire [10:0] _T_58441; // @[Modules.scala 65:57:@5711.4]
  wire [10:0] buffer_2_450; // @[Modules.scala 65:57:@5712.4]
  wire [10:0] buffer_2_130; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58461; // @[Modules.scala 65:57:@5738.4]
  wire [10:0] _T_58462; // @[Modules.scala 65:57:@5739.4]
  wire [10:0] buffer_2_457; // @[Modules.scala 65:57:@5740.4]
  wire [10:0] buffer_2_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58479; // @[Modules.scala 65:57:@5762.4]
  wire [10:0] _T_58480; // @[Modules.scala 65:57:@5763.4]
  wire [10:0] buffer_2_463; // @[Modules.scala 65:57:@5764.4]
  wire [10:0] buffer_2_144; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58482; // @[Modules.scala 65:57:@5766.4]
  wire [10:0] _T_58483; // @[Modules.scala 65:57:@5767.4]
  wire [10:0] buffer_2_464; // @[Modules.scala 65:57:@5768.4]
  wire [10:0] buffer_2_152; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58494; // @[Modules.scala 65:57:@5782.4]
  wire [10:0] _T_58495; // @[Modules.scala 65:57:@5783.4]
  wire [10:0] buffer_2_468; // @[Modules.scala 65:57:@5784.4]
  wire [10:0] buffer_2_157; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58500; // @[Modules.scala 65:57:@5790.4]
  wire [10:0] _T_58501; // @[Modules.scala 65:57:@5791.4]
  wire [10:0] buffer_2_470; // @[Modules.scala 65:57:@5792.4]
  wire [10:0] buffer_2_160; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58506; // @[Modules.scala 65:57:@5798.4]
  wire [10:0] _T_58507; // @[Modules.scala 65:57:@5799.4]
  wire [10:0] buffer_2_472; // @[Modules.scala 65:57:@5800.4]
  wire [10:0] buffer_2_166; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58515; // @[Modules.scala 65:57:@5810.4]
  wire [10:0] _T_58516; // @[Modules.scala 65:57:@5811.4]
  wire [10:0] buffer_2_475; // @[Modules.scala 65:57:@5812.4]
  wire [10:0] buffer_2_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58530; // @[Modules.scala 65:57:@5830.4]
  wire [10:0] _T_58531; // @[Modules.scala 65:57:@5831.4]
  wire [10:0] buffer_2_480; // @[Modules.scala 65:57:@5832.4]
  wire [10:0] buffer_2_180; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58536; // @[Modules.scala 65:57:@5838.4]
  wire [10:0] _T_58537; // @[Modules.scala 65:57:@5839.4]
  wire [10:0] buffer_2_482; // @[Modules.scala 65:57:@5840.4]
  wire [10:0] buffer_2_192; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58554; // @[Modules.scala 65:57:@5862.4]
  wire [10:0] _T_58555; // @[Modules.scala 65:57:@5863.4]
  wire [10:0] buffer_2_488; // @[Modules.scala 65:57:@5864.4]
  wire [10:0] buffer_2_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58572; // @[Modules.scala 65:57:@5886.4]
  wire [10:0] _T_58573; // @[Modules.scala 65:57:@5887.4]
  wire [10:0] buffer_2_494; // @[Modules.scala 65:57:@5888.4]
  wire [10:0] buffer_2_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58581; // @[Modules.scala 65:57:@5898.4]
  wire [10:0] _T_58582; // @[Modules.scala 65:57:@5899.4]
  wire [10:0] buffer_2_497; // @[Modules.scala 65:57:@5900.4]
  wire [11:0] _T_58584; // @[Modules.scala 65:57:@5902.4]
  wire [10:0] _T_58585; // @[Modules.scala 65:57:@5903.4]
  wire [10:0] buffer_2_498; // @[Modules.scala 65:57:@5904.4]
  wire [11:0] _T_58587; // @[Modules.scala 65:57:@5906.4]
  wire [10:0] _T_58588; // @[Modules.scala 65:57:@5907.4]
  wire [10:0] buffer_2_499; // @[Modules.scala 65:57:@5908.4]
  wire [11:0] _T_58596; // @[Modules.scala 65:57:@5918.4]
  wire [10:0] _T_58597; // @[Modules.scala 65:57:@5919.4]
  wire [10:0] buffer_2_502; // @[Modules.scala 65:57:@5920.4]
  wire [11:0] _T_58602; // @[Modules.scala 65:57:@5926.4]
  wire [10:0] _T_58603; // @[Modules.scala 65:57:@5927.4]
  wire [10:0] buffer_2_504; // @[Modules.scala 65:57:@5928.4]
  wire [10:0] buffer_2_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58605; // @[Modules.scala 65:57:@5930.4]
  wire [10:0] _T_58606; // @[Modules.scala 65:57:@5931.4]
  wire [10:0] buffer_2_505; // @[Modules.scala 65:57:@5932.4]
  wire [10:0] buffer_2_228; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58608; // @[Modules.scala 65:57:@5934.4]
  wire [10:0] _T_58609; // @[Modules.scala 65:57:@5935.4]
  wire [10:0] buffer_2_506; // @[Modules.scala 65:57:@5936.4]
  wire [10:0] buffer_2_230; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58611; // @[Modules.scala 65:57:@5938.4]
  wire [10:0] _T_58612; // @[Modules.scala 65:57:@5939.4]
  wire [10:0] buffer_2_507; // @[Modules.scala 65:57:@5940.4]
  wire [10:0] buffer_2_232; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58614; // @[Modules.scala 65:57:@5942.4]
  wire [10:0] _T_58615; // @[Modules.scala 65:57:@5943.4]
  wire [10:0] buffer_2_508; // @[Modules.scala 65:57:@5944.4]
  wire [11:0] _T_58617; // @[Modules.scala 65:57:@5946.4]
  wire [10:0] _T_58618; // @[Modules.scala 65:57:@5947.4]
  wire [10:0] buffer_2_509; // @[Modules.scala 65:57:@5948.4]
  wire [10:0] buffer_2_238; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58623; // @[Modules.scala 65:57:@5954.4]
  wire [10:0] _T_58624; // @[Modules.scala 65:57:@5955.4]
  wire [10:0] buffer_2_511; // @[Modules.scala 65:57:@5956.4]
  wire [10:0] buffer_2_242; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58629; // @[Modules.scala 65:57:@5962.4]
  wire [10:0] _T_58630; // @[Modules.scala 65:57:@5963.4]
  wire [10:0] buffer_2_513; // @[Modules.scala 65:57:@5964.4]
  wire [10:0] buffer_2_244; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58632; // @[Modules.scala 65:57:@5966.4]
  wire [10:0] _T_58633; // @[Modules.scala 65:57:@5967.4]
  wire [10:0] buffer_2_514; // @[Modules.scala 65:57:@5968.4]
  wire [11:0] _T_58638; // @[Modules.scala 65:57:@5974.4]
  wire [10:0] _T_58639; // @[Modules.scala 65:57:@5975.4]
  wire [10:0] buffer_2_516; // @[Modules.scala 65:57:@5976.4]
  wire [10:0] buffer_2_258; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58653; // @[Modules.scala 65:57:@5994.4]
  wire [10:0] _T_58654; // @[Modules.scala 65:57:@5995.4]
  wire [10:0] buffer_2_521; // @[Modules.scala 65:57:@5996.4]
  wire [11:0] _T_58656; // @[Modules.scala 65:57:@5998.4]
  wire [10:0] _T_58657; // @[Modules.scala 65:57:@5999.4]
  wire [10:0] buffer_2_522; // @[Modules.scala 65:57:@6000.4]
  wire [10:0] buffer_2_272; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58674; // @[Modules.scala 65:57:@6022.4]
  wire [10:0] _T_58675; // @[Modules.scala 65:57:@6023.4]
  wire [10:0] buffer_2_528; // @[Modules.scala 65:57:@6024.4]
  wire [10:0] buffer_2_274; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_275; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58677; // @[Modules.scala 65:57:@6026.4]
  wire [10:0] _T_58678; // @[Modules.scala 65:57:@6027.4]
  wire [10:0] buffer_2_529; // @[Modules.scala 65:57:@6028.4]
  wire [10:0] buffer_2_276; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58680; // @[Modules.scala 65:57:@6030.4]
  wire [10:0] _T_58681; // @[Modules.scala 65:57:@6031.4]
  wire [10:0] buffer_2_530; // @[Modules.scala 65:57:@6032.4]
  wire [11:0] _T_58683; // @[Modules.scala 65:57:@6034.4]
  wire [10:0] _T_58684; // @[Modules.scala 65:57:@6035.4]
  wire [10:0] buffer_2_531; // @[Modules.scala 65:57:@6036.4]
  wire [10:0] buffer_2_280; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58686; // @[Modules.scala 65:57:@6038.4]
  wire [10:0] _T_58687; // @[Modules.scala 65:57:@6039.4]
  wire [10:0] buffer_2_532; // @[Modules.scala 65:57:@6040.4]
  wire [11:0] _T_58695; // @[Modules.scala 65:57:@6050.4]
  wire [10:0] _T_58696; // @[Modules.scala 65:57:@6051.4]
  wire [10:0] buffer_2_535; // @[Modules.scala 65:57:@6052.4]
  wire [11:0] _T_58698; // @[Modules.scala 65:57:@6054.4]
  wire [10:0] _T_58699; // @[Modules.scala 65:57:@6055.4]
  wire [10:0] buffer_2_536; // @[Modules.scala 65:57:@6056.4]
  wire [10:0] buffer_2_294; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_295; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58707; // @[Modules.scala 65:57:@6066.4]
  wire [10:0] _T_58708; // @[Modules.scala 65:57:@6067.4]
  wire [10:0] buffer_2_539; // @[Modules.scala 65:57:@6068.4]
  wire [10:0] buffer_2_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58710; // @[Modules.scala 65:57:@6070.4]
  wire [10:0] _T_58711; // @[Modules.scala 65:57:@6071.4]
  wire [10:0] buffer_2_540; // @[Modules.scala 65:57:@6072.4]
  wire [10:0] buffer_2_298; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58713; // @[Modules.scala 65:57:@6074.4]
  wire [10:0] _T_58714; // @[Modules.scala 65:57:@6075.4]
  wire [10:0] buffer_2_541; // @[Modules.scala 65:57:@6076.4]
  wire [10:0] buffer_2_300; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58716; // @[Modules.scala 65:57:@6078.4]
  wire [10:0] _T_58717; // @[Modules.scala 65:57:@6079.4]
  wire [10:0] buffer_2_542; // @[Modules.scala 65:57:@6080.4]
  wire [10:0] buffer_2_302; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58719; // @[Modules.scala 65:57:@6082.4]
  wire [10:0] _T_58720; // @[Modules.scala 65:57:@6083.4]
  wire [10:0] buffer_2_543; // @[Modules.scala 65:57:@6084.4]
  wire [10:0] buffer_2_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58722; // @[Modules.scala 65:57:@6086.4]
  wire [10:0] _T_58723; // @[Modules.scala 65:57:@6087.4]
  wire [10:0] buffer_2_544; // @[Modules.scala 65:57:@6088.4]
  wire [10:0] buffer_2_308; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58728; // @[Modules.scala 65:57:@6094.4]
  wire [10:0] _T_58729; // @[Modules.scala 65:57:@6095.4]
  wire [10:0] buffer_2_546; // @[Modules.scala 65:57:@6096.4]
  wire [10:0] buffer_2_312; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58734; // @[Modules.scala 65:57:@6102.4]
  wire [10:0] _T_58735; // @[Modules.scala 65:57:@6103.4]
  wire [10:0] buffer_2_548; // @[Modules.scala 65:57:@6104.4]
  wire [10:0] buffer_2_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58740; // @[Modules.scala 65:57:@6110.4]
  wire [10:0] _T_58741; // @[Modules.scala 65:57:@6111.4]
  wire [10:0] buffer_2_550; // @[Modules.scala 65:57:@6112.4]
  wire [10:0] buffer_2_322; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_323; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58749; // @[Modules.scala 65:57:@6122.4]
  wire [10:0] _T_58750; // @[Modules.scala 65:57:@6123.4]
  wire [10:0] buffer_2_553; // @[Modules.scala 65:57:@6124.4]
  wire [10:0] buffer_2_324; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58752; // @[Modules.scala 65:57:@6126.4]
  wire [10:0] _T_58753; // @[Modules.scala 65:57:@6127.4]
  wire [10:0] buffer_2_554; // @[Modules.scala 65:57:@6128.4]
  wire [11:0] _T_58755; // @[Modules.scala 65:57:@6130.4]
  wire [10:0] _T_58756; // @[Modules.scala 65:57:@6131.4]
  wire [10:0] buffer_2_555; // @[Modules.scala 65:57:@6132.4]
  wire [10:0] buffer_2_328; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58758; // @[Modules.scala 65:57:@6134.4]
  wire [10:0] _T_58759; // @[Modules.scala 65:57:@6135.4]
  wire [10:0] buffer_2_556; // @[Modules.scala 65:57:@6136.4]
  wire [10:0] buffer_2_330; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58761; // @[Modules.scala 65:57:@6138.4]
  wire [10:0] _T_58762; // @[Modules.scala 65:57:@6139.4]
  wire [10:0] buffer_2_557; // @[Modules.scala 65:57:@6140.4]
  wire [10:0] buffer_2_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58767; // @[Modules.scala 65:57:@6146.4]
  wire [10:0] _T_58768; // @[Modules.scala 65:57:@6147.4]
  wire [10:0] buffer_2_559; // @[Modules.scala 65:57:@6148.4]
  wire [11:0] _T_58770; // @[Modules.scala 65:57:@6150.4]
  wire [10:0] _T_58771; // @[Modules.scala 65:57:@6151.4]
  wire [10:0] buffer_2_560; // @[Modules.scala 65:57:@6152.4]
  wire [10:0] buffer_2_342; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58779; // @[Modules.scala 65:57:@6162.4]
  wire [10:0] _T_58780; // @[Modules.scala 65:57:@6163.4]
  wire [10:0] buffer_2_563; // @[Modules.scala 65:57:@6164.4]
  wire [10:0] buffer_2_344; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58782; // @[Modules.scala 65:57:@6166.4]
  wire [10:0] _T_58783; // @[Modules.scala 65:57:@6167.4]
  wire [10:0] buffer_2_564; // @[Modules.scala 65:57:@6168.4]
  wire [11:0] _T_58788; // @[Modules.scala 65:57:@6174.4]
  wire [10:0] _T_58789; // @[Modules.scala 65:57:@6175.4]
  wire [10:0] buffer_2_566; // @[Modules.scala 65:57:@6176.4]
  wire [11:0] _T_58791; // @[Modules.scala 65:57:@6178.4]
  wire [10:0] _T_58792; // @[Modules.scala 65:57:@6179.4]
  wire [10:0] buffer_2_567; // @[Modules.scala 65:57:@6180.4]
  wire [10:0] buffer_2_364; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58812; // @[Modules.scala 65:57:@6206.4]
  wire [10:0] _T_58813; // @[Modules.scala 65:57:@6207.4]
  wire [10:0] buffer_2_574; // @[Modules.scala 65:57:@6208.4]
  wire [10:0] buffer_2_366; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58815; // @[Modules.scala 65:57:@6210.4]
  wire [10:0] _T_58816; // @[Modules.scala 65:57:@6211.4]
  wire [10:0] buffer_2_575; // @[Modules.scala 65:57:@6212.4]
  wire [10:0] buffer_2_374; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_2_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58827; // @[Modules.scala 65:57:@6226.4]
  wire [10:0] _T_58828; // @[Modules.scala 65:57:@6227.4]
  wire [10:0] buffer_2_579; // @[Modules.scala 65:57:@6228.4]
  wire [10:0] buffer_2_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58830; // @[Modules.scala 65:57:@6230.4]
  wire [10:0] _T_58831; // @[Modules.scala 65:57:@6231.4]
  wire [10:0] buffer_2_580; // @[Modules.scala 65:57:@6232.4]
  wire [11:0] _T_58833; // @[Modules.scala 65:57:@6234.4]
  wire [10:0] _T_58834; // @[Modules.scala 65:57:@6235.4]
  wire [10:0] buffer_2_581; // @[Modules.scala 65:57:@6236.4]
  wire [10:0] buffer_2_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_58851; // @[Modules.scala 65:57:@6258.4]
  wire [10:0] _T_58852; // @[Modules.scala 65:57:@6259.4]
  wire [10:0] buffer_2_587; // @[Modules.scala 65:57:@6260.4]
  wire [11:0] _T_58854; // @[Modules.scala 68:83:@6262.4]
  wire [10:0] _T_58855; // @[Modules.scala 68:83:@6263.4]
  wire [10:0] buffer_2_588; // @[Modules.scala 68:83:@6264.4]
  wire [11:0] _T_58857; // @[Modules.scala 68:83:@6266.4]
  wire [10:0] _T_58858; // @[Modules.scala 68:83:@6267.4]
  wire [10:0] buffer_2_589; // @[Modules.scala 68:83:@6268.4]
  wire [11:0] _T_58860; // @[Modules.scala 68:83:@6270.4]
  wire [10:0] _T_58861; // @[Modules.scala 68:83:@6271.4]
  wire [10:0] buffer_2_590; // @[Modules.scala 68:83:@6272.4]
  wire [11:0] _T_58863; // @[Modules.scala 68:83:@6274.4]
  wire [10:0] _T_58864; // @[Modules.scala 68:83:@6275.4]
  wire [10:0] buffer_2_591; // @[Modules.scala 68:83:@6276.4]
  wire [11:0] _T_58866; // @[Modules.scala 68:83:@6278.4]
  wire [10:0] _T_58867; // @[Modules.scala 68:83:@6279.4]
  wire [10:0] buffer_2_592; // @[Modules.scala 68:83:@6280.4]
  wire [11:0] _T_58869; // @[Modules.scala 68:83:@6282.4]
  wire [10:0] _T_58870; // @[Modules.scala 68:83:@6283.4]
  wire [10:0] buffer_2_593; // @[Modules.scala 68:83:@6284.4]
  wire [11:0] _T_58872; // @[Modules.scala 68:83:@6286.4]
  wire [10:0] _T_58873; // @[Modules.scala 68:83:@6287.4]
  wire [10:0] buffer_2_594; // @[Modules.scala 68:83:@6288.4]
  wire [11:0] _T_58875; // @[Modules.scala 68:83:@6290.4]
  wire [10:0] _T_58876; // @[Modules.scala 68:83:@6291.4]
  wire [10:0] buffer_2_595; // @[Modules.scala 68:83:@6292.4]
  wire [11:0] _T_58878; // @[Modules.scala 68:83:@6294.4]
  wire [10:0] _T_58879; // @[Modules.scala 68:83:@6295.4]
  wire [10:0] buffer_2_596; // @[Modules.scala 68:83:@6296.4]
  wire [11:0] _T_58881; // @[Modules.scala 68:83:@6298.4]
  wire [10:0] _T_58882; // @[Modules.scala 68:83:@6299.4]
  wire [10:0] buffer_2_597; // @[Modules.scala 68:83:@6300.4]
  wire [11:0] _T_58884; // @[Modules.scala 68:83:@6302.4]
  wire [10:0] _T_58885; // @[Modules.scala 68:83:@6303.4]
  wire [10:0] buffer_2_598; // @[Modules.scala 68:83:@6304.4]
  wire [11:0] _T_58887; // @[Modules.scala 68:83:@6306.4]
  wire [10:0] _T_58888; // @[Modules.scala 68:83:@6307.4]
  wire [10:0] buffer_2_599; // @[Modules.scala 68:83:@6308.4]
  wire [11:0] _T_58890; // @[Modules.scala 68:83:@6310.4]
  wire [10:0] _T_58891; // @[Modules.scala 68:83:@6311.4]
  wire [10:0] buffer_2_600; // @[Modules.scala 68:83:@6312.4]
  wire [11:0] _T_58893; // @[Modules.scala 68:83:@6314.4]
  wire [10:0] _T_58894; // @[Modules.scala 68:83:@6315.4]
  wire [10:0] buffer_2_601; // @[Modules.scala 68:83:@6316.4]
  wire [11:0] _T_58896; // @[Modules.scala 68:83:@6318.4]
  wire [10:0] _T_58897; // @[Modules.scala 68:83:@6319.4]
  wire [10:0] buffer_2_602; // @[Modules.scala 68:83:@6320.4]
  wire [11:0] _T_58902; // @[Modules.scala 68:83:@6326.4]
  wire [10:0] _T_58903; // @[Modules.scala 68:83:@6327.4]
  wire [10:0] buffer_2_604; // @[Modules.scala 68:83:@6328.4]
  wire [11:0] _T_58905; // @[Modules.scala 68:83:@6330.4]
  wire [10:0] _T_58906; // @[Modules.scala 68:83:@6331.4]
  wire [10:0] buffer_2_605; // @[Modules.scala 68:83:@6332.4]
  wire [11:0] _T_58911; // @[Modules.scala 68:83:@6338.4]
  wire [10:0] _T_58912; // @[Modules.scala 68:83:@6339.4]
  wire [10:0] buffer_2_607; // @[Modules.scala 68:83:@6340.4]
  wire [11:0] _T_58914; // @[Modules.scala 68:83:@6342.4]
  wire [10:0] _T_58915; // @[Modules.scala 68:83:@6343.4]
  wire [10:0] buffer_2_608; // @[Modules.scala 68:83:@6344.4]
  wire [11:0] _T_58917; // @[Modules.scala 68:83:@6346.4]
  wire [10:0] _T_58918; // @[Modules.scala 68:83:@6347.4]
  wire [10:0] buffer_2_609; // @[Modules.scala 68:83:@6348.4]
  wire [11:0] _T_58923; // @[Modules.scala 68:83:@6354.4]
  wire [10:0] _T_58924; // @[Modules.scala 68:83:@6355.4]
  wire [10:0] buffer_2_611; // @[Modules.scala 68:83:@6356.4]
  wire [11:0] _T_58926; // @[Modules.scala 68:83:@6358.4]
  wire [10:0] _T_58927; // @[Modules.scala 68:83:@6359.4]
  wire [10:0] buffer_2_612; // @[Modules.scala 68:83:@6360.4]
  wire [11:0] _T_58932; // @[Modules.scala 68:83:@6366.4]
  wire [10:0] _T_58933; // @[Modules.scala 68:83:@6367.4]
  wire [10:0] buffer_2_614; // @[Modules.scala 68:83:@6368.4]
  wire [11:0] _T_58935; // @[Modules.scala 68:83:@6370.4]
  wire [10:0] _T_58936; // @[Modules.scala 68:83:@6371.4]
  wire [10:0] buffer_2_615; // @[Modules.scala 68:83:@6372.4]
  wire [11:0] _T_58941; // @[Modules.scala 68:83:@6378.4]
  wire [10:0] _T_58942; // @[Modules.scala 68:83:@6379.4]
  wire [10:0] buffer_2_617; // @[Modules.scala 68:83:@6380.4]
  wire [11:0] _T_58944; // @[Modules.scala 68:83:@6382.4]
  wire [10:0] _T_58945; // @[Modules.scala 68:83:@6383.4]
  wire [10:0] buffer_2_618; // @[Modules.scala 68:83:@6384.4]
  wire [11:0] _T_58947; // @[Modules.scala 68:83:@6386.4]
  wire [10:0] _T_58948; // @[Modules.scala 68:83:@6387.4]
  wire [10:0] buffer_2_619; // @[Modules.scala 68:83:@6388.4]
  wire [11:0] _T_58950; // @[Modules.scala 68:83:@6390.4]
  wire [10:0] _T_58951; // @[Modules.scala 68:83:@6391.4]
  wire [10:0] buffer_2_620; // @[Modules.scala 68:83:@6392.4]
  wire [11:0] _T_58956; // @[Modules.scala 68:83:@6398.4]
  wire [10:0] _T_58957; // @[Modules.scala 68:83:@6399.4]
  wire [10:0] buffer_2_622; // @[Modules.scala 68:83:@6400.4]
  wire [11:0] _T_58959; // @[Modules.scala 68:83:@6402.4]
  wire [10:0] _T_58960; // @[Modules.scala 68:83:@6403.4]
  wire [10:0] buffer_2_623; // @[Modules.scala 68:83:@6404.4]
  wire [11:0] _T_58962; // @[Modules.scala 68:83:@6406.4]
  wire [10:0] _T_58963; // @[Modules.scala 68:83:@6407.4]
  wire [10:0] buffer_2_624; // @[Modules.scala 68:83:@6408.4]
  wire [11:0] _T_58968; // @[Modules.scala 68:83:@6414.4]
  wire [10:0] _T_58969; // @[Modules.scala 68:83:@6415.4]
  wire [10:0] buffer_2_626; // @[Modules.scala 68:83:@6416.4]
  wire [11:0] _T_58971; // @[Modules.scala 68:83:@6418.4]
  wire [10:0] _T_58972; // @[Modules.scala 68:83:@6419.4]
  wire [10:0] buffer_2_627; // @[Modules.scala 68:83:@6420.4]
  wire [11:0] _T_58974; // @[Modules.scala 68:83:@6422.4]
  wire [10:0] _T_58975; // @[Modules.scala 68:83:@6423.4]
  wire [10:0] buffer_2_628; // @[Modules.scala 68:83:@6424.4]
  wire [11:0] _T_58977; // @[Modules.scala 68:83:@6426.4]
  wire [10:0] _T_58978; // @[Modules.scala 68:83:@6427.4]
  wire [10:0] buffer_2_629; // @[Modules.scala 68:83:@6428.4]
  wire [11:0] _T_58986; // @[Modules.scala 68:83:@6438.4]
  wire [10:0] _T_58987; // @[Modules.scala 68:83:@6439.4]
  wire [10:0] buffer_2_632; // @[Modules.scala 68:83:@6440.4]
  wire [11:0] _T_58989; // @[Modules.scala 68:83:@6442.4]
  wire [10:0] _T_58990; // @[Modules.scala 68:83:@6443.4]
  wire [10:0] buffer_2_633; // @[Modules.scala 68:83:@6444.4]
  wire [11:0] _T_58998; // @[Modules.scala 68:83:@6454.4]
  wire [10:0] _T_58999; // @[Modules.scala 68:83:@6455.4]
  wire [10:0] buffer_2_636; // @[Modules.scala 68:83:@6456.4]
  wire [11:0] _T_59001; // @[Modules.scala 68:83:@6458.4]
  wire [10:0] _T_59002; // @[Modules.scala 68:83:@6459.4]
  wire [10:0] buffer_2_637; // @[Modules.scala 68:83:@6460.4]
  wire [11:0] _T_59007; // @[Modules.scala 68:83:@6466.4]
  wire [10:0] _T_59008; // @[Modules.scala 68:83:@6467.4]
  wire [10:0] buffer_2_639; // @[Modules.scala 68:83:@6468.4]
  wire [11:0] _T_59010; // @[Modules.scala 68:83:@6470.4]
  wire [10:0] _T_59011; // @[Modules.scala 68:83:@6471.4]
  wire [10:0] buffer_2_640; // @[Modules.scala 68:83:@6472.4]
  wire [11:0] _T_59013; // @[Modules.scala 68:83:@6474.4]
  wire [10:0] _T_59014; // @[Modules.scala 68:83:@6475.4]
  wire [10:0] buffer_2_641; // @[Modules.scala 68:83:@6476.4]
  wire [11:0] _T_59016; // @[Modules.scala 68:83:@6478.4]
  wire [10:0] _T_59017; // @[Modules.scala 68:83:@6479.4]
  wire [10:0] buffer_2_642; // @[Modules.scala 68:83:@6480.4]
  wire [11:0] _T_59019; // @[Modules.scala 68:83:@6482.4]
  wire [10:0] _T_59020; // @[Modules.scala 68:83:@6483.4]
  wire [10:0] buffer_2_643; // @[Modules.scala 68:83:@6484.4]
  wire [11:0] _T_59022; // @[Modules.scala 68:83:@6486.4]
  wire [10:0] _T_59023; // @[Modules.scala 68:83:@6487.4]
  wire [10:0] buffer_2_644; // @[Modules.scala 68:83:@6488.4]
  wire [11:0] _T_59025; // @[Modules.scala 68:83:@6490.4]
  wire [10:0] _T_59026; // @[Modules.scala 68:83:@6491.4]
  wire [10:0] buffer_2_645; // @[Modules.scala 68:83:@6492.4]
  wire [11:0] _T_59028; // @[Modules.scala 68:83:@6494.4]
  wire [10:0] _T_59029; // @[Modules.scala 68:83:@6495.4]
  wire [10:0] buffer_2_646; // @[Modules.scala 68:83:@6496.4]
  wire [11:0] _T_59031; // @[Modules.scala 68:83:@6498.4]
  wire [10:0] _T_59032; // @[Modules.scala 68:83:@6499.4]
  wire [10:0] buffer_2_647; // @[Modules.scala 68:83:@6500.4]
  wire [11:0] _T_59034; // @[Modules.scala 68:83:@6502.4]
  wire [10:0] _T_59035; // @[Modules.scala 68:83:@6503.4]
  wire [10:0] buffer_2_648; // @[Modules.scala 68:83:@6504.4]
  wire [11:0] _T_59037; // @[Modules.scala 68:83:@6506.4]
  wire [10:0] _T_59038; // @[Modules.scala 68:83:@6507.4]
  wire [10:0] buffer_2_649; // @[Modules.scala 68:83:@6508.4]
  wire [11:0] _T_59040; // @[Modules.scala 68:83:@6510.4]
  wire [10:0] _T_59041; // @[Modules.scala 68:83:@6511.4]
  wire [10:0] buffer_2_650; // @[Modules.scala 68:83:@6512.4]
  wire [11:0] _T_59046; // @[Modules.scala 68:83:@6518.4]
  wire [10:0] _T_59047; // @[Modules.scala 68:83:@6519.4]
  wire [10:0] buffer_2_652; // @[Modules.scala 68:83:@6520.4]
  wire [11:0] _T_59049; // @[Modules.scala 68:83:@6522.4]
  wire [10:0] _T_59050; // @[Modules.scala 68:83:@6523.4]
  wire [10:0] buffer_2_653; // @[Modules.scala 68:83:@6524.4]
  wire [11:0] _T_59058; // @[Modules.scala 68:83:@6534.4]
  wire [10:0] _T_59059; // @[Modules.scala 68:83:@6535.4]
  wire [10:0] buffer_2_656; // @[Modules.scala 68:83:@6536.4]
  wire [11:0] _T_59061; // @[Modules.scala 68:83:@6538.4]
  wire [10:0] _T_59062; // @[Modules.scala 68:83:@6539.4]
  wire [10:0] buffer_2_657; // @[Modules.scala 68:83:@6540.4]
  wire [11:0] _T_59064; // @[Modules.scala 68:83:@6542.4]
  wire [10:0] _T_59065; // @[Modules.scala 68:83:@6543.4]
  wire [10:0] buffer_2_658; // @[Modules.scala 68:83:@6544.4]
  wire [11:0] _T_59067; // @[Modules.scala 68:83:@6546.4]
  wire [10:0] _T_59068; // @[Modules.scala 68:83:@6547.4]
  wire [10:0] buffer_2_659; // @[Modules.scala 68:83:@6548.4]
  wire [11:0] _T_59070; // @[Modules.scala 68:83:@6550.4]
  wire [10:0] _T_59071; // @[Modules.scala 68:83:@6551.4]
  wire [10:0] buffer_2_660; // @[Modules.scala 68:83:@6552.4]
  wire [11:0] _T_59073; // @[Modules.scala 68:83:@6554.4]
  wire [10:0] _T_59074; // @[Modules.scala 68:83:@6555.4]
  wire [10:0] buffer_2_661; // @[Modules.scala 68:83:@6556.4]
  wire [11:0] _T_59076; // @[Modules.scala 68:83:@6558.4]
  wire [10:0] _T_59077; // @[Modules.scala 68:83:@6559.4]
  wire [10:0] buffer_2_662; // @[Modules.scala 68:83:@6560.4]
  wire [11:0] _T_59079; // @[Modules.scala 68:83:@6562.4]
  wire [10:0] _T_59080; // @[Modules.scala 68:83:@6563.4]
  wire [10:0] buffer_2_663; // @[Modules.scala 68:83:@6564.4]
  wire [11:0] _T_59082; // @[Modules.scala 68:83:@6566.4]
  wire [10:0] _T_59083; // @[Modules.scala 68:83:@6567.4]
  wire [10:0] buffer_2_664; // @[Modules.scala 68:83:@6568.4]
  wire [11:0] _T_59085; // @[Modules.scala 68:83:@6570.4]
  wire [10:0] _T_59086; // @[Modules.scala 68:83:@6571.4]
  wire [10:0] buffer_2_665; // @[Modules.scala 68:83:@6572.4]
  wire [11:0] _T_59088; // @[Modules.scala 68:83:@6574.4]
  wire [10:0] _T_59089; // @[Modules.scala 68:83:@6575.4]
  wire [10:0] buffer_2_666; // @[Modules.scala 68:83:@6576.4]
  wire [11:0] _T_59091; // @[Modules.scala 68:83:@6578.4]
  wire [10:0] _T_59092; // @[Modules.scala 68:83:@6579.4]
  wire [10:0] buffer_2_667; // @[Modules.scala 68:83:@6580.4]
  wire [11:0] _T_59094; // @[Modules.scala 68:83:@6582.4]
  wire [10:0] _T_59095; // @[Modules.scala 68:83:@6583.4]
  wire [10:0] buffer_2_668; // @[Modules.scala 68:83:@6584.4]
  wire [11:0] _T_59097; // @[Modules.scala 68:83:@6586.4]
  wire [10:0] _T_59098; // @[Modules.scala 68:83:@6587.4]
  wire [10:0] buffer_2_669; // @[Modules.scala 68:83:@6588.4]
  wire [11:0] _T_59100; // @[Modules.scala 68:83:@6590.4]
  wire [10:0] _T_59101; // @[Modules.scala 68:83:@6591.4]
  wire [10:0] buffer_2_670; // @[Modules.scala 68:83:@6592.4]
  wire [11:0] _T_59103; // @[Modules.scala 68:83:@6594.4]
  wire [10:0] _T_59104; // @[Modules.scala 68:83:@6595.4]
  wire [10:0] buffer_2_671; // @[Modules.scala 68:83:@6596.4]
  wire [11:0] _T_59106; // @[Modules.scala 68:83:@6598.4]
  wire [10:0] _T_59107; // @[Modules.scala 68:83:@6599.4]
  wire [10:0] buffer_2_672; // @[Modules.scala 68:83:@6600.4]
  wire [11:0] _T_59109; // @[Modules.scala 68:83:@6602.4]
  wire [10:0] _T_59110; // @[Modules.scala 68:83:@6603.4]
  wire [10:0] buffer_2_673; // @[Modules.scala 68:83:@6604.4]
  wire [11:0] _T_59112; // @[Modules.scala 68:83:@6606.4]
  wire [10:0] _T_59113; // @[Modules.scala 68:83:@6607.4]
  wire [10:0] buffer_2_674; // @[Modules.scala 68:83:@6608.4]
  wire [11:0] _T_59115; // @[Modules.scala 68:83:@6610.4]
  wire [10:0] _T_59116; // @[Modules.scala 68:83:@6611.4]
  wire [10:0] buffer_2_675; // @[Modules.scala 68:83:@6612.4]
  wire [11:0] _T_59127; // @[Modules.scala 68:83:@6626.4]
  wire [10:0] _T_59128; // @[Modules.scala 68:83:@6627.4]
  wire [10:0] buffer_2_679; // @[Modules.scala 68:83:@6628.4]
  wire [11:0] _T_59133; // @[Modules.scala 68:83:@6634.4]
  wire [10:0] _T_59134; // @[Modules.scala 68:83:@6635.4]
  wire [10:0] buffer_2_681; // @[Modules.scala 68:83:@6636.4]
  wire [11:0] _T_59136; // @[Modules.scala 68:83:@6638.4]
  wire [10:0] _T_59137; // @[Modules.scala 68:83:@6639.4]
  wire [10:0] buffer_2_682; // @[Modules.scala 68:83:@6640.4]
  wire [11:0] _T_59145; // @[Modules.scala 68:83:@6650.4]
  wire [10:0] _T_59146; // @[Modules.scala 68:83:@6651.4]
  wire [10:0] buffer_2_685; // @[Modules.scala 68:83:@6652.4]
  wire [11:0] _T_59148; // @[Modules.scala 71:109:@6654.4]
  wire [10:0] _T_59149; // @[Modules.scala 71:109:@6655.4]
  wire [10:0] buffer_2_686; // @[Modules.scala 71:109:@6656.4]
  wire [11:0] _T_59151; // @[Modules.scala 71:109:@6658.4]
  wire [10:0] _T_59152; // @[Modules.scala 71:109:@6659.4]
  wire [10:0] buffer_2_687; // @[Modules.scala 71:109:@6660.4]
  wire [11:0] _T_59154; // @[Modules.scala 71:109:@6662.4]
  wire [10:0] _T_59155; // @[Modules.scala 71:109:@6663.4]
  wire [10:0] buffer_2_688; // @[Modules.scala 71:109:@6664.4]
  wire [11:0] _T_59157; // @[Modules.scala 71:109:@6666.4]
  wire [10:0] _T_59158; // @[Modules.scala 71:109:@6667.4]
  wire [10:0] buffer_2_689; // @[Modules.scala 71:109:@6668.4]
  wire [11:0] _T_59160; // @[Modules.scala 71:109:@6670.4]
  wire [10:0] _T_59161; // @[Modules.scala 71:109:@6671.4]
  wire [10:0] buffer_2_690; // @[Modules.scala 71:109:@6672.4]
  wire [11:0] _T_59163; // @[Modules.scala 71:109:@6674.4]
  wire [10:0] _T_59164; // @[Modules.scala 71:109:@6675.4]
  wire [10:0] buffer_2_691; // @[Modules.scala 71:109:@6676.4]
  wire [11:0] _T_59166; // @[Modules.scala 71:109:@6678.4]
  wire [10:0] _T_59167; // @[Modules.scala 71:109:@6679.4]
  wire [10:0] buffer_2_692; // @[Modules.scala 71:109:@6680.4]
  wire [11:0] _T_59169; // @[Modules.scala 71:109:@6682.4]
  wire [10:0] _T_59170; // @[Modules.scala 71:109:@6683.4]
  wire [10:0] buffer_2_693; // @[Modules.scala 71:109:@6684.4]
  wire [11:0] _T_59172; // @[Modules.scala 71:109:@6686.4]
  wire [10:0] _T_59173; // @[Modules.scala 71:109:@6687.4]
  wire [10:0] buffer_2_694; // @[Modules.scala 71:109:@6688.4]
  wire [11:0] _T_59175; // @[Modules.scala 71:109:@6690.4]
  wire [10:0] _T_59176; // @[Modules.scala 71:109:@6691.4]
  wire [10:0] buffer_2_695; // @[Modules.scala 71:109:@6692.4]
  wire [11:0] _T_59178; // @[Modules.scala 71:109:@6694.4]
  wire [10:0] _T_59179; // @[Modules.scala 71:109:@6695.4]
  wire [10:0] buffer_2_696; // @[Modules.scala 71:109:@6696.4]
  wire [11:0] _T_59181; // @[Modules.scala 71:109:@6698.4]
  wire [10:0] _T_59182; // @[Modules.scala 71:109:@6699.4]
  wire [10:0] buffer_2_697; // @[Modules.scala 71:109:@6700.4]
  wire [11:0] _T_59184; // @[Modules.scala 71:109:@6702.4]
  wire [10:0] _T_59185; // @[Modules.scala 71:109:@6703.4]
  wire [10:0] buffer_2_698; // @[Modules.scala 71:109:@6704.4]
  wire [11:0] _T_59187; // @[Modules.scala 71:109:@6706.4]
  wire [10:0] _T_59188; // @[Modules.scala 71:109:@6707.4]
  wire [10:0] buffer_2_699; // @[Modules.scala 71:109:@6708.4]
  wire [11:0] _T_59190; // @[Modules.scala 71:109:@6710.4]
  wire [10:0] _T_59191; // @[Modules.scala 71:109:@6711.4]
  wire [10:0] buffer_2_700; // @[Modules.scala 71:109:@6712.4]
  wire [11:0] _T_59193; // @[Modules.scala 71:109:@6714.4]
  wire [10:0] _T_59194; // @[Modules.scala 71:109:@6715.4]
  wire [10:0] buffer_2_701; // @[Modules.scala 71:109:@6716.4]
  wire [11:0] _T_59196; // @[Modules.scala 71:109:@6718.4]
  wire [10:0] _T_59197; // @[Modules.scala 71:109:@6719.4]
  wire [10:0] buffer_2_702; // @[Modules.scala 71:109:@6720.4]
  wire [11:0] _T_59199; // @[Modules.scala 71:109:@6722.4]
  wire [10:0] _T_59200; // @[Modules.scala 71:109:@6723.4]
  wire [10:0] buffer_2_703; // @[Modules.scala 71:109:@6724.4]
  wire [11:0] _T_59202; // @[Modules.scala 71:109:@6726.4]
  wire [10:0] _T_59203; // @[Modules.scala 71:109:@6727.4]
  wire [10:0] buffer_2_704; // @[Modules.scala 71:109:@6728.4]
  wire [11:0] _T_59205; // @[Modules.scala 71:109:@6730.4]
  wire [10:0] _T_59206; // @[Modules.scala 71:109:@6731.4]
  wire [10:0] buffer_2_705; // @[Modules.scala 71:109:@6732.4]
  wire [11:0] _T_59208; // @[Modules.scala 71:109:@6734.4]
  wire [10:0] _T_59209; // @[Modules.scala 71:109:@6735.4]
  wire [10:0] buffer_2_706; // @[Modules.scala 71:109:@6736.4]
  wire [11:0] _T_59214; // @[Modules.scala 71:109:@6742.4]
  wire [10:0] _T_59215; // @[Modules.scala 71:109:@6743.4]
  wire [10:0] buffer_2_708; // @[Modules.scala 71:109:@6744.4]
  wire [11:0] _T_59217; // @[Modules.scala 71:109:@6746.4]
  wire [10:0] _T_59218; // @[Modules.scala 71:109:@6747.4]
  wire [10:0] buffer_2_709; // @[Modules.scala 71:109:@6748.4]
  wire [11:0] _T_59220; // @[Modules.scala 71:109:@6750.4]
  wire [10:0] _T_59221; // @[Modules.scala 71:109:@6751.4]
  wire [10:0] buffer_2_710; // @[Modules.scala 71:109:@6752.4]
  wire [11:0] _T_59223; // @[Modules.scala 71:109:@6754.4]
  wire [10:0] _T_59224; // @[Modules.scala 71:109:@6755.4]
  wire [10:0] buffer_2_711; // @[Modules.scala 71:109:@6756.4]
  wire [11:0] _T_59226; // @[Modules.scala 71:109:@6758.4]
  wire [10:0] _T_59227; // @[Modules.scala 71:109:@6759.4]
  wire [10:0] buffer_2_712; // @[Modules.scala 71:109:@6760.4]
  wire [11:0] _T_59229; // @[Modules.scala 71:109:@6762.4]
  wire [10:0] _T_59230; // @[Modules.scala 71:109:@6763.4]
  wire [10:0] buffer_2_713; // @[Modules.scala 71:109:@6764.4]
  wire [11:0] _T_59232; // @[Modules.scala 71:109:@6766.4]
  wire [10:0] _T_59233; // @[Modules.scala 71:109:@6767.4]
  wire [10:0] buffer_2_714; // @[Modules.scala 71:109:@6768.4]
  wire [11:0] _T_59235; // @[Modules.scala 71:109:@6770.4]
  wire [10:0] _T_59236; // @[Modules.scala 71:109:@6771.4]
  wire [10:0] buffer_2_715; // @[Modules.scala 71:109:@6772.4]
  wire [11:0] _T_59238; // @[Modules.scala 71:109:@6774.4]
  wire [10:0] _T_59239; // @[Modules.scala 71:109:@6775.4]
  wire [10:0] buffer_2_716; // @[Modules.scala 71:109:@6776.4]
  wire [11:0] _T_59241; // @[Modules.scala 71:109:@6778.4]
  wire [10:0] _T_59242; // @[Modules.scala 71:109:@6779.4]
  wire [10:0] buffer_2_717; // @[Modules.scala 71:109:@6780.4]
  wire [11:0] _T_59244; // @[Modules.scala 71:109:@6782.4]
  wire [10:0] _T_59245; // @[Modules.scala 71:109:@6783.4]
  wire [10:0] buffer_2_718; // @[Modules.scala 71:109:@6784.4]
  wire [11:0] _T_59247; // @[Modules.scala 71:109:@6786.4]
  wire [10:0] _T_59248; // @[Modules.scala 71:109:@6787.4]
  wire [10:0] buffer_2_719; // @[Modules.scala 71:109:@6788.4]
  wire [11:0] _T_59250; // @[Modules.scala 71:109:@6790.4]
  wire [10:0] _T_59251; // @[Modules.scala 71:109:@6791.4]
  wire [10:0] buffer_2_720; // @[Modules.scala 71:109:@6792.4]
  wire [11:0] _T_59253; // @[Modules.scala 71:109:@6794.4]
  wire [10:0] _T_59254; // @[Modules.scala 71:109:@6795.4]
  wire [10:0] buffer_2_721; // @[Modules.scala 71:109:@6796.4]
  wire [11:0] _T_59256; // @[Modules.scala 71:109:@6798.4]
  wire [10:0] _T_59257; // @[Modules.scala 71:109:@6799.4]
  wire [10:0] buffer_2_722; // @[Modules.scala 71:109:@6800.4]
  wire [11:0] _T_59259; // @[Modules.scala 71:109:@6802.4]
  wire [10:0] _T_59260; // @[Modules.scala 71:109:@6803.4]
  wire [10:0] buffer_2_723; // @[Modules.scala 71:109:@6804.4]
  wire [11:0] _T_59262; // @[Modules.scala 71:109:@6806.4]
  wire [10:0] _T_59263; // @[Modules.scala 71:109:@6807.4]
  wire [10:0] buffer_2_724; // @[Modules.scala 71:109:@6808.4]
  wire [11:0] _T_59265; // @[Modules.scala 71:109:@6810.4]
  wire [10:0] _T_59266; // @[Modules.scala 71:109:@6811.4]
  wire [10:0] buffer_2_725; // @[Modules.scala 71:109:@6812.4]
  wire [11:0] _T_59268; // @[Modules.scala 71:109:@6814.4]
  wire [10:0] _T_59269; // @[Modules.scala 71:109:@6815.4]
  wire [10:0] buffer_2_726; // @[Modules.scala 71:109:@6816.4]
  wire [11:0] _T_59271; // @[Modules.scala 71:109:@6818.4]
  wire [10:0] _T_59272; // @[Modules.scala 71:109:@6819.4]
  wire [10:0] buffer_2_727; // @[Modules.scala 71:109:@6820.4]
  wire [11:0] _T_59274; // @[Modules.scala 71:109:@6822.4]
  wire [10:0] _T_59275; // @[Modules.scala 71:109:@6823.4]
  wire [10:0] buffer_2_728; // @[Modules.scala 71:109:@6824.4]
  wire [11:0] _T_59277; // @[Modules.scala 71:109:@6826.4]
  wire [10:0] _T_59278; // @[Modules.scala 71:109:@6827.4]
  wire [10:0] buffer_2_729; // @[Modules.scala 71:109:@6828.4]
  wire [11:0] _T_59283; // @[Modules.scala 71:109:@6834.4]
  wire [10:0] _T_59284; // @[Modules.scala 71:109:@6835.4]
  wire [10:0] buffer_2_731; // @[Modules.scala 71:109:@6836.4]
  wire [11:0] _T_59286; // @[Modules.scala 71:109:@6838.4]
  wire [10:0] _T_59287; // @[Modules.scala 71:109:@6839.4]
  wire [10:0] buffer_2_732; // @[Modules.scala 71:109:@6840.4]
  wire [11:0] _T_59289; // @[Modules.scala 71:109:@6842.4]
  wire [10:0] _T_59290; // @[Modules.scala 71:109:@6843.4]
  wire [10:0] buffer_2_733; // @[Modules.scala 71:109:@6844.4]
  wire [11:0] _T_59292; // @[Modules.scala 71:109:@6846.4]
  wire [10:0] _T_59293; // @[Modules.scala 71:109:@6847.4]
  wire [10:0] buffer_2_734; // @[Modules.scala 71:109:@6848.4]
  wire [11:0] _T_59295; // @[Modules.scala 78:156:@6851.4]
  wire [10:0] _T_59296; // @[Modules.scala 78:156:@6852.4]
  wire [10:0] buffer_2_736; // @[Modules.scala 78:156:@6853.4]
  wire [11:0] _T_59298; // @[Modules.scala 78:156:@6855.4]
  wire [10:0] _T_59299; // @[Modules.scala 78:156:@6856.4]
  wire [10:0] buffer_2_737; // @[Modules.scala 78:156:@6857.4]
  wire [11:0] _T_59301; // @[Modules.scala 78:156:@6859.4]
  wire [10:0] _T_59302; // @[Modules.scala 78:156:@6860.4]
  wire [10:0] buffer_2_738; // @[Modules.scala 78:156:@6861.4]
  wire [11:0] _T_59304; // @[Modules.scala 78:156:@6863.4]
  wire [10:0] _T_59305; // @[Modules.scala 78:156:@6864.4]
  wire [10:0] buffer_2_739; // @[Modules.scala 78:156:@6865.4]
  wire [11:0] _T_59307; // @[Modules.scala 78:156:@6867.4]
  wire [10:0] _T_59308; // @[Modules.scala 78:156:@6868.4]
  wire [10:0] buffer_2_740; // @[Modules.scala 78:156:@6869.4]
  wire [11:0] _T_59310; // @[Modules.scala 78:156:@6871.4]
  wire [10:0] _T_59311; // @[Modules.scala 78:156:@6872.4]
  wire [10:0] buffer_2_741; // @[Modules.scala 78:156:@6873.4]
  wire [11:0] _T_59313; // @[Modules.scala 78:156:@6875.4]
  wire [10:0] _T_59314; // @[Modules.scala 78:156:@6876.4]
  wire [10:0] buffer_2_742; // @[Modules.scala 78:156:@6877.4]
  wire [11:0] _T_59316; // @[Modules.scala 78:156:@6879.4]
  wire [10:0] _T_59317; // @[Modules.scala 78:156:@6880.4]
  wire [10:0] buffer_2_743; // @[Modules.scala 78:156:@6881.4]
  wire [11:0] _T_59319; // @[Modules.scala 78:156:@6883.4]
  wire [10:0] _T_59320; // @[Modules.scala 78:156:@6884.4]
  wire [10:0] buffer_2_744; // @[Modules.scala 78:156:@6885.4]
  wire [11:0] _T_59322; // @[Modules.scala 78:156:@6887.4]
  wire [10:0] _T_59323; // @[Modules.scala 78:156:@6888.4]
  wire [10:0] buffer_2_745; // @[Modules.scala 78:156:@6889.4]
  wire [11:0] _T_59325; // @[Modules.scala 78:156:@6891.4]
  wire [10:0] _T_59326; // @[Modules.scala 78:156:@6892.4]
  wire [10:0] buffer_2_746; // @[Modules.scala 78:156:@6893.4]
  wire [11:0] _T_59328; // @[Modules.scala 78:156:@6895.4]
  wire [10:0] _T_59329; // @[Modules.scala 78:156:@6896.4]
  wire [10:0] buffer_2_747; // @[Modules.scala 78:156:@6897.4]
  wire [11:0] _T_59331; // @[Modules.scala 78:156:@6899.4]
  wire [10:0] _T_59332; // @[Modules.scala 78:156:@6900.4]
  wire [10:0] buffer_2_748; // @[Modules.scala 78:156:@6901.4]
  wire [11:0] _T_59334; // @[Modules.scala 78:156:@6903.4]
  wire [10:0] _T_59335; // @[Modules.scala 78:156:@6904.4]
  wire [10:0] buffer_2_749; // @[Modules.scala 78:156:@6905.4]
  wire [11:0] _T_59337; // @[Modules.scala 78:156:@6907.4]
  wire [10:0] _T_59338; // @[Modules.scala 78:156:@6908.4]
  wire [10:0] buffer_2_750; // @[Modules.scala 78:156:@6909.4]
  wire [11:0] _T_59340; // @[Modules.scala 78:156:@6911.4]
  wire [10:0] _T_59341; // @[Modules.scala 78:156:@6912.4]
  wire [10:0] buffer_2_751; // @[Modules.scala 78:156:@6913.4]
  wire [11:0] _T_59343; // @[Modules.scala 78:156:@6915.4]
  wire [10:0] _T_59344; // @[Modules.scala 78:156:@6916.4]
  wire [10:0] buffer_2_752; // @[Modules.scala 78:156:@6917.4]
  wire [11:0] _T_59346; // @[Modules.scala 78:156:@6919.4]
  wire [10:0] _T_59347; // @[Modules.scala 78:156:@6920.4]
  wire [10:0] buffer_2_753; // @[Modules.scala 78:156:@6921.4]
  wire [11:0] _T_59349; // @[Modules.scala 78:156:@6923.4]
  wire [10:0] _T_59350; // @[Modules.scala 78:156:@6924.4]
  wire [10:0] buffer_2_754; // @[Modules.scala 78:156:@6925.4]
  wire [11:0] _T_59352; // @[Modules.scala 78:156:@6927.4]
  wire [10:0] _T_59353; // @[Modules.scala 78:156:@6928.4]
  wire [10:0] buffer_2_755; // @[Modules.scala 78:156:@6929.4]
  wire [11:0] _T_59355; // @[Modules.scala 78:156:@6931.4]
  wire [10:0] _T_59356; // @[Modules.scala 78:156:@6932.4]
  wire [10:0] buffer_2_756; // @[Modules.scala 78:156:@6933.4]
  wire [11:0] _T_59358; // @[Modules.scala 78:156:@6935.4]
  wire [10:0] _T_59359; // @[Modules.scala 78:156:@6936.4]
  wire [10:0] buffer_2_757; // @[Modules.scala 78:156:@6937.4]
  wire [11:0] _T_59361; // @[Modules.scala 78:156:@6939.4]
  wire [10:0] _T_59362; // @[Modules.scala 78:156:@6940.4]
  wire [10:0] buffer_2_758; // @[Modules.scala 78:156:@6941.4]
  wire [11:0] _T_59364; // @[Modules.scala 78:156:@6943.4]
  wire [10:0] _T_59365; // @[Modules.scala 78:156:@6944.4]
  wire [10:0] buffer_2_759; // @[Modules.scala 78:156:@6945.4]
  wire [11:0] _T_59367; // @[Modules.scala 78:156:@6947.4]
  wire [10:0] _T_59368; // @[Modules.scala 78:156:@6948.4]
  wire [10:0] buffer_2_760; // @[Modules.scala 78:156:@6949.4]
  wire [11:0] _T_59370; // @[Modules.scala 78:156:@6951.4]
  wire [10:0] _T_59371; // @[Modules.scala 78:156:@6952.4]
  wire [10:0] buffer_2_761; // @[Modules.scala 78:156:@6953.4]
  wire [11:0] _T_59373; // @[Modules.scala 78:156:@6955.4]
  wire [10:0] _T_59374; // @[Modules.scala 78:156:@6956.4]
  wire [10:0] buffer_2_762; // @[Modules.scala 78:156:@6957.4]
  wire [11:0] _T_59376; // @[Modules.scala 78:156:@6959.4]
  wire [10:0] _T_59377; // @[Modules.scala 78:156:@6960.4]
  wire [10:0] buffer_2_763; // @[Modules.scala 78:156:@6961.4]
  wire [11:0] _T_59379; // @[Modules.scala 78:156:@6963.4]
  wire [10:0] _T_59380; // @[Modules.scala 78:156:@6964.4]
  wire [10:0] buffer_2_764; // @[Modules.scala 78:156:@6965.4]
  wire [11:0] _T_59382; // @[Modules.scala 78:156:@6967.4]
  wire [10:0] _T_59383; // @[Modules.scala 78:156:@6968.4]
  wire [10:0] buffer_2_765; // @[Modules.scala 78:156:@6969.4]
  wire [11:0] _T_59385; // @[Modules.scala 78:156:@6971.4]
  wire [10:0] _T_59386; // @[Modules.scala 78:156:@6972.4]
  wire [10:0] buffer_2_766; // @[Modules.scala 78:156:@6973.4]
  wire [11:0] _T_59388; // @[Modules.scala 78:156:@6975.4]
  wire [10:0] _T_59389; // @[Modules.scala 78:156:@6976.4]
  wire [10:0] buffer_2_767; // @[Modules.scala 78:156:@6977.4]
  wire [11:0] _T_59391; // @[Modules.scala 78:156:@6979.4]
  wire [10:0] _T_59392; // @[Modules.scala 78:156:@6980.4]
  wire [10:0] buffer_2_768; // @[Modules.scala 78:156:@6981.4]
  wire [11:0] _T_59394; // @[Modules.scala 78:156:@6983.4]
  wire [10:0] _T_59395; // @[Modules.scala 78:156:@6984.4]
  wire [10:0] buffer_2_769; // @[Modules.scala 78:156:@6985.4]
  wire [11:0] _T_59397; // @[Modules.scala 78:156:@6987.4]
  wire [10:0] _T_59398; // @[Modules.scala 78:156:@6988.4]
  wire [10:0] buffer_2_770; // @[Modules.scala 78:156:@6989.4]
  wire [11:0] _T_59400; // @[Modules.scala 78:156:@6991.4]
  wire [10:0] _T_59401; // @[Modules.scala 78:156:@6992.4]
  wire [10:0] buffer_2_771; // @[Modules.scala 78:156:@6993.4]
  wire [11:0] _T_59403; // @[Modules.scala 78:156:@6995.4]
  wire [10:0] _T_59404; // @[Modules.scala 78:156:@6996.4]
  wire [10:0] buffer_2_772; // @[Modules.scala 78:156:@6997.4]
  wire [11:0] _T_59406; // @[Modules.scala 78:156:@6999.4]
  wire [10:0] _T_59407; // @[Modules.scala 78:156:@7000.4]
  wire [10:0] buffer_2_773; // @[Modules.scala 78:156:@7001.4]
  wire [11:0] _T_59409; // @[Modules.scala 78:156:@7003.4]
  wire [10:0] _T_59410; // @[Modules.scala 78:156:@7004.4]
  wire [10:0] buffer_2_774; // @[Modules.scala 78:156:@7005.4]
  wire [11:0] _T_59412; // @[Modules.scala 78:156:@7007.4]
  wire [10:0] _T_59413; // @[Modules.scala 78:156:@7008.4]
  wire [10:0] buffer_2_775; // @[Modules.scala 78:156:@7009.4]
  wire [11:0] _T_59415; // @[Modules.scala 78:156:@7011.4]
  wire [10:0] _T_59416; // @[Modules.scala 78:156:@7012.4]
  wire [10:0] buffer_2_776; // @[Modules.scala 78:156:@7013.4]
  wire [11:0] _T_59418; // @[Modules.scala 78:156:@7015.4]
  wire [10:0] _T_59419; // @[Modules.scala 78:156:@7016.4]
  wire [10:0] buffer_2_777; // @[Modules.scala 78:156:@7017.4]
  wire [11:0] _T_59421; // @[Modules.scala 78:156:@7019.4]
  wire [10:0] _T_59422; // @[Modules.scala 78:156:@7020.4]
  wire [10:0] buffer_2_778; // @[Modules.scala 78:156:@7021.4]
  wire [11:0] _T_59424; // @[Modules.scala 78:156:@7023.4]
  wire [10:0] _T_59425; // @[Modules.scala 78:156:@7024.4]
  wire [10:0] buffer_2_779; // @[Modules.scala 78:156:@7025.4]
  wire [11:0] _T_59427; // @[Modules.scala 78:156:@7027.4]
  wire [10:0] _T_59428; // @[Modules.scala 78:156:@7028.4]
  wire [10:0] buffer_2_780; // @[Modules.scala 78:156:@7029.4]
  wire [11:0] _T_59430; // @[Modules.scala 78:156:@7031.4]
  wire [10:0] _T_59431; // @[Modules.scala 78:156:@7032.4]
  wire [10:0] buffer_2_781; // @[Modules.scala 78:156:@7033.4]
  wire [11:0] _T_59433; // @[Modules.scala 78:156:@7035.4]
  wire [10:0] _T_59434; // @[Modules.scala 78:156:@7036.4]
  wire [10:0] buffer_2_782; // @[Modules.scala 78:156:@7037.4]
  wire [11:0] _T_59436; // @[Modules.scala 78:156:@7039.4]
  wire [10:0] _T_59437; // @[Modules.scala 78:156:@7040.4]
  wire [10:0] buffer_2_783; // @[Modules.scala 78:156:@7041.4]
  wire [5:0] _T_59453; // @[Modules.scala 37:46:@7069.4]
  wire [4:0] _T_59454; // @[Modules.scala 37:46:@7070.4]
  wire [4:0] _T_59455; // @[Modules.scala 37:46:@7071.4]
  wire [5:0] _T_59456; // @[Modules.scala 37:46:@7073.4]
  wire [4:0] _T_59457; // @[Modules.scala 37:46:@7074.4]
  wire [4:0] _T_59458; // @[Modules.scala 37:46:@7075.4]
  wire [5:0] _T_59506; // @[Modules.scala 37:46:@7143.4]
  wire [4:0] _T_59507; // @[Modules.scala 37:46:@7144.4]
  wire [4:0] _T_59508; // @[Modules.scala 37:46:@7145.4]
  wire [5:0] _T_59513; // @[Modules.scala 37:46:@7152.4]
  wire [4:0] _T_59514; // @[Modules.scala 37:46:@7153.4]
  wire [4:0] _T_59515; // @[Modules.scala 37:46:@7154.4]
  wire [5:0] _T_59516; // @[Modules.scala 37:46:@7156.4]
  wire [4:0] _T_59517; // @[Modules.scala 37:46:@7157.4]
  wire [4:0] _T_59518; // @[Modules.scala 37:46:@7158.4]
  wire [5:0] _T_59519; // @[Modules.scala 37:46:@7160.4]
  wire [4:0] _T_59520; // @[Modules.scala 37:46:@7161.4]
  wire [4:0] _T_59521; // @[Modules.scala 37:46:@7162.4]
  wire [5:0] _T_59522; // @[Modules.scala 37:46:@7164.4]
  wire [4:0] _T_59523; // @[Modules.scala 37:46:@7165.4]
  wire [4:0] _T_59524; // @[Modules.scala 37:46:@7166.4]
  wire [5:0] _T_59544; // @[Modules.scala 37:46:@7197.4]
  wire [4:0] _T_59545; // @[Modules.scala 37:46:@7198.4]
  wire [4:0] _T_59546; // @[Modules.scala 37:46:@7199.4]
  wire [5:0] _T_59547; // @[Modules.scala 37:46:@7202.4]
  wire [4:0] _T_59548; // @[Modules.scala 37:46:@7203.4]
  wire [4:0] _T_59549; // @[Modules.scala 37:46:@7204.4]
  wire [5:0] _T_59550; // @[Modules.scala 37:46:@7207.4]
  wire [4:0] _T_59551; // @[Modules.scala 37:46:@7208.4]
  wire [4:0] _T_59552; // @[Modules.scala 37:46:@7209.4]
  wire [5:0] _T_59568; // @[Modules.scala 37:46:@7232.4]
  wire [4:0] _T_59569; // @[Modules.scala 37:46:@7233.4]
  wire [4:0] _T_59570; // @[Modules.scala 37:46:@7234.4]
  wire [5:0] _T_59577; // @[Modules.scala 37:46:@7244.4]
  wire [4:0] _T_59578; // @[Modules.scala 37:46:@7245.4]
  wire [4:0] _T_59579; // @[Modules.scala 37:46:@7246.4]
  wire [5:0] _T_59580; // @[Modules.scala 37:46:@7248.4]
  wire [4:0] _T_59581; // @[Modules.scala 37:46:@7249.4]
  wire [4:0] _T_59582; // @[Modules.scala 37:46:@7250.4]
  wire [5:0] _T_59590; // @[Modules.scala 37:46:@7266.4]
  wire [4:0] _T_59591; // @[Modules.scala 37:46:@7267.4]
  wire [4:0] _T_59592; // @[Modules.scala 37:46:@7268.4]
  wire [5:0] _T_59593; // @[Modules.scala 37:46:@7270.4]
  wire [4:0] _T_59594; // @[Modules.scala 37:46:@7271.4]
  wire [4:0] _T_59595; // @[Modules.scala 37:46:@7272.4]
  wire [5:0] _T_59599; // @[Modules.scala 37:46:@7279.4]
  wire [4:0] _T_59600; // @[Modules.scala 37:46:@7280.4]
  wire [4:0] _T_59601; // @[Modules.scala 37:46:@7281.4]
  wire [5:0] _T_59602; // @[Modules.scala 37:46:@7283.4]
  wire [4:0] _T_59603; // @[Modules.scala 37:46:@7284.4]
  wire [4:0] _T_59604; // @[Modules.scala 37:46:@7285.4]
  wire [5:0] _T_59605; // @[Modules.scala 37:46:@7288.4]
  wire [4:0] _T_59606; // @[Modules.scala 37:46:@7289.4]
  wire [4:0] _T_59607; // @[Modules.scala 37:46:@7290.4]
  wire [5:0] _T_59620; // @[Modules.scala 37:46:@7310.4]
  wire [4:0] _T_59621; // @[Modules.scala 37:46:@7311.4]
  wire [4:0] _T_59622; // @[Modules.scala 37:46:@7312.4]
  wire [5:0] _T_59623; // @[Modules.scala 37:46:@7314.4]
  wire [4:0] _T_59624; // @[Modules.scala 37:46:@7315.4]
  wire [4:0] _T_59625; // @[Modules.scala 37:46:@7316.4]
  wire [5:0] _T_59626; // @[Modules.scala 37:46:@7320.4]
  wire [4:0] _T_59627; // @[Modules.scala 37:46:@7321.4]
  wire [4:0] _T_59628; // @[Modules.scala 37:46:@7322.4]
  wire [5:0] _T_59629; // @[Modules.scala 37:46:@7324.4]
  wire [4:0] _T_59630; // @[Modules.scala 37:46:@7325.4]
  wire [4:0] _T_59631; // @[Modules.scala 37:46:@7326.4]
  wire [5:0] _T_59632; // @[Modules.scala 37:46:@7328.4]
  wire [4:0] _T_59633; // @[Modules.scala 37:46:@7329.4]
  wire [4:0] _T_59634; // @[Modules.scala 37:46:@7330.4]
  wire [5:0] _T_59638; // @[Modules.scala 37:46:@7336.4]
  wire [4:0] _T_59639; // @[Modules.scala 37:46:@7337.4]
  wire [4:0] _T_59640; // @[Modules.scala 37:46:@7338.4]
  wire [5:0] _T_59641; // @[Modules.scala 37:46:@7341.4]
  wire [4:0] _T_59642; // @[Modules.scala 37:46:@7342.4]
  wire [4:0] _T_59643; // @[Modules.scala 37:46:@7343.4]
  wire [5:0] _T_59650; // @[Modules.scala 37:46:@7353.4]
  wire [4:0] _T_59651; // @[Modules.scala 37:46:@7354.4]
  wire [4:0] _T_59652; // @[Modules.scala 37:46:@7355.4]
  wire [5:0] _T_59653; // @[Modules.scala 37:46:@7357.4]
  wire [4:0] _T_59654; // @[Modules.scala 37:46:@7358.4]
  wire [4:0] _T_59655; // @[Modules.scala 37:46:@7359.4]
  wire [5:0] _T_59656; // @[Modules.scala 37:46:@7361.4]
  wire [4:0] _T_59657; // @[Modules.scala 37:46:@7362.4]
  wire [4:0] _T_59658; // @[Modules.scala 37:46:@7363.4]
  wire [5:0] _T_59660; // @[Modules.scala 37:46:@7368.4]
  wire [4:0] _T_59661; // @[Modules.scala 37:46:@7369.4]
  wire [4:0] _T_59662; // @[Modules.scala 37:46:@7370.4]
  wire [5:0] _T_59666; // @[Modules.scala 37:46:@7376.4]
  wire [4:0] _T_59667; // @[Modules.scala 37:46:@7377.4]
  wire [4:0] _T_59668; // @[Modules.scala 37:46:@7378.4]
  wire [5:0] _T_59669; // @[Modules.scala 37:46:@7380.4]
  wire [4:0] _T_59670; // @[Modules.scala 37:46:@7381.4]
  wire [4:0] _T_59671; // @[Modules.scala 37:46:@7382.4]
  wire [5:0] _T_59672; // @[Modules.scala 37:46:@7384.4]
  wire [4:0] _T_59673; // @[Modules.scala 37:46:@7385.4]
  wire [4:0] _T_59674; // @[Modules.scala 37:46:@7386.4]
  wire [5:0] _T_59675; // @[Modules.scala 37:46:@7388.4]
  wire [4:0] _T_59676; // @[Modules.scala 37:46:@7389.4]
  wire [4:0] _T_59677; // @[Modules.scala 37:46:@7390.4]
  wire [5:0] _T_59684; // @[Modules.scala 37:46:@7400.4]
  wire [4:0] _T_59685; // @[Modules.scala 37:46:@7401.4]
  wire [4:0] _T_59686; // @[Modules.scala 37:46:@7402.4]
  wire [5:0] _T_59687; // @[Modules.scala 37:46:@7404.4]
  wire [4:0] _T_59688; // @[Modules.scala 37:46:@7405.4]
  wire [4:0] _T_59689; // @[Modules.scala 37:46:@7406.4]
  wire [5:0] _T_59694; // @[Modules.scala 37:46:@7414.4]
  wire [4:0] _T_59695; // @[Modules.scala 37:46:@7415.4]
  wire [4:0] _T_59696; // @[Modules.scala 37:46:@7416.4]
  wire [5:0] _T_59704; // @[Modules.scala 37:46:@7430.4]
  wire [4:0] _T_59705; // @[Modules.scala 37:46:@7431.4]
  wire [4:0] _T_59706; // @[Modules.scala 37:46:@7432.4]
  wire [5:0] _T_59738; // @[Modules.scala 37:46:@7473.4]
  wire [4:0] _T_59739; // @[Modules.scala 37:46:@7474.4]
  wire [4:0] _T_59740; // @[Modules.scala 37:46:@7475.4]
  wire [5:0] _T_59751; // @[Modules.scala 37:46:@7493.4]
  wire [4:0] _T_59752; // @[Modules.scala 37:46:@7494.4]
  wire [4:0] _T_59753; // @[Modules.scala 37:46:@7495.4]
  wire [5:0] _T_59757; // @[Modules.scala 37:46:@7502.4]
  wire [4:0] _T_59758; // @[Modules.scala 37:46:@7503.4]
  wire [4:0] _T_59759; // @[Modules.scala 37:46:@7504.4]
  wire [5:0] _T_59769; // @[Modules.scala 37:46:@7518.4]
  wire [4:0] _T_59770; // @[Modules.scala 37:46:@7519.4]
  wire [4:0] _T_59771; // @[Modules.scala 37:46:@7520.4]
  wire [5:0] _T_59772; // @[Modules.scala 37:46:@7522.4]
  wire [4:0] _T_59773; // @[Modules.scala 37:46:@7523.4]
  wire [4:0] _T_59774; // @[Modules.scala 37:46:@7524.4]
  wire [5:0] _T_59778; // @[Modules.scala 37:46:@7531.4]
  wire [4:0] _T_59779; // @[Modules.scala 37:46:@7532.4]
  wire [4:0] _T_59780; // @[Modules.scala 37:46:@7533.4]
  wire [5:0] _T_59798; // @[Modules.scala 37:46:@7556.4]
  wire [4:0] _T_59799; // @[Modules.scala 37:46:@7557.4]
  wire [4:0] _T_59800; // @[Modules.scala 37:46:@7558.4]
  wire [5:0] _T_59801; // @[Modules.scala 37:46:@7560.4]
  wire [4:0] _T_59802; // @[Modules.scala 37:46:@7561.4]
  wire [4:0] _T_59803; // @[Modules.scala 37:46:@7562.4]
  wire [5:0] _T_59808; // @[Modules.scala 37:46:@7569.4]
  wire [4:0] _T_59809; // @[Modules.scala 37:46:@7570.4]
  wire [4:0] _T_59810; // @[Modules.scala 37:46:@7571.4]
  wire [5:0] _T_59824; // @[Modules.scala 37:46:@7591.4]
  wire [4:0] _T_59825; // @[Modules.scala 37:46:@7592.4]
  wire [4:0] _T_59826; // @[Modules.scala 37:46:@7593.4]
  wire [5:0] _T_59827; // @[Modules.scala 37:46:@7595.4]
  wire [4:0] _T_59828; // @[Modules.scala 37:46:@7596.4]
  wire [4:0] _T_59829; // @[Modules.scala 37:46:@7597.4]
  wire [5:0] _T_59833; // @[Modules.scala 37:46:@7604.4]
  wire [4:0] _T_59834; // @[Modules.scala 37:46:@7605.4]
  wire [4:0] _T_59835; // @[Modules.scala 37:46:@7606.4]
  wire [5:0] _T_59855; // @[Modules.scala 37:46:@7633.4]
  wire [4:0] _T_59856; // @[Modules.scala 37:46:@7634.4]
  wire [4:0] _T_59857; // @[Modules.scala 37:46:@7635.4]
  wire [5:0] _T_59877; // @[Modules.scala 37:46:@7663.4]
  wire [4:0] _T_59878; // @[Modules.scala 37:46:@7664.4]
  wire [4:0] _T_59879; // @[Modules.scala 37:46:@7665.4]
  wire [5:0] _T_59880; // @[Modules.scala 37:46:@7667.4]
  wire [4:0] _T_59881; // @[Modules.scala 37:46:@7668.4]
  wire [4:0] _T_59882; // @[Modules.scala 37:46:@7669.4]
  wire [5:0] _T_59889; // @[Modules.scala 37:46:@7681.4]
  wire [4:0] _T_59890; // @[Modules.scala 37:46:@7682.4]
  wire [4:0] _T_59891; // @[Modules.scala 37:46:@7683.4]
  wire [5:0] _T_59898; // @[Modules.scala 37:46:@7698.4]
  wire [4:0] _T_59899; // @[Modules.scala 37:46:@7699.4]
  wire [4:0] _T_59900; // @[Modules.scala 37:46:@7700.4]
  wire [5:0] _T_59904; // @[Modules.scala 37:46:@7706.4]
  wire [4:0] _T_59905; // @[Modules.scala 37:46:@7707.4]
  wire [4:0] _T_59906; // @[Modules.scala 37:46:@7708.4]
  wire [5:0] _T_59914; // @[Modules.scala 37:46:@7719.4]
  wire [4:0] _T_59915; // @[Modules.scala 37:46:@7720.4]
  wire [4:0] _T_59916; // @[Modules.scala 37:46:@7721.4]
  wire [5:0] _T_59922; // @[Modules.scala 37:46:@7733.4]
  wire [4:0] _T_59923; // @[Modules.scala 37:46:@7734.4]
  wire [4:0] _T_59924; // @[Modules.scala 37:46:@7735.4]
  wire [5:0] _T_59932; // @[Modules.scala 37:46:@7747.4]
  wire [4:0] _T_59933; // @[Modules.scala 37:46:@7748.4]
  wire [4:0] _T_59934; // @[Modules.scala 37:46:@7749.4]
  wire [5:0] _T_59945; // @[Modules.scala 37:46:@7768.4]
  wire [4:0] _T_59946; // @[Modules.scala 37:46:@7769.4]
  wire [4:0] _T_59947; // @[Modules.scala 37:46:@7770.4]
  wire [5:0] _T_59979; // @[Modules.scala 37:46:@7822.4]
  wire [4:0] _T_59980; // @[Modules.scala 37:46:@7823.4]
  wire [4:0] _T_59981; // @[Modules.scala 37:46:@7824.4]
  wire [5:0] _T_59987; // @[Modules.scala 37:46:@7831.4]
  wire [4:0] _T_59988; // @[Modules.scala 37:46:@7832.4]
  wire [4:0] _T_59989; // @[Modules.scala 37:46:@7833.4]
  wire [5:0] _T_59999; // @[Modules.scala 37:46:@7849.4]
  wire [4:0] _T_60000; // @[Modules.scala 37:46:@7850.4]
  wire [4:0] _T_60001; // @[Modules.scala 37:46:@7851.4]
  wire [5:0] _T_60020; // @[Modules.scala 37:46:@7880.4]
  wire [4:0] _T_60021; // @[Modules.scala 37:46:@7881.4]
  wire [4:0] _T_60022; // @[Modules.scala 37:46:@7882.4]
  wire [5:0] _T_60023; // @[Modules.scala 37:46:@7884.4]
  wire [4:0] _T_60024; // @[Modules.scala 37:46:@7885.4]
  wire [4:0] _T_60025; // @[Modules.scala 37:46:@7886.4]
  wire [5:0] _T_60026; // @[Modules.scala 37:46:@7888.4]
  wire [4:0] _T_60027; // @[Modules.scala 37:46:@7889.4]
  wire [4:0] _T_60028; // @[Modules.scala 37:46:@7890.4]
  wire [5:0] _T_60029; // @[Modules.scala 37:46:@7893.4]
  wire [4:0] _T_60030; // @[Modules.scala 37:46:@7894.4]
  wire [4:0] _T_60031; // @[Modules.scala 37:46:@7895.4]
  wire [5:0] _T_60032; // @[Modules.scala 37:46:@7897.4]
  wire [4:0] _T_60033; // @[Modules.scala 37:46:@7898.4]
  wire [4:0] _T_60034; // @[Modules.scala 37:46:@7899.4]
  wire [5:0] _T_60036; // @[Modules.scala 37:46:@7905.4]
  wire [4:0] _T_60037; // @[Modules.scala 37:46:@7906.4]
  wire [4:0] _T_60038; // @[Modules.scala 37:46:@7907.4]
  wire [5:0] _T_60046; // @[Modules.scala 37:46:@7918.4]
  wire [4:0] _T_60047; // @[Modules.scala 37:46:@7919.4]
  wire [4:0] _T_60048; // @[Modules.scala 37:46:@7920.4]
  wire [5:0] _T_60052; // @[Modules.scala 37:46:@7926.4]
  wire [4:0] _T_60053; // @[Modules.scala 37:46:@7927.4]
  wire [4:0] _T_60054; // @[Modules.scala 37:46:@7928.4]
  wire [5:0] _T_60055; // @[Modules.scala 37:46:@7930.4]
  wire [4:0] _T_60056; // @[Modules.scala 37:46:@7931.4]
  wire [4:0] _T_60057; // @[Modules.scala 37:46:@7932.4]
  wire [5:0] _T_60058; // @[Modules.scala 37:46:@7934.4]
  wire [4:0] _T_60059; // @[Modules.scala 37:46:@7935.4]
  wire [4:0] _T_60060; // @[Modules.scala 37:46:@7936.4]
  wire [5:0] _T_60061; // @[Modules.scala 37:46:@7938.4]
  wire [4:0] _T_60062; // @[Modules.scala 37:46:@7939.4]
  wire [4:0] _T_60063; // @[Modules.scala 37:46:@7940.4]
  wire [10:0] buffer_3_0; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60068; // @[Modules.scala 65:57:@7949.4]
  wire [10:0] _T_60069; // @[Modules.scala 65:57:@7950.4]
  wire [10:0] buffer_3_392; // @[Modules.scala 65:57:@7951.4]
  wire [10:0] buffer_3_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60074; // @[Modules.scala 65:57:@7957.4]
  wire [10:0] _T_60075; // @[Modules.scala 65:57:@7958.4]
  wire [10:0] buffer_3_394; // @[Modules.scala 65:57:@7959.4]
  wire [11:0] _T_60080; // @[Modules.scala 65:57:@7965.4]
  wire [10:0] _T_60081; // @[Modules.scala 65:57:@7966.4]
  wire [10:0] buffer_3_396; // @[Modules.scala 65:57:@7967.4]
  wire [11:0] _T_60083; // @[Modules.scala 65:57:@7969.4]
  wire [10:0] _T_60084; // @[Modules.scala 65:57:@7970.4]
  wire [10:0] buffer_3_397; // @[Modules.scala 65:57:@7971.4]
  wire [10:0] buffer_3_12; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60086; // @[Modules.scala 65:57:@7973.4]
  wire [10:0] _T_60087; // @[Modules.scala 65:57:@7974.4]
  wire [10:0] buffer_3_398; // @[Modules.scala 65:57:@7975.4]
  wire [10:0] buffer_3_14; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60089; // @[Modules.scala 65:57:@7977.4]
  wire [10:0] _T_60090; // @[Modules.scala 65:57:@7978.4]
  wire [10:0] buffer_3_399; // @[Modules.scala 65:57:@7979.4]
  wire [10:0] buffer_3_16; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60092; // @[Modules.scala 65:57:@7981.4]
  wire [10:0] _T_60093; // @[Modules.scala 65:57:@7982.4]
  wire [10:0] buffer_3_400; // @[Modules.scala 65:57:@7983.4]
  wire [11:0] _T_60101; // @[Modules.scala 65:57:@7993.4]
  wire [10:0] _T_60102; // @[Modules.scala 65:57:@7994.4]
  wire [10:0] buffer_3_403; // @[Modules.scala 65:57:@7995.4]
  wire [11:0] _T_60104; // @[Modules.scala 65:57:@7997.4]
  wire [10:0] _T_60105; // @[Modules.scala 65:57:@7998.4]
  wire [10:0] buffer_3_404; // @[Modules.scala 65:57:@7999.4]
  wire [10:0] buffer_3_26; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60107; // @[Modules.scala 65:57:@8001.4]
  wire [10:0] _T_60108; // @[Modules.scala 65:57:@8002.4]
  wire [10:0] buffer_3_405; // @[Modules.scala 65:57:@8003.4]
  wire [10:0] buffer_3_29; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60110; // @[Modules.scala 65:57:@8005.4]
  wire [10:0] _T_60111; // @[Modules.scala 65:57:@8006.4]
  wire [10:0] buffer_3_406; // @[Modules.scala 65:57:@8007.4]
  wire [10:0] buffer_3_30; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60113; // @[Modules.scala 65:57:@8009.4]
  wire [10:0] _T_60114; // @[Modules.scala 65:57:@8010.4]
  wire [10:0] buffer_3_407; // @[Modules.scala 65:57:@8011.4]
  wire [11:0] _T_60128; // @[Modules.scala 65:57:@8029.4]
  wire [10:0] _T_60129; // @[Modules.scala 65:57:@8030.4]
  wire [10:0] buffer_3_412; // @[Modules.scala 65:57:@8031.4]
  wire [10:0] buffer_3_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60131; // @[Modules.scala 65:57:@8033.4]
  wire [10:0] _T_60132; // @[Modules.scala 65:57:@8034.4]
  wire [10:0] buffer_3_413; // @[Modules.scala 65:57:@8035.4]
  wire [11:0] _T_60137; // @[Modules.scala 65:57:@8041.4]
  wire [10:0] _T_60138; // @[Modules.scala 65:57:@8042.4]
  wire [10:0] buffer_3_415; // @[Modules.scala 65:57:@8043.4]
  wire [10:0] buffer_3_49; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60140; // @[Modules.scala 65:57:@8045.4]
  wire [10:0] _T_60141; // @[Modules.scala 65:57:@8046.4]
  wire [10:0] buffer_3_416; // @[Modules.scala 65:57:@8047.4]
  wire [11:0] _T_60143; // @[Modules.scala 65:57:@8049.4]
  wire [10:0] _T_60144; // @[Modules.scala 65:57:@8050.4]
  wire [10:0] buffer_3_417; // @[Modules.scala 65:57:@8051.4]
  wire [10:0] buffer_3_54; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60149; // @[Modules.scala 65:57:@8057.4]
  wire [10:0] _T_60150; // @[Modules.scala 65:57:@8058.4]
  wire [10:0] buffer_3_419; // @[Modules.scala 65:57:@8059.4]
  wire [10:0] buffer_3_56; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60152; // @[Modules.scala 65:57:@8061.4]
  wire [10:0] _T_60153; // @[Modules.scala 65:57:@8062.4]
  wire [10:0] buffer_3_420; // @[Modules.scala 65:57:@8063.4]
  wire [11:0] _T_60155; // @[Modules.scala 65:57:@8065.4]
  wire [10:0] _T_60156; // @[Modules.scala 65:57:@8066.4]
  wire [10:0] buffer_3_421; // @[Modules.scala 65:57:@8067.4]
  wire [10:0] buffer_3_60; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60158; // @[Modules.scala 65:57:@8069.4]
  wire [10:0] _T_60159; // @[Modules.scala 65:57:@8070.4]
  wire [10:0] buffer_3_422; // @[Modules.scala 65:57:@8071.4]
  wire [10:0] buffer_3_62; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60161; // @[Modules.scala 65:57:@8073.4]
  wire [10:0] _T_60162; // @[Modules.scala 65:57:@8074.4]
  wire [10:0] buffer_3_423; // @[Modules.scala 65:57:@8075.4]
  wire [10:0] buffer_3_67; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60167; // @[Modules.scala 65:57:@8081.4]
  wire [10:0] _T_60168; // @[Modules.scala 65:57:@8082.4]
  wire [10:0] buffer_3_425; // @[Modules.scala 65:57:@8083.4]
  wire [10:0] buffer_3_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60170; // @[Modules.scala 65:57:@8085.4]
  wire [10:0] _T_60171; // @[Modules.scala 65:57:@8086.4]
  wire [10:0] buffer_3_426; // @[Modules.scala 65:57:@8087.4]
  wire [11:0] _T_60173; // @[Modules.scala 65:57:@8089.4]
  wire [10:0] _T_60174; // @[Modules.scala 65:57:@8090.4]
  wire [10:0] buffer_3_427; // @[Modules.scala 65:57:@8091.4]
  wire [10:0] buffer_3_72; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60176; // @[Modules.scala 65:57:@8093.4]
  wire [10:0] _T_60177; // @[Modules.scala 65:57:@8094.4]
  wire [10:0] buffer_3_428; // @[Modules.scala 65:57:@8095.4]
  wire [10:0] buffer_3_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60179; // @[Modules.scala 65:57:@8097.4]
  wire [10:0] _T_60180; // @[Modules.scala 65:57:@8098.4]
  wire [10:0] buffer_3_429; // @[Modules.scala 65:57:@8099.4]
  wire [10:0] buffer_3_76; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_77; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60182; // @[Modules.scala 65:57:@8101.4]
  wire [10:0] _T_60183; // @[Modules.scala 65:57:@8102.4]
  wire [10:0] buffer_3_430; // @[Modules.scala 65:57:@8103.4]
  wire [10:0] buffer_3_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60185; // @[Modules.scala 65:57:@8105.4]
  wire [10:0] _T_60186; // @[Modules.scala 65:57:@8106.4]
  wire [10:0] buffer_3_431; // @[Modules.scala 65:57:@8107.4]
  wire [10:0] buffer_3_86; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60197; // @[Modules.scala 65:57:@8121.4]
  wire [10:0] _T_60198; // @[Modules.scala 65:57:@8122.4]
  wire [10:0] buffer_3_435; // @[Modules.scala 65:57:@8123.4]
  wire [10:0] buffer_3_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60200; // @[Modules.scala 65:57:@8125.4]
  wire [10:0] _T_60201; // @[Modules.scala 65:57:@8126.4]
  wire [10:0] buffer_3_436; // @[Modules.scala 65:57:@8127.4]
  wire [10:0] buffer_3_90; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60203; // @[Modules.scala 65:57:@8129.4]
  wire [10:0] _T_60204; // @[Modules.scala 65:57:@8130.4]
  wire [10:0] buffer_3_437; // @[Modules.scala 65:57:@8131.4]
  wire [10:0] buffer_3_92; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60206; // @[Modules.scala 65:57:@8133.4]
  wire [10:0] _T_60207; // @[Modules.scala 65:57:@8134.4]
  wire [10:0] buffer_3_438; // @[Modules.scala 65:57:@8135.4]
  wire [11:0] _T_60209; // @[Modules.scala 65:57:@8137.4]
  wire [10:0] _T_60210; // @[Modules.scala 65:57:@8138.4]
  wire [10:0] buffer_3_439; // @[Modules.scala 65:57:@8139.4]
  wire [10:0] buffer_3_98; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_99; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60215; // @[Modules.scala 65:57:@8145.4]
  wire [10:0] _T_60216; // @[Modules.scala 65:57:@8146.4]
  wire [10:0] buffer_3_441; // @[Modules.scala 65:57:@8147.4]
  wire [10:0] buffer_3_100; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60218; // @[Modules.scala 65:57:@8149.4]
  wire [10:0] _T_60219; // @[Modules.scala 65:57:@8150.4]
  wire [10:0] buffer_3_442; // @[Modules.scala 65:57:@8151.4]
  wire [10:0] buffer_3_103; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60221; // @[Modules.scala 65:57:@8153.4]
  wire [10:0] _T_60222; // @[Modules.scala 65:57:@8154.4]
  wire [10:0] buffer_3_443; // @[Modules.scala 65:57:@8155.4]
  wire [10:0] buffer_3_104; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60224; // @[Modules.scala 65:57:@8157.4]
  wire [10:0] _T_60225; // @[Modules.scala 65:57:@8158.4]
  wire [10:0] buffer_3_444; // @[Modules.scala 65:57:@8159.4]
  wire [10:0] buffer_3_106; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60227; // @[Modules.scala 65:57:@8161.4]
  wire [10:0] _T_60228; // @[Modules.scala 65:57:@8162.4]
  wire [10:0] buffer_3_445; // @[Modules.scala 65:57:@8163.4]
  wire [10:0] buffer_3_109; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60230; // @[Modules.scala 65:57:@8165.4]
  wire [10:0] _T_60231; // @[Modules.scala 65:57:@8166.4]
  wire [10:0] buffer_3_446; // @[Modules.scala 65:57:@8167.4]
  wire [10:0] buffer_3_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60236; // @[Modules.scala 65:57:@8173.4]
  wire [10:0] _T_60237; // @[Modules.scala 65:57:@8174.4]
  wire [10:0] buffer_3_448; // @[Modules.scala 65:57:@8175.4]
  wire [10:0] buffer_3_114; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60239; // @[Modules.scala 65:57:@8177.4]
  wire [10:0] _T_60240; // @[Modules.scala 65:57:@8178.4]
  wire [10:0] buffer_3_449; // @[Modules.scala 65:57:@8179.4]
  wire [10:0] buffer_3_116; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60242; // @[Modules.scala 65:57:@8181.4]
  wire [10:0] _T_60243; // @[Modules.scala 65:57:@8182.4]
  wire [10:0] buffer_3_450; // @[Modules.scala 65:57:@8183.4]
  wire [10:0] buffer_3_118; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60245; // @[Modules.scala 65:57:@8185.4]
  wire [10:0] _T_60246; // @[Modules.scala 65:57:@8186.4]
  wire [10:0] buffer_3_451; // @[Modules.scala 65:57:@8187.4]
  wire [10:0] buffer_3_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60248; // @[Modules.scala 65:57:@8189.4]
  wire [10:0] _T_60249; // @[Modules.scala 65:57:@8190.4]
  wire [10:0] buffer_3_452; // @[Modules.scala 65:57:@8191.4]
  wire [10:0] buffer_3_122; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60251; // @[Modules.scala 65:57:@8193.4]
  wire [10:0] _T_60252; // @[Modules.scala 65:57:@8194.4]
  wire [10:0] buffer_3_453; // @[Modules.scala 65:57:@8195.4]
  wire [10:0] buffer_3_126; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_127; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60257; // @[Modules.scala 65:57:@8201.4]
  wire [10:0] _T_60258; // @[Modules.scala 65:57:@8202.4]
  wire [10:0] buffer_3_455; // @[Modules.scala 65:57:@8203.4]
  wire [10:0] buffer_3_128; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60260; // @[Modules.scala 65:57:@8205.4]
  wire [10:0] _T_60261; // @[Modules.scala 65:57:@8206.4]
  wire [10:0] buffer_3_456; // @[Modules.scala 65:57:@8207.4]
  wire [10:0] buffer_3_132; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60266; // @[Modules.scala 65:57:@8213.4]
  wire [10:0] _T_60267; // @[Modules.scala 65:57:@8214.4]
  wire [10:0] buffer_3_458; // @[Modules.scala 65:57:@8215.4]
  wire [10:0] buffer_3_134; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60269; // @[Modules.scala 65:57:@8217.4]
  wire [10:0] _T_60270; // @[Modules.scala 65:57:@8218.4]
  wire [10:0] buffer_3_459; // @[Modules.scala 65:57:@8219.4]
  wire [10:0] buffer_3_136; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60272; // @[Modules.scala 65:57:@8221.4]
  wire [10:0] _T_60273; // @[Modules.scala 65:57:@8222.4]
  wire [10:0] buffer_3_460; // @[Modules.scala 65:57:@8223.4]
  wire [10:0] buffer_3_140; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60278; // @[Modules.scala 65:57:@8229.4]
  wire [10:0] _T_60279; // @[Modules.scala 65:57:@8230.4]
  wire [10:0] buffer_3_462; // @[Modules.scala 65:57:@8231.4]
  wire [10:0] buffer_3_142; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60281; // @[Modules.scala 65:57:@8233.4]
  wire [10:0] _T_60282; // @[Modules.scala 65:57:@8234.4]
  wire [10:0] buffer_3_463; // @[Modules.scala 65:57:@8235.4]
  wire [10:0] buffer_3_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60287; // @[Modules.scala 65:57:@8241.4]
  wire [10:0] _T_60288; // @[Modules.scala 65:57:@8242.4]
  wire [10:0] buffer_3_465; // @[Modules.scala 65:57:@8243.4]
  wire [10:0] buffer_3_148; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_149; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60290; // @[Modules.scala 65:57:@8245.4]
  wire [10:0] _T_60291; // @[Modules.scala 65:57:@8246.4]
  wire [10:0] buffer_3_466; // @[Modules.scala 65:57:@8247.4]
  wire [10:0] buffer_3_150; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60293; // @[Modules.scala 65:57:@8249.4]
  wire [10:0] _T_60294; // @[Modules.scala 65:57:@8250.4]
  wire [10:0] buffer_3_467; // @[Modules.scala 65:57:@8251.4]
  wire [10:0] buffer_3_154; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60299; // @[Modules.scala 65:57:@8257.4]
  wire [10:0] _T_60300; // @[Modules.scala 65:57:@8258.4]
  wire [10:0] buffer_3_469; // @[Modules.scala 65:57:@8259.4]
  wire [10:0] buffer_3_167; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60317; // @[Modules.scala 65:57:@8281.4]
  wire [10:0] _T_60318; // @[Modules.scala 65:57:@8282.4]
  wire [10:0] buffer_3_475; // @[Modules.scala 65:57:@8283.4]
  wire [10:0] buffer_3_168; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60320; // @[Modules.scala 65:57:@8285.4]
  wire [10:0] _T_60321; // @[Modules.scala 65:57:@8286.4]
  wire [10:0] buffer_3_476; // @[Modules.scala 65:57:@8287.4]
  wire [10:0] buffer_3_182; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60341; // @[Modules.scala 65:57:@8313.4]
  wire [10:0] _T_60342; // @[Modules.scala 65:57:@8314.4]
  wire [10:0] buffer_3_483; // @[Modules.scala 65:57:@8315.4]
  wire [10:0] buffer_3_187; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60347; // @[Modules.scala 65:57:@8321.4]
  wire [10:0] _T_60348; // @[Modules.scala 65:57:@8322.4]
  wire [10:0] buffer_3_485; // @[Modules.scala 65:57:@8323.4]
  wire [10:0] buffer_3_190; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60353; // @[Modules.scala 65:57:@8329.4]
  wire [10:0] _T_60354; // @[Modules.scala 65:57:@8330.4]
  wire [10:0] buffer_3_487; // @[Modules.scala 65:57:@8331.4]
  wire [10:0] buffer_3_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60359; // @[Modules.scala 65:57:@8337.4]
  wire [10:0] _T_60360; // @[Modules.scala 65:57:@8338.4]
  wire [10:0] buffer_3_489; // @[Modules.scala 65:57:@8339.4]
  wire [10:0] buffer_3_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60362; // @[Modules.scala 65:57:@8341.4]
  wire [10:0] _T_60363; // @[Modules.scala 65:57:@8342.4]
  wire [10:0] buffer_3_490; // @[Modules.scala 65:57:@8343.4]
  wire [10:0] buffer_3_200; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_201; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60368; // @[Modules.scala 65:57:@8349.4]
  wire [10:0] _T_60369; // @[Modules.scala 65:57:@8350.4]
  wire [10:0] buffer_3_492; // @[Modules.scala 65:57:@8351.4]
  wire [10:0] buffer_3_205; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60374; // @[Modules.scala 65:57:@8357.4]
  wire [10:0] _T_60375; // @[Modules.scala 65:57:@8358.4]
  wire [10:0] buffer_3_494; // @[Modules.scala 65:57:@8359.4]
  wire [10:0] buffer_3_208; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60380; // @[Modules.scala 65:57:@8365.4]
  wire [10:0] _T_60381; // @[Modules.scala 65:57:@8366.4]
  wire [10:0] buffer_3_496; // @[Modules.scala 65:57:@8367.4]
  wire [10:0] buffer_3_210; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60383; // @[Modules.scala 65:57:@8369.4]
  wire [10:0] _T_60384; // @[Modules.scala 65:57:@8370.4]
  wire [10:0] buffer_3_497; // @[Modules.scala 65:57:@8371.4]
  wire [10:0] buffer_3_212; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60386; // @[Modules.scala 65:57:@8373.4]
  wire [10:0] _T_60387; // @[Modules.scala 65:57:@8374.4]
  wire [10:0] buffer_3_498; // @[Modules.scala 65:57:@8375.4]
  wire [10:0] buffer_3_220; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60398; // @[Modules.scala 65:57:@8389.4]
  wire [10:0] _T_60399; // @[Modules.scala 65:57:@8390.4]
  wire [10:0] buffer_3_502; // @[Modules.scala 65:57:@8391.4]
  wire [10:0] buffer_3_222; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_223; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60401; // @[Modules.scala 65:57:@8393.4]
  wire [10:0] _T_60402; // @[Modules.scala 65:57:@8394.4]
  wire [10:0] buffer_3_503; // @[Modules.scala 65:57:@8395.4]
  wire [10:0] buffer_3_224; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60404; // @[Modules.scala 65:57:@8397.4]
  wire [10:0] _T_60405; // @[Modules.scala 65:57:@8398.4]
  wire [10:0] buffer_3_504; // @[Modules.scala 65:57:@8399.4]
  wire [10:0] buffer_3_226; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60407; // @[Modules.scala 65:57:@8401.4]
  wire [10:0] _T_60408; // @[Modules.scala 65:57:@8402.4]
  wire [10:0] buffer_3_505; // @[Modules.scala 65:57:@8403.4]
  wire [11:0] _T_60416; // @[Modules.scala 65:57:@8413.4]
  wire [10:0] _T_60417; // @[Modules.scala 65:57:@8414.4]
  wire [10:0] buffer_3_508; // @[Modules.scala 65:57:@8415.4]
  wire [10:0] buffer_3_236; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_237; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60422; // @[Modules.scala 65:57:@8421.4]
  wire [10:0] _T_60423; // @[Modules.scala 65:57:@8422.4]
  wire [10:0] buffer_3_510; // @[Modules.scala 65:57:@8423.4]
  wire [11:0] _T_60425; // @[Modules.scala 65:57:@8425.4]
  wire [10:0] _T_60426; // @[Modules.scala 65:57:@8426.4]
  wire [10:0] buffer_3_511; // @[Modules.scala 65:57:@8427.4]
  wire [10:0] buffer_3_240; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60428; // @[Modules.scala 65:57:@8429.4]
  wire [10:0] _T_60429; // @[Modules.scala 65:57:@8430.4]
  wire [10:0] buffer_3_512; // @[Modules.scala 65:57:@8431.4]
  wire [10:0] buffer_3_246; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60437; // @[Modules.scala 65:57:@8441.4]
  wire [10:0] _T_60438; // @[Modules.scala 65:57:@8442.4]
  wire [10:0] buffer_3_515; // @[Modules.scala 65:57:@8443.4]
  wire [10:0] buffer_3_250; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_251; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60443; // @[Modules.scala 65:57:@8449.4]
  wire [10:0] _T_60444; // @[Modules.scala 65:57:@8450.4]
  wire [10:0] buffer_3_517; // @[Modules.scala 65:57:@8451.4]
  wire [10:0] buffer_3_252; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60446; // @[Modules.scala 65:57:@8453.4]
  wire [10:0] _T_60447; // @[Modules.scala 65:57:@8454.4]
  wire [10:0] buffer_3_518; // @[Modules.scala 65:57:@8455.4]
  wire [10:0] buffer_3_254; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60449; // @[Modules.scala 65:57:@8457.4]
  wire [10:0] _T_60450; // @[Modules.scala 65:57:@8458.4]
  wire [10:0] buffer_3_519; // @[Modules.scala 65:57:@8459.4]
  wire [10:0] buffer_3_265; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60464; // @[Modules.scala 65:57:@8477.4]
  wire [10:0] _T_60465; // @[Modules.scala 65:57:@8478.4]
  wire [10:0] buffer_3_524; // @[Modules.scala 65:57:@8479.4]
  wire [10:0] buffer_3_270; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60473; // @[Modules.scala 65:57:@8489.4]
  wire [10:0] _T_60474; // @[Modules.scala 65:57:@8490.4]
  wire [10:0] buffer_3_527; // @[Modules.scala 65:57:@8491.4]
  wire [10:0] buffer_3_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60476; // @[Modules.scala 65:57:@8493.4]
  wire [10:0] _T_60477; // @[Modules.scala 65:57:@8494.4]
  wire [10:0] buffer_3_528; // @[Modules.scala 65:57:@8495.4]
  wire [10:0] buffer_3_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60482; // @[Modules.scala 65:57:@8501.4]
  wire [10:0] _T_60483; // @[Modules.scala 65:57:@8502.4]
  wire [10:0] buffer_3_530; // @[Modules.scala 65:57:@8503.4]
  wire [10:0] buffer_3_278; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60485; // @[Modules.scala 65:57:@8505.4]
  wire [10:0] _T_60486; // @[Modules.scala 65:57:@8506.4]
  wire [10:0] buffer_3_531; // @[Modules.scala 65:57:@8507.4]
  wire [11:0] _T_60488; // @[Modules.scala 65:57:@8509.4]
  wire [10:0] _T_60489; // @[Modules.scala 65:57:@8510.4]
  wire [10:0] buffer_3_532; // @[Modules.scala 65:57:@8511.4]
  wire [10:0] buffer_3_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60491; // @[Modules.scala 65:57:@8513.4]
  wire [10:0] _T_60492; // @[Modules.scala 65:57:@8514.4]
  wire [10:0] buffer_3_533; // @[Modules.scala 65:57:@8515.4]
  wire [10:0] buffer_3_286; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60497; // @[Modules.scala 65:57:@8521.4]
  wire [10:0] _T_60498; // @[Modules.scala 65:57:@8522.4]
  wire [10:0] buffer_3_535; // @[Modules.scala 65:57:@8523.4]
  wire [11:0] _T_60500; // @[Modules.scala 65:57:@8525.4]
  wire [10:0] _T_60501; // @[Modules.scala 65:57:@8526.4]
  wire [10:0] buffer_3_536; // @[Modules.scala 65:57:@8527.4]
  wire [10:0] buffer_3_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60503; // @[Modules.scala 65:57:@8529.4]
  wire [10:0] _T_60504; // @[Modules.scala 65:57:@8530.4]
  wire [10:0] buffer_3_537; // @[Modules.scala 65:57:@8531.4]
  wire [10:0] buffer_3_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60506; // @[Modules.scala 65:57:@8533.4]
  wire [10:0] _T_60507; // @[Modules.scala 65:57:@8534.4]
  wire [10:0] buffer_3_538; // @[Modules.scala 65:57:@8535.4]
  wire [10:0] buffer_3_297; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60512; // @[Modules.scala 65:57:@8541.4]
  wire [10:0] _T_60513; // @[Modules.scala 65:57:@8542.4]
  wire [10:0] buffer_3_540; // @[Modules.scala 65:57:@8543.4]
  wire [11:0] _T_60515; // @[Modules.scala 65:57:@8545.4]
  wire [10:0] _T_60516; // @[Modules.scala 65:57:@8546.4]
  wire [10:0] buffer_3_541; // @[Modules.scala 65:57:@8547.4]
  wire [11:0] _T_60518; // @[Modules.scala 65:57:@8549.4]
  wire [10:0] _T_60519; // @[Modules.scala 65:57:@8550.4]
  wire [10:0] buffer_3_542; // @[Modules.scala 65:57:@8551.4]
  wire [11:0] _T_60521; // @[Modules.scala 65:57:@8553.4]
  wire [10:0] _T_60522; // @[Modules.scala 65:57:@8554.4]
  wire [10:0] buffer_3_543; // @[Modules.scala 65:57:@8555.4]
  wire [10:0] buffer_3_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60524; // @[Modules.scala 65:57:@8557.4]
  wire [10:0] _T_60525; // @[Modules.scala 65:57:@8558.4]
  wire [10:0] buffer_3_544; // @[Modules.scala 65:57:@8559.4]
  wire [10:0] buffer_3_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60527; // @[Modules.scala 65:57:@8561.4]
  wire [10:0] _T_60528; // @[Modules.scala 65:57:@8562.4]
  wire [10:0] buffer_3_545; // @[Modules.scala 65:57:@8563.4]
  wire [10:0] buffer_3_310; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60533; // @[Modules.scala 65:57:@8569.4]
  wire [10:0] _T_60534; // @[Modules.scala 65:57:@8570.4]
  wire [10:0] buffer_3_547; // @[Modules.scala 65:57:@8571.4]
  wire [10:0] buffer_3_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60536; // @[Modules.scala 65:57:@8573.4]
  wire [10:0] _T_60537; // @[Modules.scala 65:57:@8574.4]
  wire [10:0] buffer_3_548; // @[Modules.scala 65:57:@8575.4]
  wire [10:0] buffer_3_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60539; // @[Modules.scala 65:57:@8577.4]
  wire [10:0] _T_60540; // @[Modules.scala 65:57:@8578.4]
  wire [10:0] buffer_3_549; // @[Modules.scala 65:57:@8579.4]
  wire [10:0] buffer_3_316; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_317; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60542; // @[Modules.scala 65:57:@8581.4]
  wire [10:0] _T_60543; // @[Modules.scala 65:57:@8582.4]
  wire [10:0] buffer_3_550; // @[Modules.scala 65:57:@8583.4]
  wire [10:0] buffer_3_319; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60545; // @[Modules.scala 65:57:@8585.4]
  wire [10:0] _T_60546; // @[Modules.scala 65:57:@8586.4]
  wire [10:0] buffer_3_551; // @[Modules.scala 65:57:@8587.4]
  wire [10:0] buffer_3_321; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60548; // @[Modules.scala 65:57:@8589.4]
  wire [10:0] _T_60549; // @[Modules.scala 65:57:@8590.4]
  wire [10:0] buffer_3_552; // @[Modules.scala 65:57:@8591.4]
  wire [11:0] _T_60551; // @[Modules.scala 65:57:@8593.4]
  wire [10:0] _T_60552; // @[Modules.scala 65:57:@8594.4]
  wire [10:0] buffer_3_553; // @[Modules.scala 65:57:@8595.4]
  wire [10:0] buffer_3_325; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60554; // @[Modules.scala 65:57:@8597.4]
  wire [10:0] _T_60555; // @[Modules.scala 65:57:@8598.4]
  wire [10:0] buffer_3_554; // @[Modules.scala 65:57:@8599.4]
  wire [10:0] buffer_3_326; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60557; // @[Modules.scala 65:57:@8601.4]
  wire [10:0] _T_60558; // @[Modules.scala 65:57:@8602.4]
  wire [10:0] buffer_3_555; // @[Modules.scala 65:57:@8603.4]
  wire [11:0] _T_60560; // @[Modules.scala 65:57:@8605.4]
  wire [10:0] _T_60561; // @[Modules.scala 65:57:@8606.4]
  wire [10:0] buffer_3_556; // @[Modules.scala 65:57:@8607.4]
  wire [10:0] buffer_3_333; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60566; // @[Modules.scala 65:57:@8613.4]
  wire [10:0] _T_60567; // @[Modules.scala 65:57:@8614.4]
  wire [10:0] buffer_3_558; // @[Modules.scala 65:57:@8615.4]
  wire [10:0] buffer_3_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60569; // @[Modules.scala 65:57:@8617.4]
  wire [10:0] _T_60570; // @[Modules.scala 65:57:@8618.4]
  wire [10:0] buffer_3_559; // @[Modules.scala 65:57:@8619.4]
  wire [10:0] buffer_3_336; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_337; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60572; // @[Modules.scala 65:57:@8621.4]
  wire [10:0] _T_60573; // @[Modules.scala 65:57:@8622.4]
  wire [10:0] buffer_3_560; // @[Modules.scala 65:57:@8623.4]
  wire [11:0] _T_60578; // @[Modules.scala 65:57:@8629.4]
  wire [10:0] _T_60579; // @[Modules.scala 65:57:@8630.4]
  wire [10:0] buffer_3_562; // @[Modules.scala 65:57:@8631.4]
  wire [10:0] buffer_3_342; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60581; // @[Modules.scala 65:57:@8633.4]
  wire [10:0] _T_60582; // @[Modules.scala 65:57:@8634.4]
  wire [10:0] buffer_3_563; // @[Modules.scala 65:57:@8635.4]
  wire [10:0] buffer_3_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60590; // @[Modules.scala 65:57:@8645.4]
  wire [10:0] _T_60591; // @[Modules.scala 65:57:@8646.4]
  wire [10:0] buffer_3_566; // @[Modules.scala 65:57:@8647.4]
  wire [10:0] buffer_3_351; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60593; // @[Modules.scala 65:57:@8649.4]
  wire [10:0] _T_60594; // @[Modules.scala 65:57:@8650.4]
  wire [10:0] buffer_3_567; // @[Modules.scala 65:57:@8651.4]
  wire [10:0] buffer_3_355; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60599; // @[Modules.scala 65:57:@8657.4]
  wire [10:0] _T_60600; // @[Modules.scala 65:57:@8658.4]
  wire [10:0] buffer_3_569; // @[Modules.scala 65:57:@8659.4]
  wire [11:0] _T_60611; // @[Modules.scala 65:57:@8673.4]
  wire [10:0] _T_60612; // @[Modules.scala 65:57:@8674.4]
  wire [10:0] buffer_3_573; // @[Modules.scala 65:57:@8675.4]
  wire [10:0] buffer_3_365; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60614; // @[Modules.scala 65:57:@8677.4]
  wire [10:0] _T_60615; // @[Modules.scala 65:57:@8678.4]
  wire [10:0] buffer_3_574; // @[Modules.scala 65:57:@8679.4]
  wire [10:0] buffer_3_368; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_369; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60620; // @[Modules.scala 65:57:@8685.4]
  wire [10:0] _T_60621; // @[Modules.scala 65:57:@8686.4]
  wire [10:0] buffer_3_576; // @[Modules.scala 65:57:@8687.4]
  wire [10:0] buffer_3_370; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60623; // @[Modules.scala 65:57:@8689.4]
  wire [10:0] _T_60624; // @[Modules.scala 65:57:@8690.4]
  wire [10:0] buffer_3_577; // @[Modules.scala 65:57:@8691.4]
  wire [10:0] buffer_3_372; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_373; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60626; // @[Modules.scala 65:57:@8693.4]
  wire [10:0] _T_60627; // @[Modules.scala 65:57:@8694.4]
  wire [10:0] buffer_3_578; // @[Modules.scala 65:57:@8695.4]
  wire [11:0] _T_60629; // @[Modules.scala 65:57:@8697.4]
  wire [10:0] _T_60630; // @[Modules.scala 65:57:@8698.4]
  wire [10:0] buffer_3_579; // @[Modules.scala 65:57:@8699.4]
  wire [10:0] buffer_3_376; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_377; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60632; // @[Modules.scala 65:57:@8701.4]
  wire [10:0] _T_60633; // @[Modules.scala 65:57:@8702.4]
  wire [10:0] buffer_3_580; // @[Modules.scala 65:57:@8703.4]
  wire [10:0] buffer_3_378; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60635; // @[Modules.scala 65:57:@8705.4]
  wire [10:0] _T_60636; // @[Modules.scala 65:57:@8706.4]
  wire [10:0] buffer_3_581; // @[Modules.scala 65:57:@8707.4]
  wire [10:0] buffer_3_382; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60641; // @[Modules.scala 65:57:@8713.4]
  wire [10:0] _T_60642; // @[Modules.scala 65:57:@8714.4]
  wire [10:0] buffer_3_583; // @[Modules.scala 65:57:@8715.4]
  wire [10:0] buffer_3_384; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_385; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60644; // @[Modules.scala 65:57:@8717.4]
  wire [10:0] _T_60645; // @[Modules.scala 65:57:@8718.4]
  wire [10:0] buffer_3_584; // @[Modules.scala 65:57:@8719.4]
  wire [10:0] buffer_3_386; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_3_387; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60647; // @[Modules.scala 65:57:@8721.4]
  wire [10:0] _T_60648; // @[Modules.scala 65:57:@8722.4]
  wire [10:0] buffer_3_585; // @[Modules.scala 65:57:@8723.4]
  wire [10:0] buffer_3_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_60650; // @[Modules.scala 65:57:@8725.4]
  wire [10:0] _T_60651; // @[Modules.scala 65:57:@8726.4]
  wire [10:0] buffer_3_586; // @[Modules.scala 65:57:@8727.4]
  wire [11:0] _T_60653; // @[Modules.scala 65:57:@8729.4]
  wire [10:0] _T_60654; // @[Modules.scala 65:57:@8730.4]
  wire [10:0] buffer_3_587; // @[Modules.scala 65:57:@8731.4]
  wire [11:0] _T_60656; // @[Modules.scala 68:83:@8733.4]
  wire [10:0] _T_60657; // @[Modules.scala 68:83:@8734.4]
  wire [10:0] buffer_3_588; // @[Modules.scala 68:83:@8735.4]
  wire [11:0] _T_60659; // @[Modules.scala 68:83:@8737.4]
  wire [10:0] _T_60660; // @[Modules.scala 68:83:@8738.4]
  wire [10:0] buffer_3_589; // @[Modules.scala 68:83:@8739.4]
  wire [11:0] _T_60662; // @[Modules.scala 68:83:@8741.4]
  wire [10:0] _T_60663; // @[Modules.scala 68:83:@8742.4]
  wire [10:0] buffer_3_590; // @[Modules.scala 68:83:@8743.4]
  wire [11:0] _T_60665; // @[Modules.scala 68:83:@8745.4]
  wire [10:0] _T_60666; // @[Modules.scala 68:83:@8746.4]
  wire [10:0] buffer_3_591; // @[Modules.scala 68:83:@8747.4]
  wire [11:0] _T_60668; // @[Modules.scala 68:83:@8749.4]
  wire [10:0] _T_60669; // @[Modules.scala 68:83:@8750.4]
  wire [10:0] buffer_3_592; // @[Modules.scala 68:83:@8751.4]
  wire [11:0] _T_60671; // @[Modules.scala 68:83:@8753.4]
  wire [10:0] _T_60672; // @[Modules.scala 68:83:@8754.4]
  wire [10:0] buffer_3_593; // @[Modules.scala 68:83:@8755.4]
  wire [11:0] _T_60674; // @[Modules.scala 68:83:@8757.4]
  wire [10:0] _T_60675; // @[Modules.scala 68:83:@8758.4]
  wire [10:0] buffer_3_594; // @[Modules.scala 68:83:@8759.4]
  wire [11:0] _T_60677; // @[Modules.scala 68:83:@8761.4]
  wire [10:0] _T_60678; // @[Modules.scala 68:83:@8762.4]
  wire [10:0] buffer_3_595; // @[Modules.scala 68:83:@8763.4]
  wire [11:0] _T_60686; // @[Modules.scala 68:83:@8773.4]
  wire [10:0] _T_60687; // @[Modules.scala 68:83:@8774.4]
  wire [10:0] buffer_3_598; // @[Modules.scala 68:83:@8775.4]
  wire [11:0] _T_60689; // @[Modules.scala 68:83:@8777.4]
  wire [10:0] _T_60690; // @[Modules.scala 68:83:@8778.4]
  wire [10:0] buffer_3_599; // @[Modules.scala 68:83:@8779.4]
  wire [11:0] _T_60692; // @[Modules.scala 68:83:@8781.4]
  wire [10:0] _T_60693; // @[Modules.scala 68:83:@8782.4]
  wire [10:0] buffer_3_600; // @[Modules.scala 68:83:@8783.4]
  wire [11:0] _T_60695; // @[Modules.scala 68:83:@8785.4]
  wire [10:0] _T_60696; // @[Modules.scala 68:83:@8786.4]
  wire [10:0] buffer_3_601; // @[Modules.scala 68:83:@8787.4]
  wire [11:0] _T_60698; // @[Modules.scala 68:83:@8789.4]
  wire [10:0] _T_60699; // @[Modules.scala 68:83:@8790.4]
  wire [10:0] buffer_3_602; // @[Modules.scala 68:83:@8791.4]
  wire [11:0] _T_60701; // @[Modules.scala 68:83:@8793.4]
  wire [10:0] _T_60702; // @[Modules.scala 68:83:@8794.4]
  wire [10:0] buffer_3_603; // @[Modules.scala 68:83:@8795.4]
  wire [11:0] _T_60704; // @[Modules.scala 68:83:@8797.4]
  wire [10:0] _T_60705; // @[Modules.scala 68:83:@8798.4]
  wire [10:0] buffer_3_604; // @[Modules.scala 68:83:@8799.4]
  wire [11:0] _T_60707; // @[Modules.scala 68:83:@8801.4]
  wire [10:0] _T_60708; // @[Modules.scala 68:83:@8802.4]
  wire [10:0] buffer_3_605; // @[Modules.scala 68:83:@8803.4]
  wire [11:0] _T_60710; // @[Modules.scala 68:83:@8805.4]
  wire [10:0] _T_60711; // @[Modules.scala 68:83:@8806.4]
  wire [10:0] buffer_3_606; // @[Modules.scala 68:83:@8807.4]
  wire [11:0] _T_60713; // @[Modules.scala 68:83:@8809.4]
  wire [10:0] _T_60714; // @[Modules.scala 68:83:@8810.4]
  wire [10:0] buffer_3_607; // @[Modules.scala 68:83:@8811.4]
  wire [11:0] _T_60719; // @[Modules.scala 68:83:@8817.4]
  wire [10:0] _T_60720; // @[Modules.scala 68:83:@8818.4]
  wire [10:0] buffer_3_609; // @[Modules.scala 68:83:@8819.4]
  wire [11:0] _T_60722; // @[Modules.scala 68:83:@8821.4]
  wire [10:0] _T_60723; // @[Modules.scala 68:83:@8822.4]
  wire [10:0] buffer_3_610; // @[Modules.scala 68:83:@8823.4]
  wire [11:0] _T_60725; // @[Modules.scala 68:83:@8825.4]
  wire [10:0] _T_60726; // @[Modules.scala 68:83:@8826.4]
  wire [10:0] buffer_3_611; // @[Modules.scala 68:83:@8827.4]
  wire [11:0] _T_60728; // @[Modules.scala 68:83:@8829.4]
  wire [10:0] _T_60729; // @[Modules.scala 68:83:@8830.4]
  wire [10:0] buffer_3_612; // @[Modules.scala 68:83:@8831.4]
  wire [11:0] _T_60731; // @[Modules.scala 68:83:@8833.4]
  wire [10:0] _T_60732; // @[Modules.scala 68:83:@8834.4]
  wire [10:0] buffer_3_613; // @[Modules.scala 68:83:@8835.4]
  wire [11:0] _T_60734; // @[Modules.scala 68:83:@8837.4]
  wire [10:0] _T_60735; // @[Modules.scala 68:83:@8838.4]
  wire [10:0] buffer_3_614; // @[Modules.scala 68:83:@8839.4]
  wire [11:0] _T_60737; // @[Modules.scala 68:83:@8841.4]
  wire [10:0] _T_60738; // @[Modules.scala 68:83:@8842.4]
  wire [10:0] buffer_3_615; // @[Modules.scala 68:83:@8843.4]
  wire [11:0] _T_60740; // @[Modules.scala 68:83:@8845.4]
  wire [10:0] _T_60741; // @[Modules.scala 68:83:@8846.4]
  wire [10:0] buffer_3_616; // @[Modules.scala 68:83:@8847.4]
  wire [11:0] _T_60743; // @[Modules.scala 68:83:@8849.4]
  wire [10:0] _T_60744; // @[Modules.scala 68:83:@8850.4]
  wire [10:0] buffer_3_617; // @[Modules.scala 68:83:@8851.4]
  wire [11:0] _T_60746; // @[Modules.scala 68:83:@8853.4]
  wire [10:0] _T_60747; // @[Modules.scala 68:83:@8854.4]
  wire [10:0] buffer_3_618; // @[Modules.scala 68:83:@8855.4]
  wire [11:0] _T_60749; // @[Modules.scala 68:83:@8857.4]
  wire [10:0] _T_60750; // @[Modules.scala 68:83:@8858.4]
  wire [10:0] buffer_3_619; // @[Modules.scala 68:83:@8859.4]
  wire [11:0] _T_60752; // @[Modules.scala 68:83:@8861.4]
  wire [10:0] _T_60753; // @[Modules.scala 68:83:@8862.4]
  wire [10:0] buffer_3_620; // @[Modules.scala 68:83:@8863.4]
  wire [11:0] _T_60755; // @[Modules.scala 68:83:@8865.4]
  wire [10:0] _T_60756; // @[Modules.scala 68:83:@8866.4]
  wire [10:0] buffer_3_621; // @[Modules.scala 68:83:@8867.4]
  wire [11:0] _T_60758; // @[Modules.scala 68:83:@8869.4]
  wire [10:0] _T_60759; // @[Modules.scala 68:83:@8870.4]
  wire [10:0] buffer_3_622; // @[Modules.scala 68:83:@8871.4]
  wire [11:0] _T_60761; // @[Modules.scala 68:83:@8873.4]
  wire [10:0] _T_60762; // @[Modules.scala 68:83:@8874.4]
  wire [10:0] buffer_3_623; // @[Modules.scala 68:83:@8875.4]
  wire [11:0] _T_60764; // @[Modules.scala 68:83:@8877.4]
  wire [10:0] _T_60765; // @[Modules.scala 68:83:@8878.4]
  wire [10:0] buffer_3_624; // @[Modules.scala 68:83:@8879.4]
  wire [11:0] _T_60767; // @[Modules.scala 68:83:@8881.4]
  wire [10:0] _T_60768; // @[Modules.scala 68:83:@8882.4]
  wire [10:0] buffer_3_625; // @[Modules.scala 68:83:@8883.4]
  wire [11:0] _T_60770; // @[Modules.scala 68:83:@8885.4]
  wire [10:0] _T_60771; // @[Modules.scala 68:83:@8886.4]
  wire [10:0] buffer_3_626; // @[Modules.scala 68:83:@8887.4]
  wire [11:0] _T_60779; // @[Modules.scala 68:83:@8897.4]
  wire [10:0] _T_60780; // @[Modules.scala 68:83:@8898.4]
  wire [10:0] buffer_3_629; // @[Modules.scala 68:83:@8899.4]
  wire [11:0] _T_60782; // @[Modules.scala 68:83:@8901.4]
  wire [10:0] _T_60783; // @[Modules.scala 68:83:@8902.4]
  wire [10:0] buffer_3_630; // @[Modules.scala 68:83:@8903.4]
  wire [11:0] _T_60791; // @[Modules.scala 68:83:@8913.4]
  wire [10:0] _T_60792; // @[Modules.scala 68:83:@8914.4]
  wire [10:0] buffer_3_633; // @[Modules.scala 68:83:@8915.4]
  wire [11:0] _T_60794; // @[Modules.scala 68:83:@8917.4]
  wire [10:0] _T_60795; // @[Modules.scala 68:83:@8918.4]
  wire [10:0] buffer_3_634; // @[Modules.scala 68:83:@8919.4]
  wire [11:0] _T_60797; // @[Modules.scala 68:83:@8921.4]
  wire [10:0] _T_60798; // @[Modules.scala 68:83:@8922.4]
  wire [10:0] buffer_3_635; // @[Modules.scala 68:83:@8923.4]
  wire [11:0] _T_60800; // @[Modules.scala 68:83:@8925.4]
  wire [10:0] _T_60801; // @[Modules.scala 68:83:@8926.4]
  wire [10:0] buffer_3_636; // @[Modules.scala 68:83:@8927.4]
  wire [11:0] _T_60803; // @[Modules.scala 68:83:@8929.4]
  wire [10:0] _T_60804; // @[Modules.scala 68:83:@8930.4]
  wire [10:0] buffer_3_637; // @[Modules.scala 68:83:@8931.4]
  wire [11:0] _T_60806; // @[Modules.scala 68:83:@8933.4]
  wire [10:0] _T_60807; // @[Modules.scala 68:83:@8934.4]
  wire [10:0] buffer_3_638; // @[Modules.scala 68:83:@8935.4]
  wire [11:0] _T_60809; // @[Modules.scala 68:83:@8937.4]
  wire [10:0] _T_60810; // @[Modules.scala 68:83:@8938.4]
  wire [10:0] buffer_3_639; // @[Modules.scala 68:83:@8939.4]
  wire [11:0] _T_60812; // @[Modules.scala 68:83:@8941.4]
  wire [10:0] _T_60813; // @[Modules.scala 68:83:@8942.4]
  wire [10:0] buffer_3_640; // @[Modules.scala 68:83:@8943.4]
  wire [11:0] _T_60815; // @[Modules.scala 68:83:@8945.4]
  wire [10:0] _T_60816; // @[Modules.scala 68:83:@8946.4]
  wire [10:0] buffer_3_641; // @[Modules.scala 68:83:@8947.4]
  wire [11:0] _T_60821; // @[Modules.scala 68:83:@8953.4]
  wire [10:0] _T_60822; // @[Modules.scala 68:83:@8954.4]
  wire [10:0] buffer_3_643; // @[Modules.scala 68:83:@8955.4]
  wire [11:0] _T_60824; // @[Modules.scala 68:83:@8957.4]
  wire [10:0] _T_60825; // @[Modules.scala 68:83:@8958.4]
  wire [10:0] buffer_3_644; // @[Modules.scala 68:83:@8959.4]
  wire [11:0] _T_60830; // @[Modules.scala 68:83:@8965.4]
  wire [10:0] _T_60831; // @[Modules.scala 68:83:@8966.4]
  wire [10:0] buffer_3_646; // @[Modules.scala 68:83:@8967.4]
  wire [11:0] _T_60833; // @[Modules.scala 68:83:@8969.4]
  wire [10:0] _T_60834; // @[Modules.scala 68:83:@8970.4]
  wire [10:0] buffer_3_647; // @[Modules.scala 68:83:@8971.4]
  wire [11:0] _T_60836; // @[Modules.scala 68:83:@8973.4]
  wire [10:0] _T_60837; // @[Modules.scala 68:83:@8974.4]
  wire [10:0] buffer_3_648; // @[Modules.scala 68:83:@8975.4]
  wire [11:0] _T_60839; // @[Modules.scala 68:83:@8977.4]
  wire [10:0] _T_60840; // @[Modules.scala 68:83:@8978.4]
  wire [10:0] buffer_3_649; // @[Modules.scala 68:83:@8979.4]
  wire [11:0] _T_60842; // @[Modules.scala 68:83:@8981.4]
  wire [10:0] _T_60843; // @[Modules.scala 68:83:@8982.4]
  wire [10:0] buffer_3_650; // @[Modules.scala 68:83:@8983.4]
  wire [11:0] _T_60845; // @[Modules.scala 68:83:@8985.4]
  wire [10:0] _T_60846; // @[Modules.scala 68:83:@8986.4]
  wire [10:0] buffer_3_651; // @[Modules.scala 68:83:@8987.4]
  wire [11:0] _T_60851; // @[Modules.scala 68:83:@8993.4]
  wire [10:0] _T_60852; // @[Modules.scala 68:83:@8994.4]
  wire [10:0] buffer_3_653; // @[Modules.scala 68:83:@8995.4]
  wire [11:0] _T_60854; // @[Modules.scala 68:83:@8997.4]
  wire [10:0] _T_60855; // @[Modules.scala 68:83:@8998.4]
  wire [10:0] buffer_3_654; // @[Modules.scala 68:83:@8999.4]
  wire [11:0] _T_60857; // @[Modules.scala 68:83:@9001.4]
  wire [10:0] _T_60858; // @[Modules.scala 68:83:@9002.4]
  wire [10:0] buffer_3_655; // @[Modules.scala 68:83:@9003.4]
  wire [11:0] _T_60860; // @[Modules.scala 68:83:@9005.4]
  wire [10:0] _T_60861; // @[Modules.scala 68:83:@9006.4]
  wire [10:0] buffer_3_656; // @[Modules.scala 68:83:@9007.4]
  wire [11:0] _T_60863; // @[Modules.scala 68:83:@9009.4]
  wire [10:0] _T_60864; // @[Modules.scala 68:83:@9010.4]
  wire [10:0] buffer_3_657; // @[Modules.scala 68:83:@9011.4]
  wire [11:0] _T_60866; // @[Modules.scala 68:83:@9013.4]
  wire [10:0] _T_60867; // @[Modules.scala 68:83:@9014.4]
  wire [10:0] buffer_3_658; // @[Modules.scala 68:83:@9015.4]
  wire [11:0] _T_60869; // @[Modules.scala 68:83:@9017.4]
  wire [10:0] _T_60870; // @[Modules.scala 68:83:@9018.4]
  wire [10:0] buffer_3_659; // @[Modules.scala 68:83:@9019.4]
  wire [11:0] _T_60872; // @[Modules.scala 68:83:@9021.4]
  wire [10:0] _T_60873; // @[Modules.scala 68:83:@9022.4]
  wire [10:0] buffer_3_660; // @[Modules.scala 68:83:@9023.4]
  wire [11:0] _T_60875; // @[Modules.scala 68:83:@9025.4]
  wire [10:0] _T_60876; // @[Modules.scala 68:83:@9026.4]
  wire [10:0] buffer_3_661; // @[Modules.scala 68:83:@9027.4]
  wire [11:0] _T_60878; // @[Modules.scala 68:83:@9029.4]
  wire [10:0] _T_60879; // @[Modules.scala 68:83:@9030.4]
  wire [10:0] buffer_3_662; // @[Modules.scala 68:83:@9031.4]
  wire [11:0] _T_60881; // @[Modules.scala 68:83:@9033.4]
  wire [10:0] _T_60882; // @[Modules.scala 68:83:@9034.4]
  wire [10:0] buffer_3_663; // @[Modules.scala 68:83:@9035.4]
  wire [11:0] _T_60884; // @[Modules.scala 68:83:@9037.4]
  wire [10:0] _T_60885; // @[Modules.scala 68:83:@9038.4]
  wire [10:0] buffer_3_664; // @[Modules.scala 68:83:@9039.4]
  wire [11:0] _T_60887; // @[Modules.scala 68:83:@9041.4]
  wire [10:0] _T_60888; // @[Modules.scala 68:83:@9042.4]
  wire [10:0] buffer_3_665; // @[Modules.scala 68:83:@9043.4]
  wire [11:0] _T_60890; // @[Modules.scala 68:83:@9045.4]
  wire [10:0] _T_60891; // @[Modules.scala 68:83:@9046.4]
  wire [10:0] buffer_3_666; // @[Modules.scala 68:83:@9047.4]
  wire [11:0] _T_60893; // @[Modules.scala 68:83:@9049.4]
  wire [10:0] _T_60894; // @[Modules.scala 68:83:@9050.4]
  wire [10:0] buffer_3_667; // @[Modules.scala 68:83:@9051.4]
  wire [11:0] _T_60896; // @[Modules.scala 68:83:@9053.4]
  wire [10:0] _T_60897; // @[Modules.scala 68:83:@9054.4]
  wire [10:0] buffer_3_668; // @[Modules.scala 68:83:@9055.4]
  wire [11:0] _T_60899; // @[Modules.scala 68:83:@9057.4]
  wire [10:0] _T_60900; // @[Modules.scala 68:83:@9058.4]
  wire [10:0] buffer_3_669; // @[Modules.scala 68:83:@9059.4]
  wire [11:0] _T_60902; // @[Modules.scala 68:83:@9061.4]
  wire [10:0] _T_60903; // @[Modules.scala 68:83:@9062.4]
  wire [10:0] buffer_3_670; // @[Modules.scala 68:83:@9063.4]
  wire [11:0] _T_60905; // @[Modules.scala 68:83:@9065.4]
  wire [10:0] _T_60906; // @[Modules.scala 68:83:@9066.4]
  wire [10:0] buffer_3_671; // @[Modules.scala 68:83:@9067.4]
  wire [11:0] _T_60908; // @[Modules.scala 68:83:@9069.4]
  wire [10:0] _T_60909; // @[Modules.scala 68:83:@9070.4]
  wire [10:0] buffer_3_672; // @[Modules.scala 68:83:@9071.4]
  wire [11:0] _T_60911; // @[Modules.scala 68:83:@9073.4]
  wire [10:0] _T_60912; // @[Modules.scala 68:83:@9074.4]
  wire [10:0] buffer_3_673; // @[Modules.scala 68:83:@9075.4]
  wire [11:0] _T_60917; // @[Modules.scala 68:83:@9081.4]
  wire [10:0] _T_60918; // @[Modules.scala 68:83:@9082.4]
  wire [10:0] buffer_3_675; // @[Modules.scala 68:83:@9083.4]
  wire [11:0] _T_60920; // @[Modules.scala 68:83:@9085.4]
  wire [10:0] _T_60921; // @[Modules.scala 68:83:@9086.4]
  wire [10:0] buffer_3_676; // @[Modules.scala 68:83:@9087.4]
  wire [11:0] _T_60923; // @[Modules.scala 68:83:@9089.4]
  wire [10:0] _T_60924; // @[Modules.scala 68:83:@9090.4]
  wire [10:0] buffer_3_677; // @[Modules.scala 68:83:@9091.4]
  wire [11:0] _T_60926; // @[Modules.scala 68:83:@9093.4]
  wire [10:0] _T_60927; // @[Modules.scala 68:83:@9094.4]
  wire [10:0] buffer_3_678; // @[Modules.scala 68:83:@9095.4]
  wire [11:0] _T_60929; // @[Modules.scala 68:83:@9097.4]
  wire [10:0] _T_60930; // @[Modules.scala 68:83:@9098.4]
  wire [10:0] buffer_3_679; // @[Modules.scala 68:83:@9099.4]
  wire [11:0] _T_60932; // @[Modules.scala 68:83:@9101.4]
  wire [10:0] _T_60933; // @[Modules.scala 68:83:@9102.4]
  wire [10:0] buffer_3_680; // @[Modules.scala 68:83:@9103.4]
  wire [11:0] _T_60935; // @[Modules.scala 68:83:@9105.4]
  wire [10:0] _T_60936; // @[Modules.scala 68:83:@9106.4]
  wire [10:0] buffer_3_681; // @[Modules.scala 68:83:@9107.4]
  wire [11:0] _T_60938; // @[Modules.scala 68:83:@9109.4]
  wire [10:0] _T_60939; // @[Modules.scala 68:83:@9110.4]
  wire [10:0] buffer_3_682; // @[Modules.scala 68:83:@9111.4]
  wire [11:0] _T_60941; // @[Modules.scala 68:83:@9113.4]
  wire [10:0] _T_60942; // @[Modules.scala 68:83:@9114.4]
  wire [10:0] buffer_3_683; // @[Modules.scala 68:83:@9115.4]
  wire [11:0] _T_60944; // @[Modules.scala 68:83:@9117.4]
  wire [10:0] _T_60945; // @[Modules.scala 68:83:@9118.4]
  wire [10:0] buffer_3_684; // @[Modules.scala 68:83:@9119.4]
  wire [11:0] _T_60947; // @[Modules.scala 68:83:@9121.4]
  wire [10:0] _T_60948; // @[Modules.scala 68:83:@9122.4]
  wire [10:0] buffer_3_685; // @[Modules.scala 68:83:@9123.4]
  wire [11:0] _T_60950; // @[Modules.scala 71:109:@9125.4]
  wire [10:0] _T_60951; // @[Modules.scala 71:109:@9126.4]
  wire [10:0] buffer_3_686; // @[Modules.scala 71:109:@9127.4]
  wire [11:0] _T_60953; // @[Modules.scala 71:109:@9129.4]
  wire [10:0] _T_60954; // @[Modules.scala 71:109:@9130.4]
  wire [10:0] buffer_3_687; // @[Modules.scala 71:109:@9131.4]
  wire [11:0] _T_60956; // @[Modules.scala 71:109:@9133.4]
  wire [10:0] _T_60957; // @[Modules.scala 71:109:@9134.4]
  wire [10:0] buffer_3_688; // @[Modules.scala 71:109:@9135.4]
  wire [11:0] _T_60959; // @[Modules.scala 71:109:@9137.4]
  wire [10:0] _T_60960; // @[Modules.scala 71:109:@9138.4]
  wire [10:0] buffer_3_689; // @[Modules.scala 71:109:@9139.4]
  wire [11:0] _T_60965; // @[Modules.scala 71:109:@9145.4]
  wire [10:0] _T_60966; // @[Modules.scala 71:109:@9146.4]
  wire [10:0] buffer_3_691; // @[Modules.scala 71:109:@9147.4]
  wire [11:0] _T_60968; // @[Modules.scala 71:109:@9149.4]
  wire [10:0] _T_60969; // @[Modules.scala 71:109:@9150.4]
  wire [10:0] buffer_3_692; // @[Modules.scala 71:109:@9151.4]
  wire [11:0] _T_60971; // @[Modules.scala 71:109:@9153.4]
  wire [10:0] _T_60972; // @[Modules.scala 71:109:@9154.4]
  wire [10:0] buffer_3_693; // @[Modules.scala 71:109:@9155.4]
  wire [11:0] _T_60974; // @[Modules.scala 71:109:@9157.4]
  wire [10:0] _T_60975; // @[Modules.scala 71:109:@9158.4]
  wire [10:0] buffer_3_694; // @[Modules.scala 71:109:@9159.4]
  wire [11:0] _T_60977; // @[Modules.scala 71:109:@9161.4]
  wire [10:0] _T_60978; // @[Modules.scala 71:109:@9162.4]
  wire [10:0] buffer_3_695; // @[Modules.scala 71:109:@9163.4]
  wire [11:0] _T_60980; // @[Modules.scala 71:109:@9165.4]
  wire [10:0] _T_60981; // @[Modules.scala 71:109:@9166.4]
  wire [10:0] buffer_3_696; // @[Modules.scala 71:109:@9167.4]
  wire [11:0] _T_60983; // @[Modules.scala 71:109:@9169.4]
  wire [10:0] _T_60984; // @[Modules.scala 71:109:@9170.4]
  wire [10:0] buffer_3_697; // @[Modules.scala 71:109:@9171.4]
  wire [11:0] _T_60986; // @[Modules.scala 71:109:@9173.4]
  wire [10:0] _T_60987; // @[Modules.scala 71:109:@9174.4]
  wire [10:0] buffer_3_698; // @[Modules.scala 71:109:@9175.4]
  wire [11:0] _T_60989; // @[Modules.scala 71:109:@9177.4]
  wire [10:0] _T_60990; // @[Modules.scala 71:109:@9178.4]
  wire [10:0] buffer_3_699; // @[Modules.scala 71:109:@9179.4]
  wire [11:0] _T_60992; // @[Modules.scala 71:109:@9181.4]
  wire [10:0] _T_60993; // @[Modules.scala 71:109:@9182.4]
  wire [10:0] buffer_3_700; // @[Modules.scala 71:109:@9183.4]
  wire [11:0] _T_60995; // @[Modules.scala 71:109:@9185.4]
  wire [10:0] _T_60996; // @[Modules.scala 71:109:@9186.4]
  wire [10:0] buffer_3_701; // @[Modules.scala 71:109:@9187.4]
  wire [11:0] _T_60998; // @[Modules.scala 71:109:@9189.4]
  wire [10:0] _T_60999; // @[Modules.scala 71:109:@9190.4]
  wire [10:0] buffer_3_702; // @[Modules.scala 71:109:@9191.4]
  wire [11:0] _T_61001; // @[Modules.scala 71:109:@9193.4]
  wire [10:0] _T_61002; // @[Modules.scala 71:109:@9194.4]
  wire [10:0] buffer_3_703; // @[Modules.scala 71:109:@9195.4]
  wire [11:0] _T_61004; // @[Modules.scala 71:109:@9197.4]
  wire [10:0] _T_61005; // @[Modules.scala 71:109:@9198.4]
  wire [10:0] buffer_3_704; // @[Modules.scala 71:109:@9199.4]
  wire [11:0] _T_61007; // @[Modules.scala 71:109:@9201.4]
  wire [10:0] _T_61008; // @[Modules.scala 71:109:@9202.4]
  wire [10:0] buffer_3_705; // @[Modules.scala 71:109:@9203.4]
  wire [11:0] _T_61010; // @[Modules.scala 71:109:@9205.4]
  wire [10:0] _T_61011; // @[Modules.scala 71:109:@9206.4]
  wire [10:0] buffer_3_706; // @[Modules.scala 71:109:@9207.4]
  wire [11:0] _T_61013; // @[Modules.scala 71:109:@9209.4]
  wire [10:0] _T_61014; // @[Modules.scala 71:109:@9210.4]
  wire [10:0] buffer_3_707; // @[Modules.scala 71:109:@9211.4]
  wire [11:0] _T_61016; // @[Modules.scala 71:109:@9213.4]
  wire [10:0] _T_61017; // @[Modules.scala 71:109:@9214.4]
  wire [10:0] buffer_3_708; // @[Modules.scala 71:109:@9215.4]
  wire [11:0] _T_61019; // @[Modules.scala 71:109:@9217.4]
  wire [10:0] _T_61020; // @[Modules.scala 71:109:@9218.4]
  wire [10:0] buffer_3_709; // @[Modules.scala 71:109:@9219.4]
  wire [11:0] _T_61022; // @[Modules.scala 71:109:@9221.4]
  wire [10:0] _T_61023; // @[Modules.scala 71:109:@9222.4]
  wire [10:0] buffer_3_710; // @[Modules.scala 71:109:@9223.4]
  wire [11:0] _T_61025; // @[Modules.scala 71:109:@9225.4]
  wire [10:0] _T_61026; // @[Modules.scala 71:109:@9226.4]
  wire [10:0] buffer_3_711; // @[Modules.scala 71:109:@9227.4]
  wire [11:0] _T_61028; // @[Modules.scala 71:109:@9229.4]
  wire [10:0] _T_61029; // @[Modules.scala 71:109:@9230.4]
  wire [10:0] buffer_3_712; // @[Modules.scala 71:109:@9231.4]
  wire [11:0] _T_61031; // @[Modules.scala 71:109:@9233.4]
  wire [10:0] _T_61032; // @[Modules.scala 71:109:@9234.4]
  wire [10:0] buffer_3_713; // @[Modules.scala 71:109:@9235.4]
  wire [11:0] _T_61034; // @[Modules.scala 71:109:@9237.4]
  wire [10:0] _T_61035; // @[Modules.scala 71:109:@9238.4]
  wire [10:0] buffer_3_714; // @[Modules.scala 71:109:@9239.4]
  wire [11:0] _T_61037; // @[Modules.scala 71:109:@9241.4]
  wire [10:0] _T_61038; // @[Modules.scala 71:109:@9242.4]
  wire [10:0] buffer_3_715; // @[Modules.scala 71:109:@9243.4]
  wire [11:0] _T_61040; // @[Modules.scala 71:109:@9245.4]
  wire [10:0] _T_61041; // @[Modules.scala 71:109:@9246.4]
  wire [10:0] buffer_3_716; // @[Modules.scala 71:109:@9247.4]
  wire [11:0] _T_61043; // @[Modules.scala 71:109:@9249.4]
  wire [10:0] _T_61044; // @[Modules.scala 71:109:@9250.4]
  wire [10:0] buffer_3_717; // @[Modules.scala 71:109:@9251.4]
  wire [11:0] _T_61046; // @[Modules.scala 71:109:@9253.4]
  wire [10:0] _T_61047; // @[Modules.scala 71:109:@9254.4]
  wire [10:0] buffer_3_718; // @[Modules.scala 71:109:@9255.4]
  wire [11:0] _T_61049; // @[Modules.scala 71:109:@9257.4]
  wire [10:0] _T_61050; // @[Modules.scala 71:109:@9258.4]
  wire [10:0] buffer_3_719; // @[Modules.scala 71:109:@9259.4]
  wire [11:0] _T_61052; // @[Modules.scala 71:109:@9261.4]
  wire [10:0] _T_61053; // @[Modules.scala 71:109:@9262.4]
  wire [10:0] buffer_3_720; // @[Modules.scala 71:109:@9263.4]
  wire [11:0] _T_61055; // @[Modules.scala 71:109:@9265.4]
  wire [10:0] _T_61056; // @[Modules.scala 71:109:@9266.4]
  wire [10:0] buffer_3_721; // @[Modules.scala 71:109:@9267.4]
  wire [11:0] _T_61058; // @[Modules.scala 71:109:@9269.4]
  wire [10:0] _T_61059; // @[Modules.scala 71:109:@9270.4]
  wire [10:0] buffer_3_722; // @[Modules.scala 71:109:@9271.4]
  wire [11:0] _T_61061; // @[Modules.scala 71:109:@9273.4]
  wire [10:0] _T_61062; // @[Modules.scala 71:109:@9274.4]
  wire [10:0] buffer_3_723; // @[Modules.scala 71:109:@9275.4]
  wire [11:0] _T_61064; // @[Modules.scala 71:109:@9277.4]
  wire [10:0] _T_61065; // @[Modules.scala 71:109:@9278.4]
  wire [10:0] buffer_3_724; // @[Modules.scala 71:109:@9279.4]
  wire [11:0] _T_61067; // @[Modules.scala 71:109:@9281.4]
  wire [10:0] _T_61068; // @[Modules.scala 71:109:@9282.4]
  wire [10:0] buffer_3_725; // @[Modules.scala 71:109:@9283.4]
  wire [11:0] _T_61070; // @[Modules.scala 71:109:@9285.4]
  wire [10:0] _T_61071; // @[Modules.scala 71:109:@9286.4]
  wire [10:0] buffer_3_726; // @[Modules.scala 71:109:@9287.4]
  wire [11:0] _T_61073; // @[Modules.scala 71:109:@9289.4]
  wire [10:0] _T_61074; // @[Modules.scala 71:109:@9290.4]
  wire [10:0] buffer_3_727; // @[Modules.scala 71:109:@9291.4]
  wire [11:0] _T_61076; // @[Modules.scala 71:109:@9293.4]
  wire [10:0] _T_61077; // @[Modules.scala 71:109:@9294.4]
  wire [10:0] buffer_3_728; // @[Modules.scala 71:109:@9295.4]
  wire [11:0] _T_61079; // @[Modules.scala 71:109:@9297.4]
  wire [10:0] _T_61080; // @[Modules.scala 71:109:@9298.4]
  wire [10:0] buffer_3_729; // @[Modules.scala 71:109:@9299.4]
  wire [11:0] _T_61082; // @[Modules.scala 71:109:@9301.4]
  wire [10:0] _T_61083; // @[Modules.scala 71:109:@9302.4]
  wire [10:0] buffer_3_730; // @[Modules.scala 71:109:@9303.4]
  wire [11:0] _T_61085; // @[Modules.scala 71:109:@9305.4]
  wire [10:0] _T_61086; // @[Modules.scala 71:109:@9306.4]
  wire [10:0] buffer_3_731; // @[Modules.scala 71:109:@9307.4]
  wire [11:0] _T_61088; // @[Modules.scala 71:109:@9309.4]
  wire [10:0] _T_61089; // @[Modules.scala 71:109:@9310.4]
  wire [10:0] buffer_3_732; // @[Modules.scala 71:109:@9311.4]
  wire [11:0] _T_61091; // @[Modules.scala 71:109:@9313.4]
  wire [10:0] _T_61092; // @[Modules.scala 71:109:@9314.4]
  wire [10:0] buffer_3_733; // @[Modules.scala 71:109:@9315.4]
  wire [11:0] _T_61094; // @[Modules.scala 71:109:@9317.4]
  wire [10:0] _T_61095; // @[Modules.scala 71:109:@9318.4]
  wire [10:0] buffer_3_734; // @[Modules.scala 71:109:@9319.4]
  wire [11:0] _T_61097; // @[Modules.scala 78:156:@9322.4]
  wire [10:0] _T_61098; // @[Modules.scala 78:156:@9323.4]
  wire [10:0] buffer_3_736; // @[Modules.scala 78:156:@9324.4]
  wire [11:0] _T_61100; // @[Modules.scala 78:156:@9326.4]
  wire [10:0] _T_61101; // @[Modules.scala 78:156:@9327.4]
  wire [10:0] buffer_3_737; // @[Modules.scala 78:156:@9328.4]
  wire [11:0] _T_61103; // @[Modules.scala 78:156:@9330.4]
  wire [10:0] _T_61104; // @[Modules.scala 78:156:@9331.4]
  wire [10:0] buffer_3_738; // @[Modules.scala 78:156:@9332.4]
  wire [11:0] _T_61106; // @[Modules.scala 78:156:@9334.4]
  wire [10:0] _T_61107; // @[Modules.scala 78:156:@9335.4]
  wire [10:0] buffer_3_739; // @[Modules.scala 78:156:@9336.4]
  wire [11:0] _T_61109; // @[Modules.scala 78:156:@9338.4]
  wire [10:0] _T_61110; // @[Modules.scala 78:156:@9339.4]
  wire [10:0] buffer_3_740; // @[Modules.scala 78:156:@9340.4]
  wire [11:0] _T_61112; // @[Modules.scala 78:156:@9342.4]
  wire [10:0] _T_61113; // @[Modules.scala 78:156:@9343.4]
  wire [10:0] buffer_3_741; // @[Modules.scala 78:156:@9344.4]
  wire [11:0] _T_61115; // @[Modules.scala 78:156:@9346.4]
  wire [10:0] _T_61116; // @[Modules.scala 78:156:@9347.4]
  wire [10:0] buffer_3_742; // @[Modules.scala 78:156:@9348.4]
  wire [11:0] _T_61118; // @[Modules.scala 78:156:@9350.4]
  wire [10:0] _T_61119; // @[Modules.scala 78:156:@9351.4]
  wire [10:0] buffer_3_743; // @[Modules.scala 78:156:@9352.4]
  wire [11:0] _T_61121; // @[Modules.scala 78:156:@9354.4]
  wire [10:0] _T_61122; // @[Modules.scala 78:156:@9355.4]
  wire [10:0] buffer_3_744; // @[Modules.scala 78:156:@9356.4]
  wire [11:0] _T_61124; // @[Modules.scala 78:156:@9358.4]
  wire [10:0] _T_61125; // @[Modules.scala 78:156:@9359.4]
  wire [10:0] buffer_3_745; // @[Modules.scala 78:156:@9360.4]
  wire [11:0] _T_61127; // @[Modules.scala 78:156:@9362.4]
  wire [10:0] _T_61128; // @[Modules.scala 78:156:@9363.4]
  wire [10:0] buffer_3_746; // @[Modules.scala 78:156:@9364.4]
  wire [11:0] _T_61130; // @[Modules.scala 78:156:@9366.4]
  wire [10:0] _T_61131; // @[Modules.scala 78:156:@9367.4]
  wire [10:0] buffer_3_747; // @[Modules.scala 78:156:@9368.4]
  wire [11:0] _T_61133; // @[Modules.scala 78:156:@9370.4]
  wire [10:0] _T_61134; // @[Modules.scala 78:156:@9371.4]
  wire [10:0] buffer_3_748; // @[Modules.scala 78:156:@9372.4]
  wire [11:0] _T_61136; // @[Modules.scala 78:156:@9374.4]
  wire [10:0] _T_61137; // @[Modules.scala 78:156:@9375.4]
  wire [10:0] buffer_3_749; // @[Modules.scala 78:156:@9376.4]
  wire [11:0] _T_61139; // @[Modules.scala 78:156:@9378.4]
  wire [10:0] _T_61140; // @[Modules.scala 78:156:@9379.4]
  wire [10:0] buffer_3_750; // @[Modules.scala 78:156:@9380.4]
  wire [11:0] _T_61142; // @[Modules.scala 78:156:@9382.4]
  wire [10:0] _T_61143; // @[Modules.scala 78:156:@9383.4]
  wire [10:0] buffer_3_751; // @[Modules.scala 78:156:@9384.4]
  wire [11:0] _T_61145; // @[Modules.scala 78:156:@9386.4]
  wire [10:0] _T_61146; // @[Modules.scala 78:156:@9387.4]
  wire [10:0] buffer_3_752; // @[Modules.scala 78:156:@9388.4]
  wire [11:0] _T_61148; // @[Modules.scala 78:156:@9390.4]
  wire [10:0] _T_61149; // @[Modules.scala 78:156:@9391.4]
  wire [10:0] buffer_3_753; // @[Modules.scala 78:156:@9392.4]
  wire [11:0] _T_61151; // @[Modules.scala 78:156:@9394.4]
  wire [10:0] _T_61152; // @[Modules.scala 78:156:@9395.4]
  wire [10:0] buffer_3_754; // @[Modules.scala 78:156:@9396.4]
  wire [11:0] _T_61154; // @[Modules.scala 78:156:@9398.4]
  wire [10:0] _T_61155; // @[Modules.scala 78:156:@9399.4]
  wire [10:0] buffer_3_755; // @[Modules.scala 78:156:@9400.4]
  wire [11:0] _T_61157; // @[Modules.scala 78:156:@9402.4]
  wire [10:0] _T_61158; // @[Modules.scala 78:156:@9403.4]
  wire [10:0] buffer_3_756; // @[Modules.scala 78:156:@9404.4]
  wire [11:0] _T_61160; // @[Modules.scala 78:156:@9406.4]
  wire [10:0] _T_61161; // @[Modules.scala 78:156:@9407.4]
  wire [10:0] buffer_3_757; // @[Modules.scala 78:156:@9408.4]
  wire [11:0] _T_61163; // @[Modules.scala 78:156:@9410.4]
  wire [10:0] _T_61164; // @[Modules.scala 78:156:@9411.4]
  wire [10:0] buffer_3_758; // @[Modules.scala 78:156:@9412.4]
  wire [11:0] _T_61166; // @[Modules.scala 78:156:@9414.4]
  wire [10:0] _T_61167; // @[Modules.scala 78:156:@9415.4]
  wire [10:0] buffer_3_759; // @[Modules.scala 78:156:@9416.4]
  wire [11:0] _T_61169; // @[Modules.scala 78:156:@9418.4]
  wire [10:0] _T_61170; // @[Modules.scala 78:156:@9419.4]
  wire [10:0] buffer_3_760; // @[Modules.scala 78:156:@9420.4]
  wire [11:0] _T_61172; // @[Modules.scala 78:156:@9422.4]
  wire [10:0] _T_61173; // @[Modules.scala 78:156:@9423.4]
  wire [10:0] buffer_3_761; // @[Modules.scala 78:156:@9424.4]
  wire [11:0] _T_61175; // @[Modules.scala 78:156:@9426.4]
  wire [10:0] _T_61176; // @[Modules.scala 78:156:@9427.4]
  wire [10:0] buffer_3_762; // @[Modules.scala 78:156:@9428.4]
  wire [11:0] _T_61178; // @[Modules.scala 78:156:@9430.4]
  wire [10:0] _T_61179; // @[Modules.scala 78:156:@9431.4]
  wire [10:0] buffer_3_763; // @[Modules.scala 78:156:@9432.4]
  wire [11:0] _T_61181; // @[Modules.scala 78:156:@9434.4]
  wire [10:0] _T_61182; // @[Modules.scala 78:156:@9435.4]
  wire [10:0] buffer_3_764; // @[Modules.scala 78:156:@9436.4]
  wire [11:0] _T_61184; // @[Modules.scala 78:156:@9438.4]
  wire [10:0] _T_61185; // @[Modules.scala 78:156:@9439.4]
  wire [10:0] buffer_3_765; // @[Modules.scala 78:156:@9440.4]
  wire [11:0] _T_61187; // @[Modules.scala 78:156:@9442.4]
  wire [10:0] _T_61188; // @[Modules.scala 78:156:@9443.4]
  wire [10:0] buffer_3_766; // @[Modules.scala 78:156:@9444.4]
  wire [11:0] _T_61190; // @[Modules.scala 78:156:@9446.4]
  wire [10:0] _T_61191; // @[Modules.scala 78:156:@9447.4]
  wire [10:0] buffer_3_767; // @[Modules.scala 78:156:@9448.4]
  wire [11:0] _T_61193; // @[Modules.scala 78:156:@9450.4]
  wire [10:0] _T_61194; // @[Modules.scala 78:156:@9451.4]
  wire [10:0] buffer_3_768; // @[Modules.scala 78:156:@9452.4]
  wire [11:0] _T_61196; // @[Modules.scala 78:156:@9454.4]
  wire [10:0] _T_61197; // @[Modules.scala 78:156:@9455.4]
  wire [10:0] buffer_3_769; // @[Modules.scala 78:156:@9456.4]
  wire [11:0] _T_61199; // @[Modules.scala 78:156:@9458.4]
  wire [10:0] _T_61200; // @[Modules.scala 78:156:@9459.4]
  wire [10:0] buffer_3_770; // @[Modules.scala 78:156:@9460.4]
  wire [11:0] _T_61202; // @[Modules.scala 78:156:@9462.4]
  wire [10:0] _T_61203; // @[Modules.scala 78:156:@9463.4]
  wire [10:0] buffer_3_771; // @[Modules.scala 78:156:@9464.4]
  wire [11:0] _T_61205; // @[Modules.scala 78:156:@9466.4]
  wire [10:0] _T_61206; // @[Modules.scala 78:156:@9467.4]
  wire [10:0] buffer_3_772; // @[Modules.scala 78:156:@9468.4]
  wire [11:0] _T_61208; // @[Modules.scala 78:156:@9470.4]
  wire [10:0] _T_61209; // @[Modules.scala 78:156:@9471.4]
  wire [10:0] buffer_3_773; // @[Modules.scala 78:156:@9472.4]
  wire [11:0] _T_61211; // @[Modules.scala 78:156:@9474.4]
  wire [10:0] _T_61212; // @[Modules.scala 78:156:@9475.4]
  wire [10:0] buffer_3_774; // @[Modules.scala 78:156:@9476.4]
  wire [11:0] _T_61214; // @[Modules.scala 78:156:@9478.4]
  wire [10:0] _T_61215; // @[Modules.scala 78:156:@9479.4]
  wire [10:0] buffer_3_775; // @[Modules.scala 78:156:@9480.4]
  wire [11:0] _T_61217; // @[Modules.scala 78:156:@9482.4]
  wire [10:0] _T_61218; // @[Modules.scala 78:156:@9483.4]
  wire [10:0] buffer_3_776; // @[Modules.scala 78:156:@9484.4]
  wire [11:0] _T_61220; // @[Modules.scala 78:156:@9486.4]
  wire [10:0] _T_61221; // @[Modules.scala 78:156:@9487.4]
  wire [10:0] buffer_3_777; // @[Modules.scala 78:156:@9488.4]
  wire [11:0] _T_61223; // @[Modules.scala 78:156:@9490.4]
  wire [10:0] _T_61224; // @[Modules.scala 78:156:@9491.4]
  wire [10:0] buffer_3_778; // @[Modules.scala 78:156:@9492.4]
  wire [11:0] _T_61226; // @[Modules.scala 78:156:@9494.4]
  wire [10:0] _T_61227; // @[Modules.scala 78:156:@9495.4]
  wire [10:0] buffer_3_779; // @[Modules.scala 78:156:@9496.4]
  wire [11:0] _T_61229; // @[Modules.scala 78:156:@9498.4]
  wire [10:0] _T_61230; // @[Modules.scala 78:156:@9499.4]
  wire [10:0] buffer_3_780; // @[Modules.scala 78:156:@9500.4]
  wire [11:0] _T_61232; // @[Modules.scala 78:156:@9502.4]
  wire [10:0] _T_61233; // @[Modules.scala 78:156:@9503.4]
  wire [10:0] buffer_3_781; // @[Modules.scala 78:156:@9504.4]
  wire [11:0] _T_61235; // @[Modules.scala 78:156:@9506.4]
  wire [10:0] _T_61236; // @[Modules.scala 78:156:@9507.4]
  wire [10:0] buffer_3_782; // @[Modules.scala 78:156:@9508.4]
  wire [11:0] _T_61238; // @[Modules.scala 78:156:@9510.4]
  wire [10:0] _T_61239; // @[Modules.scala 78:156:@9511.4]
  wire [10:0] buffer_3_783; // @[Modules.scala 78:156:@9512.4]
  wire [5:0] _T_61268; // @[Modules.scala 37:46:@9558.4]
  wire [4:0] _T_61269; // @[Modules.scala 37:46:@9559.4]
  wire [4:0] _T_61270; // @[Modules.scala 37:46:@9560.4]
  wire [5:0] _T_61361; // @[Modules.scala 37:46:@9686.4]
  wire [4:0] _T_61362; // @[Modules.scala 37:46:@9687.4]
  wire [4:0] _T_61363; // @[Modules.scala 37:46:@9688.4]
  wire [5:0] _T_61365; // @[Modules.scala 37:46:@9692.4]
  wire [4:0] _T_61366; // @[Modules.scala 37:46:@9693.4]
  wire [4:0] _T_61367; // @[Modules.scala 37:46:@9694.4]
  wire [5:0] _T_61377; // @[Modules.scala 37:46:@9708.4]
  wire [4:0] _T_61378; // @[Modules.scala 37:46:@9709.4]
  wire [4:0] _T_61379; // @[Modules.scala 37:46:@9710.4]
  wire [5:0] _T_61383; // @[Modules.scala 37:46:@9716.4]
  wire [4:0] _T_61384; // @[Modules.scala 37:46:@9717.4]
  wire [4:0] _T_61385; // @[Modules.scala 37:46:@9718.4]
  wire [5:0] _T_61395; // @[Modules.scala 37:46:@9734.4]
  wire [4:0] _T_61396; // @[Modules.scala 37:46:@9735.4]
  wire [4:0] _T_61397; // @[Modules.scala 37:46:@9736.4]
  wire [5:0] _T_61413; // @[Modules.scala 37:46:@9759.4]
  wire [4:0] _T_61414; // @[Modules.scala 37:46:@9760.4]
  wire [4:0] _T_61415; // @[Modules.scala 37:46:@9761.4]
  wire [5:0] _T_61447; // @[Modules.scala 37:46:@9808.4]
  wire [4:0] _T_61448; // @[Modules.scala 37:46:@9809.4]
  wire [4:0] _T_61449; // @[Modules.scala 37:46:@9810.4]
  wire [5:0] _T_61456; // @[Modules.scala 37:46:@9820.4]
  wire [4:0] _T_61457; // @[Modules.scala 37:46:@9821.4]
  wire [4:0] _T_61458; // @[Modules.scala 37:46:@9822.4]
  wire [5:0] _T_61470; // @[Modules.scala 37:46:@9839.4]
  wire [4:0] _T_61471; // @[Modules.scala 37:46:@9840.4]
  wire [4:0] _T_61472; // @[Modules.scala 37:46:@9841.4]
  wire [5:0] _T_61473; // @[Modules.scala 37:46:@9843.4]
  wire [4:0] _T_61474; // @[Modules.scala 37:46:@9844.4]
  wire [4:0] _T_61475; // @[Modules.scala 37:46:@9845.4]
  wire [5:0] _T_61496; // @[Modules.scala 37:46:@9877.4]
  wire [4:0] _T_61497; // @[Modules.scala 37:46:@9878.4]
  wire [4:0] _T_61498; // @[Modules.scala 37:46:@9879.4]
  wire [5:0] _T_61500; // @[Modules.scala 37:46:@9882.4]
  wire [4:0] _T_61501; // @[Modules.scala 37:46:@9883.4]
  wire [4:0] _T_61502; // @[Modules.scala 37:46:@9884.4]
  wire [5:0] _T_61554; // @[Modules.scala 37:46:@9961.4]
  wire [4:0] _T_61555; // @[Modules.scala 37:46:@9962.4]
  wire [4:0] _T_61556; // @[Modules.scala 37:46:@9963.4]
  wire [5:0] _T_61570; // @[Modules.scala 37:46:@9990.4]
  wire [4:0] _T_61571; // @[Modules.scala 37:46:@9991.4]
  wire [4:0] _T_61572; // @[Modules.scala 37:46:@9992.4]
  wire [5:0] _T_61573; // @[Modules.scala 37:46:@9995.4]
  wire [4:0] _T_61574; // @[Modules.scala 37:46:@9996.4]
  wire [4:0] _T_61575; // @[Modules.scala 37:46:@9997.4]
  wire [5:0] _T_61635; // @[Modules.scala 37:46:@10091.4]
  wire [4:0] _T_61636; // @[Modules.scala 37:46:@10092.4]
  wire [4:0] _T_61637; // @[Modules.scala 37:46:@10093.4]
  wire [5:0] _T_61686; // @[Modules.scala 37:46:@10166.4]
  wire [4:0] _T_61687; // @[Modules.scala 37:46:@10167.4]
  wire [4:0] _T_61688; // @[Modules.scala 37:46:@10168.4]
  wire [5:0] _T_61729; // @[Modules.scala 37:46:@10225.4]
  wire [4:0] _T_61730; // @[Modules.scala 37:46:@10226.4]
  wire [4:0] _T_61731; // @[Modules.scala 37:46:@10227.4]
  wire [5:0] _T_61766; // @[Modules.scala 37:46:@10278.4]
  wire [4:0] _T_61767; // @[Modules.scala 37:46:@10279.4]
  wire [4:0] _T_61768; // @[Modules.scala 37:46:@10280.4]
  wire [5:0] _T_61775; // @[Modules.scala 37:46:@10291.4]
  wire [4:0] _T_61776; // @[Modules.scala 37:46:@10292.4]
  wire [4:0] _T_61777; // @[Modules.scala 37:46:@10293.4]
  wire [5:0] _T_61821; // @[Modules.scala 37:46:@10358.4]
  wire [4:0] _T_61822; // @[Modules.scala 37:46:@10359.4]
  wire [4:0] _T_61823; // @[Modules.scala 37:46:@10360.4]
  wire [5:0] _T_61861; // @[Modules.scala 37:46:@10412.4]
  wire [4:0] _T_61862; // @[Modules.scala 37:46:@10413.4]
  wire [4:0] _T_61863; // @[Modules.scala 37:46:@10414.4]
  wire [10:0] buffer_4_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61887; // @[Modules.scala 65:57:@10450.4]
  wire [10:0] _T_61888; // @[Modules.scala 65:57:@10451.4]
  wire [10:0] buffer_4_392; // @[Modules.scala 65:57:@10452.4]
  wire [11:0] _T_61890; // @[Modules.scala 65:57:@10454.4]
  wire [10:0] _T_61891; // @[Modules.scala 65:57:@10455.4]
  wire [10:0] buffer_4_393; // @[Modules.scala 65:57:@10456.4]
  wire [10:0] buffer_4_5; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61893; // @[Modules.scala 65:57:@10458.4]
  wire [10:0] _T_61894; // @[Modules.scala 65:57:@10459.4]
  wire [10:0] buffer_4_394; // @[Modules.scala 65:57:@10460.4]
  wire [11:0] _T_61896; // @[Modules.scala 65:57:@10462.4]
  wire [10:0] _T_61897; // @[Modules.scala 65:57:@10463.4]
  wire [10:0] buffer_4_395; // @[Modules.scala 65:57:@10464.4]
  wire [11:0] _T_61899; // @[Modules.scala 65:57:@10466.4]
  wire [10:0] _T_61900; // @[Modules.scala 65:57:@10467.4]
  wire [10:0] buffer_4_396; // @[Modules.scala 65:57:@10468.4]
  wire [11:0] _T_61902; // @[Modules.scala 65:57:@10470.4]
  wire [10:0] _T_61903; // @[Modules.scala 65:57:@10471.4]
  wire [10:0] buffer_4_397; // @[Modules.scala 65:57:@10472.4]
  wire [10:0] buffer_4_13; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61905; // @[Modules.scala 65:57:@10474.4]
  wire [10:0] _T_61906; // @[Modules.scala 65:57:@10475.4]
  wire [10:0] buffer_4_398; // @[Modules.scala 65:57:@10476.4]
  wire [10:0] buffer_4_14; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61908; // @[Modules.scala 65:57:@10478.4]
  wire [10:0] _T_61909; // @[Modules.scala 65:57:@10479.4]
  wire [10:0] buffer_4_399; // @[Modules.scala 65:57:@10480.4]
  wire [11:0] _T_61917; // @[Modules.scala 65:57:@10490.4]
  wire [10:0] _T_61918; // @[Modules.scala 65:57:@10491.4]
  wire [10:0] buffer_4_402; // @[Modules.scala 65:57:@10492.4]
  wire [10:0] buffer_4_22; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61920; // @[Modules.scala 65:57:@10494.4]
  wire [10:0] _T_61921; // @[Modules.scala 65:57:@10495.4]
  wire [10:0] buffer_4_403; // @[Modules.scala 65:57:@10496.4]
  wire [11:0] _T_61926; // @[Modules.scala 65:57:@10502.4]
  wire [10:0] _T_61927; // @[Modules.scala 65:57:@10503.4]
  wire [10:0] buffer_4_405; // @[Modules.scala 65:57:@10504.4]
  wire [11:0] _T_61950; // @[Modules.scala 65:57:@10534.4]
  wire [10:0] _T_61951; // @[Modules.scala 65:57:@10535.4]
  wire [10:0] buffer_4_413; // @[Modules.scala 65:57:@10536.4]
  wire [10:0] buffer_4_44; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61953; // @[Modules.scala 65:57:@10538.4]
  wire [10:0] _T_61954; // @[Modules.scala 65:57:@10539.4]
  wire [10:0] buffer_4_414; // @[Modules.scala 65:57:@10540.4]
  wire [10:0] buffer_4_58; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_59; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61974; // @[Modules.scala 65:57:@10566.4]
  wire [10:0] _T_61975; // @[Modules.scala 65:57:@10567.4]
  wire [10:0] buffer_4_421; // @[Modules.scala 65:57:@10568.4]
  wire [10:0] buffer_4_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61977; // @[Modules.scala 65:57:@10570.4]
  wire [10:0] _T_61978; // @[Modules.scala 65:57:@10571.4]
  wire [10:0] buffer_4_422; // @[Modules.scala 65:57:@10572.4]
  wire [11:0] _T_61980; // @[Modules.scala 65:57:@10574.4]
  wire [10:0] _T_61981; // @[Modules.scala 65:57:@10575.4]
  wire [10:0] buffer_4_423; // @[Modules.scala 65:57:@10576.4]
  wire [10:0] buffer_4_64; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61983; // @[Modules.scala 65:57:@10578.4]
  wire [10:0] _T_61984; // @[Modules.scala 65:57:@10579.4]
  wire [10:0] buffer_4_424; // @[Modules.scala 65:57:@10580.4]
  wire [10:0] buffer_4_69; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61989; // @[Modules.scala 65:57:@10586.4]
  wire [10:0] _T_61990; // @[Modules.scala 65:57:@10587.4]
  wire [10:0] buffer_4_426; // @[Modules.scala 65:57:@10588.4]
  wire [11:0] _T_61992; // @[Modules.scala 65:57:@10590.4]
  wire [10:0] _T_61993; // @[Modules.scala 65:57:@10591.4]
  wire [10:0] buffer_4_427; // @[Modules.scala 65:57:@10592.4]
  wire [10:0] buffer_4_72; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_61995; // @[Modules.scala 65:57:@10594.4]
  wire [10:0] _T_61996; // @[Modules.scala 65:57:@10595.4]
  wire [10:0] buffer_4_428; // @[Modules.scala 65:57:@10596.4]
  wire [10:0] buffer_4_76; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62001; // @[Modules.scala 65:57:@10602.4]
  wire [10:0] _T_62002; // @[Modules.scala 65:57:@10603.4]
  wire [10:0] buffer_4_430; // @[Modules.scala 65:57:@10604.4]
  wire [10:0] buffer_4_78; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62004; // @[Modules.scala 65:57:@10606.4]
  wire [10:0] _T_62005; // @[Modules.scala 65:57:@10607.4]
  wire [10:0] buffer_4_431; // @[Modules.scala 65:57:@10608.4]
  wire [10:0] buffer_4_80; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62007; // @[Modules.scala 65:57:@10610.4]
  wire [10:0] _T_62008; // @[Modules.scala 65:57:@10611.4]
  wire [10:0] buffer_4_432; // @[Modules.scala 65:57:@10612.4]
  wire [10:0] buffer_4_84; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62013; // @[Modules.scala 65:57:@10618.4]
  wire [10:0] _T_62014; // @[Modules.scala 65:57:@10619.4]
  wire [10:0] buffer_4_434; // @[Modules.scala 65:57:@10620.4]
  wire [10:0] buffer_4_92; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62025; // @[Modules.scala 65:57:@10634.4]
  wire [10:0] _T_62026; // @[Modules.scala 65:57:@10635.4]
  wire [10:0] buffer_4_438; // @[Modules.scala 65:57:@10636.4]
  wire [10:0] buffer_4_94; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62028; // @[Modules.scala 65:57:@10638.4]
  wire [10:0] _T_62029; // @[Modules.scala 65:57:@10639.4]
  wire [10:0] buffer_4_439; // @[Modules.scala 65:57:@10640.4]
  wire [11:0] _T_62034; // @[Modules.scala 65:57:@10646.4]
  wire [10:0] _T_62035; // @[Modules.scala 65:57:@10647.4]
  wire [10:0] buffer_4_441; // @[Modules.scala 65:57:@10648.4]
  wire [10:0] buffer_4_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62037; // @[Modules.scala 65:57:@10650.4]
  wire [10:0] _T_62038; // @[Modules.scala 65:57:@10651.4]
  wire [10:0] buffer_4_442; // @[Modules.scala 65:57:@10652.4]
  wire [10:0] buffer_4_102; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62040; // @[Modules.scala 65:57:@10654.4]
  wire [10:0] _T_62041; // @[Modules.scala 65:57:@10655.4]
  wire [10:0] buffer_4_443; // @[Modules.scala 65:57:@10656.4]
  wire [10:0] buffer_4_114; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62058; // @[Modules.scala 65:57:@10678.4]
  wire [10:0] _T_62059; // @[Modules.scala 65:57:@10679.4]
  wire [10:0] buffer_4_449; // @[Modules.scala 65:57:@10680.4]
  wire [10:0] buffer_4_116; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62061; // @[Modules.scala 65:57:@10682.4]
  wire [10:0] _T_62062; // @[Modules.scala 65:57:@10683.4]
  wire [10:0] buffer_4_450; // @[Modules.scala 65:57:@10684.4]
  wire [10:0] buffer_4_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62067; // @[Modules.scala 65:57:@10690.4]
  wire [10:0] _T_62068; // @[Modules.scala 65:57:@10691.4]
  wire [10:0] buffer_4_452; // @[Modules.scala 65:57:@10692.4]
  wire [10:0] buffer_4_122; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62070; // @[Modules.scala 65:57:@10694.4]
  wire [10:0] _T_62071; // @[Modules.scala 65:57:@10695.4]
  wire [10:0] buffer_4_453; // @[Modules.scala 65:57:@10696.4]
  wire [10:0] buffer_4_128; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62079; // @[Modules.scala 65:57:@10706.4]
  wire [10:0] _T_62080; // @[Modules.scala 65:57:@10707.4]
  wire [10:0] buffer_4_456; // @[Modules.scala 65:57:@10708.4]
  wire [10:0] buffer_4_130; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62082; // @[Modules.scala 65:57:@10710.4]
  wire [10:0] _T_62083; // @[Modules.scala 65:57:@10711.4]
  wire [10:0] buffer_4_457; // @[Modules.scala 65:57:@10712.4]
  wire [11:0] _T_62097; // @[Modules.scala 65:57:@10730.4]
  wire [10:0] _T_62098; // @[Modules.scala 65:57:@10731.4]
  wire [10:0] buffer_4_462; // @[Modules.scala 65:57:@10732.4]
  wire [11:0] _T_62100; // @[Modules.scala 65:57:@10734.4]
  wire [10:0] _T_62101; // @[Modules.scala 65:57:@10735.4]
  wire [10:0] buffer_4_463; // @[Modules.scala 65:57:@10736.4]
  wire [10:0] buffer_4_148; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_149; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62109; // @[Modules.scala 65:57:@10746.4]
  wire [10:0] _T_62110; // @[Modules.scala 65:57:@10747.4]
  wire [10:0] buffer_4_466; // @[Modules.scala 65:57:@10748.4]
  wire [10:0] buffer_4_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62112; // @[Modules.scala 65:57:@10750.4]
  wire [10:0] _T_62113; // @[Modules.scala 65:57:@10751.4]
  wire [10:0] buffer_4_467; // @[Modules.scala 65:57:@10752.4]
  wire [10:0] buffer_4_154; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62118; // @[Modules.scala 65:57:@10758.4]
  wire [10:0] _T_62119; // @[Modules.scala 65:57:@10759.4]
  wire [10:0] buffer_4_469; // @[Modules.scala 65:57:@10760.4]
  wire [11:0] _T_62127; // @[Modules.scala 65:57:@10770.4]
  wire [10:0] _T_62128; // @[Modules.scala 65:57:@10771.4]
  wire [10:0] buffer_4_472; // @[Modules.scala 65:57:@10772.4]
  wire [11:0] _T_62136; // @[Modules.scala 65:57:@10782.4]
  wire [10:0] _T_62137; // @[Modules.scala 65:57:@10783.4]
  wire [10:0] buffer_4_475; // @[Modules.scala 65:57:@10784.4]
  wire [10:0] buffer_4_172; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62145; // @[Modules.scala 65:57:@10794.4]
  wire [10:0] _T_62146; // @[Modules.scala 65:57:@10795.4]
  wire [10:0] buffer_4_478; // @[Modules.scala 65:57:@10796.4]
  wire [10:0] buffer_4_176; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62151; // @[Modules.scala 65:57:@10802.4]
  wire [10:0] _T_62152; // @[Modules.scala 65:57:@10803.4]
  wire [10:0] buffer_4_480; // @[Modules.scala 65:57:@10804.4]
  wire [11:0] _T_62157; // @[Modules.scala 65:57:@10810.4]
  wire [10:0] _T_62158; // @[Modules.scala 65:57:@10811.4]
  wire [10:0] buffer_4_482; // @[Modules.scala 65:57:@10812.4]
  wire [10:0] buffer_4_182; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62160; // @[Modules.scala 65:57:@10814.4]
  wire [10:0] _T_62161; // @[Modules.scala 65:57:@10815.4]
  wire [10:0] buffer_4_483; // @[Modules.scala 65:57:@10816.4]
  wire [10:0] buffer_4_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62163; // @[Modules.scala 65:57:@10818.4]
  wire [10:0] _T_62164; // @[Modules.scala 65:57:@10819.4]
  wire [10:0] buffer_4_484; // @[Modules.scala 65:57:@10820.4]
  wire [10:0] buffer_4_190; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62172; // @[Modules.scala 65:57:@10830.4]
  wire [10:0] _T_62173; // @[Modules.scala 65:57:@10831.4]
  wire [10:0] buffer_4_487; // @[Modules.scala 65:57:@10832.4]
  wire [11:0] _T_62175; // @[Modules.scala 65:57:@10834.4]
  wire [10:0] _T_62176; // @[Modules.scala 65:57:@10835.4]
  wire [10:0] buffer_4_488; // @[Modules.scala 65:57:@10836.4]
  wire [10:0] buffer_4_194; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_195; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62178; // @[Modules.scala 65:57:@10838.4]
  wire [10:0] _T_62179; // @[Modules.scala 65:57:@10839.4]
  wire [10:0] buffer_4_489; // @[Modules.scala 65:57:@10840.4]
  wire [10:0] buffer_4_196; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62181; // @[Modules.scala 65:57:@10842.4]
  wire [10:0] _T_62182; // @[Modules.scala 65:57:@10843.4]
  wire [10:0] buffer_4_490; // @[Modules.scala 65:57:@10844.4]
  wire [10:0] buffer_4_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62184; // @[Modules.scala 65:57:@10846.4]
  wire [10:0] _T_62185; // @[Modules.scala 65:57:@10847.4]
  wire [10:0] buffer_4_491; // @[Modules.scala 65:57:@10848.4]
  wire [11:0] _T_62187; // @[Modules.scala 65:57:@10850.4]
  wire [10:0] _T_62188; // @[Modules.scala 65:57:@10851.4]
  wire [10:0] buffer_4_492; // @[Modules.scala 65:57:@10852.4]
  wire [10:0] buffer_4_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62190; // @[Modules.scala 65:57:@10854.4]
  wire [10:0] _T_62191; // @[Modules.scala 65:57:@10855.4]
  wire [10:0] buffer_4_493; // @[Modules.scala 65:57:@10856.4]
  wire [11:0] _T_62193; // @[Modules.scala 65:57:@10858.4]
  wire [10:0] _T_62194; // @[Modules.scala 65:57:@10859.4]
  wire [10:0] buffer_4_494; // @[Modules.scala 65:57:@10860.4]
  wire [10:0] buffer_4_206; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62196; // @[Modules.scala 65:57:@10862.4]
  wire [10:0] _T_62197; // @[Modules.scala 65:57:@10863.4]
  wire [10:0] buffer_4_495; // @[Modules.scala 65:57:@10864.4]
  wire [10:0] buffer_4_208; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_209; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62199; // @[Modules.scala 65:57:@10866.4]
  wire [10:0] _T_62200; // @[Modules.scala 65:57:@10867.4]
  wire [10:0] buffer_4_496; // @[Modules.scala 65:57:@10868.4]
  wire [10:0] buffer_4_210; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62202; // @[Modules.scala 65:57:@10870.4]
  wire [10:0] _T_62203; // @[Modules.scala 65:57:@10871.4]
  wire [10:0] buffer_4_497; // @[Modules.scala 65:57:@10872.4]
  wire [10:0] buffer_4_216; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62211; // @[Modules.scala 65:57:@10882.4]
  wire [10:0] _T_62212; // @[Modules.scala 65:57:@10883.4]
  wire [10:0] buffer_4_500; // @[Modules.scala 65:57:@10884.4]
  wire [10:0] buffer_4_218; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62214; // @[Modules.scala 65:57:@10886.4]
  wire [10:0] _T_62215; // @[Modules.scala 65:57:@10887.4]
  wire [10:0] buffer_4_501; // @[Modules.scala 65:57:@10888.4]
  wire [11:0] _T_62217; // @[Modules.scala 65:57:@10890.4]
  wire [10:0] _T_62218; // @[Modules.scala 65:57:@10891.4]
  wire [10:0] buffer_4_502; // @[Modules.scala 65:57:@10892.4]
  wire [10:0] buffer_4_227; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62226; // @[Modules.scala 65:57:@10902.4]
  wire [10:0] _T_62227; // @[Modules.scala 65:57:@10903.4]
  wire [10:0] buffer_4_505; // @[Modules.scala 65:57:@10904.4]
  wire [10:0] buffer_4_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62232; // @[Modules.scala 65:57:@10910.4]
  wire [10:0] _T_62233; // @[Modules.scala 65:57:@10911.4]
  wire [10:0] buffer_4_507; // @[Modules.scala 65:57:@10912.4]
  wire [11:0] _T_62235; // @[Modules.scala 65:57:@10914.4]
  wire [10:0] _T_62236; // @[Modules.scala 65:57:@10915.4]
  wire [10:0] buffer_4_508; // @[Modules.scala 65:57:@10916.4]
  wire [11:0] _T_62244; // @[Modules.scala 65:57:@10926.4]
  wire [10:0] _T_62245; // @[Modules.scala 65:57:@10927.4]
  wire [10:0] buffer_4_511; // @[Modules.scala 65:57:@10928.4]
  wire [11:0] _T_62247; // @[Modules.scala 65:57:@10930.4]
  wire [10:0] _T_62248; // @[Modules.scala 65:57:@10931.4]
  wire [10:0] buffer_4_512; // @[Modules.scala 65:57:@10932.4]
  wire [10:0] buffer_4_243; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62250; // @[Modules.scala 65:57:@10934.4]
  wire [10:0] _T_62251; // @[Modules.scala 65:57:@10935.4]
  wire [10:0] buffer_4_513; // @[Modules.scala 65:57:@10936.4]
  wire [10:0] buffer_4_246; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_247; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62256; // @[Modules.scala 65:57:@10942.4]
  wire [10:0] _T_62257; // @[Modules.scala 65:57:@10943.4]
  wire [10:0] buffer_4_515; // @[Modules.scala 65:57:@10944.4]
  wire [11:0] _T_62265; // @[Modules.scala 65:57:@10954.4]
  wire [10:0] _T_62266; // @[Modules.scala 65:57:@10955.4]
  wire [10:0] buffer_4_518; // @[Modules.scala 65:57:@10956.4]
  wire [10:0] buffer_4_256; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_257; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62271; // @[Modules.scala 65:57:@10962.4]
  wire [10:0] _T_62272; // @[Modules.scala 65:57:@10963.4]
  wire [10:0] buffer_4_520; // @[Modules.scala 65:57:@10964.4]
  wire [10:0] buffer_4_259; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62274; // @[Modules.scala 65:57:@10966.4]
  wire [10:0] _T_62275; // @[Modules.scala 65:57:@10967.4]
  wire [10:0] buffer_4_521; // @[Modules.scala 65:57:@10968.4]
  wire [10:0] buffer_4_260; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62277; // @[Modules.scala 65:57:@10970.4]
  wire [10:0] _T_62278; // @[Modules.scala 65:57:@10971.4]
  wire [10:0] buffer_4_522; // @[Modules.scala 65:57:@10972.4]
  wire [11:0] _T_62280; // @[Modules.scala 65:57:@10974.4]
  wire [10:0] _T_62281; // @[Modules.scala 65:57:@10975.4]
  wire [10:0] buffer_4_523; // @[Modules.scala 65:57:@10976.4]
  wire [11:0] _T_62286; // @[Modules.scala 65:57:@10982.4]
  wire [10:0] _T_62287; // @[Modules.scala 65:57:@10983.4]
  wire [10:0] buffer_4_525; // @[Modules.scala 65:57:@10984.4]
  wire [10:0] buffer_4_272; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_273; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62295; // @[Modules.scala 65:57:@10994.4]
  wire [10:0] _T_62296; // @[Modules.scala 65:57:@10995.4]
  wire [10:0] buffer_4_528; // @[Modules.scala 65:57:@10996.4]
  wire [11:0] _T_62304; // @[Modules.scala 65:57:@11006.4]
  wire [10:0] _T_62305; // @[Modules.scala 65:57:@11007.4]
  wire [10:0] buffer_4_531; // @[Modules.scala 65:57:@11008.4]
  wire [11:0] _T_62316; // @[Modules.scala 65:57:@11022.4]
  wire [10:0] _T_62317; // @[Modules.scala 65:57:@11023.4]
  wire [10:0] buffer_4_535; // @[Modules.scala 65:57:@11024.4]
  wire [10:0] buffer_4_290; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62322; // @[Modules.scala 65:57:@11030.4]
  wire [10:0] _T_62323; // @[Modules.scala 65:57:@11031.4]
  wire [10:0] buffer_4_537; // @[Modules.scala 65:57:@11032.4]
  wire [10:0] buffer_4_292; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62325; // @[Modules.scala 65:57:@11034.4]
  wire [10:0] _T_62326; // @[Modules.scala 65:57:@11035.4]
  wire [10:0] buffer_4_538; // @[Modules.scala 65:57:@11036.4]
  wire [11:0] _T_62328; // @[Modules.scala 65:57:@11038.4]
  wire [10:0] _T_62329; // @[Modules.scala 65:57:@11039.4]
  wire [10:0] buffer_4_539; // @[Modules.scala 65:57:@11040.4]
  wire [11:0] _T_62334; // @[Modules.scala 65:57:@11046.4]
  wire [10:0] _T_62335; // @[Modules.scala 65:57:@11047.4]
  wire [10:0] buffer_4_541; // @[Modules.scala 65:57:@11048.4]
  wire [11:0] _T_62343; // @[Modules.scala 65:57:@11058.4]
  wire [10:0] _T_62344; // @[Modules.scala 65:57:@11059.4]
  wire [10:0] buffer_4_544; // @[Modules.scala 65:57:@11060.4]
  wire [10:0] buffer_4_306; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_307; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62346; // @[Modules.scala 65:57:@11062.4]
  wire [10:0] _T_62347; // @[Modules.scala 65:57:@11063.4]
  wire [10:0] buffer_4_545; // @[Modules.scala 65:57:@11064.4]
  wire [10:0] buffer_4_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62352; // @[Modules.scala 65:57:@11070.4]
  wire [10:0] _T_62353; // @[Modules.scala 65:57:@11071.4]
  wire [10:0] buffer_4_547; // @[Modules.scala 65:57:@11072.4]
  wire [11:0] _T_62355; // @[Modules.scala 65:57:@11074.4]
  wire [10:0] _T_62356; // @[Modules.scala 65:57:@11075.4]
  wire [10:0] buffer_4_548; // @[Modules.scala 65:57:@11076.4]
  wire [10:0] buffer_4_316; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62361; // @[Modules.scala 65:57:@11082.4]
  wire [10:0] _T_62362; // @[Modules.scala 65:57:@11083.4]
  wire [10:0] buffer_4_550; // @[Modules.scala 65:57:@11084.4]
  wire [11:0] _T_62367; // @[Modules.scala 65:57:@11090.4]
  wire [10:0] _T_62368; // @[Modules.scala 65:57:@11091.4]
  wire [10:0] buffer_4_552; // @[Modules.scala 65:57:@11092.4]
  wire [10:0] buffer_4_324; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62373; // @[Modules.scala 65:57:@11098.4]
  wire [10:0] _T_62374; // @[Modules.scala 65:57:@11099.4]
  wire [10:0] buffer_4_554; // @[Modules.scala 65:57:@11100.4]
  wire [10:0] buffer_4_330; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62382; // @[Modules.scala 65:57:@11110.4]
  wire [10:0] _T_62383; // @[Modules.scala 65:57:@11111.4]
  wire [10:0] buffer_4_557; // @[Modules.scala 65:57:@11112.4]
  wire [11:0] _T_62385; // @[Modules.scala 65:57:@11114.4]
  wire [10:0] _T_62386; // @[Modules.scala 65:57:@11115.4]
  wire [10:0] buffer_4_558; // @[Modules.scala 65:57:@11116.4]
  wire [10:0] buffer_4_334; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_335; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62388; // @[Modules.scala 65:57:@11118.4]
  wire [10:0] _T_62389; // @[Modules.scala 65:57:@11119.4]
  wire [10:0] buffer_4_559; // @[Modules.scala 65:57:@11120.4]
  wire [10:0] buffer_4_336; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62391; // @[Modules.scala 65:57:@11122.4]
  wire [10:0] _T_62392; // @[Modules.scala 65:57:@11123.4]
  wire [10:0] buffer_4_560; // @[Modules.scala 65:57:@11124.4]
  wire [10:0] buffer_4_338; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62394; // @[Modules.scala 65:57:@11126.4]
  wire [10:0] _T_62395; // @[Modules.scala 65:57:@11127.4]
  wire [10:0] buffer_4_561; // @[Modules.scala 65:57:@11128.4]
  wire [11:0] _T_62400; // @[Modules.scala 65:57:@11134.4]
  wire [10:0] _T_62401; // @[Modules.scala 65:57:@11135.4]
  wire [10:0] buffer_4_563; // @[Modules.scala 65:57:@11136.4]
  wire [11:0] _T_62403; // @[Modules.scala 65:57:@11138.4]
  wire [10:0] _T_62404; // @[Modules.scala 65:57:@11139.4]
  wire [10:0] buffer_4_564; // @[Modules.scala 65:57:@11140.4]
  wire [10:0] buffer_4_348; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_4_349; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62409; // @[Modules.scala 65:57:@11146.4]
  wire [10:0] _T_62410; // @[Modules.scala 65:57:@11147.4]
  wire [10:0] buffer_4_566; // @[Modules.scala 65:57:@11148.4]
  wire [10:0] buffer_4_352; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62415; // @[Modules.scala 65:57:@11154.4]
  wire [10:0] _T_62416; // @[Modules.scala 65:57:@11155.4]
  wire [10:0] buffer_4_568; // @[Modules.scala 65:57:@11156.4]
  wire [10:0] buffer_4_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62430; // @[Modules.scala 65:57:@11174.4]
  wire [10:0] _T_62431; // @[Modules.scala 65:57:@11175.4]
  wire [10:0] buffer_4_573; // @[Modules.scala 65:57:@11176.4]
  wire [10:0] buffer_4_376; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62451; // @[Modules.scala 65:57:@11202.4]
  wire [10:0] _T_62452; // @[Modules.scala 65:57:@11203.4]
  wire [10:0] buffer_4_580; // @[Modules.scala 65:57:@11204.4]
  wire [11:0] _T_62454; // @[Modules.scala 65:57:@11206.4]
  wire [10:0] _T_62455; // @[Modules.scala 65:57:@11207.4]
  wire [10:0] buffer_4_581; // @[Modules.scala 65:57:@11208.4]
  wire [11:0] _T_62457; // @[Modules.scala 65:57:@11210.4]
  wire [10:0] _T_62458; // @[Modules.scala 65:57:@11211.4]
  wire [10:0] buffer_4_582; // @[Modules.scala 65:57:@11212.4]
  wire [10:0] buffer_4_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62460; // @[Modules.scala 65:57:@11214.4]
  wire [10:0] _T_62461; // @[Modules.scala 65:57:@11215.4]
  wire [10:0] buffer_4_583; // @[Modules.scala 65:57:@11216.4]
  wire [11:0] _T_62463; // @[Modules.scala 65:57:@11218.4]
  wire [10:0] _T_62464; // @[Modules.scala 65:57:@11219.4]
  wire [10:0] buffer_4_584; // @[Modules.scala 65:57:@11220.4]
  wire [10:0] buffer_4_386; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_62466; // @[Modules.scala 65:57:@11222.4]
  wire [10:0] _T_62467; // @[Modules.scala 65:57:@11223.4]
  wire [10:0] buffer_4_585; // @[Modules.scala 65:57:@11224.4]
  wire [11:0] _T_62472; // @[Modules.scala 65:57:@11230.4]
  wire [10:0] _T_62473; // @[Modules.scala 65:57:@11231.4]
  wire [10:0] buffer_4_587; // @[Modules.scala 65:57:@11232.4]
  wire [11:0] _T_62475; // @[Modules.scala 68:83:@11234.4]
  wire [10:0] _T_62476; // @[Modules.scala 68:83:@11235.4]
  wire [10:0] buffer_4_588; // @[Modules.scala 68:83:@11236.4]
  wire [11:0] _T_62478; // @[Modules.scala 68:83:@11238.4]
  wire [10:0] _T_62479; // @[Modules.scala 68:83:@11239.4]
  wire [10:0] buffer_4_589; // @[Modules.scala 68:83:@11240.4]
  wire [11:0] _T_62481; // @[Modules.scala 68:83:@11242.4]
  wire [10:0] _T_62482; // @[Modules.scala 68:83:@11243.4]
  wire [10:0] buffer_4_590; // @[Modules.scala 68:83:@11244.4]
  wire [11:0] _T_62484; // @[Modules.scala 68:83:@11246.4]
  wire [10:0] _T_62485; // @[Modules.scala 68:83:@11247.4]
  wire [10:0] buffer_4_591; // @[Modules.scala 68:83:@11248.4]
  wire [11:0] _T_62487; // @[Modules.scala 68:83:@11250.4]
  wire [10:0] _T_62488; // @[Modules.scala 68:83:@11251.4]
  wire [10:0] buffer_4_592; // @[Modules.scala 68:83:@11252.4]
  wire [11:0] _T_62490; // @[Modules.scala 68:83:@11254.4]
  wire [10:0] _T_62491; // @[Modules.scala 68:83:@11255.4]
  wire [10:0] buffer_4_593; // @[Modules.scala 68:83:@11256.4]
  wire [11:0] _T_62493; // @[Modules.scala 68:83:@11258.4]
  wire [10:0] _T_62494; // @[Modules.scala 68:83:@11259.4]
  wire [10:0] buffer_4_594; // @[Modules.scala 68:83:@11260.4]
  wire [11:0] _T_62496; // @[Modules.scala 68:83:@11262.4]
  wire [10:0] _T_62497; // @[Modules.scala 68:83:@11263.4]
  wire [10:0] buffer_4_595; // @[Modules.scala 68:83:@11264.4]
  wire [11:0] _T_62505; // @[Modules.scala 68:83:@11274.4]
  wire [10:0] _T_62506; // @[Modules.scala 68:83:@11275.4]
  wire [10:0] buffer_4_598; // @[Modules.scala 68:83:@11276.4]
  wire [11:0] _T_62508; // @[Modules.scala 68:83:@11278.4]
  wire [10:0] _T_62509; // @[Modules.scala 68:83:@11279.4]
  wire [10:0] buffer_4_599; // @[Modules.scala 68:83:@11280.4]
  wire [11:0] _T_62517; // @[Modules.scala 68:83:@11290.4]
  wire [10:0] _T_62518; // @[Modules.scala 68:83:@11291.4]
  wire [10:0] buffer_4_602; // @[Modules.scala 68:83:@11292.4]
  wire [11:0] _T_62520; // @[Modules.scala 68:83:@11294.4]
  wire [10:0] _T_62521; // @[Modules.scala 68:83:@11295.4]
  wire [10:0] buffer_4_603; // @[Modules.scala 68:83:@11296.4]
  wire [11:0] _T_62523; // @[Modules.scala 68:83:@11298.4]
  wire [10:0] _T_62524; // @[Modules.scala 68:83:@11299.4]
  wire [10:0] buffer_4_604; // @[Modules.scala 68:83:@11300.4]
  wire [11:0] _T_62526; // @[Modules.scala 68:83:@11302.4]
  wire [10:0] _T_62527; // @[Modules.scala 68:83:@11303.4]
  wire [10:0] buffer_4_605; // @[Modules.scala 68:83:@11304.4]
  wire [11:0] _T_62529; // @[Modules.scala 68:83:@11306.4]
  wire [10:0] _T_62530; // @[Modules.scala 68:83:@11307.4]
  wire [10:0] buffer_4_606; // @[Modules.scala 68:83:@11308.4]
  wire [11:0] _T_62532; // @[Modules.scala 68:83:@11310.4]
  wire [10:0] _T_62533; // @[Modules.scala 68:83:@11311.4]
  wire [10:0] buffer_4_607; // @[Modules.scala 68:83:@11312.4]
  wire [11:0] _T_62535; // @[Modules.scala 68:83:@11314.4]
  wire [10:0] _T_62536; // @[Modules.scala 68:83:@11315.4]
  wire [10:0] buffer_4_608; // @[Modules.scala 68:83:@11316.4]
  wire [11:0] _T_62538; // @[Modules.scala 68:83:@11318.4]
  wire [10:0] _T_62539; // @[Modules.scala 68:83:@11319.4]
  wire [10:0] buffer_4_609; // @[Modules.scala 68:83:@11320.4]
  wire [11:0] _T_62541; // @[Modules.scala 68:83:@11322.4]
  wire [10:0] _T_62542; // @[Modules.scala 68:83:@11323.4]
  wire [10:0] buffer_4_610; // @[Modules.scala 68:83:@11324.4]
  wire [11:0] _T_62544; // @[Modules.scala 68:83:@11326.4]
  wire [10:0] _T_62545; // @[Modules.scala 68:83:@11327.4]
  wire [10:0] buffer_4_611; // @[Modules.scala 68:83:@11328.4]
  wire [11:0] _T_62547; // @[Modules.scala 68:83:@11330.4]
  wire [10:0] _T_62548; // @[Modules.scala 68:83:@11331.4]
  wire [10:0] buffer_4_612; // @[Modules.scala 68:83:@11332.4]
  wire [11:0] _T_62550; // @[Modules.scala 68:83:@11334.4]
  wire [10:0] _T_62551; // @[Modules.scala 68:83:@11335.4]
  wire [10:0] buffer_4_613; // @[Modules.scala 68:83:@11336.4]
  wire [11:0] _T_62559; // @[Modules.scala 68:83:@11346.4]
  wire [10:0] _T_62560; // @[Modules.scala 68:83:@11347.4]
  wire [10:0] buffer_4_616; // @[Modules.scala 68:83:@11348.4]
  wire [11:0] _T_62562; // @[Modules.scala 68:83:@11350.4]
  wire [10:0] _T_62563; // @[Modules.scala 68:83:@11351.4]
  wire [10:0] buffer_4_617; // @[Modules.scala 68:83:@11352.4]
  wire [11:0] _T_62565; // @[Modules.scala 68:83:@11354.4]
  wire [10:0] _T_62566; // @[Modules.scala 68:83:@11355.4]
  wire [10:0] buffer_4_618; // @[Modules.scala 68:83:@11356.4]
  wire [11:0] _T_62571; // @[Modules.scala 68:83:@11362.4]
  wire [10:0] _T_62572; // @[Modules.scala 68:83:@11363.4]
  wire [10:0] buffer_4_620; // @[Modules.scala 68:83:@11364.4]
  wire [11:0] _T_62580; // @[Modules.scala 68:83:@11374.4]
  wire [10:0] _T_62581; // @[Modules.scala 68:83:@11375.4]
  wire [10:0] buffer_4_623; // @[Modules.scala 68:83:@11376.4]
  wire [11:0] _T_62586; // @[Modules.scala 68:83:@11382.4]
  wire [10:0] _T_62587; // @[Modules.scala 68:83:@11383.4]
  wire [10:0] buffer_4_625; // @[Modules.scala 68:83:@11384.4]
  wire [11:0] _T_62589; // @[Modules.scala 68:83:@11386.4]
  wire [10:0] _T_62590; // @[Modules.scala 68:83:@11387.4]
  wire [10:0] buffer_4_626; // @[Modules.scala 68:83:@11388.4]
  wire [11:0] _T_62592; // @[Modules.scala 68:83:@11390.4]
  wire [10:0] _T_62593; // @[Modules.scala 68:83:@11391.4]
  wire [10:0] buffer_4_627; // @[Modules.scala 68:83:@11392.4]
  wire [11:0] _T_62595; // @[Modules.scala 68:83:@11394.4]
  wire [10:0] _T_62596; // @[Modules.scala 68:83:@11395.4]
  wire [10:0] buffer_4_628; // @[Modules.scala 68:83:@11396.4]
  wire [11:0] _T_62598; // @[Modules.scala 68:83:@11398.4]
  wire [10:0] _T_62599; // @[Modules.scala 68:83:@11399.4]
  wire [10:0] buffer_4_629; // @[Modules.scala 68:83:@11400.4]
  wire [11:0] _T_62601; // @[Modules.scala 68:83:@11402.4]
  wire [10:0] _T_62602; // @[Modules.scala 68:83:@11403.4]
  wire [10:0] buffer_4_630; // @[Modules.scala 68:83:@11404.4]
  wire [11:0] _T_62604; // @[Modules.scala 68:83:@11406.4]
  wire [10:0] _T_62605; // @[Modules.scala 68:83:@11407.4]
  wire [10:0] buffer_4_631; // @[Modules.scala 68:83:@11408.4]
  wire [11:0] _T_62607; // @[Modules.scala 68:83:@11410.4]
  wire [10:0] _T_62608; // @[Modules.scala 68:83:@11411.4]
  wire [10:0] buffer_4_632; // @[Modules.scala 68:83:@11412.4]
  wire [11:0] _T_62610; // @[Modules.scala 68:83:@11414.4]
  wire [10:0] _T_62611; // @[Modules.scala 68:83:@11415.4]
  wire [10:0] buffer_4_633; // @[Modules.scala 68:83:@11416.4]
  wire [11:0] _T_62613; // @[Modules.scala 68:83:@11418.4]
  wire [10:0] _T_62614; // @[Modules.scala 68:83:@11419.4]
  wire [10:0] buffer_4_634; // @[Modules.scala 68:83:@11420.4]
  wire [11:0] _T_62616; // @[Modules.scala 68:83:@11422.4]
  wire [10:0] _T_62617; // @[Modules.scala 68:83:@11423.4]
  wire [10:0] buffer_4_635; // @[Modules.scala 68:83:@11424.4]
  wire [11:0] _T_62619; // @[Modules.scala 68:83:@11426.4]
  wire [10:0] _T_62620; // @[Modules.scala 68:83:@11427.4]
  wire [10:0] buffer_4_636; // @[Modules.scala 68:83:@11428.4]
  wire [11:0] _T_62622; // @[Modules.scala 68:83:@11430.4]
  wire [10:0] _T_62623; // @[Modules.scala 68:83:@11431.4]
  wire [10:0] buffer_4_637; // @[Modules.scala 68:83:@11432.4]
  wire [11:0] _T_62625; // @[Modules.scala 68:83:@11434.4]
  wire [10:0] _T_62626; // @[Modules.scala 68:83:@11435.4]
  wire [10:0] buffer_4_638; // @[Modules.scala 68:83:@11436.4]
  wire [11:0] _T_62628; // @[Modules.scala 68:83:@11438.4]
  wire [10:0] _T_62629; // @[Modules.scala 68:83:@11439.4]
  wire [10:0] buffer_4_639; // @[Modules.scala 68:83:@11440.4]
  wire [11:0] _T_62631; // @[Modules.scala 68:83:@11442.4]
  wire [10:0] _T_62632; // @[Modules.scala 68:83:@11443.4]
  wire [10:0] buffer_4_640; // @[Modules.scala 68:83:@11444.4]
  wire [11:0] _T_62634; // @[Modules.scala 68:83:@11446.4]
  wire [10:0] _T_62635; // @[Modules.scala 68:83:@11447.4]
  wire [10:0] buffer_4_641; // @[Modules.scala 68:83:@11448.4]
  wire [11:0] _T_62637; // @[Modules.scala 68:83:@11450.4]
  wire [10:0] _T_62638; // @[Modules.scala 68:83:@11451.4]
  wire [10:0] buffer_4_642; // @[Modules.scala 68:83:@11452.4]
  wire [11:0] _T_62640; // @[Modules.scala 68:83:@11454.4]
  wire [10:0] _T_62641; // @[Modules.scala 68:83:@11455.4]
  wire [10:0] buffer_4_643; // @[Modules.scala 68:83:@11456.4]
  wire [11:0] _T_62643; // @[Modules.scala 68:83:@11458.4]
  wire [10:0] _T_62644; // @[Modules.scala 68:83:@11459.4]
  wire [10:0] buffer_4_644; // @[Modules.scala 68:83:@11460.4]
  wire [11:0] _T_62646; // @[Modules.scala 68:83:@11462.4]
  wire [10:0] _T_62647; // @[Modules.scala 68:83:@11463.4]
  wire [10:0] buffer_4_645; // @[Modules.scala 68:83:@11464.4]
  wire [11:0] _T_62649; // @[Modules.scala 68:83:@11466.4]
  wire [10:0] _T_62650; // @[Modules.scala 68:83:@11467.4]
  wire [10:0] buffer_4_646; // @[Modules.scala 68:83:@11468.4]
  wire [11:0] _T_62652; // @[Modules.scala 68:83:@11470.4]
  wire [10:0] _T_62653; // @[Modules.scala 68:83:@11471.4]
  wire [10:0] buffer_4_647; // @[Modules.scala 68:83:@11472.4]
  wire [11:0] _T_62655; // @[Modules.scala 68:83:@11474.4]
  wire [10:0] _T_62656; // @[Modules.scala 68:83:@11475.4]
  wire [10:0] buffer_4_648; // @[Modules.scala 68:83:@11476.4]
  wire [11:0] _T_62658; // @[Modules.scala 68:83:@11478.4]
  wire [10:0] _T_62659; // @[Modules.scala 68:83:@11479.4]
  wire [10:0] buffer_4_649; // @[Modules.scala 68:83:@11480.4]
  wire [11:0] _T_62664; // @[Modules.scala 68:83:@11486.4]
  wire [10:0] _T_62665; // @[Modules.scala 68:83:@11487.4]
  wire [10:0] buffer_4_651; // @[Modules.scala 68:83:@11488.4]
  wire [11:0] _T_62667; // @[Modules.scala 68:83:@11490.4]
  wire [10:0] _T_62668; // @[Modules.scala 68:83:@11491.4]
  wire [10:0] buffer_4_652; // @[Modules.scala 68:83:@11492.4]
  wire [11:0] _T_62670; // @[Modules.scala 68:83:@11494.4]
  wire [10:0] _T_62671; // @[Modules.scala 68:83:@11495.4]
  wire [10:0] buffer_4_653; // @[Modules.scala 68:83:@11496.4]
  wire [11:0] _T_62673; // @[Modules.scala 68:83:@11498.4]
  wire [10:0] _T_62674; // @[Modules.scala 68:83:@11499.4]
  wire [10:0] buffer_4_654; // @[Modules.scala 68:83:@11500.4]
  wire [11:0] _T_62679; // @[Modules.scala 68:83:@11506.4]
  wire [10:0] _T_62680; // @[Modules.scala 68:83:@11507.4]
  wire [10:0] buffer_4_656; // @[Modules.scala 68:83:@11508.4]
  wire [11:0] _T_62682; // @[Modules.scala 68:83:@11510.4]
  wire [10:0] _T_62683; // @[Modules.scala 68:83:@11511.4]
  wire [10:0] buffer_4_657; // @[Modules.scala 68:83:@11512.4]
  wire [11:0] _T_62685; // @[Modules.scala 68:83:@11514.4]
  wire [10:0] _T_62686; // @[Modules.scala 68:83:@11515.4]
  wire [10:0] buffer_4_658; // @[Modules.scala 68:83:@11516.4]
  wire [11:0] _T_62688; // @[Modules.scala 68:83:@11518.4]
  wire [10:0] _T_62689; // @[Modules.scala 68:83:@11519.4]
  wire [10:0] buffer_4_659; // @[Modules.scala 68:83:@11520.4]
  wire [11:0] _T_62691; // @[Modules.scala 68:83:@11522.4]
  wire [10:0] _T_62692; // @[Modules.scala 68:83:@11523.4]
  wire [10:0] buffer_4_660; // @[Modules.scala 68:83:@11524.4]
  wire [11:0] _T_62694; // @[Modules.scala 68:83:@11526.4]
  wire [10:0] _T_62695; // @[Modules.scala 68:83:@11527.4]
  wire [10:0] buffer_4_661; // @[Modules.scala 68:83:@11528.4]
  wire [11:0] _T_62697; // @[Modules.scala 68:83:@11530.4]
  wire [10:0] _T_62698; // @[Modules.scala 68:83:@11531.4]
  wire [10:0] buffer_4_662; // @[Modules.scala 68:83:@11532.4]
  wire [11:0] _T_62703; // @[Modules.scala 68:83:@11538.4]
  wire [10:0] _T_62704; // @[Modules.scala 68:83:@11539.4]
  wire [10:0] buffer_4_664; // @[Modules.scala 68:83:@11540.4]
  wire [11:0] _T_62706; // @[Modules.scala 68:83:@11542.4]
  wire [10:0] _T_62707; // @[Modules.scala 68:83:@11543.4]
  wire [10:0] buffer_4_665; // @[Modules.scala 68:83:@11544.4]
  wire [11:0] _T_62709; // @[Modules.scala 68:83:@11546.4]
  wire [10:0] _T_62710; // @[Modules.scala 68:83:@11547.4]
  wire [10:0] buffer_4_666; // @[Modules.scala 68:83:@11548.4]
  wire [11:0] _T_62712; // @[Modules.scala 68:83:@11550.4]
  wire [10:0] _T_62713; // @[Modules.scala 68:83:@11551.4]
  wire [10:0] buffer_4_667; // @[Modules.scala 68:83:@11552.4]
  wire [11:0] _T_62715; // @[Modules.scala 68:83:@11554.4]
  wire [10:0] _T_62716; // @[Modules.scala 68:83:@11555.4]
  wire [10:0] buffer_4_668; // @[Modules.scala 68:83:@11556.4]
  wire [11:0] _T_62718; // @[Modules.scala 68:83:@11558.4]
  wire [10:0] _T_62719; // @[Modules.scala 68:83:@11559.4]
  wire [10:0] buffer_4_669; // @[Modules.scala 68:83:@11560.4]
  wire [11:0] _T_62721; // @[Modules.scala 68:83:@11562.4]
  wire [10:0] _T_62722; // @[Modules.scala 68:83:@11563.4]
  wire [10:0] buffer_4_670; // @[Modules.scala 68:83:@11564.4]
  wire [11:0] _T_62724; // @[Modules.scala 68:83:@11566.4]
  wire [10:0] _T_62725; // @[Modules.scala 68:83:@11567.4]
  wire [10:0] buffer_4_671; // @[Modules.scala 68:83:@11568.4]
  wire [11:0] _T_62727; // @[Modules.scala 68:83:@11570.4]
  wire [10:0] _T_62728; // @[Modules.scala 68:83:@11571.4]
  wire [10:0] buffer_4_672; // @[Modules.scala 68:83:@11572.4]
  wire [11:0] _T_62730; // @[Modules.scala 68:83:@11574.4]
  wire [10:0] _T_62731; // @[Modules.scala 68:83:@11575.4]
  wire [10:0] buffer_4_673; // @[Modules.scala 68:83:@11576.4]
  wire [11:0] _T_62733; // @[Modules.scala 68:83:@11578.4]
  wire [10:0] _T_62734; // @[Modules.scala 68:83:@11579.4]
  wire [10:0] buffer_4_674; // @[Modules.scala 68:83:@11580.4]
  wire [11:0] _T_62736; // @[Modules.scala 68:83:@11582.4]
  wire [10:0] _T_62737; // @[Modules.scala 68:83:@11583.4]
  wire [10:0] buffer_4_675; // @[Modules.scala 68:83:@11584.4]
  wire [11:0] _T_62739; // @[Modules.scala 68:83:@11586.4]
  wire [10:0] _T_62740; // @[Modules.scala 68:83:@11587.4]
  wire [10:0] buffer_4_676; // @[Modules.scala 68:83:@11588.4]
  wire [11:0] _T_62745; // @[Modules.scala 68:83:@11594.4]
  wire [10:0] _T_62746; // @[Modules.scala 68:83:@11595.4]
  wire [10:0] buffer_4_678; // @[Modules.scala 68:83:@11596.4]
  wire [11:0] _T_62748; // @[Modules.scala 68:83:@11598.4]
  wire [10:0] _T_62749; // @[Modules.scala 68:83:@11599.4]
  wire [10:0] buffer_4_679; // @[Modules.scala 68:83:@11600.4]
  wire [11:0] _T_62757; // @[Modules.scala 68:83:@11610.4]
  wire [10:0] _T_62758; // @[Modules.scala 68:83:@11611.4]
  wire [10:0] buffer_4_682; // @[Modules.scala 68:83:@11612.4]
  wire [11:0] _T_62760; // @[Modules.scala 68:83:@11614.4]
  wire [10:0] _T_62761; // @[Modules.scala 68:83:@11615.4]
  wire [10:0] buffer_4_683; // @[Modules.scala 68:83:@11616.4]
  wire [11:0] _T_62763; // @[Modules.scala 68:83:@11618.4]
  wire [10:0] _T_62764; // @[Modules.scala 68:83:@11619.4]
  wire [10:0] buffer_4_684; // @[Modules.scala 68:83:@11620.4]
  wire [11:0] _T_62766; // @[Modules.scala 68:83:@11622.4]
  wire [10:0] _T_62767; // @[Modules.scala 68:83:@11623.4]
  wire [10:0] buffer_4_685; // @[Modules.scala 68:83:@11624.4]
  wire [11:0] _T_62769; // @[Modules.scala 71:109:@11626.4]
  wire [10:0] _T_62770; // @[Modules.scala 71:109:@11627.4]
  wire [10:0] buffer_4_686; // @[Modules.scala 71:109:@11628.4]
  wire [11:0] _T_62772; // @[Modules.scala 71:109:@11630.4]
  wire [10:0] _T_62773; // @[Modules.scala 71:109:@11631.4]
  wire [10:0] buffer_4_687; // @[Modules.scala 71:109:@11632.4]
  wire [11:0] _T_62775; // @[Modules.scala 71:109:@11634.4]
  wire [10:0] _T_62776; // @[Modules.scala 71:109:@11635.4]
  wire [10:0] buffer_4_688; // @[Modules.scala 71:109:@11636.4]
  wire [11:0] _T_62778; // @[Modules.scala 71:109:@11638.4]
  wire [10:0] _T_62779; // @[Modules.scala 71:109:@11639.4]
  wire [10:0] buffer_4_689; // @[Modules.scala 71:109:@11640.4]
  wire [11:0] _T_62784; // @[Modules.scala 71:109:@11646.4]
  wire [10:0] _T_62785; // @[Modules.scala 71:109:@11647.4]
  wire [10:0] buffer_4_691; // @[Modules.scala 71:109:@11648.4]
  wire [11:0] _T_62790; // @[Modules.scala 71:109:@11654.4]
  wire [10:0] _T_62791; // @[Modules.scala 71:109:@11655.4]
  wire [10:0] buffer_4_693; // @[Modules.scala 71:109:@11656.4]
  wire [11:0] _T_62793; // @[Modules.scala 71:109:@11658.4]
  wire [10:0] _T_62794; // @[Modules.scala 71:109:@11659.4]
  wire [10:0] buffer_4_694; // @[Modules.scala 71:109:@11660.4]
  wire [11:0] _T_62796; // @[Modules.scala 71:109:@11662.4]
  wire [10:0] _T_62797; // @[Modules.scala 71:109:@11663.4]
  wire [10:0] buffer_4_695; // @[Modules.scala 71:109:@11664.4]
  wire [11:0] _T_62799; // @[Modules.scala 71:109:@11666.4]
  wire [10:0] _T_62800; // @[Modules.scala 71:109:@11667.4]
  wire [10:0] buffer_4_696; // @[Modules.scala 71:109:@11668.4]
  wire [11:0] _T_62802; // @[Modules.scala 71:109:@11670.4]
  wire [10:0] _T_62803; // @[Modules.scala 71:109:@11671.4]
  wire [10:0] buffer_4_697; // @[Modules.scala 71:109:@11672.4]
  wire [11:0] _T_62805; // @[Modules.scala 71:109:@11674.4]
  wire [10:0] _T_62806; // @[Modules.scala 71:109:@11675.4]
  wire [10:0] buffer_4_698; // @[Modules.scala 71:109:@11676.4]
  wire [11:0] _T_62808; // @[Modules.scala 71:109:@11678.4]
  wire [10:0] _T_62809; // @[Modules.scala 71:109:@11679.4]
  wire [10:0] buffer_4_699; // @[Modules.scala 71:109:@11680.4]
  wire [11:0] _T_62811; // @[Modules.scala 71:109:@11682.4]
  wire [10:0] _T_62812; // @[Modules.scala 71:109:@11683.4]
  wire [10:0] buffer_4_700; // @[Modules.scala 71:109:@11684.4]
  wire [11:0] _T_62814; // @[Modules.scala 71:109:@11686.4]
  wire [10:0] _T_62815; // @[Modules.scala 71:109:@11687.4]
  wire [10:0] buffer_4_701; // @[Modules.scala 71:109:@11688.4]
  wire [11:0] _T_62817; // @[Modules.scala 71:109:@11690.4]
  wire [10:0] _T_62818; // @[Modules.scala 71:109:@11691.4]
  wire [10:0] buffer_4_702; // @[Modules.scala 71:109:@11692.4]
  wire [11:0] _T_62820; // @[Modules.scala 71:109:@11694.4]
  wire [10:0] _T_62821; // @[Modules.scala 71:109:@11695.4]
  wire [10:0] buffer_4_703; // @[Modules.scala 71:109:@11696.4]
  wire [11:0] _T_62823; // @[Modules.scala 71:109:@11698.4]
  wire [10:0] _T_62824; // @[Modules.scala 71:109:@11699.4]
  wire [10:0] buffer_4_704; // @[Modules.scala 71:109:@11700.4]
  wire [11:0] _T_62826; // @[Modules.scala 71:109:@11702.4]
  wire [10:0] _T_62827; // @[Modules.scala 71:109:@11703.4]
  wire [10:0] buffer_4_705; // @[Modules.scala 71:109:@11704.4]
  wire [11:0] _T_62829; // @[Modules.scala 71:109:@11706.4]
  wire [10:0] _T_62830; // @[Modules.scala 71:109:@11707.4]
  wire [10:0] buffer_4_706; // @[Modules.scala 71:109:@11708.4]
  wire [11:0] _T_62832; // @[Modules.scala 71:109:@11710.4]
  wire [10:0] _T_62833; // @[Modules.scala 71:109:@11711.4]
  wire [10:0] buffer_4_707; // @[Modules.scala 71:109:@11712.4]
  wire [11:0] _T_62835; // @[Modules.scala 71:109:@11714.4]
  wire [10:0] _T_62836; // @[Modules.scala 71:109:@11715.4]
  wire [10:0] buffer_4_708; // @[Modules.scala 71:109:@11716.4]
  wire [11:0] _T_62838; // @[Modules.scala 71:109:@11718.4]
  wire [10:0] _T_62839; // @[Modules.scala 71:109:@11719.4]
  wire [10:0] buffer_4_709; // @[Modules.scala 71:109:@11720.4]
  wire [11:0] _T_62841; // @[Modules.scala 71:109:@11722.4]
  wire [10:0] _T_62842; // @[Modules.scala 71:109:@11723.4]
  wire [10:0] buffer_4_710; // @[Modules.scala 71:109:@11724.4]
  wire [11:0] _T_62844; // @[Modules.scala 71:109:@11726.4]
  wire [10:0] _T_62845; // @[Modules.scala 71:109:@11727.4]
  wire [10:0] buffer_4_711; // @[Modules.scala 71:109:@11728.4]
  wire [11:0] _T_62847; // @[Modules.scala 71:109:@11730.4]
  wire [10:0] _T_62848; // @[Modules.scala 71:109:@11731.4]
  wire [10:0] buffer_4_712; // @[Modules.scala 71:109:@11732.4]
  wire [11:0] _T_62850; // @[Modules.scala 71:109:@11734.4]
  wire [10:0] _T_62851; // @[Modules.scala 71:109:@11735.4]
  wire [10:0] buffer_4_713; // @[Modules.scala 71:109:@11736.4]
  wire [11:0] _T_62853; // @[Modules.scala 71:109:@11738.4]
  wire [10:0] _T_62854; // @[Modules.scala 71:109:@11739.4]
  wire [10:0] buffer_4_714; // @[Modules.scala 71:109:@11740.4]
  wire [11:0] _T_62856; // @[Modules.scala 71:109:@11742.4]
  wire [10:0] _T_62857; // @[Modules.scala 71:109:@11743.4]
  wire [10:0] buffer_4_715; // @[Modules.scala 71:109:@11744.4]
  wire [11:0] _T_62859; // @[Modules.scala 71:109:@11746.4]
  wire [10:0] _T_62860; // @[Modules.scala 71:109:@11747.4]
  wire [10:0] buffer_4_716; // @[Modules.scala 71:109:@11748.4]
  wire [11:0] _T_62862; // @[Modules.scala 71:109:@11750.4]
  wire [10:0] _T_62863; // @[Modules.scala 71:109:@11751.4]
  wire [10:0] buffer_4_717; // @[Modules.scala 71:109:@11752.4]
  wire [11:0] _T_62865; // @[Modules.scala 71:109:@11754.4]
  wire [10:0] _T_62866; // @[Modules.scala 71:109:@11755.4]
  wire [10:0] buffer_4_718; // @[Modules.scala 71:109:@11756.4]
  wire [11:0] _T_62868; // @[Modules.scala 71:109:@11758.4]
  wire [10:0] _T_62869; // @[Modules.scala 71:109:@11759.4]
  wire [10:0] buffer_4_719; // @[Modules.scala 71:109:@11760.4]
  wire [11:0] _T_62871; // @[Modules.scala 71:109:@11762.4]
  wire [10:0] _T_62872; // @[Modules.scala 71:109:@11763.4]
  wire [10:0] buffer_4_720; // @[Modules.scala 71:109:@11764.4]
  wire [11:0] _T_62874; // @[Modules.scala 71:109:@11766.4]
  wire [10:0] _T_62875; // @[Modules.scala 71:109:@11767.4]
  wire [10:0] buffer_4_721; // @[Modules.scala 71:109:@11768.4]
  wire [11:0] _T_62877; // @[Modules.scala 71:109:@11770.4]
  wire [10:0] _T_62878; // @[Modules.scala 71:109:@11771.4]
  wire [10:0] buffer_4_722; // @[Modules.scala 71:109:@11772.4]
  wire [11:0] _T_62880; // @[Modules.scala 71:109:@11774.4]
  wire [10:0] _T_62881; // @[Modules.scala 71:109:@11775.4]
  wire [10:0] buffer_4_723; // @[Modules.scala 71:109:@11776.4]
  wire [11:0] _T_62883; // @[Modules.scala 71:109:@11778.4]
  wire [10:0] _T_62884; // @[Modules.scala 71:109:@11779.4]
  wire [10:0] buffer_4_724; // @[Modules.scala 71:109:@11780.4]
  wire [11:0] _T_62886; // @[Modules.scala 71:109:@11782.4]
  wire [10:0] _T_62887; // @[Modules.scala 71:109:@11783.4]
  wire [10:0] buffer_4_725; // @[Modules.scala 71:109:@11784.4]
  wire [11:0] _T_62889; // @[Modules.scala 71:109:@11786.4]
  wire [10:0] _T_62890; // @[Modules.scala 71:109:@11787.4]
  wire [10:0] buffer_4_726; // @[Modules.scala 71:109:@11788.4]
  wire [11:0] _T_62892; // @[Modules.scala 71:109:@11790.4]
  wire [10:0] _T_62893; // @[Modules.scala 71:109:@11791.4]
  wire [10:0] buffer_4_727; // @[Modules.scala 71:109:@11792.4]
  wire [11:0] _T_62895; // @[Modules.scala 71:109:@11794.4]
  wire [10:0] _T_62896; // @[Modules.scala 71:109:@11795.4]
  wire [10:0] buffer_4_728; // @[Modules.scala 71:109:@11796.4]
  wire [11:0] _T_62898; // @[Modules.scala 71:109:@11798.4]
  wire [10:0] _T_62899; // @[Modules.scala 71:109:@11799.4]
  wire [10:0] buffer_4_729; // @[Modules.scala 71:109:@11800.4]
  wire [11:0] _T_62901; // @[Modules.scala 71:109:@11802.4]
  wire [10:0] _T_62902; // @[Modules.scala 71:109:@11803.4]
  wire [10:0] buffer_4_730; // @[Modules.scala 71:109:@11804.4]
  wire [11:0] _T_62904; // @[Modules.scala 71:109:@11806.4]
  wire [10:0] _T_62905; // @[Modules.scala 71:109:@11807.4]
  wire [10:0] buffer_4_731; // @[Modules.scala 71:109:@11808.4]
  wire [11:0] _T_62910; // @[Modules.scala 71:109:@11814.4]
  wire [10:0] _T_62911; // @[Modules.scala 71:109:@11815.4]
  wire [10:0] buffer_4_733; // @[Modules.scala 71:109:@11816.4]
  wire [11:0] _T_62913; // @[Modules.scala 71:109:@11818.4]
  wire [10:0] _T_62914; // @[Modules.scala 71:109:@11819.4]
  wire [10:0] buffer_4_734; // @[Modules.scala 71:109:@11820.4]
  wire [11:0] _T_62916; // @[Modules.scala 78:156:@11823.4]
  wire [10:0] _T_62917; // @[Modules.scala 78:156:@11824.4]
  wire [10:0] buffer_4_736; // @[Modules.scala 78:156:@11825.4]
  wire [11:0] _T_62919; // @[Modules.scala 78:156:@11827.4]
  wire [10:0] _T_62920; // @[Modules.scala 78:156:@11828.4]
  wire [10:0] buffer_4_737; // @[Modules.scala 78:156:@11829.4]
  wire [11:0] _T_62922; // @[Modules.scala 78:156:@11831.4]
  wire [10:0] _T_62923; // @[Modules.scala 78:156:@11832.4]
  wire [10:0] buffer_4_738; // @[Modules.scala 78:156:@11833.4]
  wire [11:0] _T_62925; // @[Modules.scala 78:156:@11835.4]
  wire [10:0] _T_62926; // @[Modules.scala 78:156:@11836.4]
  wire [10:0] buffer_4_739; // @[Modules.scala 78:156:@11837.4]
  wire [11:0] _T_62928; // @[Modules.scala 78:156:@11839.4]
  wire [10:0] _T_62929; // @[Modules.scala 78:156:@11840.4]
  wire [10:0] buffer_4_740; // @[Modules.scala 78:156:@11841.4]
  wire [11:0] _T_62931; // @[Modules.scala 78:156:@11843.4]
  wire [10:0] _T_62932; // @[Modules.scala 78:156:@11844.4]
  wire [10:0] buffer_4_741; // @[Modules.scala 78:156:@11845.4]
  wire [11:0] _T_62934; // @[Modules.scala 78:156:@11847.4]
  wire [10:0] _T_62935; // @[Modules.scala 78:156:@11848.4]
  wire [10:0] buffer_4_742; // @[Modules.scala 78:156:@11849.4]
  wire [11:0] _T_62937; // @[Modules.scala 78:156:@11851.4]
  wire [10:0] _T_62938; // @[Modules.scala 78:156:@11852.4]
  wire [10:0] buffer_4_743; // @[Modules.scala 78:156:@11853.4]
  wire [11:0] _T_62940; // @[Modules.scala 78:156:@11855.4]
  wire [10:0] _T_62941; // @[Modules.scala 78:156:@11856.4]
  wire [10:0] buffer_4_744; // @[Modules.scala 78:156:@11857.4]
  wire [11:0] _T_62943; // @[Modules.scala 78:156:@11859.4]
  wire [10:0] _T_62944; // @[Modules.scala 78:156:@11860.4]
  wire [10:0] buffer_4_745; // @[Modules.scala 78:156:@11861.4]
  wire [11:0] _T_62946; // @[Modules.scala 78:156:@11863.4]
  wire [10:0] _T_62947; // @[Modules.scala 78:156:@11864.4]
  wire [10:0] buffer_4_746; // @[Modules.scala 78:156:@11865.4]
  wire [11:0] _T_62949; // @[Modules.scala 78:156:@11867.4]
  wire [10:0] _T_62950; // @[Modules.scala 78:156:@11868.4]
  wire [10:0] buffer_4_747; // @[Modules.scala 78:156:@11869.4]
  wire [11:0] _T_62952; // @[Modules.scala 78:156:@11871.4]
  wire [10:0] _T_62953; // @[Modules.scala 78:156:@11872.4]
  wire [10:0] buffer_4_748; // @[Modules.scala 78:156:@11873.4]
  wire [11:0] _T_62955; // @[Modules.scala 78:156:@11875.4]
  wire [10:0] _T_62956; // @[Modules.scala 78:156:@11876.4]
  wire [10:0] buffer_4_749; // @[Modules.scala 78:156:@11877.4]
  wire [11:0] _T_62958; // @[Modules.scala 78:156:@11879.4]
  wire [10:0] _T_62959; // @[Modules.scala 78:156:@11880.4]
  wire [10:0] buffer_4_750; // @[Modules.scala 78:156:@11881.4]
  wire [11:0] _T_62961; // @[Modules.scala 78:156:@11883.4]
  wire [10:0] _T_62962; // @[Modules.scala 78:156:@11884.4]
  wire [10:0] buffer_4_751; // @[Modules.scala 78:156:@11885.4]
  wire [11:0] _T_62964; // @[Modules.scala 78:156:@11887.4]
  wire [10:0] _T_62965; // @[Modules.scala 78:156:@11888.4]
  wire [10:0] buffer_4_752; // @[Modules.scala 78:156:@11889.4]
  wire [11:0] _T_62967; // @[Modules.scala 78:156:@11891.4]
  wire [10:0] _T_62968; // @[Modules.scala 78:156:@11892.4]
  wire [10:0] buffer_4_753; // @[Modules.scala 78:156:@11893.4]
  wire [11:0] _T_62970; // @[Modules.scala 78:156:@11895.4]
  wire [10:0] _T_62971; // @[Modules.scala 78:156:@11896.4]
  wire [10:0] buffer_4_754; // @[Modules.scala 78:156:@11897.4]
  wire [11:0] _T_62973; // @[Modules.scala 78:156:@11899.4]
  wire [10:0] _T_62974; // @[Modules.scala 78:156:@11900.4]
  wire [10:0] buffer_4_755; // @[Modules.scala 78:156:@11901.4]
  wire [11:0] _T_62976; // @[Modules.scala 78:156:@11903.4]
  wire [10:0] _T_62977; // @[Modules.scala 78:156:@11904.4]
  wire [10:0] buffer_4_756; // @[Modules.scala 78:156:@11905.4]
  wire [11:0] _T_62979; // @[Modules.scala 78:156:@11907.4]
  wire [10:0] _T_62980; // @[Modules.scala 78:156:@11908.4]
  wire [10:0] buffer_4_757; // @[Modules.scala 78:156:@11909.4]
  wire [11:0] _T_62982; // @[Modules.scala 78:156:@11911.4]
  wire [10:0] _T_62983; // @[Modules.scala 78:156:@11912.4]
  wire [10:0] buffer_4_758; // @[Modules.scala 78:156:@11913.4]
  wire [11:0] _T_62985; // @[Modules.scala 78:156:@11915.4]
  wire [10:0] _T_62986; // @[Modules.scala 78:156:@11916.4]
  wire [10:0] buffer_4_759; // @[Modules.scala 78:156:@11917.4]
  wire [11:0] _T_62988; // @[Modules.scala 78:156:@11919.4]
  wire [10:0] _T_62989; // @[Modules.scala 78:156:@11920.4]
  wire [10:0] buffer_4_760; // @[Modules.scala 78:156:@11921.4]
  wire [11:0] _T_62991; // @[Modules.scala 78:156:@11923.4]
  wire [10:0] _T_62992; // @[Modules.scala 78:156:@11924.4]
  wire [10:0] buffer_4_761; // @[Modules.scala 78:156:@11925.4]
  wire [11:0] _T_62994; // @[Modules.scala 78:156:@11927.4]
  wire [10:0] _T_62995; // @[Modules.scala 78:156:@11928.4]
  wire [10:0] buffer_4_762; // @[Modules.scala 78:156:@11929.4]
  wire [11:0] _T_62997; // @[Modules.scala 78:156:@11931.4]
  wire [10:0] _T_62998; // @[Modules.scala 78:156:@11932.4]
  wire [10:0] buffer_4_763; // @[Modules.scala 78:156:@11933.4]
  wire [11:0] _T_63000; // @[Modules.scala 78:156:@11935.4]
  wire [10:0] _T_63001; // @[Modules.scala 78:156:@11936.4]
  wire [10:0] buffer_4_764; // @[Modules.scala 78:156:@11937.4]
  wire [11:0] _T_63003; // @[Modules.scala 78:156:@11939.4]
  wire [10:0] _T_63004; // @[Modules.scala 78:156:@11940.4]
  wire [10:0] buffer_4_765; // @[Modules.scala 78:156:@11941.4]
  wire [11:0] _T_63006; // @[Modules.scala 78:156:@11943.4]
  wire [10:0] _T_63007; // @[Modules.scala 78:156:@11944.4]
  wire [10:0] buffer_4_766; // @[Modules.scala 78:156:@11945.4]
  wire [11:0] _T_63009; // @[Modules.scala 78:156:@11947.4]
  wire [10:0] _T_63010; // @[Modules.scala 78:156:@11948.4]
  wire [10:0] buffer_4_767; // @[Modules.scala 78:156:@11949.4]
  wire [11:0] _T_63012; // @[Modules.scala 78:156:@11951.4]
  wire [10:0] _T_63013; // @[Modules.scala 78:156:@11952.4]
  wire [10:0] buffer_4_768; // @[Modules.scala 78:156:@11953.4]
  wire [11:0] _T_63015; // @[Modules.scala 78:156:@11955.4]
  wire [10:0] _T_63016; // @[Modules.scala 78:156:@11956.4]
  wire [10:0] buffer_4_769; // @[Modules.scala 78:156:@11957.4]
  wire [11:0] _T_63018; // @[Modules.scala 78:156:@11959.4]
  wire [10:0] _T_63019; // @[Modules.scala 78:156:@11960.4]
  wire [10:0] buffer_4_770; // @[Modules.scala 78:156:@11961.4]
  wire [11:0] _T_63021; // @[Modules.scala 78:156:@11963.4]
  wire [10:0] _T_63022; // @[Modules.scala 78:156:@11964.4]
  wire [10:0] buffer_4_771; // @[Modules.scala 78:156:@11965.4]
  wire [11:0] _T_63024; // @[Modules.scala 78:156:@11967.4]
  wire [10:0] _T_63025; // @[Modules.scala 78:156:@11968.4]
  wire [10:0] buffer_4_772; // @[Modules.scala 78:156:@11969.4]
  wire [11:0] _T_63027; // @[Modules.scala 78:156:@11971.4]
  wire [10:0] _T_63028; // @[Modules.scala 78:156:@11972.4]
  wire [10:0] buffer_4_773; // @[Modules.scala 78:156:@11973.4]
  wire [11:0] _T_63030; // @[Modules.scala 78:156:@11975.4]
  wire [10:0] _T_63031; // @[Modules.scala 78:156:@11976.4]
  wire [10:0] buffer_4_774; // @[Modules.scala 78:156:@11977.4]
  wire [11:0] _T_63033; // @[Modules.scala 78:156:@11979.4]
  wire [10:0] _T_63034; // @[Modules.scala 78:156:@11980.4]
  wire [10:0] buffer_4_775; // @[Modules.scala 78:156:@11981.4]
  wire [11:0] _T_63036; // @[Modules.scala 78:156:@11983.4]
  wire [10:0] _T_63037; // @[Modules.scala 78:156:@11984.4]
  wire [10:0] buffer_4_776; // @[Modules.scala 78:156:@11985.4]
  wire [11:0] _T_63039; // @[Modules.scala 78:156:@11987.4]
  wire [10:0] _T_63040; // @[Modules.scala 78:156:@11988.4]
  wire [10:0] buffer_4_777; // @[Modules.scala 78:156:@11989.4]
  wire [11:0] _T_63042; // @[Modules.scala 78:156:@11991.4]
  wire [10:0] _T_63043; // @[Modules.scala 78:156:@11992.4]
  wire [10:0] buffer_4_778; // @[Modules.scala 78:156:@11993.4]
  wire [11:0] _T_63045; // @[Modules.scala 78:156:@11995.4]
  wire [10:0] _T_63046; // @[Modules.scala 78:156:@11996.4]
  wire [10:0] buffer_4_779; // @[Modules.scala 78:156:@11997.4]
  wire [11:0] _T_63048; // @[Modules.scala 78:156:@11999.4]
  wire [10:0] _T_63049; // @[Modules.scala 78:156:@12000.4]
  wire [10:0] buffer_4_780; // @[Modules.scala 78:156:@12001.4]
  wire [11:0] _T_63051; // @[Modules.scala 78:156:@12003.4]
  wire [10:0] _T_63052; // @[Modules.scala 78:156:@12004.4]
  wire [10:0] buffer_4_781; // @[Modules.scala 78:156:@12005.4]
  wire [11:0] _T_63054; // @[Modules.scala 78:156:@12007.4]
  wire [10:0] _T_63055; // @[Modules.scala 78:156:@12008.4]
  wire [10:0] buffer_4_782; // @[Modules.scala 78:156:@12009.4]
  wire [11:0] _T_63057; // @[Modules.scala 78:156:@12011.4]
  wire [10:0] _T_63058; // @[Modules.scala 78:156:@12012.4]
  wire [10:0] buffer_4_783; // @[Modules.scala 78:156:@12013.4]
  wire [5:0] _T_63098; // @[Modules.scala 37:46:@12076.4]
  wire [4:0] _T_63099; // @[Modules.scala 37:46:@12077.4]
  wire [4:0] _T_63100; // @[Modules.scala 37:46:@12078.4]
  wire [5:0] _T_63118; // @[Modules.scala 37:46:@12107.4]
  wire [4:0] _T_63119; // @[Modules.scala 37:46:@12108.4]
  wire [4:0] _T_63120; // @[Modules.scala 37:46:@12109.4]
  wire [5:0] _T_63141; // @[Modules.scala 37:46:@12141.4]
  wire [4:0] _T_63142; // @[Modules.scala 37:46:@12142.4]
  wire [4:0] _T_63143; // @[Modules.scala 37:46:@12143.4]
  wire [5:0] _T_63177; // @[Modules.scala 37:46:@12194.4]
  wire [4:0] _T_63178; // @[Modules.scala 37:46:@12195.4]
  wire [4:0] _T_63179; // @[Modules.scala 37:46:@12196.4]
  wire [5:0] _T_63180; // @[Modules.scala 37:46:@12198.4]
  wire [4:0] _T_63181; // @[Modules.scala 37:46:@12199.4]
  wire [4:0] _T_63182; // @[Modules.scala 37:46:@12200.4]
  wire [5:0] _T_63206; // @[Modules.scala 37:46:@12242.4]
  wire [4:0] _T_63207; // @[Modules.scala 37:46:@12243.4]
  wire [4:0] _T_63208; // @[Modules.scala 37:46:@12244.4]
  wire [5:0] _T_63253; // @[Modules.scala 37:46:@12310.4]
  wire [4:0] _T_63254; // @[Modules.scala 37:46:@12311.4]
  wire [4:0] _T_63255; // @[Modules.scala 37:46:@12312.4]
  wire [5:0] _T_63259; // @[Modules.scala 37:46:@12319.4]
  wire [4:0] _T_63260; // @[Modules.scala 37:46:@12320.4]
  wire [4:0] _T_63261; // @[Modules.scala 37:46:@12321.4]
  wire [5:0] _T_63269; // @[Modules.scala 37:46:@12333.4]
  wire [4:0] _T_63270; // @[Modules.scala 37:46:@12334.4]
  wire [4:0] _T_63271; // @[Modules.scala 37:46:@12335.4]
  wire [5:0] _T_63272; // @[Modules.scala 37:46:@12338.4]
  wire [4:0] _T_63273; // @[Modules.scala 37:46:@12339.4]
  wire [4:0] _T_63274; // @[Modules.scala 37:46:@12340.4]
  wire [5:0] _T_63278; // @[Modules.scala 37:46:@12346.4]
  wire [4:0] _T_63279; // @[Modules.scala 37:46:@12347.4]
  wire [4:0] _T_63280; // @[Modules.scala 37:46:@12348.4]
  wire [5:0] _T_63282; // @[Modules.scala 37:46:@12352.4]
  wire [4:0] _T_63283; // @[Modules.scala 37:46:@12353.4]
  wire [4:0] _T_63284; // @[Modules.scala 37:46:@12354.4]
  wire [5:0] _T_63425; // @[Modules.scala 37:46:@12568.4]
  wire [4:0] _T_63426; // @[Modules.scala 37:46:@12569.4]
  wire [4:0] _T_63427; // @[Modules.scala 37:46:@12570.4]
  wire [5:0] _T_63560; // @[Modules.scala 37:46:@12777.4]
  wire [4:0] _T_63561; // @[Modules.scala 37:46:@12778.4]
  wire [4:0] _T_63562; // @[Modules.scala 37:46:@12779.4]
  wire [5:0] _T_63572; // @[Modules.scala 37:46:@12793.4]
  wire [4:0] _T_63573; // @[Modules.scala 37:46:@12794.4]
  wire [4:0] _T_63574; // @[Modules.scala 37:46:@12795.4]
  wire [5:0] _T_63596; // @[Modules.scala 37:46:@12828.4]
  wire [4:0] _T_63597; // @[Modules.scala 37:46:@12829.4]
  wire [4:0] _T_63598; // @[Modules.scala 37:46:@12830.4]
  wire [11:0] _T_63602; // @[Modules.scala 65:57:@12837.4]
  wire [10:0] _T_63603; // @[Modules.scala 65:57:@12838.4]
  wire [10:0] buffer_5_392; // @[Modules.scala 65:57:@12839.4]
  wire [11:0] _T_63605; // @[Modules.scala 65:57:@12841.4]
  wire [10:0] _T_63606; // @[Modules.scala 65:57:@12842.4]
  wire [10:0] buffer_5_393; // @[Modules.scala 65:57:@12843.4]
  wire [11:0] _T_63608; // @[Modules.scala 65:57:@12845.4]
  wire [10:0] _T_63609; // @[Modules.scala 65:57:@12846.4]
  wire [10:0] buffer_5_394; // @[Modules.scala 65:57:@12847.4]
  wire [10:0] buffer_5_10; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63617; // @[Modules.scala 65:57:@12857.4]
  wire [10:0] _T_63618; // @[Modules.scala 65:57:@12858.4]
  wire [10:0] buffer_5_397; // @[Modules.scala 65:57:@12859.4]
  wire [11:0] _T_63623; // @[Modules.scala 65:57:@12865.4]
  wire [10:0] _T_63624; // @[Modules.scala 65:57:@12866.4]
  wire [10:0] buffer_5_399; // @[Modules.scala 65:57:@12867.4]
  wire [10:0] buffer_5_16; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63626; // @[Modules.scala 65:57:@12869.4]
  wire [10:0] _T_63627; // @[Modules.scala 65:57:@12870.4]
  wire [10:0] buffer_5_400; // @[Modules.scala 65:57:@12871.4]
  wire [10:0] buffer_5_21; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63632; // @[Modules.scala 65:57:@12877.4]
  wire [10:0] _T_63633; // @[Modules.scala 65:57:@12878.4]
  wire [10:0] buffer_5_402; // @[Modules.scala 65:57:@12879.4]
  wire [11:0] _T_63644; // @[Modules.scala 65:57:@12893.4]
  wire [10:0] _T_63645; // @[Modules.scala 65:57:@12894.4]
  wire [10:0] buffer_5_406; // @[Modules.scala 65:57:@12895.4]
  wire [11:0] _T_63653; // @[Modules.scala 65:57:@12905.4]
  wire [10:0] _T_63654; // @[Modules.scala 65:57:@12906.4]
  wire [10:0] buffer_5_409; // @[Modules.scala 65:57:@12907.4]
  wire [10:0] buffer_5_36; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63656; // @[Modules.scala 65:57:@12909.4]
  wire [10:0] _T_63657; // @[Modules.scala 65:57:@12910.4]
  wire [10:0] buffer_5_410; // @[Modules.scala 65:57:@12911.4]
  wire [11:0] _T_63662; // @[Modules.scala 65:57:@12917.4]
  wire [10:0] _T_63663; // @[Modules.scala 65:57:@12918.4]
  wire [10:0] buffer_5_412; // @[Modules.scala 65:57:@12919.4]
  wire [10:0] buffer_5_42; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63665; // @[Modules.scala 65:57:@12921.4]
  wire [10:0] _T_63666; // @[Modules.scala 65:57:@12922.4]
  wire [10:0] buffer_5_413; // @[Modules.scala 65:57:@12923.4]
  wire [11:0] _T_63677; // @[Modules.scala 65:57:@12937.4]
  wire [10:0] _T_63678; // @[Modules.scala 65:57:@12938.4]
  wire [10:0] buffer_5_417; // @[Modules.scala 65:57:@12939.4]
  wire [11:0] _T_63683; // @[Modules.scala 65:57:@12945.4]
  wire [10:0] _T_63684; // @[Modules.scala 65:57:@12946.4]
  wire [10:0] buffer_5_419; // @[Modules.scala 65:57:@12947.4]
  wire [10:0] buffer_5_57; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63686; // @[Modules.scala 65:57:@12949.4]
  wire [10:0] _T_63687; // @[Modules.scala 65:57:@12950.4]
  wire [10:0] buffer_5_420; // @[Modules.scala 65:57:@12951.4]
  wire [10:0] buffer_5_58; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63689; // @[Modules.scala 65:57:@12953.4]
  wire [10:0] _T_63690; // @[Modules.scala 65:57:@12954.4]
  wire [10:0] buffer_5_421; // @[Modules.scala 65:57:@12955.4]
  wire [11:0] _T_63698; // @[Modules.scala 65:57:@12965.4]
  wire [10:0] _T_63699; // @[Modules.scala 65:57:@12966.4]
  wire [10:0] buffer_5_424; // @[Modules.scala 65:57:@12967.4]
  wire [10:0] buffer_5_66; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63701; // @[Modules.scala 65:57:@12969.4]
  wire [10:0] _T_63702; // @[Modules.scala 65:57:@12970.4]
  wire [10:0] buffer_5_425; // @[Modules.scala 65:57:@12971.4]
  wire [10:0] buffer_5_68; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63704; // @[Modules.scala 65:57:@12973.4]
  wire [10:0] _T_63705; // @[Modules.scala 65:57:@12974.4]
  wire [10:0] buffer_5_426; // @[Modules.scala 65:57:@12975.4]
  wire [10:0] buffer_5_71; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63707; // @[Modules.scala 65:57:@12977.4]
  wire [10:0] _T_63708; // @[Modules.scala 65:57:@12978.4]
  wire [10:0] buffer_5_427; // @[Modules.scala 65:57:@12979.4]
  wire [10:0] buffer_5_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63710; // @[Modules.scala 65:57:@12981.4]
  wire [10:0] _T_63711; // @[Modules.scala 65:57:@12982.4]
  wire [10:0] buffer_5_428; // @[Modules.scala 65:57:@12983.4]
  wire [10:0] buffer_5_80; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63722; // @[Modules.scala 65:57:@12997.4]
  wire [10:0] _T_63723; // @[Modules.scala 65:57:@12998.4]
  wire [10:0] buffer_5_432; // @[Modules.scala 65:57:@12999.4]
  wire [10:0] buffer_5_82; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_83; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63725; // @[Modules.scala 65:57:@13001.4]
  wire [10:0] _T_63726; // @[Modules.scala 65:57:@13002.4]
  wire [10:0] buffer_5_433; // @[Modules.scala 65:57:@13003.4]
  wire [11:0] _T_63728; // @[Modules.scala 65:57:@13005.4]
  wire [10:0] _T_63729; // @[Modules.scala 65:57:@13006.4]
  wire [10:0] buffer_5_434; // @[Modules.scala 65:57:@13007.4]
  wire [10:0] buffer_5_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63731; // @[Modules.scala 65:57:@13009.4]
  wire [10:0] _T_63732; // @[Modules.scala 65:57:@13010.4]
  wire [10:0] buffer_5_435; // @[Modules.scala 65:57:@13011.4]
  wire [10:0] buffer_5_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63737; // @[Modules.scala 65:57:@13017.4]
  wire [10:0] _T_63738; // @[Modules.scala 65:57:@13018.4]
  wire [10:0] buffer_5_437; // @[Modules.scala 65:57:@13019.4]
  wire [10:0] buffer_5_92; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63740; // @[Modules.scala 65:57:@13021.4]
  wire [10:0] _T_63741; // @[Modules.scala 65:57:@13022.4]
  wire [10:0] buffer_5_438; // @[Modules.scala 65:57:@13023.4]
  wire [11:0] _T_63743; // @[Modules.scala 65:57:@13025.4]
  wire [10:0] _T_63744; // @[Modules.scala 65:57:@13026.4]
  wire [10:0] buffer_5_439; // @[Modules.scala 65:57:@13027.4]
  wire [11:0] _T_63746; // @[Modules.scala 65:57:@13029.4]
  wire [10:0] _T_63747; // @[Modules.scala 65:57:@13030.4]
  wire [10:0] buffer_5_440; // @[Modules.scala 65:57:@13031.4]
  wire [10:0] buffer_5_101; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63752; // @[Modules.scala 65:57:@13037.4]
  wire [10:0] _T_63753; // @[Modules.scala 65:57:@13038.4]
  wire [10:0] buffer_5_442; // @[Modules.scala 65:57:@13039.4]
  wire [11:0] _T_63755; // @[Modules.scala 65:57:@13041.4]
  wire [10:0] _T_63756; // @[Modules.scala 65:57:@13042.4]
  wire [10:0] buffer_5_443; // @[Modules.scala 65:57:@13043.4]
  wire [11:0] _T_63758; // @[Modules.scala 65:57:@13045.4]
  wire [10:0] _T_63759; // @[Modules.scala 65:57:@13046.4]
  wire [10:0] buffer_5_444; // @[Modules.scala 65:57:@13047.4]
  wire [11:0] _T_63761; // @[Modules.scala 65:57:@13049.4]
  wire [10:0] _T_63762; // @[Modules.scala 65:57:@13050.4]
  wire [10:0] buffer_5_445; // @[Modules.scala 65:57:@13051.4]
  wire [10:0] buffer_5_108; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63764; // @[Modules.scala 65:57:@13053.4]
  wire [10:0] _T_63765; // @[Modules.scala 65:57:@13054.4]
  wire [10:0] buffer_5_446; // @[Modules.scala 65:57:@13055.4]
  wire [10:0] buffer_5_111; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63767; // @[Modules.scala 65:57:@13057.4]
  wire [10:0] _T_63768; // @[Modules.scala 65:57:@13058.4]
  wire [10:0] buffer_5_447; // @[Modules.scala 65:57:@13059.4]
  wire [10:0] buffer_5_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63770; // @[Modules.scala 65:57:@13061.4]
  wire [10:0] _T_63771; // @[Modules.scala 65:57:@13062.4]
  wire [10:0] buffer_5_448; // @[Modules.scala 65:57:@13063.4]
  wire [10:0] buffer_5_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63773; // @[Modules.scala 65:57:@13065.4]
  wire [10:0] _T_63774; // @[Modules.scala 65:57:@13066.4]
  wire [10:0] buffer_5_449; // @[Modules.scala 65:57:@13067.4]
  wire [11:0] _T_63785; // @[Modules.scala 65:57:@13081.4]
  wire [10:0] _T_63786; // @[Modules.scala 65:57:@13082.4]
  wire [10:0] buffer_5_453; // @[Modules.scala 65:57:@13083.4]
  wire [11:0] _T_63788; // @[Modules.scala 65:57:@13085.4]
  wire [10:0] _T_63789; // @[Modules.scala 65:57:@13086.4]
  wire [10:0] buffer_5_454; // @[Modules.scala 65:57:@13087.4]
  wire [10:0] buffer_5_126; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63791; // @[Modules.scala 65:57:@13089.4]
  wire [10:0] _T_63792; // @[Modules.scala 65:57:@13090.4]
  wire [10:0] buffer_5_455; // @[Modules.scala 65:57:@13091.4]
  wire [11:0] _T_63797; // @[Modules.scala 65:57:@13097.4]
  wire [10:0] _T_63798; // @[Modules.scala 65:57:@13098.4]
  wire [10:0] buffer_5_457; // @[Modules.scala 65:57:@13099.4]
  wire [10:0] buffer_5_132; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63800; // @[Modules.scala 65:57:@13101.4]
  wire [10:0] _T_63801; // @[Modules.scala 65:57:@13102.4]
  wire [10:0] buffer_5_458; // @[Modules.scala 65:57:@13103.4]
  wire [10:0] buffer_5_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63803; // @[Modules.scala 65:57:@13105.4]
  wire [10:0] _T_63804; // @[Modules.scala 65:57:@13106.4]
  wire [10:0] buffer_5_459; // @[Modules.scala 65:57:@13107.4]
  wire [10:0] buffer_5_136; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_137; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63806; // @[Modules.scala 65:57:@13109.4]
  wire [10:0] _T_63807; // @[Modules.scala 65:57:@13110.4]
  wire [10:0] buffer_5_460; // @[Modules.scala 65:57:@13111.4]
  wire [10:0] buffer_5_139; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63809; // @[Modules.scala 65:57:@13113.4]
  wire [10:0] _T_63810; // @[Modules.scala 65:57:@13114.4]
  wire [10:0] buffer_5_461; // @[Modules.scala 65:57:@13115.4]
  wire [10:0] buffer_5_140; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63812; // @[Modules.scala 65:57:@13117.4]
  wire [10:0] _T_63813; // @[Modules.scala 65:57:@13118.4]
  wire [10:0] buffer_5_462; // @[Modules.scala 65:57:@13119.4]
  wire [10:0] buffer_5_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63815; // @[Modules.scala 65:57:@13121.4]
  wire [10:0] _T_63816; // @[Modules.scala 65:57:@13122.4]
  wire [10:0] buffer_5_463; // @[Modules.scala 65:57:@13123.4]
  wire [10:0] buffer_5_147; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63821; // @[Modules.scala 65:57:@13129.4]
  wire [10:0] _T_63822; // @[Modules.scala 65:57:@13130.4]
  wire [10:0] buffer_5_465; // @[Modules.scala 65:57:@13131.4]
  wire [10:0] buffer_5_148; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63824; // @[Modules.scala 65:57:@13133.4]
  wire [10:0] _T_63825; // @[Modules.scala 65:57:@13134.4]
  wire [10:0] buffer_5_466; // @[Modules.scala 65:57:@13135.4]
  wire [10:0] buffer_5_150; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_151; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63827; // @[Modules.scala 65:57:@13137.4]
  wire [10:0] _T_63828; // @[Modules.scala 65:57:@13138.4]
  wire [10:0] buffer_5_467; // @[Modules.scala 65:57:@13139.4]
  wire [10:0] buffer_5_153; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63830; // @[Modules.scala 65:57:@13141.4]
  wire [10:0] _T_63831; // @[Modules.scala 65:57:@13142.4]
  wire [10:0] buffer_5_468; // @[Modules.scala 65:57:@13143.4]
  wire [11:0] _T_63833; // @[Modules.scala 65:57:@13145.4]
  wire [10:0] _T_63834; // @[Modules.scala 65:57:@13146.4]
  wire [10:0] buffer_5_469; // @[Modules.scala 65:57:@13147.4]
  wire [10:0] buffer_5_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63842; // @[Modules.scala 65:57:@13157.4]
  wire [10:0] _T_63843; // @[Modules.scala 65:57:@13158.4]
  wire [10:0] buffer_5_472; // @[Modules.scala 65:57:@13159.4]
  wire [10:0] buffer_5_162; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_163; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63845; // @[Modules.scala 65:57:@13161.4]
  wire [10:0] _T_63846; // @[Modules.scala 65:57:@13162.4]
  wire [10:0] buffer_5_473; // @[Modules.scala 65:57:@13163.4]
  wire [10:0] buffer_5_165; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63848; // @[Modules.scala 65:57:@13165.4]
  wire [10:0] _T_63849; // @[Modules.scala 65:57:@13166.4]
  wire [10:0] buffer_5_474; // @[Modules.scala 65:57:@13167.4]
  wire [10:0] buffer_5_168; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63854; // @[Modules.scala 65:57:@13173.4]
  wire [10:0] _T_63855; // @[Modules.scala 65:57:@13174.4]
  wire [10:0] buffer_5_476; // @[Modules.scala 65:57:@13175.4]
  wire [10:0] buffer_5_170; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63857; // @[Modules.scala 65:57:@13177.4]
  wire [10:0] _T_63858; // @[Modules.scala 65:57:@13178.4]
  wire [10:0] buffer_5_477; // @[Modules.scala 65:57:@13179.4]
  wire [11:0] _T_63863; // @[Modules.scala 65:57:@13185.4]
  wire [10:0] _T_63864; // @[Modules.scala 65:57:@13186.4]
  wire [10:0] buffer_5_479; // @[Modules.scala 65:57:@13187.4]
  wire [10:0] buffer_5_177; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63866; // @[Modules.scala 65:57:@13189.4]
  wire [10:0] _T_63867; // @[Modules.scala 65:57:@13190.4]
  wire [10:0] buffer_5_480; // @[Modules.scala 65:57:@13191.4]
  wire [10:0] buffer_5_178; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63869; // @[Modules.scala 65:57:@13193.4]
  wire [10:0] _T_63870; // @[Modules.scala 65:57:@13194.4]
  wire [10:0] buffer_5_481; // @[Modules.scala 65:57:@13195.4]
  wire [10:0] buffer_5_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63875; // @[Modules.scala 65:57:@13201.4]
  wire [10:0] _T_63876; // @[Modules.scala 65:57:@13202.4]
  wire [10:0] buffer_5_483; // @[Modules.scala 65:57:@13203.4]
  wire [10:0] buffer_5_186; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63881; // @[Modules.scala 65:57:@13209.4]
  wire [10:0] _T_63882; // @[Modules.scala 65:57:@13210.4]
  wire [10:0] buffer_5_485; // @[Modules.scala 65:57:@13211.4]
  wire [10:0] buffer_5_188; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63884; // @[Modules.scala 65:57:@13213.4]
  wire [10:0] _T_63885; // @[Modules.scala 65:57:@13214.4]
  wire [10:0] buffer_5_486; // @[Modules.scala 65:57:@13215.4]
  wire [10:0] buffer_5_194; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63893; // @[Modules.scala 65:57:@13225.4]
  wire [10:0] _T_63894; // @[Modules.scala 65:57:@13226.4]
  wire [10:0] buffer_5_489; // @[Modules.scala 65:57:@13227.4]
  wire [10:0] buffer_5_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63896; // @[Modules.scala 65:57:@13229.4]
  wire [10:0] _T_63897; // @[Modules.scala 65:57:@13230.4]
  wire [10:0] buffer_5_490; // @[Modules.scala 65:57:@13231.4]
  wire [11:0] _T_63914; // @[Modules.scala 65:57:@13253.4]
  wire [10:0] _T_63915; // @[Modules.scala 65:57:@13254.4]
  wire [10:0] buffer_5_496; // @[Modules.scala 65:57:@13255.4]
  wire [10:0] buffer_5_211; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63917; // @[Modules.scala 65:57:@13257.4]
  wire [10:0] _T_63918; // @[Modules.scala 65:57:@13258.4]
  wire [10:0] buffer_5_497; // @[Modules.scala 65:57:@13259.4]
  wire [10:0] buffer_5_212; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63920; // @[Modules.scala 65:57:@13261.4]
  wire [10:0] _T_63921; // @[Modules.scala 65:57:@13262.4]
  wire [10:0] buffer_5_498; // @[Modules.scala 65:57:@13263.4]
  wire [10:0] buffer_5_218; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63929; // @[Modules.scala 65:57:@13273.4]
  wire [10:0] _T_63930; // @[Modules.scala 65:57:@13274.4]
  wire [10:0] buffer_5_501; // @[Modules.scala 65:57:@13275.4]
  wire [10:0] buffer_5_222; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63935; // @[Modules.scala 65:57:@13281.4]
  wire [10:0] _T_63936; // @[Modules.scala 65:57:@13282.4]
  wire [10:0] buffer_5_503; // @[Modules.scala 65:57:@13283.4]
  wire [11:0] _T_63941; // @[Modules.scala 65:57:@13289.4]
  wire [10:0] _T_63942; // @[Modules.scala 65:57:@13290.4]
  wire [10:0] buffer_5_505; // @[Modules.scala 65:57:@13291.4]
  wire [10:0] buffer_5_231; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63947; // @[Modules.scala 65:57:@13297.4]
  wire [10:0] _T_63948; // @[Modules.scala 65:57:@13298.4]
  wire [10:0] buffer_5_507; // @[Modules.scala 65:57:@13299.4]
  wire [10:0] buffer_5_232; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63950; // @[Modules.scala 65:57:@13301.4]
  wire [10:0] _T_63951; // @[Modules.scala 65:57:@13302.4]
  wire [10:0] buffer_5_508; // @[Modules.scala 65:57:@13303.4]
  wire [10:0] buffer_5_236; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63956; // @[Modules.scala 65:57:@13309.4]
  wire [10:0] _T_63957; // @[Modules.scala 65:57:@13310.4]
  wire [10:0] buffer_5_510; // @[Modules.scala 65:57:@13311.4]
  wire [11:0] _T_63962; // @[Modules.scala 65:57:@13317.4]
  wire [10:0] _T_63963; // @[Modules.scala 65:57:@13318.4]
  wire [10:0] buffer_5_512; // @[Modules.scala 65:57:@13319.4]
  wire [10:0] buffer_5_242; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63965; // @[Modules.scala 65:57:@13321.4]
  wire [10:0] _T_63966; // @[Modules.scala 65:57:@13322.4]
  wire [10:0] buffer_5_513; // @[Modules.scala 65:57:@13323.4]
  wire [11:0] _T_63971; // @[Modules.scala 65:57:@13329.4]
  wire [10:0] _T_63972; // @[Modules.scala 65:57:@13330.4]
  wire [10:0] buffer_5_515; // @[Modules.scala 65:57:@13331.4]
  wire [10:0] buffer_5_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63983; // @[Modules.scala 65:57:@13345.4]
  wire [10:0] _T_63984; // @[Modules.scala 65:57:@13346.4]
  wire [10:0] buffer_5_519; // @[Modules.scala 65:57:@13347.4]
  wire [10:0] buffer_5_256; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_63986; // @[Modules.scala 65:57:@13349.4]
  wire [10:0] _T_63987; // @[Modules.scala 65:57:@13350.4]
  wire [10:0] buffer_5_520; // @[Modules.scala 65:57:@13351.4]
  wire [11:0] _T_63989; // @[Modules.scala 65:57:@13353.4]
  wire [10:0] _T_63990; // @[Modules.scala 65:57:@13354.4]
  wire [10:0] buffer_5_521; // @[Modules.scala 65:57:@13355.4]
  wire [11:0] _T_63992; // @[Modules.scala 65:57:@13357.4]
  wire [10:0] _T_63993; // @[Modules.scala 65:57:@13358.4]
  wire [10:0] buffer_5_522; // @[Modules.scala 65:57:@13359.4]
  wire [10:0] buffer_5_268; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64004; // @[Modules.scala 65:57:@13373.4]
  wire [10:0] _T_64005; // @[Modules.scala 65:57:@13374.4]
  wire [10:0] buffer_5_526; // @[Modules.scala 65:57:@13375.4]
  wire [10:0] buffer_5_270; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64007; // @[Modules.scala 65:57:@13377.4]
  wire [10:0] _T_64008; // @[Modules.scala 65:57:@13378.4]
  wire [10:0] buffer_5_527; // @[Modules.scala 65:57:@13379.4]
  wire [11:0] _T_64010; // @[Modules.scala 65:57:@13381.4]
  wire [10:0] _T_64011; // @[Modules.scala 65:57:@13382.4]
  wire [10:0] buffer_5_528; // @[Modules.scala 65:57:@13383.4]
  wire [11:0] _T_64013; // @[Modules.scala 65:57:@13385.4]
  wire [10:0] _T_64014; // @[Modules.scala 65:57:@13386.4]
  wire [10:0] buffer_5_529; // @[Modules.scala 65:57:@13387.4]
  wire [10:0] buffer_5_277; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64016; // @[Modules.scala 65:57:@13389.4]
  wire [10:0] _T_64017; // @[Modules.scala 65:57:@13390.4]
  wire [10:0] buffer_5_530; // @[Modules.scala 65:57:@13391.4]
  wire [10:0] buffer_5_279; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64019; // @[Modules.scala 65:57:@13393.4]
  wire [10:0] _T_64020; // @[Modules.scala 65:57:@13394.4]
  wire [10:0] buffer_5_531; // @[Modules.scala 65:57:@13395.4]
  wire [10:0] buffer_5_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64022; // @[Modules.scala 65:57:@13397.4]
  wire [10:0] _T_64023; // @[Modules.scala 65:57:@13398.4]
  wire [10:0] buffer_5_532; // @[Modules.scala 65:57:@13399.4]
  wire [10:0] buffer_5_282; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64025; // @[Modules.scala 65:57:@13401.4]
  wire [10:0] _T_64026; // @[Modules.scala 65:57:@13402.4]
  wire [10:0] buffer_5_533; // @[Modules.scala 65:57:@13403.4]
  wire [10:0] buffer_5_289; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64034; // @[Modules.scala 65:57:@13413.4]
  wire [10:0] _T_64035; // @[Modules.scala 65:57:@13414.4]
  wire [10:0] buffer_5_536; // @[Modules.scala 65:57:@13415.4]
  wire [10:0] buffer_5_290; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_291; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64037; // @[Modules.scala 65:57:@13417.4]
  wire [10:0] _T_64038; // @[Modules.scala 65:57:@13418.4]
  wire [10:0] buffer_5_537; // @[Modules.scala 65:57:@13419.4]
  wire [11:0] _T_64049; // @[Modules.scala 65:57:@13433.4]
  wire [10:0] _T_64050; // @[Modules.scala 65:57:@13434.4]
  wire [10:0] buffer_5_541; // @[Modules.scala 65:57:@13435.4]
  wire [10:0] buffer_5_302; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64055; // @[Modules.scala 65:57:@13441.4]
  wire [10:0] _T_64056; // @[Modules.scala 65:57:@13442.4]
  wire [10:0] buffer_5_543; // @[Modules.scala 65:57:@13443.4]
  wire [10:0] buffer_5_313; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64070; // @[Modules.scala 65:57:@13461.4]
  wire [10:0] _T_64071; // @[Modules.scala 65:57:@13462.4]
  wire [10:0] buffer_5_548; // @[Modules.scala 65:57:@13463.4]
  wire [10:0] buffer_5_314; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64073; // @[Modules.scala 65:57:@13465.4]
  wire [10:0] _T_64074; // @[Modules.scala 65:57:@13466.4]
  wire [10:0] buffer_5_549; // @[Modules.scala 65:57:@13467.4]
  wire [11:0] _T_64076; // @[Modules.scala 65:57:@13469.4]
  wire [10:0] _T_64077; // @[Modules.scala 65:57:@13470.4]
  wire [10:0] buffer_5_550; // @[Modules.scala 65:57:@13471.4]
  wire [10:0] buffer_5_320; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64082; // @[Modules.scala 65:57:@13477.4]
  wire [10:0] _T_64083; // @[Modules.scala 65:57:@13478.4]
  wire [10:0] buffer_5_552; // @[Modules.scala 65:57:@13479.4]
  wire [11:0] _T_64088; // @[Modules.scala 65:57:@13485.4]
  wire [10:0] _T_64089; // @[Modules.scala 65:57:@13486.4]
  wire [10:0] buffer_5_554; // @[Modules.scala 65:57:@13487.4]
  wire [10:0] buffer_5_326; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64091; // @[Modules.scala 65:57:@13489.4]
  wire [10:0] _T_64092; // @[Modules.scala 65:57:@13490.4]
  wire [10:0] buffer_5_555; // @[Modules.scala 65:57:@13491.4]
  wire [10:0] buffer_5_328; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64094; // @[Modules.scala 65:57:@13493.4]
  wire [10:0] _T_64095; // @[Modules.scala 65:57:@13494.4]
  wire [10:0] buffer_5_556; // @[Modules.scala 65:57:@13495.4]
  wire [11:0] _T_64097; // @[Modules.scala 65:57:@13497.4]
  wire [10:0] _T_64098; // @[Modules.scala 65:57:@13498.4]
  wire [10:0] buffer_5_557; // @[Modules.scala 65:57:@13499.4]
  wire [10:0] buffer_5_332; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64100; // @[Modules.scala 65:57:@13501.4]
  wire [10:0] _T_64101; // @[Modules.scala 65:57:@13502.4]
  wire [10:0] buffer_5_558; // @[Modules.scala 65:57:@13503.4]
  wire [11:0] _T_64106; // @[Modules.scala 65:57:@13509.4]
  wire [10:0] _T_64107; // @[Modules.scala 65:57:@13510.4]
  wire [10:0] buffer_5_560; // @[Modules.scala 65:57:@13511.4]
  wire [10:0] buffer_5_339; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64109; // @[Modules.scala 65:57:@13513.4]
  wire [10:0] _T_64110; // @[Modules.scala 65:57:@13514.4]
  wire [10:0] buffer_5_561; // @[Modules.scala 65:57:@13515.4]
  wire [10:0] buffer_5_340; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_5_341; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64112; // @[Modules.scala 65:57:@13517.4]
  wire [10:0] _T_64113; // @[Modules.scala 65:57:@13518.4]
  wire [10:0] buffer_5_562; // @[Modules.scala 65:57:@13519.4]
  wire [10:0] buffer_5_343; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64115; // @[Modules.scala 65:57:@13521.4]
  wire [10:0] _T_64116; // @[Modules.scala 65:57:@13522.4]
  wire [10:0] buffer_5_563; // @[Modules.scala 65:57:@13523.4]
  wire [11:0] _T_64124; // @[Modules.scala 65:57:@13533.4]
  wire [10:0] _T_64125; // @[Modules.scala 65:57:@13534.4]
  wire [10:0] buffer_5_566; // @[Modules.scala 65:57:@13535.4]
  wire [10:0] buffer_5_350; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64127; // @[Modules.scala 65:57:@13537.4]
  wire [10:0] _T_64128; // @[Modules.scala 65:57:@13538.4]
  wire [10:0] buffer_5_567; // @[Modules.scala 65:57:@13539.4]
  wire [10:0] buffer_5_352; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64130; // @[Modules.scala 65:57:@13541.4]
  wire [10:0] _T_64131; // @[Modules.scala 65:57:@13542.4]
  wire [10:0] buffer_5_568; // @[Modules.scala 65:57:@13543.4]
  wire [10:0] buffer_5_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64142; // @[Modules.scala 65:57:@13557.4]
  wire [10:0] _T_64143; // @[Modules.scala 65:57:@13558.4]
  wire [10:0] buffer_5_572; // @[Modules.scala 65:57:@13559.4]
  wire [10:0] buffer_5_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64151; // @[Modules.scala 65:57:@13569.4]
  wire [10:0] _T_64152; // @[Modules.scala 65:57:@13570.4]
  wire [10:0] buffer_5_575; // @[Modules.scala 65:57:@13571.4]
  wire [10:0] buffer_5_371; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64157; // @[Modules.scala 65:57:@13577.4]
  wire [10:0] _T_64158; // @[Modules.scala 65:57:@13578.4]
  wire [10:0] buffer_5_577; // @[Modules.scala 65:57:@13579.4]
  wire [10:0] buffer_5_375; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64163; // @[Modules.scala 65:57:@13585.4]
  wire [10:0] _T_64164; // @[Modules.scala 65:57:@13586.4]
  wire [10:0] buffer_5_579; // @[Modules.scala 65:57:@13587.4]
  wire [10:0] buffer_5_383; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64175; // @[Modules.scala 65:57:@13601.4]
  wire [10:0] _T_64176; // @[Modules.scala 65:57:@13602.4]
  wire [10:0] buffer_5_583; // @[Modules.scala 65:57:@13603.4]
  wire [10:0] buffer_5_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_64184; // @[Modules.scala 65:57:@13613.4]
  wire [10:0] _T_64185; // @[Modules.scala 65:57:@13614.4]
  wire [10:0] buffer_5_586; // @[Modules.scala 65:57:@13615.4]
  wire [11:0] _T_64190; // @[Modules.scala 68:83:@13621.4]
  wire [10:0] _T_64191; // @[Modules.scala 68:83:@13622.4]
  wire [10:0] buffer_5_588; // @[Modules.scala 68:83:@13623.4]
  wire [11:0] _T_64193; // @[Modules.scala 68:83:@13625.4]
  wire [10:0] _T_64194; // @[Modules.scala 68:83:@13626.4]
  wire [10:0] buffer_5_589; // @[Modules.scala 68:83:@13627.4]
  wire [11:0] _T_64196; // @[Modules.scala 68:83:@13629.4]
  wire [10:0] _T_64197; // @[Modules.scala 68:83:@13630.4]
  wire [10:0] buffer_5_590; // @[Modules.scala 68:83:@13631.4]
  wire [11:0] _T_64199; // @[Modules.scala 68:83:@13633.4]
  wire [10:0] _T_64200; // @[Modules.scala 68:83:@13634.4]
  wire [10:0] buffer_5_591; // @[Modules.scala 68:83:@13635.4]
  wire [11:0] _T_64202; // @[Modules.scala 68:83:@13637.4]
  wire [10:0] _T_64203; // @[Modules.scala 68:83:@13638.4]
  wire [10:0] buffer_5_592; // @[Modules.scala 68:83:@13639.4]
  wire [11:0] _T_64205; // @[Modules.scala 68:83:@13641.4]
  wire [10:0] _T_64206; // @[Modules.scala 68:83:@13642.4]
  wire [10:0] buffer_5_593; // @[Modules.scala 68:83:@13643.4]
  wire [11:0] _T_64208; // @[Modules.scala 68:83:@13645.4]
  wire [10:0] _T_64209; // @[Modules.scala 68:83:@13646.4]
  wire [10:0] buffer_5_594; // @[Modules.scala 68:83:@13647.4]
  wire [11:0] _T_64211; // @[Modules.scala 68:83:@13649.4]
  wire [10:0] _T_64212; // @[Modules.scala 68:83:@13650.4]
  wire [10:0] buffer_5_595; // @[Modules.scala 68:83:@13651.4]
  wire [11:0] _T_64214; // @[Modules.scala 68:83:@13653.4]
  wire [10:0] _T_64215; // @[Modules.scala 68:83:@13654.4]
  wire [10:0] buffer_5_596; // @[Modules.scala 68:83:@13655.4]
  wire [11:0] _T_64217; // @[Modules.scala 68:83:@13657.4]
  wire [10:0] _T_64218; // @[Modules.scala 68:83:@13658.4]
  wire [10:0] buffer_5_597; // @[Modules.scala 68:83:@13659.4]
  wire [11:0] _T_64220; // @[Modules.scala 68:83:@13661.4]
  wire [10:0] _T_64221; // @[Modules.scala 68:83:@13662.4]
  wire [10:0] buffer_5_598; // @[Modules.scala 68:83:@13663.4]
  wire [11:0] _T_64226; // @[Modules.scala 68:83:@13669.4]
  wire [10:0] _T_64227; // @[Modules.scala 68:83:@13670.4]
  wire [10:0] buffer_5_600; // @[Modules.scala 68:83:@13671.4]
  wire [11:0] _T_64229; // @[Modules.scala 68:83:@13673.4]
  wire [10:0] _T_64230; // @[Modules.scala 68:83:@13674.4]
  wire [10:0] buffer_5_601; // @[Modules.scala 68:83:@13675.4]
  wire [11:0] _T_64232; // @[Modules.scala 68:83:@13677.4]
  wire [10:0] _T_64233; // @[Modules.scala 68:83:@13678.4]
  wire [10:0] buffer_5_602; // @[Modules.scala 68:83:@13679.4]
  wire [11:0] _T_64238; // @[Modules.scala 68:83:@13685.4]
  wire [10:0] _T_64239; // @[Modules.scala 68:83:@13686.4]
  wire [10:0] buffer_5_604; // @[Modules.scala 68:83:@13687.4]
  wire [11:0] _T_64241; // @[Modules.scala 68:83:@13689.4]
  wire [10:0] _T_64242; // @[Modules.scala 68:83:@13690.4]
  wire [10:0] buffer_5_605; // @[Modules.scala 68:83:@13691.4]
  wire [11:0] _T_64244; // @[Modules.scala 68:83:@13693.4]
  wire [10:0] _T_64245; // @[Modules.scala 68:83:@13694.4]
  wire [10:0] buffer_5_606; // @[Modules.scala 68:83:@13695.4]
  wire [11:0] _T_64247; // @[Modules.scala 68:83:@13697.4]
  wire [10:0] _T_64248; // @[Modules.scala 68:83:@13698.4]
  wire [10:0] buffer_5_607; // @[Modules.scala 68:83:@13699.4]
  wire [11:0] _T_64250; // @[Modules.scala 68:83:@13701.4]
  wire [10:0] _T_64251; // @[Modules.scala 68:83:@13702.4]
  wire [10:0] buffer_5_608; // @[Modules.scala 68:83:@13703.4]
  wire [11:0] _T_64253; // @[Modules.scala 68:83:@13705.4]
  wire [10:0] _T_64254; // @[Modules.scala 68:83:@13706.4]
  wire [10:0] buffer_5_609; // @[Modules.scala 68:83:@13707.4]
  wire [11:0] _T_64256; // @[Modules.scala 68:83:@13709.4]
  wire [10:0] _T_64257; // @[Modules.scala 68:83:@13710.4]
  wire [10:0] buffer_5_610; // @[Modules.scala 68:83:@13711.4]
  wire [11:0] _T_64259; // @[Modules.scala 68:83:@13713.4]
  wire [10:0] _T_64260; // @[Modules.scala 68:83:@13714.4]
  wire [10:0] buffer_5_611; // @[Modules.scala 68:83:@13715.4]
  wire [11:0] _T_64262; // @[Modules.scala 68:83:@13717.4]
  wire [10:0] _T_64263; // @[Modules.scala 68:83:@13718.4]
  wire [10:0] buffer_5_612; // @[Modules.scala 68:83:@13719.4]
  wire [11:0] _T_64265; // @[Modules.scala 68:83:@13721.4]
  wire [10:0] _T_64266; // @[Modules.scala 68:83:@13722.4]
  wire [10:0] buffer_5_613; // @[Modules.scala 68:83:@13723.4]
  wire [11:0] _T_64268; // @[Modules.scala 68:83:@13725.4]
  wire [10:0] _T_64269; // @[Modules.scala 68:83:@13726.4]
  wire [10:0] buffer_5_614; // @[Modules.scala 68:83:@13727.4]
  wire [11:0] _T_64271; // @[Modules.scala 68:83:@13729.4]
  wire [10:0] _T_64272; // @[Modules.scala 68:83:@13730.4]
  wire [10:0] buffer_5_615; // @[Modules.scala 68:83:@13731.4]
  wire [11:0] _T_64274; // @[Modules.scala 68:83:@13733.4]
  wire [10:0] _T_64275; // @[Modules.scala 68:83:@13734.4]
  wire [10:0] buffer_5_616; // @[Modules.scala 68:83:@13735.4]
  wire [11:0] _T_64277; // @[Modules.scala 68:83:@13737.4]
  wire [10:0] _T_64278; // @[Modules.scala 68:83:@13738.4]
  wire [10:0] buffer_5_617; // @[Modules.scala 68:83:@13739.4]
  wire [11:0] _T_64280; // @[Modules.scala 68:83:@13741.4]
  wire [10:0] _T_64281; // @[Modules.scala 68:83:@13742.4]
  wire [10:0] buffer_5_618; // @[Modules.scala 68:83:@13743.4]
  wire [11:0] _T_64283; // @[Modules.scala 68:83:@13745.4]
  wire [10:0] _T_64284; // @[Modules.scala 68:83:@13746.4]
  wire [10:0] buffer_5_619; // @[Modules.scala 68:83:@13747.4]
  wire [11:0] _T_64286; // @[Modules.scala 68:83:@13749.4]
  wire [10:0] _T_64287; // @[Modules.scala 68:83:@13750.4]
  wire [10:0] buffer_5_620; // @[Modules.scala 68:83:@13751.4]
  wire [11:0] _T_64289; // @[Modules.scala 68:83:@13753.4]
  wire [10:0] _T_64290; // @[Modules.scala 68:83:@13754.4]
  wire [10:0] buffer_5_621; // @[Modules.scala 68:83:@13755.4]
  wire [11:0] _T_64292; // @[Modules.scala 68:83:@13757.4]
  wire [10:0] _T_64293; // @[Modules.scala 68:83:@13758.4]
  wire [10:0] buffer_5_622; // @[Modules.scala 68:83:@13759.4]
  wire [11:0] _T_64295; // @[Modules.scala 68:83:@13761.4]
  wire [10:0] _T_64296; // @[Modules.scala 68:83:@13762.4]
  wire [10:0] buffer_5_623; // @[Modules.scala 68:83:@13763.4]
  wire [11:0] _T_64298; // @[Modules.scala 68:83:@13765.4]
  wire [10:0] _T_64299; // @[Modules.scala 68:83:@13766.4]
  wire [10:0] buffer_5_624; // @[Modules.scala 68:83:@13767.4]
  wire [11:0] _T_64301; // @[Modules.scala 68:83:@13769.4]
  wire [10:0] _T_64302; // @[Modules.scala 68:83:@13770.4]
  wire [10:0] buffer_5_625; // @[Modules.scala 68:83:@13771.4]
  wire [11:0] _T_64304; // @[Modules.scala 68:83:@13773.4]
  wire [10:0] _T_64305; // @[Modules.scala 68:83:@13774.4]
  wire [10:0] buffer_5_626; // @[Modules.scala 68:83:@13775.4]
  wire [11:0] _T_64310; // @[Modules.scala 68:83:@13781.4]
  wire [10:0] _T_64311; // @[Modules.scala 68:83:@13782.4]
  wire [10:0] buffer_5_628; // @[Modules.scala 68:83:@13783.4]
  wire [11:0] _T_64313; // @[Modules.scala 68:83:@13785.4]
  wire [10:0] _T_64314; // @[Modules.scala 68:83:@13786.4]
  wire [10:0] buffer_5_629; // @[Modules.scala 68:83:@13787.4]
  wire [11:0] _T_64316; // @[Modules.scala 68:83:@13789.4]
  wire [10:0] _T_64317; // @[Modules.scala 68:83:@13790.4]
  wire [10:0] buffer_5_630; // @[Modules.scala 68:83:@13791.4]
  wire [11:0] _T_64319; // @[Modules.scala 68:83:@13793.4]
  wire [10:0] _T_64320; // @[Modules.scala 68:83:@13794.4]
  wire [10:0] buffer_5_631; // @[Modules.scala 68:83:@13795.4]
  wire [11:0] _T_64322; // @[Modules.scala 68:83:@13797.4]
  wire [10:0] _T_64323; // @[Modules.scala 68:83:@13798.4]
  wire [10:0] buffer_5_632; // @[Modules.scala 68:83:@13799.4]
  wire [11:0] _T_64325; // @[Modules.scala 68:83:@13801.4]
  wire [10:0] _T_64326; // @[Modules.scala 68:83:@13802.4]
  wire [10:0] buffer_5_633; // @[Modules.scala 68:83:@13803.4]
  wire [11:0] _T_64328; // @[Modules.scala 68:83:@13805.4]
  wire [10:0] _T_64329; // @[Modules.scala 68:83:@13806.4]
  wire [10:0] buffer_5_634; // @[Modules.scala 68:83:@13807.4]
  wire [11:0] _T_64331; // @[Modules.scala 68:83:@13809.4]
  wire [10:0] _T_64332; // @[Modules.scala 68:83:@13810.4]
  wire [10:0] buffer_5_635; // @[Modules.scala 68:83:@13811.4]
  wire [11:0] _T_64334; // @[Modules.scala 68:83:@13813.4]
  wire [10:0] _T_64335; // @[Modules.scala 68:83:@13814.4]
  wire [10:0] buffer_5_636; // @[Modules.scala 68:83:@13815.4]
  wire [11:0] _T_64337; // @[Modules.scala 68:83:@13817.4]
  wire [10:0] _T_64338; // @[Modules.scala 68:83:@13818.4]
  wire [10:0] buffer_5_637; // @[Modules.scala 68:83:@13819.4]
  wire [11:0] _T_64340; // @[Modules.scala 68:83:@13821.4]
  wire [10:0] _T_64341; // @[Modules.scala 68:83:@13822.4]
  wire [10:0] buffer_5_638; // @[Modules.scala 68:83:@13823.4]
  wire [11:0] _T_64343; // @[Modules.scala 68:83:@13825.4]
  wire [10:0] _T_64344; // @[Modules.scala 68:83:@13826.4]
  wire [10:0] buffer_5_639; // @[Modules.scala 68:83:@13827.4]
  wire [11:0] _T_64346; // @[Modules.scala 68:83:@13829.4]
  wire [10:0] _T_64347; // @[Modules.scala 68:83:@13830.4]
  wire [10:0] buffer_5_640; // @[Modules.scala 68:83:@13831.4]
  wire [11:0] _T_64349; // @[Modules.scala 68:83:@13833.4]
  wire [10:0] _T_64350; // @[Modules.scala 68:83:@13834.4]
  wire [10:0] buffer_5_641; // @[Modules.scala 68:83:@13835.4]
  wire [11:0] _T_64352; // @[Modules.scala 68:83:@13837.4]
  wire [10:0] _T_64353; // @[Modules.scala 68:83:@13838.4]
  wire [10:0] buffer_5_642; // @[Modules.scala 68:83:@13839.4]
  wire [11:0] _T_64355; // @[Modules.scala 68:83:@13841.4]
  wire [10:0] _T_64356; // @[Modules.scala 68:83:@13842.4]
  wire [10:0] buffer_5_643; // @[Modules.scala 68:83:@13843.4]
  wire [11:0] _T_64358; // @[Modules.scala 68:83:@13845.4]
  wire [10:0] _T_64359; // @[Modules.scala 68:83:@13846.4]
  wire [10:0] buffer_5_644; // @[Modules.scala 68:83:@13847.4]
  wire [11:0] _T_64361; // @[Modules.scala 68:83:@13849.4]
  wire [10:0] _T_64362; // @[Modules.scala 68:83:@13850.4]
  wire [10:0] buffer_5_645; // @[Modules.scala 68:83:@13851.4]
  wire [11:0] _T_64364; // @[Modules.scala 68:83:@13853.4]
  wire [10:0] _T_64365; // @[Modules.scala 68:83:@13854.4]
  wire [10:0] buffer_5_646; // @[Modules.scala 68:83:@13855.4]
  wire [11:0] _T_64367; // @[Modules.scala 68:83:@13857.4]
  wire [10:0] _T_64368; // @[Modules.scala 68:83:@13858.4]
  wire [10:0] buffer_5_647; // @[Modules.scala 68:83:@13859.4]
  wire [11:0] _T_64370; // @[Modules.scala 68:83:@13861.4]
  wire [10:0] _T_64371; // @[Modules.scala 68:83:@13862.4]
  wire [10:0] buffer_5_648; // @[Modules.scala 68:83:@13863.4]
  wire [11:0] _T_64373; // @[Modules.scala 68:83:@13865.4]
  wire [10:0] _T_64374; // @[Modules.scala 68:83:@13866.4]
  wire [10:0] buffer_5_649; // @[Modules.scala 68:83:@13867.4]
  wire [11:0] _T_64376; // @[Modules.scala 68:83:@13869.4]
  wire [10:0] _T_64377; // @[Modules.scala 68:83:@13870.4]
  wire [10:0] buffer_5_650; // @[Modules.scala 68:83:@13871.4]
  wire [11:0] _T_64379; // @[Modules.scala 68:83:@13873.4]
  wire [10:0] _T_64380; // @[Modules.scala 68:83:@13874.4]
  wire [10:0] buffer_5_651; // @[Modules.scala 68:83:@13875.4]
  wire [11:0] _T_64382; // @[Modules.scala 68:83:@13877.4]
  wire [10:0] _T_64383; // @[Modules.scala 68:83:@13878.4]
  wire [10:0] buffer_5_652; // @[Modules.scala 68:83:@13879.4]
  wire [11:0] _T_64385; // @[Modules.scala 68:83:@13881.4]
  wire [10:0] _T_64386; // @[Modules.scala 68:83:@13882.4]
  wire [10:0] buffer_5_653; // @[Modules.scala 68:83:@13883.4]
  wire [11:0] _T_64388; // @[Modules.scala 68:83:@13885.4]
  wire [10:0] _T_64389; // @[Modules.scala 68:83:@13886.4]
  wire [10:0] buffer_5_654; // @[Modules.scala 68:83:@13887.4]
  wire [11:0] _T_64391; // @[Modules.scala 68:83:@13889.4]
  wire [10:0] _T_64392; // @[Modules.scala 68:83:@13890.4]
  wire [10:0] buffer_5_655; // @[Modules.scala 68:83:@13891.4]
  wire [11:0] _T_64394; // @[Modules.scala 68:83:@13893.4]
  wire [10:0] _T_64395; // @[Modules.scala 68:83:@13894.4]
  wire [10:0] buffer_5_656; // @[Modules.scala 68:83:@13895.4]
  wire [11:0] _T_64397; // @[Modules.scala 68:83:@13897.4]
  wire [10:0] _T_64398; // @[Modules.scala 68:83:@13898.4]
  wire [10:0] buffer_5_657; // @[Modules.scala 68:83:@13899.4]
  wire [11:0] _T_64400; // @[Modules.scala 68:83:@13901.4]
  wire [10:0] _T_64401; // @[Modules.scala 68:83:@13902.4]
  wire [10:0] buffer_5_658; // @[Modules.scala 68:83:@13903.4]
  wire [11:0] _T_64406; // @[Modules.scala 68:83:@13909.4]
  wire [10:0] _T_64407; // @[Modules.scala 68:83:@13910.4]
  wire [10:0] buffer_5_660; // @[Modules.scala 68:83:@13911.4]
  wire [11:0] _T_64409; // @[Modules.scala 68:83:@13913.4]
  wire [10:0] _T_64410; // @[Modules.scala 68:83:@13914.4]
  wire [10:0] buffer_5_661; // @[Modules.scala 68:83:@13915.4]
  wire [11:0] _T_64412; // @[Modules.scala 68:83:@13917.4]
  wire [10:0] _T_64413; // @[Modules.scala 68:83:@13918.4]
  wire [10:0] buffer_5_662; // @[Modules.scala 68:83:@13919.4]
  wire [11:0] _T_64415; // @[Modules.scala 68:83:@13921.4]
  wire [10:0] _T_64416; // @[Modules.scala 68:83:@13922.4]
  wire [10:0] buffer_5_663; // @[Modules.scala 68:83:@13923.4]
  wire [11:0] _T_64418; // @[Modules.scala 68:83:@13925.4]
  wire [10:0] _T_64419; // @[Modules.scala 68:83:@13926.4]
  wire [10:0] buffer_5_664; // @[Modules.scala 68:83:@13927.4]
  wire [11:0] _T_64421; // @[Modules.scala 68:83:@13929.4]
  wire [10:0] _T_64422; // @[Modules.scala 68:83:@13930.4]
  wire [10:0] buffer_5_665; // @[Modules.scala 68:83:@13931.4]
  wire [11:0] _T_64424; // @[Modules.scala 68:83:@13933.4]
  wire [10:0] _T_64425; // @[Modules.scala 68:83:@13934.4]
  wire [10:0] buffer_5_666; // @[Modules.scala 68:83:@13935.4]
  wire [11:0] _T_64427; // @[Modules.scala 68:83:@13937.4]
  wire [10:0] _T_64428; // @[Modules.scala 68:83:@13938.4]
  wire [10:0] buffer_5_667; // @[Modules.scala 68:83:@13939.4]
  wire [11:0] _T_64430; // @[Modules.scala 68:83:@13941.4]
  wire [10:0] _T_64431; // @[Modules.scala 68:83:@13942.4]
  wire [10:0] buffer_5_668; // @[Modules.scala 68:83:@13943.4]
  wire [11:0] _T_64433; // @[Modules.scala 68:83:@13945.4]
  wire [10:0] _T_64434; // @[Modules.scala 68:83:@13946.4]
  wire [10:0] buffer_5_669; // @[Modules.scala 68:83:@13947.4]
  wire [11:0] _T_64436; // @[Modules.scala 68:83:@13949.4]
  wire [10:0] _T_64437; // @[Modules.scala 68:83:@13950.4]
  wire [10:0] buffer_5_670; // @[Modules.scala 68:83:@13951.4]
  wire [11:0] _T_64439; // @[Modules.scala 68:83:@13953.4]
  wire [10:0] _T_64440; // @[Modules.scala 68:83:@13954.4]
  wire [10:0] buffer_5_671; // @[Modules.scala 68:83:@13955.4]
  wire [11:0] _T_64442; // @[Modules.scala 68:83:@13957.4]
  wire [10:0] _T_64443; // @[Modules.scala 68:83:@13958.4]
  wire [10:0] buffer_5_672; // @[Modules.scala 68:83:@13959.4]
  wire [11:0] _T_64445; // @[Modules.scala 68:83:@13961.4]
  wire [10:0] _T_64446; // @[Modules.scala 68:83:@13962.4]
  wire [10:0] buffer_5_673; // @[Modules.scala 68:83:@13963.4]
  wire [11:0] _T_64451; // @[Modules.scala 68:83:@13969.4]
  wire [10:0] _T_64452; // @[Modules.scala 68:83:@13970.4]
  wire [10:0] buffer_5_675; // @[Modules.scala 68:83:@13971.4]
  wire [11:0] _T_64454; // @[Modules.scala 68:83:@13973.4]
  wire [10:0] _T_64455; // @[Modules.scala 68:83:@13974.4]
  wire [10:0] buffer_5_676; // @[Modules.scala 68:83:@13975.4]
  wire [11:0] _T_64460; // @[Modules.scala 68:83:@13981.4]
  wire [10:0] _T_64461; // @[Modules.scala 68:83:@13982.4]
  wire [10:0] buffer_5_678; // @[Modules.scala 68:83:@13983.4]
  wire [11:0] _T_64463; // @[Modules.scala 68:83:@13985.4]
  wire [10:0] _T_64464; // @[Modules.scala 68:83:@13986.4]
  wire [10:0] buffer_5_679; // @[Modules.scala 68:83:@13987.4]
  wire [11:0] _T_64466; // @[Modules.scala 68:83:@13989.4]
  wire [10:0] _T_64467; // @[Modules.scala 68:83:@13990.4]
  wire [10:0] buffer_5_680; // @[Modules.scala 68:83:@13991.4]
  wire [11:0] _T_64469; // @[Modules.scala 68:83:@13993.4]
  wire [10:0] _T_64470; // @[Modules.scala 68:83:@13994.4]
  wire [10:0] buffer_5_681; // @[Modules.scala 68:83:@13995.4]
  wire [11:0] _T_64472; // @[Modules.scala 68:83:@13997.4]
  wire [10:0] _T_64473; // @[Modules.scala 68:83:@13998.4]
  wire [10:0] buffer_5_682; // @[Modules.scala 68:83:@13999.4]
  wire [11:0] _T_64475; // @[Modules.scala 68:83:@14001.4]
  wire [10:0] _T_64476; // @[Modules.scala 68:83:@14002.4]
  wire [10:0] buffer_5_683; // @[Modules.scala 68:83:@14003.4]
  wire [11:0] _T_64481; // @[Modules.scala 68:83:@14009.4]
  wire [10:0] _T_64482; // @[Modules.scala 68:83:@14010.4]
  wire [10:0] buffer_5_685; // @[Modules.scala 68:83:@14011.4]
  wire [11:0] _T_64484; // @[Modules.scala 71:109:@14013.4]
  wire [10:0] _T_64485; // @[Modules.scala 71:109:@14014.4]
  wire [10:0] buffer_5_686; // @[Modules.scala 71:109:@14015.4]
  wire [11:0] _T_64487; // @[Modules.scala 71:109:@14017.4]
  wire [10:0] _T_64488; // @[Modules.scala 71:109:@14018.4]
  wire [10:0] buffer_5_687; // @[Modules.scala 71:109:@14019.4]
  wire [11:0] _T_64490; // @[Modules.scala 71:109:@14021.4]
  wire [10:0] _T_64491; // @[Modules.scala 71:109:@14022.4]
  wire [10:0] buffer_5_688; // @[Modules.scala 71:109:@14023.4]
  wire [11:0] _T_64493; // @[Modules.scala 71:109:@14025.4]
  wire [10:0] _T_64494; // @[Modules.scala 71:109:@14026.4]
  wire [10:0] buffer_5_689; // @[Modules.scala 71:109:@14027.4]
  wire [11:0] _T_64496; // @[Modules.scala 71:109:@14029.4]
  wire [10:0] _T_64497; // @[Modules.scala 71:109:@14030.4]
  wire [10:0] buffer_5_690; // @[Modules.scala 71:109:@14031.4]
  wire [11:0] _T_64499; // @[Modules.scala 71:109:@14033.4]
  wire [10:0] _T_64500; // @[Modules.scala 71:109:@14034.4]
  wire [10:0] buffer_5_691; // @[Modules.scala 71:109:@14035.4]
  wire [11:0] _T_64502; // @[Modules.scala 71:109:@14037.4]
  wire [10:0] _T_64503; // @[Modules.scala 71:109:@14038.4]
  wire [10:0] buffer_5_692; // @[Modules.scala 71:109:@14039.4]
  wire [11:0] _T_64505; // @[Modules.scala 71:109:@14041.4]
  wire [10:0] _T_64506; // @[Modules.scala 71:109:@14042.4]
  wire [10:0] buffer_5_693; // @[Modules.scala 71:109:@14043.4]
  wire [11:0] _T_64508; // @[Modules.scala 71:109:@14045.4]
  wire [10:0] _T_64509; // @[Modules.scala 71:109:@14046.4]
  wire [10:0] buffer_5_694; // @[Modules.scala 71:109:@14047.4]
  wire [11:0] _T_64511; // @[Modules.scala 71:109:@14049.4]
  wire [10:0] _T_64512; // @[Modules.scala 71:109:@14050.4]
  wire [10:0] buffer_5_695; // @[Modules.scala 71:109:@14051.4]
  wire [11:0] _T_64514; // @[Modules.scala 71:109:@14053.4]
  wire [10:0] _T_64515; // @[Modules.scala 71:109:@14054.4]
  wire [10:0] buffer_5_696; // @[Modules.scala 71:109:@14055.4]
  wire [11:0] _T_64517; // @[Modules.scala 71:109:@14057.4]
  wire [10:0] _T_64518; // @[Modules.scala 71:109:@14058.4]
  wire [10:0] buffer_5_697; // @[Modules.scala 71:109:@14059.4]
  wire [11:0] _T_64520; // @[Modules.scala 71:109:@14061.4]
  wire [10:0] _T_64521; // @[Modules.scala 71:109:@14062.4]
  wire [10:0] buffer_5_698; // @[Modules.scala 71:109:@14063.4]
  wire [11:0] _T_64523; // @[Modules.scala 71:109:@14065.4]
  wire [10:0] _T_64524; // @[Modules.scala 71:109:@14066.4]
  wire [10:0] buffer_5_699; // @[Modules.scala 71:109:@14067.4]
  wire [11:0] _T_64526; // @[Modules.scala 71:109:@14069.4]
  wire [10:0] _T_64527; // @[Modules.scala 71:109:@14070.4]
  wire [10:0] buffer_5_700; // @[Modules.scala 71:109:@14071.4]
  wire [11:0] _T_64529; // @[Modules.scala 71:109:@14073.4]
  wire [10:0] _T_64530; // @[Modules.scala 71:109:@14074.4]
  wire [10:0] buffer_5_701; // @[Modules.scala 71:109:@14075.4]
  wire [11:0] _T_64532; // @[Modules.scala 71:109:@14077.4]
  wire [10:0] _T_64533; // @[Modules.scala 71:109:@14078.4]
  wire [10:0] buffer_5_702; // @[Modules.scala 71:109:@14079.4]
  wire [11:0] _T_64535; // @[Modules.scala 71:109:@14081.4]
  wire [10:0] _T_64536; // @[Modules.scala 71:109:@14082.4]
  wire [10:0] buffer_5_703; // @[Modules.scala 71:109:@14083.4]
  wire [11:0] _T_64538; // @[Modules.scala 71:109:@14085.4]
  wire [10:0] _T_64539; // @[Modules.scala 71:109:@14086.4]
  wire [10:0] buffer_5_704; // @[Modules.scala 71:109:@14087.4]
  wire [11:0] _T_64541; // @[Modules.scala 71:109:@14089.4]
  wire [10:0] _T_64542; // @[Modules.scala 71:109:@14090.4]
  wire [10:0] buffer_5_705; // @[Modules.scala 71:109:@14091.4]
  wire [11:0] _T_64544; // @[Modules.scala 71:109:@14093.4]
  wire [10:0] _T_64545; // @[Modules.scala 71:109:@14094.4]
  wire [10:0] buffer_5_706; // @[Modules.scala 71:109:@14095.4]
  wire [11:0] _T_64547; // @[Modules.scala 71:109:@14097.4]
  wire [10:0] _T_64548; // @[Modules.scala 71:109:@14098.4]
  wire [10:0] buffer_5_707; // @[Modules.scala 71:109:@14099.4]
  wire [11:0] _T_64550; // @[Modules.scala 71:109:@14101.4]
  wire [10:0] _T_64551; // @[Modules.scala 71:109:@14102.4]
  wire [10:0] buffer_5_708; // @[Modules.scala 71:109:@14103.4]
  wire [11:0] _T_64553; // @[Modules.scala 71:109:@14105.4]
  wire [10:0] _T_64554; // @[Modules.scala 71:109:@14106.4]
  wire [10:0] buffer_5_709; // @[Modules.scala 71:109:@14107.4]
  wire [11:0] _T_64556; // @[Modules.scala 71:109:@14109.4]
  wire [10:0] _T_64557; // @[Modules.scala 71:109:@14110.4]
  wire [10:0] buffer_5_710; // @[Modules.scala 71:109:@14111.4]
  wire [11:0] _T_64559; // @[Modules.scala 71:109:@14113.4]
  wire [10:0] _T_64560; // @[Modules.scala 71:109:@14114.4]
  wire [10:0] buffer_5_711; // @[Modules.scala 71:109:@14115.4]
  wire [11:0] _T_64562; // @[Modules.scala 71:109:@14117.4]
  wire [10:0] _T_64563; // @[Modules.scala 71:109:@14118.4]
  wire [10:0] buffer_5_712; // @[Modules.scala 71:109:@14119.4]
  wire [11:0] _T_64565; // @[Modules.scala 71:109:@14121.4]
  wire [10:0] _T_64566; // @[Modules.scala 71:109:@14122.4]
  wire [10:0] buffer_5_713; // @[Modules.scala 71:109:@14123.4]
  wire [11:0] _T_64568; // @[Modules.scala 71:109:@14125.4]
  wire [10:0] _T_64569; // @[Modules.scala 71:109:@14126.4]
  wire [10:0] buffer_5_714; // @[Modules.scala 71:109:@14127.4]
  wire [11:0] _T_64571; // @[Modules.scala 71:109:@14129.4]
  wire [10:0] _T_64572; // @[Modules.scala 71:109:@14130.4]
  wire [10:0] buffer_5_715; // @[Modules.scala 71:109:@14131.4]
  wire [11:0] _T_64574; // @[Modules.scala 71:109:@14133.4]
  wire [10:0] _T_64575; // @[Modules.scala 71:109:@14134.4]
  wire [10:0] buffer_5_716; // @[Modules.scala 71:109:@14135.4]
  wire [11:0] _T_64577; // @[Modules.scala 71:109:@14137.4]
  wire [10:0] _T_64578; // @[Modules.scala 71:109:@14138.4]
  wire [10:0] buffer_5_717; // @[Modules.scala 71:109:@14139.4]
  wire [11:0] _T_64580; // @[Modules.scala 71:109:@14141.4]
  wire [10:0] _T_64581; // @[Modules.scala 71:109:@14142.4]
  wire [10:0] buffer_5_718; // @[Modules.scala 71:109:@14143.4]
  wire [11:0] _T_64583; // @[Modules.scala 71:109:@14145.4]
  wire [10:0] _T_64584; // @[Modules.scala 71:109:@14146.4]
  wire [10:0] buffer_5_719; // @[Modules.scala 71:109:@14147.4]
  wire [11:0] _T_64586; // @[Modules.scala 71:109:@14149.4]
  wire [10:0] _T_64587; // @[Modules.scala 71:109:@14150.4]
  wire [10:0] buffer_5_720; // @[Modules.scala 71:109:@14151.4]
  wire [11:0] _T_64589; // @[Modules.scala 71:109:@14153.4]
  wire [10:0] _T_64590; // @[Modules.scala 71:109:@14154.4]
  wire [10:0] buffer_5_721; // @[Modules.scala 71:109:@14155.4]
  wire [11:0] _T_64592; // @[Modules.scala 71:109:@14157.4]
  wire [10:0] _T_64593; // @[Modules.scala 71:109:@14158.4]
  wire [10:0] buffer_5_722; // @[Modules.scala 71:109:@14159.4]
  wire [11:0] _T_64595; // @[Modules.scala 71:109:@14161.4]
  wire [10:0] _T_64596; // @[Modules.scala 71:109:@14162.4]
  wire [10:0] buffer_5_723; // @[Modules.scala 71:109:@14163.4]
  wire [11:0] _T_64598; // @[Modules.scala 71:109:@14165.4]
  wire [10:0] _T_64599; // @[Modules.scala 71:109:@14166.4]
  wire [10:0] buffer_5_724; // @[Modules.scala 71:109:@14167.4]
  wire [11:0] _T_64601; // @[Modules.scala 71:109:@14169.4]
  wire [10:0] _T_64602; // @[Modules.scala 71:109:@14170.4]
  wire [10:0] buffer_5_725; // @[Modules.scala 71:109:@14171.4]
  wire [11:0] _T_64604; // @[Modules.scala 71:109:@14173.4]
  wire [10:0] _T_64605; // @[Modules.scala 71:109:@14174.4]
  wire [10:0] buffer_5_726; // @[Modules.scala 71:109:@14175.4]
  wire [11:0] _T_64607; // @[Modules.scala 71:109:@14177.4]
  wire [10:0] _T_64608; // @[Modules.scala 71:109:@14178.4]
  wire [10:0] buffer_5_727; // @[Modules.scala 71:109:@14179.4]
  wire [11:0] _T_64610; // @[Modules.scala 71:109:@14181.4]
  wire [10:0] _T_64611; // @[Modules.scala 71:109:@14182.4]
  wire [10:0] buffer_5_728; // @[Modules.scala 71:109:@14183.4]
  wire [11:0] _T_64613; // @[Modules.scala 71:109:@14185.4]
  wire [10:0] _T_64614; // @[Modules.scala 71:109:@14186.4]
  wire [10:0] buffer_5_729; // @[Modules.scala 71:109:@14187.4]
  wire [11:0] _T_64616; // @[Modules.scala 71:109:@14189.4]
  wire [10:0] _T_64617; // @[Modules.scala 71:109:@14190.4]
  wire [10:0] buffer_5_730; // @[Modules.scala 71:109:@14191.4]
  wire [11:0] _T_64619; // @[Modules.scala 71:109:@14193.4]
  wire [10:0] _T_64620; // @[Modules.scala 71:109:@14194.4]
  wire [10:0] buffer_5_731; // @[Modules.scala 71:109:@14195.4]
  wire [11:0] _T_64622; // @[Modules.scala 71:109:@14197.4]
  wire [10:0] _T_64623; // @[Modules.scala 71:109:@14198.4]
  wire [10:0] buffer_5_732; // @[Modules.scala 71:109:@14199.4]
  wire [11:0] _T_64625; // @[Modules.scala 71:109:@14201.4]
  wire [10:0] _T_64626; // @[Modules.scala 71:109:@14202.4]
  wire [10:0] buffer_5_733; // @[Modules.scala 71:109:@14203.4]
  wire [11:0] _T_64628; // @[Modules.scala 71:109:@14205.4]
  wire [10:0] _T_64629; // @[Modules.scala 71:109:@14206.4]
  wire [10:0] buffer_5_734; // @[Modules.scala 71:109:@14207.4]
  wire [11:0] _T_64631; // @[Modules.scala 78:156:@14210.4]
  wire [10:0] _T_64632; // @[Modules.scala 78:156:@14211.4]
  wire [10:0] buffer_5_736; // @[Modules.scala 78:156:@14212.4]
  wire [11:0] _T_64634; // @[Modules.scala 78:156:@14214.4]
  wire [10:0] _T_64635; // @[Modules.scala 78:156:@14215.4]
  wire [10:0] buffer_5_737; // @[Modules.scala 78:156:@14216.4]
  wire [11:0] _T_64637; // @[Modules.scala 78:156:@14218.4]
  wire [10:0] _T_64638; // @[Modules.scala 78:156:@14219.4]
  wire [10:0] buffer_5_738; // @[Modules.scala 78:156:@14220.4]
  wire [11:0] _T_64640; // @[Modules.scala 78:156:@14222.4]
  wire [10:0] _T_64641; // @[Modules.scala 78:156:@14223.4]
  wire [10:0] buffer_5_739; // @[Modules.scala 78:156:@14224.4]
  wire [11:0] _T_64643; // @[Modules.scala 78:156:@14226.4]
  wire [10:0] _T_64644; // @[Modules.scala 78:156:@14227.4]
  wire [10:0] buffer_5_740; // @[Modules.scala 78:156:@14228.4]
  wire [11:0] _T_64646; // @[Modules.scala 78:156:@14230.4]
  wire [10:0] _T_64647; // @[Modules.scala 78:156:@14231.4]
  wire [10:0] buffer_5_741; // @[Modules.scala 78:156:@14232.4]
  wire [11:0] _T_64649; // @[Modules.scala 78:156:@14234.4]
  wire [10:0] _T_64650; // @[Modules.scala 78:156:@14235.4]
  wire [10:0] buffer_5_742; // @[Modules.scala 78:156:@14236.4]
  wire [11:0] _T_64652; // @[Modules.scala 78:156:@14238.4]
  wire [10:0] _T_64653; // @[Modules.scala 78:156:@14239.4]
  wire [10:0] buffer_5_743; // @[Modules.scala 78:156:@14240.4]
  wire [11:0] _T_64655; // @[Modules.scala 78:156:@14242.4]
  wire [10:0] _T_64656; // @[Modules.scala 78:156:@14243.4]
  wire [10:0] buffer_5_744; // @[Modules.scala 78:156:@14244.4]
  wire [11:0] _T_64658; // @[Modules.scala 78:156:@14246.4]
  wire [10:0] _T_64659; // @[Modules.scala 78:156:@14247.4]
  wire [10:0] buffer_5_745; // @[Modules.scala 78:156:@14248.4]
  wire [11:0] _T_64661; // @[Modules.scala 78:156:@14250.4]
  wire [10:0] _T_64662; // @[Modules.scala 78:156:@14251.4]
  wire [10:0] buffer_5_746; // @[Modules.scala 78:156:@14252.4]
  wire [11:0] _T_64664; // @[Modules.scala 78:156:@14254.4]
  wire [10:0] _T_64665; // @[Modules.scala 78:156:@14255.4]
  wire [10:0] buffer_5_747; // @[Modules.scala 78:156:@14256.4]
  wire [11:0] _T_64667; // @[Modules.scala 78:156:@14258.4]
  wire [10:0] _T_64668; // @[Modules.scala 78:156:@14259.4]
  wire [10:0] buffer_5_748; // @[Modules.scala 78:156:@14260.4]
  wire [11:0] _T_64670; // @[Modules.scala 78:156:@14262.4]
  wire [10:0] _T_64671; // @[Modules.scala 78:156:@14263.4]
  wire [10:0] buffer_5_749; // @[Modules.scala 78:156:@14264.4]
  wire [11:0] _T_64673; // @[Modules.scala 78:156:@14266.4]
  wire [10:0] _T_64674; // @[Modules.scala 78:156:@14267.4]
  wire [10:0] buffer_5_750; // @[Modules.scala 78:156:@14268.4]
  wire [11:0] _T_64676; // @[Modules.scala 78:156:@14270.4]
  wire [10:0] _T_64677; // @[Modules.scala 78:156:@14271.4]
  wire [10:0] buffer_5_751; // @[Modules.scala 78:156:@14272.4]
  wire [11:0] _T_64679; // @[Modules.scala 78:156:@14274.4]
  wire [10:0] _T_64680; // @[Modules.scala 78:156:@14275.4]
  wire [10:0] buffer_5_752; // @[Modules.scala 78:156:@14276.4]
  wire [11:0] _T_64682; // @[Modules.scala 78:156:@14278.4]
  wire [10:0] _T_64683; // @[Modules.scala 78:156:@14279.4]
  wire [10:0] buffer_5_753; // @[Modules.scala 78:156:@14280.4]
  wire [11:0] _T_64685; // @[Modules.scala 78:156:@14282.4]
  wire [10:0] _T_64686; // @[Modules.scala 78:156:@14283.4]
  wire [10:0] buffer_5_754; // @[Modules.scala 78:156:@14284.4]
  wire [11:0] _T_64688; // @[Modules.scala 78:156:@14286.4]
  wire [10:0] _T_64689; // @[Modules.scala 78:156:@14287.4]
  wire [10:0] buffer_5_755; // @[Modules.scala 78:156:@14288.4]
  wire [11:0] _T_64691; // @[Modules.scala 78:156:@14290.4]
  wire [10:0] _T_64692; // @[Modules.scala 78:156:@14291.4]
  wire [10:0] buffer_5_756; // @[Modules.scala 78:156:@14292.4]
  wire [11:0] _T_64694; // @[Modules.scala 78:156:@14294.4]
  wire [10:0] _T_64695; // @[Modules.scala 78:156:@14295.4]
  wire [10:0] buffer_5_757; // @[Modules.scala 78:156:@14296.4]
  wire [11:0] _T_64697; // @[Modules.scala 78:156:@14298.4]
  wire [10:0] _T_64698; // @[Modules.scala 78:156:@14299.4]
  wire [10:0] buffer_5_758; // @[Modules.scala 78:156:@14300.4]
  wire [11:0] _T_64700; // @[Modules.scala 78:156:@14302.4]
  wire [10:0] _T_64701; // @[Modules.scala 78:156:@14303.4]
  wire [10:0] buffer_5_759; // @[Modules.scala 78:156:@14304.4]
  wire [11:0] _T_64703; // @[Modules.scala 78:156:@14306.4]
  wire [10:0] _T_64704; // @[Modules.scala 78:156:@14307.4]
  wire [10:0] buffer_5_760; // @[Modules.scala 78:156:@14308.4]
  wire [11:0] _T_64706; // @[Modules.scala 78:156:@14310.4]
  wire [10:0] _T_64707; // @[Modules.scala 78:156:@14311.4]
  wire [10:0] buffer_5_761; // @[Modules.scala 78:156:@14312.4]
  wire [11:0] _T_64709; // @[Modules.scala 78:156:@14314.4]
  wire [10:0] _T_64710; // @[Modules.scala 78:156:@14315.4]
  wire [10:0] buffer_5_762; // @[Modules.scala 78:156:@14316.4]
  wire [11:0] _T_64712; // @[Modules.scala 78:156:@14318.4]
  wire [10:0] _T_64713; // @[Modules.scala 78:156:@14319.4]
  wire [10:0] buffer_5_763; // @[Modules.scala 78:156:@14320.4]
  wire [11:0] _T_64715; // @[Modules.scala 78:156:@14322.4]
  wire [10:0] _T_64716; // @[Modules.scala 78:156:@14323.4]
  wire [10:0] buffer_5_764; // @[Modules.scala 78:156:@14324.4]
  wire [11:0] _T_64718; // @[Modules.scala 78:156:@14326.4]
  wire [10:0] _T_64719; // @[Modules.scala 78:156:@14327.4]
  wire [10:0] buffer_5_765; // @[Modules.scala 78:156:@14328.4]
  wire [11:0] _T_64721; // @[Modules.scala 78:156:@14330.4]
  wire [10:0] _T_64722; // @[Modules.scala 78:156:@14331.4]
  wire [10:0] buffer_5_766; // @[Modules.scala 78:156:@14332.4]
  wire [11:0] _T_64724; // @[Modules.scala 78:156:@14334.4]
  wire [10:0] _T_64725; // @[Modules.scala 78:156:@14335.4]
  wire [10:0] buffer_5_767; // @[Modules.scala 78:156:@14336.4]
  wire [11:0] _T_64727; // @[Modules.scala 78:156:@14338.4]
  wire [10:0] _T_64728; // @[Modules.scala 78:156:@14339.4]
  wire [10:0] buffer_5_768; // @[Modules.scala 78:156:@14340.4]
  wire [11:0] _T_64730; // @[Modules.scala 78:156:@14342.4]
  wire [10:0] _T_64731; // @[Modules.scala 78:156:@14343.4]
  wire [10:0] buffer_5_769; // @[Modules.scala 78:156:@14344.4]
  wire [11:0] _T_64733; // @[Modules.scala 78:156:@14346.4]
  wire [10:0] _T_64734; // @[Modules.scala 78:156:@14347.4]
  wire [10:0] buffer_5_770; // @[Modules.scala 78:156:@14348.4]
  wire [11:0] _T_64736; // @[Modules.scala 78:156:@14350.4]
  wire [10:0] _T_64737; // @[Modules.scala 78:156:@14351.4]
  wire [10:0] buffer_5_771; // @[Modules.scala 78:156:@14352.4]
  wire [11:0] _T_64739; // @[Modules.scala 78:156:@14354.4]
  wire [10:0] _T_64740; // @[Modules.scala 78:156:@14355.4]
  wire [10:0] buffer_5_772; // @[Modules.scala 78:156:@14356.4]
  wire [11:0] _T_64742; // @[Modules.scala 78:156:@14358.4]
  wire [10:0] _T_64743; // @[Modules.scala 78:156:@14359.4]
  wire [10:0] buffer_5_773; // @[Modules.scala 78:156:@14360.4]
  wire [11:0] _T_64745; // @[Modules.scala 78:156:@14362.4]
  wire [10:0] _T_64746; // @[Modules.scala 78:156:@14363.4]
  wire [10:0] buffer_5_774; // @[Modules.scala 78:156:@14364.4]
  wire [11:0] _T_64748; // @[Modules.scala 78:156:@14366.4]
  wire [10:0] _T_64749; // @[Modules.scala 78:156:@14367.4]
  wire [10:0] buffer_5_775; // @[Modules.scala 78:156:@14368.4]
  wire [11:0] _T_64751; // @[Modules.scala 78:156:@14370.4]
  wire [10:0] _T_64752; // @[Modules.scala 78:156:@14371.4]
  wire [10:0] buffer_5_776; // @[Modules.scala 78:156:@14372.4]
  wire [11:0] _T_64754; // @[Modules.scala 78:156:@14374.4]
  wire [10:0] _T_64755; // @[Modules.scala 78:156:@14375.4]
  wire [10:0] buffer_5_777; // @[Modules.scala 78:156:@14376.4]
  wire [11:0] _T_64757; // @[Modules.scala 78:156:@14378.4]
  wire [10:0] _T_64758; // @[Modules.scala 78:156:@14379.4]
  wire [10:0] buffer_5_778; // @[Modules.scala 78:156:@14380.4]
  wire [11:0] _T_64760; // @[Modules.scala 78:156:@14382.4]
  wire [10:0] _T_64761; // @[Modules.scala 78:156:@14383.4]
  wire [10:0] buffer_5_779; // @[Modules.scala 78:156:@14384.4]
  wire [11:0] _T_64763; // @[Modules.scala 78:156:@14386.4]
  wire [10:0] _T_64764; // @[Modules.scala 78:156:@14387.4]
  wire [10:0] buffer_5_780; // @[Modules.scala 78:156:@14388.4]
  wire [11:0] _T_64766; // @[Modules.scala 78:156:@14390.4]
  wire [10:0] _T_64767; // @[Modules.scala 78:156:@14391.4]
  wire [10:0] buffer_5_781; // @[Modules.scala 78:156:@14392.4]
  wire [11:0] _T_64769; // @[Modules.scala 78:156:@14394.4]
  wire [10:0] _T_64770; // @[Modules.scala 78:156:@14395.4]
  wire [10:0] buffer_5_782; // @[Modules.scala 78:156:@14396.4]
  wire [11:0] _T_64772; // @[Modules.scala 78:156:@14398.4]
  wire [10:0] _T_64773; // @[Modules.scala 78:156:@14399.4]
  wire [10:0] buffer_5_783; // @[Modules.scala 78:156:@14400.4]
  wire [5:0] _T_64873; // @[Modules.scala 37:46:@14544.4]
  wire [4:0] _T_64874; // @[Modules.scala 37:46:@14545.4]
  wire [4:0] _T_64875; // @[Modules.scala 37:46:@14546.4]
  wire [5:0] _T_64909; // @[Modules.scala 37:46:@14603.4]
  wire [4:0] _T_64910; // @[Modules.scala 37:46:@14604.4]
  wire [4:0] _T_64911; // @[Modules.scala 37:46:@14605.4]
  wire [5:0] _T_64948; // @[Modules.scala 37:46:@14664.4]
  wire [4:0] _T_64949; // @[Modules.scala 37:46:@14665.4]
  wire [4:0] _T_64950; // @[Modules.scala 37:46:@14666.4]
  wire [5:0] _T_64960; // @[Modules.scala 37:46:@14680.4]
  wire [4:0] _T_64961; // @[Modules.scala 37:46:@14681.4]
  wire [4:0] _T_64962; // @[Modules.scala 37:46:@14682.4]
  wire [5:0] _T_64963; // @[Modules.scala 37:46:@14684.4]
  wire [4:0] _T_64964; // @[Modules.scala 37:46:@14685.4]
  wire [4:0] _T_64965; // @[Modules.scala 37:46:@14686.4]
  wire [5:0] _T_65020; // @[Modules.scala 37:46:@14784.4]
  wire [4:0] _T_65021; // @[Modules.scala 37:46:@14785.4]
  wire [4:0] _T_65022; // @[Modules.scala 37:46:@14786.4]
  wire [5:0] _T_65058; // @[Modules.scala 37:46:@14844.4]
  wire [4:0] _T_65059; // @[Modules.scala 37:46:@14845.4]
  wire [4:0] _T_65060; // @[Modules.scala 37:46:@14846.4]
  wire [5:0] _T_65102; // @[Modules.scala 37:46:@14892.4]
  wire [4:0] _T_65103; // @[Modules.scala 37:46:@14893.4]
  wire [4:0] _T_65104; // @[Modules.scala 37:46:@14894.4]
  wire [11:0] _T_65226; // @[Modules.scala 65:57:@15066.4]
  wire [10:0] _T_65227; // @[Modules.scala 65:57:@15067.4]
  wire [10:0] buffer_6_393; // @[Modules.scala 65:57:@15068.4]
  wire [11:0] _T_65229; // @[Modules.scala 65:57:@15070.4]
  wire [10:0] _T_65230; // @[Modules.scala 65:57:@15071.4]
  wire [10:0] buffer_6_394; // @[Modules.scala 65:57:@15072.4]
  wire [11:0] _T_65262; // @[Modules.scala 65:57:@15114.4]
  wire [10:0] _T_65263; // @[Modules.scala 65:57:@15115.4]
  wire [10:0] buffer_6_405; // @[Modules.scala 65:57:@15116.4]
  wire [11:0] _T_65265; // @[Modules.scala 65:57:@15118.4]
  wire [10:0] _T_65266; // @[Modules.scala 65:57:@15119.4]
  wire [10:0] buffer_6_406; // @[Modules.scala 65:57:@15120.4]
  wire [11:0] _T_65286; // @[Modules.scala 65:57:@15146.4]
  wire [10:0] _T_65287; // @[Modules.scala 65:57:@15147.4]
  wire [10:0] buffer_6_413; // @[Modules.scala 65:57:@15148.4]
  wire [10:0] buffer_6_53; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65301; // @[Modules.scala 65:57:@15166.4]
  wire [10:0] _T_65302; // @[Modules.scala 65:57:@15167.4]
  wire [10:0] buffer_6_418; // @[Modules.scala 65:57:@15168.4]
  wire [11:0] _T_65304; // @[Modules.scala 65:57:@15170.4]
  wire [10:0] _T_65305; // @[Modules.scala 65:57:@15171.4]
  wire [10:0] buffer_6_419; // @[Modules.scala 65:57:@15172.4]
  wire [10:0] buffer_6_73; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65331; // @[Modules.scala 65:57:@15206.4]
  wire [10:0] _T_65332; // @[Modules.scala 65:57:@15207.4]
  wire [10:0] buffer_6_428; // @[Modules.scala 65:57:@15208.4]
  wire [10:0] buffer_6_74; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65334; // @[Modules.scala 65:57:@15210.4]
  wire [10:0] _T_65335; // @[Modules.scala 65:57:@15211.4]
  wire [10:0] buffer_6_429; // @[Modules.scala 65:57:@15212.4]
  wire [11:0] _T_65346; // @[Modules.scala 65:57:@15226.4]
  wire [10:0] _T_65347; // @[Modules.scala 65:57:@15227.4]
  wire [10:0] buffer_6_433; // @[Modules.scala 65:57:@15228.4]
  wire [10:0] buffer_6_86; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65352; // @[Modules.scala 65:57:@15234.4]
  wire [10:0] _T_65353; // @[Modules.scala 65:57:@15235.4]
  wire [10:0] buffer_6_435; // @[Modules.scala 65:57:@15236.4]
  wire [11:0] _T_65355; // @[Modules.scala 65:57:@15238.4]
  wire [10:0] _T_65356; // @[Modules.scala 65:57:@15239.4]
  wire [10:0] buffer_6_436; // @[Modules.scala 65:57:@15240.4]
  wire [10:0] buffer_6_94; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65364; // @[Modules.scala 65:57:@15250.4]
  wire [10:0] _T_65365; // @[Modules.scala 65:57:@15251.4]
  wire [10:0] buffer_6_439; // @[Modules.scala 65:57:@15252.4]
  wire [10:0] buffer_6_97; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65367; // @[Modules.scala 65:57:@15254.4]
  wire [10:0] _T_65368; // @[Modules.scala 65:57:@15255.4]
  wire [10:0] buffer_6_440; // @[Modules.scala 65:57:@15256.4]
  wire [11:0] _T_65370; // @[Modules.scala 65:57:@15258.4]
  wire [10:0] _T_65371; // @[Modules.scala 65:57:@15259.4]
  wire [10:0] buffer_6_441; // @[Modules.scala 65:57:@15260.4]
  wire [11:0] _T_65373; // @[Modules.scala 65:57:@15262.4]
  wire [10:0] _T_65374; // @[Modules.scala 65:57:@15263.4]
  wire [10:0] buffer_6_442; // @[Modules.scala 65:57:@15264.4]
  wire [10:0] buffer_6_102; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65376; // @[Modules.scala 65:57:@15266.4]
  wire [10:0] _T_65377; // @[Modules.scala 65:57:@15267.4]
  wire [10:0] buffer_6_443; // @[Modules.scala 65:57:@15268.4]
  wire [11:0] _T_65379; // @[Modules.scala 65:57:@15270.4]
  wire [10:0] _T_65380; // @[Modules.scala 65:57:@15271.4]
  wire [10:0] buffer_6_444; // @[Modules.scala 65:57:@15272.4]
  wire [10:0] buffer_6_107; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65382; // @[Modules.scala 65:57:@15274.4]
  wire [10:0] _T_65383; // @[Modules.scala 65:57:@15275.4]
  wire [10:0] buffer_6_445; // @[Modules.scala 65:57:@15276.4]
  wire [11:0] _T_65385; // @[Modules.scala 65:57:@15278.4]
  wire [10:0] _T_65386; // @[Modules.scala 65:57:@15279.4]
  wire [10:0] buffer_6_446; // @[Modules.scala 65:57:@15280.4]
  wire [11:0] _T_65391; // @[Modules.scala 65:57:@15286.4]
  wire [10:0] _T_65392; // @[Modules.scala 65:57:@15287.4]
  wire [10:0] buffer_6_448; // @[Modules.scala 65:57:@15288.4]
  wire [11:0] _T_65397; // @[Modules.scala 65:57:@15294.4]
  wire [10:0] _T_65398; // @[Modules.scala 65:57:@15295.4]
  wire [10:0] buffer_6_450; // @[Modules.scala 65:57:@15296.4]
  wire [10:0] buffer_6_120; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_121; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65403; // @[Modules.scala 65:57:@15302.4]
  wire [10:0] _T_65404; // @[Modules.scala 65:57:@15303.4]
  wire [10:0] buffer_6_452; // @[Modules.scala 65:57:@15304.4]
  wire [10:0] buffer_6_123; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65406; // @[Modules.scala 65:57:@15306.4]
  wire [10:0] _T_65407; // @[Modules.scala 65:57:@15307.4]
  wire [10:0] buffer_6_453; // @[Modules.scala 65:57:@15308.4]
  wire [11:0] _T_65412; // @[Modules.scala 65:57:@15314.4]
  wire [10:0] _T_65413; // @[Modules.scala 65:57:@15315.4]
  wire [10:0] buffer_6_455; // @[Modules.scala 65:57:@15316.4]
  wire [10:0] buffer_6_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65415; // @[Modules.scala 65:57:@15318.4]
  wire [10:0] _T_65416; // @[Modules.scala 65:57:@15319.4]
  wire [10:0] buffer_6_456; // @[Modules.scala 65:57:@15320.4]
  wire [10:0] buffer_6_131; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65418; // @[Modules.scala 65:57:@15322.4]
  wire [10:0] _T_65419; // @[Modules.scala 65:57:@15323.4]
  wire [10:0] buffer_6_457; // @[Modules.scala 65:57:@15324.4]
  wire [11:0] _T_65427; // @[Modules.scala 65:57:@15334.4]
  wire [10:0] _T_65428; // @[Modules.scala 65:57:@15335.4]
  wire [10:0] buffer_6_460; // @[Modules.scala 65:57:@15336.4]
  wire [11:0] _T_65433; // @[Modules.scala 65:57:@15342.4]
  wire [10:0] _T_65434; // @[Modules.scala 65:57:@15343.4]
  wire [10:0] buffer_6_462; // @[Modules.scala 65:57:@15344.4]
  wire [10:0] buffer_6_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65439; // @[Modules.scala 65:57:@15350.4]
  wire [10:0] _T_65440; // @[Modules.scala 65:57:@15351.4]
  wire [10:0] buffer_6_464; // @[Modules.scala 65:57:@15352.4]
  wire [11:0] _T_65442; // @[Modules.scala 65:57:@15354.4]
  wire [10:0] _T_65443; // @[Modules.scala 65:57:@15355.4]
  wire [10:0] buffer_6_465; // @[Modules.scala 65:57:@15356.4]
  wire [11:0] _T_65445; // @[Modules.scala 65:57:@15358.4]
  wire [10:0] _T_65446; // @[Modules.scala 65:57:@15359.4]
  wire [10:0] buffer_6_466; // @[Modules.scala 65:57:@15360.4]
  wire [10:0] buffer_6_150; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65448; // @[Modules.scala 65:57:@15362.4]
  wire [10:0] _T_65449; // @[Modules.scala 65:57:@15363.4]
  wire [10:0] buffer_6_467; // @[Modules.scala 65:57:@15364.4]
  wire [11:0] _T_65454; // @[Modules.scala 65:57:@15370.4]
  wire [10:0] _T_65455; // @[Modules.scala 65:57:@15371.4]
  wire [10:0] buffer_6_469; // @[Modules.scala 65:57:@15372.4]
  wire [10:0] buffer_6_156; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65457; // @[Modules.scala 65:57:@15374.4]
  wire [10:0] _T_65458; // @[Modules.scala 65:57:@15375.4]
  wire [10:0] buffer_6_470; // @[Modules.scala 65:57:@15376.4]
  wire [10:0] buffer_6_158; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65460; // @[Modules.scala 65:57:@15378.4]
  wire [10:0] _T_65461; // @[Modules.scala 65:57:@15379.4]
  wire [10:0] buffer_6_471; // @[Modules.scala 65:57:@15380.4]
  wire [10:0] buffer_6_161; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65463; // @[Modules.scala 65:57:@15382.4]
  wire [10:0] _T_65464; // @[Modules.scala 65:57:@15383.4]
  wire [10:0] buffer_6_472; // @[Modules.scala 65:57:@15384.4]
  wire [10:0] buffer_6_162; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65466; // @[Modules.scala 65:57:@15386.4]
  wire [10:0] _T_65467; // @[Modules.scala 65:57:@15387.4]
  wire [10:0] buffer_6_473; // @[Modules.scala 65:57:@15388.4]
  wire [10:0] buffer_6_169; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65475; // @[Modules.scala 65:57:@15398.4]
  wire [10:0] _T_65476; // @[Modules.scala 65:57:@15399.4]
  wire [10:0] buffer_6_476; // @[Modules.scala 65:57:@15400.4]
  wire [10:0] buffer_6_170; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65478; // @[Modules.scala 65:57:@15402.4]
  wire [10:0] _T_65479; // @[Modules.scala 65:57:@15403.4]
  wire [10:0] buffer_6_477; // @[Modules.scala 65:57:@15404.4]
  wire [10:0] buffer_6_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65481; // @[Modules.scala 65:57:@15406.4]
  wire [10:0] _T_65482; // @[Modules.scala 65:57:@15407.4]
  wire [10:0] buffer_6_478; // @[Modules.scala 65:57:@15408.4]
  wire [10:0] buffer_6_175; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65484; // @[Modules.scala 65:57:@15410.4]
  wire [10:0] _T_65485; // @[Modules.scala 65:57:@15411.4]
  wire [10:0] buffer_6_479; // @[Modules.scala 65:57:@15412.4]
  wire [10:0] buffer_6_178; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_179; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65490; // @[Modules.scala 65:57:@15418.4]
  wire [10:0] _T_65491; // @[Modules.scala 65:57:@15419.4]
  wire [10:0] buffer_6_481; // @[Modules.scala 65:57:@15420.4]
  wire [11:0] _T_65496; // @[Modules.scala 65:57:@15426.4]
  wire [10:0] _T_65497; // @[Modules.scala 65:57:@15427.4]
  wire [10:0] buffer_6_483; // @[Modules.scala 65:57:@15428.4]
  wire [11:0] _T_65502; // @[Modules.scala 65:57:@15434.4]
  wire [10:0] _T_65503; // @[Modules.scala 65:57:@15435.4]
  wire [10:0] buffer_6_485; // @[Modules.scala 65:57:@15436.4]
  wire [10:0] buffer_6_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65505; // @[Modules.scala 65:57:@15438.4]
  wire [10:0] _T_65506; // @[Modules.scala 65:57:@15439.4]
  wire [10:0] buffer_6_486; // @[Modules.scala 65:57:@15440.4]
  wire [10:0] buffer_6_196; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65517; // @[Modules.scala 65:57:@15454.4]
  wire [10:0] _T_65518; // @[Modules.scala 65:57:@15455.4]
  wire [10:0] buffer_6_490; // @[Modules.scala 65:57:@15456.4]
  wire [11:0] _T_65523; // @[Modules.scala 65:57:@15462.4]
  wire [10:0] _T_65524; // @[Modules.scala 65:57:@15463.4]
  wire [10:0] buffer_6_492; // @[Modules.scala 65:57:@15464.4]
  wire [11:0] _T_65526; // @[Modules.scala 65:57:@15466.4]
  wire [10:0] _T_65527; // @[Modules.scala 65:57:@15467.4]
  wire [10:0] buffer_6_493; // @[Modules.scala 65:57:@15468.4]
  wire [10:0] buffer_6_207; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65532; // @[Modules.scala 65:57:@15474.4]
  wire [10:0] _T_65533; // @[Modules.scala 65:57:@15475.4]
  wire [10:0] buffer_6_495; // @[Modules.scala 65:57:@15476.4]
  wire [11:0] _T_65535; // @[Modules.scala 65:57:@15478.4]
  wire [10:0] _T_65536; // @[Modules.scala 65:57:@15479.4]
  wire [10:0] buffer_6_496; // @[Modules.scala 65:57:@15480.4]
  wire [11:0] _T_65538; // @[Modules.scala 65:57:@15482.4]
  wire [10:0] _T_65539; // @[Modules.scala 65:57:@15483.4]
  wire [10:0] buffer_6_497; // @[Modules.scala 65:57:@15484.4]
  wire [10:0] buffer_6_213; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65541; // @[Modules.scala 65:57:@15486.4]
  wire [10:0] _T_65542; // @[Modules.scala 65:57:@15487.4]
  wire [10:0] buffer_6_498; // @[Modules.scala 65:57:@15488.4]
  wire [10:0] buffer_6_214; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65544; // @[Modules.scala 65:57:@15490.4]
  wire [10:0] _T_65545; // @[Modules.scala 65:57:@15491.4]
  wire [10:0] buffer_6_499; // @[Modules.scala 65:57:@15492.4]
  wire [10:0] buffer_6_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65547; // @[Modules.scala 65:57:@15494.4]
  wire [10:0] _T_65548; // @[Modules.scala 65:57:@15495.4]
  wire [10:0] buffer_6_500; // @[Modules.scala 65:57:@15496.4]
  wire [10:0] buffer_6_219; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65550; // @[Modules.scala 65:57:@15498.4]
  wire [10:0] _T_65551; // @[Modules.scala 65:57:@15499.4]
  wire [10:0] buffer_6_501; // @[Modules.scala 65:57:@15500.4]
  wire [10:0] buffer_6_221; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65553; // @[Modules.scala 65:57:@15502.4]
  wire [10:0] _T_65554; // @[Modules.scala 65:57:@15503.4]
  wire [10:0] buffer_6_502; // @[Modules.scala 65:57:@15504.4]
  wire [11:0] _T_65559; // @[Modules.scala 65:57:@15510.4]
  wire [10:0] _T_65560; // @[Modules.scala 65:57:@15511.4]
  wire [10:0] buffer_6_504; // @[Modules.scala 65:57:@15512.4]
  wire [10:0] buffer_6_229; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65565; // @[Modules.scala 65:57:@15518.4]
  wire [10:0] _T_65566; // @[Modules.scala 65:57:@15519.4]
  wire [10:0] buffer_6_506; // @[Modules.scala 65:57:@15520.4]
  wire [11:0] _T_65568; // @[Modules.scala 65:57:@15522.4]
  wire [10:0] _T_65569; // @[Modules.scala 65:57:@15523.4]
  wire [10:0] buffer_6_507; // @[Modules.scala 65:57:@15524.4]
  wire [10:0] buffer_6_233; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65571; // @[Modules.scala 65:57:@15526.4]
  wire [10:0] _T_65572; // @[Modules.scala 65:57:@15527.4]
  wire [10:0] buffer_6_508; // @[Modules.scala 65:57:@15528.4]
  wire [10:0] buffer_6_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65574; // @[Modules.scala 65:57:@15530.4]
  wire [10:0] _T_65575; // @[Modules.scala 65:57:@15531.4]
  wire [10:0] buffer_6_509; // @[Modules.scala 65:57:@15532.4]
  wire [11:0] _T_65580; // @[Modules.scala 65:57:@15538.4]
  wire [10:0] _T_65581; // @[Modules.scala 65:57:@15539.4]
  wire [10:0] buffer_6_511; // @[Modules.scala 65:57:@15540.4]
  wire [10:0] buffer_6_241; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65583; // @[Modules.scala 65:57:@15542.4]
  wire [10:0] _T_65584; // @[Modules.scala 65:57:@15543.4]
  wire [10:0] buffer_6_512; // @[Modules.scala 65:57:@15544.4]
  wire [11:0] _T_65586; // @[Modules.scala 65:57:@15546.4]
  wire [10:0] _T_65587; // @[Modules.scala 65:57:@15547.4]
  wire [10:0] buffer_6_513; // @[Modules.scala 65:57:@15548.4]
  wire [11:0] _T_65592; // @[Modules.scala 65:57:@15554.4]
  wire [10:0] _T_65593; // @[Modules.scala 65:57:@15555.4]
  wire [10:0] buffer_6_515; // @[Modules.scala 65:57:@15556.4]
  wire [10:0] buffer_6_252; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_6_253; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65601; // @[Modules.scala 65:57:@15566.4]
  wire [10:0] _T_65602; // @[Modules.scala 65:57:@15567.4]
  wire [10:0] buffer_6_518; // @[Modules.scala 65:57:@15568.4]
  wire [11:0] _T_65610; // @[Modules.scala 65:57:@15578.4]
  wire [10:0] _T_65611; // @[Modules.scala 65:57:@15579.4]
  wire [10:0] buffer_6_521; // @[Modules.scala 65:57:@15580.4]
  wire [10:0] buffer_6_294; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65664; // @[Modules.scala 65:57:@15650.4]
  wire [10:0] _T_65665; // @[Modules.scala 65:57:@15651.4]
  wire [10:0] buffer_6_539; // @[Modules.scala 65:57:@15652.4]
  wire [10:0] buffer_6_306; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65682; // @[Modules.scala 65:57:@15674.4]
  wire [10:0] _T_65683; // @[Modules.scala 65:57:@15675.4]
  wire [10:0] buffer_6_545; // @[Modules.scala 65:57:@15676.4]
  wire [10:0] buffer_6_312; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65691; // @[Modules.scala 65:57:@15686.4]
  wire [10:0] _T_65692; // @[Modules.scala 65:57:@15687.4]
  wire [10:0] buffer_6_548; // @[Modules.scala 65:57:@15688.4]
  wire [10:0] buffer_6_315; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65694; // @[Modules.scala 65:57:@15690.4]
  wire [10:0] _T_65695; // @[Modules.scala 65:57:@15691.4]
  wire [10:0] buffer_6_549; // @[Modules.scala 65:57:@15692.4]
  wire [11:0] _T_65709; // @[Modules.scala 65:57:@15710.4]
  wire [10:0] _T_65710; // @[Modules.scala 65:57:@15711.4]
  wire [10:0] buffer_6_554; // @[Modules.scala 65:57:@15712.4]
  wire [10:0] buffer_6_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65712; // @[Modules.scala 65:57:@15714.4]
  wire [10:0] _T_65713; // @[Modules.scala 65:57:@15715.4]
  wire [10:0] buffer_6_555; // @[Modules.scala 65:57:@15716.4]
  wire [11:0] _T_65724; // @[Modules.scala 65:57:@15730.4]
  wire [10:0] _T_65725; // @[Modules.scala 65:57:@15731.4]
  wire [10:0] buffer_6_559; // @[Modules.scala 65:57:@15732.4]
  wire [11:0] _T_65727; // @[Modules.scala 65:57:@15734.4]
  wire [10:0] _T_65728; // @[Modules.scala 65:57:@15735.4]
  wire [10:0] buffer_6_560; // @[Modules.scala 65:57:@15736.4]
  wire [11:0] _T_65739; // @[Modules.scala 65:57:@15750.4]
  wire [10:0] _T_65740; // @[Modules.scala 65:57:@15751.4]
  wire [10:0] buffer_6_564; // @[Modules.scala 65:57:@15752.4]
  wire [11:0] _T_65742; // @[Modules.scala 65:57:@15754.4]
  wire [10:0] _T_65743; // @[Modules.scala 65:57:@15755.4]
  wire [10:0] buffer_6_565; // @[Modules.scala 65:57:@15756.4]
  wire [11:0] _T_65754; // @[Modules.scala 65:57:@15770.4]
  wire [10:0] _T_65755; // @[Modules.scala 65:57:@15771.4]
  wire [10:0] buffer_6_569; // @[Modules.scala 65:57:@15772.4]
  wire [10:0] buffer_6_357; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65757; // @[Modules.scala 65:57:@15774.4]
  wire [10:0] _T_65758; // @[Modules.scala 65:57:@15775.4]
  wire [10:0] buffer_6_570; // @[Modules.scala 65:57:@15776.4]
  wire [10:0] buffer_6_359; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65760; // @[Modules.scala 65:57:@15778.4]
  wire [10:0] _T_65761; // @[Modules.scala 65:57:@15779.4]
  wire [10:0] buffer_6_571; // @[Modules.scala 65:57:@15780.4]
  wire [11:0] _T_65769; // @[Modules.scala 65:57:@15790.4]
  wire [10:0] _T_65770; // @[Modules.scala 65:57:@15791.4]
  wire [10:0] buffer_6_574; // @[Modules.scala 65:57:@15792.4]
  wire [11:0] _T_65784; // @[Modules.scala 65:57:@15810.4]
  wire [10:0] _T_65785; // @[Modules.scala 65:57:@15811.4]
  wire [10:0] buffer_6_579; // @[Modules.scala 65:57:@15812.4]
  wire [10:0] buffer_6_384; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65799; // @[Modules.scala 65:57:@15830.4]
  wire [10:0] _T_65800; // @[Modules.scala 65:57:@15831.4]
  wire [10:0] buffer_6_584; // @[Modules.scala 65:57:@15832.4]
  wire [10:0] buffer_6_388; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_65805; // @[Modules.scala 65:57:@15838.4]
  wire [10:0] _T_65806; // @[Modules.scala 65:57:@15839.4]
  wire [10:0] buffer_6_586; // @[Modules.scala 65:57:@15840.4]
  wire [11:0] _T_65811; // @[Modules.scala 68:83:@15846.4]
  wire [10:0] _T_65812; // @[Modules.scala 68:83:@15847.4]
  wire [10:0] buffer_6_588; // @[Modules.scala 68:83:@15848.4]
  wire [11:0] _T_65814; // @[Modules.scala 68:83:@15850.4]
  wire [10:0] _T_65815; // @[Modules.scala 68:83:@15851.4]
  wire [10:0] buffer_6_589; // @[Modules.scala 68:83:@15852.4]
  wire [11:0] _T_65817; // @[Modules.scala 68:83:@15854.4]
  wire [10:0] _T_65818; // @[Modules.scala 68:83:@15855.4]
  wire [10:0] buffer_6_590; // @[Modules.scala 68:83:@15856.4]
  wire [11:0] _T_65820; // @[Modules.scala 68:83:@15858.4]
  wire [10:0] _T_65821; // @[Modules.scala 68:83:@15859.4]
  wire [10:0] buffer_6_591; // @[Modules.scala 68:83:@15860.4]
  wire [11:0] _T_65823; // @[Modules.scala 68:83:@15862.4]
  wire [10:0] _T_65824; // @[Modules.scala 68:83:@15863.4]
  wire [10:0] buffer_6_592; // @[Modules.scala 68:83:@15864.4]
  wire [11:0] _T_65829; // @[Modules.scala 68:83:@15870.4]
  wire [10:0] _T_65830; // @[Modules.scala 68:83:@15871.4]
  wire [10:0] buffer_6_594; // @[Modules.scala 68:83:@15872.4]
  wire [11:0] _T_65832; // @[Modules.scala 68:83:@15874.4]
  wire [10:0] _T_65833; // @[Modules.scala 68:83:@15875.4]
  wire [10:0] buffer_6_595; // @[Modules.scala 68:83:@15876.4]
  wire [11:0] _T_65841; // @[Modules.scala 68:83:@15886.4]
  wire [10:0] _T_65842; // @[Modules.scala 68:83:@15887.4]
  wire [10:0] buffer_6_598; // @[Modules.scala 68:83:@15888.4]
  wire [11:0] _T_65850; // @[Modules.scala 68:83:@15898.4]
  wire [10:0] _T_65851; // @[Modules.scala 68:83:@15899.4]
  wire [10:0] buffer_6_601; // @[Modules.scala 68:83:@15900.4]
  wire [11:0] _T_65853; // @[Modules.scala 68:83:@15902.4]
  wire [10:0] _T_65854; // @[Modules.scala 68:83:@15903.4]
  wire [10:0] buffer_6_602; // @[Modules.scala 68:83:@15904.4]
  wire [11:0] _T_65859; // @[Modules.scala 68:83:@15910.4]
  wire [10:0] _T_65860; // @[Modules.scala 68:83:@15911.4]
  wire [10:0] buffer_6_604; // @[Modules.scala 68:83:@15912.4]
  wire [11:0] _T_65862; // @[Modules.scala 68:83:@15914.4]
  wire [10:0] _T_65863; // @[Modules.scala 68:83:@15915.4]
  wire [10:0] buffer_6_605; // @[Modules.scala 68:83:@15916.4]
  wire [11:0] _T_65865; // @[Modules.scala 68:83:@15918.4]
  wire [10:0] _T_65866; // @[Modules.scala 68:83:@15919.4]
  wire [10:0] buffer_6_606; // @[Modules.scala 68:83:@15920.4]
  wire [11:0] _T_65871; // @[Modules.scala 68:83:@15926.4]
  wire [10:0] _T_65872; // @[Modules.scala 68:83:@15927.4]
  wire [10:0] buffer_6_608; // @[Modules.scala 68:83:@15928.4]
  wire [11:0] _T_65874; // @[Modules.scala 68:83:@15930.4]
  wire [10:0] _T_65875; // @[Modules.scala 68:83:@15931.4]
  wire [10:0] buffer_6_609; // @[Modules.scala 68:83:@15932.4]
  wire [11:0] _T_65877; // @[Modules.scala 68:83:@15934.4]
  wire [10:0] _T_65878; // @[Modules.scala 68:83:@15935.4]
  wire [10:0] buffer_6_610; // @[Modules.scala 68:83:@15936.4]
  wire [11:0] _T_65880; // @[Modules.scala 68:83:@15938.4]
  wire [10:0] _T_65881; // @[Modules.scala 68:83:@15939.4]
  wire [10:0] buffer_6_611; // @[Modules.scala 68:83:@15940.4]
  wire [11:0] _T_65883; // @[Modules.scala 68:83:@15942.4]
  wire [10:0] _T_65884; // @[Modules.scala 68:83:@15943.4]
  wire [10:0] buffer_6_612; // @[Modules.scala 68:83:@15944.4]
  wire [11:0] _T_65886; // @[Modules.scala 68:83:@15946.4]
  wire [10:0] _T_65887; // @[Modules.scala 68:83:@15947.4]
  wire [10:0] buffer_6_613; // @[Modules.scala 68:83:@15948.4]
  wire [11:0] _T_65889; // @[Modules.scala 68:83:@15950.4]
  wire [10:0] _T_65890; // @[Modules.scala 68:83:@15951.4]
  wire [10:0] buffer_6_614; // @[Modules.scala 68:83:@15952.4]
  wire [11:0] _T_65892; // @[Modules.scala 68:83:@15954.4]
  wire [10:0] _T_65893; // @[Modules.scala 68:83:@15955.4]
  wire [10:0] buffer_6_615; // @[Modules.scala 68:83:@15956.4]
  wire [11:0] _T_65895; // @[Modules.scala 68:83:@15958.4]
  wire [10:0] _T_65896; // @[Modules.scala 68:83:@15959.4]
  wire [10:0] buffer_6_616; // @[Modules.scala 68:83:@15960.4]
  wire [11:0] _T_65898; // @[Modules.scala 68:83:@15962.4]
  wire [10:0] _T_65899; // @[Modules.scala 68:83:@15963.4]
  wire [10:0] buffer_6_617; // @[Modules.scala 68:83:@15964.4]
  wire [11:0] _T_65901; // @[Modules.scala 68:83:@15966.4]
  wire [10:0] _T_65902; // @[Modules.scala 68:83:@15967.4]
  wire [10:0] buffer_6_618; // @[Modules.scala 68:83:@15968.4]
  wire [11:0] _T_65904; // @[Modules.scala 68:83:@15970.4]
  wire [10:0] _T_65905; // @[Modules.scala 68:83:@15971.4]
  wire [10:0] buffer_6_619; // @[Modules.scala 68:83:@15972.4]
  wire [11:0] _T_65907; // @[Modules.scala 68:83:@15974.4]
  wire [10:0] _T_65908; // @[Modules.scala 68:83:@15975.4]
  wire [10:0] buffer_6_620; // @[Modules.scala 68:83:@15976.4]
  wire [11:0] _T_65913; // @[Modules.scala 68:83:@15982.4]
  wire [10:0] _T_65914; // @[Modules.scala 68:83:@15983.4]
  wire [10:0] buffer_6_622; // @[Modules.scala 68:83:@15984.4]
  wire [11:0] _T_65916; // @[Modules.scala 68:83:@15986.4]
  wire [10:0] _T_65917; // @[Modules.scala 68:83:@15987.4]
  wire [10:0] buffer_6_623; // @[Modules.scala 68:83:@15988.4]
  wire [11:0] _T_65919; // @[Modules.scala 68:83:@15990.4]
  wire [10:0] _T_65920; // @[Modules.scala 68:83:@15991.4]
  wire [10:0] buffer_6_624; // @[Modules.scala 68:83:@15992.4]
  wire [11:0] _T_65922; // @[Modules.scala 68:83:@15994.4]
  wire [10:0] _T_65923; // @[Modules.scala 68:83:@15995.4]
  wire [10:0] buffer_6_625; // @[Modules.scala 68:83:@15996.4]
  wire [11:0] _T_65925; // @[Modules.scala 68:83:@15998.4]
  wire [10:0] _T_65926; // @[Modules.scala 68:83:@15999.4]
  wire [10:0] buffer_6_626; // @[Modules.scala 68:83:@16000.4]
  wire [11:0] _T_65928; // @[Modules.scala 68:83:@16002.4]
  wire [10:0] _T_65929; // @[Modules.scala 68:83:@16003.4]
  wire [10:0] buffer_6_627; // @[Modules.scala 68:83:@16004.4]
  wire [11:0] _T_65931; // @[Modules.scala 68:83:@16006.4]
  wire [10:0] _T_65932; // @[Modules.scala 68:83:@16007.4]
  wire [10:0] buffer_6_628; // @[Modules.scala 68:83:@16008.4]
  wire [11:0] _T_65934; // @[Modules.scala 68:83:@16010.4]
  wire [10:0] _T_65935; // @[Modules.scala 68:83:@16011.4]
  wire [10:0] buffer_6_629; // @[Modules.scala 68:83:@16012.4]
  wire [11:0] _T_65937; // @[Modules.scala 68:83:@16014.4]
  wire [10:0] _T_65938; // @[Modules.scala 68:83:@16015.4]
  wire [10:0] buffer_6_630; // @[Modules.scala 68:83:@16016.4]
  wire [11:0] _T_65940; // @[Modules.scala 68:83:@16018.4]
  wire [10:0] _T_65941; // @[Modules.scala 68:83:@16019.4]
  wire [10:0] buffer_6_631; // @[Modules.scala 68:83:@16020.4]
  wire [11:0] _T_65943; // @[Modules.scala 68:83:@16022.4]
  wire [10:0] _T_65944; // @[Modules.scala 68:83:@16023.4]
  wire [10:0] buffer_6_632; // @[Modules.scala 68:83:@16024.4]
  wire [11:0] _T_65946; // @[Modules.scala 68:83:@16026.4]
  wire [10:0] _T_65947; // @[Modules.scala 68:83:@16027.4]
  wire [10:0] buffer_6_633; // @[Modules.scala 68:83:@16028.4]
  wire [11:0] _T_65949; // @[Modules.scala 68:83:@16030.4]
  wire [10:0] _T_65950; // @[Modules.scala 68:83:@16031.4]
  wire [10:0] buffer_6_634; // @[Modules.scala 68:83:@16032.4]
  wire [11:0] _T_65952; // @[Modules.scala 68:83:@16034.4]
  wire [10:0] _T_65953; // @[Modules.scala 68:83:@16035.4]
  wire [10:0] buffer_6_635; // @[Modules.scala 68:83:@16036.4]
  wire [11:0] _T_65955; // @[Modules.scala 68:83:@16038.4]
  wire [10:0] _T_65956; // @[Modules.scala 68:83:@16039.4]
  wire [10:0] buffer_6_636; // @[Modules.scala 68:83:@16040.4]
  wire [11:0] _T_65958; // @[Modules.scala 68:83:@16042.4]
  wire [10:0] _T_65959; // @[Modules.scala 68:83:@16043.4]
  wire [10:0] buffer_6_637; // @[Modules.scala 68:83:@16044.4]
  wire [11:0] _T_65961; // @[Modules.scala 68:83:@16046.4]
  wire [10:0] _T_65962; // @[Modules.scala 68:83:@16047.4]
  wire [10:0] buffer_6_638; // @[Modules.scala 68:83:@16048.4]
  wire [11:0] _T_65964; // @[Modules.scala 68:83:@16050.4]
  wire [10:0] _T_65965; // @[Modules.scala 68:83:@16051.4]
  wire [10:0] buffer_6_639; // @[Modules.scala 68:83:@16052.4]
  wire [11:0] _T_65967; // @[Modules.scala 68:83:@16054.4]
  wire [10:0] _T_65968; // @[Modules.scala 68:83:@16055.4]
  wire [10:0] buffer_6_640; // @[Modules.scala 68:83:@16056.4]
  wire [11:0] _T_65970; // @[Modules.scala 68:83:@16058.4]
  wire [10:0] _T_65971; // @[Modules.scala 68:83:@16059.4]
  wire [10:0] buffer_6_641; // @[Modules.scala 68:83:@16060.4]
  wire [11:0] _T_65973; // @[Modules.scala 68:83:@16062.4]
  wire [10:0] _T_65974; // @[Modules.scala 68:83:@16063.4]
  wire [10:0] buffer_6_642; // @[Modules.scala 68:83:@16064.4]
  wire [11:0] _T_65976; // @[Modules.scala 68:83:@16066.4]
  wire [10:0] _T_65977; // @[Modules.scala 68:83:@16067.4]
  wire [10:0] buffer_6_643; // @[Modules.scala 68:83:@16068.4]
  wire [11:0] _T_65979; // @[Modules.scala 68:83:@16070.4]
  wire [10:0] _T_65980; // @[Modules.scala 68:83:@16071.4]
  wire [10:0] buffer_6_644; // @[Modules.scala 68:83:@16072.4]
  wire [11:0] _T_65982; // @[Modules.scala 68:83:@16074.4]
  wire [10:0] _T_65983; // @[Modules.scala 68:83:@16075.4]
  wire [10:0] buffer_6_645; // @[Modules.scala 68:83:@16076.4]
  wire [11:0] _T_65985; // @[Modules.scala 68:83:@16078.4]
  wire [10:0] _T_65986; // @[Modules.scala 68:83:@16079.4]
  wire [10:0] buffer_6_646; // @[Modules.scala 68:83:@16080.4]
  wire [11:0] _T_65988; // @[Modules.scala 68:83:@16082.4]
  wire [10:0] _T_65989; // @[Modules.scala 68:83:@16083.4]
  wire [10:0] buffer_6_647; // @[Modules.scala 68:83:@16084.4]
  wire [11:0] _T_65991; // @[Modules.scala 68:83:@16086.4]
  wire [10:0] _T_65992; // @[Modules.scala 68:83:@16087.4]
  wire [10:0] buffer_6_648; // @[Modules.scala 68:83:@16088.4]
  wire [11:0] _T_65994; // @[Modules.scala 68:83:@16090.4]
  wire [10:0] _T_65995; // @[Modules.scala 68:83:@16091.4]
  wire [10:0] buffer_6_649; // @[Modules.scala 68:83:@16092.4]
  wire [11:0] _T_66000; // @[Modules.scala 68:83:@16098.4]
  wire [10:0] _T_66001; // @[Modules.scala 68:83:@16099.4]
  wire [10:0] buffer_6_651; // @[Modules.scala 68:83:@16100.4]
  wire [11:0] _T_66003; // @[Modules.scala 68:83:@16102.4]
  wire [10:0] _T_66004; // @[Modules.scala 68:83:@16103.4]
  wire [10:0] buffer_6_652; // @[Modules.scala 68:83:@16104.4]
  wire [11:0] _T_66018; // @[Modules.scala 68:83:@16122.4]
  wire [10:0] _T_66019; // @[Modules.scala 68:83:@16123.4]
  wire [10:0] buffer_6_657; // @[Modules.scala 68:83:@16124.4]
  wire [11:0] _T_66030; // @[Modules.scala 68:83:@16138.4]
  wire [10:0] _T_66031; // @[Modules.scala 68:83:@16139.4]
  wire [10:0] buffer_6_661; // @[Modules.scala 68:83:@16140.4]
  wire [11:0] _T_66039; // @[Modules.scala 68:83:@16150.4]
  wire [10:0] _T_66040; // @[Modules.scala 68:83:@16151.4]
  wire [10:0] buffer_6_664; // @[Modules.scala 68:83:@16152.4]
  wire [11:0] _T_66045; // @[Modules.scala 68:83:@16158.4]
  wire [10:0] _T_66046; // @[Modules.scala 68:83:@16159.4]
  wire [10:0] buffer_6_666; // @[Modules.scala 68:83:@16160.4]
  wire [11:0] _T_66051; // @[Modules.scala 68:83:@16166.4]
  wire [10:0] _T_66052; // @[Modules.scala 68:83:@16167.4]
  wire [10:0] buffer_6_668; // @[Modules.scala 68:83:@16168.4]
  wire [11:0] _T_66054; // @[Modules.scala 68:83:@16170.4]
  wire [10:0] _T_66055; // @[Modules.scala 68:83:@16171.4]
  wire [10:0] buffer_6_669; // @[Modules.scala 68:83:@16172.4]
  wire [11:0] _T_66060; // @[Modules.scala 68:83:@16178.4]
  wire [10:0] _T_66061; // @[Modules.scala 68:83:@16179.4]
  wire [10:0] buffer_6_671; // @[Modules.scala 68:83:@16180.4]
  wire [11:0] _T_66063; // @[Modules.scala 68:83:@16182.4]
  wire [10:0] _T_66064; // @[Modules.scala 68:83:@16183.4]
  wire [10:0] buffer_6_672; // @[Modules.scala 68:83:@16184.4]
  wire [11:0] _T_66069; // @[Modules.scala 68:83:@16190.4]
  wire [10:0] _T_66070; // @[Modules.scala 68:83:@16191.4]
  wire [10:0] buffer_6_674; // @[Modules.scala 68:83:@16192.4]
  wire [11:0] _T_66072; // @[Modules.scala 68:83:@16194.4]
  wire [10:0] _T_66073; // @[Modules.scala 68:83:@16195.4]
  wire [10:0] buffer_6_675; // @[Modules.scala 68:83:@16196.4]
  wire [11:0] _T_66075; // @[Modules.scala 68:83:@16198.4]
  wire [10:0] _T_66076; // @[Modules.scala 68:83:@16199.4]
  wire [10:0] buffer_6_676; // @[Modules.scala 68:83:@16200.4]
  wire [11:0] _T_66078; // @[Modules.scala 68:83:@16202.4]
  wire [10:0] _T_66079; // @[Modules.scala 68:83:@16203.4]
  wire [10:0] buffer_6_677; // @[Modules.scala 68:83:@16204.4]
  wire [11:0] _T_66081; // @[Modules.scala 68:83:@16206.4]
  wire [10:0] _T_66082; // @[Modules.scala 68:83:@16207.4]
  wire [10:0] buffer_6_678; // @[Modules.scala 68:83:@16208.4]
  wire [11:0] _T_66084; // @[Modules.scala 68:83:@16210.4]
  wire [10:0] _T_66085; // @[Modules.scala 68:83:@16211.4]
  wire [10:0] buffer_6_679; // @[Modules.scala 68:83:@16212.4]
  wire [11:0] _T_66090; // @[Modules.scala 68:83:@16218.4]
  wire [10:0] _T_66091; // @[Modules.scala 68:83:@16219.4]
  wire [10:0] buffer_6_681; // @[Modules.scala 68:83:@16220.4]
  wire [11:0] _T_66093; // @[Modules.scala 68:83:@16222.4]
  wire [10:0] _T_66094; // @[Modules.scala 68:83:@16223.4]
  wire [10:0] buffer_6_682; // @[Modules.scala 68:83:@16224.4]
  wire [11:0] _T_66099; // @[Modules.scala 68:83:@16230.4]
  wire [10:0] _T_66100; // @[Modules.scala 68:83:@16231.4]
  wire [10:0] buffer_6_684; // @[Modules.scala 68:83:@16232.4]
  wire [11:0] _T_66102; // @[Modules.scala 68:83:@16234.4]
  wire [10:0] _T_66103; // @[Modules.scala 68:83:@16235.4]
  wire [10:0] buffer_6_685; // @[Modules.scala 68:83:@16236.4]
  wire [11:0] _T_66105; // @[Modules.scala 71:109:@16238.4]
  wire [10:0] _T_66106; // @[Modules.scala 71:109:@16239.4]
  wire [10:0] buffer_6_686; // @[Modules.scala 71:109:@16240.4]
  wire [11:0] _T_66108; // @[Modules.scala 71:109:@16242.4]
  wire [10:0] _T_66109; // @[Modules.scala 71:109:@16243.4]
  wire [10:0] buffer_6_687; // @[Modules.scala 71:109:@16244.4]
  wire [11:0] _T_66111; // @[Modules.scala 71:109:@16246.4]
  wire [10:0] _T_66112; // @[Modules.scala 71:109:@16247.4]
  wire [10:0] buffer_6_688; // @[Modules.scala 71:109:@16248.4]
  wire [11:0] _T_66114; // @[Modules.scala 71:109:@16250.4]
  wire [10:0] _T_66115; // @[Modules.scala 71:109:@16251.4]
  wire [10:0] buffer_6_689; // @[Modules.scala 71:109:@16252.4]
  wire [11:0] _T_66120; // @[Modules.scala 71:109:@16258.4]
  wire [10:0] _T_66121; // @[Modules.scala 71:109:@16259.4]
  wire [10:0] buffer_6_691; // @[Modules.scala 71:109:@16260.4]
  wire [11:0] _T_66123; // @[Modules.scala 71:109:@16262.4]
  wire [10:0] _T_66124; // @[Modules.scala 71:109:@16263.4]
  wire [10:0] buffer_6_692; // @[Modules.scala 71:109:@16264.4]
  wire [11:0] _T_66126; // @[Modules.scala 71:109:@16266.4]
  wire [10:0] _T_66127; // @[Modules.scala 71:109:@16267.4]
  wire [10:0] buffer_6_693; // @[Modules.scala 71:109:@16268.4]
  wire [11:0] _T_66129; // @[Modules.scala 71:109:@16270.4]
  wire [10:0] _T_66130; // @[Modules.scala 71:109:@16271.4]
  wire [10:0] buffer_6_694; // @[Modules.scala 71:109:@16272.4]
  wire [11:0] _T_66132; // @[Modules.scala 71:109:@16274.4]
  wire [10:0] _T_66133; // @[Modules.scala 71:109:@16275.4]
  wire [10:0] buffer_6_695; // @[Modules.scala 71:109:@16276.4]
  wire [11:0] _T_66135; // @[Modules.scala 71:109:@16278.4]
  wire [10:0] _T_66136; // @[Modules.scala 71:109:@16279.4]
  wire [10:0] buffer_6_696; // @[Modules.scala 71:109:@16280.4]
  wire [11:0] _T_66138; // @[Modules.scala 71:109:@16282.4]
  wire [10:0] _T_66139; // @[Modules.scala 71:109:@16283.4]
  wire [10:0] buffer_6_697; // @[Modules.scala 71:109:@16284.4]
  wire [11:0] _T_66141; // @[Modules.scala 71:109:@16286.4]
  wire [10:0] _T_66142; // @[Modules.scala 71:109:@16287.4]
  wire [10:0] buffer_6_698; // @[Modules.scala 71:109:@16288.4]
  wire [11:0] _T_66144; // @[Modules.scala 71:109:@16290.4]
  wire [10:0] _T_66145; // @[Modules.scala 71:109:@16291.4]
  wire [10:0] buffer_6_699; // @[Modules.scala 71:109:@16292.4]
  wire [11:0] _T_66147; // @[Modules.scala 71:109:@16294.4]
  wire [10:0] _T_66148; // @[Modules.scala 71:109:@16295.4]
  wire [10:0] buffer_6_700; // @[Modules.scala 71:109:@16296.4]
  wire [11:0] _T_66150; // @[Modules.scala 71:109:@16298.4]
  wire [10:0] _T_66151; // @[Modules.scala 71:109:@16299.4]
  wire [10:0] buffer_6_701; // @[Modules.scala 71:109:@16300.4]
  wire [11:0] _T_66153; // @[Modules.scala 71:109:@16302.4]
  wire [10:0] _T_66154; // @[Modules.scala 71:109:@16303.4]
  wire [10:0] buffer_6_702; // @[Modules.scala 71:109:@16304.4]
  wire [11:0] _T_66156; // @[Modules.scala 71:109:@16306.4]
  wire [10:0] _T_66157; // @[Modules.scala 71:109:@16307.4]
  wire [10:0] buffer_6_703; // @[Modules.scala 71:109:@16308.4]
  wire [11:0] _T_66159; // @[Modules.scala 71:109:@16310.4]
  wire [10:0] _T_66160; // @[Modules.scala 71:109:@16311.4]
  wire [10:0] buffer_6_704; // @[Modules.scala 71:109:@16312.4]
  wire [11:0] _T_66162; // @[Modules.scala 71:109:@16314.4]
  wire [10:0] _T_66163; // @[Modules.scala 71:109:@16315.4]
  wire [10:0] buffer_6_705; // @[Modules.scala 71:109:@16316.4]
  wire [11:0] _T_66165; // @[Modules.scala 71:109:@16318.4]
  wire [10:0] _T_66166; // @[Modules.scala 71:109:@16319.4]
  wire [10:0] buffer_6_706; // @[Modules.scala 71:109:@16320.4]
  wire [11:0] _T_66168; // @[Modules.scala 71:109:@16322.4]
  wire [10:0] _T_66169; // @[Modules.scala 71:109:@16323.4]
  wire [10:0] buffer_6_707; // @[Modules.scala 71:109:@16324.4]
  wire [11:0] _T_66171; // @[Modules.scala 71:109:@16326.4]
  wire [10:0] _T_66172; // @[Modules.scala 71:109:@16327.4]
  wire [10:0] buffer_6_708; // @[Modules.scala 71:109:@16328.4]
  wire [11:0] _T_66174; // @[Modules.scala 71:109:@16330.4]
  wire [10:0] _T_66175; // @[Modules.scala 71:109:@16331.4]
  wire [10:0] buffer_6_709; // @[Modules.scala 71:109:@16332.4]
  wire [11:0] _T_66177; // @[Modules.scala 71:109:@16334.4]
  wire [10:0] _T_66178; // @[Modules.scala 71:109:@16335.4]
  wire [10:0] buffer_6_710; // @[Modules.scala 71:109:@16336.4]
  wire [11:0] _T_66180; // @[Modules.scala 71:109:@16338.4]
  wire [10:0] _T_66181; // @[Modules.scala 71:109:@16339.4]
  wire [10:0] buffer_6_711; // @[Modules.scala 71:109:@16340.4]
  wire [11:0] _T_66183; // @[Modules.scala 71:109:@16342.4]
  wire [10:0] _T_66184; // @[Modules.scala 71:109:@16343.4]
  wire [10:0] buffer_6_712; // @[Modules.scala 71:109:@16344.4]
  wire [11:0] _T_66186; // @[Modules.scala 71:109:@16346.4]
  wire [10:0] _T_66187; // @[Modules.scala 71:109:@16347.4]
  wire [10:0] buffer_6_713; // @[Modules.scala 71:109:@16348.4]
  wire [11:0] _T_66189; // @[Modules.scala 71:109:@16350.4]
  wire [10:0] _T_66190; // @[Modules.scala 71:109:@16351.4]
  wire [10:0] buffer_6_714; // @[Modules.scala 71:109:@16352.4]
  wire [11:0] _T_66192; // @[Modules.scala 71:109:@16354.4]
  wire [10:0] _T_66193; // @[Modules.scala 71:109:@16355.4]
  wire [10:0] buffer_6_715; // @[Modules.scala 71:109:@16356.4]
  wire [11:0] _T_66195; // @[Modules.scala 71:109:@16358.4]
  wire [10:0] _T_66196; // @[Modules.scala 71:109:@16359.4]
  wire [10:0] buffer_6_716; // @[Modules.scala 71:109:@16360.4]
  wire [11:0] _T_66198; // @[Modules.scala 71:109:@16362.4]
  wire [10:0] _T_66199; // @[Modules.scala 71:109:@16363.4]
  wire [10:0] buffer_6_717; // @[Modules.scala 71:109:@16364.4]
  wire [11:0] _T_66201; // @[Modules.scala 71:109:@16366.4]
  wire [10:0] _T_66202; // @[Modules.scala 71:109:@16367.4]
  wire [10:0] buffer_6_718; // @[Modules.scala 71:109:@16368.4]
  wire [11:0] _T_66207; // @[Modules.scala 71:109:@16374.4]
  wire [10:0] _T_66208; // @[Modules.scala 71:109:@16375.4]
  wire [10:0] buffer_6_720; // @[Modules.scala 71:109:@16376.4]
  wire [11:0] _T_66213; // @[Modules.scala 71:109:@16382.4]
  wire [10:0] _T_66214; // @[Modules.scala 71:109:@16383.4]
  wire [10:0] buffer_6_722; // @[Modules.scala 71:109:@16384.4]
  wire [11:0] _T_66219; // @[Modules.scala 71:109:@16390.4]
  wire [10:0] _T_66220; // @[Modules.scala 71:109:@16391.4]
  wire [10:0] buffer_6_724; // @[Modules.scala 71:109:@16392.4]
  wire [11:0] _T_66222; // @[Modules.scala 71:109:@16394.4]
  wire [10:0] _T_66223; // @[Modules.scala 71:109:@16395.4]
  wire [10:0] buffer_6_725; // @[Modules.scala 71:109:@16396.4]
  wire [11:0] _T_66225; // @[Modules.scala 71:109:@16398.4]
  wire [10:0] _T_66226; // @[Modules.scala 71:109:@16399.4]
  wire [10:0] buffer_6_726; // @[Modules.scala 71:109:@16400.4]
  wire [11:0] _T_66228; // @[Modules.scala 71:109:@16402.4]
  wire [10:0] _T_66229; // @[Modules.scala 71:109:@16403.4]
  wire [10:0] buffer_6_727; // @[Modules.scala 71:109:@16404.4]
  wire [11:0] _T_66231; // @[Modules.scala 71:109:@16406.4]
  wire [10:0] _T_66232; // @[Modules.scala 71:109:@16407.4]
  wire [10:0] buffer_6_728; // @[Modules.scala 71:109:@16408.4]
  wire [11:0] _T_66234; // @[Modules.scala 71:109:@16410.4]
  wire [10:0] _T_66235; // @[Modules.scala 71:109:@16411.4]
  wire [10:0] buffer_6_729; // @[Modules.scala 71:109:@16412.4]
  wire [11:0] _T_66237; // @[Modules.scala 71:109:@16414.4]
  wire [10:0] _T_66238; // @[Modules.scala 71:109:@16415.4]
  wire [10:0] buffer_6_730; // @[Modules.scala 71:109:@16416.4]
  wire [11:0] _T_66240; // @[Modules.scala 71:109:@16418.4]
  wire [10:0] _T_66241; // @[Modules.scala 71:109:@16419.4]
  wire [10:0] buffer_6_731; // @[Modules.scala 71:109:@16420.4]
  wire [11:0] _T_66243; // @[Modules.scala 71:109:@16422.4]
  wire [10:0] _T_66244; // @[Modules.scala 71:109:@16423.4]
  wire [10:0] buffer_6_732; // @[Modules.scala 71:109:@16424.4]
  wire [11:0] _T_66246; // @[Modules.scala 71:109:@16426.4]
  wire [10:0] _T_66247; // @[Modules.scala 71:109:@16427.4]
  wire [10:0] buffer_6_733; // @[Modules.scala 71:109:@16428.4]
  wire [11:0] _T_66249; // @[Modules.scala 71:109:@16430.4]
  wire [10:0] _T_66250; // @[Modules.scala 71:109:@16431.4]
  wire [10:0] buffer_6_734; // @[Modules.scala 71:109:@16432.4]
  wire [11:0] _T_66252; // @[Modules.scala 78:156:@16435.4]
  wire [10:0] _T_66253; // @[Modules.scala 78:156:@16436.4]
  wire [10:0] buffer_6_736; // @[Modules.scala 78:156:@16437.4]
  wire [11:0] _T_66255; // @[Modules.scala 78:156:@16439.4]
  wire [10:0] _T_66256; // @[Modules.scala 78:156:@16440.4]
  wire [10:0] buffer_6_737; // @[Modules.scala 78:156:@16441.4]
  wire [11:0] _T_66258; // @[Modules.scala 78:156:@16443.4]
  wire [10:0] _T_66259; // @[Modules.scala 78:156:@16444.4]
  wire [10:0] buffer_6_738; // @[Modules.scala 78:156:@16445.4]
  wire [11:0] _T_66261; // @[Modules.scala 78:156:@16447.4]
  wire [10:0] _T_66262; // @[Modules.scala 78:156:@16448.4]
  wire [10:0] buffer_6_739; // @[Modules.scala 78:156:@16449.4]
  wire [11:0] _T_66264; // @[Modules.scala 78:156:@16451.4]
  wire [10:0] _T_66265; // @[Modules.scala 78:156:@16452.4]
  wire [10:0] buffer_6_740; // @[Modules.scala 78:156:@16453.4]
  wire [11:0] _T_66267; // @[Modules.scala 78:156:@16455.4]
  wire [10:0] _T_66268; // @[Modules.scala 78:156:@16456.4]
  wire [10:0] buffer_6_741; // @[Modules.scala 78:156:@16457.4]
  wire [11:0] _T_66270; // @[Modules.scala 78:156:@16459.4]
  wire [10:0] _T_66271; // @[Modules.scala 78:156:@16460.4]
  wire [10:0] buffer_6_742; // @[Modules.scala 78:156:@16461.4]
  wire [11:0] _T_66273; // @[Modules.scala 78:156:@16463.4]
  wire [10:0] _T_66274; // @[Modules.scala 78:156:@16464.4]
  wire [10:0] buffer_6_743; // @[Modules.scala 78:156:@16465.4]
  wire [11:0] _T_66276; // @[Modules.scala 78:156:@16467.4]
  wire [10:0] _T_66277; // @[Modules.scala 78:156:@16468.4]
  wire [10:0] buffer_6_744; // @[Modules.scala 78:156:@16469.4]
  wire [11:0] _T_66279; // @[Modules.scala 78:156:@16471.4]
  wire [10:0] _T_66280; // @[Modules.scala 78:156:@16472.4]
  wire [10:0] buffer_6_745; // @[Modules.scala 78:156:@16473.4]
  wire [11:0] _T_66282; // @[Modules.scala 78:156:@16475.4]
  wire [10:0] _T_66283; // @[Modules.scala 78:156:@16476.4]
  wire [10:0] buffer_6_746; // @[Modules.scala 78:156:@16477.4]
  wire [11:0] _T_66285; // @[Modules.scala 78:156:@16479.4]
  wire [10:0] _T_66286; // @[Modules.scala 78:156:@16480.4]
  wire [10:0] buffer_6_747; // @[Modules.scala 78:156:@16481.4]
  wire [11:0] _T_66288; // @[Modules.scala 78:156:@16483.4]
  wire [10:0] _T_66289; // @[Modules.scala 78:156:@16484.4]
  wire [10:0] buffer_6_748; // @[Modules.scala 78:156:@16485.4]
  wire [11:0] _T_66291; // @[Modules.scala 78:156:@16487.4]
  wire [10:0] _T_66292; // @[Modules.scala 78:156:@16488.4]
  wire [10:0] buffer_6_749; // @[Modules.scala 78:156:@16489.4]
  wire [11:0] _T_66294; // @[Modules.scala 78:156:@16491.4]
  wire [10:0] _T_66295; // @[Modules.scala 78:156:@16492.4]
  wire [10:0] buffer_6_750; // @[Modules.scala 78:156:@16493.4]
  wire [11:0] _T_66297; // @[Modules.scala 78:156:@16495.4]
  wire [10:0] _T_66298; // @[Modules.scala 78:156:@16496.4]
  wire [10:0] buffer_6_751; // @[Modules.scala 78:156:@16497.4]
  wire [11:0] _T_66300; // @[Modules.scala 78:156:@16499.4]
  wire [10:0] _T_66301; // @[Modules.scala 78:156:@16500.4]
  wire [10:0] buffer_6_752; // @[Modules.scala 78:156:@16501.4]
  wire [11:0] _T_66303; // @[Modules.scala 78:156:@16503.4]
  wire [10:0] _T_66304; // @[Modules.scala 78:156:@16504.4]
  wire [10:0] buffer_6_753; // @[Modules.scala 78:156:@16505.4]
  wire [11:0] _T_66306; // @[Modules.scala 78:156:@16507.4]
  wire [10:0] _T_66307; // @[Modules.scala 78:156:@16508.4]
  wire [10:0] buffer_6_754; // @[Modules.scala 78:156:@16509.4]
  wire [11:0] _T_66309; // @[Modules.scala 78:156:@16511.4]
  wire [10:0] _T_66310; // @[Modules.scala 78:156:@16512.4]
  wire [10:0] buffer_6_755; // @[Modules.scala 78:156:@16513.4]
  wire [11:0] _T_66312; // @[Modules.scala 78:156:@16515.4]
  wire [10:0] _T_66313; // @[Modules.scala 78:156:@16516.4]
  wire [10:0] buffer_6_756; // @[Modules.scala 78:156:@16517.4]
  wire [11:0] _T_66315; // @[Modules.scala 78:156:@16519.4]
  wire [10:0] _T_66316; // @[Modules.scala 78:156:@16520.4]
  wire [10:0] buffer_6_757; // @[Modules.scala 78:156:@16521.4]
  wire [11:0] _T_66318; // @[Modules.scala 78:156:@16523.4]
  wire [10:0] _T_66319; // @[Modules.scala 78:156:@16524.4]
  wire [10:0] buffer_6_758; // @[Modules.scala 78:156:@16525.4]
  wire [11:0] _T_66321; // @[Modules.scala 78:156:@16527.4]
  wire [10:0] _T_66322; // @[Modules.scala 78:156:@16528.4]
  wire [10:0] buffer_6_759; // @[Modules.scala 78:156:@16529.4]
  wire [11:0] _T_66324; // @[Modules.scala 78:156:@16531.4]
  wire [10:0] _T_66325; // @[Modules.scala 78:156:@16532.4]
  wire [10:0] buffer_6_760; // @[Modules.scala 78:156:@16533.4]
  wire [11:0] _T_66327; // @[Modules.scala 78:156:@16535.4]
  wire [10:0] _T_66328; // @[Modules.scala 78:156:@16536.4]
  wire [10:0] buffer_6_761; // @[Modules.scala 78:156:@16537.4]
  wire [11:0] _T_66330; // @[Modules.scala 78:156:@16539.4]
  wire [10:0] _T_66331; // @[Modules.scala 78:156:@16540.4]
  wire [10:0] buffer_6_762; // @[Modules.scala 78:156:@16541.4]
  wire [11:0] _T_66333; // @[Modules.scala 78:156:@16543.4]
  wire [10:0] _T_66334; // @[Modules.scala 78:156:@16544.4]
  wire [10:0] buffer_6_763; // @[Modules.scala 78:156:@16545.4]
  wire [11:0] _T_66336; // @[Modules.scala 78:156:@16547.4]
  wire [10:0] _T_66337; // @[Modules.scala 78:156:@16548.4]
  wire [10:0] buffer_6_764; // @[Modules.scala 78:156:@16549.4]
  wire [11:0] _T_66339; // @[Modules.scala 78:156:@16551.4]
  wire [10:0] _T_66340; // @[Modules.scala 78:156:@16552.4]
  wire [10:0] buffer_6_765; // @[Modules.scala 78:156:@16553.4]
  wire [11:0] _T_66342; // @[Modules.scala 78:156:@16555.4]
  wire [10:0] _T_66343; // @[Modules.scala 78:156:@16556.4]
  wire [10:0] buffer_6_766; // @[Modules.scala 78:156:@16557.4]
  wire [11:0] _T_66345; // @[Modules.scala 78:156:@16559.4]
  wire [10:0] _T_66346; // @[Modules.scala 78:156:@16560.4]
  wire [10:0] buffer_6_767; // @[Modules.scala 78:156:@16561.4]
  wire [11:0] _T_66348; // @[Modules.scala 78:156:@16563.4]
  wire [10:0] _T_66349; // @[Modules.scala 78:156:@16564.4]
  wire [10:0] buffer_6_768; // @[Modules.scala 78:156:@16565.4]
  wire [11:0] _T_66351; // @[Modules.scala 78:156:@16567.4]
  wire [10:0] _T_66352; // @[Modules.scala 78:156:@16568.4]
  wire [10:0] buffer_6_769; // @[Modules.scala 78:156:@16569.4]
  wire [11:0] _T_66354; // @[Modules.scala 78:156:@16571.4]
  wire [10:0] _T_66355; // @[Modules.scala 78:156:@16572.4]
  wire [10:0] buffer_6_770; // @[Modules.scala 78:156:@16573.4]
  wire [11:0] _T_66357; // @[Modules.scala 78:156:@16575.4]
  wire [10:0] _T_66358; // @[Modules.scala 78:156:@16576.4]
  wire [10:0] buffer_6_771; // @[Modules.scala 78:156:@16577.4]
  wire [11:0] _T_66360; // @[Modules.scala 78:156:@16579.4]
  wire [10:0] _T_66361; // @[Modules.scala 78:156:@16580.4]
  wire [10:0] buffer_6_772; // @[Modules.scala 78:156:@16581.4]
  wire [11:0] _T_66363; // @[Modules.scala 78:156:@16583.4]
  wire [10:0] _T_66364; // @[Modules.scala 78:156:@16584.4]
  wire [10:0] buffer_6_773; // @[Modules.scala 78:156:@16585.4]
  wire [11:0] _T_66366; // @[Modules.scala 78:156:@16587.4]
  wire [10:0] _T_66367; // @[Modules.scala 78:156:@16588.4]
  wire [10:0] buffer_6_774; // @[Modules.scala 78:156:@16589.4]
  wire [11:0] _T_66369; // @[Modules.scala 78:156:@16591.4]
  wire [10:0] _T_66370; // @[Modules.scala 78:156:@16592.4]
  wire [10:0] buffer_6_775; // @[Modules.scala 78:156:@16593.4]
  wire [11:0] _T_66372; // @[Modules.scala 78:156:@16595.4]
  wire [10:0] _T_66373; // @[Modules.scala 78:156:@16596.4]
  wire [10:0] buffer_6_776; // @[Modules.scala 78:156:@16597.4]
  wire [11:0] _T_66375; // @[Modules.scala 78:156:@16599.4]
  wire [10:0] _T_66376; // @[Modules.scala 78:156:@16600.4]
  wire [10:0] buffer_6_777; // @[Modules.scala 78:156:@16601.4]
  wire [11:0] _T_66378; // @[Modules.scala 78:156:@16603.4]
  wire [10:0] _T_66379; // @[Modules.scala 78:156:@16604.4]
  wire [10:0] buffer_6_778; // @[Modules.scala 78:156:@16605.4]
  wire [11:0] _T_66381; // @[Modules.scala 78:156:@16607.4]
  wire [10:0] _T_66382; // @[Modules.scala 78:156:@16608.4]
  wire [10:0] buffer_6_779; // @[Modules.scala 78:156:@16609.4]
  wire [11:0] _T_66384; // @[Modules.scala 78:156:@16611.4]
  wire [10:0] _T_66385; // @[Modules.scala 78:156:@16612.4]
  wire [10:0] buffer_6_780; // @[Modules.scala 78:156:@16613.4]
  wire [11:0] _T_66387; // @[Modules.scala 78:156:@16615.4]
  wire [10:0] _T_66388; // @[Modules.scala 78:156:@16616.4]
  wire [10:0] buffer_6_781; // @[Modules.scala 78:156:@16617.4]
  wire [11:0] _T_66390; // @[Modules.scala 78:156:@16619.4]
  wire [10:0] _T_66391; // @[Modules.scala 78:156:@16620.4]
  wire [10:0] buffer_6_782; // @[Modules.scala 78:156:@16621.4]
  wire [11:0] _T_66393; // @[Modules.scala 78:156:@16623.4]
  wire [10:0] _T_66394; // @[Modules.scala 78:156:@16624.4]
  wire [10:0] buffer_6_783; // @[Modules.scala 78:156:@16625.4]
  wire [5:0] _T_66396; // @[Modules.scala 37:46:@16628.4]
  wire [4:0] _T_66397; // @[Modules.scala 37:46:@16629.4]
  wire [4:0] _T_66398; // @[Modules.scala 37:46:@16630.4]
  wire [5:0] _T_66427; // @[Modules.scala 37:46:@16679.4]
  wire [4:0] _T_66428; // @[Modules.scala 37:46:@16680.4]
  wire [4:0] _T_66429; // @[Modules.scala 37:46:@16681.4]
  wire [5:0] _T_66557; // @[Modules.scala 37:46:@16871.4]
  wire [4:0] _T_66558; // @[Modules.scala 37:46:@16872.4]
  wire [4:0] _T_66559; // @[Modules.scala 37:46:@16873.4]
  wire [5:0] _T_66599; // @[Modules.scala 37:46:@16932.4]
  wire [4:0] _T_66600; // @[Modules.scala 37:46:@16933.4]
  wire [4:0] _T_66601; // @[Modules.scala 37:46:@16934.4]
  wire [5:0] _T_66602; // @[Modules.scala 37:46:@16936.4]
  wire [4:0] _T_66603; // @[Modules.scala 37:46:@16937.4]
  wire [4:0] _T_66604; // @[Modules.scala 37:46:@16938.4]
  wire [5:0] _T_66618; // @[Modules.scala 37:46:@16958.4]
  wire [4:0] _T_66619; // @[Modules.scala 37:46:@16959.4]
  wire [4:0] _T_66620; // @[Modules.scala 37:46:@16960.4]
  wire [5:0] _T_66648; // @[Modules.scala 37:46:@17002.4]
  wire [4:0] _T_66649; // @[Modules.scala 37:46:@17003.4]
  wire [4:0] _T_66650; // @[Modules.scala 37:46:@17004.4]
  wire [5:0] _T_66927; // @[Modules.scala 37:46:@17405.4]
  wire [4:0] _T_66928; // @[Modules.scala 37:46:@17406.4]
  wire [4:0] _T_66929; // @[Modules.scala 37:46:@17407.4]
  wire [10:0] buffer_7_0; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66930; // @[Modules.scala 65:57:@17410.4]
  wire [10:0] _T_66931; // @[Modules.scala 65:57:@17411.4]
  wire [10:0] buffer_7_392; // @[Modules.scala 65:57:@17412.4]
  wire [11:0] _T_66933; // @[Modules.scala 65:57:@17414.4]
  wire [10:0] _T_66934; // @[Modules.scala 65:57:@17415.4]
  wire [10:0] buffer_7_393; // @[Modules.scala 65:57:@17416.4]
  wire [10:0] buffer_7_8; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66942; // @[Modules.scala 65:57:@17426.4]
  wire [10:0] _T_66943; // @[Modules.scala 65:57:@17427.4]
  wire [10:0] buffer_7_396; // @[Modules.scala 65:57:@17428.4]
  wire [11:0] _T_66945; // @[Modules.scala 65:57:@17430.4]
  wire [10:0] _T_66946; // @[Modules.scala 65:57:@17431.4]
  wire [10:0] buffer_7_397; // @[Modules.scala 65:57:@17432.4]
  wire [11:0] _T_66951; // @[Modules.scala 65:57:@17438.4]
  wire [10:0] _T_66952; // @[Modules.scala 65:57:@17439.4]
  wire [10:0] buffer_7_399; // @[Modules.scala 65:57:@17440.4]
  wire [10:0] buffer_7_17; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66954; // @[Modules.scala 65:57:@17442.4]
  wire [10:0] _T_66955; // @[Modules.scala 65:57:@17443.4]
  wire [10:0] buffer_7_400; // @[Modules.scala 65:57:@17444.4]
  wire [10:0] buffer_7_27; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_66969; // @[Modules.scala 65:57:@17462.4]
  wire [10:0] _T_66970; // @[Modules.scala 65:57:@17463.4]
  wire [10:0] buffer_7_405; // @[Modules.scala 65:57:@17464.4]
  wire [11:0] _T_66975; // @[Modules.scala 65:57:@17470.4]
  wire [10:0] _T_66976; // @[Modules.scala 65:57:@17471.4]
  wire [10:0] buffer_7_407; // @[Modules.scala 65:57:@17472.4]
  wire [11:0] _T_67002; // @[Modules.scala 65:57:@17506.4]
  wire [10:0] _T_67003; // @[Modules.scala 65:57:@17507.4]
  wire [10:0] buffer_7_416; // @[Modules.scala 65:57:@17508.4]
  wire [11:0] _T_67017; // @[Modules.scala 65:57:@17526.4]
  wire [10:0] _T_67018; // @[Modules.scala 65:57:@17527.4]
  wire [10:0] buffer_7_421; // @[Modules.scala 65:57:@17528.4]
  wire [11:0] _T_67020; // @[Modules.scala 65:57:@17530.4]
  wire [10:0] _T_67021; // @[Modules.scala 65:57:@17531.4]
  wire [10:0] buffer_7_422; // @[Modules.scala 65:57:@17532.4]
  wire [10:0] buffer_7_63; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67023; // @[Modules.scala 65:57:@17534.4]
  wire [10:0] _T_67024; // @[Modules.scala 65:57:@17535.4]
  wire [10:0] buffer_7_423; // @[Modules.scala 65:57:@17536.4]
  wire [11:0] _T_67029; // @[Modules.scala 65:57:@17542.4]
  wire [10:0] _T_67030; // @[Modules.scala 65:57:@17543.4]
  wire [10:0] buffer_7_425; // @[Modules.scala 65:57:@17544.4]
  wire [11:0] _T_67038; // @[Modules.scala 65:57:@17554.4]
  wire [10:0] _T_67039; // @[Modules.scala 65:57:@17555.4]
  wire [10:0] buffer_7_428; // @[Modules.scala 65:57:@17556.4]
  wire [11:0] _T_67041; // @[Modules.scala 65:57:@17558.4]
  wire [10:0] _T_67042; // @[Modules.scala 65:57:@17559.4]
  wire [10:0] buffer_7_429; // @[Modules.scala 65:57:@17560.4]
  wire [10:0] buffer_7_76; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67044; // @[Modules.scala 65:57:@17562.4]
  wire [10:0] _T_67045; // @[Modules.scala 65:57:@17563.4]
  wire [10:0] buffer_7_430; // @[Modules.scala 65:57:@17564.4]
  wire [10:0] buffer_7_87; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67059; // @[Modules.scala 65:57:@17582.4]
  wire [10:0] _T_67060; // @[Modules.scala 65:57:@17583.4]
  wire [10:0] buffer_7_435; // @[Modules.scala 65:57:@17584.4]
  wire [10:0] buffer_7_89; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67062; // @[Modules.scala 65:57:@17586.4]
  wire [10:0] _T_67063; // @[Modules.scala 65:57:@17587.4]
  wire [10:0] buffer_7_436; // @[Modules.scala 65:57:@17588.4]
  wire [11:0] _T_67071; // @[Modules.scala 65:57:@17598.4]
  wire [10:0] _T_67072; // @[Modules.scala 65:57:@17599.4]
  wire [10:0] buffer_7_439; // @[Modules.scala 65:57:@17600.4]
  wire [10:0] buffer_7_108; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67092; // @[Modules.scala 65:57:@17626.4]
  wire [10:0] _T_67093; // @[Modules.scala 65:57:@17627.4]
  wire [10:0] buffer_7_446; // @[Modules.scala 65:57:@17628.4]
  wire [11:0] _T_67101; // @[Modules.scala 65:57:@17638.4]
  wire [10:0] _T_67102; // @[Modules.scala 65:57:@17639.4]
  wire [10:0] buffer_7_449; // @[Modules.scala 65:57:@17640.4]
  wire [10:0] buffer_7_116; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_117; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67104; // @[Modules.scala 65:57:@17642.4]
  wire [10:0] _T_67105; // @[Modules.scala 65:57:@17643.4]
  wire [10:0] buffer_7_450; // @[Modules.scala 65:57:@17644.4]
  wire [11:0] _T_67113; // @[Modules.scala 65:57:@17654.4]
  wire [10:0] _T_67114; // @[Modules.scala 65:57:@17655.4]
  wire [10:0] buffer_7_453; // @[Modules.scala 65:57:@17656.4]
  wire [11:0] _T_67131; // @[Modules.scala 65:57:@17678.4]
  wire [10:0] _T_67132; // @[Modules.scala 65:57:@17679.4]
  wire [10:0] buffer_7_459; // @[Modules.scala 65:57:@17680.4]
  wire [10:0] buffer_7_136; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67134; // @[Modules.scala 65:57:@17682.4]
  wire [10:0] _T_67135; // @[Modules.scala 65:57:@17683.4]
  wire [10:0] buffer_7_460; // @[Modules.scala 65:57:@17684.4]
  wire [10:0] buffer_7_142; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_143; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67143; // @[Modules.scala 65:57:@17694.4]
  wire [10:0] _T_67144; // @[Modules.scala 65:57:@17695.4]
  wire [10:0] buffer_7_463; // @[Modules.scala 65:57:@17696.4]
  wire [10:0] buffer_7_144; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67146; // @[Modules.scala 65:57:@17698.4]
  wire [10:0] _T_67147; // @[Modules.scala 65:57:@17699.4]
  wire [10:0] buffer_7_464; // @[Modules.scala 65:57:@17700.4]
  wire [10:0] buffer_7_146; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67149; // @[Modules.scala 65:57:@17702.4]
  wire [10:0] _T_67150; // @[Modules.scala 65:57:@17703.4]
  wire [10:0] buffer_7_465; // @[Modules.scala 65:57:@17704.4]
  wire [10:0] buffer_7_156; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67164; // @[Modules.scala 65:57:@17722.4]
  wire [10:0] _T_67165; // @[Modules.scala 65:57:@17723.4]
  wire [10:0] buffer_7_470; // @[Modules.scala 65:57:@17724.4]
  wire [11:0] _T_67167; // @[Modules.scala 65:57:@17726.4]
  wire [10:0] _T_67168; // @[Modules.scala 65:57:@17727.4]
  wire [10:0] buffer_7_471; // @[Modules.scala 65:57:@17728.4]
  wire [11:0] _T_67197; // @[Modules.scala 65:57:@17766.4]
  wire [10:0] _T_67198; // @[Modules.scala 65:57:@17767.4]
  wire [10:0] buffer_7_481; // @[Modules.scala 65:57:@17768.4]
  wire [10:0] buffer_7_182; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67203; // @[Modules.scala 65:57:@17774.4]
  wire [10:0] _T_67204; // @[Modules.scala 65:57:@17775.4]
  wire [10:0] buffer_7_483; // @[Modules.scala 65:57:@17776.4]
  wire [10:0] buffer_7_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67215; // @[Modules.scala 65:57:@17790.4]
  wire [10:0] _T_67216; // @[Modules.scala 65:57:@17791.4]
  wire [10:0] buffer_7_487; // @[Modules.scala 65:57:@17792.4]
  wire [11:0] _T_67224; // @[Modules.scala 65:57:@17802.4]
  wire [10:0] _T_67225; // @[Modules.scala 65:57:@17803.4]
  wire [10:0] buffer_7_490; // @[Modules.scala 65:57:@17804.4]
  wire [10:0] buffer_7_198; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_199; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67227; // @[Modules.scala 65:57:@17806.4]
  wire [10:0] _T_67228; // @[Modules.scala 65:57:@17807.4]
  wire [10:0] buffer_7_491; // @[Modules.scala 65:57:@17808.4]
  wire [11:0] _T_67230; // @[Modules.scala 65:57:@17810.4]
  wire [10:0] _T_67231; // @[Modules.scala 65:57:@17811.4]
  wire [10:0] buffer_7_492; // @[Modules.scala 65:57:@17812.4]
  wire [11:0] _T_67236; // @[Modules.scala 65:57:@17818.4]
  wire [10:0] _T_67237; // @[Modules.scala 65:57:@17819.4]
  wire [10:0] buffer_7_494; // @[Modules.scala 65:57:@17820.4]
  wire [11:0] _T_67245; // @[Modules.scala 65:57:@17830.4]
  wire [10:0] _T_67246; // @[Modules.scala 65:57:@17831.4]
  wire [10:0] buffer_7_497; // @[Modules.scala 65:57:@17832.4]
  wire [11:0] _T_67248; // @[Modules.scala 65:57:@17834.4]
  wire [10:0] _T_67249; // @[Modules.scala 65:57:@17835.4]
  wire [10:0] buffer_7_498; // @[Modules.scala 65:57:@17836.4]
  wire [11:0] _T_67251; // @[Modules.scala 65:57:@17838.4]
  wire [10:0] _T_67252; // @[Modules.scala 65:57:@17839.4]
  wire [10:0] buffer_7_499; // @[Modules.scala 65:57:@17840.4]
  wire [11:0] _T_67257; // @[Modules.scala 65:57:@17846.4]
  wire [10:0] _T_67258; // @[Modules.scala 65:57:@17847.4]
  wire [10:0] buffer_7_501; // @[Modules.scala 65:57:@17848.4]
  wire [10:0] buffer_7_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67266; // @[Modules.scala 65:57:@17858.4]
  wire [10:0] _T_67267; // @[Modules.scala 65:57:@17859.4]
  wire [10:0] buffer_7_504; // @[Modules.scala 65:57:@17860.4]
  wire [11:0] _T_67272; // @[Modules.scala 65:57:@17866.4]
  wire [10:0] _T_67273; // @[Modules.scala 65:57:@17867.4]
  wire [10:0] buffer_7_506; // @[Modules.scala 65:57:@17868.4]
  wire [10:0] buffer_7_234; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67281; // @[Modules.scala 65:57:@17878.4]
  wire [10:0] _T_67282; // @[Modules.scala 65:57:@17879.4]
  wire [10:0] buffer_7_509; // @[Modules.scala 65:57:@17880.4]
  wire [10:0] buffer_7_240; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67290; // @[Modules.scala 65:57:@17890.4]
  wire [10:0] _T_67291; // @[Modules.scala 65:57:@17891.4]
  wire [10:0] buffer_7_512; // @[Modules.scala 65:57:@17892.4]
  wire [11:0] _T_67299; // @[Modules.scala 65:57:@17902.4]
  wire [10:0] _T_67300; // @[Modules.scala 65:57:@17903.4]
  wire [10:0] buffer_7_515; // @[Modules.scala 65:57:@17904.4]
  wire [10:0] buffer_7_251; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67305; // @[Modules.scala 65:57:@17910.4]
  wire [10:0] _T_67306; // @[Modules.scala 65:57:@17911.4]
  wire [10:0] buffer_7_517; // @[Modules.scala 65:57:@17912.4]
  wire [11:0] _T_67320; // @[Modules.scala 65:57:@17930.4]
  wire [10:0] _T_67321; // @[Modules.scala 65:57:@17931.4]
  wire [10:0] buffer_7_522; // @[Modules.scala 65:57:@17932.4]
  wire [10:0] buffer_7_262; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_7_263; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67323; // @[Modules.scala 65:57:@17934.4]
  wire [10:0] _T_67324; // @[Modules.scala 65:57:@17935.4]
  wire [10:0] buffer_7_523; // @[Modules.scala 65:57:@17936.4]
  wire [10:0] buffer_7_269; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67332; // @[Modules.scala 65:57:@17946.4]
  wire [10:0] _T_67333; // @[Modules.scala 65:57:@17947.4]
  wire [10:0] buffer_7_526; // @[Modules.scala 65:57:@17948.4]
  wire [11:0] _T_67338; // @[Modules.scala 65:57:@17954.4]
  wire [10:0] _T_67339; // @[Modules.scala 65:57:@17955.4]
  wire [10:0] buffer_7_528; // @[Modules.scala 65:57:@17956.4]
  wire [11:0] _T_67341; // @[Modules.scala 65:57:@17958.4]
  wire [10:0] _T_67342; // @[Modules.scala 65:57:@17959.4]
  wire [10:0] buffer_7_529; // @[Modules.scala 65:57:@17960.4]
  wire [10:0] buffer_7_276; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67344; // @[Modules.scala 65:57:@17962.4]
  wire [10:0] _T_67345; // @[Modules.scala 65:57:@17963.4]
  wire [10:0] buffer_7_530; // @[Modules.scala 65:57:@17964.4]
  wire [11:0] _T_67353; // @[Modules.scala 65:57:@17974.4]
  wire [10:0] _T_67354; // @[Modules.scala 65:57:@17975.4]
  wire [10:0] buffer_7_533; // @[Modules.scala 65:57:@17976.4]
  wire [10:0] buffer_7_293; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67368; // @[Modules.scala 65:57:@17994.4]
  wire [10:0] _T_67369; // @[Modules.scala 65:57:@17995.4]
  wire [10:0] buffer_7_538; // @[Modules.scala 65:57:@17996.4]
  wire [10:0] buffer_7_299; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67377; // @[Modules.scala 65:57:@18006.4]
  wire [10:0] _T_67378; // @[Modules.scala 65:57:@18007.4]
  wire [10:0] buffer_7_541; // @[Modules.scala 65:57:@18008.4]
  wire [10:0] buffer_7_301; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67380; // @[Modules.scala 65:57:@18010.4]
  wire [10:0] _T_67381; // @[Modules.scala 65:57:@18011.4]
  wire [10:0] buffer_7_542; // @[Modules.scala 65:57:@18012.4]
  wire [11:0] _T_67389; // @[Modules.scala 65:57:@18022.4]
  wire [10:0] _T_67390; // @[Modules.scala 65:57:@18023.4]
  wire [10:0] buffer_7_545; // @[Modules.scala 65:57:@18024.4]
  wire [10:0] buffer_7_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67395; // @[Modules.scala 65:57:@18030.4]
  wire [10:0] _T_67396; // @[Modules.scala 65:57:@18031.4]
  wire [10:0] buffer_7_547; // @[Modules.scala 65:57:@18032.4]
  wire [11:0] _T_67398; // @[Modules.scala 65:57:@18034.4]
  wire [10:0] _T_67399; // @[Modules.scala 65:57:@18035.4]
  wire [10:0] buffer_7_548; // @[Modules.scala 65:57:@18036.4]
  wire [11:0] _T_67404; // @[Modules.scala 65:57:@18042.4]
  wire [10:0] _T_67405; // @[Modules.scala 65:57:@18043.4]
  wire [10:0] buffer_7_550; // @[Modules.scala 65:57:@18044.4]
  wire [11:0] _T_67413; // @[Modules.scala 65:57:@18054.4]
  wire [10:0] _T_67414; // @[Modules.scala 65:57:@18055.4]
  wire [10:0] buffer_7_553; // @[Modules.scala 65:57:@18056.4]
  wire [11:0] _T_67422; // @[Modules.scala 65:57:@18066.4]
  wire [10:0] _T_67423; // @[Modules.scala 65:57:@18067.4]
  wire [10:0] buffer_7_556; // @[Modules.scala 65:57:@18068.4]
  wire [11:0] _T_67428; // @[Modules.scala 65:57:@18074.4]
  wire [10:0] _T_67429; // @[Modules.scala 65:57:@18075.4]
  wire [10:0] buffer_7_558; // @[Modules.scala 65:57:@18076.4]
  wire [11:0] _T_67431; // @[Modules.scala 65:57:@18078.4]
  wire [10:0] _T_67432; // @[Modules.scala 65:57:@18079.4]
  wire [10:0] buffer_7_559; // @[Modules.scala 65:57:@18080.4]
  wire [11:0] _T_67434; // @[Modules.scala 65:57:@18082.4]
  wire [10:0] _T_67435; // @[Modules.scala 65:57:@18083.4]
  wire [10:0] buffer_7_560; // @[Modules.scala 65:57:@18084.4]
  wire [11:0] _T_67443; // @[Modules.scala 65:57:@18094.4]
  wire [10:0] _T_67444; // @[Modules.scala 65:57:@18095.4]
  wire [10:0] buffer_7_563; // @[Modules.scala 65:57:@18096.4]
  wire [10:0] buffer_7_345; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67446; // @[Modules.scala 65:57:@18098.4]
  wire [10:0] _T_67447; // @[Modules.scala 65:57:@18099.4]
  wire [10:0] buffer_7_564; // @[Modules.scala 65:57:@18100.4]
  wire [11:0] _T_67452; // @[Modules.scala 65:57:@18106.4]
  wire [10:0] _T_67453; // @[Modules.scala 65:57:@18107.4]
  wire [10:0] buffer_7_566; // @[Modules.scala 65:57:@18108.4]
  wire [11:0] _T_67473; // @[Modules.scala 65:57:@18134.4]
  wire [10:0] _T_67474; // @[Modules.scala 65:57:@18135.4]
  wire [10:0] buffer_7_573; // @[Modules.scala 65:57:@18136.4]
  wire [11:0] _T_67494; // @[Modules.scala 65:57:@18162.4]
  wire [10:0] _T_67495; // @[Modules.scala 65:57:@18163.4]
  wire [10:0] buffer_7_580; // @[Modules.scala 65:57:@18164.4]
  wire [10:0] buffer_7_380; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67500; // @[Modules.scala 65:57:@18170.4]
  wire [10:0] _T_67501; // @[Modules.scala 65:57:@18171.4]
  wire [10:0] buffer_7_582; // @[Modules.scala 65:57:@18172.4]
  wire [10:0] buffer_7_390; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_67515; // @[Modules.scala 65:57:@18190.4]
  wire [10:0] _T_67516; // @[Modules.scala 65:57:@18191.4]
  wire [10:0] buffer_7_587; // @[Modules.scala 65:57:@18192.4]
  wire [11:0] _T_67518; // @[Modules.scala 68:83:@18194.4]
  wire [10:0] _T_67519; // @[Modules.scala 68:83:@18195.4]
  wire [10:0] buffer_7_588; // @[Modules.scala 68:83:@18196.4]
  wire [11:0] _T_67524; // @[Modules.scala 68:83:@18202.4]
  wire [10:0] _T_67525; // @[Modules.scala 68:83:@18203.4]
  wire [10:0] buffer_7_590; // @[Modules.scala 68:83:@18204.4]
  wire [11:0] _T_67527; // @[Modules.scala 68:83:@18206.4]
  wire [10:0] _T_67528; // @[Modules.scala 68:83:@18207.4]
  wire [10:0] buffer_7_591; // @[Modules.scala 68:83:@18208.4]
  wire [11:0] _T_67530; // @[Modules.scala 68:83:@18210.4]
  wire [10:0] _T_67531; // @[Modules.scala 68:83:@18211.4]
  wire [10:0] buffer_7_592; // @[Modules.scala 68:83:@18212.4]
  wire [11:0] _T_67533; // @[Modules.scala 68:83:@18214.4]
  wire [10:0] _T_67534; // @[Modules.scala 68:83:@18215.4]
  wire [10:0] buffer_7_593; // @[Modules.scala 68:83:@18216.4]
  wire [11:0] _T_67536; // @[Modules.scala 68:83:@18218.4]
  wire [10:0] _T_67537; // @[Modules.scala 68:83:@18219.4]
  wire [10:0] buffer_7_594; // @[Modules.scala 68:83:@18220.4]
  wire [11:0] _T_67539; // @[Modules.scala 68:83:@18222.4]
  wire [10:0] _T_67540; // @[Modules.scala 68:83:@18223.4]
  wire [10:0] buffer_7_595; // @[Modules.scala 68:83:@18224.4]
  wire [11:0] _T_67548; // @[Modules.scala 68:83:@18234.4]
  wire [10:0] _T_67549; // @[Modules.scala 68:83:@18235.4]
  wire [10:0] buffer_7_598; // @[Modules.scala 68:83:@18236.4]
  wire [11:0] _T_67551; // @[Modules.scala 68:83:@18238.4]
  wire [10:0] _T_67552; // @[Modules.scala 68:83:@18239.4]
  wire [10:0] buffer_7_599; // @[Modules.scala 68:83:@18240.4]
  wire [11:0] _T_67554; // @[Modules.scala 68:83:@18242.4]
  wire [10:0] _T_67555; // @[Modules.scala 68:83:@18243.4]
  wire [10:0] buffer_7_600; // @[Modules.scala 68:83:@18244.4]
  wire [11:0] _T_67557; // @[Modules.scala 68:83:@18246.4]
  wire [10:0] _T_67558; // @[Modules.scala 68:83:@18247.4]
  wire [10:0] buffer_7_601; // @[Modules.scala 68:83:@18248.4]
  wire [11:0] _T_67560; // @[Modules.scala 68:83:@18250.4]
  wire [10:0] _T_67561; // @[Modules.scala 68:83:@18251.4]
  wire [10:0] buffer_7_602; // @[Modules.scala 68:83:@18252.4]
  wire [11:0] _T_67563; // @[Modules.scala 68:83:@18254.4]
  wire [10:0] _T_67564; // @[Modules.scala 68:83:@18255.4]
  wire [10:0] buffer_7_603; // @[Modules.scala 68:83:@18256.4]
  wire [11:0] _T_67566; // @[Modules.scala 68:83:@18258.4]
  wire [10:0] _T_67567; // @[Modules.scala 68:83:@18259.4]
  wire [10:0] buffer_7_604; // @[Modules.scala 68:83:@18260.4]
  wire [11:0] _T_67569; // @[Modules.scala 68:83:@18262.4]
  wire [10:0] _T_67570; // @[Modules.scala 68:83:@18263.4]
  wire [10:0] buffer_7_605; // @[Modules.scala 68:83:@18264.4]
  wire [11:0] _T_67572; // @[Modules.scala 68:83:@18266.4]
  wire [10:0] _T_67573; // @[Modules.scala 68:83:@18267.4]
  wire [10:0] buffer_7_606; // @[Modules.scala 68:83:@18268.4]
  wire [11:0] _T_67575; // @[Modules.scala 68:83:@18270.4]
  wire [10:0] _T_67576; // @[Modules.scala 68:83:@18271.4]
  wire [10:0] buffer_7_607; // @[Modules.scala 68:83:@18272.4]
  wire [11:0] _T_67581; // @[Modules.scala 68:83:@18278.4]
  wire [10:0] _T_67582; // @[Modules.scala 68:83:@18279.4]
  wire [10:0] buffer_7_609; // @[Modules.scala 68:83:@18280.4]
  wire [11:0] _T_67584; // @[Modules.scala 68:83:@18282.4]
  wire [10:0] _T_67585; // @[Modules.scala 68:83:@18283.4]
  wire [10:0] buffer_7_610; // @[Modules.scala 68:83:@18284.4]
  wire [11:0] _T_67587; // @[Modules.scala 68:83:@18286.4]
  wire [10:0] _T_67588; // @[Modules.scala 68:83:@18287.4]
  wire [10:0] buffer_7_611; // @[Modules.scala 68:83:@18288.4]
  wire [11:0] _T_67590; // @[Modules.scala 68:83:@18290.4]
  wire [10:0] _T_67591; // @[Modules.scala 68:83:@18291.4]
  wire [10:0] buffer_7_612; // @[Modules.scala 68:83:@18292.4]
  wire [11:0] _T_67593; // @[Modules.scala 68:83:@18294.4]
  wire [10:0] _T_67594; // @[Modules.scala 68:83:@18295.4]
  wire [10:0] buffer_7_613; // @[Modules.scala 68:83:@18296.4]
  wire [11:0] _T_67599; // @[Modules.scala 68:83:@18302.4]
  wire [10:0] _T_67600; // @[Modules.scala 68:83:@18303.4]
  wire [10:0] buffer_7_615; // @[Modules.scala 68:83:@18304.4]
  wire [11:0] _T_67602; // @[Modules.scala 68:83:@18306.4]
  wire [10:0] _T_67603; // @[Modules.scala 68:83:@18307.4]
  wire [10:0] buffer_7_616; // @[Modules.scala 68:83:@18308.4]
  wire [11:0] _T_67605; // @[Modules.scala 68:83:@18310.4]
  wire [10:0] _T_67606; // @[Modules.scala 68:83:@18311.4]
  wire [10:0] buffer_7_617; // @[Modules.scala 68:83:@18312.4]
  wire [11:0] _T_67608; // @[Modules.scala 68:83:@18314.4]
  wire [10:0] _T_67609; // @[Modules.scala 68:83:@18315.4]
  wire [10:0] buffer_7_618; // @[Modules.scala 68:83:@18316.4]
  wire [11:0] _T_67617; // @[Modules.scala 68:83:@18326.4]
  wire [10:0] _T_67618; // @[Modules.scala 68:83:@18327.4]
  wire [10:0] buffer_7_621; // @[Modules.scala 68:83:@18328.4]
  wire [11:0] _T_67620; // @[Modules.scala 68:83:@18330.4]
  wire [10:0] _T_67621; // @[Modules.scala 68:83:@18331.4]
  wire [10:0] buffer_7_622; // @[Modules.scala 68:83:@18332.4]
  wire [11:0] _T_67623; // @[Modules.scala 68:83:@18334.4]
  wire [10:0] _T_67624; // @[Modules.scala 68:83:@18335.4]
  wire [10:0] buffer_7_623; // @[Modules.scala 68:83:@18336.4]
  wire [11:0] _T_67626; // @[Modules.scala 68:83:@18338.4]
  wire [10:0] _T_67627; // @[Modules.scala 68:83:@18339.4]
  wire [10:0] buffer_7_624; // @[Modules.scala 68:83:@18340.4]
  wire [11:0] _T_67635; // @[Modules.scala 68:83:@18350.4]
  wire [10:0] _T_67636; // @[Modules.scala 68:83:@18351.4]
  wire [10:0] buffer_7_627; // @[Modules.scala 68:83:@18352.4]
  wire [11:0] _T_67644; // @[Modules.scala 68:83:@18362.4]
  wire [10:0] _T_67645; // @[Modules.scala 68:83:@18363.4]
  wire [10:0] buffer_7_630; // @[Modules.scala 68:83:@18364.4]
  wire [11:0] _T_67650; // @[Modules.scala 68:83:@18370.4]
  wire [10:0] _T_67651; // @[Modules.scala 68:83:@18371.4]
  wire [10:0] buffer_7_632; // @[Modules.scala 68:83:@18372.4]
  wire [11:0] _T_67653; // @[Modules.scala 68:83:@18374.4]
  wire [10:0] _T_67654; // @[Modules.scala 68:83:@18375.4]
  wire [10:0] buffer_7_633; // @[Modules.scala 68:83:@18376.4]
  wire [11:0] _T_67659; // @[Modules.scala 68:83:@18382.4]
  wire [10:0] _T_67660; // @[Modules.scala 68:83:@18383.4]
  wire [10:0] buffer_7_635; // @[Modules.scala 68:83:@18384.4]
  wire [11:0] _T_67665; // @[Modules.scala 68:83:@18390.4]
  wire [10:0] _T_67666; // @[Modules.scala 68:83:@18391.4]
  wire [10:0] buffer_7_637; // @[Modules.scala 68:83:@18392.4]
  wire [11:0] _T_67668; // @[Modules.scala 68:83:@18394.4]
  wire [10:0] _T_67669; // @[Modules.scala 68:83:@18395.4]
  wire [10:0] buffer_7_638; // @[Modules.scala 68:83:@18396.4]
  wire [11:0] _T_67671; // @[Modules.scala 68:83:@18398.4]
  wire [10:0] _T_67672; // @[Modules.scala 68:83:@18399.4]
  wire [10:0] buffer_7_639; // @[Modules.scala 68:83:@18400.4]
  wire [11:0] _T_67674; // @[Modules.scala 68:83:@18402.4]
  wire [10:0] _T_67675; // @[Modules.scala 68:83:@18403.4]
  wire [10:0] buffer_7_640; // @[Modules.scala 68:83:@18404.4]
  wire [11:0] _T_67677; // @[Modules.scala 68:83:@18406.4]
  wire [10:0] _T_67678; // @[Modules.scala 68:83:@18407.4]
  wire [10:0] buffer_7_641; // @[Modules.scala 68:83:@18408.4]
  wire [11:0] _T_67680; // @[Modules.scala 68:83:@18410.4]
  wire [10:0] _T_67681; // @[Modules.scala 68:83:@18411.4]
  wire [10:0] buffer_7_642; // @[Modules.scala 68:83:@18412.4]
  wire [11:0] _T_67683; // @[Modules.scala 68:83:@18414.4]
  wire [10:0] _T_67684; // @[Modules.scala 68:83:@18415.4]
  wire [10:0] buffer_7_643; // @[Modules.scala 68:83:@18416.4]
  wire [11:0] _T_67686; // @[Modules.scala 68:83:@18418.4]
  wire [10:0] _T_67687; // @[Modules.scala 68:83:@18419.4]
  wire [10:0] buffer_7_644; // @[Modules.scala 68:83:@18420.4]
  wire [11:0] _T_67689; // @[Modules.scala 68:83:@18422.4]
  wire [10:0] _T_67690; // @[Modules.scala 68:83:@18423.4]
  wire [10:0] buffer_7_645; // @[Modules.scala 68:83:@18424.4]
  wire [11:0] _T_67692; // @[Modules.scala 68:83:@18426.4]
  wire [10:0] _T_67693; // @[Modules.scala 68:83:@18427.4]
  wire [10:0] buffer_7_646; // @[Modules.scala 68:83:@18428.4]
  wire [11:0] _T_67695; // @[Modules.scala 68:83:@18430.4]
  wire [10:0] _T_67696; // @[Modules.scala 68:83:@18431.4]
  wire [10:0] buffer_7_647; // @[Modules.scala 68:83:@18432.4]
  wire [11:0] _T_67698; // @[Modules.scala 68:83:@18434.4]
  wire [10:0] _T_67699; // @[Modules.scala 68:83:@18435.4]
  wire [10:0] buffer_7_648; // @[Modules.scala 68:83:@18436.4]
  wire [11:0] _T_67701; // @[Modules.scala 68:83:@18438.4]
  wire [10:0] _T_67702; // @[Modules.scala 68:83:@18439.4]
  wire [10:0] buffer_7_649; // @[Modules.scala 68:83:@18440.4]
  wire [11:0] _T_67704; // @[Modules.scala 68:83:@18442.4]
  wire [10:0] _T_67705; // @[Modules.scala 68:83:@18443.4]
  wire [10:0] buffer_7_650; // @[Modules.scala 68:83:@18444.4]
  wire [11:0] _T_67707; // @[Modules.scala 68:83:@18446.4]
  wire [10:0] _T_67708; // @[Modules.scala 68:83:@18447.4]
  wire [10:0] buffer_7_651; // @[Modules.scala 68:83:@18448.4]
  wire [11:0] _T_67710; // @[Modules.scala 68:83:@18450.4]
  wire [10:0] _T_67711; // @[Modules.scala 68:83:@18451.4]
  wire [10:0] buffer_7_652; // @[Modules.scala 68:83:@18452.4]
  wire [11:0] _T_67713; // @[Modules.scala 68:83:@18454.4]
  wire [10:0] _T_67714; // @[Modules.scala 68:83:@18455.4]
  wire [10:0] buffer_7_653; // @[Modules.scala 68:83:@18456.4]
  wire [11:0] _T_67716; // @[Modules.scala 68:83:@18458.4]
  wire [10:0] _T_67717; // @[Modules.scala 68:83:@18459.4]
  wire [10:0] buffer_7_654; // @[Modules.scala 68:83:@18460.4]
  wire [11:0] _T_67719; // @[Modules.scala 68:83:@18462.4]
  wire [10:0] _T_67720; // @[Modules.scala 68:83:@18463.4]
  wire [10:0] buffer_7_655; // @[Modules.scala 68:83:@18464.4]
  wire [11:0] _T_67722; // @[Modules.scala 68:83:@18466.4]
  wire [10:0] _T_67723; // @[Modules.scala 68:83:@18467.4]
  wire [10:0] buffer_7_656; // @[Modules.scala 68:83:@18468.4]
  wire [11:0] _T_67725; // @[Modules.scala 68:83:@18470.4]
  wire [10:0] _T_67726; // @[Modules.scala 68:83:@18471.4]
  wire [10:0] buffer_7_657; // @[Modules.scala 68:83:@18472.4]
  wire [11:0] _T_67728; // @[Modules.scala 68:83:@18474.4]
  wire [10:0] _T_67729; // @[Modules.scala 68:83:@18475.4]
  wire [10:0] buffer_7_658; // @[Modules.scala 68:83:@18476.4]
  wire [11:0] _T_67734; // @[Modules.scala 68:83:@18482.4]
  wire [10:0] _T_67735; // @[Modules.scala 68:83:@18483.4]
  wire [10:0] buffer_7_660; // @[Modules.scala 68:83:@18484.4]
  wire [11:0] _T_67737; // @[Modules.scala 68:83:@18486.4]
  wire [10:0] _T_67738; // @[Modules.scala 68:83:@18487.4]
  wire [10:0] buffer_7_661; // @[Modules.scala 68:83:@18488.4]
  wire [11:0] _T_67740; // @[Modules.scala 68:83:@18490.4]
  wire [10:0] _T_67741; // @[Modules.scala 68:83:@18491.4]
  wire [10:0] buffer_7_662; // @[Modules.scala 68:83:@18492.4]
  wire [11:0] _T_67743; // @[Modules.scala 68:83:@18494.4]
  wire [10:0] _T_67744; // @[Modules.scala 68:83:@18495.4]
  wire [10:0] buffer_7_663; // @[Modules.scala 68:83:@18496.4]
  wire [11:0] _T_67746; // @[Modules.scala 68:83:@18498.4]
  wire [10:0] _T_67747; // @[Modules.scala 68:83:@18499.4]
  wire [10:0] buffer_7_664; // @[Modules.scala 68:83:@18500.4]
  wire [11:0] _T_67749; // @[Modules.scala 68:83:@18502.4]
  wire [10:0] _T_67750; // @[Modules.scala 68:83:@18503.4]
  wire [10:0] buffer_7_665; // @[Modules.scala 68:83:@18504.4]
  wire [11:0] _T_67752; // @[Modules.scala 68:83:@18506.4]
  wire [10:0] _T_67753; // @[Modules.scala 68:83:@18507.4]
  wire [10:0] buffer_7_666; // @[Modules.scala 68:83:@18508.4]
  wire [11:0] _T_67755; // @[Modules.scala 68:83:@18510.4]
  wire [10:0] _T_67756; // @[Modules.scala 68:83:@18511.4]
  wire [10:0] buffer_7_667; // @[Modules.scala 68:83:@18512.4]
  wire [11:0] _T_67758; // @[Modules.scala 68:83:@18514.4]
  wire [10:0] _T_67759; // @[Modules.scala 68:83:@18515.4]
  wire [10:0] buffer_7_668; // @[Modules.scala 68:83:@18516.4]
  wire [11:0] _T_67761; // @[Modules.scala 68:83:@18518.4]
  wire [10:0] _T_67762; // @[Modules.scala 68:83:@18519.4]
  wire [10:0] buffer_7_669; // @[Modules.scala 68:83:@18520.4]
  wire [11:0] _T_67764; // @[Modules.scala 68:83:@18522.4]
  wire [10:0] _T_67765; // @[Modules.scala 68:83:@18523.4]
  wire [10:0] buffer_7_670; // @[Modules.scala 68:83:@18524.4]
  wire [11:0] _T_67767; // @[Modules.scala 68:83:@18526.4]
  wire [10:0] _T_67768; // @[Modules.scala 68:83:@18527.4]
  wire [10:0] buffer_7_671; // @[Modules.scala 68:83:@18528.4]
  wire [11:0] _T_67770; // @[Modules.scala 68:83:@18530.4]
  wire [10:0] _T_67771; // @[Modules.scala 68:83:@18531.4]
  wire [10:0] buffer_7_672; // @[Modules.scala 68:83:@18532.4]
  wire [11:0] _T_67773; // @[Modules.scala 68:83:@18534.4]
  wire [10:0] _T_67774; // @[Modules.scala 68:83:@18535.4]
  wire [10:0] buffer_7_673; // @[Modules.scala 68:83:@18536.4]
  wire [11:0] _T_67776; // @[Modules.scala 68:83:@18538.4]
  wire [10:0] _T_67777; // @[Modules.scala 68:83:@18539.4]
  wire [10:0] buffer_7_674; // @[Modules.scala 68:83:@18540.4]
  wire [11:0] _T_67779; // @[Modules.scala 68:83:@18542.4]
  wire [10:0] _T_67780; // @[Modules.scala 68:83:@18543.4]
  wire [10:0] buffer_7_675; // @[Modules.scala 68:83:@18544.4]
  wire [11:0] _T_67788; // @[Modules.scala 68:83:@18554.4]
  wire [10:0] _T_67789; // @[Modules.scala 68:83:@18555.4]
  wire [10:0] buffer_7_678; // @[Modules.scala 68:83:@18556.4]
  wire [11:0] _T_67800; // @[Modules.scala 68:83:@18570.4]
  wire [10:0] _T_67801; // @[Modules.scala 68:83:@18571.4]
  wire [10:0] buffer_7_682; // @[Modules.scala 68:83:@18572.4]
  wire [11:0] _T_67803; // @[Modules.scala 68:83:@18574.4]
  wire [10:0] _T_67804; // @[Modules.scala 68:83:@18575.4]
  wire [10:0] buffer_7_683; // @[Modules.scala 68:83:@18576.4]
  wire [11:0] _T_67809; // @[Modules.scala 68:83:@18582.4]
  wire [10:0] _T_67810; // @[Modules.scala 68:83:@18583.4]
  wire [10:0] buffer_7_685; // @[Modules.scala 68:83:@18584.4]
  wire [11:0] _T_67812; // @[Modules.scala 71:109:@18586.4]
  wire [10:0] _T_67813; // @[Modules.scala 71:109:@18587.4]
  wire [10:0] buffer_7_686; // @[Modules.scala 71:109:@18588.4]
  wire [11:0] _T_67815; // @[Modules.scala 71:109:@18590.4]
  wire [10:0] _T_67816; // @[Modules.scala 71:109:@18591.4]
  wire [10:0] buffer_7_687; // @[Modules.scala 71:109:@18592.4]
  wire [11:0] _T_67818; // @[Modules.scala 71:109:@18594.4]
  wire [10:0] _T_67819; // @[Modules.scala 71:109:@18595.4]
  wire [10:0] buffer_7_688; // @[Modules.scala 71:109:@18596.4]
  wire [11:0] _T_67821; // @[Modules.scala 71:109:@18598.4]
  wire [10:0] _T_67822; // @[Modules.scala 71:109:@18599.4]
  wire [10:0] buffer_7_689; // @[Modules.scala 71:109:@18600.4]
  wire [11:0] _T_67827; // @[Modules.scala 71:109:@18606.4]
  wire [10:0] _T_67828; // @[Modules.scala 71:109:@18607.4]
  wire [10:0] buffer_7_691; // @[Modules.scala 71:109:@18608.4]
  wire [11:0] _T_67830; // @[Modules.scala 71:109:@18610.4]
  wire [10:0] _T_67831; // @[Modules.scala 71:109:@18611.4]
  wire [10:0] buffer_7_692; // @[Modules.scala 71:109:@18612.4]
  wire [11:0] _T_67833; // @[Modules.scala 71:109:@18614.4]
  wire [10:0] _T_67834; // @[Modules.scala 71:109:@18615.4]
  wire [10:0] buffer_7_693; // @[Modules.scala 71:109:@18616.4]
  wire [11:0] _T_67836; // @[Modules.scala 71:109:@18618.4]
  wire [10:0] _T_67837; // @[Modules.scala 71:109:@18619.4]
  wire [10:0] buffer_7_694; // @[Modules.scala 71:109:@18620.4]
  wire [11:0] _T_67839; // @[Modules.scala 71:109:@18622.4]
  wire [10:0] _T_67840; // @[Modules.scala 71:109:@18623.4]
  wire [10:0] buffer_7_695; // @[Modules.scala 71:109:@18624.4]
  wire [11:0] _T_67842; // @[Modules.scala 71:109:@18626.4]
  wire [10:0] _T_67843; // @[Modules.scala 71:109:@18627.4]
  wire [10:0] buffer_7_696; // @[Modules.scala 71:109:@18628.4]
  wire [11:0] _T_67845; // @[Modules.scala 71:109:@18630.4]
  wire [10:0] _T_67846; // @[Modules.scala 71:109:@18631.4]
  wire [10:0] buffer_7_697; // @[Modules.scala 71:109:@18632.4]
  wire [11:0] _T_67848; // @[Modules.scala 71:109:@18634.4]
  wire [10:0] _T_67849; // @[Modules.scala 71:109:@18635.4]
  wire [10:0] buffer_7_698; // @[Modules.scala 71:109:@18636.4]
  wire [11:0] _T_67851; // @[Modules.scala 71:109:@18638.4]
  wire [10:0] _T_67852; // @[Modules.scala 71:109:@18639.4]
  wire [10:0] buffer_7_699; // @[Modules.scala 71:109:@18640.4]
  wire [11:0] _T_67854; // @[Modules.scala 71:109:@18642.4]
  wire [10:0] _T_67855; // @[Modules.scala 71:109:@18643.4]
  wire [10:0] buffer_7_700; // @[Modules.scala 71:109:@18644.4]
  wire [11:0] _T_67857; // @[Modules.scala 71:109:@18646.4]
  wire [10:0] _T_67858; // @[Modules.scala 71:109:@18647.4]
  wire [10:0] buffer_7_701; // @[Modules.scala 71:109:@18648.4]
  wire [11:0] _T_67860; // @[Modules.scala 71:109:@18650.4]
  wire [10:0] _T_67861; // @[Modules.scala 71:109:@18651.4]
  wire [10:0] buffer_7_702; // @[Modules.scala 71:109:@18652.4]
  wire [11:0] _T_67863; // @[Modules.scala 71:109:@18654.4]
  wire [10:0] _T_67864; // @[Modules.scala 71:109:@18655.4]
  wire [10:0] buffer_7_703; // @[Modules.scala 71:109:@18656.4]
  wire [11:0] _T_67866; // @[Modules.scala 71:109:@18658.4]
  wire [10:0] _T_67867; // @[Modules.scala 71:109:@18659.4]
  wire [10:0] buffer_7_704; // @[Modules.scala 71:109:@18660.4]
  wire [11:0] _T_67869; // @[Modules.scala 71:109:@18662.4]
  wire [10:0] _T_67870; // @[Modules.scala 71:109:@18663.4]
  wire [10:0] buffer_7_705; // @[Modules.scala 71:109:@18664.4]
  wire [11:0] _T_67872; // @[Modules.scala 71:109:@18666.4]
  wire [10:0] _T_67873; // @[Modules.scala 71:109:@18667.4]
  wire [10:0] buffer_7_706; // @[Modules.scala 71:109:@18668.4]
  wire [11:0] _T_67875; // @[Modules.scala 71:109:@18670.4]
  wire [10:0] _T_67876; // @[Modules.scala 71:109:@18671.4]
  wire [10:0] buffer_7_707; // @[Modules.scala 71:109:@18672.4]
  wire [11:0] _T_67878; // @[Modules.scala 71:109:@18674.4]
  wire [10:0] _T_67879; // @[Modules.scala 71:109:@18675.4]
  wire [10:0] buffer_7_708; // @[Modules.scala 71:109:@18676.4]
  wire [11:0] _T_67881; // @[Modules.scala 71:109:@18678.4]
  wire [10:0] _T_67882; // @[Modules.scala 71:109:@18679.4]
  wire [10:0] buffer_7_709; // @[Modules.scala 71:109:@18680.4]
  wire [11:0] _T_67884; // @[Modules.scala 71:109:@18682.4]
  wire [10:0] _T_67885; // @[Modules.scala 71:109:@18683.4]
  wire [10:0] buffer_7_710; // @[Modules.scala 71:109:@18684.4]
  wire [11:0] _T_67887; // @[Modules.scala 71:109:@18686.4]
  wire [10:0] _T_67888; // @[Modules.scala 71:109:@18687.4]
  wire [10:0] buffer_7_711; // @[Modules.scala 71:109:@18688.4]
  wire [11:0] _T_67890; // @[Modules.scala 71:109:@18690.4]
  wire [10:0] _T_67891; // @[Modules.scala 71:109:@18691.4]
  wire [10:0] buffer_7_712; // @[Modules.scala 71:109:@18692.4]
  wire [11:0] _T_67893; // @[Modules.scala 71:109:@18694.4]
  wire [10:0] _T_67894; // @[Modules.scala 71:109:@18695.4]
  wire [10:0] buffer_7_713; // @[Modules.scala 71:109:@18696.4]
  wire [11:0] _T_67896; // @[Modules.scala 71:109:@18698.4]
  wire [10:0] _T_67897; // @[Modules.scala 71:109:@18699.4]
  wire [10:0] buffer_7_714; // @[Modules.scala 71:109:@18700.4]
  wire [11:0] _T_67899; // @[Modules.scala 71:109:@18702.4]
  wire [10:0] _T_67900; // @[Modules.scala 71:109:@18703.4]
  wire [10:0] buffer_7_715; // @[Modules.scala 71:109:@18704.4]
  wire [11:0] _T_67902; // @[Modules.scala 71:109:@18706.4]
  wire [10:0] _T_67903; // @[Modules.scala 71:109:@18707.4]
  wire [10:0] buffer_7_716; // @[Modules.scala 71:109:@18708.4]
  wire [11:0] _T_67905; // @[Modules.scala 71:109:@18710.4]
  wire [10:0] _T_67906; // @[Modules.scala 71:109:@18711.4]
  wire [10:0] buffer_7_717; // @[Modules.scala 71:109:@18712.4]
  wire [11:0] _T_67908; // @[Modules.scala 71:109:@18714.4]
  wire [10:0] _T_67909; // @[Modules.scala 71:109:@18715.4]
  wire [10:0] buffer_7_718; // @[Modules.scala 71:109:@18716.4]
  wire [11:0] _T_67911; // @[Modules.scala 71:109:@18718.4]
  wire [10:0] _T_67912; // @[Modules.scala 71:109:@18719.4]
  wire [10:0] buffer_7_719; // @[Modules.scala 71:109:@18720.4]
  wire [11:0] _T_67914; // @[Modules.scala 71:109:@18722.4]
  wire [10:0] _T_67915; // @[Modules.scala 71:109:@18723.4]
  wire [10:0] buffer_7_720; // @[Modules.scala 71:109:@18724.4]
  wire [11:0] _T_67917; // @[Modules.scala 71:109:@18726.4]
  wire [10:0] _T_67918; // @[Modules.scala 71:109:@18727.4]
  wire [10:0] buffer_7_721; // @[Modules.scala 71:109:@18728.4]
  wire [11:0] _T_67920; // @[Modules.scala 71:109:@18730.4]
  wire [10:0] _T_67921; // @[Modules.scala 71:109:@18731.4]
  wire [10:0] buffer_7_722; // @[Modules.scala 71:109:@18732.4]
  wire [11:0] _T_67923; // @[Modules.scala 71:109:@18734.4]
  wire [10:0] _T_67924; // @[Modules.scala 71:109:@18735.4]
  wire [10:0] buffer_7_723; // @[Modules.scala 71:109:@18736.4]
  wire [11:0] _T_67926; // @[Modules.scala 71:109:@18738.4]
  wire [10:0] _T_67927; // @[Modules.scala 71:109:@18739.4]
  wire [10:0] buffer_7_724; // @[Modules.scala 71:109:@18740.4]
  wire [11:0] _T_67929; // @[Modules.scala 71:109:@18742.4]
  wire [10:0] _T_67930; // @[Modules.scala 71:109:@18743.4]
  wire [10:0] buffer_7_725; // @[Modules.scala 71:109:@18744.4]
  wire [11:0] _T_67932; // @[Modules.scala 71:109:@18746.4]
  wire [10:0] _T_67933; // @[Modules.scala 71:109:@18747.4]
  wire [10:0] buffer_7_726; // @[Modules.scala 71:109:@18748.4]
  wire [11:0] _T_67935; // @[Modules.scala 71:109:@18750.4]
  wire [10:0] _T_67936; // @[Modules.scala 71:109:@18751.4]
  wire [10:0] buffer_7_727; // @[Modules.scala 71:109:@18752.4]
  wire [11:0] _T_67938; // @[Modules.scala 71:109:@18754.4]
  wire [10:0] _T_67939; // @[Modules.scala 71:109:@18755.4]
  wire [10:0] buffer_7_728; // @[Modules.scala 71:109:@18756.4]
  wire [11:0] _T_67941; // @[Modules.scala 71:109:@18758.4]
  wire [10:0] _T_67942; // @[Modules.scala 71:109:@18759.4]
  wire [10:0] buffer_7_729; // @[Modules.scala 71:109:@18760.4]
  wire [11:0] _T_67947; // @[Modules.scala 71:109:@18766.4]
  wire [10:0] _T_67948; // @[Modules.scala 71:109:@18767.4]
  wire [10:0] buffer_7_731; // @[Modules.scala 71:109:@18768.4]
  wire [11:0] _T_67953; // @[Modules.scala 71:109:@18774.4]
  wire [10:0] _T_67954; // @[Modules.scala 71:109:@18775.4]
  wire [10:0] buffer_7_733; // @[Modules.scala 71:109:@18776.4]
  wire [11:0] _T_67956; // @[Modules.scala 71:109:@18778.4]
  wire [10:0] _T_67957; // @[Modules.scala 71:109:@18779.4]
  wire [10:0] buffer_7_734; // @[Modules.scala 71:109:@18780.4]
  wire [11:0] _T_67959; // @[Modules.scala 78:156:@18783.4]
  wire [10:0] _T_67960; // @[Modules.scala 78:156:@18784.4]
  wire [10:0] buffer_7_736; // @[Modules.scala 78:156:@18785.4]
  wire [11:0] _T_67962; // @[Modules.scala 78:156:@18787.4]
  wire [10:0] _T_67963; // @[Modules.scala 78:156:@18788.4]
  wire [10:0] buffer_7_737; // @[Modules.scala 78:156:@18789.4]
  wire [11:0] _T_67965; // @[Modules.scala 78:156:@18791.4]
  wire [10:0] _T_67966; // @[Modules.scala 78:156:@18792.4]
  wire [10:0] buffer_7_738; // @[Modules.scala 78:156:@18793.4]
  wire [11:0] _T_67968; // @[Modules.scala 78:156:@18795.4]
  wire [10:0] _T_67969; // @[Modules.scala 78:156:@18796.4]
  wire [10:0] buffer_7_739; // @[Modules.scala 78:156:@18797.4]
  wire [11:0] _T_67971; // @[Modules.scala 78:156:@18799.4]
  wire [10:0] _T_67972; // @[Modules.scala 78:156:@18800.4]
  wire [10:0] buffer_7_740; // @[Modules.scala 78:156:@18801.4]
  wire [11:0] _T_67974; // @[Modules.scala 78:156:@18803.4]
  wire [10:0] _T_67975; // @[Modules.scala 78:156:@18804.4]
  wire [10:0] buffer_7_741; // @[Modules.scala 78:156:@18805.4]
  wire [11:0] _T_67977; // @[Modules.scala 78:156:@18807.4]
  wire [10:0] _T_67978; // @[Modules.scala 78:156:@18808.4]
  wire [10:0] buffer_7_742; // @[Modules.scala 78:156:@18809.4]
  wire [11:0] _T_67980; // @[Modules.scala 78:156:@18811.4]
  wire [10:0] _T_67981; // @[Modules.scala 78:156:@18812.4]
  wire [10:0] buffer_7_743; // @[Modules.scala 78:156:@18813.4]
  wire [11:0] _T_67983; // @[Modules.scala 78:156:@18815.4]
  wire [10:0] _T_67984; // @[Modules.scala 78:156:@18816.4]
  wire [10:0] buffer_7_744; // @[Modules.scala 78:156:@18817.4]
  wire [11:0] _T_67986; // @[Modules.scala 78:156:@18819.4]
  wire [10:0] _T_67987; // @[Modules.scala 78:156:@18820.4]
  wire [10:0] buffer_7_745; // @[Modules.scala 78:156:@18821.4]
  wire [11:0] _T_67989; // @[Modules.scala 78:156:@18823.4]
  wire [10:0] _T_67990; // @[Modules.scala 78:156:@18824.4]
  wire [10:0] buffer_7_746; // @[Modules.scala 78:156:@18825.4]
  wire [11:0] _T_67992; // @[Modules.scala 78:156:@18827.4]
  wire [10:0] _T_67993; // @[Modules.scala 78:156:@18828.4]
  wire [10:0] buffer_7_747; // @[Modules.scala 78:156:@18829.4]
  wire [11:0] _T_67995; // @[Modules.scala 78:156:@18831.4]
  wire [10:0] _T_67996; // @[Modules.scala 78:156:@18832.4]
  wire [10:0] buffer_7_748; // @[Modules.scala 78:156:@18833.4]
  wire [11:0] _T_67998; // @[Modules.scala 78:156:@18835.4]
  wire [10:0] _T_67999; // @[Modules.scala 78:156:@18836.4]
  wire [10:0] buffer_7_749; // @[Modules.scala 78:156:@18837.4]
  wire [11:0] _T_68001; // @[Modules.scala 78:156:@18839.4]
  wire [10:0] _T_68002; // @[Modules.scala 78:156:@18840.4]
  wire [10:0] buffer_7_750; // @[Modules.scala 78:156:@18841.4]
  wire [11:0] _T_68004; // @[Modules.scala 78:156:@18843.4]
  wire [10:0] _T_68005; // @[Modules.scala 78:156:@18844.4]
  wire [10:0] buffer_7_751; // @[Modules.scala 78:156:@18845.4]
  wire [11:0] _T_68007; // @[Modules.scala 78:156:@18847.4]
  wire [10:0] _T_68008; // @[Modules.scala 78:156:@18848.4]
  wire [10:0] buffer_7_752; // @[Modules.scala 78:156:@18849.4]
  wire [11:0] _T_68010; // @[Modules.scala 78:156:@18851.4]
  wire [10:0] _T_68011; // @[Modules.scala 78:156:@18852.4]
  wire [10:0] buffer_7_753; // @[Modules.scala 78:156:@18853.4]
  wire [11:0] _T_68013; // @[Modules.scala 78:156:@18855.4]
  wire [10:0] _T_68014; // @[Modules.scala 78:156:@18856.4]
  wire [10:0] buffer_7_754; // @[Modules.scala 78:156:@18857.4]
  wire [11:0] _T_68016; // @[Modules.scala 78:156:@18859.4]
  wire [10:0] _T_68017; // @[Modules.scala 78:156:@18860.4]
  wire [10:0] buffer_7_755; // @[Modules.scala 78:156:@18861.4]
  wire [11:0] _T_68019; // @[Modules.scala 78:156:@18863.4]
  wire [10:0] _T_68020; // @[Modules.scala 78:156:@18864.4]
  wire [10:0] buffer_7_756; // @[Modules.scala 78:156:@18865.4]
  wire [11:0] _T_68022; // @[Modules.scala 78:156:@18867.4]
  wire [10:0] _T_68023; // @[Modules.scala 78:156:@18868.4]
  wire [10:0] buffer_7_757; // @[Modules.scala 78:156:@18869.4]
  wire [11:0] _T_68025; // @[Modules.scala 78:156:@18871.4]
  wire [10:0] _T_68026; // @[Modules.scala 78:156:@18872.4]
  wire [10:0] buffer_7_758; // @[Modules.scala 78:156:@18873.4]
  wire [11:0] _T_68028; // @[Modules.scala 78:156:@18875.4]
  wire [10:0] _T_68029; // @[Modules.scala 78:156:@18876.4]
  wire [10:0] buffer_7_759; // @[Modules.scala 78:156:@18877.4]
  wire [11:0] _T_68031; // @[Modules.scala 78:156:@18879.4]
  wire [10:0] _T_68032; // @[Modules.scala 78:156:@18880.4]
  wire [10:0] buffer_7_760; // @[Modules.scala 78:156:@18881.4]
  wire [11:0] _T_68034; // @[Modules.scala 78:156:@18883.4]
  wire [10:0] _T_68035; // @[Modules.scala 78:156:@18884.4]
  wire [10:0] buffer_7_761; // @[Modules.scala 78:156:@18885.4]
  wire [11:0] _T_68037; // @[Modules.scala 78:156:@18887.4]
  wire [10:0] _T_68038; // @[Modules.scala 78:156:@18888.4]
  wire [10:0] buffer_7_762; // @[Modules.scala 78:156:@18889.4]
  wire [11:0] _T_68040; // @[Modules.scala 78:156:@18891.4]
  wire [10:0] _T_68041; // @[Modules.scala 78:156:@18892.4]
  wire [10:0] buffer_7_763; // @[Modules.scala 78:156:@18893.4]
  wire [11:0] _T_68043; // @[Modules.scala 78:156:@18895.4]
  wire [10:0] _T_68044; // @[Modules.scala 78:156:@18896.4]
  wire [10:0] buffer_7_764; // @[Modules.scala 78:156:@18897.4]
  wire [11:0] _T_68046; // @[Modules.scala 78:156:@18899.4]
  wire [10:0] _T_68047; // @[Modules.scala 78:156:@18900.4]
  wire [10:0] buffer_7_765; // @[Modules.scala 78:156:@18901.4]
  wire [11:0] _T_68049; // @[Modules.scala 78:156:@18903.4]
  wire [10:0] _T_68050; // @[Modules.scala 78:156:@18904.4]
  wire [10:0] buffer_7_766; // @[Modules.scala 78:156:@18905.4]
  wire [11:0] _T_68052; // @[Modules.scala 78:156:@18907.4]
  wire [10:0] _T_68053; // @[Modules.scala 78:156:@18908.4]
  wire [10:0] buffer_7_767; // @[Modules.scala 78:156:@18909.4]
  wire [11:0] _T_68055; // @[Modules.scala 78:156:@18911.4]
  wire [10:0] _T_68056; // @[Modules.scala 78:156:@18912.4]
  wire [10:0] buffer_7_768; // @[Modules.scala 78:156:@18913.4]
  wire [11:0] _T_68058; // @[Modules.scala 78:156:@18915.4]
  wire [10:0] _T_68059; // @[Modules.scala 78:156:@18916.4]
  wire [10:0] buffer_7_769; // @[Modules.scala 78:156:@18917.4]
  wire [11:0] _T_68061; // @[Modules.scala 78:156:@18919.4]
  wire [10:0] _T_68062; // @[Modules.scala 78:156:@18920.4]
  wire [10:0] buffer_7_770; // @[Modules.scala 78:156:@18921.4]
  wire [11:0] _T_68064; // @[Modules.scala 78:156:@18923.4]
  wire [10:0] _T_68065; // @[Modules.scala 78:156:@18924.4]
  wire [10:0] buffer_7_771; // @[Modules.scala 78:156:@18925.4]
  wire [11:0] _T_68067; // @[Modules.scala 78:156:@18927.4]
  wire [10:0] _T_68068; // @[Modules.scala 78:156:@18928.4]
  wire [10:0] buffer_7_772; // @[Modules.scala 78:156:@18929.4]
  wire [11:0] _T_68070; // @[Modules.scala 78:156:@18931.4]
  wire [10:0] _T_68071; // @[Modules.scala 78:156:@18932.4]
  wire [10:0] buffer_7_773; // @[Modules.scala 78:156:@18933.4]
  wire [11:0] _T_68073; // @[Modules.scala 78:156:@18935.4]
  wire [10:0] _T_68074; // @[Modules.scala 78:156:@18936.4]
  wire [10:0] buffer_7_774; // @[Modules.scala 78:156:@18937.4]
  wire [11:0] _T_68076; // @[Modules.scala 78:156:@18939.4]
  wire [10:0] _T_68077; // @[Modules.scala 78:156:@18940.4]
  wire [10:0] buffer_7_775; // @[Modules.scala 78:156:@18941.4]
  wire [11:0] _T_68079; // @[Modules.scala 78:156:@18943.4]
  wire [10:0] _T_68080; // @[Modules.scala 78:156:@18944.4]
  wire [10:0] buffer_7_776; // @[Modules.scala 78:156:@18945.4]
  wire [11:0] _T_68082; // @[Modules.scala 78:156:@18947.4]
  wire [10:0] _T_68083; // @[Modules.scala 78:156:@18948.4]
  wire [10:0] buffer_7_777; // @[Modules.scala 78:156:@18949.4]
  wire [11:0] _T_68085; // @[Modules.scala 78:156:@18951.4]
  wire [10:0] _T_68086; // @[Modules.scala 78:156:@18952.4]
  wire [10:0] buffer_7_778; // @[Modules.scala 78:156:@18953.4]
  wire [11:0] _T_68088; // @[Modules.scala 78:156:@18955.4]
  wire [10:0] _T_68089; // @[Modules.scala 78:156:@18956.4]
  wire [10:0] buffer_7_779; // @[Modules.scala 78:156:@18957.4]
  wire [11:0] _T_68091; // @[Modules.scala 78:156:@18959.4]
  wire [10:0] _T_68092; // @[Modules.scala 78:156:@18960.4]
  wire [10:0] buffer_7_780; // @[Modules.scala 78:156:@18961.4]
  wire [11:0] _T_68094; // @[Modules.scala 78:156:@18963.4]
  wire [10:0] _T_68095; // @[Modules.scala 78:156:@18964.4]
  wire [10:0] buffer_7_781; // @[Modules.scala 78:156:@18965.4]
  wire [11:0] _T_68097; // @[Modules.scala 78:156:@18967.4]
  wire [10:0] _T_68098; // @[Modules.scala 78:156:@18968.4]
  wire [10:0] buffer_7_782; // @[Modules.scala 78:156:@18969.4]
  wire [11:0] _T_68100; // @[Modules.scala 78:156:@18971.4]
  wire [10:0] _T_68101; // @[Modules.scala 78:156:@18972.4]
  wire [10:0] buffer_7_783; // @[Modules.scala 78:156:@18973.4]
  wire [5:0] _T_68334; // @[Modules.scala 37:46:@19298.4]
  wire [4:0] _T_68335; // @[Modules.scala 37:46:@19299.4]
  wire [4:0] _T_68336; // @[Modules.scala 37:46:@19300.4]
  wire [5:0] _T_68355; // @[Modules.scala 37:46:@19329.4]
  wire [4:0] _T_68356; // @[Modules.scala 37:46:@19330.4]
  wire [4:0] _T_68357; // @[Modules.scala 37:46:@19331.4]
  wire [11:0] _T_68626; // @[Modules.scala 65:57:@19724.4]
  wire [10:0] _T_68627; // @[Modules.scala 65:57:@19725.4]
  wire [10:0] buffer_8_394; // @[Modules.scala 65:57:@19726.4]
  wire [11:0] _T_68635; // @[Modules.scala 65:57:@19736.4]
  wire [10:0] _T_68636; // @[Modules.scala 65:57:@19737.4]
  wire [10:0] buffer_8_397; // @[Modules.scala 65:57:@19738.4]
  wire [11:0] _T_68641; // @[Modules.scala 65:57:@19744.4]
  wire [10:0] _T_68642; // @[Modules.scala 65:57:@19745.4]
  wire [10:0] buffer_8_399; // @[Modules.scala 65:57:@19746.4]
  wire [11:0] _T_68686; // @[Modules.scala 65:57:@19804.4]
  wire [10:0] _T_68687; // @[Modules.scala 65:57:@19805.4]
  wire [10:0] buffer_8_414; // @[Modules.scala 65:57:@19806.4]
  wire [10:0] buffer_8_55; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68701; // @[Modules.scala 65:57:@19824.4]
  wire [10:0] _T_68702; // @[Modules.scala 65:57:@19825.4]
  wire [10:0] buffer_8_419; // @[Modules.scala 65:57:@19826.4]
  wire [11:0] _T_68704; // @[Modules.scala 65:57:@19828.4]
  wire [10:0] _T_68705; // @[Modules.scala 65:57:@19829.4]
  wire [10:0] buffer_8_420; // @[Modules.scala 65:57:@19830.4]
  wire [10:0] buffer_8_60; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_8_61; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68710; // @[Modules.scala 65:57:@19836.4]
  wire [10:0] _T_68711; // @[Modules.scala 65:57:@19837.4]
  wire [10:0] buffer_8_422; // @[Modules.scala 65:57:@19838.4]
  wire [10:0] buffer_8_62; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68713; // @[Modules.scala 65:57:@19840.4]
  wire [10:0] _T_68714; // @[Modules.scala 65:57:@19841.4]
  wire [10:0] buffer_8_423; // @[Modules.scala 65:57:@19842.4]
  wire [11:0] _T_68725; // @[Modules.scala 65:57:@19856.4]
  wire [10:0] _T_68726; // @[Modules.scala 65:57:@19857.4]
  wire [10:0] buffer_8_427; // @[Modules.scala 65:57:@19858.4]
  wire [11:0] _T_68743; // @[Modules.scala 65:57:@19880.4]
  wire [10:0] _T_68744; // @[Modules.scala 65:57:@19881.4]
  wire [10:0] buffer_8_433; // @[Modules.scala 65:57:@19882.4]
  wire [10:0] buffer_8_96; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68764; // @[Modules.scala 65:57:@19908.4]
  wire [10:0] _T_68765; // @[Modules.scala 65:57:@19909.4]
  wire [10:0] buffer_8_440; // @[Modules.scala 65:57:@19910.4]
  wire [11:0] _T_68773; // @[Modules.scala 65:57:@19920.4]
  wire [10:0] _T_68774; // @[Modules.scala 65:57:@19921.4]
  wire [10:0] buffer_8_443; // @[Modules.scala 65:57:@19922.4]
  wire [11:0] _T_68779; // @[Modules.scala 65:57:@19928.4]
  wire [10:0] _T_68780; // @[Modules.scala 65:57:@19929.4]
  wire [10:0] buffer_8_445; // @[Modules.scala 65:57:@19930.4]
  wire [10:0] buffer_8_112; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68788; // @[Modules.scala 65:57:@19940.4]
  wire [10:0] _T_68789; // @[Modules.scala 65:57:@19941.4]
  wire [10:0] buffer_8_448; // @[Modules.scala 65:57:@19942.4]
  wire [10:0] buffer_8_115; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68791; // @[Modules.scala 65:57:@19944.4]
  wire [10:0] _T_68792; // @[Modules.scala 65:57:@19945.4]
  wire [10:0] buffer_8_449; // @[Modules.scala 65:57:@19946.4]
  wire [10:0] buffer_8_118; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68797; // @[Modules.scala 65:57:@19952.4]
  wire [10:0] _T_68798; // @[Modules.scala 65:57:@19953.4]
  wire [10:0] buffer_8_451; // @[Modules.scala 65:57:@19954.4]
  wire [11:0] _T_68800; // @[Modules.scala 65:57:@19956.4]
  wire [10:0] _T_68801; // @[Modules.scala 65:57:@19957.4]
  wire [10:0] buffer_8_452; // @[Modules.scala 65:57:@19958.4]
  wire [11:0] _T_68803; // @[Modules.scala 65:57:@19960.4]
  wire [10:0] _T_68804; // @[Modules.scala 65:57:@19961.4]
  wire [10:0] buffer_8_453; // @[Modules.scala 65:57:@19962.4]
  wire [10:0] buffer_8_127; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68809; // @[Modules.scala 65:57:@19968.4]
  wire [10:0] _T_68810; // @[Modules.scala 65:57:@19969.4]
  wire [10:0] buffer_8_455; // @[Modules.scala 65:57:@19970.4]
  wire [10:0] buffer_8_128; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68812; // @[Modules.scala 65:57:@19972.4]
  wire [10:0] _T_68813; // @[Modules.scala 65:57:@19973.4]
  wire [10:0] buffer_8_456; // @[Modules.scala 65:57:@19974.4]
  wire [11:0] _T_68824; // @[Modules.scala 65:57:@19988.4]
  wire [10:0] _T_68825; // @[Modules.scala 65:57:@19989.4]
  wire [10:0] buffer_8_460; // @[Modules.scala 65:57:@19990.4]
  wire [10:0] buffer_8_141; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68830; // @[Modules.scala 65:57:@19996.4]
  wire [10:0] _T_68831; // @[Modules.scala 65:57:@19997.4]
  wire [10:0] buffer_8_462; // @[Modules.scala 65:57:@19998.4]
  wire [11:0] _T_68851; // @[Modules.scala 65:57:@20024.4]
  wire [10:0] _T_68852; // @[Modules.scala 65:57:@20025.4]
  wire [10:0] buffer_8_469; // @[Modules.scala 65:57:@20026.4]
  wire [11:0] _T_68863; // @[Modules.scala 65:57:@20040.4]
  wire [10:0] _T_68864; // @[Modules.scala 65:57:@20041.4]
  wire [10:0] buffer_8_473; // @[Modules.scala 65:57:@20042.4]
  wire [11:0] _T_68872; // @[Modules.scala 65:57:@20052.4]
  wire [10:0] _T_68873; // @[Modules.scala 65:57:@20053.4]
  wire [10:0] buffer_8_476; // @[Modules.scala 65:57:@20054.4]
  wire [11:0] _T_68884; // @[Modules.scala 65:57:@20068.4]
  wire [10:0] _T_68885; // @[Modules.scala 65:57:@20069.4]
  wire [10:0] buffer_8_480; // @[Modules.scala 65:57:@20070.4]
  wire [10:0] buffer_8_181; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68890; // @[Modules.scala 65:57:@20076.4]
  wire [10:0] _T_68891; // @[Modules.scala 65:57:@20077.4]
  wire [10:0] buffer_8_482; // @[Modules.scala 65:57:@20078.4]
  wire [10:0] buffer_8_189; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68902; // @[Modules.scala 65:57:@20092.4]
  wire [10:0] _T_68903; // @[Modules.scala 65:57:@20093.4]
  wire [10:0] buffer_8_486; // @[Modules.scala 65:57:@20094.4]
  wire [10:0] buffer_8_192; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68908; // @[Modules.scala 65:57:@20100.4]
  wire [10:0] _T_68909; // @[Modules.scala 65:57:@20101.4]
  wire [10:0] buffer_8_488; // @[Modules.scala 65:57:@20102.4]
  wire [10:0] buffer_8_197; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68914; // @[Modules.scala 65:57:@20108.4]
  wire [10:0] _T_68915; // @[Modules.scala 65:57:@20109.4]
  wire [10:0] buffer_8_490; // @[Modules.scala 65:57:@20110.4]
  wire [11:0] _T_68920; // @[Modules.scala 65:57:@20116.4]
  wire [10:0] _T_68921; // @[Modules.scala 65:57:@20117.4]
  wire [10:0] buffer_8_492; // @[Modules.scala 65:57:@20118.4]
  wire [10:0] buffer_8_204; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68926; // @[Modules.scala 65:57:@20124.4]
  wire [10:0] _T_68927; // @[Modules.scala 65:57:@20125.4]
  wire [10:0] buffer_8_494; // @[Modules.scala 65:57:@20126.4]
  wire [11:0] _T_68929; // @[Modules.scala 65:57:@20128.4]
  wire [10:0] _T_68930; // @[Modules.scala 65:57:@20129.4]
  wire [10:0] buffer_8_495; // @[Modules.scala 65:57:@20130.4]
  wire [11:0] _T_68950; // @[Modules.scala 65:57:@20156.4]
  wire [10:0] _T_68951; // @[Modules.scala 65:57:@20157.4]
  wire [10:0] buffer_8_502; // @[Modules.scala 65:57:@20158.4]
  wire [11:0] _T_68953; // @[Modules.scala 65:57:@20160.4]
  wire [10:0] _T_68954; // @[Modules.scala 65:57:@20161.4]
  wire [10:0] buffer_8_503; // @[Modules.scala 65:57:@20162.4]
  wire [11:0] _T_68956; // @[Modules.scala 65:57:@20164.4]
  wire [10:0] _T_68957; // @[Modules.scala 65:57:@20165.4]
  wire [10:0] buffer_8_504; // @[Modules.scala 65:57:@20166.4]
  wire [10:0] buffer_8_239; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68977; // @[Modules.scala 65:57:@20192.4]
  wire [10:0] _T_68978; // @[Modules.scala 65:57:@20193.4]
  wire [10:0] buffer_8_511; // @[Modules.scala 65:57:@20194.4]
  wire [11:0] _T_68989; // @[Modules.scala 65:57:@20208.4]
  wire [10:0] _T_68990; // @[Modules.scala 65:57:@20209.4]
  wire [10:0] buffer_8_515; // @[Modules.scala 65:57:@20210.4]
  wire [10:0] buffer_8_248; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_68992; // @[Modules.scala 65:57:@20212.4]
  wire [10:0] _T_68993; // @[Modules.scala 65:57:@20213.4]
  wire [10:0] buffer_8_516; // @[Modules.scala 65:57:@20214.4]
  wire [11:0] _T_68998; // @[Modules.scala 65:57:@20220.4]
  wire [10:0] _T_68999; // @[Modules.scala 65:57:@20221.4]
  wire [10:0] buffer_8_518; // @[Modules.scala 65:57:@20222.4]
  wire [10:0] buffer_8_254; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69001; // @[Modules.scala 65:57:@20224.4]
  wire [10:0] _T_69002; // @[Modules.scala 65:57:@20225.4]
  wire [10:0] buffer_8_519; // @[Modules.scala 65:57:@20226.4]
  wire [11:0] _T_69019; // @[Modules.scala 65:57:@20248.4]
  wire [10:0] _T_69020; // @[Modules.scala 65:57:@20249.4]
  wire [10:0] buffer_8_525; // @[Modules.scala 65:57:@20250.4]
  wire [11:0] _T_69022; // @[Modules.scala 65:57:@20252.4]
  wire [10:0] _T_69023; // @[Modules.scala 65:57:@20253.4]
  wire [10:0] buffer_8_526; // @[Modules.scala 65:57:@20254.4]
  wire [11:0] _T_69028; // @[Modules.scala 65:57:@20260.4]
  wire [10:0] _T_69029; // @[Modules.scala 65:57:@20261.4]
  wire [10:0] buffer_8_528; // @[Modules.scala 65:57:@20262.4]
  wire [11:0] _T_69034; // @[Modules.scala 65:57:@20268.4]
  wire [10:0] _T_69035; // @[Modules.scala 65:57:@20269.4]
  wire [10:0] buffer_8_530; // @[Modules.scala 65:57:@20270.4]
  wire [11:0] _T_69040; // @[Modules.scala 65:57:@20276.4]
  wire [10:0] _T_69041; // @[Modules.scala 65:57:@20277.4]
  wire [10:0] buffer_8_532; // @[Modules.scala 65:57:@20278.4]
  wire [11:0] _T_69043; // @[Modules.scala 65:57:@20280.4]
  wire [10:0] _T_69044; // @[Modules.scala 65:57:@20281.4]
  wire [10:0] buffer_8_533; // @[Modules.scala 65:57:@20282.4]
  wire [10:0] buffer_8_284; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69046; // @[Modules.scala 65:57:@20284.4]
  wire [10:0] _T_69047; // @[Modules.scala 65:57:@20285.4]
  wire [10:0] buffer_8_534; // @[Modules.scala 65:57:@20286.4]
  wire [11:0] _T_69058; // @[Modules.scala 65:57:@20300.4]
  wire [10:0] _T_69059; // @[Modules.scala 65:57:@20301.4]
  wire [10:0] buffer_8_538; // @[Modules.scala 65:57:@20302.4]
  wire [10:0] buffer_8_298; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69067; // @[Modules.scala 65:57:@20312.4]
  wire [10:0] _T_69068; // @[Modules.scala 65:57:@20313.4]
  wire [10:0] buffer_8_541; // @[Modules.scala 65:57:@20314.4]
  wire [11:0] _T_69070; // @[Modules.scala 65:57:@20316.4]
  wire [10:0] _T_69071; // @[Modules.scala 65:57:@20317.4]
  wire [10:0] buffer_8_542; // @[Modules.scala 65:57:@20318.4]
  wire [10:0] buffer_8_303; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69073; // @[Modules.scala 65:57:@20320.4]
  wire [10:0] _T_69074; // @[Modules.scala 65:57:@20321.4]
  wire [10:0] buffer_8_543; // @[Modules.scala 65:57:@20322.4]
  wire [10:0] buffer_8_311; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69085; // @[Modules.scala 65:57:@20336.4]
  wire [10:0] _T_69086; // @[Modules.scala 65:57:@20337.4]
  wire [10:0] buffer_8_547; // @[Modules.scala 65:57:@20338.4]
  wire [11:0] _T_69088; // @[Modules.scala 65:57:@20340.4]
  wire [10:0] _T_69089; // @[Modules.scala 65:57:@20341.4]
  wire [10:0] buffer_8_548; // @[Modules.scala 65:57:@20342.4]
  wire [11:0] _T_69091; // @[Modules.scala 65:57:@20344.4]
  wire [10:0] _T_69092; // @[Modules.scala 65:57:@20345.4]
  wire [10:0] buffer_8_549; // @[Modules.scala 65:57:@20346.4]
  wire [11:0] _T_69106; // @[Modules.scala 65:57:@20364.4]
  wire [10:0] _T_69107; // @[Modules.scala 65:57:@20365.4]
  wire [10:0] buffer_8_554; // @[Modules.scala 65:57:@20366.4]
  wire [10:0] buffer_8_327; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69109; // @[Modules.scala 65:57:@20368.4]
  wire [10:0] _T_69110; // @[Modules.scala 65:57:@20369.4]
  wire [10:0] buffer_8_555; // @[Modules.scala 65:57:@20370.4]
  wire [11:0] _T_69115; // @[Modules.scala 65:57:@20376.4]
  wire [10:0] _T_69116; // @[Modules.scala 65:57:@20377.4]
  wire [10:0] buffer_8_557; // @[Modules.scala 65:57:@20378.4]
  wire [11:0] _T_69121; // @[Modules.scala 65:57:@20384.4]
  wire [10:0] _T_69122; // @[Modules.scala 65:57:@20385.4]
  wire [10:0] buffer_8_559; // @[Modules.scala 65:57:@20386.4]
  wire [11:0] _T_69127; // @[Modules.scala 65:57:@20392.4]
  wire [10:0] _T_69128; // @[Modules.scala 65:57:@20393.4]
  wire [10:0] buffer_8_561; // @[Modules.scala 65:57:@20394.4]
  wire [11:0] _T_69145; // @[Modules.scala 65:57:@20416.4]
  wire [10:0] _T_69146; // @[Modules.scala 65:57:@20417.4]
  wire [10:0] buffer_8_567; // @[Modules.scala 65:57:@20418.4]
  wire [11:0] _T_69184; // @[Modules.scala 65:57:@20468.4]
  wire [10:0] _T_69185; // @[Modules.scala 65:57:@20469.4]
  wire [10:0] buffer_8_580; // @[Modules.scala 65:57:@20470.4]
  wire [10:0] buffer_8_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69187; // @[Modules.scala 65:57:@20472.4]
  wire [10:0] _T_69188; // @[Modules.scala 65:57:@20473.4]
  wire [10:0] buffer_8_581; // @[Modules.scala 65:57:@20474.4]
  wire [10:0] buffer_8_382; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_69193; // @[Modules.scala 65:57:@20480.4]
  wire [10:0] _T_69194; // @[Modules.scala 65:57:@20481.4]
  wire [10:0] buffer_8_583; // @[Modules.scala 65:57:@20482.4]
  wire [11:0] _T_69202; // @[Modules.scala 65:57:@20492.4]
  wire [10:0] _T_69203; // @[Modules.scala 65:57:@20493.4]
  wire [10:0] buffer_8_586; // @[Modules.scala 65:57:@20494.4]
  wire [11:0] _T_69211; // @[Modules.scala 68:83:@20504.4]
  wire [10:0] _T_69212; // @[Modules.scala 68:83:@20505.4]
  wire [10:0] buffer_8_589; // @[Modules.scala 68:83:@20506.4]
  wire [11:0] _T_69214; // @[Modules.scala 68:83:@20508.4]
  wire [10:0] _T_69215; // @[Modules.scala 68:83:@20509.4]
  wire [10:0] buffer_8_590; // @[Modules.scala 68:83:@20510.4]
  wire [11:0] _T_69217; // @[Modules.scala 68:83:@20512.4]
  wire [10:0] _T_69218; // @[Modules.scala 68:83:@20513.4]
  wire [10:0] buffer_8_591; // @[Modules.scala 68:83:@20514.4]
  wire [11:0] _T_69226; // @[Modules.scala 68:83:@20524.4]
  wire [10:0] _T_69227; // @[Modules.scala 68:83:@20525.4]
  wire [10:0] buffer_8_594; // @[Modules.scala 68:83:@20526.4]
  wire [11:0] _T_69238; // @[Modules.scala 68:83:@20540.4]
  wire [10:0] _T_69239; // @[Modules.scala 68:83:@20541.4]
  wire [10:0] buffer_8_598; // @[Modules.scala 68:83:@20542.4]
  wire [11:0] _T_69241; // @[Modules.scala 68:83:@20544.4]
  wire [10:0] _T_69242; // @[Modules.scala 68:83:@20545.4]
  wire [10:0] buffer_8_599; // @[Modules.scala 68:83:@20546.4]
  wire [11:0] _T_69247; // @[Modules.scala 68:83:@20552.4]
  wire [10:0] _T_69248; // @[Modules.scala 68:83:@20553.4]
  wire [10:0] buffer_8_601; // @[Modules.scala 68:83:@20554.4]
  wire [11:0] _T_69250; // @[Modules.scala 68:83:@20556.4]
  wire [10:0] _T_69251; // @[Modules.scala 68:83:@20557.4]
  wire [10:0] buffer_8_602; // @[Modules.scala 68:83:@20558.4]
  wire [11:0] _T_69253; // @[Modules.scala 68:83:@20560.4]
  wire [10:0] _T_69254; // @[Modules.scala 68:83:@20561.4]
  wire [10:0] buffer_8_603; // @[Modules.scala 68:83:@20562.4]
  wire [11:0] _T_69259; // @[Modules.scala 68:83:@20568.4]
  wire [10:0] _T_69260; // @[Modules.scala 68:83:@20569.4]
  wire [10:0] buffer_8_605; // @[Modules.scala 68:83:@20570.4]
  wire [11:0] _T_69268; // @[Modules.scala 68:83:@20580.4]
  wire [10:0] _T_69269; // @[Modules.scala 68:83:@20581.4]
  wire [10:0] buffer_8_608; // @[Modules.scala 68:83:@20582.4]
  wire [11:0] _T_69274; // @[Modules.scala 68:83:@20588.4]
  wire [10:0] _T_69275; // @[Modules.scala 68:83:@20589.4]
  wire [10:0] buffer_8_610; // @[Modules.scala 68:83:@20590.4]
  wire [11:0] _T_69277; // @[Modules.scala 68:83:@20592.4]
  wire [10:0] _T_69278; // @[Modules.scala 68:83:@20593.4]
  wire [10:0] buffer_8_611; // @[Modules.scala 68:83:@20594.4]
  wire [11:0] _T_69280; // @[Modules.scala 68:83:@20596.4]
  wire [10:0] _T_69281; // @[Modules.scala 68:83:@20597.4]
  wire [10:0] buffer_8_612; // @[Modules.scala 68:83:@20598.4]
  wire [11:0] _T_69283; // @[Modules.scala 68:83:@20600.4]
  wire [10:0] _T_69284; // @[Modules.scala 68:83:@20601.4]
  wire [10:0] buffer_8_613; // @[Modules.scala 68:83:@20602.4]
  wire [11:0] _T_69286; // @[Modules.scala 68:83:@20604.4]
  wire [10:0] _T_69287; // @[Modules.scala 68:83:@20605.4]
  wire [10:0] buffer_8_614; // @[Modules.scala 68:83:@20606.4]
  wire [11:0] _T_69289; // @[Modules.scala 68:83:@20608.4]
  wire [10:0] _T_69290; // @[Modules.scala 68:83:@20609.4]
  wire [10:0] buffer_8_615; // @[Modules.scala 68:83:@20610.4]
  wire [11:0] _T_69292; // @[Modules.scala 68:83:@20612.4]
  wire [10:0] _T_69293; // @[Modules.scala 68:83:@20613.4]
  wire [10:0] buffer_8_616; // @[Modules.scala 68:83:@20614.4]
  wire [11:0] _T_69295; // @[Modules.scala 68:83:@20616.4]
  wire [10:0] _T_69296; // @[Modules.scala 68:83:@20617.4]
  wire [10:0] buffer_8_617; // @[Modules.scala 68:83:@20618.4]
  wire [11:0] _T_69298; // @[Modules.scala 68:83:@20620.4]
  wire [10:0] _T_69299; // @[Modules.scala 68:83:@20621.4]
  wire [10:0] buffer_8_618; // @[Modules.scala 68:83:@20622.4]
  wire [11:0] _T_69301; // @[Modules.scala 68:83:@20624.4]
  wire [10:0] _T_69302; // @[Modules.scala 68:83:@20625.4]
  wire [10:0] buffer_8_619; // @[Modules.scala 68:83:@20626.4]
  wire [11:0] _T_69304; // @[Modules.scala 68:83:@20628.4]
  wire [10:0] _T_69305; // @[Modules.scala 68:83:@20629.4]
  wire [10:0] buffer_8_620; // @[Modules.scala 68:83:@20630.4]
  wire [11:0] _T_69307; // @[Modules.scala 68:83:@20632.4]
  wire [10:0] _T_69308; // @[Modules.scala 68:83:@20633.4]
  wire [10:0] buffer_8_621; // @[Modules.scala 68:83:@20634.4]
  wire [11:0] _T_69310; // @[Modules.scala 68:83:@20636.4]
  wire [10:0] _T_69311; // @[Modules.scala 68:83:@20637.4]
  wire [10:0] buffer_8_622; // @[Modules.scala 68:83:@20638.4]
  wire [11:0] _T_69313; // @[Modules.scala 68:83:@20640.4]
  wire [10:0] _T_69314; // @[Modules.scala 68:83:@20641.4]
  wire [10:0] buffer_8_623; // @[Modules.scala 68:83:@20642.4]
  wire [11:0] _T_69319; // @[Modules.scala 68:83:@20648.4]
  wire [10:0] _T_69320; // @[Modules.scala 68:83:@20649.4]
  wire [10:0] buffer_8_625; // @[Modules.scala 68:83:@20650.4]
  wire [11:0] _T_69322; // @[Modules.scala 68:83:@20652.4]
  wire [10:0] _T_69323; // @[Modules.scala 68:83:@20653.4]
  wire [10:0] buffer_8_626; // @[Modules.scala 68:83:@20654.4]
  wire [11:0] _T_69328; // @[Modules.scala 68:83:@20660.4]
  wire [10:0] _T_69329; // @[Modules.scala 68:83:@20661.4]
  wire [10:0] buffer_8_628; // @[Modules.scala 68:83:@20662.4]
  wire [11:0] _T_69331; // @[Modules.scala 68:83:@20664.4]
  wire [10:0] _T_69332; // @[Modules.scala 68:83:@20665.4]
  wire [10:0] buffer_8_629; // @[Modules.scala 68:83:@20666.4]
  wire [11:0] _T_69334; // @[Modules.scala 68:83:@20668.4]
  wire [10:0] _T_69335; // @[Modules.scala 68:83:@20669.4]
  wire [10:0] buffer_8_630; // @[Modules.scala 68:83:@20670.4]
  wire [11:0] _T_69340; // @[Modules.scala 68:83:@20676.4]
  wire [10:0] _T_69341; // @[Modules.scala 68:83:@20677.4]
  wire [10:0] buffer_8_632; // @[Modules.scala 68:83:@20678.4]
  wire [11:0] _T_69343; // @[Modules.scala 68:83:@20680.4]
  wire [10:0] _T_69344; // @[Modules.scala 68:83:@20681.4]
  wire [10:0] buffer_8_633; // @[Modules.scala 68:83:@20682.4]
  wire [11:0] _T_69346; // @[Modules.scala 68:83:@20684.4]
  wire [10:0] _T_69347; // @[Modules.scala 68:83:@20685.4]
  wire [10:0] buffer_8_634; // @[Modules.scala 68:83:@20686.4]
  wire [11:0] _T_69349; // @[Modules.scala 68:83:@20688.4]
  wire [10:0] _T_69350; // @[Modules.scala 68:83:@20689.4]
  wire [10:0] buffer_8_635; // @[Modules.scala 68:83:@20690.4]
  wire [11:0] _T_69352; // @[Modules.scala 68:83:@20692.4]
  wire [10:0] _T_69353; // @[Modules.scala 68:83:@20693.4]
  wire [10:0] buffer_8_636; // @[Modules.scala 68:83:@20694.4]
  wire [11:0] _T_69355; // @[Modules.scala 68:83:@20696.4]
  wire [10:0] _T_69356; // @[Modules.scala 68:83:@20697.4]
  wire [10:0] buffer_8_637; // @[Modules.scala 68:83:@20698.4]
  wire [11:0] _T_69358; // @[Modules.scala 68:83:@20700.4]
  wire [10:0] _T_69359; // @[Modules.scala 68:83:@20701.4]
  wire [10:0] buffer_8_638; // @[Modules.scala 68:83:@20702.4]
  wire [11:0] _T_69361; // @[Modules.scala 68:83:@20704.4]
  wire [10:0] _T_69362; // @[Modules.scala 68:83:@20705.4]
  wire [10:0] buffer_8_639; // @[Modules.scala 68:83:@20706.4]
  wire [11:0] _T_69367; // @[Modules.scala 68:83:@20712.4]
  wire [10:0] _T_69368; // @[Modules.scala 68:83:@20713.4]
  wire [10:0] buffer_8_641; // @[Modules.scala 68:83:@20714.4]
  wire [11:0] _T_69370; // @[Modules.scala 68:83:@20716.4]
  wire [10:0] _T_69371; // @[Modules.scala 68:83:@20717.4]
  wire [10:0] buffer_8_642; // @[Modules.scala 68:83:@20718.4]
  wire [11:0] _T_69373; // @[Modules.scala 68:83:@20720.4]
  wire [10:0] _T_69374; // @[Modules.scala 68:83:@20721.4]
  wire [10:0] buffer_8_643; // @[Modules.scala 68:83:@20722.4]
  wire [11:0] _T_69376; // @[Modules.scala 68:83:@20724.4]
  wire [10:0] _T_69377; // @[Modules.scala 68:83:@20725.4]
  wire [10:0] buffer_8_644; // @[Modules.scala 68:83:@20726.4]
  wire [11:0] _T_69382; // @[Modules.scala 68:83:@20732.4]
  wire [10:0] _T_69383; // @[Modules.scala 68:83:@20733.4]
  wire [10:0] buffer_8_646; // @[Modules.scala 68:83:@20734.4]
  wire [11:0] _T_69385; // @[Modules.scala 68:83:@20736.4]
  wire [10:0] _T_69386; // @[Modules.scala 68:83:@20737.4]
  wire [10:0] buffer_8_647; // @[Modules.scala 68:83:@20738.4]
  wire [11:0] _T_69388; // @[Modules.scala 68:83:@20740.4]
  wire [10:0] _T_69389; // @[Modules.scala 68:83:@20741.4]
  wire [10:0] buffer_8_648; // @[Modules.scala 68:83:@20742.4]
  wire [11:0] _T_69391; // @[Modules.scala 68:83:@20744.4]
  wire [10:0] _T_69392; // @[Modules.scala 68:83:@20745.4]
  wire [10:0] buffer_8_649; // @[Modules.scala 68:83:@20746.4]
  wire [11:0] _T_69394; // @[Modules.scala 68:83:@20748.4]
  wire [10:0] _T_69395; // @[Modules.scala 68:83:@20749.4]
  wire [10:0] buffer_8_650; // @[Modules.scala 68:83:@20750.4]
  wire [11:0] _T_69397; // @[Modules.scala 68:83:@20752.4]
  wire [10:0] _T_69398; // @[Modules.scala 68:83:@20753.4]
  wire [10:0] buffer_8_651; // @[Modules.scala 68:83:@20754.4]
  wire [11:0] _T_69400; // @[Modules.scala 68:83:@20756.4]
  wire [10:0] _T_69401; // @[Modules.scala 68:83:@20757.4]
  wire [10:0] buffer_8_652; // @[Modules.scala 68:83:@20758.4]
  wire [11:0] _T_69403; // @[Modules.scala 68:83:@20760.4]
  wire [10:0] _T_69404; // @[Modules.scala 68:83:@20761.4]
  wire [10:0] buffer_8_653; // @[Modules.scala 68:83:@20762.4]
  wire [11:0] _T_69406; // @[Modules.scala 68:83:@20764.4]
  wire [10:0] _T_69407; // @[Modules.scala 68:83:@20765.4]
  wire [10:0] buffer_8_654; // @[Modules.scala 68:83:@20766.4]
  wire [11:0] _T_69409; // @[Modules.scala 68:83:@20768.4]
  wire [10:0] _T_69410; // @[Modules.scala 68:83:@20769.4]
  wire [10:0] buffer_8_655; // @[Modules.scala 68:83:@20770.4]
  wire [11:0] _T_69412; // @[Modules.scala 68:83:@20772.4]
  wire [10:0] _T_69413; // @[Modules.scala 68:83:@20773.4]
  wire [10:0] buffer_8_656; // @[Modules.scala 68:83:@20774.4]
  wire [11:0] _T_69415; // @[Modules.scala 68:83:@20776.4]
  wire [10:0] _T_69416; // @[Modules.scala 68:83:@20777.4]
  wire [10:0] buffer_8_657; // @[Modules.scala 68:83:@20778.4]
  wire [11:0] _T_69418; // @[Modules.scala 68:83:@20780.4]
  wire [10:0] _T_69419; // @[Modules.scala 68:83:@20781.4]
  wire [10:0] buffer_8_658; // @[Modules.scala 68:83:@20782.4]
  wire [11:0] _T_69421; // @[Modules.scala 68:83:@20784.4]
  wire [10:0] _T_69422; // @[Modules.scala 68:83:@20785.4]
  wire [10:0] buffer_8_659; // @[Modules.scala 68:83:@20786.4]
  wire [11:0] _T_69424; // @[Modules.scala 68:83:@20788.4]
  wire [10:0] _T_69425; // @[Modules.scala 68:83:@20789.4]
  wire [10:0] buffer_8_660; // @[Modules.scala 68:83:@20790.4]
  wire [11:0] _T_69427; // @[Modules.scala 68:83:@20792.4]
  wire [10:0] _T_69428; // @[Modules.scala 68:83:@20793.4]
  wire [10:0] buffer_8_661; // @[Modules.scala 68:83:@20794.4]
  wire [11:0] _T_69430; // @[Modules.scala 68:83:@20796.4]
  wire [10:0] _T_69431; // @[Modules.scala 68:83:@20797.4]
  wire [10:0] buffer_8_662; // @[Modules.scala 68:83:@20798.4]
  wire [11:0] _T_69433; // @[Modules.scala 68:83:@20800.4]
  wire [10:0] _T_69434; // @[Modules.scala 68:83:@20801.4]
  wire [10:0] buffer_8_663; // @[Modules.scala 68:83:@20802.4]
  wire [11:0] _T_69439; // @[Modules.scala 68:83:@20808.4]
  wire [10:0] _T_69440; // @[Modules.scala 68:83:@20809.4]
  wire [10:0] buffer_8_665; // @[Modules.scala 68:83:@20810.4]
  wire [11:0] _T_69442; // @[Modules.scala 68:83:@20812.4]
  wire [10:0] _T_69443; // @[Modules.scala 68:83:@20813.4]
  wire [10:0] buffer_8_666; // @[Modules.scala 68:83:@20814.4]
  wire [11:0] _T_69451; // @[Modules.scala 68:83:@20824.4]
  wire [10:0] _T_69452; // @[Modules.scala 68:83:@20825.4]
  wire [10:0] buffer_8_669; // @[Modules.scala 68:83:@20826.4]
  wire [11:0] _T_69454; // @[Modules.scala 68:83:@20828.4]
  wire [10:0] _T_69455; // @[Modules.scala 68:83:@20829.4]
  wire [10:0] buffer_8_670; // @[Modules.scala 68:83:@20830.4]
  wire [11:0] _T_69457; // @[Modules.scala 68:83:@20832.4]
  wire [10:0] _T_69458; // @[Modules.scala 68:83:@20833.4]
  wire [10:0] buffer_8_671; // @[Modules.scala 68:83:@20834.4]
  wire [11:0] _T_69460; // @[Modules.scala 68:83:@20836.4]
  wire [10:0] _T_69461; // @[Modules.scala 68:83:@20837.4]
  wire [10:0] buffer_8_672; // @[Modules.scala 68:83:@20838.4]
  wire [11:0] _T_69469; // @[Modules.scala 68:83:@20848.4]
  wire [10:0] _T_69470; // @[Modules.scala 68:83:@20849.4]
  wire [10:0] buffer_8_675; // @[Modules.scala 68:83:@20850.4]
  wire [11:0] _T_69490; // @[Modules.scala 68:83:@20876.4]
  wire [10:0] _T_69491; // @[Modules.scala 68:83:@20877.4]
  wire [10:0] buffer_8_682; // @[Modules.scala 68:83:@20878.4]
  wire [11:0] _T_69493; // @[Modules.scala 68:83:@20880.4]
  wire [10:0] _T_69494; // @[Modules.scala 68:83:@20881.4]
  wire [10:0] buffer_8_683; // @[Modules.scala 68:83:@20882.4]
  wire [11:0] _T_69499; // @[Modules.scala 68:83:@20888.4]
  wire [10:0] _T_69500; // @[Modules.scala 68:83:@20889.4]
  wire [10:0] buffer_8_685; // @[Modules.scala 68:83:@20890.4]
  wire [11:0] _T_69502; // @[Modules.scala 71:109:@20892.4]
  wire [10:0] _T_69503; // @[Modules.scala 71:109:@20893.4]
  wire [10:0] buffer_8_686; // @[Modules.scala 71:109:@20894.4]
  wire [11:0] _T_69505; // @[Modules.scala 71:109:@20896.4]
  wire [10:0] _T_69506; // @[Modules.scala 71:109:@20897.4]
  wire [10:0] buffer_8_687; // @[Modules.scala 71:109:@20898.4]
  wire [11:0] _T_69511; // @[Modules.scala 71:109:@20904.4]
  wire [10:0] _T_69512; // @[Modules.scala 71:109:@20905.4]
  wire [10:0] buffer_8_689; // @[Modules.scala 71:109:@20906.4]
  wire [11:0] _T_69517; // @[Modules.scala 71:109:@20912.4]
  wire [10:0] _T_69518; // @[Modules.scala 71:109:@20913.4]
  wire [10:0] buffer_8_691; // @[Modules.scala 71:109:@20914.4]
  wire [11:0] _T_69520; // @[Modules.scala 71:109:@20916.4]
  wire [10:0] _T_69521; // @[Modules.scala 71:109:@20917.4]
  wire [10:0] buffer_8_692; // @[Modules.scala 71:109:@20918.4]
  wire [11:0] _T_69523; // @[Modules.scala 71:109:@20920.4]
  wire [10:0] _T_69524; // @[Modules.scala 71:109:@20921.4]
  wire [10:0] buffer_8_693; // @[Modules.scala 71:109:@20922.4]
  wire [11:0] _T_69526; // @[Modules.scala 71:109:@20924.4]
  wire [10:0] _T_69527; // @[Modules.scala 71:109:@20925.4]
  wire [10:0] buffer_8_694; // @[Modules.scala 71:109:@20926.4]
  wire [11:0] _T_69532; // @[Modules.scala 71:109:@20932.4]
  wire [10:0] _T_69533; // @[Modules.scala 71:109:@20933.4]
  wire [10:0] buffer_8_696; // @[Modules.scala 71:109:@20934.4]
  wire [11:0] _T_69535; // @[Modules.scala 71:109:@20936.4]
  wire [10:0] _T_69536; // @[Modules.scala 71:109:@20937.4]
  wire [10:0] buffer_8_697; // @[Modules.scala 71:109:@20938.4]
  wire [11:0] _T_69538; // @[Modules.scala 71:109:@20940.4]
  wire [10:0] _T_69539; // @[Modules.scala 71:109:@20941.4]
  wire [10:0] buffer_8_698; // @[Modules.scala 71:109:@20942.4]
  wire [11:0] _T_69541; // @[Modules.scala 71:109:@20944.4]
  wire [10:0] _T_69542; // @[Modules.scala 71:109:@20945.4]
  wire [10:0] buffer_8_699; // @[Modules.scala 71:109:@20946.4]
  wire [11:0] _T_69544; // @[Modules.scala 71:109:@20948.4]
  wire [10:0] _T_69545; // @[Modules.scala 71:109:@20949.4]
  wire [10:0] buffer_8_700; // @[Modules.scala 71:109:@20950.4]
  wire [11:0] _T_69547; // @[Modules.scala 71:109:@20952.4]
  wire [10:0] _T_69548; // @[Modules.scala 71:109:@20953.4]
  wire [10:0] buffer_8_701; // @[Modules.scala 71:109:@20954.4]
  wire [11:0] _T_69550; // @[Modules.scala 71:109:@20956.4]
  wire [10:0] _T_69551; // @[Modules.scala 71:109:@20957.4]
  wire [10:0] buffer_8_702; // @[Modules.scala 71:109:@20958.4]
  wire [11:0] _T_69553; // @[Modules.scala 71:109:@20960.4]
  wire [10:0] _T_69554; // @[Modules.scala 71:109:@20961.4]
  wire [10:0] buffer_8_703; // @[Modules.scala 71:109:@20962.4]
  wire [11:0] _T_69556; // @[Modules.scala 71:109:@20964.4]
  wire [10:0] _T_69557; // @[Modules.scala 71:109:@20965.4]
  wire [10:0] buffer_8_704; // @[Modules.scala 71:109:@20966.4]
  wire [11:0] _T_69559; // @[Modules.scala 71:109:@20968.4]
  wire [10:0] _T_69560; // @[Modules.scala 71:109:@20969.4]
  wire [10:0] buffer_8_705; // @[Modules.scala 71:109:@20970.4]
  wire [11:0] _T_69562; // @[Modules.scala 71:109:@20972.4]
  wire [10:0] _T_69563; // @[Modules.scala 71:109:@20973.4]
  wire [10:0] buffer_8_706; // @[Modules.scala 71:109:@20974.4]
  wire [11:0] _T_69565; // @[Modules.scala 71:109:@20976.4]
  wire [10:0] _T_69566; // @[Modules.scala 71:109:@20977.4]
  wire [10:0] buffer_8_707; // @[Modules.scala 71:109:@20978.4]
  wire [11:0] _T_69568; // @[Modules.scala 71:109:@20980.4]
  wire [10:0] _T_69569; // @[Modules.scala 71:109:@20981.4]
  wire [10:0] buffer_8_708; // @[Modules.scala 71:109:@20982.4]
  wire [11:0] _T_69571; // @[Modules.scala 71:109:@20984.4]
  wire [10:0] _T_69572; // @[Modules.scala 71:109:@20985.4]
  wire [10:0] buffer_8_709; // @[Modules.scala 71:109:@20986.4]
  wire [11:0] _T_69574; // @[Modules.scala 71:109:@20988.4]
  wire [10:0] _T_69575; // @[Modules.scala 71:109:@20989.4]
  wire [10:0] buffer_8_710; // @[Modules.scala 71:109:@20990.4]
  wire [11:0] _T_69577; // @[Modules.scala 71:109:@20992.4]
  wire [10:0] _T_69578; // @[Modules.scala 71:109:@20993.4]
  wire [10:0] buffer_8_711; // @[Modules.scala 71:109:@20994.4]
  wire [11:0] _T_69580; // @[Modules.scala 71:109:@20996.4]
  wire [10:0] _T_69581; // @[Modules.scala 71:109:@20997.4]
  wire [10:0] buffer_8_712; // @[Modules.scala 71:109:@20998.4]
  wire [11:0] _T_69583; // @[Modules.scala 71:109:@21000.4]
  wire [10:0] _T_69584; // @[Modules.scala 71:109:@21001.4]
  wire [10:0] buffer_8_713; // @[Modules.scala 71:109:@21002.4]
  wire [11:0] _T_69586; // @[Modules.scala 71:109:@21004.4]
  wire [10:0] _T_69587; // @[Modules.scala 71:109:@21005.4]
  wire [10:0] buffer_8_714; // @[Modules.scala 71:109:@21006.4]
  wire [11:0] _T_69589; // @[Modules.scala 71:109:@21008.4]
  wire [10:0] _T_69590; // @[Modules.scala 71:109:@21009.4]
  wire [10:0] buffer_8_715; // @[Modules.scala 71:109:@21010.4]
  wire [11:0] _T_69592; // @[Modules.scala 71:109:@21012.4]
  wire [10:0] _T_69593; // @[Modules.scala 71:109:@21013.4]
  wire [10:0] buffer_8_716; // @[Modules.scala 71:109:@21014.4]
  wire [11:0] _T_69595; // @[Modules.scala 71:109:@21016.4]
  wire [10:0] _T_69596; // @[Modules.scala 71:109:@21017.4]
  wire [10:0] buffer_8_717; // @[Modules.scala 71:109:@21018.4]
  wire [11:0] _T_69598; // @[Modules.scala 71:109:@21020.4]
  wire [10:0] _T_69599; // @[Modules.scala 71:109:@21021.4]
  wire [10:0] buffer_8_718; // @[Modules.scala 71:109:@21022.4]
  wire [11:0] _T_69601; // @[Modules.scala 71:109:@21024.4]
  wire [10:0] _T_69602; // @[Modules.scala 71:109:@21025.4]
  wire [10:0] buffer_8_719; // @[Modules.scala 71:109:@21026.4]
  wire [11:0] _T_69604; // @[Modules.scala 71:109:@21028.4]
  wire [10:0] _T_69605; // @[Modules.scala 71:109:@21029.4]
  wire [10:0] buffer_8_720; // @[Modules.scala 71:109:@21030.4]
  wire [11:0] _T_69607; // @[Modules.scala 71:109:@21032.4]
  wire [10:0] _T_69608; // @[Modules.scala 71:109:@21033.4]
  wire [10:0] buffer_8_721; // @[Modules.scala 71:109:@21034.4]
  wire [11:0] _T_69610; // @[Modules.scala 71:109:@21036.4]
  wire [10:0] _T_69611; // @[Modules.scala 71:109:@21037.4]
  wire [10:0] buffer_8_722; // @[Modules.scala 71:109:@21038.4]
  wire [11:0] _T_69613; // @[Modules.scala 71:109:@21040.4]
  wire [10:0] _T_69614; // @[Modules.scala 71:109:@21041.4]
  wire [10:0] buffer_8_723; // @[Modules.scala 71:109:@21042.4]
  wire [11:0] _T_69616; // @[Modules.scala 71:109:@21044.4]
  wire [10:0] _T_69617; // @[Modules.scala 71:109:@21045.4]
  wire [10:0] buffer_8_724; // @[Modules.scala 71:109:@21046.4]
  wire [11:0] _T_69619; // @[Modules.scala 71:109:@21048.4]
  wire [10:0] _T_69620; // @[Modules.scala 71:109:@21049.4]
  wire [10:0] buffer_8_725; // @[Modules.scala 71:109:@21050.4]
  wire [11:0] _T_69622; // @[Modules.scala 71:109:@21052.4]
  wire [10:0] _T_69623; // @[Modules.scala 71:109:@21053.4]
  wire [10:0] buffer_8_726; // @[Modules.scala 71:109:@21054.4]
  wire [11:0] _T_69625; // @[Modules.scala 71:109:@21056.4]
  wire [10:0] _T_69626; // @[Modules.scala 71:109:@21057.4]
  wire [10:0] buffer_8_727; // @[Modules.scala 71:109:@21058.4]
  wire [11:0] _T_69628; // @[Modules.scala 71:109:@21060.4]
  wire [10:0] _T_69629; // @[Modules.scala 71:109:@21061.4]
  wire [10:0] buffer_8_728; // @[Modules.scala 71:109:@21062.4]
  wire [11:0] _T_69631; // @[Modules.scala 71:109:@21064.4]
  wire [10:0] _T_69632; // @[Modules.scala 71:109:@21065.4]
  wire [10:0] buffer_8_729; // @[Modules.scala 71:109:@21066.4]
  wire [11:0] _T_69637; // @[Modules.scala 71:109:@21072.4]
  wire [10:0] _T_69638; // @[Modules.scala 71:109:@21073.4]
  wire [10:0] buffer_8_731; // @[Modules.scala 71:109:@21074.4]
  wire [11:0] _T_69643; // @[Modules.scala 71:109:@21080.4]
  wire [10:0] _T_69644; // @[Modules.scala 71:109:@21081.4]
  wire [10:0] buffer_8_733; // @[Modules.scala 71:109:@21082.4]
  wire [11:0] _T_69646; // @[Modules.scala 71:109:@21084.4]
  wire [10:0] _T_69647; // @[Modules.scala 71:109:@21085.4]
  wire [10:0] buffer_8_734; // @[Modules.scala 71:109:@21086.4]
  wire [11:0] _T_69649; // @[Modules.scala 78:156:@21089.4]
  wire [10:0] _T_69650; // @[Modules.scala 78:156:@21090.4]
  wire [10:0] buffer_8_736; // @[Modules.scala 78:156:@21091.4]
  wire [11:0] _T_69652; // @[Modules.scala 78:156:@21093.4]
  wire [10:0] _T_69653; // @[Modules.scala 78:156:@21094.4]
  wire [10:0] buffer_8_737; // @[Modules.scala 78:156:@21095.4]
  wire [11:0] _T_69655; // @[Modules.scala 78:156:@21097.4]
  wire [10:0] _T_69656; // @[Modules.scala 78:156:@21098.4]
  wire [10:0] buffer_8_738; // @[Modules.scala 78:156:@21099.4]
  wire [11:0] _T_69658; // @[Modules.scala 78:156:@21101.4]
  wire [10:0] _T_69659; // @[Modules.scala 78:156:@21102.4]
  wire [10:0] buffer_8_739; // @[Modules.scala 78:156:@21103.4]
  wire [11:0] _T_69661; // @[Modules.scala 78:156:@21105.4]
  wire [10:0] _T_69662; // @[Modules.scala 78:156:@21106.4]
  wire [10:0] buffer_8_740; // @[Modules.scala 78:156:@21107.4]
  wire [11:0] _T_69664; // @[Modules.scala 78:156:@21109.4]
  wire [10:0] _T_69665; // @[Modules.scala 78:156:@21110.4]
  wire [10:0] buffer_8_741; // @[Modules.scala 78:156:@21111.4]
  wire [11:0] _T_69667; // @[Modules.scala 78:156:@21113.4]
  wire [10:0] _T_69668; // @[Modules.scala 78:156:@21114.4]
  wire [10:0] buffer_8_742; // @[Modules.scala 78:156:@21115.4]
  wire [11:0] _T_69670; // @[Modules.scala 78:156:@21117.4]
  wire [10:0] _T_69671; // @[Modules.scala 78:156:@21118.4]
  wire [10:0] buffer_8_743; // @[Modules.scala 78:156:@21119.4]
  wire [11:0] _T_69673; // @[Modules.scala 78:156:@21121.4]
  wire [10:0] _T_69674; // @[Modules.scala 78:156:@21122.4]
  wire [10:0] buffer_8_744; // @[Modules.scala 78:156:@21123.4]
  wire [11:0] _T_69676; // @[Modules.scala 78:156:@21125.4]
  wire [10:0] _T_69677; // @[Modules.scala 78:156:@21126.4]
  wire [10:0] buffer_8_745; // @[Modules.scala 78:156:@21127.4]
  wire [11:0] _T_69679; // @[Modules.scala 78:156:@21129.4]
  wire [10:0] _T_69680; // @[Modules.scala 78:156:@21130.4]
  wire [10:0] buffer_8_746; // @[Modules.scala 78:156:@21131.4]
  wire [11:0] _T_69682; // @[Modules.scala 78:156:@21133.4]
  wire [10:0] _T_69683; // @[Modules.scala 78:156:@21134.4]
  wire [10:0] buffer_8_747; // @[Modules.scala 78:156:@21135.4]
  wire [11:0] _T_69685; // @[Modules.scala 78:156:@21137.4]
  wire [10:0] _T_69686; // @[Modules.scala 78:156:@21138.4]
  wire [10:0] buffer_8_748; // @[Modules.scala 78:156:@21139.4]
  wire [11:0] _T_69688; // @[Modules.scala 78:156:@21141.4]
  wire [10:0] _T_69689; // @[Modules.scala 78:156:@21142.4]
  wire [10:0] buffer_8_749; // @[Modules.scala 78:156:@21143.4]
  wire [11:0] _T_69691; // @[Modules.scala 78:156:@21145.4]
  wire [10:0] _T_69692; // @[Modules.scala 78:156:@21146.4]
  wire [10:0] buffer_8_750; // @[Modules.scala 78:156:@21147.4]
  wire [11:0] _T_69694; // @[Modules.scala 78:156:@21149.4]
  wire [10:0] _T_69695; // @[Modules.scala 78:156:@21150.4]
  wire [10:0] buffer_8_751; // @[Modules.scala 78:156:@21151.4]
  wire [11:0] _T_69697; // @[Modules.scala 78:156:@21153.4]
  wire [10:0] _T_69698; // @[Modules.scala 78:156:@21154.4]
  wire [10:0] buffer_8_752; // @[Modules.scala 78:156:@21155.4]
  wire [11:0] _T_69700; // @[Modules.scala 78:156:@21157.4]
  wire [10:0] _T_69701; // @[Modules.scala 78:156:@21158.4]
  wire [10:0] buffer_8_753; // @[Modules.scala 78:156:@21159.4]
  wire [11:0] _T_69703; // @[Modules.scala 78:156:@21161.4]
  wire [10:0] _T_69704; // @[Modules.scala 78:156:@21162.4]
  wire [10:0] buffer_8_754; // @[Modules.scala 78:156:@21163.4]
  wire [11:0] _T_69706; // @[Modules.scala 78:156:@21165.4]
  wire [10:0] _T_69707; // @[Modules.scala 78:156:@21166.4]
  wire [10:0] buffer_8_755; // @[Modules.scala 78:156:@21167.4]
  wire [11:0] _T_69709; // @[Modules.scala 78:156:@21169.4]
  wire [10:0] _T_69710; // @[Modules.scala 78:156:@21170.4]
  wire [10:0] buffer_8_756; // @[Modules.scala 78:156:@21171.4]
  wire [11:0] _T_69712; // @[Modules.scala 78:156:@21173.4]
  wire [10:0] _T_69713; // @[Modules.scala 78:156:@21174.4]
  wire [10:0] buffer_8_757; // @[Modules.scala 78:156:@21175.4]
  wire [11:0] _T_69715; // @[Modules.scala 78:156:@21177.4]
  wire [10:0] _T_69716; // @[Modules.scala 78:156:@21178.4]
  wire [10:0] buffer_8_758; // @[Modules.scala 78:156:@21179.4]
  wire [11:0] _T_69718; // @[Modules.scala 78:156:@21181.4]
  wire [10:0] _T_69719; // @[Modules.scala 78:156:@21182.4]
  wire [10:0] buffer_8_759; // @[Modules.scala 78:156:@21183.4]
  wire [11:0] _T_69721; // @[Modules.scala 78:156:@21185.4]
  wire [10:0] _T_69722; // @[Modules.scala 78:156:@21186.4]
  wire [10:0] buffer_8_760; // @[Modules.scala 78:156:@21187.4]
  wire [11:0] _T_69724; // @[Modules.scala 78:156:@21189.4]
  wire [10:0] _T_69725; // @[Modules.scala 78:156:@21190.4]
  wire [10:0] buffer_8_761; // @[Modules.scala 78:156:@21191.4]
  wire [11:0] _T_69727; // @[Modules.scala 78:156:@21193.4]
  wire [10:0] _T_69728; // @[Modules.scala 78:156:@21194.4]
  wire [10:0] buffer_8_762; // @[Modules.scala 78:156:@21195.4]
  wire [11:0] _T_69730; // @[Modules.scala 78:156:@21197.4]
  wire [10:0] _T_69731; // @[Modules.scala 78:156:@21198.4]
  wire [10:0] buffer_8_763; // @[Modules.scala 78:156:@21199.4]
  wire [11:0] _T_69733; // @[Modules.scala 78:156:@21201.4]
  wire [10:0] _T_69734; // @[Modules.scala 78:156:@21202.4]
  wire [10:0] buffer_8_764; // @[Modules.scala 78:156:@21203.4]
  wire [11:0] _T_69736; // @[Modules.scala 78:156:@21205.4]
  wire [10:0] _T_69737; // @[Modules.scala 78:156:@21206.4]
  wire [10:0] buffer_8_765; // @[Modules.scala 78:156:@21207.4]
  wire [11:0] _T_69739; // @[Modules.scala 78:156:@21209.4]
  wire [10:0] _T_69740; // @[Modules.scala 78:156:@21210.4]
  wire [10:0] buffer_8_766; // @[Modules.scala 78:156:@21211.4]
  wire [11:0] _T_69742; // @[Modules.scala 78:156:@21213.4]
  wire [10:0] _T_69743; // @[Modules.scala 78:156:@21214.4]
  wire [10:0] buffer_8_767; // @[Modules.scala 78:156:@21215.4]
  wire [11:0] _T_69745; // @[Modules.scala 78:156:@21217.4]
  wire [10:0] _T_69746; // @[Modules.scala 78:156:@21218.4]
  wire [10:0] buffer_8_768; // @[Modules.scala 78:156:@21219.4]
  wire [11:0] _T_69748; // @[Modules.scala 78:156:@21221.4]
  wire [10:0] _T_69749; // @[Modules.scala 78:156:@21222.4]
  wire [10:0] buffer_8_769; // @[Modules.scala 78:156:@21223.4]
  wire [11:0] _T_69751; // @[Modules.scala 78:156:@21225.4]
  wire [10:0] _T_69752; // @[Modules.scala 78:156:@21226.4]
  wire [10:0] buffer_8_770; // @[Modules.scala 78:156:@21227.4]
  wire [11:0] _T_69754; // @[Modules.scala 78:156:@21229.4]
  wire [10:0] _T_69755; // @[Modules.scala 78:156:@21230.4]
  wire [10:0] buffer_8_771; // @[Modules.scala 78:156:@21231.4]
  wire [11:0] _T_69757; // @[Modules.scala 78:156:@21233.4]
  wire [10:0] _T_69758; // @[Modules.scala 78:156:@21234.4]
  wire [10:0] buffer_8_772; // @[Modules.scala 78:156:@21235.4]
  wire [11:0] _T_69760; // @[Modules.scala 78:156:@21237.4]
  wire [10:0] _T_69761; // @[Modules.scala 78:156:@21238.4]
  wire [10:0] buffer_8_773; // @[Modules.scala 78:156:@21239.4]
  wire [11:0] _T_69763; // @[Modules.scala 78:156:@21241.4]
  wire [10:0] _T_69764; // @[Modules.scala 78:156:@21242.4]
  wire [10:0] buffer_8_774; // @[Modules.scala 78:156:@21243.4]
  wire [11:0] _T_69766; // @[Modules.scala 78:156:@21245.4]
  wire [10:0] _T_69767; // @[Modules.scala 78:156:@21246.4]
  wire [10:0] buffer_8_775; // @[Modules.scala 78:156:@21247.4]
  wire [11:0] _T_69769; // @[Modules.scala 78:156:@21249.4]
  wire [10:0] _T_69770; // @[Modules.scala 78:156:@21250.4]
  wire [10:0] buffer_8_776; // @[Modules.scala 78:156:@21251.4]
  wire [11:0] _T_69772; // @[Modules.scala 78:156:@21253.4]
  wire [10:0] _T_69773; // @[Modules.scala 78:156:@21254.4]
  wire [10:0] buffer_8_777; // @[Modules.scala 78:156:@21255.4]
  wire [11:0] _T_69775; // @[Modules.scala 78:156:@21257.4]
  wire [10:0] _T_69776; // @[Modules.scala 78:156:@21258.4]
  wire [10:0] buffer_8_778; // @[Modules.scala 78:156:@21259.4]
  wire [11:0] _T_69778; // @[Modules.scala 78:156:@21261.4]
  wire [10:0] _T_69779; // @[Modules.scala 78:156:@21262.4]
  wire [10:0] buffer_8_779; // @[Modules.scala 78:156:@21263.4]
  wire [11:0] _T_69781; // @[Modules.scala 78:156:@21265.4]
  wire [10:0] _T_69782; // @[Modules.scala 78:156:@21266.4]
  wire [10:0] buffer_8_780; // @[Modules.scala 78:156:@21267.4]
  wire [11:0] _T_69784; // @[Modules.scala 78:156:@21269.4]
  wire [10:0] _T_69785; // @[Modules.scala 78:156:@21270.4]
  wire [10:0] buffer_8_781; // @[Modules.scala 78:156:@21271.4]
  wire [11:0] _T_69787; // @[Modules.scala 78:156:@21273.4]
  wire [10:0] _T_69788; // @[Modules.scala 78:156:@21274.4]
  wire [10:0] buffer_8_782; // @[Modules.scala 78:156:@21275.4]
  wire [11:0] _T_69790; // @[Modules.scala 78:156:@21277.4]
  wire [10:0] _T_69791; // @[Modules.scala 78:156:@21278.4]
  wire [10:0] buffer_8_783; // @[Modules.scala 78:156:@21279.4]
  wire [5:0] _T_69794; // @[Modules.scala 37:46:@21283.4]
  wire [4:0] _T_69795; // @[Modules.scala 37:46:@21284.4]
  wire [4:0] _T_69796; // @[Modules.scala 37:46:@21285.4]
  wire [5:0] _T_69803; // @[Modules.scala 37:46:@21294.4]
  wire [4:0] _T_69804; // @[Modules.scala 37:46:@21295.4]
  wire [4:0] _T_69805; // @[Modules.scala 37:46:@21296.4]
  wire [10:0] buffer_9_1; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70417; // @[Modules.scala 65:57:@22199.4]
  wire [10:0] _T_70418; // @[Modules.scala 65:57:@22200.4]
  wire [10:0] buffer_9_392; // @[Modules.scala 65:57:@22201.4]
  wire [11:0] _T_70420; // @[Modules.scala 65:57:@22203.4]
  wire [10:0] _T_70421; // @[Modules.scala 65:57:@22204.4]
  wire [10:0] buffer_9_393; // @[Modules.scala 65:57:@22205.4]
  wire [10:0] buffer_9_9; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70429; // @[Modules.scala 65:57:@22215.4]
  wire [10:0] _T_70430; // @[Modules.scala 65:57:@22216.4]
  wire [10:0] buffer_9_396; // @[Modules.scala 65:57:@22217.4]
  wire [11:0] _T_70435; // @[Modules.scala 65:57:@22223.4]
  wire [10:0] _T_70436; // @[Modules.scala 65:57:@22224.4]
  wire [10:0] buffer_9_398; // @[Modules.scala 65:57:@22225.4]
  wire [11:0] _T_70450; // @[Modules.scala 65:57:@22243.4]
  wire [10:0] _T_70451; // @[Modules.scala 65:57:@22244.4]
  wire [10:0] buffer_9_403; // @[Modules.scala 65:57:@22245.4]
  wire [10:0] buffer_9_41; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70477; // @[Modules.scala 65:57:@22279.4]
  wire [10:0] _T_70478; // @[Modules.scala 65:57:@22280.4]
  wire [10:0] buffer_9_412; // @[Modules.scala 65:57:@22281.4]
  wire [11:0] _T_70501; // @[Modules.scala 65:57:@22311.4]
  wire [10:0] _T_70502; // @[Modules.scala 65:57:@22312.4]
  wire [10:0] buffer_9_420; // @[Modules.scala 65:57:@22313.4]
  wire [11:0] _T_70519; // @[Modules.scala 65:57:@22335.4]
  wire [10:0] _T_70520; // @[Modules.scala 65:57:@22336.4]
  wire [10:0] buffer_9_426; // @[Modules.scala 65:57:@22337.4]
  wire [10:0] buffer_9_75; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70528; // @[Modules.scala 65:57:@22347.4]
  wire [10:0] _T_70529; // @[Modules.scala 65:57:@22348.4]
  wire [10:0] buffer_9_429; // @[Modules.scala 65:57:@22349.4]
  wire [11:0] _T_70531; // @[Modules.scala 65:57:@22351.4]
  wire [10:0] _T_70532; // @[Modules.scala 65:57:@22352.4]
  wire [10:0] buffer_9_430; // @[Modules.scala 65:57:@22353.4]
  wire [10:0] buffer_9_78; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70534; // @[Modules.scala 65:57:@22355.4]
  wire [10:0] _T_70535; // @[Modules.scala 65:57:@22356.4]
  wire [10:0] buffer_9_431; // @[Modules.scala 65:57:@22357.4]
  wire [10:0] buffer_9_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70543; // @[Modules.scala 65:57:@22367.4]
  wire [10:0] _T_70544; // @[Modules.scala 65:57:@22368.4]
  wire [10:0] buffer_9_434; // @[Modules.scala 65:57:@22369.4]
  wire [10:0] buffer_9_91; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70552; // @[Modules.scala 65:57:@22379.4]
  wire [10:0] _T_70553; // @[Modules.scala 65:57:@22380.4]
  wire [10:0] buffer_9_437; // @[Modules.scala 65:57:@22381.4]
  wire [11:0] _T_70561; // @[Modules.scala 65:57:@22391.4]
  wire [10:0] _T_70562; // @[Modules.scala 65:57:@22392.4]
  wire [10:0] buffer_9_440; // @[Modules.scala 65:57:@22393.4]
  wire [11:0] _T_70570; // @[Modules.scala 65:57:@22403.4]
  wire [10:0] _T_70571; // @[Modules.scala 65:57:@22404.4]
  wire [10:0] buffer_9_443; // @[Modules.scala 65:57:@22405.4]
  wire [11:0] _T_70576; // @[Modules.scala 65:57:@22411.4]
  wire [10:0] _T_70577; // @[Modules.scala 65:57:@22412.4]
  wire [10:0] buffer_9_445; // @[Modules.scala 65:57:@22413.4]
  wire [11:0] _T_70579; // @[Modules.scala 65:57:@22415.4]
  wire [10:0] _T_70580; // @[Modules.scala 65:57:@22416.4]
  wire [10:0] buffer_9_446; // @[Modules.scala 65:57:@22417.4]
  wire [11:0] _T_70582; // @[Modules.scala 65:57:@22419.4]
  wire [10:0] _T_70583; // @[Modules.scala 65:57:@22420.4]
  wire [10:0] buffer_9_447; // @[Modules.scala 65:57:@22421.4]
  wire [11:0] _T_70585; // @[Modules.scala 65:57:@22423.4]
  wire [10:0] _T_70586; // @[Modules.scala 65:57:@22424.4]
  wire [10:0] buffer_9_448; // @[Modules.scala 65:57:@22425.4]
  wire [10:0] buffer_9_114; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70588; // @[Modules.scala 65:57:@22427.4]
  wire [10:0] _T_70589; // @[Modules.scala 65:57:@22428.4]
  wire [10:0] buffer_9_449; // @[Modules.scala 65:57:@22429.4]
  wire [11:0] _T_70594; // @[Modules.scala 65:57:@22435.4]
  wire [10:0] _T_70595; // @[Modules.scala 65:57:@22436.4]
  wire [10:0] buffer_9_451; // @[Modules.scala 65:57:@22437.4]
  wire [10:0] buffer_9_122; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70600; // @[Modules.scala 65:57:@22443.4]
  wire [10:0] _T_70601; // @[Modules.scala 65:57:@22444.4]
  wire [10:0] buffer_9_453; // @[Modules.scala 65:57:@22445.4]
  wire [11:0] _T_70609; // @[Modules.scala 65:57:@22455.4]
  wire [10:0] _T_70610; // @[Modules.scala 65:57:@22456.4]
  wire [10:0] buffer_9_456; // @[Modules.scala 65:57:@22457.4]
  wire [10:0] buffer_9_133; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70615; // @[Modules.scala 65:57:@22463.4]
  wire [10:0] _T_70616; // @[Modules.scala 65:57:@22464.4]
  wire [10:0] buffer_9_458; // @[Modules.scala 65:57:@22465.4]
  wire [11:0] _T_70624; // @[Modules.scala 65:57:@22475.4]
  wire [10:0] _T_70625; // @[Modules.scala 65:57:@22476.4]
  wire [10:0] buffer_9_461; // @[Modules.scala 65:57:@22477.4]
  wire [11:0] _T_70627; // @[Modules.scala 65:57:@22479.4]
  wire [10:0] _T_70628; // @[Modules.scala 65:57:@22480.4]
  wire [10:0] buffer_9_462; // @[Modules.scala 65:57:@22481.4]
  wire [11:0] _T_70630; // @[Modules.scala 65:57:@22483.4]
  wire [10:0] _T_70631; // @[Modules.scala 65:57:@22484.4]
  wire [10:0] buffer_9_463; // @[Modules.scala 65:57:@22485.4]
  wire [11:0] _T_70642; // @[Modules.scala 65:57:@22499.4]
  wire [10:0] _T_70643; // @[Modules.scala 65:57:@22500.4]
  wire [10:0] buffer_9_467; // @[Modules.scala 65:57:@22501.4]
  wire [10:0] buffer_9_152; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70645; // @[Modules.scala 65:57:@22503.4]
  wire [10:0] _T_70646; // @[Modules.scala 65:57:@22504.4]
  wire [10:0] buffer_9_468; // @[Modules.scala 65:57:@22505.4]
  wire [10:0] buffer_9_156; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70651; // @[Modules.scala 65:57:@22511.4]
  wire [10:0] _T_70652; // @[Modules.scala 65:57:@22512.4]
  wire [10:0] buffer_9_470; // @[Modules.scala 65:57:@22513.4]
  wire [10:0] buffer_9_160; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70657; // @[Modules.scala 65:57:@22519.4]
  wire [10:0] _T_70658; // @[Modules.scala 65:57:@22520.4]
  wire [10:0] buffer_9_472; // @[Modules.scala 65:57:@22521.4]
  wire [10:0] buffer_9_174; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70678; // @[Modules.scala 65:57:@22547.4]
  wire [10:0] _T_70679; // @[Modules.scala 65:57:@22548.4]
  wire [10:0] buffer_9_479; // @[Modules.scala 65:57:@22549.4]
  wire [11:0] _T_70681; // @[Modules.scala 65:57:@22551.4]
  wire [10:0] _T_70682; // @[Modules.scala 65:57:@22552.4]
  wire [10:0] buffer_9_480; // @[Modules.scala 65:57:@22553.4]
  wire [11:0] _T_70684; // @[Modules.scala 65:57:@22555.4]
  wire [10:0] _T_70685; // @[Modules.scala 65:57:@22556.4]
  wire [10:0] buffer_9_481; // @[Modules.scala 65:57:@22557.4]
  wire [10:0] buffer_9_191; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70702; // @[Modules.scala 65:57:@22579.4]
  wire [10:0] _T_70703; // @[Modules.scala 65:57:@22580.4]
  wire [10:0] buffer_9_487; // @[Modules.scala 65:57:@22581.4]
  wire [11:0] _T_70708; // @[Modules.scala 65:57:@22587.4]
  wire [10:0] _T_70709; // @[Modules.scala 65:57:@22588.4]
  wire [10:0] buffer_9_489; // @[Modules.scala 65:57:@22589.4]
  wire [11:0] _T_70711; // @[Modules.scala 65:57:@22591.4]
  wire [10:0] _T_70712; // @[Modules.scala 65:57:@22592.4]
  wire [10:0] buffer_9_490; // @[Modules.scala 65:57:@22593.4]
  wire [10:0] buffer_9_200; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70717; // @[Modules.scala 65:57:@22599.4]
  wire [10:0] _T_70718; // @[Modules.scala 65:57:@22600.4]
  wire [10:0] buffer_9_492; // @[Modules.scala 65:57:@22601.4]
  wire [11:0] _T_70738; // @[Modules.scala 65:57:@22627.4]
  wire [10:0] _T_70739; // @[Modules.scala 65:57:@22628.4]
  wire [10:0] buffer_9_499; // @[Modules.scala 65:57:@22629.4]
  wire [11:0] _T_70753; // @[Modules.scala 65:57:@22647.4]
  wire [10:0] _T_70754; // @[Modules.scala 65:57:@22648.4]
  wire [10:0] buffer_9_504; // @[Modules.scala 65:57:@22649.4]
  wire [10:0] buffer_9_226; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70756; // @[Modules.scala 65:57:@22651.4]
  wire [10:0] _T_70757; // @[Modules.scala 65:57:@22652.4]
  wire [10:0] buffer_9_505; // @[Modules.scala 65:57:@22653.4]
  wire [11:0] _T_70759; // @[Modules.scala 65:57:@22655.4]
  wire [10:0] _T_70760; // @[Modules.scala 65:57:@22656.4]
  wire [10:0] buffer_9_506; // @[Modules.scala 65:57:@22657.4]
  wire [11:0] _T_70777; // @[Modules.scala 65:57:@22679.4]
  wire [10:0] _T_70778; // @[Modules.scala 65:57:@22680.4]
  wire [10:0] buffer_9_512; // @[Modules.scala 65:57:@22681.4]
  wire [10:0] buffer_9_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70783; // @[Modules.scala 65:57:@22687.4]
  wire [10:0] _T_70784; // @[Modules.scala 65:57:@22688.4]
  wire [10:0] buffer_9_514; // @[Modules.scala 65:57:@22689.4]
  wire [11:0] _T_70798; // @[Modules.scala 65:57:@22707.4]
  wire [10:0] _T_70799; // @[Modules.scala 65:57:@22708.4]
  wire [10:0] buffer_9_519; // @[Modules.scala 65:57:@22709.4]
  wire [11:0] _T_70819; // @[Modules.scala 65:57:@22735.4]
  wire [10:0] _T_70820; // @[Modules.scala 65:57:@22736.4]
  wire [10:0] buffer_9_526; // @[Modules.scala 65:57:@22737.4]
  wire [10:0] buffer_9_283; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70840; // @[Modules.scala 65:57:@22763.4]
  wire [10:0] _T_70841; // @[Modules.scala 65:57:@22764.4]
  wire [10:0] buffer_9_533; // @[Modules.scala 65:57:@22765.4]
  wire [11:0] _T_70843; // @[Modules.scala 65:57:@22767.4]
  wire [10:0] _T_70844; // @[Modules.scala 65:57:@22768.4]
  wire [10:0] buffer_9_534; // @[Modules.scala 65:57:@22769.4]
  wire [11:0] _T_70846; // @[Modules.scala 65:57:@22771.4]
  wire [10:0] _T_70847; // @[Modules.scala 65:57:@22772.4]
  wire [10:0] buffer_9_535; // @[Modules.scala 65:57:@22773.4]
  wire [11:0] _T_70864; // @[Modules.scala 65:57:@22795.4]
  wire [10:0] _T_70865; // @[Modules.scala 65:57:@22796.4]
  wire [10:0] buffer_9_541; // @[Modules.scala 65:57:@22797.4]
  wire [10:0] buffer_9_300; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70867; // @[Modules.scala 65:57:@22799.4]
  wire [10:0] _T_70868; // @[Modules.scala 65:57:@22800.4]
  wire [10:0] buffer_9_542; // @[Modules.scala 65:57:@22801.4]
  wire [10:0] buffer_9_304; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_9_305; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70873; // @[Modules.scala 65:57:@22807.4]
  wire [10:0] _T_70874; // @[Modules.scala 65:57:@22808.4]
  wire [10:0] buffer_9_544; // @[Modules.scala 65:57:@22809.4]
  wire [11:0] _T_70885; // @[Modules.scala 65:57:@22823.4]
  wire [10:0] _T_70886; // @[Modules.scala 65:57:@22824.4]
  wire [10:0] buffer_9_548; // @[Modules.scala 65:57:@22825.4]
  wire [11:0] _T_70891; // @[Modules.scala 65:57:@22831.4]
  wire [10:0] _T_70892; // @[Modules.scala 65:57:@22832.4]
  wire [10:0] buffer_9_550; // @[Modules.scala 65:57:@22833.4]
  wire [11:0] _T_70894; // @[Modules.scala 65:57:@22835.4]
  wire [10:0] _T_70895; // @[Modules.scala 65:57:@22836.4]
  wire [10:0] buffer_9_551; // @[Modules.scala 65:57:@22837.4]
  wire [10:0] buffer_9_320; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70897; // @[Modules.scala 65:57:@22839.4]
  wire [10:0] _T_70898; // @[Modules.scala 65:57:@22840.4]
  wire [10:0] buffer_9_552; // @[Modules.scala 65:57:@22841.4]
  wire [11:0] _T_70906; // @[Modules.scala 65:57:@22851.4]
  wire [10:0] _T_70907; // @[Modules.scala 65:57:@22852.4]
  wire [10:0] buffer_9_555; // @[Modules.scala 65:57:@22853.4]
  wire [11:0] _T_70915; // @[Modules.scala 65:57:@22863.4]
  wire [10:0] _T_70916; // @[Modules.scala 65:57:@22864.4]
  wire [10:0] buffer_9_558; // @[Modules.scala 65:57:@22865.4]
  wire [10:0] buffer_9_346; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_9_347; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70936; // @[Modules.scala 65:57:@22891.4]
  wire [10:0] _T_70937; // @[Modules.scala 65:57:@22892.4]
  wire [10:0] buffer_9_565; // @[Modules.scala 65:57:@22893.4]
  wire [11:0] _T_70939; // @[Modules.scala 65:57:@22895.4]
  wire [10:0] _T_70940; // @[Modules.scala 65:57:@22896.4]
  wire [10:0] buffer_9_566; // @[Modules.scala 65:57:@22897.4]
  wire [11:0] _T_70942; // @[Modules.scala 65:57:@22899.4]
  wire [10:0] _T_70943; // @[Modules.scala 65:57:@22900.4]
  wire [10:0] buffer_9_567; // @[Modules.scala 65:57:@22901.4]
  wire [10:0] buffer_9_354; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70948; // @[Modules.scala 65:57:@22907.4]
  wire [10:0] _T_70949; // @[Modules.scala 65:57:@22908.4]
  wire [10:0] buffer_9_569; // @[Modules.scala 65:57:@22909.4]
  wire [10:0] buffer_9_356; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70951; // @[Modules.scala 65:57:@22911.4]
  wire [10:0] _T_70952; // @[Modules.scala 65:57:@22912.4]
  wire [10:0] buffer_9_570; // @[Modules.scala 65:57:@22913.4]
  wire [10:0] buffer_9_358; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70954; // @[Modules.scala 65:57:@22915.4]
  wire [10:0] _T_70955; // @[Modules.scala 65:57:@22916.4]
  wire [10:0] buffer_9_571; // @[Modules.scala 65:57:@22917.4]
  wire [10:0] buffer_9_362; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70960; // @[Modules.scala 65:57:@22923.4]
  wire [10:0] _T_70961; // @[Modules.scala 65:57:@22924.4]
  wire [10:0] buffer_9_573; // @[Modules.scala 65:57:@22925.4]
  wire [10:0] buffer_9_364; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70963; // @[Modules.scala 65:57:@22927.4]
  wire [10:0] _T_70964; // @[Modules.scala 65:57:@22928.4]
  wire [10:0] buffer_9_574; // @[Modules.scala 65:57:@22929.4]
  wire [11:0] _T_70975; // @[Modules.scala 65:57:@22943.4]
  wire [10:0] _T_70976; // @[Modules.scala 65:57:@22944.4]
  wire [10:0] buffer_9_578; // @[Modules.scala 65:57:@22945.4]
  wire [11:0] _T_70978; // @[Modules.scala 65:57:@22947.4]
  wire [10:0] _T_70979; // @[Modules.scala 65:57:@22948.4]
  wire [10:0] buffer_9_579; // @[Modules.scala 65:57:@22949.4]
  wire [11:0] _T_70981; // @[Modules.scala 65:57:@22951.4]
  wire [10:0] _T_70982; // @[Modules.scala 65:57:@22952.4]
  wire [10:0] buffer_9_580; // @[Modules.scala 65:57:@22953.4]
  wire [10:0] buffer_9_379; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70984; // @[Modules.scala 65:57:@22955.4]
  wire [10:0] _T_70985; // @[Modules.scala 65:57:@22956.4]
  wire [10:0] buffer_9_581; // @[Modules.scala 65:57:@22957.4]
  wire [10:0] buffer_9_381; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70987; // @[Modules.scala 65:57:@22959.4]
  wire [10:0] _T_70988; // @[Modules.scala 65:57:@22960.4]
  wire [10:0] buffer_9_582; // @[Modules.scala 65:57:@22961.4]
  wire [11:0] _T_70990; // @[Modules.scala 65:57:@22963.4]
  wire [10:0] _T_70991; // @[Modules.scala 65:57:@22964.4]
  wire [10:0] buffer_9_583; // @[Modules.scala 65:57:@22965.4]
  wire [10:0] buffer_9_387; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_70996; // @[Modules.scala 65:57:@22971.4]
  wire [10:0] _T_70997; // @[Modules.scala 65:57:@22972.4]
  wire [10:0] buffer_9_585; // @[Modules.scala 65:57:@22973.4]
  wire [11:0] _T_71005; // @[Modules.scala 68:83:@22983.4]
  wire [10:0] _T_71006; // @[Modules.scala 68:83:@22984.4]
  wire [10:0] buffer_9_588; // @[Modules.scala 68:83:@22985.4]
  wire [11:0] _T_71011; // @[Modules.scala 68:83:@22991.4]
  wire [10:0] _T_71012; // @[Modules.scala 68:83:@22992.4]
  wire [10:0] buffer_9_590; // @[Modules.scala 68:83:@22993.4]
  wire [11:0] _T_71014; // @[Modules.scala 68:83:@22995.4]
  wire [10:0] _T_71015; // @[Modules.scala 68:83:@22996.4]
  wire [10:0] buffer_9_591; // @[Modules.scala 68:83:@22997.4]
  wire [11:0] _T_71020; // @[Modules.scala 68:83:@23003.4]
  wire [10:0] _T_71021; // @[Modules.scala 68:83:@23004.4]
  wire [10:0] buffer_9_593; // @[Modules.scala 68:83:@23005.4]
  wire [11:0] _T_71023; // @[Modules.scala 68:83:@23007.4]
  wire [10:0] _T_71024; // @[Modules.scala 68:83:@23008.4]
  wire [10:0] buffer_9_594; // @[Modules.scala 68:83:@23009.4]
  wire [11:0] _T_71026; // @[Modules.scala 68:83:@23011.4]
  wire [10:0] _T_71027; // @[Modules.scala 68:83:@23012.4]
  wire [10:0] buffer_9_595; // @[Modules.scala 68:83:@23013.4]
  wire [11:0] _T_71035; // @[Modules.scala 68:83:@23023.4]
  wire [10:0] _T_71036; // @[Modules.scala 68:83:@23024.4]
  wire [10:0] buffer_9_598; // @[Modules.scala 68:83:@23025.4]
  wire [11:0] _T_71047; // @[Modules.scala 68:83:@23039.4]
  wire [10:0] _T_71048; // @[Modules.scala 68:83:@23040.4]
  wire [10:0] buffer_9_602; // @[Modules.scala 68:83:@23041.4]
  wire [11:0] _T_71053; // @[Modules.scala 68:83:@23047.4]
  wire [10:0] _T_71054; // @[Modules.scala 68:83:@23048.4]
  wire [10:0] buffer_9_604; // @[Modules.scala 68:83:@23049.4]
  wire [11:0] _T_71056; // @[Modules.scala 68:83:@23051.4]
  wire [10:0] _T_71057; // @[Modules.scala 68:83:@23052.4]
  wire [10:0] buffer_9_605; // @[Modules.scala 68:83:@23053.4]
  wire [11:0] _T_71059; // @[Modules.scala 68:83:@23055.4]
  wire [10:0] _T_71060; // @[Modules.scala 68:83:@23056.4]
  wire [10:0] buffer_9_606; // @[Modules.scala 68:83:@23057.4]
  wire [11:0] _T_71062; // @[Modules.scala 68:83:@23059.4]
  wire [10:0] _T_71063; // @[Modules.scala 68:83:@23060.4]
  wire [10:0] buffer_9_607; // @[Modules.scala 68:83:@23061.4]
  wire [11:0] _T_71065; // @[Modules.scala 68:83:@23063.4]
  wire [10:0] _T_71066; // @[Modules.scala 68:83:@23064.4]
  wire [10:0] buffer_9_608; // @[Modules.scala 68:83:@23065.4]
  wire [11:0] _T_71068; // @[Modules.scala 68:83:@23067.4]
  wire [10:0] _T_71069; // @[Modules.scala 68:83:@23068.4]
  wire [10:0] buffer_9_609; // @[Modules.scala 68:83:@23069.4]
  wire [11:0] _T_71071; // @[Modules.scala 68:83:@23071.4]
  wire [10:0] _T_71072; // @[Modules.scala 68:83:@23072.4]
  wire [10:0] buffer_9_610; // @[Modules.scala 68:83:@23073.4]
  wire [11:0] _T_71074; // @[Modules.scala 68:83:@23075.4]
  wire [10:0] _T_71075; // @[Modules.scala 68:83:@23076.4]
  wire [10:0] buffer_9_611; // @[Modules.scala 68:83:@23077.4]
  wire [11:0] _T_71077; // @[Modules.scala 68:83:@23079.4]
  wire [10:0] _T_71078; // @[Modules.scala 68:83:@23080.4]
  wire [10:0] buffer_9_612; // @[Modules.scala 68:83:@23081.4]
  wire [11:0] _T_71080; // @[Modules.scala 68:83:@23083.4]
  wire [10:0] _T_71081; // @[Modules.scala 68:83:@23084.4]
  wire [10:0] buffer_9_613; // @[Modules.scala 68:83:@23085.4]
  wire [11:0] _T_71083; // @[Modules.scala 68:83:@23087.4]
  wire [10:0] _T_71084; // @[Modules.scala 68:83:@23088.4]
  wire [10:0] buffer_9_614; // @[Modules.scala 68:83:@23089.4]
  wire [11:0] _T_71086; // @[Modules.scala 68:83:@23091.4]
  wire [10:0] _T_71087; // @[Modules.scala 68:83:@23092.4]
  wire [10:0] buffer_9_615; // @[Modules.scala 68:83:@23093.4]
  wire [11:0] _T_71089; // @[Modules.scala 68:83:@23095.4]
  wire [10:0] _T_71090; // @[Modules.scala 68:83:@23096.4]
  wire [10:0] buffer_9_616; // @[Modules.scala 68:83:@23097.4]
  wire [11:0] _T_71092; // @[Modules.scala 68:83:@23099.4]
  wire [10:0] _T_71093; // @[Modules.scala 68:83:@23100.4]
  wire [10:0] buffer_9_617; // @[Modules.scala 68:83:@23101.4]
  wire [11:0] _T_71095; // @[Modules.scala 68:83:@23103.4]
  wire [10:0] _T_71096; // @[Modules.scala 68:83:@23104.4]
  wire [10:0] buffer_9_618; // @[Modules.scala 68:83:@23105.4]
  wire [11:0] _T_71101; // @[Modules.scala 68:83:@23111.4]
  wire [10:0] _T_71102; // @[Modules.scala 68:83:@23112.4]
  wire [10:0] buffer_9_620; // @[Modules.scala 68:83:@23113.4]
  wire [11:0] _T_71104; // @[Modules.scala 68:83:@23115.4]
  wire [10:0] _T_71105; // @[Modules.scala 68:83:@23116.4]
  wire [10:0] buffer_9_621; // @[Modules.scala 68:83:@23117.4]
  wire [11:0] _T_71107; // @[Modules.scala 68:83:@23119.4]
  wire [10:0] _T_71108; // @[Modules.scala 68:83:@23120.4]
  wire [10:0] buffer_9_622; // @[Modules.scala 68:83:@23121.4]
  wire [11:0] _T_71110; // @[Modules.scala 68:83:@23123.4]
  wire [10:0] _T_71111; // @[Modules.scala 68:83:@23124.4]
  wire [10:0] buffer_9_623; // @[Modules.scala 68:83:@23125.4]
  wire [11:0] _T_71116; // @[Modules.scala 68:83:@23131.4]
  wire [10:0] _T_71117; // @[Modules.scala 68:83:@23132.4]
  wire [10:0] buffer_9_625; // @[Modules.scala 68:83:@23133.4]
  wire [11:0] _T_71119; // @[Modules.scala 68:83:@23135.4]
  wire [10:0] _T_71120; // @[Modules.scala 68:83:@23136.4]
  wire [10:0] buffer_9_626; // @[Modules.scala 68:83:@23137.4]
  wire [11:0] _T_71122; // @[Modules.scala 68:83:@23139.4]
  wire [10:0] _T_71123; // @[Modules.scala 68:83:@23140.4]
  wire [10:0] buffer_9_627; // @[Modules.scala 68:83:@23141.4]
  wire [11:0] _T_71125; // @[Modules.scala 68:83:@23143.4]
  wire [10:0] _T_71126; // @[Modules.scala 68:83:@23144.4]
  wire [10:0] buffer_9_628; // @[Modules.scala 68:83:@23145.4]
  wire [11:0] _T_71128; // @[Modules.scala 68:83:@23147.4]
  wire [10:0] _T_71129; // @[Modules.scala 68:83:@23148.4]
  wire [10:0] buffer_9_629; // @[Modules.scala 68:83:@23149.4]
  wire [11:0] _T_71134; // @[Modules.scala 68:83:@23155.4]
  wire [10:0] _T_71135; // @[Modules.scala 68:83:@23156.4]
  wire [10:0] buffer_9_631; // @[Modules.scala 68:83:@23157.4]
  wire [11:0] _T_71137; // @[Modules.scala 68:83:@23159.4]
  wire [10:0] _T_71138; // @[Modules.scala 68:83:@23160.4]
  wire [10:0] buffer_9_632; // @[Modules.scala 68:83:@23161.4]
  wire [11:0] _T_71146; // @[Modules.scala 68:83:@23171.4]
  wire [10:0] _T_71147; // @[Modules.scala 68:83:@23172.4]
  wire [10:0] buffer_9_635; // @[Modules.scala 68:83:@23173.4]
  wire [11:0] _T_71149; // @[Modules.scala 68:83:@23175.4]
  wire [10:0] _T_71150; // @[Modules.scala 68:83:@23176.4]
  wire [10:0] buffer_9_636; // @[Modules.scala 68:83:@23177.4]
  wire [11:0] _T_71152; // @[Modules.scala 68:83:@23179.4]
  wire [10:0] _T_71153; // @[Modules.scala 68:83:@23180.4]
  wire [10:0] buffer_9_637; // @[Modules.scala 68:83:@23181.4]
  wire [11:0] _T_71155; // @[Modules.scala 68:83:@23183.4]
  wire [10:0] _T_71156; // @[Modules.scala 68:83:@23184.4]
  wire [10:0] buffer_9_638; // @[Modules.scala 68:83:@23185.4]
  wire [11:0] _T_71161; // @[Modules.scala 68:83:@23191.4]
  wire [10:0] _T_71162; // @[Modules.scala 68:83:@23192.4]
  wire [10:0] buffer_9_640; // @[Modules.scala 68:83:@23193.4]
  wire [11:0] _T_71164; // @[Modules.scala 68:83:@23195.4]
  wire [10:0] _T_71165; // @[Modules.scala 68:83:@23196.4]
  wire [10:0] buffer_9_641; // @[Modules.scala 68:83:@23197.4]
  wire [11:0] _T_71173; // @[Modules.scala 68:83:@23207.4]
  wire [10:0] _T_71174; // @[Modules.scala 68:83:@23208.4]
  wire [10:0] buffer_9_644; // @[Modules.scala 68:83:@23209.4]
  wire [11:0] _T_71176; // @[Modules.scala 68:83:@23211.4]
  wire [10:0] _T_71177; // @[Modules.scala 68:83:@23212.4]
  wire [10:0] buffer_9_645; // @[Modules.scala 68:83:@23213.4]
  wire [11:0] _T_71185; // @[Modules.scala 68:83:@23223.4]
  wire [10:0] _T_71186; // @[Modules.scala 68:83:@23224.4]
  wire [10:0] buffer_9_648; // @[Modules.scala 68:83:@23225.4]
  wire [11:0] _T_71188; // @[Modules.scala 68:83:@23227.4]
  wire [10:0] _T_71189; // @[Modules.scala 68:83:@23228.4]
  wire [10:0] buffer_9_649; // @[Modules.scala 68:83:@23229.4]
  wire [11:0] _T_71194; // @[Modules.scala 68:83:@23235.4]
  wire [10:0] _T_71195; // @[Modules.scala 68:83:@23236.4]
  wire [10:0] buffer_9_651; // @[Modules.scala 68:83:@23237.4]
  wire [11:0] _T_71206; // @[Modules.scala 68:83:@23251.4]
  wire [10:0] _T_71207; // @[Modules.scala 68:83:@23252.4]
  wire [10:0] buffer_9_655; // @[Modules.scala 68:83:@23253.4]
  wire [11:0] _T_71215; // @[Modules.scala 68:83:@23263.4]
  wire [10:0] _T_71216; // @[Modules.scala 68:83:@23264.4]
  wire [10:0] buffer_9_658; // @[Modules.scala 68:83:@23265.4]
  wire [11:0] _T_71218; // @[Modules.scala 68:83:@23267.4]
  wire [10:0] _T_71219; // @[Modules.scala 68:83:@23268.4]
  wire [10:0] buffer_9_659; // @[Modules.scala 68:83:@23269.4]
  wire [11:0] _T_71224; // @[Modules.scala 68:83:@23275.4]
  wire [10:0] _T_71225; // @[Modules.scala 68:83:@23276.4]
  wire [10:0] buffer_9_661; // @[Modules.scala 68:83:@23277.4]
  wire [11:0] _T_71227; // @[Modules.scala 68:83:@23279.4]
  wire [10:0] _T_71228; // @[Modules.scala 68:83:@23280.4]
  wire [10:0] buffer_9_662; // @[Modules.scala 68:83:@23281.4]
  wire [11:0] _T_71230; // @[Modules.scala 68:83:@23283.4]
  wire [10:0] _T_71231; // @[Modules.scala 68:83:@23284.4]
  wire [10:0] buffer_9_663; // @[Modules.scala 68:83:@23285.4]
  wire [11:0] _T_71233; // @[Modules.scala 68:83:@23287.4]
  wire [10:0] _T_71234; // @[Modules.scala 68:83:@23288.4]
  wire [10:0] buffer_9_664; // @[Modules.scala 68:83:@23289.4]
  wire [11:0] _T_71239; // @[Modules.scala 68:83:@23295.4]
  wire [10:0] _T_71240; // @[Modules.scala 68:83:@23296.4]
  wire [10:0] buffer_9_666; // @[Modules.scala 68:83:@23297.4]
  wire [11:0] _T_71242; // @[Modules.scala 68:83:@23299.4]
  wire [10:0] _T_71243; // @[Modules.scala 68:83:@23300.4]
  wire [10:0] buffer_9_667; // @[Modules.scala 68:83:@23301.4]
  wire [11:0] _T_71245; // @[Modules.scala 68:83:@23303.4]
  wire [10:0] _T_71246; // @[Modules.scala 68:83:@23304.4]
  wire [10:0] buffer_9_668; // @[Modules.scala 68:83:@23305.4]
  wire [11:0] _T_71248; // @[Modules.scala 68:83:@23307.4]
  wire [10:0] _T_71249; // @[Modules.scala 68:83:@23308.4]
  wire [10:0] buffer_9_669; // @[Modules.scala 68:83:@23309.4]
  wire [11:0] _T_71254; // @[Modules.scala 68:83:@23315.4]
  wire [10:0] _T_71255; // @[Modules.scala 68:83:@23316.4]
  wire [10:0] buffer_9_671; // @[Modules.scala 68:83:@23317.4]
  wire [11:0] _T_71257; // @[Modules.scala 68:83:@23319.4]
  wire [10:0] _T_71258; // @[Modules.scala 68:83:@23320.4]
  wire [10:0] buffer_9_672; // @[Modules.scala 68:83:@23321.4]
  wire [11:0] _T_71263; // @[Modules.scala 68:83:@23327.4]
  wire [10:0] _T_71264; // @[Modules.scala 68:83:@23328.4]
  wire [10:0] buffer_9_674; // @[Modules.scala 68:83:@23329.4]
  wire [11:0] _T_71266; // @[Modules.scala 68:83:@23331.4]
  wire [10:0] _T_71267; // @[Modules.scala 68:83:@23332.4]
  wire [10:0] buffer_9_675; // @[Modules.scala 68:83:@23333.4]
  wire [11:0] _T_71269; // @[Modules.scala 68:83:@23335.4]
  wire [10:0] _T_71270; // @[Modules.scala 68:83:@23336.4]
  wire [10:0] buffer_9_676; // @[Modules.scala 68:83:@23337.4]
  wire [11:0] _T_71272; // @[Modules.scala 68:83:@23339.4]
  wire [10:0] _T_71273; // @[Modules.scala 68:83:@23340.4]
  wire [10:0] buffer_9_677; // @[Modules.scala 68:83:@23341.4]
  wire [11:0] _T_71275; // @[Modules.scala 68:83:@23343.4]
  wire [10:0] _T_71276; // @[Modules.scala 68:83:@23344.4]
  wire [10:0] buffer_9_678; // @[Modules.scala 68:83:@23345.4]
  wire [11:0] _T_71278; // @[Modules.scala 68:83:@23347.4]
  wire [10:0] _T_71279; // @[Modules.scala 68:83:@23348.4]
  wire [10:0] buffer_9_679; // @[Modules.scala 68:83:@23349.4]
  wire [11:0] _T_71284; // @[Modules.scala 68:83:@23355.4]
  wire [10:0] _T_71285; // @[Modules.scala 68:83:@23356.4]
  wire [10:0] buffer_9_681; // @[Modules.scala 68:83:@23357.4]
  wire [11:0] _T_71287; // @[Modules.scala 68:83:@23359.4]
  wire [10:0] _T_71288; // @[Modules.scala 68:83:@23360.4]
  wire [10:0] buffer_9_682; // @[Modules.scala 68:83:@23361.4]
  wire [11:0] _T_71290; // @[Modules.scala 68:83:@23363.4]
  wire [10:0] _T_71291; // @[Modules.scala 68:83:@23364.4]
  wire [10:0] buffer_9_683; // @[Modules.scala 68:83:@23365.4]
  wire [11:0] _T_71293; // @[Modules.scala 68:83:@23367.4]
  wire [10:0] _T_71294; // @[Modules.scala 68:83:@23368.4]
  wire [10:0] buffer_9_684; // @[Modules.scala 68:83:@23369.4]
  wire [11:0] _T_71299; // @[Modules.scala 71:109:@23375.4]
  wire [10:0] _T_71300; // @[Modules.scala 71:109:@23376.4]
  wire [10:0] buffer_9_686; // @[Modules.scala 71:109:@23377.4]
  wire [11:0] _T_71302; // @[Modules.scala 71:109:@23379.4]
  wire [10:0] _T_71303; // @[Modules.scala 71:109:@23380.4]
  wire [10:0] buffer_9_687; // @[Modules.scala 71:109:@23381.4]
  wire [11:0] _T_71305; // @[Modules.scala 71:109:@23383.4]
  wire [10:0] _T_71306; // @[Modules.scala 71:109:@23384.4]
  wire [10:0] buffer_9_688; // @[Modules.scala 71:109:@23385.4]
  wire [11:0] _T_71308; // @[Modules.scala 71:109:@23387.4]
  wire [10:0] _T_71309; // @[Modules.scala 71:109:@23388.4]
  wire [10:0] buffer_9_689; // @[Modules.scala 71:109:@23389.4]
  wire [11:0] _T_71314; // @[Modules.scala 71:109:@23395.4]
  wire [10:0] _T_71315; // @[Modules.scala 71:109:@23396.4]
  wire [10:0] buffer_9_691; // @[Modules.scala 71:109:@23397.4]
  wire [11:0] _T_71320; // @[Modules.scala 71:109:@23403.4]
  wire [10:0] _T_71321; // @[Modules.scala 71:109:@23404.4]
  wire [10:0] buffer_9_693; // @[Modules.scala 71:109:@23405.4]
  wire [11:0] _T_71323; // @[Modules.scala 71:109:@23407.4]
  wire [10:0] _T_71324; // @[Modules.scala 71:109:@23408.4]
  wire [10:0] buffer_9_694; // @[Modules.scala 71:109:@23409.4]
  wire [11:0] _T_71326; // @[Modules.scala 71:109:@23411.4]
  wire [10:0] _T_71327; // @[Modules.scala 71:109:@23412.4]
  wire [10:0] buffer_9_695; // @[Modules.scala 71:109:@23413.4]
  wire [11:0] _T_71329; // @[Modules.scala 71:109:@23415.4]
  wire [10:0] _T_71330; // @[Modules.scala 71:109:@23416.4]
  wire [10:0] buffer_9_696; // @[Modules.scala 71:109:@23417.4]
  wire [11:0] _T_71332; // @[Modules.scala 71:109:@23419.4]
  wire [10:0] _T_71333; // @[Modules.scala 71:109:@23420.4]
  wire [10:0] buffer_9_697; // @[Modules.scala 71:109:@23421.4]
  wire [11:0] _T_71335; // @[Modules.scala 71:109:@23423.4]
  wire [10:0] _T_71336; // @[Modules.scala 71:109:@23424.4]
  wire [10:0] buffer_9_698; // @[Modules.scala 71:109:@23425.4]
  wire [11:0] _T_71338; // @[Modules.scala 71:109:@23427.4]
  wire [10:0] _T_71339; // @[Modules.scala 71:109:@23428.4]
  wire [10:0] buffer_9_699; // @[Modules.scala 71:109:@23429.4]
  wire [11:0] _T_71341; // @[Modules.scala 71:109:@23431.4]
  wire [10:0] _T_71342; // @[Modules.scala 71:109:@23432.4]
  wire [10:0] buffer_9_700; // @[Modules.scala 71:109:@23433.4]
  wire [11:0] _T_71344; // @[Modules.scala 71:109:@23435.4]
  wire [10:0] _T_71345; // @[Modules.scala 71:109:@23436.4]
  wire [10:0] buffer_9_701; // @[Modules.scala 71:109:@23437.4]
  wire [11:0] _T_71347; // @[Modules.scala 71:109:@23439.4]
  wire [10:0] _T_71348; // @[Modules.scala 71:109:@23440.4]
  wire [10:0] buffer_9_702; // @[Modules.scala 71:109:@23441.4]
  wire [11:0] _T_71350; // @[Modules.scala 71:109:@23443.4]
  wire [10:0] _T_71351; // @[Modules.scala 71:109:@23444.4]
  wire [10:0] buffer_9_703; // @[Modules.scala 71:109:@23445.4]
  wire [11:0] _T_71353; // @[Modules.scala 71:109:@23447.4]
  wire [10:0] _T_71354; // @[Modules.scala 71:109:@23448.4]
  wire [10:0] buffer_9_704; // @[Modules.scala 71:109:@23449.4]
  wire [11:0] _T_71356; // @[Modules.scala 71:109:@23451.4]
  wire [10:0] _T_71357; // @[Modules.scala 71:109:@23452.4]
  wire [10:0] buffer_9_705; // @[Modules.scala 71:109:@23453.4]
  wire [11:0] _T_71359; // @[Modules.scala 71:109:@23455.4]
  wire [10:0] _T_71360; // @[Modules.scala 71:109:@23456.4]
  wire [10:0] buffer_9_706; // @[Modules.scala 71:109:@23457.4]
  wire [11:0] _T_71362; // @[Modules.scala 71:109:@23459.4]
  wire [10:0] _T_71363; // @[Modules.scala 71:109:@23460.4]
  wire [10:0] buffer_9_707; // @[Modules.scala 71:109:@23461.4]
  wire [11:0] _T_71365; // @[Modules.scala 71:109:@23463.4]
  wire [10:0] _T_71366; // @[Modules.scala 71:109:@23464.4]
  wire [10:0] buffer_9_708; // @[Modules.scala 71:109:@23465.4]
  wire [11:0] _T_71368; // @[Modules.scala 71:109:@23467.4]
  wire [10:0] _T_71369; // @[Modules.scala 71:109:@23468.4]
  wire [10:0] buffer_9_709; // @[Modules.scala 71:109:@23469.4]
  wire [11:0] _T_71371; // @[Modules.scala 71:109:@23471.4]
  wire [10:0] _T_71372; // @[Modules.scala 71:109:@23472.4]
  wire [10:0] buffer_9_710; // @[Modules.scala 71:109:@23473.4]
  wire [11:0] _T_71374; // @[Modules.scala 71:109:@23475.4]
  wire [10:0] _T_71375; // @[Modules.scala 71:109:@23476.4]
  wire [10:0] buffer_9_711; // @[Modules.scala 71:109:@23477.4]
  wire [11:0] _T_71377; // @[Modules.scala 71:109:@23479.4]
  wire [10:0] _T_71378; // @[Modules.scala 71:109:@23480.4]
  wire [10:0] buffer_9_712; // @[Modules.scala 71:109:@23481.4]
  wire [11:0] _T_71380; // @[Modules.scala 71:109:@23483.4]
  wire [10:0] _T_71381; // @[Modules.scala 71:109:@23484.4]
  wire [10:0] buffer_9_713; // @[Modules.scala 71:109:@23485.4]
  wire [11:0] _T_71383; // @[Modules.scala 71:109:@23487.4]
  wire [10:0] _T_71384; // @[Modules.scala 71:109:@23488.4]
  wire [10:0] buffer_9_714; // @[Modules.scala 71:109:@23489.4]
  wire [11:0] _T_71386; // @[Modules.scala 71:109:@23491.4]
  wire [10:0] _T_71387; // @[Modules.scala 71:109:@23492.4]
  wire [10:0] buffer_9_715; // @[Modules.scala 71:109:@23493.4]
  wire [11:0] _T_71389; // @[Modules.scala 71:109:@23495.4]
  wire [10:0] _T_71390; // @[Modules.scala 71:109:@23496.4]
  wire [10:0] buffer_9_716; // @[Modules.scala 71:109:@23497.4]
  wire [11:0] _T_71392; // @[Modules.scala 71:109:@23499.4]
  wire [10:0] _T_71393; // @[Modules.scala 71:109:@23500.4]
  wire [10:0] buffer_9_717; // @[Modules.scala 71:109:@23501.4]
  wire [11:0] _T_71395; // @[Modules.scala 71:109:@23503.4]
  wire [10:0] _T_71396; // @[Modules.scala 71:109:@23504.4]
  wire [10:0] buffer_9_718; // @[Modules.scala 71:109:@23505.4]
  wire [11:0] _T_71398; // @[Modules.scala 71:109:@23507.4]
  wire [10:0] _T_71399; // @[Modules.scala 71:109:@23508.4]
  wire [10:0] buffer_9_719; // @[Modules.scala 71:109:@23509.4]
  wire [11:0] _T_71401; // @[Modules.scala 71:109:@23511.4]
  wire [10:0] _T_71402; // @[Modules.scala 71:109:@23512.4]
  wire [10:0] buffer_9_720; // @[Modules.scala 71:109:@23513.4]
  wire [11:0] _T_71404; // @[Modules.scala 71:109:@23515.4]
  wire [10:0] _T_71405; // @[Modules.scala 71:109:@23516.4]
  wire [10:0] buffer_9_721; // @[Modules.scala 71:109:@23517.4]
  wire [11:0] _T_71407; // @[Modules.scala 71:109:@23519.4]
  wire [10:0] _T_71408; // @[Modules.scala 71:109:@23520.4]
  wire [10:0] buffer_9_722; // @[Modules.scala 71:109:@23521.4]
  wire [11:0] _T_71410; // @[Modules.scala 71:109:@23523.4]
  wire [10:0] _T_71411; // @[Modules.scala 71:109:@23524.4]
  wire [10:0] buffer_9_723; // @[Modules.scala 71:109:@23525.4]
  wire [11:0] _T_71413; // @[Modules.scala 71:109:@23527.4]
  wire [10:0] _T_71414; // @[Modules.scala 71:109:@23528.4]
  wire [10:0] buffer_9_724; // @[Modules.scala 71:109:@23529.4]
  wire [11:0] _T_71416; // @[Modules.scala 71:109:@23531.4]
  wire [10:0] _T_71417; // @[Modules.scala 71:109:@23532.4]
  wire [10:0] buffer_9_725; // @[Modules.scala 71:109:@23533.4]
  wire [11:0] _T_71419; // @[Modules.scala 71:109:@23535.4]
  wire [10:0] _T_71420; // @[Modules.scala 71:109:@23536.4]
  wire [10:0] buffer_9_726; // @[Modules.scala 71:109:@23537.4]
  wire [11:0] _T_71422; // @[Modules.scala 71:109:@23539.4]
  wire [10:0] _T_71423; // @[Modules.scala 71:109:@23540.4]
  wire [10:0] buffer_9_727; // @[Modules.scala 71:109:@23541.4]
  wire [11:0] _T_71425; // @[Modules.scala 71:109:@23543.4]
  wire [10:0] _T_71426; // @[Modules.scala 71:109:@23544.4]
  wire [10:0] buffer_9_728; // @[Modules.scala 71:109:@23545.4]
  wire [11:0] _T_71428; // @[Modules.scala 71:109:@23547.4]
  wire [10:0] _T_71429; // @[Modules.scala 71:109:@23548.4]
  wire [10:0] buffer_9_729; // @[Modules.scala 71:109:@23549.4]
  wire [11:0] _T_71431; // @[Modules.scala 71:109:@23551.4]
  wire [10:0] _T_71432; // @[Modules.scala 71:109:@23552.4]
  wire [10:0] buffer_9_730; // @[Modules.scala 71:109:@23553.4]
  wire [11:0] _T_71434; // @[Modules.scala 71:109:@23555.4]
  wire [10:0] _T_71435; // @[Modules.scala 71:109:@23556.4]
  wire [10:0] buffer_9_731; // @[Modules.scala 71:109:@23557.4]
  wire [11:0] _T_71437; // @[Modules.scala 71:109:@23559.4]
  wire [10:0] _T_71438; // @[Modules.scala 71:109:@23560.4]
  wire [10:0] buffer_9_732; // @[Modules.scala 71:109:@23561.4]
  wire [11:0] _T_71440; // @[Modules.scala 71:109:@23563.4]
  wire [10:0] _T_71441; // @[Modules.scala 71:109:@23564.4]
  wire [10:0] buffer_9_733; // @[Modules.scala 71:109:@23565.4]
  wire [11:0] _T_71443; // @[Modules.scala 71:109:@23567.4]
  wire [10:0] _T_71444; // @[Modules.scala 71:109:@23568.4]
  wire [10:0] buffer_9_734; // @[Modules.scala 71:109:@23569.4]
  wire [11:0] _T_71446; // @[Modules.scala 78:156:@23572.4]
  wire [10:0] _T_71447; // @[Modules.scala 78:156:@23573.4]
  wire [10:0] buffer_9_736; // @[Modules.scala 78:156:@23574.4]
  wire [11:0] _T_71449; // @[Modules.scala 78:156:@23576.4]
  wire [10:0] _T_71450; // @[Modules.scala 78:156:@23577.4]
  wire [10:0] buffer_9_737; // @[Modules.scala 78:156:@23578.4]
  wire [11:0] _T_71452; // @[Modules.scala 78:156:@23580.4]
  wire [10:0] _T_71453; // @[Modules.scala 78:156:@23581.4]
  wire [10:0] buffer_9_738; // @[Modules.scala 78:156:@23582.4]
  wire [11:0] _T_71455; // @[Modules.scala 78:156:@23584.4]
  wire [10:0] _T_71456; // @[Modules.scala 78:156:@23585.4]
  wire [10:0] buffer_9_739; // @[Modules.scala 78:156:@23586.4]
  wire [11:0] _T_71458; // @[Modules.scala 78:156:@23588.4]
  wire [10:0] _T_71459; // @[Modules.scala 78:156:@23589.4]
  wire [10:0] buffer_9_740; // @[Modules.scala 78:156:@23590.4]
  wire [11:0] _T_71461; // @[Modules.scala 78:156:@23592.4]
  wire [10:0] _T_71462; // @[Modules.scala 78:156:@23593.4]
  wire [10:0] buffer_9_741; // @[Modules.scala 78:156:@23594.4]
  wire [11:0] _T_71464; // @[Modules.scala 78:156:@23596.4]
  wire [10:0] _T_71465; // @[Modules.scala 78:156:@23597.4]
  wire [10:0] buffer_9_742; // @[Modules.scala 78:156:@23598.4]
  wire [11:0] _T_71467; // @[Modules.scala 78:156:@23600.4]
  wire [10:0] _T_71468; // @[Modules.scala 78:156:@23601.4]
  wire [10:0] buffer_9_743; // @[Modules.scala 78:156:@23602.4]
  wire [11:0] _T_71470; // @[Modules.scala 78:156:@23604.4]
  wire [10:0] _T_71471; // @[Modules.scala 78:156:@23605.4]
  wire [10:0] buffer_9_744; // @[Modules.scala 78:156:@23606.4]
  wire [11:0] _T_71473; // @[Modules.scala 78:156:@23608.4]
  wire [10:0] _T_71474; // @[Modules.scala 78:156:@23609.4]
  wire [10:0] buffer_9_745; // @[Modules.scala 78:156:@23610.4]
  wire [11:0] _T_71476; // @[Modules.scala 78:156:@23612.4]
  wire [10:0] _T_71477; // @[Modules.scala 78:156:@23613.4]
  wire [10:0] buffer_9_746; // @[Modules.scala 78:156:@23614.4]
  wire [11:0] _T_71479; // @[Modules.scala 78:156:@23616.4]
  wire [10:0] _T_71480; // @[Modules.scala 78:156:@23617.4]
  wire [10:0] buffer_9_747; // @[Modules.scala 78:156:@23618.4]
  wire [11:0] _T_71482; // @[Modules.scala 78:156:@23620.4]
  wire [10:0] _T_71483; // @[Modules.scala 78:156:@23621.4]
  wire [10:0] buffer_9_748; // @[Modules.scala 78:156:@23622.4]
  wire [11:0] _T_71485; // @[Modules.scala 78:156:@23624.4]
  wire [10:0] _T_71486; // @[Modules.scala 78:156:@23625.4]
  wire [10:0] buffer_9_749; // @[Modules.scala 78:156:@23626.4]
  wire [11:0] _T_71488; // @[Modules.scala 78:156:@23628.4]
  wire [10:0] _T_71489; // @[Modules.scala 78:156:@23629.4]
  wire [10:0] buffer_9_750; // @[Modules.scala 78:156:@23630.4]
  wire [11:0] _T_71491; // @[Modules.scala 78:156:@23632.4]
  wire [10:0] _T_71492; // @[Modules.scala 78:156:@23633.4]
  wire [10:0] buffer_9_751; // @[Modules.scala 78:156:@23634.4]
  wire [11:0] _T_71494; // @[Modules.scala 78:156:@23636.4]
  wire [10:0] _T_71495; // @[Modules.scala 78:156:@23637.4]
  wire [10:0] buffer_9_752; // @[Modules.scala 78:156:@23638.4]
  wire [11:0] _T_71497; // @[Modules.scala 78:156:@23640.4]
  wire [10:0] _T_71498; // @[Modules.scala 78:156:@23641.4]
  wire [10:0] buffer_9_753; // @[Modules.scala 78:156:@23642.4]
  wire [11:0] _T_71500; // @[Modules.scala 78:156:@23644.4]
  wire [10:0] _T_71501; // @[Modules.scala 78:156:@23645.4]
  wire [10:0] buffer_9_754; // @[Modules.scala 78:156:@23646.4]
  wire [11:0] _T_71503; // @[Modules.scala 78:156:@23648.4]
  wire [10:0] _T_71504; // @[Modules.scala 78:156:@23649.4]
  wire [10:0] buffer_9_755; // @[Modules.scala 78:156:@23650.4]
  wire [11:0] _T_71506; // @[Modules.scala 78:156:@23652.4]
  wire [10:0] _T_71507; // @[Modules.scala 78:156:@23653.4]
  wire [10:0] buffer_9_756; // @[Modules.scala 78:156:@23654.4]
  wire [11:0] _T_71509; // @[Modules.scala 78:156:@23656.4]
  wire [10:0] _T_71510; // @[Modules.scala 78:156:@23657.4]
  wire [10:0] buffer_9_757; // @[Modules.scala 78:156:@23658.4]
  wire [11:0] _T_71512; // @[Modules.scala 78:156:@23660.4]
  wire [10:0] _T_71513; // @[Modules.scala 78:156:@23661.4]
  wire [10:0] buffer_9_758; // @[Modules.scala 78:156:@23662.4]
  wire [11:0] _T_71515; // @[Modules.scala 78:156:@23664.4]
  wire [10:0] _T_71516; // @[Modules.scala 78:156:@23665.4]
  wire [10:0] buffer_9_759; // @[Modules.scala 78:156:@23666.4]
  wire [11:0] _T_71518; // @[Modules.scala 78:156:@23668.4]
  wire [10:0] _T_71519; // @[Modules.scala 78:156:@23669.4]
  wire [10:0] buffer_9_760; // @[Modules.scala 78:156:@23670.4]
  wire [11:0] _T_71521; // @[Modules.scala 78:156:@23672.4]
  wire [10:0] _T_71522; // @[Modules.scala 78:156:@23673.4]
  wire [10:0] buffer_9_761; // @[Modules.scala 78:156:@23674.4]
  wire [11:0] _T_71524; // @[Modules.scala 78:156:@23676.4]
  wire [10:0] _T_71525; // @[Modules.scala 78:156:@23677.4]
  wire [10:0] buffer_9_762; // @[Modules.scala 78:156:@23678.4]
  wire [11:0] _T_71527; // @[Modules.scala 78:156:@23680.4]
  wire [10:0] _T_71528; // @[Modules.scala 78:156:@23681.4]
  wire [10:0] buffer_9_763; // @[Modules.scala 78:156:@23682.4]
  wire [11:0] _T_71530; // @[Modules.scala 78:156:@23684.4]
  wire [10:0] _T_71531; // @[Modules.scala 78:156:@23685.4]
  wire [10:0] buffer_9_764; // @[Modules.scala 78:156:@23686.4]
  wire [11:0] _T_71533; // @[Modules.scala 78:156:@23688.4]
  wire [10:0] _T_71534; // @[Modules.scala 78:156:@23689.4]
  wire [10:0] buffer_9_765; // @[Modules.scala 78:156:@23690.4]
  wire [11:0] _T_71536; // @[Modules.scala 78:156:@23692.4]
  wire [10:0] _T_71537; // @[Modules.scala 78:156:@23693.4]
  wire [10:0] buffer_9_766; // @[Modules.scala 78:156:@23694.4]
  wire [11:0] _T_71539; // @[Modules.scala 78:156:@23696.4]
  wire [10:0] _T_71540; // @[Modules.scala 78:156:@23697.4]
  wire [10:0] buffer_9_767; // @[Modules.scala 78:156:@23698.4]
  wire [11:0] _T_71542; // @[Modules.scala 78:156:@23700.4]
  wire [10:0] _T_71543; // @[Modules.scala 78:156:@23701.4]
  wire [10:0] buffer_9_768; // @[Modules.scala 78:156:@23702.4]
  wire [11:0] _T_71545; // @[Modules.scala 78:156:@23704.4]
  wire [10:0] _T_71546; // @[Modules.scala 78:156:@23705.4]
  wire [10:0] buffer_9_769; // @[Modules.scala 78:156:@23706.4]
  wire [11:0] _T_71548; // @[Modules.scala 78:156:@23708.4]
  wire [10:0] _T_71549; // @[Modules.scala 78:156:@23709.4]
  wire [10:0] buffer_9_770; // @[Modules.scala 78:156:@23710.4]
  wire [11:0] _T_71551; // @[Modules.scala 78:156:@23712.4]
  wire [10:0] _T_71552; // @[Modules.scala 78:156:@23713.4]
  wire [10:0] buffer_9_771; // @[Modules.scala 78:156:@23714.4]
  wire [11:0] _T_71554; // @[Modules.scala 78:156:@23716.4]
  wire [10:0] _T_71555; // @[Modules.scala 78:156:@23717.4]
  wire [10:0] buffer_9_772; // @[Modules.scala 78:156:@23718.4]
  wire [11:0] _T_71557; // @[Modules.scala 78:156:@23720.4]
  wire [10:0] _T_71558; // @[Modules.scala 78:156:@23721.4]
  wire [10:0] buffer_9_773; // @[Modules.scala 78:156:@23722.4]
  wire [11:0] _T_71560; // @[Modules.scala 78:156:@23724.4]
  wire [10:0] _T_71561; // @[Modules.scala 78:156:@23725.4]
  wire [10:0] buffer_9_774; // @[Modules.scala 78:156:@23726.4]
  wire [11:0] _T_71563; // @[Modules.scala 78:156:@23728.4]
  wire [10:0] _T_71564; // @[Modules.scala 78:156:@23729.4]
  wire [10:0] buffer_9_775; // @[Modules.scala 78:156:@23730.4]
  wire [11:0] _T_71566; // @[Modules.scala 78:156:@23732.4]
  wire [10:0] _T_71567; // @[Modules.scala 78:156:@23733.4]
  wire [10:0] buffer_9_776; // @[Modules.scala 78:156:@23734.4]
  wire [11:0] _T_71569; // @[Modules.scala 78:156:@23736.4]
  wire [10:0] _T_71570; // @[Modules.scala 78:156:@23737.4]
  wire [10:0] buffer_9_777; // @[Modules.scala 78:156:@23738.4]
  wire [11:0] _T_71572; // @[Modules.scala 78:156:@23740.4]
  wire [10:0] _T_71573; // @[Modules.scala 78:156:@23741.4]
  wire [10:0] buffer_9_778; // @[Modules.scala 78:156:@23742.4]
  wire [11:0] _T_71575; // @[Modules.scala 78:156:@23744.4]
  wire [10:0] _T_71576; // @[Modules.scala 78:156:@23745.4]
  wire [10:0] buffer_9_779; // @[Modules.scala 78:156:@23746.4]
  wire [11:0] _T_71578; // @[Modules.scala 78:156:@23748.4]
  wire [10:0] _T_71579; // @[Modules.scala 78:156:@23749.4]
  wire [10:0] buffer_9_780; // @[Modules.scala 78:156:@23750.4]
  wire [11:0] _T_71581; // @[Modules.scala 78:156:@23752.4]
  wire [10:0] _T_71582; // @[Modules.scala 78:156:@23753.4]
  wire [10:0] buffer_9_781; // @[Modules.scala 78:156:@23754.4]
  wire [11:0] _T_71584; // @[Modules.scala 78:156:@23756.4]
  wire [10:0] _T_71585; // @[Modules.scala 78:156:@23757.4]
  wire [10:0] buffer_9_782; // @[Modules.scala 78:156:@23758.4]
  wire [11:0] _T_71587; // @[Modules.scala 78:156:@23760.4]
  wire [10:0] _T_71588; // @[Modules.scala 78:156:@23761.4]
  wire [10:0] buffer_9_783; // @[Modules.scala 78:156:@23762.4]
  wire [5:0] _T_71705; // @[Modules.scala 37:46:@23929.4]
  wire [4:0] _T_71706; // @[Modules.scala 37:46:@23930.4]
  wire [4:0] _T_71707; // @[Modules.scala 37:46:@23931.4]
  wire [5:0] _T_71839; // @[Modules.scala 37:46:@24117.4]
  wire [4:0] _T_71840; // @[Modules.scala 37:46:@24118.4]
  wire [4:0] _T_71841; // @[Modules.scala 37:46:@24119.4]
  wire [5:0] _T_72129; // @[Modules.scala 37:46:@24534.4]
  wire [4:0] _T_72130; // @[Modules.scala 37:46:@24535.4]
  wire [4:0] _T_72131; // @[Modules.scala 37:46:@24536.4]
  wire [11:0] _T_72240; // @[Modules.scala 65:57:@24686.4]
  wire [10:0] _T_72241; // @[Modules.scala 65:57:@24687.4]
  wire [10:0] buffer_10_393; // @[Modules.scala 65:57:@24688.4]
  wire [11:0] _T_72243; // @[Modules.scala 65:57:@24690.4]
  wire [10:0] _T_72244; // @[Modules.scala 65:57:@24691.4]
  wire [10:0] buffer_10_394; // @[Modules.scala 65:57:@24692.4]
  wire [11:0] _T_72255; // @[Modules.scala 65:57:@24706.4]
  wire [10:0] _T_72256; // @[Modules.scala 65:57:@24707.4]
  wire [10:0] buffer_10_398; // @[Modules.scala 65:57:@24708.4]
  wire [11:0] _T_72276; // @[Modules.scala 65:57:@24734.4]
  wire [10:0] _T_72277; // @[Modules.scala 65:57:@24735.4]
  wire [10:0] buffer_10_405; // @[Modules.scala 65:57:@24736.4]
  wire [11:0] _T_72282; // @[Modules.scala 65:57:@24742.4]
  wire [10:0] _T_72283; // @[Modules.scala 65:57:@24743.4]
  wire [10:0] buffer_10_407; // @[Modules.scala 65:57:@24744.4]
  wire [11:0] _T_72300; // @[Modules.scala 65:57:@24766.4]
  wire [10:0] _T_72301; // @[Modules.scala 65:57:@24767.4]
  wire [10:0] buffer_10_413; // @[Modules.scala 65:57:@24768.4]
  wire [11:0] _T_72318; // @[Modules.scala 65:57:@24790.4]
  wire [10:0] _T_72319; // @[Modules.scala 65:57:@24791.4]
  wire [10:0] buffer_10_419; // @[Modules.scala 65:57:@24792.4]
  wire [10:0] buffer_10_56; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72321; // @[Modules.scala 65:57:@24794.4]
  wire [10:0] _T_72322; // @[Modules.scala 65:57:@24795.4]
  wire [10:0] buffer_10_420; // @[Modules.scala 65:57:@24796.4]
  wire [11:0] _T_72333; // @[Modules.scala 65:57:@24810.4]
  wire [10:0] _T_72334; // @[Modules.scala 65:57:@24811.4]
  wire [10:0] buffer_10_424; // @[Modules.scala 65:57:@24812.4]
  wire [11:0] _T_72339; // @[Modules.scala 65:57:@24818.4]
  wire [10:0] _T_72340; // @[Modules.scala 65:57:@24819.4]
  wire [10:0] buffer_10_426; // @[Modules.scala 65:57:@24820.4]
  wire [11:0] _T_72342; // @[Modules.scala 65:57:@24822.4]
  wire [10:0] _T_72343; // @[Modules.scala 65:57:@24823.4]
  wire [10:0] buffer_10_427; // @[Modules.scala 65:57:@24824.4]
  wire [11:0] _T_72348; // @[Modules.scala 65:57:@24830.4]
  wire [10:0] _T_72349; // @[Modules.scala 65:57:@24831.4]
  wire [10:0] buffer_10_429; // @[Modules.scala 65:57:@24832.4]
  wire [10:0] buffer_10_77; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72351; // @[Modules.scala 65:57:@24834.4]
  wire [10:0] _T_72352; // @[Modules.scala 65:57:@24835.4]
  wire [10:0] buffer_10_430; // @[Modules.scala 65:57:@24836.4]
  wire [11:0] _T_72354; // @[Modules.scala 65:57:@24838.4]
  wire [10:0] _T_72355; // @[Modules.scala 65:57:@24839.4]
  wire [10:0] buffer_10_431; // @[Modules.scala 65:57:@24840.4]
  wire [11:0] _T_72357; // @[Modules.scala 65:57:@24842.4]
  wire [10:0] _T_72358; // @[Modules.scala 65:57:@24843.4]
  wire [10:0] buffer_10_432; // @[Modules.scala 65:57:@24844.4]
  wire [11:0] _T_72360; // @[Modules.scala 65:57:@24846.4]
  wire [10:0] _T_72361; // @[Modules.scala 65:57:@24847.4]
  wire [10:0] buffer_10_433; // @[Modules.scala 65:57:@24848.4]
  wire [11:0] _T_72363; // @[Modules.scala 65:57:@24850.4]
  wire [10:0] _T_72364; // @[Modules.scala 65:57:@24851.4]
  wire [10:0] buffer_10_434; // @[Modules.scala 65:57:@24852.4]
  wire [11:0] _T_72366; // @[Modules.scala 65:57:@24854.4]
  wire [10:0] _T_72367; // @[Modules.scala 65:57:@24855.4]
  wire [10:0] buffer_10_435; // @[Modules.scala 65:57:@24856.4]
  wire [10:0] buffer_10_88; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72369; // @[Modules.scala 65:57:@24858.4]
  wire [10:0] _T_72370; // @[Modules.scala 65:57:@24859.4]
  wire [10:0] buffer_10_436; // @[Modules.scala 65:57:@24860.4]
  wire [11:0] _T_72381; // @[Modules.scala 65:57:@24874.4]
  wire [10:0] _T_72382; // @[Modules.scala 65:57:@24875.4]
  wire [10:0] buffer_10_440; // @[Modules.scala 65:57:@24876.4]
  wire [10:0] buffer_10_100; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72387; // @[Modules.scala 65:57:@24882.4]
  wire [10:0] _T_72388; // @[Modules.scala 65:57:@24883.4]
  wire [10:0] buffer_10_442; // @[Modules.scala 65:57:@24884.4]
  wire [11:0] _T_72390; // @[Modules.scala 65:57:@24886.4]
  wire [10:0] _T_72391; // @[Modules.scala 65:57:@24887.4]
  wire [10:0] buffer_10_443; // @[Modules.scala 65:57:@24888.4]
  wire [11:0] _T_72393; // @[Modules.scala 65:57:@24890.4]
  wire [10:0] _T_72394; // @[Modules.scala 65:57:@24891.4]
  wire [10:0] buffer_10_444; // @[Modules.scala 65:57:@24892.4]
  wire [11:0] _T_72408; // @[Modules.scala 65:57:@24910.4]
  wire [10:0] _T_72409; // @[Modules.scala 65:57:@24911.4]
  wire [10:0] buffer_10_449; // @[Modules.scala 65:57:@24912.4]
  wire [10:0] buffer_10_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72414; // @[Modules.scala 65:57:@24918.4]
  wire [10:0] _T_72415; // @[Modules.scala 65:57:@24919.4]
  wire [10:0] buffer_10_451; // @[Modules.scala 65:57:@24920.4]
  wire [10:0] buffer_10_154; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72468; // @[Modules.scala 65:57:@24990.4]
  wire [10:0] _T_72469; // @[Modules.scala 65:57:@24991.4]
  wire [10:0] buffer_10_469; // @[Modules.scala 65:57:@24992.4]
  wire [11:0] _T_72480; // @[Modules.scala 65:57:@25006.4]
  wire [10:0] _T_72481; // @[Modules.scala 65:57:@25007.4]
  wire [10:0] buffer_10_473; // @[Modules.scala 65:57:@25008.4]
  wire [11:0] _T_72486; // @[Modules.scala 65:57:@25014.4]
  wire [10:0] _T_72487; // @[Modules.scala 65:57:@25015.4]
  wire [10:0] buffer_10_475; // @[Modules.scala 65:57:@25016.4]
  wire [11:0] _T_72501; // @[Modules.scala 65:57:@25034.4]
  wire [10:0] _T_72502; // @[Modules.scala 65:57:@25035.4]
  wire [10:0] buffer_10_480; // @[Modules.scala 65:57:@25036.4]
  wire [11:0] _T_72522; // @[Modules.scala 65:57:@25062.4]
  wire [10:0] _T_72523; // @[Modules.scala 65:57:@25063.4]
  wire [10:0] buffer_10_487; // @[Modules.scala 65:57:@25064.4]
  wire [10:0] buffer_10_193; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72525; // @[Modules.scala 65:57:@25066.4]
  wire [10:0] _T_72526; // @[Modules.scala 65:57:@25067.4]
  wire [10:0] buffer_10_488; // @[Modules.scala 65:57:@25068.4]
  wire [10:0] buffer_10_203; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72540; // @[Modules.scala 65:57:@25086.4]
  wire [10:0] _T_72541; // @[Modules.scala 65:57:@25087.4]
  wire [10:0] buffer_10_493; // @[Modules.scala 65:57:@25088.4]
  wire [11:0] _T_72546; // @[Modules.scala 65:57:@25094.4]
  wire [10:0] _T_72547; // @[Modules.scala 65:57:@25095.4]
  wire [10:0] buffer_10_495; // @[Modules.scala 65:57:@25096.4]
  wire [11:0] _T_72549; // @[Modules.scala 65:57:@25098.4]
  wire [10:0] _T_72550; // @[Modules.scala 65:57:@25099.4]
  wire [10:0] buffer_10_496; // @[Modules.scala 65:57:@25100.4]
  wire [11:0] _T_72567; // @[Modules.scala 65:57:@25122.4]
  wire [10:0] _T_72568; // @[Modules.scala 65:57:@25123.4]
  wire [10:0] buffer_10_502; // @[Modules.scala 65:57:@25124.4]
  wire [11:0] _T_72576; // @[Modules.scala 65:57:@25134.4]
  wire [10:0] _T_72577; // @[Modules.scala 65:57:@25135.4]
  wire [10:0] buffer_10_505; // @[Modules.scala 65:57:@25136.4]
  wire [10:0] buffer_10_230; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72582; // @[Modules.scala 65:57:@25142.4]
  wire [10:0] _T_72583; // @[Modules.scala 65:57:@25143.4]
  wire [10:0] buffer_10_507; // @[Modules.scala 65:57:@25144.4]
  wire [11:0] _T_72588; // @[Modules.scala 65:57:@25150.4]
  wire [10:0] _T_72589; // @[Modules.scala 65:57:@25151.4]
  wire [10:0] buffer_10_509; // @[Modules.scala 65:57:@25152.4]
  wire [11:0] _T_72603; // @[Modules.scala 65:57:@25170.4]
  wire [10:0] _T_72604; // @[Modules.scala 65:57:@25171.4]
  wire [10:0] buffer_10_514; // @[Modules.scala 65:57:@25172.4]
  wire [11:0] _T_72606; // @[Modules.scala 65:57:@25174.4]
  wire [10:0] _T_72607; // @[Modules.scala 65:57:@25175.4]
  wire [10:0] buffer_10_515; // @[Modules.scala 65:57:@25176.4]
  wire [10:0] buffer_10_255; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72618; // @[Modules.scala 65:57:@25190.4]
  wire [10:0] _T_72619; // @[Modules.scala 65:57:@25191.4]
  wire [10:0] buffer_10_519; // @[Modules.scala 65:57:@25192.4]
  wire [11:0] _T_72621; // @[Modules.scala 65:57:@25194.4]
  wire [10:0] _T_72622; // @[Modules.scala 65:57:@25195.4]
  wire [10:0] buffer_10_520; // @[Modules.scala 65:57:@25196.4]
  wire [11:0] _T_72624; // @[Modules.scala 65:57:@25198.4]
  wire [10:0] _T_72625; // @[Modules.scala 65:57:@25199.4]
  wire [10:0] buffer_10_521; // @[Modules.scala 65:57:@25200.4]
  wire [11:0] _T_72642; // @[Modules.scala 65:57:@25222.4]
  wire [10:0] _T_72643; // @[Modules.scala 65:57:@25223.4]
  wire [10:0] buffer_10_527; // @[Modules.scala 65:57:@25224.4]
  wire [11:0] _T_72663; // @[Modules.scala 65:57:@25250.4]
  wire [10:0] _T_72664; // @[Modules.scala 65:57:@25251.4]
  wire [10:0] buffer_10_534; // @[Modules.scala 65:57:@25252.4]
  wire [11:0] _T_72672; // @[Modules.scala 65:57:@25262.4]
  wire [10:0] _T_72673; // @[Modules.scala 65:57:@25263.4]
  wire [10:0] buffer_10_537; // @[Modules.scala 65:57:@25264.4]
  wire [11:0] _T_72693; // @[Modules.scala 65:57:@25290.4]
  wire [10:0] _T_72694; // @[Modules.scala 65:57:@25291.4]
  wire [10:0] buffer_10_544; // @[Modules.scala 65:57:@25292.4]
  wire [11:0] _T_72696; // @[Modules.scala 65:57:@25294.4]
  wire [10:0] _T_72697; // @[Modules.scala 65:57:@25295.4]
  wire [10:0] buffer_10_545; // @[Modules.scala 65:57:@25296.4]
  wire [10:0] buffer_10_318; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72714; // @[Modules.scala 65:57:@25318.4]
  wire [10:0] _T_72715; // @[Modules.scala 65:57:@25319.4]
  wire [10:0] buffer_10_551; // @[Modules.scala 65:57:@25320.4]
  wire [11:0] _T_72717; // @[Modules.scala 65:57:@25322.4]
  wire [10:0] _T_72718; // @[Modules.scala 65:57:@25323.4]
  wire [10:0] buffer_10_552; // @[Modules.scala 65:57:@25324.4]
  wire [10:0] buffer_10_322; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72720; // @[Modules.scala 65:57:@25326.4]
  wire [10:0] _T_72721; // @[Modules.scala 65:57:@25327.4]
  wire [10:0] buffer_10_553; // @[Modules.scala 65:57:@25328.4]
  wire [11:0] _T_72726; // @[Modules.scala 65:57:@25334.4]
  wire [10:0] _T_72727; // @[Modules.scala 65:57:@25335.4]
  wire [10:0] buffer_10_555; // @[Modules.scala 65:57:@25336.4]
  wire [11:0] _T_72750; // @[Modules.scala 65:57:@25366.4]
  wire [10:0] _T_72751; // @[Modules.scala 65:57:@25367.4]
  wire [10:0] buffer_10_563; // @[Modules.scala 65:57:@25368.4]
  wire [10:0] buffer_10_353; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72765; // @[Modules.scala 65:57:@25386.4]
  wire [10:0] _T_72766; // @[Modules.scala 65:57:@25387.4]
  wire [10:0] buffer_10_568; // @[Modules.scala 65:57:@25388.4]
  wire [10:0] buffer_10_368; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_72789; // @[Modules.scala 65:57:@25418.4]
  wire [10:0] _T_72790; // @[Modules.scala 65:57:@25419.4]
  wire [10:0] buffer_10_576; // @[Modules.scala 65:57:@25420.4]
  wire [11:0] _T_72801; // @[Modules.scala 65:57:@25434.4]
  wire [10:0] _T_72802; // @[Modules.scala 65:57:@25435.4]
  wire [10:0] buffer_10_580; // @[Modules.scala 65:57:@25436.4]
  wire [11:0] _T_72804; // @[Modules.scala 65:57:@25438.4]
  wire [10:0] _T_72805; // @[Modules.scala 65:57:@25439.4]
  wire [10:0] buffer_10_581; // @[Modules.scala 65:57:@25440.4]
  wire [11:0] _T_72807; // @[Modules.scala 65:57:@25442.4]
  wire [10:0] _T_72808; // @[Modules.scala 65:57:@25443.4]
  wire [10:0] buffer_10_582; // @[Modules.scala 65:57:@25444.4]
  wire [11:0] _T_72822; // @[Modules.scala 65:57:@25462.4]
  wire [10:0] _T_72823; // @[Modules.scala 65:57:@25463.4]
  wire [10:0] buffer_10_587; // @[Modules.scala 65:57:@25464.4]
  wire [11:0] _T_72825; // @[Modules.scala 68:83:@25466.4]
  wire [10:0] _T_72826; // @[Modules.scala 68:83:@25467.4]
  wire [10:0] buffer_10_588; // @[Modules.scala 68:83:@25468.4]
  wire [11:0] _T_72828; // @[Modules.scala 68:83:@25470.4]
  wire [10:0] _T_72829; // @[Modules.scala 68:83:@25471.4]
  wire [10:0] buffer_10_589; // @[Modules.scala 68:83:@25472.4]
  wire [11:0] _T_72834; // @[Modules.scala 68:83:@25478.4]
  wire [10:0] _T_72835; // @[Modules.scala 68:83:@25479.4]
  wire [10:0] buffer_10_591; // @[Modules.scala 68:83:@25480.4]
  wire [11:0] _T_72843; // @[Modules.scala 68:83:@25490.4]
  wire [10:0] _T_72844; // @[Modules.scala 68:83:@25491.4]
  wire [10:0] buffer_10_594; // @[Modules.scala 68:83:@25492.4]
  wire [11:0] _T_72846; // @[Modules.scala 68:83:@25494.4]
  wire [10:0] _T_72847; // @[Modules.scala 68:83:@25495.4]
  wire [10:0] buffer_10_595; // @[Modules.scala 68:83:@25496.4]
  wire [11:0] _T_72855; // @[Modules.scala 68:83:@25506.4]
  wire [10:0] _T_72856; // @[Modules.scala 68:83:@25507.4]
  wire [10:0] buffer_10_598; // @[Modules.scala 68:83:@25508.4]
  wire [11:0] _T_72864; // @[Modules.scala 68:83:@25518.4]
  wire [10:0] _T_72865; // @[Modules.scala 68:83:@25519.4]
  wire [10:0] buffer_10_601; // @[Modules.scala 68:83:@25520.4]
  wire [11:0] _T_72867; // @[Modules.scala 68:83:@25522.4]
  wire [10:0] _T_72868; // @[Modules.scala 68:83:@25523.4]
  wire [10:0] buffer_10_602; // @[Modules.scala 68:83:@25524.4]
  wire [11:0] _T_72870; // @[Modules.scala 68:83:@25526.4]
  wire [10:0] _T_72871; // @[Modules.scala 68:83:@25527.4]
  wire [10:0] buffer_10_603; // @[Modules.scala 68:83:@25528.4]
  wire [11:0] _T_72873; // @[Modules.scala 68:83:@25530.4]
  wire [10:0] _T_72874; // @[Modules.scala 68:83:@25531.4]
  wire [10:0] buffer_10_604; // @[Modules.scala 68:83:@25532.4]
  wire [11:0] _T_72876; // @[Modules.scala 68:83:@25534.4]
  wire [10:0] _T_72877; // @[Modules.scala 68:83:@25535.4]
  wire [10:0] buffer_10_605; // @[Modules.scala 68:83:@25536.4]
  wire [11:0] _T_72879; // @[Modules.scala 68:83:@25538.4]
  wire [10:0] _T_72880; // @[Modules.scala 68:83:@25539.4]
  wire [10:0] buffer_10_606; // @[Modules.scala 68:83:@25540.4]
  wire [11:0] _T_72882; // @[Modules.scala 68:83:@25542.4]
  wire [10:0] _T_72883; // @[Modules.scala 68:83:@25543.4]
  wire [10:0] buffer_10_607; // @[Modules.scala 68:83:@25544.4]
  wire [11:0] _T_72885; // @[Modules.scala 68:83:@25546.4]
  wire [10:0] _T_72886; // @[Modules.scala 68:83:@25547.4]
  wire [10:0] buffer_10_608; // @[Modules.scala 68:83:@25548.4]
  wire [11:0] _T_72888; // @[Modules.scala 68:83:@25550.4]
  wire [10:0] _T_72889; // @[Modules.scala 68:83:@25551.4]
  wire [10:0] buffer_10_609; // @[Modules.scala 68:83:@25552.4]
  wire [11:0] _T_72891; // @[Modules.scala 68:83:@25554.4]
  wire [10:0] _T_72892; // @[Modules.scala 68:83:@25555.4]
  wire [10:0] buffer_10_610; // @[Modules.scala 68:83:@25556.4]
  wire [11:0] _T_72897; // @[Modules.scala 68:83:@25562.4]
  wire [10:0] _T_72898; // @[Modules.scala 68:83:@25563.4]
  wire [10:0] buffer_10_612; // @[Modules.scala 68:83:@25564.4]
  wire [11:0] _T_72900; // @[Modules.scala 68:83:@25566.4]
  wire [10:0] _T_72901; // @[Modules.scala 68:83:@25567.4]
  wire [10:0] buffer_10_613; // @[Modules.scala 68:83:@25568.4]
  wire [11:0] _T_72903; // @[Modules.scala 68:83:@25570.4]
  wire [10:0] _T_72904; // @[Modules.scala 68:83:@25571.4]
  wire [10:0] buffer_10_614; // @[Modules.scala 68:83:@25572.4]
  wire [11:0] _T_72906; // @[Modules.scala 68:83:@25574.4]
  wire [10:0] _T_72907; // @[Modules.scala 68:83:@25575.4]
  wire [10:0] buffer_10_615; // @[Modules.scala 68:83:@25576.4]
  wire [11:0] _T_72909; // @[Modules.scala 68:83:@25578.4]
  wire [10:0] _T_72910; // @[Modules.scala 68:83:@25579.4]
  wire [10:0] buffer_10_616; // @[Modules.scala 68:83:@25580.4]
  wire [11:0] _T_72912; // @[Modules.scala 68:83:@25582.4]
  wire [10:0] _T_72913; // @[Modules.scala 68:83:@25583.4]
  wire [10:0] buffer_10_617; // @[Modules.scala 68:83:@25584.4]
  wire [11:0] _T_72918; // @[Modules.scala 68:83:@25590.4]
  wire [10:0] _T_72919; // @[Modules.scala 68:83:@25591.4]
  wire [10:0] buffer_10_619; // @[Modules.scala 68:83:@25592.4]
  wire [11:0] _T_72921; // @[Modules.scala 68:83:@25594.4]
  wire [10:0] _T_72922; // @[Modules.scala 68:83:@25595.4]
  wire [10:0] buffer_10_620; // @[Modules.scala 68:83:@25596.4]
  wire [11:0] _T_72930; // @[Modules.scala 68:83:@25606.4]
  wire [10:0] _T_72931; // @[Modules.scala 68:83:@25607.4]
  wire [10:0] buffer_10_623; // @[Modules.scala 68:83:@25608.4]
  wire [11:0] _T_72939; // @[Modules.scala 68:83:@25618.4]
  wire [10:0] _T_72940; // @[Modules.scala 68:83:@25619.4]
  wire [10:0] buffer_10_626; // @[Modules.scala 68:83:@25620.4]
  wire [11:0] _T_72945; // @[Modules.scala 68:83:@25626.4]
  wire [10:0] _T_72946; // @[Modules.scala 68:83:@25627.4]
  wire [10:0] buffer_10_628; // @[Modules.scala 68:83:@25628.4]
  wire [11:0] _T_72948; // @[Modules.scala 68:83:@25630.4]
  wire [10:0] _T_72949; // @[Modules.scala 68:83:@25631.4]
  wire [10:0] buffer_10_629; // @[Modules.scala 68:83:@25632.4]
  wire [11:0] _T_72957; // @[Modules.scala 68:83:@25642.4]
  wire [10:0] _T_72958; // @[Modules.scala 68:83:@25643.4]
  wire [10:0] buffer_10_632; // @[Modules.scala 68:83:@25644.4]
  wire [11:0] _T_72960; // @[Modules.scala 68:83:@25646.4]
  wire [10:0] _T_72961; // @[Modules.scala 68:83:@25647.4]
  wire [10:0] buffer_10_633; // @[Modules.scala 68:83:@25648.4]
  wire [11:0] _T_72966; // @[Modules.scala 68:83:@25654.4]
  wire [10:0] _T_72967; // @[Modules.scala 68:83:@25655.4]
  wire [10:0] buffer_10_635; // @[Modules.scala 68:83:@25656.4]
  wire [11:0] _T_72969; // @[Modules.scala 68:83:@25658.4]
  wire [10:0] _T_72970; // @[Modules.scala 68:83:@25659.4]
  wire [10:0] buffer_10_636; // @[Modules.scala 68:83:@25660.4]
  wire [11:0] _T_72972; // @[Modules.scala 68:83:@25662.4]
  wire [10:0] _T_72973; // @[Modules.scala 68:83:@25663.4]
  wire [10:0] buffer_10_637; // @[Modules.scala 68:83:@25664.4]
  wire [11:0] _T_72975; // @[Modules.scala 68:83:@25666.4]
  wire [10:0] _T_72976; // @[Modules.scala 68:83:@25667.4]
  wire [10:0] buffer_10_638; // @[Modules.scala 68:83:@25668.4]
  wire [11:0] _T_72978; // @[Modules.scala 68:83:@25670.4]
  wire [10:0] _T_72979; // @[Modules.scala 68:83:@25671.4]
  wire [10:0] buffer_10_639; // @[Modules.scala 68:83:@25672.4]
  wire [11:0] _T_72981; // @[Modules.scala 68:83:@25674.4]
  wire [10:0] _T_72982; // @[Modules.scala 68:83:@25675.4]
  wire [10:0] buffer_10_640; // @[Modules.scala 68:83:@25676.4]
  wire [11:0] _T_72987; // @[Modules.scala 68:83:@25682.4]
  wire [10:0] _T_72988; // @[Modules.scala 68:83:@25683.4]
  wire [10:0] buffer_10_642; // @[Modules.scala 68:83:@25684.4]
  wire [11:0] _T_72990; // @[Modules.scala 68:83:@25686.4]
  wire [10:0] _T_72991; // @[Modules.scala 68:83:@25687.4]
  wire [10:0] buffer_10_643; // @[Modules.scala 68:83:@25688.4]
  wire [11:0] _T_72993; // @[Modules.scala 68:83:@25690.4]
  wire [10:0] _T_72994; // @[Modules.scala 68:83:@25691.4]
  wire [10:0] buffer_10_644; // @[Modules.scala 68:83:@25692.4]
  wire [11:0] _T_72996; // @[Modules.scala 68:83:@25694.4]
  wire [10:0] _T_72997; // @[Modules.scala 68:83:@25695.4]
  wire [10:0] buffer_10_645; // @[Modules.scala 68:83:@25696.4]
  wire [11:0] _T_72999; // @[Modules.scala 68:83:@25698.4]
  wire [10:0] _T_73000; // @[Modules.scala 68:83:@25699.4]
  wire [10:0] buffer_10_646; // @[Modules.scala 68:83:@25700.4]
  wire [11:0] _T_73005; // @[Modules.scala 68:83:@25706.4]
  wire [10:0] _T_73006; // @[Modules.scala 68:83:@25707.4]
  wire [10:0] buffer_10_648; // @[Modules.scala 68:83:@25708.4]
  wire [11:0] _T_73008; // @[Modules.scala 68:83:@25710.4]
  wire [10:0] _T_73009; // @[Modules.scala 68:83:@25711.4]
  wire [10:0] buffer_10_649; // @[Modules.scala 68:83:@25712.4]
  wire [11:0] _T_73014; // @[Modules.scala 68:83:@25718.4]
  wire [10:0] _T_73015; // @[Modules.scala 68:83:@25719.4]
  wire [10:0] buffer_10_651; // @[Modules.scala 68:83:@25720.4]
  wire [11:0] _T_73017; // @[Modules.scala 68:83:@25722.4]
  wire [10:0] _T_73018; // @[Modules.scala 68:83:@25723.4]
  wire [10:0] buffer_10_652; // @[Modules.scala 68:83:@25724.4]
  wire [11:0] _T_73020; // @[Modules.scala 68:83:@25726.4]
  wire [10:0] _T_73021; // @[Modules.scala 68:83:@25727.4]
  wire [10:0] buffer_10_653; // @[Modules.scala 68:83:@25728.4]
  wire [11:0] _T_73026; // @[Modules.scala 68:83:@25734.4]
  wire [10:0] _T_73027; // @[Modules.scala 68:83:@25735.4]
  wire [10:0] buffer_10_655; // @[Modules.scala 68:83:@25736.4]
  wire [11:0] _T_73029; // @[Modules.scala 68:83:@25738.4]
  wire [10:0] _T_73030; // @[Modules.scala 68:83:@25739.4]
  wire [10:0] buffer_10_656; // @[Modules.scala 68:83:@25740.4]
  wire [11:0] _T_73032; // @[Modules.scala 68:83:@25742.4]
  wire [10:0] _T_73033; // @[Modules.scala 68:83:@25743.4]
  wire [10:0] buffer_10_657; // @[Modules.scala 68:83:@25744.4]
  wire [11:0] _T_73035; // @[Modules.scala 68:83:@25746.4]
  wire [10:0] _T_73036; // @[Modules.scala 68:83:@25747.4]
  wire [10:0] buffer_10_658; // @[Modules.scala 68:83:@25748.4]
  wire [11:0] _T_73038; // @[Modules.scala 68:83:@25750.4]
  wire [10:0] _T_73039; // @[Modules.scala 68:83:@25751.4]
  wire [10:0] buffer_10_659; // @[Modules.scala 68:83:@25752.4]
  wire [11:0] _T_73041; // @[Modules.scala 68:83:@25754.4]
  wire [10:0] _T_73042; // @[Modules.scala 68:83:@25755.4]
  wire [10:0] buffer_10_660; // @[Modules.scala 68:83:@25756.4]
  wire [11:0] _T_73053; // @[Modules.scala 68:83:@25770.4]
  wire [10:0] _T_73054; // @[Modules.scala 68:83:@25771.4]
  wire [10:0] buffer_10_664; // @[Modules.scala 68:83:@25772.4]
  wire [11:0] _T_73059; // @[Modules.scala 68:83:@25778.4]
  wire [10:0] _T_73060; // @[Modules.scala 68:83:@25779.4]
  wire [10:0] buffer_10_666; // @[Modules.scala 68:83:@25780.4]
  wire [11:0] _T_73062; // @[Modules.scala 68:83:@25782.4]
  wire [10:0] _T_73063; // @[Modules.scala 68:83:@25783.4]
  wire [10:0] buffer_10_667; // @[Modules.scala 68:83:@25784.4]
  wire [11:0] _T_73065; // @[Modules.scala 68:83:@25786.4]
  wire [10:0] _T_73066; // @[Modules.scala 68:83:@25787.4]
  wire [10:0] buffer_10_668; // @[Modules.scala 68:83:@25788.4]
  wire [11:0] _T_73068; // @[Modules.scala 68:83:@25790.4]
  wire [10:0] _T_73069; // @[Modules.scala 68:83:@25791.4]
  wire [10:0] buffer_10_669; // @[Modules.scala 68:83:@25792.4]
  wire [11:0] _T_73080; // @[Modules.scala 68:83:@25806.4]
  wire [10:0] _T_73081; // @[Modules.scala 68:83:@25807.4]
  wire [10:0] buffer_10_673; // @[Modules.scala 68:83:@25808.4]
  wire [11:0] _T_73089; // @[Modules.scala 68:83:@25818.4]
  wire [10:0] _T_73090; // @[Modules.scala 68:83:@25819.4]
  wire [10:0] buffer_10_676; // @[Modules.scala 68:83:@25820.4]
  wire [11:0] _T_73095; // @[Modules.scala 68:83:@25826.4]
  wire [10:0] _T_73096; // @[Modules.scala 68:83:@25827.4]
  wire [10:0] buffer_10_678; // @[Modules.scala 68:83:@25828.4]
  wire [11:0] _T_73098; // @[Modules.scala 68:83:@25830.4]
  wire [10:0] _T_73099; // @[Modules.scala 68:83:@25831.4]
  wire [10:0] buffer_10_679; // @[Modules.scala 68:83:@25832.4]
  wire [11:0] _T_73101; // @[Modules.scala 68:83:@25834.4]
  wire [10:0] _T_73102; // @[Modules.scala 68:83:@25835.4]
  wire [10:0] buffer_10_680; // @[Modules.scala 68:83:@25836.4]
  wire [11:0] _T_73107; // @[Modules.scala 68:83:@25842.4]
  wire [10:0] _T_73108; // @[Modules.scala 68:83:@25843.4]
  wire [10:0] buffer_10_682; // @[Modules.scala 68:83:@25844.4]
  wire [11:0] _T_73110; // @[Modules.scala 68:83:@25846.4]
  wire [10:0] _T_73111; // @[Modules.scala 68:83:@25847.4]
  wire [10:0] buffer_10_683; // @[Modules.scala 68:83:@25848.4]
  wire [11:0] _T_73116; // @[Modules.scala 68:83:@25854.4]
  wire [10:0] _T_73117; // @[Modules.scala 68:83:@25855.4]
  wire [10:0] buffer_10_685; // @[Modules.scala 68:83:@25856.4]
  wire [11:0] _T_73119; // @[Modules.scala 71:109:@25858.4]
  wire [10:0] _T_73120; // @[Modules.scala 71:109:@25859.4]
  wire [10:0] buffer_10_686; // @[Modules.scala 71:109:@25860.4]
  wire [11:0] _T_73122; // @[Modules.scala 71:109:@25862.4]
  wire [10:0] _T_73123; // @[Modules.scala 71:109:@25863.4]
  wire [10:0] buffer_10_687; // @[Modules.scala 71:109:@25864.4]
  wire [11:0] _T_73128; // @[Modules.scala 71:109:@25870.4]
  wire [10:0] _T_73129; // @[Modules.scala 71:109:@25871.4]
  wire [10:0] buffer_10_689; // @[Modules.scala 71:109:@25872.4]
  wire [11:0] _T_73134; // @[Modules.scala 71:109:@25878.4]
  wire [10:0] _T_73135; // @[Modules.scala 71:109:@25879.4]
  wire [10:0] buffer_10_691; // @[Modules.scala 71:109:@25880.4]
  wire [11:0] _T_73137; // @[Modules.scala 71:109:@25882.4]
  wire [10:0] _T_73138; // @[Modules.scala 71:109:@25883.4]
  wire [10:0] buffer_10_692; // @[Modules.scala 71:109:@25884.4]
  wire [11:0] _T_73140; // @[Modules.scala 71:109:@25886.4]
  wire [10:0] _T_73141; // @[Modules.scala 71:109:@25887.4]
  wire [10:0] buffer_10_693; // @[Modules.scala 71:109:@25888.4]
  wire [11:0] _T_73143; // @[Modules.scala 71:109:@25890.4]
  wire [10:0] _T_73144; // @[Modules.scala 71:109:@25891.4]
  wire [10:0] buffer_10_694; // @[Modules.scala 71:109:@25892.4]
  wire [11:0] _T_73146; // @[Modules.scala 71:109:@25894.4]
  wire [10:0] _T_73147; // @[Modules.scala 71:109:@25895.4]
  wire [10:0] buffer_10_695; // @[Modules.scala 71:109:@25896.4]
  wire [11:0] _T_73149; // @[Modules.scala 71:109:@25898.4]
  wire [10:0] _T_73150; // @[Modules.scala 71:109:@25899.4]
  wire [10:0] buffer_10_696; // @[Modules.scala 71:109:@25900.4]
  wire [11:0] _T_73152; // @[Modules.scala 71:109:@25902.4]
  wire [10:0] _T_73153; // @[Modules.scala 71:109:@25903.4]
  wire [10:0] buffer_10_697; // @[Modules.scala 71:109:@25904.4]
  wire [11:0] _T_73155; // @[Modules.scala 71:109:@25906.4]
  wire [10:0] _T_73156; // @[Modules.scala 71:109:@25907.4]
  wire [10:0] buffer_10_698; // @[Modules.scala 71:109:@25908.4]
  wire [11:0] _T_73158; // @[Modules.scala 71:109:@25910.4]
  wire [10:0] _T_73159; // @[Modules.scala 71:109:@25911.4]
  wire [10:0] buffer_10_699; // @[Modules.scala 71:109:@25912.4]
  wire [11:0] _T_73161; // @[Modules.scala 71:109:@25914.4]
  wire [10:0] _T_73162; // @[Modules.scala 71:109:@25915.4]
  wire [10:0] buffer_10_700; // @[Modules.scala 71:109:@25916.4]
  wire [11:0] _T_73164; // @[Modules.scala 71:109:@25918.4]
  wire [10:0] _T_73165; // @[Modules.scala 71:109:@25919.4]
  wire [10:0] buffer_10_701; // @[Modules.scala 71:109:@25920.4]
  wire [11:0] _T_73167; // @[Modules.scala 71:109:@25922.4]
  wire [10:0] _T_73168; // @[Modules.scala 71:109:@25923.4]
  wire [10:0] buffer_10_702; // @[Modules.scala 71:109:@25924.4]
  wire [11:0] _T_73170; // @[Modules.scala 71:109:@25926.4]
  wire [10:0] _T_73171; // @[Modules.scala 71:109:@25927.4]
  wire [10:0] buffer_10_703; // @[Modules.scala 71:109:@25928.4]
  wire [11:0] _T_73173; // @[Modules.scala 71:109:@25930.4]
  wire [10:0] _T_73174; // @[Modules.scala 71:109:@25931.4]
  wire [10:0] buffer_10_704; // @[Modules.scala 71:109:@25932.4]
  wire [11:0] _T_73176; // @[Modules.scala 71:109:@25934.4]
  wire [10:0] _T_73177; // @[Modules.scala 71:109:@25935.4]
  wire [10:0] buffer_10_705; // @[Modules.scala 71:109:@25936.4]
  wire [11:0] _T_73179; // @[Modules.scala 71:109:@25938.4]
  wire [10:0] _T_73180; // @[Modules.scala 71:109:@25939.4]
  wire [10:0] buffer_10_706; // @[Modules.scala 71:109:@25940.4]
  wire [11:0] _T_73185; // @[Modules.scala 71:109:@25946.4]
  wire [10:0] _T_73186; // @[Modules.scala 71:109:@25947.4]
  wire [10:0] buffer_10_708; // @[Modules.scala 71:109:@25948.4]
  wire [11:0] _T_73188; // @[Modules.scala 71:109:@25950.4]
  wire [10:0] _T_73189; // @[Modules.scala 71:109:@25951.4]
  wire [10:0] buffer_10_709; // @[Modules.scala 71:109:@25952.4]
  wire [11:0] _T_73191; // @[Modules.scala 71:109:@25954.4]
  wire [10:0] _T_73192; // @[Modules.scala 71:109:@25955.4]
  wire [10:0] buffer_10_710; // @[Modules.scala 71:109:@25956.4]
  wire [11:0] _T_73194; // @[Modules.scala 71:109:@25958.4]
  wire [10:0] _T_73195; // @[Modules.scala 71:109:@25959.4]
  wire [10:0] buffer_10_711; // @[Modules.scala 71:109:@25960.4]
  wire [11:0] _T_73197; // @[Modules.scala 71:109:@25962.4]
  wire [10:0] _T_73198; // @[Modules.scala 71:109:@25963.4]
  wire [10:0] buffer_10_712; // @[Modules.scala 71:109:@25964.4]
  wire [11:0] _T_73200; // @[Modules.scala 71:109:@25966.4]
  wire [10:0] _T_73201; // @[Modules.scala 71:109:@25967.4]
  wire [10:0] buffer_10_713; // @[Modules.scala 71:109:@25968.4]
  wire [11:0] _T_73203; // @[Modules.scala 71:109:@25970.4]
  wire [10:0] _T_73204; // @[Modules.scala 71:109:@25971.4]
  wire [10:0] buffer_10_714; // @[Modules.scala 71:109:@25972.4]
  wire [11:0] _T_73206; // @[Modules.scala 71:109:@25974.4]
  wire [10:0] _T_73207; // @[Modules.scala 71:109:@25975.4]
  wire [10:0] buffer_10_715; // @[Modules.scala 71:109:@25976.4]
  wire [11:0] _T_73209; // @[Modules.scala 71:109:@25978.4]
  wire [10:0] _T_73210; // @[Modules.scala 71:109:@25979.4]
  wire [10:0] buffer_10_716; // @[Modules.scala 71:109:@25980.4]
  wire [11:0] _T_73212; // @[Modules.scala 71:109:@25982.4]
  wire [10:0] _T_73213; // @[Modules.scala 71:109:@25983.4]
  wire [10:0] buffer_10_717; // @[Modules.scala 71:109:@25984.4]
  wire [11:0] _T_73215; // @[Modules.scala 71:109:@25986.4]
  wire [10:0] _T_73216; // @[Modules.scala 71:109:@25987.4]
  wire [10:0] buffer_10_718; // @[Modules.scala 71:109:@25988.4]
  wire [11:0] _T_73218; // @[Modules.scala 71:109:@25990.4]
  wire [10:0] _T_73219; // @[Modules.scala 71:109:@25991.4]
  wire [10:0] buffer_10_719; // @[Modules.scala 71:109:@25992.4]
  wire [11:0] _T_73221; // @[Modules.scala 71:109:@25994.4]
  wire [10:0] _T_73222; // @[Modules.scala 71:109:@25995.4]
  wire [10:0] buffer_10_720; // @[Modules.scala 71:109:@25996.4]
  wire [11:0] _T_73224; // @[Modules.scala 71:109:@25998.4]
  wire [10:0] _T_73225; // @[Modules.scala 71:109:@25999.4]
  wire [10:0] buffer_10_721; // @[Modules.scala 71:109:@26000.4]
  wire [11:0] _T_73227; // @[Modules.scala 71:109:@26002.4]
  wire [10:0] _T_73228; // @[Modules.scala 71:109:@26003.4]
  wire [10:0] buffer_10_722; // @[Modules.scala 71:109:@26004.4]
  wire [11:0] _T_73230; // @[Modules.scala 71:109:@26006.4]
  wire [10:0] _T_73231; // @[Modules.scala 71:109:@26007.4]
  wire [10:0] buffer_10_723; // @[Modules.scala 71:109:@26008.4]
  wire [11:0] _T_73233; // @[Modules.scala 71:109:@26010.4]
  wire [10:0] _T_73234; // @[Modules.scala 71:109:@26011.4]
  wire [10:0] buffer_10_724; // @[Modules.scala 71:109:@26012.4]
  wire [11:0] _T_73236; // @[Modules.scala 71:109:@26014.4]
  wire [10:0] _T_73237; // @[Modules.scala 71:109:@26015.4]
  wire [10:0] buffer_10_725; // @[Modules.scala 71:109:@26016.4]
  wire [11:0] _T_73239; // @[Modules.scala 71:109:@26018.4]
  wire [10:0] _T_73240; // @[Modules.scala 71:109:@26019.4]
  wire [10:0] buffer_10_726; // @[Modules.scala 71:109:@26020.4]
  wire [11:0] _T_73242; // @[Modules.scala 71:109:@26022.4]
  wire [10:0] _T_73243; // @[Modules.scala 71:109:@26023.4]
  wire [10:0] buffer_10_727; // @[Modules.scala 71:109:@26024.4]
  wire [11:0] _T_73245; // @[Modules.scala 71:109:@26026.4]
  wire [10:0] _T_73246; // @[Modules.scala 71:109:@26027.4]
  wire [10:0] buffer_10_728; // @[Modules.scala 71:109:@26028.4]
  wire [11:0] _T_73248; // @[Modules.scala 71:109:@26030.4]
  wire [10:0] _T_73249; // @[Modules.scala 71:109:@26031.4]
  wire [10:0] buffer_10_729; // @[Modules.scala 71:109:@26032.4]
  wire [11:0] _T_73251; // @[Modules.scala 71:109:@26034.4]
  wire [10:0] _T_73252; // @[Modules.scala 71:109:@26035.4]
  wire [10:0] buffer_10_730; // @[Modules.scala 71:109:@26036.4]
  wire [11:0] _T_73254; // @[Modules.scala 71:109:@26038.4]
  wire [10:0] _T_73255; // @[Modules.scala 71:109:@26039.4]
  wire [10:0] buffer_10_731; // @[Modules.scala 71:109:@26040.4]
  wire [11:0] _T_73257; // @[Modules.scala 71:109:@26042.4]
  wire [10:0] _T_73258; // @[Modules.scala 71:109:@26043.4]
  wire [10:0] buffer_10_732; // @[Modules.scala 71:109:@26044.4]
  wire [11:0] _T_73260; // @[Modules.scala 71:109:@26046.4]
  wire [10:0] _T_73261; // @[Modules.scala 71:109:@26047.4]
  wire [10:0] buffer_10_733; // @[Modules.scala 71:109:@26048.4]
  wire [11:0] _T_73263; // @[Modules.scala 71:109:@26050.4]
  wire [10:0] _T_73264; // @[Modules.scala 71:109:@26051.4]
  wire [10:0] buffer_10_734; // @[Modules.scala 71:109:@26052.4]
  wire [11:0] _T_73266; // @[Modules.scala 78:156:@26055.4]
  wire [10:0] _T_73267; // @[Modules.scala 78:156:@26056.4]
  wire [10:0] buffer_10_736; // @[Modules.scala 78:156:@26057.4]
  wire [11:0] _T_73269; // @[Modules.scala 78:156:@26059.4]
  wire [10:0] _T_73270; // @[Modules.scala 78:156:@26060.4]
  wire [10:0] buffer_10_737; // @[Modules.scala 78:156:@26061.4]
  wire [11:0] _T_73272; // @[Modules.scala 78:156:@26063.4]
  wire [10:0] _T_73273; // @[Modules.scala 78:156:@26064.4]
  wire [10:0] buffer_10_738; // @[Modules.scala 78:156:@26065.4]
  wire [11:0] _T_73275; // @[Modules.scala 78:156:@26067.4]
  wire [10:0] _T_73276; // @[Modules.scala 78:156:@26068.4]
  wire [10:0] buffer_10_739; // @[Modules.scala 78:156:@26069.4]
  wire [11:0] _T_73278; // @[Modules.scala 78:156:@26071.4]
  wire [10:0] _T_73279; // @[Modules.scala 78:156:@26072.4]
  wire [10:0] buffer_10_740; // @[Modules.scala 78:156:@26073.4]
  wire [11:0] _T_73281; // @[Modules.scala 78:156:@26075.4]
  wire [10:0] _T_73282; // @[Modules.scala 78:156:@26076.4]
  wire [10:0] buffer_10_741; // @[Modules.scala 78:156:@26077.4]
  wire [11:0] _T_73284; // @[Modules.scala 78:156:@26079.4]
  wire [10:0] _T_73285; // @[Modules.scala 78:156:@26080.4]
  wire [10:0] buffer_10_742; // @[Modules.scala 78:156:@26081.4]
  wire [11:0] _T_73287; // @[Modules.scala 78:156:@26083.4]
  wire [10:0] _T_73288; // @[Modules.scala 78:156:@26084.4]
  wire [10:0] buffer_10_743; // @[Modules.scala 78:156:@26085.4]
  wire [11:0] _T_73290; // @[Modules.scala 78:156:@26087.4]
  wire [10:0] _T_73291; // @[Modules.scala 78:156:@26088.4]
  wire [10:0] buffer_10_744; // @[Modules.scala 78:156:@26089.4]
  wire [11:0] _T_73293; // @[Modules.scala 78:156:@26091.4]
  wire [10:0] _T_73294; // @[Modules.scala 78:156:@26092.4]
  wire [10:0] buffer_10_745; // @[Modules.scala 78:156:@26093.4]
  wire [11:0] _T_73296; // @[Modules.scala 78:156:@26095.4]
  wire [10:0] _T_73297; // @[Modules.scala 78:156:@26096.4]
  wire [10:0] buffer_10_746; // @[Modules.scala 78:156:@26097.4]
  wire [11:0] _T_73299; // @[Modules.scala 78:156:@26099.4]
  wire [10:0] _T_73300; // @[Modules.scala 78:156:@26100.4]
  wire [10:0] buffer_10_747; // @[Modules.scala 78:156:@26101.4]
  wire [11:0] _T_73302; // @[Modules.scala 78:156:@26103.4]
  wire [10:0] _T_73303; // @[Modules.scala 78:156:@26104.4]
  wire [10:0] buffer_10_748; // @[Modules.scala 78:156:@26105.4]
  wire [11:0] _T_73305; // @[Modules.scala 78:156:@26107.4]
  wire [10:0] _T_73306; // @[Modules.scala 78:156:@26108.4]
  wire [10:0] buffer_10_749; // @[Modules.scala 78:156:@26109.4]
  wire [11:0] _T_73308; // @[Modules.scala 78:156:@26111.4]
  wire [10:0] _T_73309; // @[Modules.scala 78:156:@26112.4]
  wire [10:0] buffer_10_750; // @[Modules.scala 78:156:@26113.4]
  wire [11:0] _T_73311; // @[Modules.scala 78:156:@26115.4]
  wire [10:0] _T_73312; // @[Modules.scala 78:156:@26116.4]
  wire [10:0] buffer_10_751; // @[Modules.scala 78:156:@26117.4]
  wire [11:0] _T_73314; // @[Modules.scala 78:156:@26119.4]
  wire [10:0] _T_73315; // @[Modules.scala 78:156:@26120.4]
  wire [10:0] buffer_10_752; // @[Modules.scala 78:156:@26121.4]
  wire [11:0] _T_73317; // @[Modules.scala 78:156:@26123.4]
  wire [10:0] _T_73318; // @[Modules.scala 78:156:@26124.4]
  wire [10:0] buffer_10_753; // @[Modules.scala 78:156:@26125.4]
  wire [11:0] _T_73320; // @[Modules.scala 78:156:@26127.4]
  wire [10:0] _T_73321; // @[Modules.scala 78:156:@26128.4]
  wire [10:0] buffer_10_754; // @[Modules.scala 78:156:@26129.4]
  wire [11:0] _T_73323; // @[Modules.scala 78:156:@26131.4]
  wire [10:0] _T_73324; // @[Modules.scala 78:156:@26132.4]
  wire [10:0] buffer_10_755; // @[Modules.scala 78:156:@26133.4]
  wire [11:0] _T_73326; // @[Modules.scala 78:156:@26135.4]
  wire [10:0] _T_73327; // @[Modules.scala 78:156:@26136.4]
  wire [10:0] buffer_10_756; // @[Modules.scala 78:156:@26137.4]
  wire [11:0] _T_73329; // @[Modules.scala 78:156:@26139.4]
  wire [10:0] _T_73330; // @[Modules.scala 78:156:@26140.4]
  wire [10:0] buffer_10_757; // @[Modules.scala 78:156:@26141.4]
  wire [11:0] _T_73332; // @[Modules.scala 78:156:@26143.4]
  wire [10:0] _T_73333; // @[Modules.scala 78:156:@26144.4]
  wire [10:0] buffer_10_758; // @[Modules.scala 78:156:@26145.4]
  wire [11:0] _T_73335; // @[Modules.scala 78:156:@26147.4]
  wire [10:0] _T_73336; // @[Modules.scala 78:156:@26148.4]
  wire [10:0] buffer_10_759; // @[Modules.scala 78:156:@26149.4]
  wire [11:0] _T_73338; // @[Modules.scala 78:156:@26151.4]
  wire [10:0] _T_73339; // @[Modules.scala 78:156:@26152.4]
  wire [10:0] buffer_10_760; // @[Modules.scala 78:156:@26153.4]
  wire [11:0] _T_73341; // @[Modules.scala 78:156:@26155.4]
  wire [10:0] _T_73342; // @[Modules.scala 78:156:@26156.4]
  wire [10:0] buffer_10_761; // @[Modules.scala 78:156:@26157.4]
  wire [11:0] _T_73344; // @[Modules.scala 78:156:@26159.4]
  wire [10:0] _T_73345; // @[Modules.scala 78:156:@26160.4]
  wire [10:0] buffer_10_762; // @[Modules.scala 78:156:@26161.4]
  wire [11:0] _T_73347; // @[Modules.scala 78:156:@26163.4]
  wire [10:0] _T_73348; // @[Modules.scala 78:156:@26164.4]
  wire [10:0] buffer_10_763; // @[Modules.scala 78:156:@26165.4]
  wire [11:0] _T_73350; // @[Modules.scala 78:156:@26167.4]
  wire [10:0] _T_73351; // @[Modules.scala 78:156:@26168.4]
  wire [10:0] buffer_10_764; // @[Modules.scala 78:156:@26169.4]
  wire [11:0] _T_73353; // @[Modules.scala 78:156:@26171.4]
  wire [10:0] _T_73354; // @[Modules.scala 78:156:@26172.4]
  wire [10:0] buffer_10_765; // @[Modules.scala 78:156:@26173.4]
  wire [11:0] _T_73356; // @[Modules.scala 78:156:@26175.4]
  wire [10:0] _T_73357; // @[Modules.scala 78:156:@26176.4]
  wire [10:0] buffer_10_766; // @[Modules.scala 78:156:@26177.4]
  wire [11:0] _T_73359; // @[Modules.scala 78:156:@26179.4]
  wire [10:0] _T_73360; // @[Modules.scala 78:156:@26180.4]
  wire [10:0] buffer_10_767; // @[Modules.scala 78:156:@26181.4]
  wire [11:0] _T_73362; // @[Modules.scala 78:156:@26183.4]
  wire [10:0] _T_73363; // @[Modules.scala 78:156:@26184.4]
  wire [10:0] buffer_10_768; // @[Modules.scala 78:156:@26185.4]
  wire [11:0] _T_73365; // @[Modules.scala 78:156:@26187.4]
  wire [10:0] _T_73366; // @[Modules.scala 78:156:@26188.4]
  wire [10:0] buffer_10_769; // @[Modules.scala 78:156:@26189.4]
  wire [11:0] _T_73368; // @[Modules.scala 78:156:@26191.4]
  wire [10:0] _T_73369; // @[Modules.scala 78:156:@26192.4]
  wire [10:0] buffer_10_770; // @[Modules.scala 78:156:@26193.4]
  wire [11:0] _T_73371; // @[Modules.scala 78:156:@26195.4]
  wire [10:0] _T_73372; // @[Modules.scala 78:156:@26196.4]
  wire [10:0] buffer_10_771; // @[Modules.scala 78:156:@26197.4]
  wire [11:0] _T_73374; // @[Modules.scala 78:156:@26199.4]
  wire [10:0] _T_73375; // @[Modules.scala 78:156:@26200.4]
  wire [10:0] buffer_10_772; // @[Modules.scala 78:156:@26201.4]
  wire [11:0] _T_73377; // @[Modules.scala 78:156:@26203.4]
  wire [10:0] _T_73378; // @[Modules.scala 78:156:@26204.4]
  wire [10:0] buffer_10_773; // @[Modules.scala 78:156:@26205.4]
  wire [11:0] _T_73380; // @[Modules.scala 78:156:@26207.4]
  wire [10:0] _T_73381; // @[Modules.scala 78:156:@26208.4]
  wire [10:0] buffer_10_774; // @[Modules.scala 78:156:@26209.4]
  wire [11:0] _T_73383; // @[Modules.scala 78:156:@26211.4]
  wire [10:0] _T_73384; // @[Modules.scala 78:156:@26212.4]
  wire [10:0] buffer_10_775; // @[Modules.scala 78:156:@26213.4]
  wire [11:0] _T_73386; // @[Modules.scala 78:156:@26215.4]
  wire [10:0] _T_73387; // @[Modules.scala 78:156:@26216.4]
  wire [10:0] buffer_10_776; // @[Modules.scala 78:156:@26217.4]
  wire [11:0] _T_73389; // @[Modules.scala 78:156:@26219.4]
  wire [10:0] _T_73390; // @[Modules.scala 78:156:@26220.4]
  wire [10:0] buffer_10_777; // @[Modules.scala 78:156:@26221.4]
  wire [11:0] _T_73392; // @[Modules.scala 78:156:@26223.4]
  wire [10:0] _T_73393; // @[Modules.scala 78:156:@26224.4]
  wire [10:0] buffer_10_778; // @[Modules.scala 78:156:@26225.4]
  wire [11:0] _T_73395; // @[Modules.scala 78:156:@26227.4]
  wire [10:0] _T_73396; // @[Modules.scala 78:156:@26228.4]
  wire [10:0] buffer_10_779; // @[Modules.scala 78:156:@26229.4]
  wire [11:0] _T_73398; // @[Modules.scala 78:156:@26231.4]
  wire [10:0] _T_73399; // @[Modules.scala 78:156:@26232.4]
  wire [10:0] buffer_10_780; // @[Modules.scala 78:156:@26233.4]
  wire [11:0] _T_73401; // @[Modules.scala 78:156:@26235.4]
  wire [10:0] _T_73402; // @[Modules.scala 78:156:@26236.4]
  wire [10:0] buffer_10_781; // @[Modules.scala 78:156:@26237.4]
  wire [11:0] _T_73404; // @[Modules.scala 78:156:@26239.4]
  wire [10:0] _T_73405; // @[Modules.scala 78:156:@26240.4]
  wire [10:0] buffer_10_782; // @[Modules.scala 78:156:@26241.4]
  wire [11:0] _T_73407; // @[Modules.scala 78:156:@26243.4]
  wire [10:0] _T_73408; // @[Modules.scala 78:156:@26244.4]
  wire [10:0] buffer_10_783; // @[Modules.scala 78:156:@26245.4]
  wire [5:0] _T_73466; // @[Modules.scala 37:46:@26333.4]
  wire [4:0] _T_73467; // @[Modules.scala 37:46:@26334.4]
  wire [4:0] _T_73468; // @[Modules.scala 37:46:@26335.4]
  wire [11:0] _T_73916; // @[Modules.scala 65:57:@26968.4]
  wire [10:0] _T_73917; // @[Modules.scala 65:57:@26969.4]
  wire [10:0] buffer_11_396; // @[Modules.scala 65:57:@26970.4]
  wire [11:0] _T_73925; // @[Modules.scala 65:57:@26980.4]
  wire [10:0] _T_73926; // @[Modules.scala 65:57:@26981.4]
  wire [10:0] buffer_11_399; // @[Modules.scala 65:57:@26982.4]
  wire [10:0] buffer_11_19; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_73931; // @[Modules.scala 65:57:@26988.4]
  wire [10:0] _T_73932; // @[Modules.scala 65:57:@26989.4]
  wire [10:0] buffer_11_401; // @[Modules.scala 65:57:@26990.4]
  wire [10:0] buffer_11_22; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_11_23; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_73937; // @[Modules.scala 65:57:@26996.4]
  wire [10:0] _T_73938; // @[Modules.scala 65:57:@26997.4]
  wire [10:0] buffer_11_403; // @[Modules.scala 65:57:@26998.4]
  wire [11:0] _T_73943; // @[Modules.scala 65:57:@27004.4]
  wire [10:0] _T_73944; // @[Modules.scala 65:57:@27005.4]
  wire [10:0] buffer_11_405; // @[Modules.scala 65:57:@27006.4]
  wire [11:0] _T_73946; // @[Modules.scala 65:57:@27008.4]
  wire [10:0] _T_73947; // @[Modules.scala 65:57:@27009.4]
  wire [10:0] buffer_11_406; // @[Modules.scala 65:57:@27010.4]
  wire [11:0] _T_73955; // @[Modules.scala 65:57:@27020.4]
  wire [10:0] _T_73956; // @[Modules.scala 65:57:@27021.4]
  wire [10:0] buffer_11_409; // @[Modules.scala 65:57:@27022.4]
  wire [10:0] buffer_11_43; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_73967; // @[Modules.scala 65:57:@27036.4]
  wire [10:0] _T_73968; // @[Modules.scala 65:57:@27037.4]
  wire [10:0] buffer_11_413; // @[Modules.scala 65:57:@27038.4]
  wire [11:0] _T_73970; // @[Modules.scala 65:57:@27040.4]
  wire [10:0] _T_73971; // @[Modules.scala 65:57:@27041.4]
  wire [10:0] buffer_11_414; // @[Modules.scala 65:57:@27042.4]
  wire [11:0] _T_74006; // @[Modules.scala 65:57:@27088.4]
  wire [10:0] _T_74007; // @[Modules.scala 65:57:@27089.4]
  wire [10:0] buffer_11_426; // @[Modules.scala 65:57:@27090.4]
  wire [11:0] _T_74009; // @[Modules.scala 65:57:@27092.4]
  wire [10:0] _T_74010; // @[Modules.scala 65:57:@27093.4]
  wire [10:0] buffer_11_427; // @[Modules.scala 65:57:@27094.4]
  wire [11:0] _T_74027; // @[Modules.scala 65:57:@27116.4]
  wire [10:0] _T_74028; // @[Modules.scala 65:57:@27117.4]
  wire [10:0] buffer_11_433; // @[Modules.scala 65:57:@27118.4]
  wire [10:0] buffer_11_90; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74039; // @[Modules.scala 65:57:@27132.4]
  wire [10:0] _T_74040; // @[Modules.scala 65:57:@27133.4]
  wire [10:0] buffer_11_437; // @[Modules.scala 65:57:@27134.4]
  wire [11:0] _T_74042; // @[Modules.scala 65:57:@27136.4]
  wire [10:0] _T_74043; // @[Modules.scala 65:57:@27137.4]
  wire [10:0] buffer_11_438; // @[Modules.scala 65:57:@27138.4]
  wire [11:0] _T_74045; // @[Modules.scala 65:57:@27140.4]
  wire [10:0] _T_74046; // @[Modules.scala 65:57:@27141.4]
  wire [10:0] buffer_11_439; // @[Modules.scala 65:57:@27142.4]
  wire [10:0] buffer_11_105; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74060; // @[Modules.scala 65:57:@27160.4]
  wire [10:0] _T_74061; // @[Modules.scala 65:57:@27161.4]
  wire [10:0] buffer_11_444; // @[Modules.scala 65:57:@27162.4]
  wire [11:0] _T_74063; // @[Modules.scala 65:57:@27164.4]
  wire [10:0] _T_74064; // @[Modules.scala 65:57:@27165.4]
  wire [10:0] buffer_11_445; // @[Modules.scala 65:57:@27166.4]
  wire [10:0] buffer_11_112; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74072; // @[Modules.scala 65:57:@27176.4]
  wire [10:0] _T_74073; // @[Modules.scala 65:57:@27177.4]
  wire [10:0] buffer_11_448; // @[Modules.scala 65:57:@27178.4]
  wire [11:0] _T_74078; // @[Modules.scala 65:57:@27184.4]
  wire [10:0] _T_74079; // @[Modules.scala 65:57:@27185.4]
  wire [10:0] buffer_11_450; // @[Modules.scala 65:57:@27186.4]
  wire [10:0] buffer_11_119; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74081; // @[Modules.scala 65:57:@27188.4]
  wire [10:0] _T_74082; // @[Modules.scala 65:57:@27189.4]
  wire [10:0] buffer_11_451; // @[Modules.scala 65:57:@27190.4]
  wire [11:0] _T_74084; // @[Modules.scala 65:57:@27192.4]
  wire [10:0] _T_74085; // @[Modules.scala 65:57:@27193.4]
  wire [10:0] buffer_11_452; // @[Modules.scala 65:57:@27194.4]
  wire [11:0] _T_74087; // @[Modules.scala 65:57:@27196.4]
  wire [10:0] _T_74088; // @[Modules.scala 65:57:@27197.4]
  wire [10:0] buffer_11_453; // @[Modules.scala 65:57:@27198.4]
  wire [11:0] _T_74096; // @[Modules.scala 65:57:@27208.4]
  wire [10:0] _T_74097; // @[Modules.scala 65:57:@27209.4]
  wire [10:0] buffer_11_456; // @[Modules.scala 65:57:@27210.4]
  wire [11:0] _T_74102; // @[Modules.scala 65:57:@27216.4]
  wire [10:0] _T_74103; // @[Modules.scala 65:57:@27217.4]
  wire [10:0] buffer_11_458; // @[Modules.scala 65:57:@27218.4]
  wire [10:0] buffer_11_135; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74105; // @[Modules.scala 65:57:@27220.4]
  wire [10:0] _T_74106; // @[Modules.scala 65:57:@27221.4]
  wire [10:0] buffer_11_459; // @[Modules.scala 65:57:@27222.4]
  wire [11:0] _T_74114; // @[Modules.scala 65:57:@27232.4]
  wire [10:0] _T_74115; // @[Modules.scala 65:57:@27233.4]
  wire [10:0] buffer_11_462; // @[Modules.scala 65:57:@27234.4]
  wire [11:0] _T_74117; // @[Modules.scala 65:57:@27236.4]
  wire [10:0] _T_74118; // @[Modules.scala 65:57:@27237.4]
  wire [10:0] buffer_11_463; // @[Modules.scala 65:57:@27238.4]
  wire [11:0] _T_74138; // @[Modules.scala 65:57:@27264.4]
  wire [10:0] _T_74139; // @[Modules.scala 65:57:@27265.4]
  wire [10:0] buffer_11_470; // @[Modules.scala 65:57:@27266.4]
  wire [11:0] _T_74144; // @[Modules.scala 65:57:@27272.4]
  wire [10:0] _T_74145; // @[Modules.scala 65:57:@27273.4]
  wire [10:0] buffer_11_472; // @[Modules.scala 65:57:@27274.4]
  wire [11:0] _T_74174; // @[Modules.scala 65:57:@27312.4]
  wire [10:0] _T_74175; // @[Modules.scala 65:57:@27313.4]
  wire [10:0] buffer_11_482; // @[Modules.scala 65:57:@27314.4]
  wire [10:0] buffer_11_185; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74180; // @[Modules.scala 65:57:@27320.4]
  wire [10:0] _T_74181; // @[Modules.scala 65:57:@27321.4]
  wire [10:0] buffer_11_484; // @[Modules.scala 65:57:@27322.4]
  wire [10:0] buffer_11_186; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74183; // @[Modules.scala 65:57:@27324.4]
  wire [10:0] _T_74184; // @[Modules.scala 65:57:@27325.4]
  wire [10:0] buffer_11_485; // @[Modules.scala 65:57:@27326.4]
  wire [11:0] _T_74195; // @[Modules.scala 65:57:@27340.4]
  wire [10:0] _T_74196; // @[Modules.scala 65:57:@27341.4]
  wire [10:0] buffer_11_489; // @[Modules.scala 65:57:@27342.4]
  wire [11:0] _T_74204; // @[Modules.scala 65:57:@27352.4]
  wire [10:0] _T_74205; // @[Modules.scala 65:57:@27353.4]
  wire [10:0] buffer_11_492; // @[Modules.scala 65:57:@27354.4]
  wire [11:0] _T_74219; // @[Modules.scala 65:57:@27372.4]
  wire [10:0] _T_74220; // @[Modules.scala 65:57:@27373.4]
  wire [10:0] buffer_11_497; // @[Modules.scala 65:57:@27374.4]
  wire [10:0] buffer_11_214; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74225; // @[Modules.scala 65:57:@27380.4]
  wire [10:0] _T_74226; // @[Modules.scala 65:57:@27381.4]
  wire [10:0] buffer_11_499; // @[Modules.scala 65:57:@27382.4]
  wire [10:0] buffer_11_217; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74228; // @[Modules.scala 65:57:@27384.4]
  wire [10:0] _T_74229; // @[Modules.scala 65:57:@27385.4]
  wire [10:0] buffer_11_500; // @[Modules.scala 65:57:@27386.4]
  wire [10:0] buffer_11_225; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74240; // @[Modules.scala 65:57:@27400.4]
  wire [10:0] _T_74241; // @[Modules.scala 65:57:@27401.4]
  wire [10:0] buffer_11_504; // @[Modules.scala 65:57:@27402.4]
  wire [11:0] _T_74246; // @[Modules.scala 65:57:@27408.4]
  wire [10:0] _T_74247; // @[Modules.scala 65:57:@27409.4]
  wire [10:0] buffer_11_506; // @[Modules.scala 65:57:@27410.4]
  wire [10:0] buffer_11_235; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74255; // @[Modules.scala 65:57:@27420.4]
  wire [10:0] _T_74256; // @[Modules.scala 65:57:@27421.4]
  wire [10:0] buffer_11_509; // @[Modules.scala 65:57:@27422.4]
  wire [11:0] _T_74261; // @[Modules.scala 65:57:@27428.4]
  wire [10:0] _T_74262; // @[Modules.scala 65:57:@27429.4]
  wire [10:0] buffer_11_511; // @[Modules.scala 65:57:@27430.4]
  wire [10:0] buffer_11_240; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74264; // @[Modules.scala 65:57:@27432.4]
  wire [10:0] _T_74265; // @[Modules.scala 65:57:@27433.4]
  wire [10:0] buffer_11_512; // @[Modules.scala 65:57:@27434.4]
  wire [10:0] buffer_11_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74276; // @[Modules.scala 65:57:@27448.4]
  wire [10:0] _T_74277; // @[Modules.scala 65:57:@27449.4]
  wire [10:0] buffer_11_516; // @[Modules.scala 65:57:@27450.4]
  wire [11:0] _T_74288; // @[Modules.scala 65:57:@27464.4]
  wire [10:0] _T_74289; // @[Modules.scala 65:57:@27465.4]
  wire [10:0] buffer_11_520; // @[Modules.scala 65:57:@27466.4]
  wire [10:0] buffer_11_258; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74291; // @[Modules.scala 65:57:@27468.4]
  wire [10:0] _T_74292; // @[Modules.scala 65:57:@27469.4]
  wire [10:0] buffer_11_521; // @[Modules.scala 65:57:@27470.4]
  wire [11:0] _T_74297; // @[Modules.scala 65:57:@27476.4]
  wire [10:0] _T_74298; // @[Modules.scala 65:57:@27477.4]
  wire [10:0] buffer_11_523; // @[Modules.scala 65:57:@27478.4]
  wire [11:0] _T_74309; // @[Modules.scala 65:57:@27492.4]
  wire [10:0] _T_74310; // @[Modules.scala 65:57:@27493.4]
  wire [10:0] buffer_11_527; // @[Modules.scala 65:57:@27494.4]
  wire [11:0] _T_74312; // @[Modules.scala 65:57:@27496.4]
  wire [10:0] _T_74313; // @[Modules.scala 65:57:@27497.4]
  wire [10:0] buffer_11_528; // @[Modules.scala 65:57:@27498.4]
  wire [11:0] _T_74318; // @[Modules.scala 65:57:@27504.4]
  wire [10:0] _T_74319; // @[Modules.scala 65:57:@27505.4]
  wire [10:0] buffer_11_530; // @[Modules.scala 65:57:@27506.4]
  wire [10:0] buffer_11_281; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74324; // @[Modules.scala 65:57:@27512.4]
  wire [10:0] _T_74325; // @[Modules.scala 65:57:@27513.4]
  wire [10:0] buffer_11_532; // @[Modules.scala 65:57:@27514.4]
  wire [11:0] _T_74333; // @[Modules.scala 65:57:@27524.4]
  wire [10:0] _T_74334; // @[Modules.scala 65:57:@27525.4]
  wire [10:0] buffer_11_535; // @[Modules.scala 65:57:@27526.4]
  wire [11:0] _T_74339; // @[Modules.scala 65:57:@27532.4]
  wire [10:0] _T_74340; // @[Modules.scala 65:57:@27533.4]
  wire [10:0] buffer_11_537; // @[Modules.scala 65:57:@27534.4]
  wire [11:0] _T_74348; // @[Modules.scala 65:57:@27544.4]
  wire [10:0] _T_74349; // @[Modules.scala 65:57:@27545.4]
  wire [10:0] buffer_11_540; // @[Modules.scala 65:57:@27546.4]
  wire [11:0] _T_74357; // @[Modules.scala 65:57:@27556.4]
  wire [10:0] _T_74358; // @[Modules.scala 65:57:@27557.4]
  wire [10:0] buffer_11_543; // @[Modules.scala 65:57:@27558.4]
  wire [10:0] buffer_11_310; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74369; // @[Modules.scala 65:57:@27572.4]
  wire [10:0] _T_74370; // @[Modules.scala 65:57:@27573.4]
  wire [10:0] buffer_11_547; // @[Modules.scala 65:57:@27574.4]
  wire [11:0] _T_74372; // @[Modules.scala 65:57:@27576.4]
  wire [10:0] _T_74373; // @[Modules.scala 65:57:@27577.4]
  wire [10:0] buffer_11_548; // @[Modules.scala 65:57:@27578.4]
  wire [11:0] _T_74384; // @[Modules.scala 65:57:@27592.4]
  wire [10:0] _T_74385; // @[Modules.scala 65:57:@27593.4]
  wire [10:0] buffer_11_552; // @[Modules.scala 65:57:@27594.4]
  wire [11:0] _T_74393; // @[Modules.scala 65:57:@27604.4]
  wire [10:0] _T_74394; // @[Modules.scala 65:57:@27605.4]
  wire [10:0] buffer_11_555; // @[Modules.scala 65:57:@27606.4]
  wire [11:0] _T_74423; // @[Modules.scala 65:57:@27644.4]
  wire [10:0] _T_74424; // @[Modules.scala 65:57:@27645.4]
  wire [10:0] buffer_11_565; // @[Modules.scala 65:57:@27646.4]
  wire [11:0] _T_74429; // @[Modules.scala 65:57:@27652.4]
  wire [10:0] _T_74430; // @[Modules.scala 65:57:@27653.4]
  wire [10:0] buffer_11_567; // @[Modules.scala 65:57:@27654.4]
  wire [10:0] buffer_11_361; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_74444; // @[Modules.scala 65:57:@27672.4]
  wire [10:0] _T_74445; // @[Modules.scala 65:57:@27673.4]
  wire [10:0] buffer_11_572; // @[Modules.scala 65:57:@27674.4]
  wire [11:0] _T_74471; // @[Modules.scala 65:57:@27708.4]
  wire [10:0] _T_74472; // @[Modules.scala 65:57:@27709.4]
  wire [10:0] buffer_11_581; // @[Modules.scala 65:57:@27710.4]
  wire [11:0] _T_74492; // @[Modules.scala 68:83:@27736.4]
  wire [10:0] _T_74493; // @[Modules.scala 68:83:@27737.4]
  wire [10:0] buffer_11_588; // @[Modules.scala 68:83:@27738.4]
  wire [11:0] _T_74495; // @[Modules.scala 68:83:@27740.4]
  wire [10:0] _T_74496; // @[Modules.scala 68:83:@27741.4]
  wire [10:0] buffer_11_589; // @[Modules.scala 68:83:@27742.4]
  wire [11:0] _T_74498; // @[Modules.scala 68:83:@27744.4]
  wire [10:0] _T_74499; // @[Modules.scala 68:83:@27745.4]
  wire [10:0] buffer_11_590; // @[Modules.scala 68:83:@27746.4]
  wire [11:0] _T_74501; // @[Modules.scala 68:83:@27748.4]
  wire [10:0] _T_74502; // @[Modules.scala 68:83:@27749.4]
  wire [10:0] buffer_11_591; // @[Modules.scala 68:83:@27750.4]
  wire [11:0] _T_74504; // @[Modules.scala 68:83:@27752.4]
  wire [10:0] _T_74505; // @[Modules.scala 68:83:@27753.4]
  wire [10:0] buffer_11_592; // @[Modules.scala 68:83:@27754.4]
  wire [11:0] _T_74507; // @[Modules.scala 68:83:@27756.4]
  wire [10:0] _T_74508; // @[Modules.scala 68:83:@27757.4]
  wire [10:0] buffer_11_593; // @[Modules.scala 68:83:@27758.4]
  wire [11:0] _T_74510; // @[Modules.scala 68:83:@27760.4]
  wire [10:0] _T_74511; // @[Modules.scala 68:83:@27761.4]
  wire [10:0] buffer_11_594; // @[Modules.scala 68:83:@27762.4]
  wire [11:0] _T_74513; // @[Modules.scala 68:83:@27764.4]
  wire [10:0] _T_74514; // @[Modules.scala 68:83:@27765.4]
  wire [10:0] buffer_11_595; // @[Modules.scala 68:83:@27766.4]
  wire [11:0] _T_74516; // @[Modules.scala 68:83:@27768.4]
  wire [10:0] _T_74517; // @[Modules.scala 68:83:@27769.4]
  wire [10:0] buffer_11_596; // @[Modules.scala 68:83:@27770.4]
  wire [11:0] _T_74522; // @[Modules.scala 68:83:@27776.4]
  wire [10:0] _T_74523; // @[Modules.scala 68:83:@27777.4]
  wire [10:0] buffer_11_598; // @[Modules.scala 68:83:@27778.4]
  wire [11:0] _T_74525; // @[Modules.scala 68:83:@27780.4]
  wire [10:0] _T_74526; // @[Modules.scala 68:83:@27781.4]
  wire [10:0] buffer_11_599; // @[Modules.scala 68:83:@27782.4]
  wire [11:0] _T_74537; // @[Modules.scala 68:83:@27796.4]
  wire [10:0] _T_74538; // @[Modules.scala 68:83:@27797.4]
  wire [10:0] buffer_11_603; // @[Modules.scala 68:83:@27798.4]
  wire [11:0] _T_74540; // @[Modules.scala 68:83:@27800.4]
  wire [10:0] _T_74541; // @[Modules.scala 68:83:@27801.4]
  wire [10:0] buffer_11_604; // @[Modules.scala 68:83:@27802.4]
  wire [11:0] _T_74543; // @[Modules.scala 68:83:@27804.4]
  wire [10:0] _T_74544; // @[Modules.scala 68:83:@27805.4]
  wire [10:0] buffer_11_605; // @[Modules.scala 68:83:@27806.4]
  wire [11:0] _T_74549; // @[Modules.scala 68:83:@27812.4]
  wire [10:0] _T_74550; // @[Modules.scala 68:83:@27813.4]
  wire [10:0] buffer_11_607; // @[Modules.scala 68:83:@27814.4]
  wire [11:0] _T_74552; // @[Modules.scala 68:83:@27816.4]
  wire [10:0] _T_74553; // @[Modules.scala 68:83:@27817.4]
  wire [10:0] buffer_11_608; // @[Modules.scala 68:83:@27818.4]
  wire [11:0] _T_74555; // @[Modules.scala 68:83:@27820.4]
  wire [10:0] _T_74556; // @[Modules.scala 68:83:@27821.4]
  wire [10:0] buffer_11_609; // @[Modules.scala 68:83:@27822.4]
  wire [11:0] _T_74558; // @[Modules.scala 68:83:@27824.4]
  wire [10:0] _T_74559; // @[Modules.scala 68:83:@27825.4]
  wire [10:0] buffer_11_610; // @[Modules.scala 68:83:@27826.4]
  wire [11:0] _T_74561; // @[Modules.scala 68:83:@27828.4]
  wire [10:0] _T_74562; // @[Modules.scala 68:83:@27829.4]
  wire [10:0] buffer_11_611; // @[Modules.scala 68:83:@27830.4]
  wire [11:0] _T_74564; // @[Modules.scala 68:83:@27832.4]
  wire [10:0] _T_74565; // @[Modules.scala 68:83:@27833.4]
  wire [10:0] buffer_11_612; // @[Modules.scala 68:83:@27834.4]
  wire [11:0] _T_74567; // @[Modules.scala 68:83:@27836.4]
  wire [10:0] _T_74568; // @[Modules.scala 68:83:@27837.4]
  wire [10:0] buffer_11_613; // @[Modules.scala 68:83:@27838.4]
  wire [11:0] _T_74570; // @[Modules.scala 68:83:@27840.4]
  wire [10:0] _T_74571; // @[Modules.scala 68:83:@27841.4]
  wire [10:0] buffer_11_614; // @[Modules.scala 68:83:@27842.4]
  wire [11:0] _T_74576; // @[Modules.scala 68:83:@27848.4]
  wire [10:0] _T_74577; // @[Modules.scala 68:83:@27849.4]
  wire [10:0] buffer_11_616; // @[Modules.scala 68:83:@27850.4]
  wire [11:0] _T_74579; // @[Modules.scala 68:83:@27852.4]
  wire [10:0] _T_74580; // @[Modules.scala 68:83:@27853.4]
  wire [10:0] buffer_11_617; // @[Modules.scala 68:83:@27854.4]
  wire [11:0] _T_74582; // @[Modules.scala 68:83:@27856.4]
  wire [10:0] _T_74583; // @[Modules.scala 68:83:@27857.4]
  wire [10:0] buffer_11_618; // @[Modules.scala 68:83:@27858.4]
  wire [11:0] _T_74585; // @[Modules.scala 68:83:@27860.4]
  wire [10:0] _T_74586; // @[Modules.scala 68:83:@27861.4]
  wire [10:0] buffer_11_619; // @[Modules.scala 68:83:@27862.4]
  wire [11:0] _T_74588; // @[Modules.scala 68:83:@27864.4]
  wire [10:0] _T_74589; // @[Modules.scala 68:83:@27865.4]
  wire [10:0] buffer_11_620; // @[Modules.scala 68:83:@27866.4]
  wire [11:0] _T_74591; // @[Modules.scala 68:83:@27868.4]
  wire [10:0] _T_74592; // @[Modules.scala 68:83:@27869.4]
  wire [10:0] buffer_11_621; // @[Modules.scala 68:83:@27870.4]
  wire [11:0] _T_74597; // @[Modules.scala 68:83:@27876.4]
  wire [10:0] _T_74598; // @[Modules.scala 68:83:@27877.4]
  wire [10:0] buffer_11_623; // @[Modules.scala 68:83:@27878.4]
  wire [11:0] _T_74600; // @[Modules.scala 68:83:@27880.4]
  wire [10:0] _T_74601; // @[Modules.scala 68:83:@27881.4]
  wire [10:0] buffer_11_624; // @[Modules.scala 68:83:@27882.4]
  wire [11:0] _T_74609; // @[Modules.scala 68:83:@27892.4]
  wire [10:0] _T_74610; // @[Modules.scala 68:83:@27893.4]
  wire [10:0] buffer_11_627; // @[Modules.scala 68:83:@27894.4]
  wire [11:0] _T_74612; // @[Modules.scala 68:83:@27896.4]
  wire [10:0] _T_74613; // @[Modules.scala 68:83:@27897.4]
  wire [10:0] buffer_11_628; // @[Modules.scala 68:83:@27898.4]
  wire [11:0] _T_74624; // @[Modules.scala 68:83:@27912.4]
  wire [10:0] _T_74625; // @[Modules.scala 68:83:@27913.4]
  wire [10:0] buffer_11_632; // @[Modules.scala 68:83:@27914.4]
  wire [11:0] _T_74627; // @[Modules.scala 68:83:@27916.4]
  wire [10:0] _T_74628; // @[Modules.scala 68:83:@27917.4]
  wire [10:0] buffer_11_633; // @[Modules.scala 68:83:@27918.4]
  wire [11:0] _T_74630; // @[Modules.scala 68:83:@27920.4]
  wire [10:0] _T_74631; // @[Modules.scala 68:83:@27921.4]
  wire [10:0] buffer_11_634; // @[Modules.scala 68:83:@27922.4]
  wire [11:0] _T_74633; // @[Modules.scala 68:83:@27924.4]
  wire [10:0] _T_74634; // @[Modules.scala 68:83:@27925.4]
  wire [10:0] buffer_11_635; // @[Modules.scala 68:83:@27926.4]
  wire [11:0] _T_74636; // @[Modules.scala 68:83:@27928.4]
  wire [10:0] _T_74637; // @[Modules.scala 68:83:@27929.4]
  wire [10:0] buffer_11_636; // @[Modules.scala 68:83:@27930.4]
  wire [11:0] _T_74642; // @[Modules.scala 68:83:@27936.4]
  wire [10:0] _T_74643; // @[Modules.scala 68:83:@27937.4]
  wire [10:0] buffer_11_638; // @[Modules.scala 68:83:@27938.4]
  wire [11:0] _T_74648; // @[Modules.scala 68:83:@27944.4]
  wire [10:0] _T_74649; // @[Modules.scala 68:83:@27945.4]
  wire [10:0] buffer_11_640; // @[Modules.scala 68:83:@27946.4]
  wire [11:0] _T_74651; // @[Modules.scala 68:83:@27948.4]
  wire [10:0] _T_74652; // @[Modules.scala 68:83:@27949.4]
  wire [10:0] buffer_11_641; // @[Modules.scala 68:83:@27950.4]
  wire [11:0] _T_74654; // @[Modules.scala 68:83:@27952.4]
  wire [10:0] _T_74655; // @[Modules.scala 68:83:@27953.4]
  wire [10:0] buffer_11_642; // @[Modules.scala 68:83:@27954.4]
  wire [11:0] _T_74660; // @[Modules.scala 68:83:@27960.4]
  wire [10:0] _T_74661; // @[Modules.scala 68:83:@27961.4]
  wire [10:0] buffer_11_644; // @[Modules.scala 68:83:@27962.4]
  wire [11:0] _T_74663; // @[Modules.scala 68:83:@27964.4]
  wire [10:0] _T_74664; // @[Modules.scala 68:83:@27965.4]
  wire [10:0] buffer_11_645; // @[Modules.scala 68:83:@27966.4]
  wire [11:0] _T_74666; // @[Modules.scala 68:83:@27968.4]
  wire [10:0] _T_74667; // @[Modules.scala 68:83:@27969.4]
  wire [10:0] buffer_11_646; // @[Modules.scala 68:83:@27970.4]
  wire [11:0] _T_74669; // @[Modules.scala 68:83:@27972.4]
  wire [10:0] _T_74670; // @[Modules.scala 68:83:@27973.4]
  wire [10:0] buffer_11_647; // @[Modules.scala 68:83:@27974.4]
  wire [11:0] _T_74672; // @[Modules.scala 68:83:@27976.4]
  wire [10:0] _T_74673; // @[Modules.scala 68:83:@27977.4]
  wire [10:0] buffer_11_648; // @[Modules.scala 68:83:@27978.4]
  wire [11:0] _T_74675; // @[Modules.scala 68:83:@27980.4]
  wire [10:0] _T_74676; // @[Modules.scala 68:83:@27981.4]
  wire [10:0] buffer_11_649; // @[Modules.scala 68:83:@27982.4]
  wire [11:0] _T_74678; // @[Modules.scala 68:83:@27984.4]
  wire [10:0] _T_74679; // @[Modules.scala 68:83:@27985.4]
  wire [10:0] buffer_11_650; // @[Modules.scala 68:83:@27986.4]
  wire [11:0] _T_74681; // @[Modules.scala 68:83:@27988.4]
  wire [10:0] _T_74682; // @[Modules.scala 68:83:@27989.4]
  wire [10:0] buffer_11_651; // @[Modules.scala 68:83:@27990.4]
  wire [11:0] _T_74684; // @[Modules.scala 68:83:@27992.4]
  wire [10:0] _T_74685; // @[Modules.scala 68:83:@27993.4]
  wire [10:0] buffer_11_652; // @[Modules.scala 68:83:@27994.4]
  wire [11:0] _T_74687; // @[Modules.scala 68:83:@27996.4]
  wire [10:0] _T_74688; // @[Modules.scala 68:83:@27997.4]
  wire [10:0] buffer_11_653; // @[Modules.scala 68:83:@27998.4]
  wire [11:0] _T_74693; // @[Modules.scala 68:83:@28004.4]
  wire [10:0] _T_74694; // @[Modules.scala 68:83:@28005.4]
  wire [10:0] buffer_11_655; // @[Modules.scala 68:83:@28006.4]
  wire [11:0] _T_74696; // @[Modules.scala 68:83:@28008.4]
  wire [10:0] _T_74697; // @[Modules.scala 68:83:@28009.4]
  wire [10:0] buffer_11_656; // @[Modules.scala 68:83:@28010.4]
  wire [11:0] _T_74699; // @[Modules.scala 68:83:@28012.4]
  wire [10:0] _T_74700; // @[Modules.scala 68:83:@28013.4]
  wire [10:0] buffer_11_657; // @[Modules.scala 68:83:@28014.4]
  wire [11:0] _T_74702; // @[Modules.scala 68:83:@28016.4]
  wire [10:0] _T_74703; // @[Modules.scala 68:83:@28017.4]
  wire [10:0] buffer_11_658; // @[Modules.scala 68:83:@28018.4]
  wire [11:0] _T_74705; // @[Modules.scala 68:83:@28020.4]
  wire [10:0] _T_74706; // @[Modules.scala 68:83:@28021.4]
  wire [10:0] buffer_11_659; // @[Modules.scala 68:83:@28022.4]
  wire [11:0] _T_74708; // @[Modules.scala 68:83:@28024.4]
  wire [10:0] _T_74709; // @[Modules.scala 68:83:@28025.4]
  wire [10:0] buffer_11_660; // @[Modules.scala 68:83:@28026.4]
  wire [11:0] _T_74711; // @[Modules.scala 68:83:@28028.4]
  wire [10:0] _T_74712; // @[Modules.scala 68:83:@28029.4]
  wire [10:0] buffer_11_661; // @[Modules.scala 68:83:@28030.4]
  wire [11:0] _T_74714; // @[Modules.scala 68:83:@28032.4]
  wire [10:0] _T_74715; // @[Modules.scala 68:83:@28033.4]
  wire [10:0] buffer_11_662; // @[Modules.scala 68:83:@28034.4]
  wire [11:0] _T_74717; // @[Modules.scala 68:83:@28036.4]
  wire [10:0] _T_74718; // @[Modules.scala 68:83:@28037.4]
  wire [10:0] buffer_11_663; // @[Modules.scala 68:83:@28038.4]
  wire [11:0] _T_74720; // @[Modules.scala 68:83:@28040.4]
  wire [10:0] _T_74721; // @[Modules.scala 68:83:@28041.4]
  wire [10:0] buffer_11_664; // @[Modules.scala 68:83:@28042.4]
  wire [11:0] _T_74723; // @[Modules.scala 68:83:@28044.4]
  wire [10:0] _T_74724; // @[Modules.scala 68:83:@28045.4]
  wire [10:0] buffer_11_665; // @[Modules.scala 68:83:@28046.4]
  wire [11:0] _T_74726; // @[Modules.scala 68:83:@28048.4]
  wire [10:0] _T_74727; // @[Modules.scala 68:83:@28049.4]
  wire [10:0] buffer_11_666; // @[Modules.scala 68:83:@28050.4]
  wire [11:0] _T_74732; // @[Modules.scala 68:83:@28056.4]
  wire [10:0] _T_74733; // @[Modules.scala 68:83:@28057.4]
  wire [10:0] buffer_11_668; // @[Modules.scala 68:83:@28058.4]
  wire [11:0] _T_74735; // @[Modules.scala 68:83:@28060.4]
  wire [10:0] _T_74736; // @[Modules.scala 68:83:@28061.4]
  wire [10:0] buffer_11_669; // @[Modules.scala 68:83:@28062.4]
  wire [11:0] _T_74738; // @[Modules.scala 68:83:@28064.4]
  wire [10:0] _T_74739; // @[Modules.scala 68:83:@28065.4]
  wire [10:0] buffer_11_670; // @[Modules.scala 68:83:@28066.4]
  wire [11:0] _T_74741; // @[Modules.scala 68:83:@28068.4]
  wire [10:0] _T_74742; // @[Modules.scala 68:83:@28069.4]
  wire [10:0] buffer_11_671; // @[Modules.scala 68:83:@28070.4]
  wire [11:0] _T_74750; // @[Modules.scala 68:83:@28080.4]
  wire [10:0] _T_74751; // @[Modules.scala 68:83:@28081.4]
  wire [10:0] buffer_11_674; // @[Modules.scala 68:83:@28082.4]
  wire [11:0] _T_74753; // @[Modules.scala 68:83:@28084.4]
  wire [10:0] _T_74754; // @[Modules.scala 68:83:@28085.4]
  wire [10:0] buffer_11_675; // @[Modules.scala 68:83:@28086.4]
  wire [11:0] _T_74762; // @[Modules.scala 68:83:@28096.4]
  wire [10:0] _T_74763; // @[Modules.scala 68:83:@28097.4]
  wire [10:0] buffer_11_678; // @[Modules.scala 68:83:@28098.4]
  wire [11:0] _T_74774; // @[Modules.scala 68:83:@28112.4]
  wire [10:0] _T_74775; // @[Modules.scala 68:83:@28113.4]
  wire [10:0] buffer_11_682; // @[Modules.scala 68:83:@28114.4]
  wire [11:0] _T_74786; // @[Modules.scala 71:109:@28128.4]
  wire [10:0] _T_74787; // @[Modules.scala 71:109:@28129.4]
  wire [10:0] buffer_11_686; // @[Modules.scala 71:109:@28130.4]
  wire [11:0] _T_74789; // @[Modules.scala 71:109:@28132.4]
  wire [10:0] _T_74790; // @[Modules.scala 71:109:@28133.4]
  wire [10:0] buffer_11_687; // @[Modules.scala 71:109:@28134.4]
  wire [11:0] _T_74792; // @[Modules.scala 71:109:@28136.4]
  wire [10:0] _T_74793; // @[Modules.scala 71:109:@28137.4]
  wire [10:0] buffer_11_688; // @[Modules.scala 71:109:@28138.4]
  wire [11:0] _T_74795; // @[Modules.scala 71:109:@28140.4]
  wire [10:0] _T_74796; // @[Modules.scala 71:109:@28141.4]
  wire [10:0] buffer_11_689; // @[Modules.scala 71:109:@28142.4]
  wire [11:0] _T_74798; // @[Modules.scala 71:109:@28144.4]
  wire [10:0] _T_74799; // @[Modules.scala 71:109:@28145.4]
  wire [10:0] buffer_11_690; // @[Modules.scala 71:109:@28146.4]
  wire [11:0] _T_74801; // @[Modules.scala 71:109:@28148.4]
  wire [10:0] _T_74802; // @[Modules.scala 71:109:@28149.4]
  wire [10:0] buffer_11_691; // @[Modules.scala 71:109:@28150.4]
  wire [11:0] _T_74807; // @[Modules.scala 71:109:@28156.4]
  wire [10:0] _T_74808; // @[Modules.scala 71:109:@28157.4]
  wire [10:0] buffer_11_693; // @[Modules.scala 71:109:@28158.4]
  wire [11:0] _T_74810; // @[Modules.scala 71:109:@28160.4]
  wire [10:0] _T_74811; // @[Modules.scala 71:109:@28161.4]
  wire [10:0] buffer_11_694; // @[Modules.scala 71:109:@28162.4]
  wire [11:0] _T_74813; // @[Modules.scala 71:109:@28164.4]
  wire [10:0] _T_74814; // @[Modules.scala 71:109:@28165.4]
  wire [10:0] buffer_11_695; // @[Modules.scala 71:109:@28166.4]
  wire [11:0] _T_74816; // @[Modules.scala 71:109:@28168.4]
  wire [10:0] _T_74817; // @[Modules.scala 71:109:@28169.4]
  wire [10:0] buffer_11_696; // @[Modules.scala 71:109:@28170.4]
  wire [11:0] _T_74819; // @[Modules.scala 71:109:@28172.4]
  wire [10:0] _T_74820; // @[Modules.scala 71:109:@28173.4]
  wire [10:0] buffer_11_697; // @[Modules.scala 71:109:@28174.4]
  wire [11:0] _T_74822; // @[Modules.scala 71:109:@28176.4]
  wire [10:0] _T_74823; // @[Modules.scala 71:109:@28177.4]
  wire [10:0] buffer_11_698; // @[Modules.scala 71:109:@28178.4]
  wire [11:0] _T_74825; // @[Modules.scala 71:109:@28180.4]
  wire [10:0] _T_74826; // @[Modules.scala 71:109:@28181.4]
  wire [10:0] buffer_11_699; // @[Modules.scala 71:109:@28182.4]
  wire [11:0] _T_74828; // @[Modules.scala 71:109:@28184.4]
  wire [10:0] _T_74829; // @[Modules.scala 71:109:@28185.4]
  wire [10:0] buffer_11_700; // @[Modules.scala 71:109:@28186.4]
  wire [11:0] _T_74831; // @[Modules.scala 71:109:@28188.4]
  wire [10:0] _T_74832; // @[Modules.scala 71:109:@28189.4]
  wire [10:0] buffer_11_701; // @[Modules.scala 71:109:@28190.4]
  wire [11:0] _T_74834; // @[Modules.scala 71:109:@28192.4]
  wire [10:0] _T_74835; // @[Modules.scala 71:109:@28193.4]
  wire [10:0] buffer_11_702; // @[Modules.scala 71:109:@28194.4]
  wire [11:0] _T_74837; // @[Modules.scala 71:109:@28196.4]
  wire [10:0] _T_74838; // @[Modules.scala 71:109:@28197.4]
  wire [10:0] buffer_11_703; // @[Modules.scala 71:109:@28198.4]
  wire [11:0] _T_74840; // @[Modules.scala 71:109:@28200.4]
  wire [10:0] _T_74841; // @[Modules.scala 71:109:@28201.4]
  wire [10:0] buffer_11_704; // @[Modules.scala 71:109:@28202.4]
  wire [11:0] _T_74843; // @[Modules.scala 71:109:@28204.4]
  wire [10:0] _T_74844; // @[Modules.scala 71:109:@28205.4]
  wire [10:0] buffer_11_705; // @[Modules.scala 71:109:@28206.4]
  wire [11:0] _T_74846; // @[Modules.scala 71:109:@28208.4]
  wire [10:0] _T_74847; // @[Modules.scala 71:109:@28209.4]
  wire [10:0] buffer_11_706; // @[Modules.scala 71:109:@28210.4]
  wire [11:0] _T_74852; // @[Modules.scala 71:109:@28216.4]
  wire [10:0] _T_74853; // @[Modules.scala 71:109:@28217.4]
  wire [10:0] buffer_11_708; // @[Modules.scala 71:109:@28218.4]
  wire [11:0] _T_74855; // @[Modules.scala 71:109:@28220.4]
  wire [10:0] _T_74856; // @[Modules.scala 71:109:@28221.4]
  wire [10:0] buffer_11_709; // @[Modules.scala 71:109:@28222.4]
  wire [11:0] _T_74858; // @[Modules.scala 71:109:@28224.4]
  wire [10:0] _T_74859; // @[Modules.scala 71:109:@28225.4]
  wire [10:0] buffer_11_710; // @[Modules.scala 71:109:@28226.4]
  wire [11:0] _T_74861; // @[Modules.scala 71:109:@28228.4]
  wire [10:0] _T_74862; // @[Modules.scala 71:109:@28229.4]
  wire [10:0] buffer_11_711; // @[Modules.scala 71:109:@28230.4]
  wire [11:0] _T_74864; // @[Modules.scala 71:109:@28232.4]
  wire [10:0] _T_74865; // @[Modules.scala 71:109:@28233.4]
  wire [10:0] buffer_11_712; // @[Modules.scala 71:109:@28234.4]
  wire [11:0] _T_74867; // @[Modules.scala 71:109:@28236.4]
  wire [10:0] _T_74868; // @[Modules.scala 71:109:@28237.4]
  wire [10:0] buffer_11_713; // @[Modules.scala 71:109:@28238.4]
  wire [11:0] _T_74870; // @[Modules.scala 71:109:@28240.4]
  wire [10:0] _T_74871; // @[Modules.scala 71:109:@28241.4]
  wire [10:0] buffer_11_714; // @[Modules.scala 71:109:@28242.4]
  wire [11:0] _T_74873; // @[Modules.scala 71:109:@28244.4]
  wire [10:0] _T_74874; // @[Modules.scala 71:109:@28245.4]
  wire [10:0] buffer_11_715; // @[Modules.scala 71:109:@28246.4]
  wire [11:0] _T_74876; // @[Modules.scala 71:109:@28248.4]
  wire [10:0] _T_74877; // @[Modules.scala 71:109:@28249.4]
  wire [10:0] buffer_11_716; // @[Modules.scala 71:109:@28250.4]
  wire [11:0] _T_74879; // @[Modules.scala 71:109:@28252.4]
  wire [10:0] _T_74880; // @[Modules.scala 71:109:@28253.4]
  wire [10:0] buffer_11_717; // @[Modules.scala 71:109:@28254.4]
  wire [11:0] _T_74882; // @[Modules.scala 71:109:@28256.4]
  wire [10:0] _T_74883; // @[Modules.scala 71:109:@28257.4]
  wire [10:0] buffer_11_718; // @[Modules.scala 71:109:@28258.4]
  wire [11:0] _T_74885; // @[Modules.scala 71:109:@28260.4]
  wire [10:0] _T_74886; // @[Modules.scala 71:109:@28261.4]
  wire [10:0] buffer_11_719; // @[Modules.scala 71:109:@28262.4]
  wire [11:0] _T_74888; // @[Modules.scala 71:109:@28264.4]
  wire [10:0] _T_74889; // @[Modules.scala 71:109:@28265.4]
  wire [10:0] buffer_11_720; // @[Modules.scala 71:109:@28266.4]
  wire [11:0] _T_74891; // @[Modules.scala 71:109:@28268.4]
  wire [10:0] _T_74892; // @[Modules.scala 71:109:@28269.4]
  wire [10:0] buffer_11_721; // @[Modules.scala 71:109:@28270.4]
  wire [11:0] _T_74894; // @[Modules.scala 71:109:@28272.4]
  wire [10:0] _T_74895; // @[Modules.scala 71:109:@28273.4]
  wire [10:0] buffer_11_722; // @[Modules.scala 71:109:@28274.4]
  wire [11:0] _T_74897; // @[Modules.scala 71:109:@28276.4]
  wire [10:0] _T_74898; // @[Modules.scala 71:109:@28277.4]
  wire [10:0] buffer_11_723; // @[Modules.scala 71:109:@28278.4]
  wire [11:0] _T_74900; // @[Modules.scala 71:109:@28280.4]
  wire [10:0] _T_74901; // @[Modules.scala 71:109:@28281.4]
  wire [10:0] buffer_11_724; // @[Modules.scala 71:109:@28282.4]
  wire [11:0] _T_74903; // @[Modules.scala 71:109:@28284.4]
  wire [10:0] _T_74904; // @[Modules.scala 71:109:@28285.4]
  wire [10:0] buffer_11_725; // @[Modules.scala 71:109:@28286.4]
  wire [11:0] _T_74906; // @[Modules.scala 71:109:@28288.4]
  wire [10:0] _T_74907; // @[Modules.scala 71:109:@28289.4]
  wire [10:0] buffer_11_726; // @[Modules.scala 71:109:@28290.4]
  wire [11:0] _T_74909; // @[Modules.scala 71:109:@28292.4]
  wire [10:0] _T_74910; // @[Modules.scala 71:109:@28293.4]
  wire [10:0] buffer_11_727; // @[Modules.scala 71:109:@28294.4]
  wire [11:0] _T_74912; // @[Modules.scala 71:109:@28296.4]
  wire [10:0] _T_74913; // @[Modules.scala 71:109:@28297.4]
  wire [10:0] buffer_11_728; // @[Modules.scala 71:109:@28298.4]
  wire [11:0] _T_74915; // @[Modules.scala 71:109:@28300.4]
  wire [10:0] _T_74916; // @[Modules.scala 71:109:@28301.4]
  wire [10:0] buffer_11_729; // @[Modules.scala 71:109:@28302.4]
  wire [11:0] _T_74921; // @[Modules.scala 71:109:@28308.4]
  wire [10:0] _T_74922; // @[Modules.scala 71:109:@28309.4]
  wire [10:0] buffer_11_731; // @[Modules.scala 71:109:@28310.4]
  wire [11:0] _T_74927; // @[Modules.scala 71:109:@28316.4]
  wire [10:0] _T_74928; // @[Modules.scala 71:109:@28317.4]
  wire [10:0] buffer_11_733; // @[Modules.scala 71:109:@28318.4]
  wire [11:0] _T_74933; // @[Modules.scala 78:156:@28325.4]
  wire [10:0] _T_74934; // @[Modules.scala 78:156:@28326.4]
  wire [10:0] buffer_11_736; // @[Modules.scala 78:156:@28327.4]
  wire [11:0] _T_74936; // @[Modules.scala 78:156:@28329.4]
  wire [10:0] _T_74937; // @[Modules.scala 78:156:@28330.4]
  wire [10:0] buffer_11_737; // @[Modules.scala 78:156:@28331.4]
  wire [11:0] _T_74939; // @[Modules.scala 78:156:@28333.4]
  wire [10:0] _T_74940; // @[Modules.scala 78:156:@28334.4]
  wire [10:0] buffer_11_738; // @[Modules.scala 78:156:@28335.4]
  wire [11:0] _T_74942; // @[Modules.scala 78:156:@28337.4]
  wire [10:0] _T_74943; // @[Modules.scala 78:156:@28338.4]
  wire [10:0] buffer_11_739; // @[Modules.scala 78:156:@28339.4]
  wire [11:0] _T_74945; // @[Modules.scala 78:156:@28341.4]
  wire [10:0] _T_74946; // @[Modules.scala 78:156:@28342.4]
  wire [10:0] buffer_11_740; // @[Modules.scala 78:156:@28343.4]
  wire [11:0] _T_74948; // @[Modules.scala 78:156:@28345.4]
  wire [10:0] _T_74949; // @[Modules.scala 78:156:@28346.4]
  wire [10:0] buffer_11_741; // @[Modules.scala 78:156:@28347.4]
  wire [11:0] _T_74951; // @[Modules.scala 78:156:@28349.4]
  wire [10:0] _T_74952; // @[Modules.scala 78:156:@28350.4]
  wire [10:0] buffer_11_742; // @[Modules.scala 78:156:@28351.4]
  wire [11:0] _T_74954; // @[Modules.scala 78:156:@28353.4]
  wire [10:0] _T_74955; // @[Modules.scala 78:156:@28354.4]
  wire [10:0] buffer_11_743; // @[Modules.scala 78:156:@28355.4]
  wire [11:0] _T_74957; // @[Modules.scala 78:156:@28357.4]
  wire [10:0] _T_74958; // @[Modules.scala 78:156:@28358.4]
  wire [10:0] buffer_11_744; // @[Modules.scala 78:156:@28359.4]
  wire [11:0] _T_74960; // @[Modules.scala 78:156:@28361.4]
  wire [10:0] _T_74961; // @[Modules.scala 78:156:@28362.4]
  wire [10:0] buffer_11_745; // @[Modules.scala 78:156:@28363.4]
  wire [11:0] _T_74963; // @[Modules.scala 78:156:@28365.4]
  wire [10:0] _T_74964; // @[Modules.scala 78:156:@28366.4]
  wire [10:0] buffer_11_746; // @[Modules.scala 78:156:@28367.4]
  wire [11:0] _T_74966; // @[Modules.scala 78:156:@28369.4]
  wire [10:0] _T_74967; // @[Modules.scala 78:156:@28370.4]
  wire [10:0] buffer_11_747; // @[Modules.scala 78:156:@28371.4]
  wire [11:0] _T_74969; // @[Modules.scala 78:156:@28373.4]
  wire [10:0] _T_74970; // @[Modules.scala 78:156:@28374.4]
  wire [10:0] buffer_11_748; // @[Modules.scala 78:156:@28375.4]
  wire [11:0] _T_74972; // @[Modules.scala 78:156:@28377.4]
  wire [10:0] _T_74973; // @[Modules.scala 78:156:@28378.4]
  wire [10:0] buffer_11_749; // @[Modules.scala 78:156:@28379.4]
  wire [11:0] _T_74975; // @[Modules.scala 78:156:@28381.4]
  wire [10:0] _T_74976; // @[Modules.scala 78:156:@28382.4]
  wire [10:0] buffer_11_750; // @[Modules.scala 78:156:@28383.4]
  wire [11:0] _T_74978; // @[Modules.scala 78:156:@28385.4]
  wire [10:0] _T_74979; // @[Modules.scala 78:156:@28386.4]
  wire [10:0] buffer_11_751; // @[Modules.scala 78:156:@28387.4]
  wire [11:0] _T_74981; // @[Modules.scala 78:156:@28389.4]
  wire [10:0] _T_74982; // @[Modules.scala 78:156:@28390.4]
  wire [10:0] buffer_11_752; // @[Modules.scala 78:156:@28391.4]
  wire [11:0] _T_74984; // @[Modules.scala 78:156:@28393.4]
  wire [10:0] _T_74985; // @[Modules.scala 78:156:@28394.4]
  wire [10:0] buffer_11_753; // @[Modules.scala 78:156:@28395.4]
  wire [11:0] _T_74987; // @[Modules.scala 78:156:@28397.4]
  wire [10:0] _T_74988; // @[Modules.scala 78:156:@28398.4]
  wire [10:0] buffer_11_754; // @[Modules.scala 78:156:@28399.4]
  wire [11:0] _T_74990; // @[Modules.scala 78:156:@28401.4]
  wire [10:0] _T_74991; // @[Modules.scala 78:156:@28402.4]
  wire [10:0] buffer_11_755; // @[Modules.scala 78:156:@28403.4]
  wire [11:0] _T_74993; // @[Modules.scala 78:156:@28405.4]
  wire [10:0] _T_74994; // @[Modules.scala 78:156:@28406.4]
  wire [10:0] buffer_11_756; // @[Modules.scala 78:156:@28407.4]
  wire [11:0] _T_74996; // @[Modules.scala 78:156:@28409.4]
  wire [10:0] _T_74997; // @[Modules.scala 78:156:@28410.4]
  wire [10:0] buffer_11_757; // @[Modules.scala 78:156:@28411.4]
  wire [11:0] _T_74999; // @[Modules.scala 78:156:@28413.4]
  wire [10:0] _T_75000; // @[Modules.scala 78:156:@28414.4]
  wire [10:0] buffer_11_758; // @[Modules.scala 78:156:@28415.4]
  wire [11:0] _T_75002; // @[Modules.scala 78:156:@28417.4]
  wire [10:0] _T_75003; // @[Modules.scala 78:156:@28418.4]
  wire [10:0] buffer_11_759; // @[Modules.scala 78:156:@28419.4]
  wire [11:0] _T_75005; // @[Modules.scala 78:156:@28421.4]
  wire [10:0] _T_75006; // @[Modules.scala 78:156:@28422.4]
  wire [10:0] buffer_11_760; // @[Modules.scala 78:156:@28423.4]
  wire [11:0] _T_75008; // @[Modules.scala 78:156:@28425.4]
  wire [10:0] _T_75009; // @[Modules.scala 78:156:@28426.4]
  wire [10:0] buffer_11_761; // @[Modules.scala 78:156:@28427.4]
  wire [11:0] _T_75011; // @[Modules.scala 78:156:@28429.4]
  wire [10:0] _T_75012; // @[Modules.scala 78:156:@28430.4]
  wire [10:0] buffer_11_762; // @[Modules.scala 78:156:@28431.4]
  wire [11:0] _T_75014; // @[Modules.scala 78:156:@28433.4]
  wire [10:0] _T_75015; // @[Modules.scala 78:156:@28434.4]
  wire [10:0] buffer_11_763; // @[Modules.scala 78:156:@28435.4]
  wire [11:0] _T_75017; // @[Modules.scala 78:156:@28437.4]
  wire [10:0] _T_75018; // @[Modules.scala 78:156:@28438.4]
  wire [10:0] buffer_11_764; // @[Modules.scala 78:156:@28439.4]
  wire [11:0] _T_75020; // @[Modules.scala 78:156:@28441.4]
  wire [10:0] _T_75021; // @[Modules.scala 78:156:@28442.4]
  wire [10:0] buffer_11_765; // @[Modules.scala 78:156:@28443.4]
  wire [11:0] _T_75023; // @[Modules.scala 78:156:@28445.4]
  wire [10:0] _T_75024; // @[Modules.scala 78:156:@28446.4]
  wire [10:0] buffer_11_766; // @[Modules.scala 78:156:@28447.4]
  wire [11:0] _T_75026; // @[Modules.scala 78:156:@28449.4]
  wire [10:0] _T_75027; // @[Modules.scala 78:156:@28450.4]
  wire [10:0] buffer_11_767; // @[Modules.scala 78:156:@28451.4]
  wire [11:0] _T_75029; // @[Modules.scala 78:156:@28453.4]
  wire [10:0] _T_75030; // @[Modules.scala 78:156:@28454.4]
  wire [10:0] buffer_11_768; // @[Modules.scala 78:156:@28455.4]
  wire [11:0] _T_75032; // @[Modules.scala 78:156:@28457.4]
  wire [10:0] _T_75033; // @[Modules.scala 78:156:@28458.4]
  wire [10:0] buffer_11_769; // @[Modules.scala 78:156:@28459.4]
  wire [11:0] _T_75035; // @[Modules.scala 78:156:@28461.4]
  wire [10:0] _T_75036; // @[Modules.scala 78:156:@28462.4]
  wire [10:0] buffer_11_770; // @[Modules.scala 78:156:@28463.4]
  wire [11:0] _T_75038; // @[Modules.scala 78:156:@28465.4]
  wire [10:0] _T_75039; // @[Modules.scala 78:156:@28466.4]
  wire [10:0] buffer_11_771; // @[Modules.scala 78:156:@28467.4]
  wire [11:0] _T_75041; // @[Modules.scala 78:156:@28469.4]
  wire [10:0] _T_75042; // @[Modules.scala 78:156:@28470.4]
  wire [10:0] buffer_11_772; // @[Modules.scala 78:156:@28471.4]
  wire [11:0] _T_75044; // @[Modules.scala 78:156:@28473.4]
  wire [10:0] _T_75045; // @[Modules.scala 78:156:@28474.4]
  wire [10:0] buffer_11_773; // @[Modules.scala 78:156:@28475.4]
  wire [11:0] _T_75047; // @[Modules.scala 78:156:@28477.4]
  wire [10:0] _T_75048; // @[Modules.scala 78:156:@28478.4]
  wire [10:0] buffer_11_774; // @[Modules.scala 78:156:@28479.4]
  wire [11:0] _T_75050; // @[Modules.scala 78:156:@28481.4]
  wire [10:0] _T_75051; // @[Modules.scala 78:156:@28482.4]
  wire [10:0] buffer_11_775; // @[Modules.scala 78:156:@28483.4]
  wire [11:0] _T_75053; // @[Modules.scala 78:156:@28485.4]
  wire [10:0] _T_75054; // @[Modules.scala 78:156:@28486.4]
  wire [10:0] buffer_11_776; // @[Modules.scala 78:156:@28487.4]
  wire [11:0] _T_75056; // @[Modules.scala 78:156:@28489.4]
  wire [10:0] _T_75057; // @[Modules.scala 78:156:@28490.4]
  wire [10:0] buffer_11_777; // @[Modules.scala 78:156:@28491.4]
  wire [11:0] _T_75059; // @[Modules.scala 78:156:@28493.4]
  wire [10:0] _T_75060; // @[Modules.scala 78:156:@28494.4]
  wire [10:0] buffer_11_778; // @[Modules.scala 78:156:@28495.4]
  wire [11:0] _T_75062; // @[Modules.scala 78:156:@28497.4]
  wire [10:0] _T_75063; // @[Modules.scala 78:156:@28498.4]
  wire [10:0] buffer_11_779; // @[Modules.scala 78:156:@28499.4]
  wire [11:0] _T_75065; // @[Modules.scala 78:156:@28501.4]
  wire [10:0] _T_75066; // @[Modules.scala 78:156:@28502.4]
  wire [10:0] buffer_11_780; // @[Modules.scala 78:156:@28503.4]
  wire [11:0] _T_75068; // @[Modules.scala 78:156:@28505.4]
  wire [10:0] _T_75069; // @[Modules.scala 78:156:@28506.4]
  wire [10:0] buffer_11_781; // @[Modules.scala 78:156:@28507.4]
  wire [11:0] _T_75071; // @[Modules.scala 78:156:@28509.4]
  wire [10:0] _T_75072; // @[Modules.scala 78:156:@28510.4]
  wire [10:0] buffer_11_782; // @[Modules.scala 78:156:@28511.4]
  wire [11:0] _T_75074; // @[Modules.scala 78:156:@28513.4]
  wire [10:0] _T_75075; // @[Modules.scala 78:156:@28514.4]
  wire [10:0] buffer_11_783; // @[Modules.scala 78:156:@28515.4]
  wire [5:0] _T_75490; // @[Modules.scala 37:46:@29119.4]
  wire [4:0] _T_75491; // @[Modules.scala 37:46:@29120.4]
  wire [4:0] _T_75492; // @[Modules.scala 37:46:@29121.4]
  wire [11:0] _T_75665; // @[Modules.scala 65:57:@29366.4]
  wire [10:0] _T_75666; // @[Modules.scala 65:57:@29367.4]
  wire [10:0] buffer_12_392; // @[Modules.scala 65:57:@29368.4]
  wire [10:0] buffer_12_7; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75674; // @[Modules.scala 65:57:@29378.4]
  wire [10:0] _T_75675; // @[Modules.scala 65:57:@29379.4]
  wire [10:0] buffer_12_395; // @[Modules.scala 65:57:@29380.4]
  wire [11:0] _T_75677; // @[Modules.scala 65:57:@29382.4]
  wire [10:0] _T_75678; // @[Modules.scala 65:57:@29383.4]
  wire [10:0] buffer_12_396; // @[Modules.scala 65:57:@29384.4]
  wire [11:0] _T_75680; // @[Modules.scala 65:57:@29386.4]
  wire [10:0] _T_75681; // @[Modules.scala 65:57:@29387.4]
  wire [10:0] buffer_12_397; // @[Modules.scala 65:57:@29388.4]
  wire [11:0] _T_75683; // @[Modules.scala 65:57:@29390.4]
  wire [10:0] _T_75684; // @[Modules.scala 65:57:@29391.4]
  wire [10:0] buffer_12_398; // @[Modules.scala 65:57:@29392.4]
  wire [11:0] _T_75686; // @[Modules.scala 65:57:@29394.4]
  wire [10:0] _T_75687; // @[Modules.scala 65:57:@29395.4]
  wire [10:0] buffer_12_399; // @[Modules.scala 65:57:@29396.4]
  wire [11:0] _T_75746; // @[Modules.scala 65:57:@29474.4]
  wire [10:0] _T_75747; // @[Modules.scala 65:57:@29475.4]
  wire [10:0] buffer_12_419; // @[Modules.scala 65:57:@29476.4]
  wire [11:0] _T_75752; // @[Modules.scala 65:57:@29482.4]
  wire [10:0] _T_75753; // @[Modules.scala 65:57:@29483.4]
  wire [10:0] buffer_12_421; // @[Modules.scala 65:57:@29484.4]
  wire [11:0] _T_75758; // @[Modules.scala 65:57:@29490.4]
  wire [10:0] _T_75759; // @[Modules.scala 65:57:@29491.4]
  wire [10:0] buffer_12_423; // @[Modules.scala 65:57:@29492.4]
  wire [11:0] _T_75764; // @[Modules.scala 65:57:@29498.4]
  wire [10:0] _T_75765; // @[Modules.scala 65:57:@29499.4]
  wire [10:0] buffer_12_425; // @[Modules.scala 65:57:@29500.4]
  wire [11:0] _T_75767; // @[Modules.scala 65:57:@29502.4]
  wire [10:0] _T_75768; // @[Modules.scala 65:57:@29503.4]
  wire [10:0] buffer_12_426; // @[Modules.scala 65:57:@29504.4]
  wire [11:0] _T_75773; // @[Modules.scala 65:57:@29510.4]
  wire [10:0] _T_75774; // @[Modules.scala 65:57:@29511.4]
  wire [10:0] buffer_12_428; // @[Modules.scala 65:57:@29512.4]
  wire [11:0] _T_75776; // @[Modules.scala 65:57:@29514.4]
  wire [10:0] _T_75777; // @[Modules.scala 65:57:@29515.4]
  wire [10:0] buffer_12_429; // @[Modules.scala 65:57:@29516.4]
  wire [11:0] _T_75782; // @[Modules.scala 65:57:@29522.4]
  wire [10:0] _T_75783; // @[Modules.scala 65:57:@29523.4]
  wire [10:0] buffer_12_431; // @[Modules.scala 65:57:@29524.4]
  wire [11:0] _T_75788; // @[Modules.scala 65:57:@29530.4]
  wire [10:0] _T_75789; // @[Modules.scala 65:57:@29531.4]
  wire [10:0] buffer_12_433; // @[Modules.scala 65:57:@29532.4]
  wire [11:0] _T_75803; // @[Modules.scala 65:57:@29550.4]
  wire [10:0] _T_75804; // @[Modules.scala 65:57:@29551.4]
  wire [10:0] buffer_12_438; // @[Modules.scala 65:57:@29552.4]
  wire [11:0] _T_75815; // @[Modules.scala 65:57:@29566.4]
  wire [10:0] _T_75816; // @[Modules.scala 65:57:@29567.4]
  wire [10:0] buffer_12_442; // @[Modules.scala 65:57:@29568.4]
  wire [11:0] _T_75818; // @[Modules.scala 65:57:@29570.4]
  wire [10:0] _T_75819; // @[Modules.scala 65:57:@29571.4]
  wire [10:0] buffer_12_443; // @[Modules.scala 65:57:@29572.4]
  wire [11:0] _T_75824; // @[Modules.scala 65:57:@29578.4]
  wire [10:0] _T_75825; // @[Modules.scala 65:57:@29579.4]
  wire [10:0] buffer_12_445; // @[Modules.scala 65:57:@29580.4]
  wire [10:0] buffer_12_113; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75833; // @[Modules.scala 65:57:@29590.4]
  wire [10:0] _T_75834; // @[Modules.scala 65:57:@29591.4]
  wire [10:0] buffer_12_448; // @[Modules.scala 65:57:@29592.4]
  wire [11:0] _T_75839; // @[Modules.scala 65:57:@29598.4]
  wire [10:0] _T_75840; // @[Modules.scala 65:57:@29599.4]
  wire [10:0] buffer_12_450; // @[Modules.scala 65:57:@29600.4]
  wire [11:0] _T_75842; // @[Modules.scala 65:57:@29602.4]
  wire [10:0] _T_75843; // @[Modules.scala 65:57:@29603.4]
  wire [10:0] buffer_12_451; // @[Modules.scala 65:57:@29604.4]
  wire [11:0] _T_75854; // @[Modules.scala 65:57:@29618.4]
  wire [10:0] _T_75855; // @[Modules.scala 65:57:@29619.4]
  wire [10:0] buffer_12_455; // @[Modules.scala 65:57:@29620.4]
  wire [11:0] _T_75857; // @[Modules.scala 65:57:@29622.4]
  wire [10:0] _T_75858; // @[Modules.scala 65:57:@29623.4]
  wire [10:0] buffer_12_456; // @[Modules.scala 65:57:@29624.4]
  wire [11:0] _T_75860; // @[Modules.scala 65:57:@29626.4]
  wire [10:0] _T_75861; // @[Modules.scala 65:57:@29627.4]
  wire [10:0] buffer_12_457; // @[Modules.scala 65:57:@29628.4]
  wire [11:0] _T_75863; // @[Modules.scala 65:57:@29630.4]
  wire [10:0] _T_75864; // @[Modules.scala 65:57:@29631.4]
  wire [10:0] buffer_12_458; // @[Modules.scala 65:57:@29632.4]
  wire [11:0] _T_75866; // @[Modules.scala 65:57:@29634.4]
  wire [10:0] _T_75867; // @[Modules.scala 65:57:@29635.4]
  wire [10:0] buffer_12_459; // @[Modules.scala 65:57:@29636.4]
  wire [11:0] _T_75875; // @[Modules.scala 65:57:@29646.4]
  wire [10:0] _T_75876; // @[Modules.scala 65:57:@29647.4]
  wire [10:0] buffer_12_462; // @[Modules.scala 65:57:@29648.4]
  wire [11:0] _T_75887; // @[Modules.scala 65:57:@29662.4]
  wire [10:0] _T_75888; // @[Modules.scala 65:57:@29663.4]
  wire [10:0] buffer_12_466; // @[Modules.scala 65:57:@29664.4]
  wire [11:0] _T_75890; // @[Modules.scala 65:57:@29666.4]
  wire [10:0] _T_75891; // @[Modules.scala 65:57:@29667.4]
  wire [10:0] buffer_12_467; // @[Modules.scala 65:57:@29668.4]
  wire [10:0] buffer_12_155; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75896; // @[Modules.scala 65:57:@29674.4]
  wire [10:0] _T_75897; // @[Modules.scala 65:57:@29675.4]
  wire [10:0] buffer_12_469; // @[Modules.scala 65:57:@29676.4]
  wire [10:0] buffer_12_163; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75908; // @[Modules.scala 65:57:@29690.4]
  wire [10:0] _T_75909; // @[Modules.scala 65:57:@29691.4]
  wire [10:0] buffer_12_473; // @[Modules.scala 65:57:@29692.4]
  wire [10:0] buffer_12_164; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75911; // @[Modules.scala 65:57:@29694.4]
  wire [10:0] _T_75912; // @[Modules.scala 65:57:@29695.4]
  wire [10:0] buffer_12_474; // @[Modules.scala 65:57:@29696.4]
  wire [10:0] buffer_12_166; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75914; // @[Modules.scala 65:57:@29698.4]
  wire [10:0] _T_75915; // @[Modules.scala 65:57:@29699.4]
  wire [10:0] buffer_12_475; // @[Modules.scala 65:57:@29700.4]
  wire [11:0] _T_75917; // @[Modules.scala 65:57:@29702.4]
  wire [10:0] _T_75918; // @[Modules.scala 65:57:@29703.4]
  wire [10:0] buffer_12_476; // @[Modules.scala 65:57:@29704.4]
  wire [11:0] _T_75959; // @[Modules.scala 65:57:@29758.4]
  wire [10:0] _T_75960; // @[Modules.scala 65:57:@29759.4]
  wire [10:0] buffer_12_490; // @[Modules.scala 65:57:@29760.4]
  wire [11:0] _T_75962; // @[Modules.scala 65:57:@29762.4]
  wire [10:0] _T_75963; // @[Modules.scala 65:57:@29763.4]
  wire [10:0] buffer_12_491; // @[Modules.scala 65:57:@29764.4]
  wire [10:0] buffer_12_206; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_75974; // @[Modules.scala 65:57:@29778.4]
  wire [10:0] _T_75975; // @[Modules.scala 65:57:@29779.4]
  wire [10:0] buffer_12_495; // @[Modules.scala 65:57:@29780.4]
  wire [11:0] _T_75980; // @[Modules.scala 65:57:@29786.4]
  wire [10:0] _T_75981; // @[Modules.scala 65:57:@29787.4]
  wire [10:0] buffer_12_497; // @[Modules.scala 65:57:@29788.4]
  wire [11:0] _T_75995; // @[Modules.scala 65:57:@29806.4]
  wire [10:0] _T_75996; // @[Modules.scala 65:57:@29807.4]
  wire [10:0] buffer_12_502; // @[Modules.scala 65:57:@29808.4]
  wire [11:0] _T_76010; // @[Modules.scala 65:57:@29826.4]
  wire [10:0] _T_76011; // @[Modules.scala 65:57:@29827.4]
  wire [10:0] buffer_12_507; // @[Modules.scala 65:57:@29828.4]
  wire [11:0] _T_76016; // @[Modules.scala 65:57:@29834.4]
  wire [10:0] _T_76017; // @[Modules.scala 65:57:@29835.4]
  wire [10:0] buffer_12_509; // @[Modules.scala 65:57:@29836.4]
  wire [10:0] buffer_12_238; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76022; // @[Modules.scala 65:57:@29842.4]
  wire [10:0] _T_76023; // @[Modules.scala 65:57:@29843.4]
  wire [10:0] buffer_12_511; // @[Modules.scala 65:57:@29844.4]
  wire [10:0] buffer_12_244; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_12_245; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76031; // @[Modules.scala 65:57:@29854.4]
  wire [10:0] _T_76032; // @[Modules.scala 65:57:@29855.4]
  wire [10:0] buffer_12_514; // @[Modules.scala 65:57:@29856.4]
  wire [11:0] _T_76043; // @[Modules.scala 65:57:@29870.4]
  wire [10:0] _T_76044; // @[Modules.scala 65:57:@29871.4]
  wire [10:0] buffer_12_518; // @[Modules.scala 65:57:@29872.4]
  wire [11:0] _T_76046; // @[Modules.scala 65:57:@29874.4]
  wire [10:0] _T_76047; // @[Modules.scala 65:57:@29875.4]
  wire [10:0] buffer_12_519; // @[Modules.scala 65:57:@29876.4]
  wire [11:0] _T_76052; // @[Modules.scala 65:57:@29882.4]
  wire [10:0] _T_76053; // @[Modules.scala 65:57:@29883.4]
  wire [10:0] buffer_12_521; // @[Modules.scala 65:57:@29884.4]
  wire [11:0] _T_76058; // @[Modules.scala 65:57:@29890.4]
  wire [10:0] _T_76059; // @[Modules.scala 65:57:@29891.4]
  wire [10:0] buffer_12_523; // @[Modules.scala 65:57:@29892.4]
  wire [11:0] _T_76064; // @[Modules.scala 65:57:@29898.4]
  wire [10:0] _T_76065; // @[Modules.scala 65:57:@29899.4]
  wire [10:0] buffer_12_525; // @[Modules.scala 65:57:@29900.4]
  wire [11:0] _T_76076; // @[Modules.scala 65:57:@29914.4]
  wire [10:0] _T_76077; // @[Modules.scala 65:57:@29915.4]
  wire [10:0] buffer_12_529; // @[Modules.scala 65:57:@29916.4]
  wire [10:0] buffer_12_280; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76085; // @[Modules.scala 65:57:@29926.4]
  wire [10:0] _T_76086; // @[Modules.scala 65:57:@29927.4]
  wire [10:0] buffer_12_532; // @[Modules.scala 65:57:@29928.4]
  wire [10:0] buffer_12_288; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76097; // @[Modules.scala 65:57:@29942.4]
  wire [10:0] _T_76098; // @[Modules.scala 65:57:@29943.4]
  wire [10:0] buffer_12_536; // @[Modules.scala 65:57:@29944.4]
  wire [11:0] _T_76106; // @[Modules.scala 65:57:@29954.4]
  wire [10:0] _T_76107; // @[Modules.scala 65:57:@29955.4]
  wire [10:0] buffer_12_539; // @[Modules.scala 65:57:@29956.4]
  wire [10:0] buffer_12_296; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76109; // @[Modules.scala 65:57:@29958.4]
  wire [10:0] _T_76110; // @[Modules.scala 65:57:@29959.4]
  wire [10:0] buffer_12_540; // @[Modules.scala 65:57:@29960.4]
  wire [11:0] _T_76112; // @[Modules.scala 65:57:@29962.4]
  wire [10:0] _T_76113; // @[Modules.scala 65:57:@29963.4]
  wire [10:0] buffer_12_541; // @[Modules.scala 65:57:@29964.4]
  wire [10:0] buffer_12_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76127; // @[Modules.scala 65:57:@29982.4]
  wire [10:0] _T_76128; // @[Modules.scala 65:57:@29983.4]
  wire [10:0] buffer_12_546; // @[Modules.scala 65:57:@29984.4]
  wire [11:0] _T_76148; // @[Modules.scala 65:57:@30010.4]
  wire [10:0] _T_76149; // @[Modules.scala 65:57:@30011.4]
  wire [10:0] buffer_12_553; // @[Modules.scala 65:57:@30012.4]
  wire [11:0] _T_76166; // @[Modules.scala 65:57:@30034.4]
  wire [10:0] _T_76167; // @[Modules.scala 65:57:@30035.4]
  wire [10:0] buffer_12_559; // @[Modules.scala 65:57:@30036.4]
  wire [11:0] _T_76175; // @[Modules.scala 65:57:@30046.4]
  wire [10:0] _T_76176; // @[Modules.scala 65:57:@30047.4]
  wire [10:0] buffer_12_562; // @[Modules.scala 65:57:@30048.4]
  wire [11:0] _T_76178; // @[Modules.scala 65:57:@30050.4]
  wire [10:0] _T_76179; // @[Modules.scala 65:57:@30051.4]
  wire [10:0] buffer_12_563; // @[Modules.scala 65:57:@30052.4]
  wire [11:0] _T_76187; // @[Modules.scala 65:57:@30062.4]
  wire [10:0] _T_76188; // @[Modules.scala 65:57:@30063.4]
  wire [10:0] buffer_12_566; // @[Modules.scala 65:57:@30064.4]
  wire [11:0] _T_76190; // @[Modules.scala 65:57:@30066.4]
  wire [10:0] _T_76191; // @[Modules.scala 65:57:@30067.4]
  wire [10:0] buffer_12_567; // @[Modules.scala 65:57:@30068.4]
  wire [11:0] _T_76211; // @[Modules.scala 65:57:@30094.4]
  wire [10:0] _T_76212; // @[Modules.scala 65:57:@30095.4]
  wire [10:0] buffer_12_574; // @[Modules.scala 65:57:@30096.4]
  wire [11:0] _T_76229; // @[Modules.scala 65:57:@30118.4]
  wire [10:0] _T_76230; // @[Modules.scala 65:57:@30119.4]
  wire [10:0] buffer_12_580; // @[Modules.scala 65:57:@30120.4]
  wire [11:0] _T_76232; // @[Modules.scala 65:57:@30122.4]
  wire [10:0] _T_76233; // @[Modules.scala 65:57:@30123.4]
  wire [10:0] buffer_12_581; // @[Modules.scala 65:57:@30124.4]
  wire [11:0] _T_76238; // @[Modules.scala 65:57:@30130.4]
  wire [10:0] _T_76239; // @[Modules.scala 65:57:@30131.4]
  wire [10:0] buffer_12_583; // @[Modules.scala 65:57:@30132.4]
  wire [10:0] buffer_12_388; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_76247; // @[Modules.scala 65:57:@30142.4]
  wire [10:0] _T_76248; // @[Modules.scala 65:57:@30143.4]
  wire [10:0] buffer_12_586; // @[Modules.scala 65:57:@30144.4]
  wire [11:0] _T_76253; // @[Modules.scala 68:83:@30150.4]
  wire [10:0] _T_76254; // @[Modules.scala 68:83:@30151.4]
  wire [10:0] buffer_12_588; // @[Modules.scala 68:83:@30152.4]
  wire [11:0] _T_76256; // @[Modules.scala 68:83:@30154.4]
  wire [10:0] _T_76257; // @[Modules.scala 68:83:@30155.4]
  wire [10:0] buffer_12_589; // @[Modules.scala 68:83:@30156.4]
  wire [11:0] _T_76259; // @[Modules.scala 68:83:@30158.4]
  wire [10:0] _T_76260; // @[Modules.scala 68:83:@30159.4]
  wire [10:0] buffer_12_590; // @[Modules.scala 68:83:@30160.4]
  wire [11:0] _T_76262; // @[Modules.scala 68:83:@30162.4]
  wire [10:0] _T_76263; // @[Modules.scala 68:83:@30163.4]
  wire [10:0] buffer_12_591; // @[Modules.scala 68:83:@30164.4]
  wire [11:0] _T_76274; // @[Modules.scala 68:83:@30178.4]
  wire [10:0] _T_76275; // @[Modules.scala 68:83:@30179.4]
  wire [10:0] buffer_12_595; // @[Modules.scala 68:83:@30180.4]
  wire [11:0] _T_76283; // @[Modules.scala 68:83:@30190.4]
  wire [10:0] _T_76284; // @[Modules.scala 68:83:@30191.4]
  wire [10:0] buffer_12_598; // @[Modules.scala 68:83:@30192.4]
  wire [11:0] _T_76292; // @[Modules.scala 68:83:@30202.4]
  wire [10:0] _T_76293; // @[Modules.scala 68:83:@30203.4]
  wire [10:0] buffer_12_601; // @[Modules.scala 68:83:@30204.4]
  wire [11:0] _T_76295; // @[Modules.scala 68:83:@30206.4]
  wire [10:0] _T_76296; // @[Modules.scala 68:83:@30207.4]
  wire [10:0] buffer_12_602; // @[Modules.scala 68:83:@30208.4]
  wire [11:0] _T_76298; // @[Modules.scala 68:83:@30210.4]
  wire [10:0] _T_76299; // @[Modules.scala 68:83:@30211.4]
  wire [10:0] buffer_12_603; // @[Modules.scala 68:83:@30212.4]
  wire [11:0] _T_76301; // @[Modules.scala 68:83:@30214.4]
  wire [10:0] _T_76302; // @[Modules.scala 68:83:@30215.4]
  wire [10:0] buffer_12_604; // @[Modules.scala 68:83:@30216.4]
  wire [11:0] _T_76304; // @[Modules.scala 68:83:@30218.4]
  wire [10:0] _T_76305; // @[Modules.scala 68:83:@30219.4]
  wire [10:0] buffer_12_605; // @[Modules.scala 68:83:@30220.4]
  wire [11:0] _T_76307; // @[Modules.scala 68:83:@30222.4]
  wire [10:0] _T_76308; // @[Modules.scala 68:83:@30223.4]
  wire [10:0] buffer_12_606; // @[Modules.scala 68:83:@30224.4]
  wire [11:0] _T_76310; // @[Modules.scala 68:83:@30226.4]
  wire [10:0] _T_76311; // @[Modules.scala 68:83:@30227.4]
  wire [10:0] buffer_12_607; // @[Modules.scala 68:83:@30228.4]
  wire [11:0] _T_76313; // @[Modules.scala 68:83:@30230.4]
  wire [10:0] _T_76314; // @[Modules.scala 68:83:@30231.4]
  wire [10:0] buffer_12_608; // @[Modules.scala 68:83:@30232.4]
  wire [11:0] _T_76319; // @[Modules.scala 68:83:@30238.4]
  wire [10:0] _T_76320; // @[Modules.scala 68:83:@30239.4]
  wire [10:0] buffer_12_610; // @[Modules.scala 68:83:@30240.4]
  wire [11:0] _T_76322; // @[Modules.scala 68:83:@30242.4]
  wire [10:0] _T_76323; // @[Modules.scala 68:83:@30243.4]
  wire [10:0] buffer_12_611; // @[Modules.scala 68:83:@30244.4]
  wire [11:0] _T_76328; // @[Modules.scala 68:83:@30250.4]
  wire [10:0] _T_76329; // @[Modules.scala 68:83:@30251.4]
  wire [10:0] buffer_12_613; // @[Modules.scala 68:83:@30252.4]
  wire [11:0] _T_76331; // @[Modules.scala 68:83:@30254.4]
  wire [10:0] _T_76332; // @[Modules.scala 68:83:@30255.4]
  wire [10:0] buffer_12_614; // @[Modules.scala 68:83:@30256.4]
  wire [11:0] _T_76337; // @[Modules.scala 68:83:@30262.4]
  wire [10:0] _T_76338; // @[Modules.scala 68:83:@30263.4]
  wire [10:0] buffer_12_616; // @[Modules.scala 68:83:@30264.4]
  wire [11:0] _T_76340; // @[Modules.scala 68:83:@30266.4]
  wire [10:0] _T_76341; // @[Modules.scala 68:83:@30267.4]
  wire [10:0] buffer_12_617; // @[Modules.scala 68:83:@30268.4]
  wire [11:0] _T_76343; // @[Modules.scala 68:83:@30270.4]
  wire [10:0] _T_76344; // @[Modules.scala 68:83:@30271.4]
  wire [10:0] buffer_12_618; // @[Modules.scala 68:83:@30272.4]
  wire [11:0] _T_76346; // @[Modules.scala 68:83:@30274.4]
  wire [10:0] _T_76347; // @[Modules.scala 68:83:@30275.4]
  wire [10:0] buffer_12_619; // @[Modules.scala 68:83:@30276.4]
  wire [11:0] _T_76349; // @[Modules.scala 68:83:@30278.4]
  wire [10:0] _T_76350; // @[Modules.scala 68:83:@30279.4]
  wire [10:0] buffer_12_620; // @[Modules.scala 68:83:@30280.4]
  wire [11:0] _T_76352; // @[Modules.scala 68:83:@30282.4]
  wire [10:0] _T_76353; // @[Modules.scala 68:83:@30283.4]
  wire [10:0] buffer_12_621; // @[Modules.scala 68:83:@30284.4]
  wire [11:0] _T_76358; // @[Modules.scala 68:83:@30290.4]
  wire [10:0] _T_76359; // @[Modules.scala 68:83:@30291.4]
  wire [10:0] buffer_12_623; // @[Modules.scala 68:83:@30292.4]
  wire [11:0] _T_76361; // @[Modules.scala 68:83:@30294.4]
  wire [10:0] _T_76362; // @[Modules.scala 68:83:@30295.4]
  wire [10:0] buffer_12_624; // @[Modules.scala 68:83:@30296.4]
  wire [11:0] _T_76364; // @[Modules.scala 68:83:@30298.4]
  wire [10:0] _T_76365; // @[Modules.scala 68:83:@30299.4]
  wire [10:0] buffer_12_625; // @[Modules.scala 68:83:@30300.4]
  wire [11:0] _T_76367; // @[Modules.scala 68:83:@30302.4]
  wire [10:0] _T_76368; // @[Modules.scala 68:83:@30303.4]
  wire [10:0] buffer_12_626; // @[Modules.scala 68:83:@30304.4]
  wire [11:0] _T_76373; // @[Modules.scala 68:83:@30310.4]
  wire [10:0] _T_76374; // @[Modules.scala 68:83:@30311.4]
  wire [10:0] buffer_12_628; // @[Modules.scala 68:83:@30312.4]
  wire [11:0] _T_76376; // @[Modules.scala 68:83:@30314.4]
  wire [10:0] _T_76377; // @[Modules.scala 68:83:@30315.4]
  wire [10:0] buffer_12_629; // @[Modules.scala 68:83:@30316.4]
  wire [11:0] _T_76379; // @[Modules.scala 68:83:@30318.4]
  wire [10:0] _T_76380; // @[Modules.scala 68:83:@30319.4]
  wire [10:0] buffer_12_630; // @[Modules.scala 68:83:@30320.4]
  wire [11:0] _T_76385; // @[Modules.scala 68:83:@30326.4]
  wire [10:0] _T_76386; // @[Modules.scala 68:83:@30327.4]
  wire [10:0] buffer_12_632; // @[Modules.scala 68:83:@30328.4]
  wire [11:0] _T_76388; // @[Modules.scala 68:83:@30330.4]
  wire [10:0] _T_76389; // @[Modules.scala 68:83:@30331.4]
  wire [10:0] buffer_12_633; // @[Modules.scala 68:83:@30332.4]
  wire [11:0] _T_76397; // @[Modules.scala 68:83:@30342.4]
  wire [10:0] _T_76398; // @[Modules.scala 68:83:@30343.4]
  wire [10:0] buffer_12_636; // @[Modules.scala 68:83:@30344.4]
  wire [11:0] _T_76400; // @[Modules.scala 68:83:@30346.4]
  wire [10:0] _T_76401; // @[Modules.scala 68:83:@30347.4]
  wire [10:0] buffer_12_637; // @[Modules.scala 68:83:@30348.4]
  wire [11:0] _T_76403; // @[Modules.scala 68:83:@30350.4]
  wire [10:0] _T_76404; // @[Modules.scala 68:83:@30351.4]
  wire [10:0] buffer_12_638; // @[Modules.scala 68:83:@30352.4]
  wire [11:0] _T_76406; // @[Modules.scala 68:83:@30354.4]
  wire [10:0] _T_76407; // @[Modules.scala 68:83:@30355.4]
  wire [10:0] buffer_12_639; // @[Modules.scala 68:83:@30356.4]
  wire [11:0] _T_76409; // @[Modules.scala 68:83:@30358.4]
  wire [10:0] _T_76410; // @[Modules.scala 68:83:@30359.4]
  wire [10:0] buffer_12_640; // @[Modules.scala 68:83:@30360.4]
  wire [11:0] _T_76418; // @[Modules.scala 68:83:@30370.4]
  wire [10:0] _T_76419; // @[Modules.scala 68:83:@30371.4]
  wire [10:0] buffer_12_643; // @[Modules.scala 68:83:@30372.4]
  wire [11:0] _T_76424; // @[Modules.scala 68:83:@30378.4]
  wire [10:0] _T_76425; // @[Modules.scala 68:83:@30379.4]
  wire [10:0] buffer_12_645; // @[Modules.scala 68:83:@30380.4]
  wire [11:0] _T_76427; // @[Modules.scala 68:83:@30382.4]
  wire [10:0] _T_76428; // @[Modules.scala 68:83:@30383.4]
  wire [10:0] buffer_12_646; // @[Modules.scala 68:83:@30384.4]
  wire [11:0] _T_76430; // @[Modules.scala 68:83:@30386.4]
  wire [10:0] _T_76431; // @[Modules.scala 68:83:@30387.4]
  wire [10:0] buffer_12_647; // @[Modules.scala 68:83:@30388.4]
  wire [11:0] _T_76433; // @[Modules.scala 68:83:@30390.4]
  wire [10:0] _T_76434; // @[Modules.scala 68:83:@30391.4]
  wire [10:0] buffer_12_648; // @[Modules.scala 68:83:@30392.4]
  wire [11:0] _T_76436; // @[Modules.scala 68:83:@30394.4]
  wire [10:0] _T_76437; // @[Modules.scala 68:83:@30395.4]
  wire [10:0] buffer_12_649; // @[Modules.scala 68:83:@30396.4]
  wire [11:0] _T_76442; // @[Modules.scala 68:83:@30402.4]
  wire [10:0] _T_76443; // @[Modules.scala 68:83:@30403.4]
  wire [10:0] buffer_12_651; // @[Modules.scala 68:83:@30404.4]
  wire [11:0] _T_76445; // @[Modules.scala 68:83:@30406.4]
  wire [10:0] _T_76446; // @[Modules.scala 68:83:@30407.4]
  wire [10:0] buffer_12_652; // @[Modules.scala 68:83:@30408.4]
  wire [11:0] _T_76448; // @[Modules.scala 68:83:@30410.4]
  wire [10:0] _T_76449; // @[Modules.scala 68:83:@30411.4]
  wire [10:0] buffer_12_653; // @[Modules.scala 68:83:@30412.4]
  wire [11:0] _T_76451; // @[Modules.scala 68:83:@30414.4]
  wire [10:0] _T_76452; // @[Modules.scala 68:83:@30415.4]
  wire [10:0] buffer_12_654; // @[Modules.scala 68:83:@30416.4]
  wire [11:0] _T_76457; // @[Modules.scala 68:83:@30422.4]
  wire [10:0] _T_76458; // @[Modules.scala 68:83:@30423.4]
  wire [10:0] buffer_12_656; // @[Modules.scala 68:83:@30424.4]
  wire [11:0] _T_76463; // @[Modules.scala 68:83:@30430.4]
  wire [10:0] _T_76464; // @[Modules.scala 68:83:@30431.4]
  wire [10:0] buffer_12_658; // @[Modules.scala 68:83:@30432.4]
  wire [11:0] _T_76469; // @[Modules.scala 68:83:@30438.4]
  wire [10:0] _T_76470; // @[Modules.scala 68:83:@30439.4]
  wire [10:0] buffer_12_660; // @[Modules.scala 68:83:@30440.4]
  wire [11:0] _T_76472; // @[Modules.scala 68:83:@30442.4]
  wire [10:0] _T_76473; // @[Modules.scala 68:83:@30443.4]
  wire [10:0] buffer_12_661; // @[Modules.scala 68:83:@30444.4]
  wire [11:0] _T_76475; // @[Modules.scala 68:83:@30446.4]
  wire [10:0] _T_76476; // @[Modules.scala 68:83:@30447.4]
  wire [10:0] buffer_12_662; // @[Modules.scala 68:83:@30448.4]
  wire [11:0] _T_76481; // @[Modules.scala 68:83:@30454.4]
  wire [10:0] _T_76482; // @[Modules.scala 68:83:@30455.4]
  wire [10:0] buffer_12_664; // @[Modules.scala 68:83:@30456.4]
  wire [11:0] _T_76484; // @[Modules.scala 68:83:@30458.4]
  wire [10:0] _T_76485; // @[Modules.scala 68:83:@30459.4]
  wire [10:0] buffer_12_665; // @[Modules.scala 68:83:@30460.4]
  wire [11:0] _T_76487; // @[Modules.scala 68:83:@30462.4]
  wire [10:0] _T_76488; // @[Modules.scala 68:83:@30463.4]
  wire [10:0] buffer_12_666; // @[Modules.scala 68:83:@30464.4]
  wire [11:0] _T_76490; // @[Modules.scala 68:83:@30466.4]
  wire [10:0] _T_76491; // @[Modules.scala 68:83:@30467.4]
  wire [10:0] buffer_12_667; // @[Modules.scala 68:83:@30468.4]
  wire [11:0] _T_76493; // @[Modules.scala 68:83:@30470.4]
  wire [10:0] _T_76494; // @[Modules.scala 68:83:@30471.4]
  wire [10:0] buffer_12_668; // @[Modules.scala 68:83:@30472.4]
  wire [11:0] _T_76496; // @[Modules.scala 68:83:@30474.4]
  wire [10:0] _T_76497; // @[Modules.scala 68:83:@30475.4]
  wire [10:0] buffer_12_669; // @[Modules.scala 68:83:@30476.4]
  wire [11:0] _T_76502; // @[Modules.scala 68:83:@30482.4]
  wire [10:0] _T_76503; // @[Modules.scala 68:83:@30483.4]
  wire [10:0] buffer_12_671; // @[Modules.scala 68:83:@30484.4]
  wire [11:0] _T_76508; // @[Modules.scala 68:83:@30490.4]
  wire [10:0] _T_76509; // @[Modules.scala 68:83:@30491.4]
  wire [10:0] buffer_12_673; // @[Modules.scala 68:83:@30492.4]
  wire [11:0] _T_76514; // @[Modules.scala 68:83:@30498.4]
  wire [10:0] _T_76515; // @[Modules.scala 68:83:@30499.4]
  wire [10:0] buffer_12_675; // @[Modules.scala 68:83:@30500.4]
  wire [11:0] _T_76526; // @[Modules.scala 68:83:@30514.4]
  wire [10:0] _T_76527; // @[Modules.scala 68:83:@30515.4]
  wire [10:0] buffer_12_679; // @[Modules.scala 68:83:@30516.4]
  wire [11:0] _T_76535; // @[Modules.scala 68:83:@30526.4]
  wire [10:0] _T_76536; // @[Modules.scala 68:83:@30527.4]
  wire [10:0] buffer_12_682; // @[Modules.scala 68:83:@30528.4]
  wire [11:0] _T_76538; // @[Modules.scala 68:83:@30530.4]
  wire [10:0] _T_76539; // @[Modules.scala 68:83:@30531.4]
  wire [10:0] buffer_12_683; // @[Modules.scala 68:83:@30532.4]
  wire [11:0] _T_76544; // @[Modules.scala 68:83:@30538.4]
  wire [10:0] _T_76545; // @[Modules.scala 68:83:@30539.4]
  wire [10:0] buffer_12_685; // @[Modules.scala 68:83:@30540.4]
  wire [11:0] _T_76547; // @[Modules.scala 71:109:@30542.4]
  wire [10:0] _T_76548; // @[Modules.scala 71:109:@30543.4]
  wire [10:0] buffer_12_686; // @[Modules.scala 71:109:@30544.4]
  wire [11:0] _T_76550; // @[Modules.scala 71:109:@30546.4]
  wire [10:0] _T_76551; // @[Modules.scala 71:109:@30547.4]
  wire [10:0] buffer_12_687; // @[Modules.scala 71:109:@30548.4]
  wire [11:0] _T_76553; // @[Modules.scala 71:109:@30550.4]
  wire [10:0] _T_76554; // @[Modules.scala 71:109:@30551.4]
  wire [10:0] buffer_12_688; // @[Modules.scala 71:109:@30552.4]
  wire [11:0] _T_76556; // @[Modules.scala 71:109:@30554.4]
  wire [10:0] _T_76557; // @[Modules.scala 71:109:@30555.4]
  wire [10:0] buffer_12_689; // @[Modules.scala 71:109:@30556.4]
  wire [11:0] _T_76562; // @[Modules.scala 71:109:@30562.4]
  wire [10:0] _T_76563; // @[Modules.scala 71:109:@30563.4]
  wire [10:0] buffer_12_691; // @[Modules.scala 71:109:@30564.4]
  wire [11:0] _T_76565; // @[Modules.scala 71:109:@30566.4]
  wire [10:0] _T_76566; // @[Modules.scala 71:109:@30567.4]
  wire [10:0] buffer_12_692; // @[Modules.scala 71:109:@30568.4]
  wire [11:0] _T_76568; // @[Modules.scala 71:109:@30570.4]
  wire [10:0] _T_76569; // @[Modules.scala 71:109:@30571.4]
  wire [10:0] buffer_12_693; // @[Modules.scala 71:109:@30572.4]
  wire [11:0] _T_76571; // @[Modules.scala 71:109:@30574.4]
  wire [10:0] _T_76572; // @[Modules.scala 71:109:@30575.4]
  wire [10:0] buffer_12_694; // @[Modules.scala 71:109:@30576.4]
  wire [11:0] _T_76574; // @[Modules.scala 71:109:@30578.4]
  wire [10:0] _T_76575; // @[Modules.scala 71:109:@30579.4]
  wire [10:0] buffer_12_695; // @[Modules.scala 71:109:@30580.4]
  wire [11:0] _T_76577; // @[Modules.scala 71:109:@30582.4]
  wire [10:0] _T_76578; // @[Modules.scala 71:109:@30583.4]
  wire [10:0] buffer_12_696; // @[Modules.scala 71:109:@30584.4]
  wire [11:0] _T_76580; // @[Modules.scala 71:109:@30586.4]
  wire [10:0] _T_76581; // @[Modules.scala 71:109:@30587.4]
  wire [10:0] buffer_12_697; // @[Modules.scala 71:109:@30588.4]
  wire [11:0] _T_76583; // @[Modules.scala 71:109:@30590.4]
  wire [10:0] _T_76584; // @[Modules.scala 71:109:@30591.4]
  wire [10:0] buffer_12_698; // @[Modules.scala 71:109:@30592.4]
  wire [11:0] _T_76586; // @[Modules.scala 71:109:@30594.4]
  wire [10:0] _T_76587; // @[Modules.scala 71:109:@30595.4]
  wire [10:0] buffer_12_699; // @[Modules.scala 71:109:@30596.4]
  wire [11:0] _T_76589; // @[Modules.scala 71:109:@30598.4]
  wire [10:0] _T_76590; // @[Modules.scala 71:109:@30599.4]
  wire [10:0] buffer_12_700; // @[Modules.scala 71:109:@30600.4]
  wire [11:0] _T_76592; // @[Modules.scala 71:109:@30602.4]
  wire [10:0] _T_76593; // @[Modules.scala 71:109:@30603.4]
  wire [10:0] buffer_12_701; // @[Modules.scala 71:109:@30604.4]
  wire [11:0] _T_76595; // @[Modules.scala 71:109:@30606.4]
  wire [10:0] _T_76596; // @[Modules.scala 71:109:@30607.4]
  wire [10:0] buffer_12_702; // @[Modules.scala 71:109:@30608.4]
  wire [11:0] _T_76598; // @[Modules.scala 71:109:@30610.4]
  wire [10:0] _T_76599; // @[Modules.scala 71:109:@30611.4]
  wire [10:0] buffer_12_703; // @[Modules.scala 71:109:@30612.4]
  wire [11:0] _T_76601; // @[Modules.scala 71:109:@30614.4]
  wire [10:0] _T_76602; // @[Modules.scala 71:109:@30615.4]
  wire [10:0] buffer_12_704; // @[Modules.scala 71:109:@30616.4]
  wire [11:0] _T_76604; // @[Modules.scala 71:109:@30618.4]
  wire [10:0] _T_76605; // @[Modules.scala 71:109:@30619.4]
  wire [10:0] buffer_12_705; // @[Modules.scala 71:109:@30620.4]
  wire [11:0] _T_76607; // @[Modules.scala 71:109:@30622.4]
  wire [10:0] _T_76608; // @[Modules.scala 71:109:@30623.4]
  wire [10:0] buffer_12_706; // @[Modules.scala 71:109:@30624.4]
  wire [11:0] _T_76610; // @[Modules.scala 71:109:@30626.4]
  wire [10:0] _T_76611; // @[Modules.scala 71:109:@30627.4]
  wire [10:0] buffer_12_707; // @[Modules.scala 71:109:@30628.4]
  wire [11:0] _T_76613; // @[Modules.scala 71:109:@30630.4]
  wire [10:0] _T_76614; // @[Modules.scala 71:109:@30631.4]
  wire [10:0] buffer_12_708; // @[Modules.scala 71:109:@30632.4]
  wire [11:0] _T_76619; // @[Modules.scala 71:109:@30638.4]
  wire [10:0] _T_76620; // @[Modules.scala 71:109:@30639.4]
  wire [10:0] buffer_12_710; // @[Modules.scala 71:109:@30640.4]
  wire [11:0] _T_76622; // @[Modules.scala 71:109:@30642.4]
  wire [10:0] _T_76623; // @[Modules.scala 71:109:@30643.4]
  wire [10:0] buffer_12_711; // @[Modules.scala 71:109:@30644.4]
  wire [11:0] _T_76625; // @[Modules.scala 71:109:@30646.4]
  wire [10:0] _T_76626; // @[Modules.scala 71:109:@30647.4]
  wire [10:0] buffer_12_712; // @[Modules.scala 71:109:@30648.4]
  wire [11:0] _T_76628; // @[Modules.scala 71:109:@30650.4]
  wire [10:0] _T_76629; // @[Modules.scala 71:109:@30651.4]
  wire [10:0] buffer_12_713; // @[Modules.scala 71:109:@30652.4]
  wire [11:0] _T_76631; // @[Modules.scala 71:109:@30654.4]
  wire [10:0] _T_76632; // @[Modules.scala 71:109:@30655.4]
  wire [10:0] buffer_12_714; // @[Modules.scala 71:109:@30656.4]
  wire [11:0] _T_76634; // @[Modules.scala 71:109:@30658.4]
  wire [10:0] _T_76635; // @[Modules.scala 71:109:@30659.4]
  wire [10:0] buffer_12_715; // @[Modules.scala 71:109:@30660.4]
  wire [11:0] _T_76637; // @[Modules.scala 71:109:@30662.4]
  wire [10:0] _T_76638; // @[Modules.scala 71:109:@30663.4]
  wire [10:0] buffer_12_716; // @[Modules.scala 71:109:@30664.4]
  wire [11:0] _T_76640; // @[Modules.scala 71:109:@30666.4]
  wire [10:0] _T_76641; // @[Modules.scala 71:109:@30667.4]
  wire [10:0] buffer_12_717; // @[Modules.scala 71:109:@30668.4]
  wire [11:0] _T_76643; // @[Modules.scala 71:109:@30670.4]
  wire [10:0] _T_76644; // @[Modules.scala 71:109:@30671.4]
  wire [10:0] buffer_12_718; // @[Modules.scala 71:109:@30672.4]
  wire [11:0] _T_76646; // @[Modules.scala 71:109:@30674.4]
  wire [10:0] _T_76647; // @[Modules.scala 71:109:@30675.4]
  wire [10:0] buffer_12_719; // @[Modules.scala 71:109:@30676.4]
  wire [11:0] _T_76649; // @[Modules.scala 71:109:@30678.4]
  wire [10:0] _T_76650; // @[Modules.scala 71:109:@30679.4]
  wire [10:0] buffer_12_720; // @[Modules.scala 71:109:@30680.4]
  wire [11:0] _T_76652; // @[Modules.scala 71:109:@30682.4]
  wire [10:0] _T_76653; // @[Modules.scala 71:109:@30683.4]
  wire [10:0] buffer_12_721; // @[Modules.scala 71:109:@30684.4]
  wire [11:0] _T_76655; // @[Modules.scala 71:109:@30686.4]
  wire [10:0] _T_76656; // @[Modules.scala 71:109:@30687.4]
  wire [10:0] buffer_12_722; // @[Modules.scala 71:109:@30688.4]
  wire [11:0] _T_76658; // @[Modules.scala 71:109:@30690.4]
  wire [10:0] _T_76659; // @[Modules.scala 71:109:@30691.4]
  wire [10:0] buffer_12_723; // @[Modules.scala 71:109:@30692.4]
  wire [11:0] _T_76661; // @[Modules.scala 71:109:@30694.4]
  wire [10:0] _T_76662; // @[Modules.scala 71:109:@30695.4]
  wire [10:0] buffer_12_724; // @[Modules.scala 71:109:@30696.4]
  wire [11:0] _T_76664; // @[Modules.scala 71:109:@30698.4]
  wire [10:0] _T_76665; // @[Modules.scala 71:109:@30699.4]
  wire [10:0] buffer_12_725; // @[Modules.scala 71:109:@30700.4]
  wire [11:0] _T_76667; // @[Modules.scala 71:109:@30702.4]
  wire [10:0] _T_76668; // @[Modules.scala 71:109:@30703.4]
  wire [10:0] buffer_12_726; // @[Modules.scala 71:109:@30704.4]
  wire [11:0] _T_76670; // @[Modules.scala 71:109:@30706.4]
  wire [10:0] _T_76671; // @[Modules.scala 71:109:@30707.4]
  wire [10:0] buffer_12_727; // @[Modules.scala 71:109:@30708.4]
  wire [11:0] _T_76673; // @[Modules.scala 71:109:@30710.4]
  wire [10:0] _T_76674; // @[Modules.scala 71:109:@30711.4]
  wire [10:0] buffer_12_728; // @[Modules.scala 71:109:@30712.4]
  wire [11:0] _T_76676; // @[Modules.scala 71:109:@30714.4]
  wire [10:0] _T_76677; // @[Modules.scala 71:109:@30715.4]
  wire [10:0] buffer_12_729; // @[Modules.scala 71:109:@30716.4]
  wire [11:0] _T_76682; // @[Modules.scala 71:109:@30722.4]
  wire [10:0] _T_76683; // @[Modules.scala 71:109:@30723.4]
  wire [10:0] buffer_12_731; // @[Modules.scala 71:109:@30724.4]
  wire [11:0] _T_76688; // @[Modules.scala 71:109:@30730.4]
  wire [10:0] _T_76689; // @[Modules.scala 71:109:@30731.4]
  wire [10:0] buffer_12_733; // @[Modules.scala 71:109:@30732.4]
  wire [11:0] _T_76691; // @[Modules.scala 71:109:@30734.4]
  wire [10:0] _T_76692; // @[Modules.scala 71:109:@30735.4]
  wire [10:0] buffer_12_734; // @[Modules.scala 71:109:@30736.4]
  wire [11:0] _T_76694; // @[Modules.scala 78:156:@30739.4]
  wire [10:0] _T_76695; // @[Modules.scala 78:156:@30740.4]
  wire [10:0] buffer_12_736; // @[Modules.scala 78:156:@30741.4]
  wire [11:0] _T_76697; // @[Modules.scala 78:156:@30743.4]
  wire [10:0] _T_76698; // @[Modules.scala 78:156:@30744.4]
  wire [10:0] buffer_12_737; // @[Modules.scala 78:156:@30745.4]
  wire [11:0] _T_76700; // @[Modules.scala 78:156:@30747.4]
  wire [10:0] _T_76701; // @[Modules.scala 78:156:@30748.4]
  wire [10:0] buffer_12_738; // @[Modules.scala 78:156:@30749.4]
  wire [11:0] _T_76703; // @[Modules.scala 78:156:@30751.4]
  wire [10:0] _T_76704; // @[Modules.scala 78:156:@30752.4]
  wire [10:0] buffer_12_739; // @[Modules.scala 78:156:@30753.4]
  wire [11:0] _T_76706; // @[Modules.scala 78:156:@30755.4]
  wire [10:0] _T_76707; // @[Modules.scala 78:156:@30756.4]
  wire [10:0] buffer_12_740; // @[Modules.scala 78:156:@30757.4]
  wire [11:0] _T_76709; // @[Modules.scala 78:156:@30759.4]
  wire [10:0] _T_76710; // @[Modules.scala 78:156:@30760.4]
  wire [10:0] buffer_12_741; // @[Modules.scala 78:156:@30761.4]
  wire [11:0] _T_76712; // @[Modules.scala 78:156:@30763.4]
  wire [10:0] _T_76713; // @[Modules.scala 78:156:@30764.4]
  wire [10:0] buffer_12_742; // @[Modules.scala 78:156:@30765.4]
  wire [11:0] _T_76715; // @[Modules.scala 78:156:@30767.4]
  wire [10:0] _T_76716; // @[Modules.scala 78:156:@30768.4]
  wire [10:0] buffer_12_743; // @[Modules.scala 78:156:@30769.4]
  wire [11:0] _T_76718; // @[Modules.scala 78:156:@30771.4]
  wire [10:0] _T_76719; // @[Modules.scala 78:156:@30772.4]
  wire [10:0] buffer_12_744; // @[Modules.scala 78:156:@30773.4]
  wire [11:0] _T_76721; // @[Modules.scala 78:156:@30775.4]
  wire [10:0] _T_76722; // @[Modules.scala 78:156:@30776.4]
  wire [10:0] buffer_12_745; // @[Modules.scala 78:156:@30777.4]
  wire [11:0] _T_76724; // @[Modules.scala 78:156:@30779.4]
  wire [10:0] _T_76725; // @[Modules.scala 78:156:@30780.4]
  wire [10:0] buffer_12_746; // @[Modules.scala 78:156:@30781.4]
  wire [11:0] _T_76727; // @[Modules.scala 78:156:@30783.4]
  wire [10:0] _T_76728; // @[Modules.scala 78:156:@30784.4]
  wire [10:0] buffer_12_747; // @[Modules.scala 78:156:@30785.4]
  wire [11:0] _T_76730; // @[Modules.scala 78:156:@30787.4]
  wire [10:0] _T_76731; // @[Modules.scala 78:156:@30788.4]
  wire [10:0] buffer_12_748; // @[Modules.scala 78:156:@30789.4]
  wire [11:0] _T_76733; // @[Modules.scala 78:156:@30791.4]
  wire [10:0] _T_76734; // @[Modules.scala 78:156:@30792.4]
  wire [10:0] buffer_12_749; // @[Modules.scala 78:156:@30793.4]
  wire [11:0] _T_76736; // @[Modules.scala 78:156:@30795.4]
  wire [10:0] _T_76737; // @[Modules.scala 78:156:@30796.4]
  wire [10:0] buffer_12_750; // @[Modules.scala 78:156:@30797.4]
  wire [11:0] _T_76739; // @[Modules.scala 78:156:@30799.4]
  wire [10:0] _T_76740; // @[Modules.scala 78:156:@30800.4]
  wire [10:0] buffer_12_751; // @[Modules.scala 78:156:@30801.4]
  wire [11:0] _T_76742; // @[Modules.scala 78:156:@30803.4]
  wire [10:0] _T_76743; // @[Modules.scala 78:156:@30804.4]
  wire [10:0] buffer_12_752; // @[Modules.scala 78:156:@30805.4]
  wire [11:0] _T_76745; // @[Modules.scala 78:156:@30807.4]
  wire [10:0] _T_76746; // @[Modules.scala 78:156:@30808.4]
  wire [10:0] buffer_12_753; // @[Modules.scala 78:156:@30809.4]
  wire [11:0] _T_76748; // @[Modules.scala 78:156:@30811.4]
  wire [10:0] _T_76749; // @[Modules.scala 78:156:@30812.4]
  wire [10:0] buffer_12_754; // @[Modules.scala 78:156:@30813.4]
  wire [11:0] _T_76751; // @[Modules.scala 78:156:@30815.4]
  wire [10:0] _T_76752; // @[Modules.scala 78:156:@30816.4]
  wire [10:0] buffer_12_755; // @[Modules.scala 78:156:@30817.4]
  wire [11:0] _T_76754; // @[Modules.scala 78:156:@30819.4]
  wire [10:0] _T_76755; // @[Modules.scala 78:156:@30820.4]
  wire [10:0] buffer_12_756; // @[Modules.scala 78:156:@30821.4]
  wire [11:0] _T_76757; // @[Modules.scala 78:156:@30823.4]
  wire [10:0] _T_76758; // @[Modules.scala 78:156:@30824.4]
  wire [10:0] buffer_12_757; // @[Modules.scala 78:156:@30825.4]
  wire [11:0] _T_76760; // @[Modules.scala 78:156:@30827.4]
  wire [10:0] _T_76761; // @[Modules.scala 78:156:@30828.4]
  wire [10:0] buffer_12_758; // @[Modules.scala 78:156:@30829.4]
  wire [11:0] _T_76763; // @[Modules.scala 78:156:@30831.4]
  wire [10:0] _T_76764; // @[Modules.scala 78:156:@30832.4]
  wire [10:0] buffer_12_759; // @[Modules.scala 78:156:@30833.4]
  wire [11:0] _T_76766; // @[Modules.scala 78:156:@30835.4]
  wire [10:0] _T_76767; // @[Modules.scala 78:156:@30836.4]
  wire [10:0] buffer_12_760; // @[Modules.scala 78:156:@30837.4]
  wire [11:0] _T_76769; // @[Modules.scala 78:156:@30839.4]
  wire [10:0] _T_76770; // @[Modules.scala 78:156:@30840.4]
  wire [10:0] buffer_12_761; // @[Modules.scala 78:156:@30841.4]
  wire [11:0] _T_76772; // @[Modules.scala 78:156:@30843.4]
  wire [10:0] _T_76773; // @[Modules.scala 78:156:@30844.4]
  wire [10:0] buffer_12_762; // @[Modules.scala 78:156:@30845.4]
  wire [11:0] _T_76775; // @[Modules.scala 78:156:@30847.4]
  wire [10:0] _T_76776; // @[Modules.scala 78:156:@30848.4]
  wire [10:0] buffer_12_763; // @[Modules.scala 78:156:@30849.4]
  wire [11:0] _T_76778; // @[Modules.scala 78:156:@30851.4]
  wire [10:0] _T_76779; // @[Modules.scala 78:156:@30852.4]
  wire [10:0] buffer_12_764; // @[Modules.scala 78:156:@30853.4]
  wire [11:0] _T_76781; // @[Modules.scala 78:156:@30855.4]
  wire [10:0] _T_76782; // @[Modules.scala 78:156:@30856.4]
  wire [10:0] buffer_12_765; // @[Modules.scala 78:156:@30857.4]
  wire [11:0] _T_76784; // @[Modules.scala 78:156:@30859.4]
  wire [10:0] _T_76785; // @[Modules.scala 78:156:@30860.4]
  wire [10:0] buffer_12_766; // @[Modules.scala 78:156:@30861.4]
  wire [11:0] _T_76787; // @[Modules.scala 78:156:@30863.4]
  wire [10:0] _T_76788; // @[Modules.scala 78:156:@30864.4]
  wire [10:0] buffer_12_767; // @[Modules.scala 78:156:@30865.4]
  wire [11:0] _T_76790; // @[Modules.scala 78:156:@30867.4]
  wire [10:0] _T_76791; // @[Modules.scala 78:156:@30868.4]
  wire [10:0] buffer_12_768; // @[Modules.scala 78:156:@30869.4]
  wire [11:0] _T_76793; // @[Modules.scala 78:156:@30871.4]
  wire [10:0] _T_76794; // @[Modules.scala 78:156:@30872.4]
  wire [10:0] buffer_12_769; // @[Modules.scala 78:156:@30873.4]
  wire [11:0] _T_76796; // @[Modules.scala 78:156:@30875.4]
  wire [10:0] _T_76797; // @[Modules.scala 78:156:@30876.4]
  wire [10:0] buffer_12_770; // @[Modules.scala 78:156:@30877.4]
  wire [11:0] _T_76799; // @[Modules.scala 78:156:@30879.4]
  wire [10:0] _T_76800; // @[Modules.scala 78:156:@30880.4]
  wire [10:0] buffer_12_771; // @[Modules.scala 78:156:@30881.4]
  wire [11:0] _T_76802; // @[Modules.scala 78:156:@30883.4]
  wire [10:0] _T_76803; // @[Modules.scala 78:156:@30884.4]
  wire [10:0] buffer_12_772; // @[Modules.scala 78:156:@30885.4]
  wire [11:0] _T_76805; // @[Modules.scala 78:156:@30887.4]
  wire [10:0] _T_76806; // @[Modules.scala 78:156:@30888.4]
  wire [10:0] buffer_12_773; // @[Modules.scala 78:156:@30889.4]
  wire [11:0] _T_76808; // @[Modules.scala 78:156:@30891.4]
  wire [10:0] _T_76809; // @[Modules.scala 78:156:@30892.4]
  wire [10:0] buffer_12_774; // @[Modules.scala 78:156:@30893.4]
  wire [11:0] _T_76811; // @[Modules.scala 78:156:@30895.4]
  wire [10:0] _T_76812; // @[Modules.scala 78:156:@30896.4]
  wire [10:0] buffer_12_775; // @[Modules.scala 78:156:@30897.4]
  wire [11:0] _T_76814; // @[Modules.scala 78:156:@30899.4]
  wire [10:0] _T_76815; // @[Modules.scala 78:156:@30900.4]
  wire [10:0] buffer_12_776; // @[Modules.scala 78:156:@30901.4]
  wire [11:0] _T_76817; // @[Modules.scala 78:156:@30903.4]
  wire [10:0] _T_76818; // @[Modules.scala 78:156:@30904.4]
  wire [10:0] buffer_12_777; // @[Modules.scala 78:156:@30905.4]
  wire [11:0] _T_76820; // @[Modules.scala 78:156:@30907.4]
  wire [10:0] _T_76821; // @[Modules.scala 78:156:@30908.4]
  wire [10:0] buffer_12_778; // @[Modules.scala 78:156:@30909.4]
  wire [11:0] _T_76823; // @[Modules.scala 78:156:@30911.4]
  wire [10:0] _T_76824; // @[Modules.scala 78:156:@30912.4]
  wire [10:0] buffer_12_779; // @[Modules.scala 78:156:@30913.4]
  wire [11:0] _T_76826; // @[Modules.scala 78:156:@30915.4]
  wire [10:0] _T_76827; // @[Modules.scala 78:156:@30916.4]
  wire [10:0] buffer_12_780; // @[Modules.scala 78:156:@30917.4]
  wire [11:0] _T_76829; // @[Modules.scala 78:156:@30919.4]
  wire [10:0] _T_76830; // @[Modules.scala 78:156:@30920.4]
  wire [10:0] buffer_12_781; // @[Modules.scala 78:156:@30921.4]
  wire [11:0] _T_76832; // @[Modules.scala 78:156:@30923.4]
  wire [10:0] _T_76833; // @[Modules.scala 78:156:@30924.4]
  wire [10:0] buffer_12_782; // @[Modules.scala 78:156:@30925.4]
  wire [11:0] _T_76835; // @[Modules.scala 78:156:@30927.4]
  wire [10:0] _T_76836; // @[Modules.scala 78:156:@30928.4]
  wire [10:0] buffer_12_783; // @[Modules.scala 78:156:@30929.4]
  wire [11:0] _T_77356; // @[Modules.scala 65:57:@31693.4]
  wire [10:0] _T_77357; // @[Modules.scala 65:57:@31694.4]
  wire [10:0] buffer_13_392; // @[Modules.scala 65:57:@31695.4]
  wire [10:0] buffer_13_6; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77365; // @[Modules.scala 65:57:@31705.4]
  wire [10:0] _T_77366; // @[Modules.scala 65:57:@31706.4]
  wire [10:0] buffer_13_395; // @[Modules.scala 65:57:@31707.4]
  wire [11:0] _T_77377; // @[Modules.scala 65:57:@31721.4]
  wire [10:0] _T_77378; // @[Modules.scala 65:57:@31722.4]
  wire [10:0] buffer_13_399; // @[Modules.scala 65:57:@31723.4]
  wire [10:0] buffer_13_18; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77383; // @[Modules.scala 65:57:@31729.4]
  wire [10:0] _T_77384; // @[Modules.scala 65:57:@31730.4]
  wire [10:0] buffer_13_401; // @[Modules.scala 65:57:@31731.4]
  wire [11:0] _T_77395; // @[Modules.scala 65:57:@31745.4]
  wire [10:0] _T_77396; // @[Modules.scala 65:57:@31746.4]
  wire [10:0] buffer_13_405; // @[Modules.scala 65:57:@31747.4]
  wire [10:0] buffer_13_35; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77407; // @[Modules.scala 65:57:@31761.4]
  wire [10:0] _T_77408; // @[Modules.scala 65:57:@31762.4]
  wire [10:0] buffer_13_409; // @[Modules.scala 65:57:@31763.4]
  wire [11:0] _T_77410; // @[Modules.scala 65:57:@31765.4]
  wire [10:0] _T_77411; // @[Modules.scala 65:57:@31766.4]
  wire [10:0] buffer_13_410; // @[Modules.scala 65:57:@31767.4]
  wire [10:0] buffer_13_40; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77416; // @[Modules.scala 65:57:@31773.4]
  wire [10:0] _T_77417; // @[Modules.scala 65:57:@31774.4]
  wire [10:0] buffer_13_412; // @[Modules.scala 65:57:@31775.4]
  wire [11:0] _T_77428; // @[Modules.scala 65:57:@31789.4]
  wire [10:0] _T_77429; // @[Modules.scala 65:57:@31790.4]
  wire [10:0] buffer_13_416; // @[Modules.scala 65:57:@31791.4]
  wire [11:0] _T_77446; // @[Modules.scala 65:57:@31813.4]
  wire [10:0] _T_77447; // @[Modules.scala 65:57:@31814.4]
  wire [10:0] buffer_13_422; // @[Modules.scala 65:57:@31815.4]
  wire [10:0] buffer_13_79; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77473; // @[Modules.scala 65:57:@31849.4]
  wire [10:0] _T_77474; // @[Modules.scala 65:57:@31850.4]
  wire [10:0] buffer_13_431; // @[Modules.scala 65:57:@31851.4]
  wire [11:0] _T_77476; // @[Modules.scala 65:57:@31853.4]
  wire [10:0] _T_77477; // @[Modules.scala 65:57:@31854.4]
  wire [10:0] buffer_13_432; // @[Modules.scala 65:57:@31855.4]
  wire [10:0] buffer_13_85; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77482; // @[Modules.scala 65:57:@31861.4]
  wire [10:0] _T_77483; // @[Modules.scala 65:57:@31862.4]
  wire [10:0] buffer_13_434; // @[Modules.scala 65:57:@31863.4]
  wire [10:0] buffer_13_90; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77491; // @[Modules.scala 65:57:@31873.4]
  wire [10:0] _T_77492; // @[Modules.scala 65:57:@31874.4]
  wire [10:0] buffer_13_437; // @[Modules.scala 65:57:@31875.4]
  wire [10:0] buffer_13_93; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77494; // @[Modules.scala 65:57:@31877.4]
  wire [10:0] _T_77495; // @[Modules.scala 65:57:@31878.4]
  wire [10:0] buffer_13_438; // @[Modules.scala 65:57:@31879.4]
  wire [11:0] _T_77497; // @[Modules.scala 65:57:@31881.4]
  wire [10:0] _T_77498; // @[Modules.scala 65:57:@31882.4]
  wire [10:0] buffer_13_439; // @[Modules.scala 65:57:@31883.4]
  wire [11:0] _T_77503; // @[Modules.scala 65:57:@31889.4]
  wire [10:0] _T_77504; // @[Modules.scala 65:57:@31890.4]
  wire [10:0] buffer_13_441; // @[Modules.scala 65:57:@31891.4]
  wire [11:0] _T_77506; // @[Modules.scala 65:57:@31893.4]
  wire [10:0] _T_77507; // @[Modules.scala 65:57:@31894.4]
  wire [10:0] buffer_13_442; // @[Modules.scala 65:57:@31895.4]
  wire [11:0] _T_77512; // @[Modules.scala 65:57:@31901.4]
  wire [10:0] _T_77513; // @[Modules.scala 65:57:@31902.4]
  wire [10:0] buffer_13_444; // @[Modules.scala 65:57:@31903.4]
  wire [11:0] _T_77524; // @[Modules.scala 65:57:@31917.4]
  wire [10:0] _T_77525; // @[Modules.scala 65:57:@31918.4]
  wire [10:0] buffer_13_448; // @[Modules.scala 65:57:@31919.4]
  wire [11:0] _T_77527; // @[Modules.scala 65:57:@31921.4]
  wire [10:0] _T_77528; // @[Modules.scala 65:57:@31922.4]
  wire [10:0] buffer_13_449; // @[Modules.scala 65:57:@31923.4]
  wire [10:0] buffer_13_120; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77536; // @[Modules.scala 65:57:@31933.4]
  wire [10:0] _T_77537; // @[Modules.scala 65:57:@31934.4]
  wire [10:0] buffer_13_452; // @[Modules.scala 65:57:@31935.4]
  wire [11:0] _T_77551; // @[Modules.scala 65:57:@31953.4]
  wire [10:0] _T_77552; // @[Modules.scala 65:57:@31954.4]
  wire [10:0] buffer_13_457; // @[Modules.scala 65:57:@31955.4]
  wire [10:0] buffer_13_132; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77554; // @[Modules.scala 65:57:@31957.4]
  wire [10:0] _T_77555; // @[Modules.scala 65:57:@31958.4]
  wire [10:0] buffer_13_458; // @[Modules.scala 65:57:@31959.4]
  wire [11:0] _T_77560; // @[Modules.scala 65:57:@31965.4]
  wire [10:0] _T_77561; // @[Modules.scala 65:57:@31966.4]
  wire [10:0] buffer_13_460; // @[Modules.scala 65:57:@31967.4]
  wire [10:0] buffer_13_145; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77572; // @[Modules.scala 65:57:@31981.4]
  wire [10:0] _T_77573; // @[Modules.scala 65:57:@31982.4]
  wire [10:0] buffer_13_464; // @[Modules.scala 65:57:@31983.4]
  wire [11:0] _T_77578; // @[Modules.scala 65:57:@31989.4]
  wire [10:0] _T_77579; // @[Modules.scala 65:57:@31990.4]
  wire [10:0] buffer_13_466; // @[Modules.scala 65:57:@31991.4]
  wire [11:0] _T_77581; // @[Modules.scala 65:57:@31993.4]
  wire [10:0] _T_77582; // @[Modules.scala 65:57:@31994.4]
  wire [10:0] buffer_13_467; // @[Modules.scala 65:57:@31995.4]
  wire [11:0] _T_77590; // @[Modules.scala 65:57:@32005.4]
  wire [10:0] _T_77591; // @[Modules.scala 65:57:@32006.4]
  wire [10:0] buffer_13_470; // @[Modules.scala 65:57:@32007.4]
  wire [10:0] buffer_13_158; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77593; // @[Modules.scala 65:57:@32009.4]
  wire [10:0] _T_77594; // @[Modules.scala 65:57:@32010.4]
  wire [10:0] buffer_13_471; // @[Modules.scala 65:57:@32011.4]
  wire [11:0] _T_77599; // @[Modules.scala 65:57:@32017.4]
  wire [10:0] _T_77600; // @[Modules.scala 65:57:@32018.4]
  wire [10:0] buffer_13_473; // @[Modules.scala 65:57:@32019.4]
  wire [11:0] _T_77608; // @[Modules.scala 65:57:@32029.4]
  wire [10:0] _T_77609; // @[Modules.scala 65:57:@32030.4]
  wire [10:0] buffer_13_476; // @[Modules.scala 65:57:@32031.4]
  wire [10:0] buffer_13_171; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77611; // @[Modules.scala 65:57:@32033.4]
  wire [10:0] _T_77612; // @[Modules.scala 65:57:@32034.4]
  wire [10:0] buffer_13_477; // @[Modules.scala 65:57:@32035.4]
  wire [10:0] buffer_13_172; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77614; // @[Modules.scala 65:57:@32037.4]
  wire [10:0] _T_77615; // @[Modules.scala 65:57:@32038.4]
  wire [10:0] buffer_13_478; // @[Modules.scala 65:57:@32039.4]
  wire [10:0] buffer_13_174; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77617; // @[Modules.scala 65:57:@32041.4]
  wire [10:0] _T_77618; // @[Modules.scala 65:57:@32042.4]
  wire [10:0] buffer_13_479; // @[Modules.scala 65:57:@32043.4]
  wire [10:0] buffer_13_176; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77620; // @[Modules.scala 65:57:@32045.4]
  wire [10:0] _T_77621; // @[Modules.scala 65:57:@32046.4]
  wire [10:0] buffer_13_480; // @[Modules.scala 65:57:@32047.4]
  wire [11:0] _T_77629; // @[Modules.scala 65:57:@32057.4]
  wire [10:0] _T_77630; // @[Modules.scala 65:57:@32058.4]
  wire [10:0] buffer_13_483; // @[Modules.scala 65:57:@32059.4]
  wire [11:0] _T_77635; // @[Modules.scala 65:57:@32065.4]
  wire [10:0] _T_77636; // @[Modules.scala 65:57:@32066.4]
  wire [10:0] buffer_13_485; // @[Modules.scala 65:57:@32067.4]
  wire [11:0] _T_77641; // @[Modules.scala 65:57:@32073.4]
  wire [10:0] _T_77642; // @[Modules.scala 65:57:@32074.4]
  wire [10:0] buffer_13_487; // @[Modules.scala 65:57:@32075.4]
  wire [11:0] _T_77644; // @[Modules.scala 65:57:@32077.4]
  wire [10:0] _T_77645; // @[Modules.scala 65:57:@32078.4]
  wire [10:0] buffer_13_488; // @[Modules.scala 65:57:@32079.4]
  wire [11:0] _T_77659; // @[Modules.scala 65:57:@32097.4]
  wire [10:0] _T_77660; // @[Modules.scala 65:57:@32098.4]
  wire [10:0] buffer_13_493; // @[Modules.scala 65:57:@32099.4]
  wire [11:0] _T_77662; // @[Modules.scala 65:57:@32101.4]
  wire [10:0] _T_77663; // @[Modules.scala 65:57:@32102.4]
  wire [10:0] buffer_13_494; // @[Modules.scala 65:57:@32103.4]
  wire [11:0] _T_77701; // @[Modules.scala 65:57:@32153.4]
  wire [10:0] _T_77702; // @[Modules.scala 65:57:@32154.4]
  wire [10:0] buffer_13_507; // @[Modules.scala 65:57:@32155.4]
  wire [11:0] _T_77704; // @[Modules.scala 65:57:@32157.4]
  wire [10:0] _T_77705; // @[Modules.scala 65:57:@32158.4]
  wire [10:0] buffer_13_508; // @[Modules.scala 65:57:@32159.4]
  wire [11:0] _T_77707; // @[Modules.scala 65:57:@32161.4]
  wire [10:0] _T_77708; // @[Modules.scala 65:57:@32162.4]
  wire [10:0] buffer_13_509; // @[Modules.scala 65:57:@32163.4]
  wire [11:0] _T_77716; // @[Modules.scala 65:57:@32173.4]
  wire [10:0] _T_77717; // @[Modules.scala 65:57:@32174.4]
  wire [10:0] buffer_13_512; // @[Modules.scala 65:57:@32175.4]
  wire [11:0] _T_77725; // @[Modules.scala 65:57:@32185.4]
  wire [10:0] _T_77726; // @[Modules.scala 65:57:@32186.4]
  wire [10:0] buffer_13_515; // @[Modules.scala 65:57:@32187.4]
  wire [10:0] buffer_13_248; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77728; // @[Modules.scala 65:57:@32189.4]
  wire [10:0] _T_77729; // @[Modules.scala 65:57:@32190.4]
  wire [10:0] buffer_13_516; // @[Modules.scala 65:57:@32191.4]
  wire [11:0] _T_77746; // @[Modules.scala 65:57:@32213.4]
  wire [10:0] _T_77747; // @[Modules.scala 65:57:@32214.4]
  wire [10:0] buffer_13_522; // @[Modules.scala 65:57:@32215.4]
  wire [11:0] _T_77749; // @[Modules.scala 65:57:@32217.4]
  wire [10:0] _T_77750; // @[Modules.scala 65:57:@32218.4]
  wire [10:0] buffer_13_523; // @[Modules.scala 65:57:@32219.4]
  wire [10:0] buffer_13_265; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77752; // @[Modules.scala 65:57:@32221.4]
  wire [10:0] _T_77753; // @[Modules.scala 65:57:@32222.4]
  wire [10:0] buffer_13_524; // @[Modules.scala 65:57:@32223.4]
  wire [11:0] _T_77758; // @[Modules.scala 65:57:@32229.4]
  wire [10:0] _T_77759; // @[Modules.scala 65:57:@32230.4]
  wire [10:0] buffer_13_526; // @[Modules.scala 65:57:@32231.4]
  wire [11:0] _T_77764; // @[Modules.scala 65:57:@32237.4]
  wire [10:0] _T_77765; // @[Modules.scala 65:57:@32238.4]
  wire [10:0] buffer_13_528; // @[Modules.scala 65:57:@32239.4]
  wire [11:0] _T_77776; // @[Modules.scala 65:57:@32253.4]
  wire [10:0] _T_77777; // @[Modules.scala 65:57:@32254.4]
  wire [10:0] buffer_13_532; // @[Modules.scala 65:57:@32255.4]
  wire [10:0] buffer_13_282; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77779; // @[Modules.scala 65:57:@32257.4]
  wire [10:0] _T_77780; // @[Modules.scala 65:57:@32258.4]
  wire [10:0] buffer_13_533; // @[Modules.scala 65:57:@32259.4]
  wire [11:0] _T_77791; // @[Modules.scala 65:57:@32273.4]
  wire [10:0] _T_77792; // @[Modules.scala 65:57:@32274.4]
  wire [10:0] buffer_13_537; // @[Modules.scala 65:57:@32275.4]
  wire [11:0] _T_77794; // @[Modules.scala 65:57:@32277.4]
  wire [10:0] _T_77795; // @[Modules.scala 65:57:@32278.4]
  wire [10:0] buffer_13_538; // @[Modules.scala 65:57:@32279.4]
  wire [11:0] _T_77800; // @[Modules.scala 65:57:@32285.4]
  wire [10:0] _T_77801; // @[Modules.scala 65:57:@32286.4]
  wire [10:0] buffer_13_540; // @[Modules.scala 65:57:@32287.4]
  wire [10:0] buffer_13_309; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77818; // @[Modules.scala 65:57:@32309.4]
  wire [10:0] _T_77819; // @[Modules.scala 65:57:@32310.4]
  wire [10:0] buffer_13_546; // @[Modules.scala 65:57:@32311.4]
  wire [11:0] _T_77821; // @[Modules.scala 65:57:@32313.4]
  wire [10:0] _T_77822; // @[Modules.scala 65:57:@32314.4]
  wire [10:0] buffer_13_547; // @[Modules.scala 65:57:@32315.4]
  wire [11:0] _T_77824; // @[Modules.scala 65:57:@32317.4]
  wire [10:0] _T_77825; // @[Modules.scala 65:57:@32318.4]
  wire [10:0] buffer_13_548; // @[Modules.scala 65:57:@32319.4]
  wire [11:0] _T_77827; // @[Modules.scala 65:57:@32321.4]
  wire [10:0] _T_77828; // @[Modules.scala 65:57:@32322.4]
  wire [10:0] buffer_13_549; // @[Modules.scala 65:57:@32323.4]
  wire [11:0] _T_77830; // @[Modules.scala 65:57:@32325.4]
  wire [10:0] _T_77831; // @[Modules.scala 65:57:@32326.4]
  wire [10:0] buffer_13_550; // @[Modules.scala 65:57:@32327.4]
  wire [11:0] _T_77836; // @[Modules.scala 65:57:@32333.4]
  wire [10:0] _T_77837; // @[Modules.scala 65:57:@32334.4]
  wire [10:0] buffer_13_552; // @[Modules.scala 65:57:@32335.4]
  wire [10:0] buffer_13_329; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77848; // @[Modules.scala 65:57:@32349.4]
  wire [10:0] _T_77849; // @[Modules.scala 65:57:@32350.4]
  wire [10:0] buffer_13_556; // @[Modules.scala 65:57:@32351.4]
  wire [11:0] _T_77860; // @[Modules.scala 65:57:@32365.4]
  wire [10:0] _T_77861; // @[Modules.scala 65:57:@32366.4]
  wire [10:0] buffer_13_560; // @[Modules.scala 65:57:@32367.4]
  wire [11:0] _T_77869; // @[Modules.scala 65:57:@32377.4]
  wire [10:0] _T_77870; // @[Modules.scala 65:57:@32378.4]
  wire [10:0] buffer_13_563; // @[Modules.scala 65:57:@32379.4]
  wire [11:0] _T_77881; // @[Modules.scala 65:57:@32393.4]
  wire [10:0] _T_77882; // @[Modules.scala 65:57:@32394.4]
  wire [10:0] buffer_13_567; // @[Modules.scala 65:57:@32395.4]
  wire [11:0] _T_77902; // @[Modules.scala 65:57:@32421.4]
  wire [10:0] _T_77903; // @[Modules.scala 65:57:@32422.4]
  wire [10:0] buffer_13_574; // @[Modules.scala 65:57:@32423.4]
  wire [11:0] _T_77923; // @[Modules.scala 65:57:@32449.4]
  wire [10:0] _T_77924; // @[Modules.scala 65:57:@32450.4]
  wire [10:0] buffer_13_581; // @[Modules.scala 65:57:@32451.4]
  wire [10:0] buffer_13_391; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_77941; // @[Modules.scala 65:57:@32473.4]
  wire [10:0] _T_77942; // @[Modules.scala 65:57:@32474.4]
  wire [10:0] buffer_13_587; // @[Modules.scala 65:57:@32475.4]
  wire [11:0] _T_77944; // @[Modules.scala 68:83:@32477.4]
  wire [10:0] _T_77945; // @[Modules.scala 68:83:@32478.4]
  wire [10:0] buffer_13_588; // @[Modules.scala 68:83:@32479.4]
  wire [11:0] _T_77947; // @[Modules.scala 68:83:@32481.4]
  wire [10:0] _T_77948; // @[Modules.scala 68:83:@32482.4]
  wire [10:0] buffer_13_589; // @[Modules.scala 68:83:@32483.4]
  wire [11:0] _T_77950; // @[Modules.scala 68:83:@32485.4]
  wire [10:0] _T_77951; // @[Modules.scala 68:83:@32486.4]
  wire [10:0] buffer_13_590; // @[Modules.scala 68:83:@32487.4]
  wire [11:0] _T_77953; // @[Modules.scala 68:83:@32489.4]
  wire [10:0] _T_77954; // @[Modules.scala 68:83:@32490.4]
  wire [10:0] buffer_13_591; // @[Modules.scala 68:83:@32491.4]
  wire [11:0] _T_77956; // @[Modules.scala 68:83:@32493.4]
  wire [10:0] _T_77957; // @[Modules.scala 68:83:@32494.4]
  wire [10:0] buffer_13_592; // @[Modules.scala 68:83:@32495.4]
  wire [11:0] _T_77959; // @[Modules.scala 68:83:@32497.4]
  wire [10:0] _T_77960; // @[Modules.scala 68:83:@32498.4]
  wire [10:0] buffer_13_593; // @[Modules.scala 68:83:@32499.4]
  wire [11:0] _T_77962; // @[Modules.scala 68:83:@32501.4]
  wire [10:0] _T_77963; // @[Modules.scala 68:83:@32502.4]
  wire [10:0] buffer_13_594; // @[Modules.scala 68:83:@32503.4]
  wire [11:0] _T_77965; // @[Modules.scala 68:83:@32505.4]
  wire [10:0] _T_77966; // @[Modules.scala 68:83:@32506.4]
  wire [10:0] buffer_13_595; // @[Modules.scala 68:83:@32507.4]
  wire [11:0] _T_77968; // @[Modules.scala 68:83:@32509.4]
  wire [10:0] _T_77969; // @[Modules.scala 68:83:@32510.4]
  wire [10:0] buffer_13_596; // @[Modules.scala 68:83:@32511.4]
  wire [11:0] _T_77971; // @[Modules.scala 68:83:@32513.4]
  wire [10:0] _T_77972; // @[Modules.scala 68:83:@32514.4]
  wire [10:0] buffer_13_597; // @[Modules.scala 68:83:@32515.4]
  wire [11:0] _T_77974; // @[Modules.scala 68:83:@32517.4]
  wire [10:0] _T_77975; // @[Modules.scala 68:83:@32518.4]
  wire [10:0] buffer_13_598; // @[Modules.scala 68:83:@32519.4]
  wire [11:0] _T_77980; // @[Modules.scala 68:83:@32525.4]
  wire [10:0] _T_77981; // @[Modules.scala 68:83:@32526.4]
  wire [10:0] buffer_13_600; // @[Modules.scala 68:83:@32527.4]
  wire [11:0] _T_77986; // @[Modules.scala 68:83:@32533.4]
  wire [10:0] _T_77987; // @[Modules.scala 68:83:@32534.4]
  wire [10:0] buffer_13_602; // @[Modules.scala 68:83:@32535.4]
  wire [11:0] _T_77989; // @[Modules.scala 68:83:@32537.4]
  wire [10:0] _T_77990; // @[Modules.scala 68:83:@32538.4]
  wire [10:0] buffer_13_603; // @[Modules.scala 68:83:@32539.4]
  wire [11:0] _T_77995; // @[Modules.scala 68:83:@32545.4]
  wire [10:0] _T_77996; // @[Modules.scala 68:83:@32546.4]
  wire [10:0] buffer_13_605; // @[Modules.scala 68:83:@32547.4]
  wire [11:0] _T_77998; // @[Modules.scala 68:83:@32549.4]
  wire [10:0] _T_77999; // @[Modules.scala 68:83:@32550.4]
  wire [10:0] buffer_13_606; // @[Modules.scala 68:83:@32551.4]
  wire [11:0] _T_78001; // @[Modules.scala 68:83:@32553.4]
  wire [10:0] _T_78002; // @[Modules.scala 68:83:@32554.4]
  wire [10:0] buffer_13_607; // @[Modules.scala 68:83:@32555.4]
  wire [11:0] _T_78004; // @[Modules.scala 68:83:@32557.4]
  wire [10:0] _T_78005; // @[Modules.scala 68:83:@32558.4]
  wire [10:0] buffer_13_608; // @[Modules.scala 68:83:@32559.4]
  wire [11:0] _T_78007; // @[Modules.scala 68:83:@32561.4]
  wire [10:0] _T_78008; // @[Modules.scala 68:83:@32562.4]
  wire [10:0] buffer_13_609; // @[Modules.scala 68:83:@32563.4]
  wire [11:0] _T_78010; // @[Modules.scala 68:83:@32565.4]
  wire [10:0] _T_78011; // @[Modules.scala 68:83:@32566.4]
  wire [10:0] buffer_13_610; // @[Modules.scala 68:83:@32567.4]
  wire [11:0] _T_78013; // @[Modules.scala 68:83:@32569.4]
  wire [10:0] _T_78014; // @[Modules.scala 68:83:@32570.4]
  wire [10:0] buffer_13_611; // @[Modules.scala 68:83:@32571.4]
  wire [11:0] _T_78016; // @[Modules.scala 68:83:@32573.4]
  wire [10:0] _T_78017; // @[Modules.scala 68:83:@32574.4]
  wire [10:0] buffer_13_612; // @[Modules.scala 68:83:@32575.4]
  wire [11:0] _T_78019; // @[Modules.scala 68:83:@32577.4]
  wire [10:0] _T_78020; // @[Modules.scala 68:83:@32578.4]
  wire [10:0] buffer_13_613; // @[Modules.scala 68:83:@32579.4]
  wire [11:0] _T_78022; // @[Modules.scala 68:83:@32581.4]
  wire [10:0] _T_78023; // @[Modules.scala 68:83:@32582.4]
  wire [10:0] buffer_13_614; // @[Modules.scala 68:83:@32583.4]
  wire [11:0] _T_78025; // @[Modules.scala 68:83:@32585.4]
  wire [10:0] _T_78026; // @[Modules.scala 68:83:@32586.4]
  wire [10:0] buffer_13_615; // @[Modules.scala 68:83:@32587.4]
  wire [11:0] _T_78028; // @[Modules.scala 68:83:@32589.4]
  wire [10:0] _T_78029; // @[Modules.scala 68:83:@32590.4]
  wire [10:0] buffer_13_616; // @[Modules.scala 68:83:@32591.4]
  wire [11:0] _T_78031; // @[Modules.scala 68:83:@32593.4]
  wire [10:0] _T_78032; // @[Modules.scala 68:83:@32594.4]
  wire [10:0] buffer_13_617; // @[Modules.scala 68:83:@32595.4]
  wire [11:0] _T_78034; // @[Modules.scala 68:83:@32597.4]
  wire [10:0] _T_78035; // @[Modules.scala 68:83:@32598.4]
  wire [10:0] buffer_13_618; // @[Modules.scala 68:83:@32599.4]
  wire [11:0] _T_78040; // @[Modules.scala 68:83:@32605.4]
  wire [10:0] _T_78041; // @[Modules.scala 68:83:@32606.4]
  wire [10:0] buffer_13_620; // @[Modules.scala 68:83:@32607.4]
  wire [11:0] _T_78043; // @[Modules.scala 68:83:@32609.4]
  wire [10:0] _T_78044; // @[Modules.scala 68:83:@32610.4]
  wire [10:0] buffer_13_621; // @[Modules.scala 68:83:@32611.4]
  wire [11:0] _T_78046; // @[Modules.scala 68:83:@32613.4]
  wire [10:0] _T_78047; // @[Modules.scala 68:83:@32614.4]
  wire [10:0] buffer_13_622; // @[Modules.scala 68:83:@32615.4]
  wire [11:0] _T_78049; // @[Modules.scala 68:83:@32617.4]
  wire [10:0] _T_78050; // @[Modules.scala 68:83:@32618.4]
  wire [10:0] buffer_13_623; // @[Modules.scala 68:83:@32619.4]
  wire [11:0] _T_78052; // @[Modules.scala 68:83:@32621.4]
  wire [10:0] _T_78053; // @[Modules.scala 68:83:@32622.4]
  wire [10:0] buffer_13_624; // @[Modules.scala 68:83:@32623.4]
  wire [11:0] _T_78055; // @[Modules.scala 68:83:@32625.4]
  wire [10:0] _T_78056; // @[Modules.scala 68:83:@32626.4]
  wire [10:0] buffer_13_625; // @[Modules.scala 68:83:@32627.4]
  wire [11:0] _T_78061; // @[Modules.scala 68:83:@32633.4]
  wire [10:0] _T_78062; // @[Modules.scala 68:83:@32634.4]
  wire [10:0] buffer_13_627; // @[Modules.scala 68:83:@32635.4]
  wire [11:0] _T_78064; // @[Modules.scala 68:83:@32637.4]
  wire [10:0] _T_78065; // @[Modules.scala 68:83:@32638.4]
  wire [10:0] buffer_13_628; // @[Modules.scala 68:83:@32639.4]
  wire [11:0] _T_78067; // @[Modules.scala 68:83:@32641.4]
  wire [10:0] _T_78068; // @[Modules.scala 68:83:@32642.4]
  wire [10:0] buffer_13_629; // @[Modules.scala 68:83:@32643.4]
  wire [11:0] _T_78070; // @[Modules.scala 68:83:@32645.4]
  wire [10:0] _T_78071; // @[Modules.scala 68:83:@32646.4]
  wire [10:0] buffer_13_630; // @[Modules.scala 68:83:@32647.4]
  wire [11:0] _T_78073; // @[Modules.scala 68:83:@32649.4]
  wire [10:0] _T_78074; // @[Modules.scala 68:83:@32650.4]
  wire [10:0] buffer_13_631; // @[Modules.scala 68:83:@32651.4]
  wire [11:0] _T_78076; // @[Modules.scala 68:83:@32653.4]
  wire [10:0] _T_78077; // @[Modules.scala 68:83:@32654.4]
  wire [10:0] buffer_13_632; // @[Modules.scala 68:83:@32655.4]
  wire [11:0] _T_78079; // @[Modules.scala 68:83:@32657.4]
  wire [10:0] _T_78080; // @[Modules.scala 68:83:@32658.4]
  wire [10:0] buffer_13_633; // @[Modules.scala 68:83:@32659.4]
  wire [11:0] _T_78082; // @[Modules.scala 68:83:@32661.4]
  wire [10:0] _T_78083; // @[Modules.scala 68:83:@32662.4]
  wire [10:0] buffer_13_634; // @[Modules.scala 68:83:@32663.4]
  wire [11:0] _T_78085; // @[Modules.scala 68:83:@32665.4]
  wire [10:0] _T_78086; // @[Modules.scala 68:83:@32666.4]
  wire [10:0] buffer_13_635; // @[Modules.scala 68:83:@32667.4]
  wire [11:0] _T_78088; // @[Modules.scala 68:83:@32669.4]
  wire [10:0] _T_78089; // @[Modules.scala 68:83:@32670.4]
  wire [10:0] buffer_13_636; // @[Modules.scala 68:83:@32671.4]
  wire [11:0] _T_78091; // @[Modules.scala 68:83:@32673.4]
  wire [10:0] _T_78092; // @[Modules.scala 68:83:@32674.4]
  wire [10:0] buffer_13_637; // @[Modules.scala 68:83:@32675.4]
  wire [11:0] _T_78094; // @[Modules.scala 68:83:@32677.4]
  wire [10:0] _T_78095; // @[Modules.scala 68:83:@32678.4]
  wire [10:0] buffer_13_638; // @[Modules.scala 68:83:@32679.4]
  wire [11:0] _T_78097; // @[Modules.scala 68:83:@32681.4]
  wire [10:0] _T_78098; // @[Modules.scala 68:83:@32682.4]
  wire [10:0] buffer_13_639; // @[Modules.scala 68:83:@32683.4]
  wire [11:0] _T_78100; // @[Modules.scala 68:83:@32685.4]
  wire [10:0] _T_78101; // @[Modules.scala 68:83:@32686.4]
  wire [10:0] buffer_13_640; // @[Modules.scala 68:83:@32687.4]
  wire [11:0] _T_78103; // @[Modules.scala 68:83:@32689.4]
  wire [10:0] _T_78104; // @[Modules.scala 68:83:@32690.4]
  wire [10:0] buffer_13_641; // @[Modules.scala 68:83:@32691.4]
  wire [11:0] _T_78106; // @[Modules.scala 68:83:@32693.4]
  wire [10:0] _T_78107; // @[Modules.scala 68:83:@32694.4]
  wire [10:0] buffer_13_642; // @[Modules.scala 68:83:@32695.4]
  wire [11:0] _T_78109; // @[Modules.scala 68:83:@32697.4]
  wire [10:0] _T_78110; // @[Modules.scala 68:83:@32698.4]
  wire [10:0] buffer_13_643; // @[Modules.scala 68:83:@32699.4]
  wire [11:0] _T_78112; // @[Modules.scala 68:83:@32701.4]
  wire [10:0] _T_78113; // @[Modules.scala 68:83:@32702.4]
  wire [10:0] buffer_13_644; // @[Modules.scala 68:83:@32703.4]
  wire [11:0] _T_78115; // @[Modules.scala 68:83:@32705.4]
  wire [10:0] _T_78116; // @[Modules.scala 68:83:@32706.4]
  wire [10:0] buffer_13_645; // @[Modules.scala 68:83:@32707.4]
  wire [11:0] _T_78118; // @[Modules.scala 68:83:@32709.4]
  wire [10:0] _T_78119; // @[Modules.scala 68:83:@32710.4]
  wire [10:0] buffer_13_646; // @[Modules.scala 68:83:@32711.4]
  wire [11:0] _T_78124; // @[Modules.scala 68:83:@32717.4]
  wire [10:0] _T_78125; // @[Modules.scala 68:83:@32718.4]
  wire [10:0] buffer_13_648; // @[Modules.scala 68:83:@32719.4]
  wire [11:0] _T_78127; // @[Modules.scala 68:83:@32721.4]
  wire [10:0] _T_78128; // @[Modules.scala 68:83:@32722.4]
  wire [10:0] buffer_13_649; // @[Modules.scala 68:83:@32723.4]
  wire [11:0] _T_78130; // @[Modules.scala 68:83:@32725.4]
  wire [10:0] _T_78131; // @[Modules.scala 68:83:@32726.4]
  wire [10:0] buffer_13_650; // @[Modules.scala 68:83:@32727.4]
  wire [11:0] _T_78139; // @[Modules.scala 68:83:@32737.4]
  wire [10:0] _T_78140; // @[Modules.scala 68:83:@32738.4]
  wire [10:0] buffer_13_653; // @[Modules.scala 68:83:@32739.4]
  wire [11:0] _T_78142; // @[Modules.scala 68:83:@32741.4]
  wire [10:0] _T_78143; // @[Modules.scala 68:83:@32742.4]
  wire [10:0] buffer_13_654; // @[Modules.scala 68:83:@32743.4]
  wire [11:0] _T_78145; // @[Modules.scala 68:83:@32745.4]
  wire [10:0] _T_78146; // @[Modules.scala 68:83:@32746.4]
  wire [10:0] buffer_13_655; // @[Modules.scala 68:83:@32747.4]
  wire [11:0] _T_78148; // @[Modules.scala 68:83:@32749.4]
  wire [10:0] _T_78149; // @[Modules.scala 68:83:@32750.4]
  wire [10:0] buffer_13_656; // @[Modules.scala 68:83:@32751.4]
  wire [11:0] _T_78154; // @[Modules.scala 68:83:@32757.4]
  wire [10:0] _T_78155; // @[Modules.scala 68:83:@32758.4]
  wire [10:0] buffer_13_658; // @[Modules.scala 68:83:@32759.4]
  wire [11:0] _T_78160; // @[Modules.scala 68:83:@32765.4]
  wire [10:0] _T_78161; // @[Modules.scala 68:83:@32766.4]
  wire [10:0] buffer_13_660; // @[Modules.scala 68:83:@32767.4]
  wire [11:0] _T_78163; // @[Modules.scala 68:83:@32769.4]
  wire [10:0] _T_78164; // @[Modules.scala 68:83:@32770.4]
  wire [10:0] buffer_13_661; // @[Modules.scala 68:83:@32771.4]
  wire [11:0] _T_78166; // @[Modules.scala 68:83:@32773.4]
  wire [10:0] _T_78167; // @[Modules.scala 68:83:@32774.4]
  wire [10:0] buffer_13_662; // @[Modules.scala 68:83:@32775.4]
  wire [11:0] _T_78175; // @[Modules.scala 68:83:@32785.4]
  wire [10:0] _T_78176; // @[Modules.scala 68:83:@32786.4]
  wire [10:0] buffer_13_665; // @[Modules.scala 68:83:@32787.4]
  wire [11:0] _T_78178; // @[Modules.scala 68:83:@32789.4]
  wire [10:0] _T_78179; // @[Modules.scala 68:83:@32790.4]
  wire [10:0] buffer_13_666; // @[Modules.scala 68:83:@32791.4]
  wire [11:0] _T_78181; // @[Modules.scala 68:83:@32793.4]
  wire [10:0] _T_78182; // @[Modules.scala 68:83:@32794.4]
  wire [10:0] buffer_13_667; // @[Modules.scala 68:83:@32795.4]
  wire [11:0] _T_78184; // @[Modules.scala 68:83:@32797.4]
  wire [10:0] _T_78185; // @[Modules.scala 68:83:@32798.4]
  wire [10:0] buffer_13_668; // @[Modules.scala 68:83:@32799.4]
  wire [11:0] _T_78190; // @[Modules.scala 68:83:@32805.4]
  wire [10:0] _T_78191; // @[Modules.scala 68:83:@32806.4]
  wire [10:0] buffer_13_670; // @[Modules.scala 68:83:@32807.4]
  wire [11:0] _T_78196; // @[Modules.scala 68:83:@32813.4]
  wire [10:0] _T_78197; // @[Modules.scala 68:83:@32814.4]
  wire [10:0] buffer_13_672; // @[Modules.scala 68:83:@32815.4]
  wire [11:0] _T_78199; // @[Modules.scala 68:83:@32817.4]
  wire [10:0] _T_78200; // @[Modules.scala 68:83:@32818.4]
  wire [10:0] buffer_13_673; // @[Modules.scala 68:83:@32819.4]
  wire [11:0] _T_78205; // @[Modules.scala 68:83:@32825.4]
  wire [10:0] _T_78206; // @[Modules.scala 68:83:@32826.4]
  wire [10:0] buffer_13_675; // @[Modules.scala 68:83:@32827.4]
  wire [11:0] _T_78217; // @[Modules.scala 68:83:@32841.4]
  wire [10:0] _T_78218; // @[Modules.scala 68:83:@32842.4]
  wire [10:0] buffer_13_679; // @[Modules.scala 68:83:@32843.4]
  wire [11:0] _T_78226; // @[Modules.scala 68:83:@32853.4]
  wire [10:0] _T_78227; // @[Modules.scala 68:83:@32854.4]
  wire [10:0] buffer_13_682; // @[Modules.scala 68:83:@32855.4]
  wire [11:0] _T_78235; // @[Modules.scala 68:83:@32865.4]
  wire [10:0] _T_78236; // @[Modules.scala 68:83:@32866.4]
  wire [10:0] buffer_13_685; // @[Modules.scala 68:83:@32867.4]
  wire [11:0] _T_78238; // @[Modules.scala 71:109:@32869.4]
  wire [10:0] _T_78239; // @[Modules.scala 71:109:@32870.4]
  wire [10:0] buffer_13_686; // @[Modules.scala 71:109:@32871.4]
  wire [11:0] _T_78241; // @[Modules.scala 71:109:@32873.4]
  wire [10:0] _T_78242; // @[Modules.scala 71:109:@32874.4]
  wire [10:0] buffer_13_687; // @[Modules.scala 71:109:@32875.4]
  wire [11:0] _T_78244; // @[Modules.scala 71:109:@32877.4]
  wire [10:0] _T_78245; // @[Modules.scala 71:109:@32878.4]
  wire [10:0] buffer_13_688; // @[Modules.scala 71:109:@32879.4]
  wire [11:0] _T_78247; // @[Modules.scala 71:109:@32881.4]
  wire [10:0] _T_78248; // @[Modules.scala 71:109:@32882.4]
  wire [10:0] buffer_13_689; // @[Modules.scala 71:109:@32883.4]
  wire [11:0] _T_78250; // @[Modules.scala 71:109:@32885.4]
  wire [10:0] _T_78251; // @[Modules.scala 71:109:@32886.4]
  wire [10:0] buffer_13_690; // @[Modules.scala 71:109:@32887.4]
  wire [11:0] _T_78253; // @[Modules.scala 71:109:@32889.4]
  wire [10:0] _T_78254; // @[Modules.scala 71:109:@32890.4]
  wire [10:0] buffer_13_691; // @[Modules.scala 71:109:@32891.4]
  wire [11:0] _T_78256; // @[Modules.scala 71:109:@32893.4]
  wire [10:0] _T_78257; // @[Modules.scala 71:109:@32894.4]
  wire [10:0] buffer_13_692; // @[Modules.scala 71:109:@32895.4]
  wire [11:0] _T_78259; // @[Modules.scala 71:109:@32897.4]
  wire [10:0] _T_78260; // @[Modules.scala 71:109:@32898.4]
  wire [10:0] buffer_13_693; // @[Modules.scala 71:109:@32899.4]
  wire [11:0] _T_78262; // @[Modules.scala 71:109:@32901.4]
  wire [10:0] _T_78263; // @[Modules.scala 71:109:@32902.4]
  wire [10:0] buffer_13_694; // @[Modules.scala 71:109:@32903.4]
  wire [11:0] _T_78265; // @[Modules.scala 71:109:@32905.4]
  wire [10:0] _T_78266; // @[Modules.scala 71:109:@32906.4]
  wire [10:0] buffer_13_695; // @[Modules.scala 71:109:@32907.4]
  wire [11:0] _T_78268; // @[Modules.scala 71:109:@32909.4]
  wire [10:0] _T_78269; // @[Modules.scala 71:109:@32910.4]
  wire [10:0] buffer_13_696; // @[Modules.scala 71:109:@32911.4]
  wire [11:0] _T_78271; // @[Modules.scala 71:109:@32913.4]
  wire [10:0] _T_78272; // @[Modules.scala 71:109:@32914.4]
  wire [10:0] buffer_13_697; // @[Modules.scala 71:109:@32915.4]
  wire [11:0] _T_78274; // @[Modules.scala 71:109:@32917.4]
  wire [10:0] _T_78275; // @[Modules.scala 71:109:@32918.4]
  wire [10:0] buffer_13_698; // @[Modules.scala 71:109:@32919.4]
  wire [11:0] _T_78277; // @[Modules.scala 71:109:@32921.4]
  wire [10:0] _T_78278; // @[Modules.scala 71:109:@32922.4]
  wire [10:0] buffer_13_699; // @[Modules.scala 71:109:@32923.4]
  wire [11:0] _T_78280; // @[Modules.scala 71:109:@32925.4]
  wire [10:0] _T_78281; // @[Modules.scala 71:109:@32926.4]
  wire [10:0] buffer_13_700; // @[Modules.scala 71:109:@32927.4]
  wire [11:0] _T_78283; // @[Modules.scala 71:109:@32929.4]
  wire [10:0] _T_78284; // @[Modules.scala 71:109:@32930.4]
  wire [10:0] buffer_13_701; // @[Modules.scala 71:109:@32931.4]
  wire [11:0] _T_78286; // @[Modules.scala 71:109:@32933.4]
  wire [10:0] _T_78287; // @[Modules.scala 71:109:@32934.4]
  wire [10:0] buffer_13_702; // @[Modules.scala 71:109:@32935.4]
  wire [11:0] _T_78289; // @[Modules.scala 71:109:@32937.4]
  wire [10:0] _T_78290; // @[Modules.scala 71:109:@32938.4]
  wire [10:0] buffer_13_703; // @[Modules.scala 71:109:@32939.4]
  wire [11:0] _T_78292; // @[Modules.scala 71:109:@32941.4]
  wire [10:0] _T_78293; // @[Modules.scala 71:109:@32942.4]
  wire [10:0] buffer_13_704; // @[Modules.scala 71:109:@32943.4]
  wire [11:0] _T_78295; // @[Modules.scala 71:109:@32945.4]
  wire [10:0] _T_78296; // @[Modules.scala 71:109:@32946.4]
  wire [10:0] buffer_13_705; // @[Modules.scala 71:109:@32947.4]
  wire [11:0] _T_78298; // @[Modules.scala 71:109:@32949.4]
  wire [10:0] _T_78299; // @[Modules.scala 71:109:@32950.4]
  wire [10:0] buffer_13_706; // @[Modules.scala 71:109:@32951.4]
  wire [11:0] _T_78301; // @[Modules.scala 71:109:@32953.4]
  wire [10:0] _T_78302; // @[Modules.scala 71:109:@32954.4]
  wire [10:0] buffer_13_707; // @[Modules.scala 71:109:@32955.4]
  wire [11:0] _T_78304; // @[Modules.scala 71:109:@32957.4]
  wire [10:0] _T_78305; // @[Modules.scala 71:109:@32958.4]
  wire [10:0] buffer_13_708; // @[Modules.scala 71:109:@32959.4]
  wire [11:0] _T_78307; // @[Modules.scala 71:109:@32961.4]
  wire [10:0] _T_78308; // @[Modules.scala 71:109:@32962.4]
  wire [10:0] buffer_13_709; // @[Modules.scala 71:109:@32963.4]
  wire [11:0] _T_78310; // @[Modules.scala 71:109:@32965.4]
  wire [10:0] _T_78311; // @[Modules.scala 71:109:@32966.4]
  wire [10:0] buffer_13_710; // @[Modules.scala 71:109:@32967.4]
  wire [11:0] _T_78313; // @[Modules.scala 71:109:@32969.4]
  wire [10:0] _T_78314; // @[Modules.scala 71:109:@32970.4]
  wire [10:0] buffer_13_711; // @[Modules.scala 71:109:@32971.4]
  wire [11:0] _T_78316; // @[Modules.scala 71:109:@32973.4]
  wire [10:0] _T_78317; // @[Modules.scala 71:109:@32974.4]
  wire [10:0] buffer_13_712; // @[Modules.scala 71:109:@32975.4]
  wire [11:0] _T_78319; // @[Modules.scala 71:109:@32977.4]
  wire [10:0] _T_78320; // @[Modules.scala 71:109:@32978.4]
  wire [10:0] buffer_13_713; // @[Modules.scala 71:109:@32979.4]
  wire [11:0] _T_78322; // @[Modules.scala 71:109:@32981.4]
  wire [10:0] _T_78323; // @[Modules.scala 71:109:@32982.4]
  wire [10:0] buffer_13_714; // @[Modules.scala 71:109:@32983.4]
  wire [11:0] _T_78325; // @[Modules.scala 71:109:@32985.4]
  wire [10:0] _T_78326; // @[Modules.scala 71:109:@32986.4]
  wire [10:0] buffer_13_715; // @[Modules.scala 71:109:@32987.4]
  wire [11:0] _T_78328; // @[Modules.scala 71:109:@32989.4]
  wire [10:0] _T_78329; // @[Modules.scala 71:109:@32990.4]
  wire [10:0] buffer_13_716; // @[Modules.scala 71:109:@32991.4]
  wire [11:0] _T_78331; // @[Modules.scala 71:109:@32993.4]
  wire [10:0] _T_78332; // @[Modules.scala 71:109:@32994.4]
  wire [10:0] buffer_13_717; // @[Modules.scala 71:109:@32995.4]
  wire [11:0] _T_78334; // @[Modules.scala 71:109:@32997.4]
  wire [10:0] _T_78335; // @[Modules.scala 71:109:@32998.4]
  wire [10:0] buffer_13_718; // @[Modules.scala 71:109:@32999.4]
  wire [11:0] _T_78337; // @[Modules.scala 71:109:@33001.4]
  wire [10:0] _T_78338; // @[Modules.scala 71:109:@33002.4]
  wire [10:0] buffer_13_719; // @[Modules.scala 71:109:@33003.4]
  wire [11:0] _T_78340; // @[Modules.scala 71:109:@33005.4]
  wire [10:0] _T_78341; // @[Modules.scala 71:109:@33006.4]
  wire [10:0] buffer_13_720; // @[Modules.scala 71:109:@33007.4]
  wire [11:0] _T_78343; // @[Modules.scala 71:109:@33009.4]
  wire [10:0] _T_78344; // @[Modules.scala 71:109:@33010.4]
  wire [10:0] buffer_13_721; // @[Modules.scala 71:109:@33011.4]
  wire [11:0] _T_78346; // @[Modules.scala 71:109:@33013.4]
  wire [10:0] _T_78347; // @[Modules.scala 71:109:@33014.4]
  wire [10:0] buffer_13_722; // @[Modules.scala 71:109:@33015.4]
  wire [11:0] _T_78349; // @[Modules.scala 71:109:@33017.4]
  wire [10:0] _T_78350; // @[Modules.scala 71:109:@33018.4]
  wire [10:0] buffer_13_723; // @[Modules.scala 71:109:@33019.4]
  wire [11:0] _T_78352; // @[Modules.scala 71:109:@33021.4]
  wire [10:0] _T_78353; // @[Modules.scala 71:109:@33022.4]
  wire [10:0] buffer_13_724; // @[Modules.scala 71:109:@33023.4]
  wire [11:0] _T_78355; // @[Modules.scala 71:109:@33025.4]
  wire [10:0] _T_78356; // @[Modules.scala 71:109:@33026.4]
  wire [10:0] buffer_13_725; // @[Modules.scala 71:109:@33027.4]
  wire [11:0] _T_78358; // @[Modules.scala 71:109:@33029.4]
  wire [10:0] _T_78359; // @[Modules.scala 71:109:@33030.4]
  wire [10:0] buffer_13_726; // @[Modules.scala 71:109:@33031.4]
  wire [11:0] _T_78361; // @[Modules.scala 71:109:@33033.4]
  wire [10:0] _T_78362; // @[Modules.scala 71:109:@33034.4]
  wire [10:0] buffer_13_727; // @[Modules.scala 71:109:@33035.4]
  wire [11:0] _T_78364; // @[Modules.scala 71:109:@33037.4]
  wire [10:0] _T_78365; // @[Modules.scala 71:109:@33038.4]
  wire [10:0] buffer_13_728; // @[Modules.scala 71:109:@33039.4]
  wire [11:0] _T_78367; // @[Modules.scala 71:109:@33041.4]
  wire [10:0] _T_78368; // @[Modules.scala 71:109:@33042.4]
  wire [10:0] buffer_13_729; // @[Modules.scala 71:109:@33043.4]
  wire [11:0] _T_78373; // @[Modules.scala 71:109:@33049.4]
  wire [10:0] _T_78374; // @[Modules.scala 71:109:@33050.4]
  wire [10:0] buffer_13_731; // @[Modules.scala 71:109:@33051.4]
  wire [11:0] _T_78379; // @[Modules.scala 71:109:@33057.4]
  wire [10:0] _T_78380; // @[Modules.scala 71:109:@33058.4]
  wire [10:0] buffer_13_733; // @[Modules.scala 71:109:@33059.4]
  wire [11:0] _T_78382; // @[Modules.scala 71:109:@33061.4]
  wire [10:0] _T_78383; // @[Modules.scala 71:109:@33062.4]
  wire [10:0] buffer_13_734; // @[Modules.scala 71:109:@33063.4]
  wire [11:0] _T_78385; // @[Modules.scala 78:156:@33066.4]
  wire [10:0] _T_78386; // @[Modules.scala 78:156:@33067.4]
  wire [10:0] buffer_13_736; // @[Modules.scala 78:156:@33068.4]
  wire [11:0] _T_78388; // @[Modules.scala 78:156:@33070.4]
  wire [10:0] _T_78389; // @[Modules.scala 78:156:@33071.4]
  wire [10:0] buffer_13_737; // @[Modules.scala 78:156:@33072.4]
  wire [11:0] _T_78391; // @[Modules.scala 78:156:@33074.4]
  wire [10:0] _T_78392; // @[Modules.scala 78:156:@33075.4]
  wire [10:0] buffer_13_738; // @[Modules.scala 78:156:@33076.4]
  wire [11:0] _T_78394; // @[Modules.scala 78:156:@33078.4]
  wire [10:0] _T_78395; // @[Modules.scala 78:156:@33079.4]
  wire [10:0] buffer_13_739; // @[Modules.scala 78:156:@33080.4]
  wire [11:0] _T_78397; // @[Modules.scala 78:156:@33082.4]
  wire [10:0] _T_78398; // @[Modules.scala 78:156:@33083.4]
  wire [10:0] buffer_13_740; // @[Modules.scala 78:156:@33084.4]
  wire [11:0] _T_78400; // @[Modules.scala 78:156:@33086.4]
  wire [10:0] _T_78401; // @[Modules.scala 78:156:@33087.4]
  wire [10:0] buffer_13_741; // @[Modules.scala 78:156:@33088.4]
  wire [11:0] _T_78403; // @[Modules.scala 78:156:@33090.4]
  wire [10:0] _T_78404; // @[Modules.scala 78:156:@33091.4]
  wire [10:0] buffer_13_742; // @[Modules.scala 78:156:@33092.4]
  wire [11:0] _T_78406; // @[Modules.scala 78:156:@33094.4]
  wire [10:0] _T_78407; // @[Modules.scala 78:156:@33095.4]
  wire [10:0] buffer_13_743; // @[Modules.scala 78:156:@33096.4]
  wire [11:0] _T_78409; // @[Modules.scala 78:156:@33098.4]
  wire [10:0] _T_78410; // @[Modules.scala 78:156:@33099.4]
  wire [10:0] buffer_13_744; // @[Modules.scala 78:156:@33100.4]
  wire [11:0] _T_78412; // @[Modules.scala 78:156:@33102.4]
  wire [10:0] _T_78413; // @[Modules.scala 78:156:@33103.4]
  wire [10:0] buffer_13_745; // @[Modules.scala 78:156:@33104.4]
  wire [11:0] _T_78415; // @[Modules.scala 78:156:@33106.4]
  wire [10:0] _T_78416; // @[Modules.scala 78:156:@33107.4]
  wire [10:0] buffer_13_746; // @[Modules.scala 78:156:@33108.4]
  wire [11:0] _T_78418; // @[Modules.scala 78:156:@33110.4]
  wire [10:0] _T_78419; // @[Modules.scala 78:156:@33111.4]
  wire [10:0] buffer_13_747; // @[Modules.scala 78:156:@33112.4]
  wire [11:0] _T_78421; // @[Modules.scala 78:156:@33114.4]
  wire [10:0] _T_78422; // @[Modules.scala 78:156:@33115.4]
  wire [10:0] buffer_13_748; // @[Modules.scala 78:156:@33116.4]
  wire [11:0] _T_78424; // @[Modules.scala 78:156:@33118.4]
  wire [10:0] _T_78425; // @[Modules.scala 78:156:@33119.4]
  wire [10:0] buffer_13_749; // @[Modules.scala 78:156:@33120.4]
  wire [11:0] _T_78427; // @[Modules.scala 78:156:@33122.4]
  wire [10:0] _T_78428; // @[Modules.scala 78:156:@33123.4]
  wire [10:0] buffer_13_750; // @[Modules.scala 78:156:@33124.4]
  wire [11:0] _T_78430; // @[Modules.scala 78:156:@33126.4]
  wire [10:0] _T_78431; // @[Modules.scala 78:156:@33127.4]
  wire [10:0] buffer_13_751; // @[Modules.scala 78:156:@33128.4]
  wire [11:0] _T_78433; // @[Modules.scala 78:156:@33130.4]
  wire [10:0] _T_78434; // @[Modules.scala 78:156:@33131.4]
  wire [10:0] buffer_13_752; // @[Modules.scala 78:156:@33132.4]
  wire [11:0] _T_78436; // @[Modules.scala 78:156:@33134.4]
  wire [10:0] _T_78437; // @[Modules.scala 78:156:@33135.4]
  wire [10:0] buffer_13_753; // @[Modules.scala 78:156:@33136.4]
  wire [11:0] _T_78439; // @[Modules.scala 78:156:@33138.4]
  wire [10:0] _T_78440; // @[Modules.scala 78:156:@33139.4]
  wire [10:0] buffer_13_754; // @[Modules.scala 78:156:@33140.4]
  wire [11:0] _T_78442; // @[Modules.scala 78:156:@33142.4]
  wire [10:0] _T_78443; // @[Modules.scala 78:156:@33143.4]
  wire [10:0] buffer_13_755; // @[Modules.scala 78:156:@33144.4]
  wire [11:0] _T_78445; // @[Modules.scala 78:156:@33146.4]
  wire [10:0] _T_78446; // @[Modules.scala 78:156:@33147.4]
  wire [10:0] buffer_13_756; // @[Modules.scala 78:156:@33148.4]
  wire [11:0] _T_78448; // @[Modules.scala 78:156:@33150.4]
  wire [10:0] _T_78449; // @[Modules.scala 78:156:@33151.4]
  wire [10:0] buffer_13_757; // @[Modules.scala 78:156:@33152.4]
  wire [11:0] _T_78451; // @[Modules.scala 78:156:@33154.4]
  wire [10:0] _T_78452; // @[Modules.scala 78:156:@33155.4]
  wire [10:0] buffer_13_758; // @[Modules.scala 78:156:@33156.4]
  wire [11:0] _T_78454; // @[Modules.scala 78:156:@33158.4]
  wire [10:0] _T_78455; // @[Modules.scala 78:156:@33159.4]
  wire [10:0] buffer_13_759; // @[Modules.scala 78:156:@33160.4]
  wire [11:0] _T_78457; // @[Modules.scala 78:156:@33162.4]
  wire [10:0] _T_78458; // @[Modules.scala 78:156:@33163.4]
  wire [10:0] buffer_13_760; // @[Modules.scala 78:156:@33164.4]
  wire [11:0] _T_78460; // @[Modules.scala 78:156:@33166.4]
  wire [10:0] _T_78461; // @[Modules.scala 78:156:@33167.4]
  wire [10:0] buffer_13_761; // @[Modules.scala 78:156:@33168.4]
  wire [11:0] _T_78463; // @[Modules.scala 78:156:@33170.4]
  wire [10:0] _T_78464; // @[Modules.scala 78:156:@33171.4]
  wire [10:0] buffer_13_762; // @[Modules.scala 78:156:@33172.4]
  wire [11:0] _T_78466; // @[Modules.scala 78:156:@33174.4]
  wire [10:0] _T_78467; // @[Modules.scala 78:156:@33175.4]
  wire [10:0] buffer_13_763; // @[Modules.scala 78:156:@33176.4]
  wire [11:0] _T_78469; // @[Modules.scala 78:156:@33178.4]
  wire [10:0] _T_78470; // @[Modules.scala 78:156:@33179.4]
  wire [10:0] buffer_13_764; // @[Modules.scala 78:156:@33180.4]
  wire [11:0] _T_78472; // @[Modules.scala 78:156:@33182.4]
  wire [10:0] _T_78473; // @[Modules.scala 78:156:@33183.4]
  wire [10:0] buffer_13_765; // @[Modules.scala 78:156:@33184.4]
  wire [11:0] _T_78475; // @[Modules.scala 78:156:@33186.4]
  wire [10:0] _T_78476; // @[Modules.scala 78:156:@33187.4]
  wire [10:0] buffer_13_766; // @[Modules.scala 78:156:@33188.4]
  wire [11:0] _T_78478; // @[Modules.scala 78:156:@33190.4]
  wire [10:0] _T_78479; // @[Modules.scala 78:156:@33191.4]
  wire [10:0] buffer_13_767; // @[Modules.scala 78:156:@33192.4]
  wire [11:0] _T_78481; // @[Modules.scala 78:156:@33194.4]
  wire [10:0] _T_78482; // @[Modules.scala 78:156:@33195.4]
  wire [10:0] buffer_13_768; // @[Modules.scala 78:156:@33196.4]
  wire [11:0] _T_78484; // @[Modules.scala 78:156:@33198.4]
  wire [10:0] _T_78485; // @[Modules.scala 78:156:@33199.4]
  wire [10:0] buffer_13_769; // @[Modules.scala 78:156:@33200.4]
  wire [11:0] _T_78487; // @[Modules.scala 78:156:@33202.4]
  wire [10:0] _T_78488; // @[Modules.scala 78:156:@33203.4]
  wire [10:0] buffer_13_770; // @[Modules.scala 78:156:@33204.4]
  wire [11:0] _T_78490; // @[Modules.scala 78:156:@33206.4]
  wire [10:0] _T_78491; // @[Modules.scala 78:156:@33207.4]
  wire [10:0] buffer_13_771; // @[Modules.scala 78:156:@33208.4]
  wire [11:0] _T_78493; // @[Modules.scala 78:156:@33210.4]
  wire [10:0] _T_78494; // @[Modules.scala 78:156:@33211.4]
  wire [10:0] buffer_13_772; // @[Modules.scala 78:156:@33212.4]
  wire [11:0] _T_78496; // @[Modules.scala 78:156:@33214.4]
  wire [10:0] _T_78497; // @[Modules.scala 78:156:@33215.4]
  wire [10:0] buffer_13_773; // @[Modules.scala 78:156:@33216.4]
  wire [11:0] _T_78499; // @[Modules.scala 78:156:@33218.4]
  wire [10:0] _T_78500; // @[Modules.scala 78:156:@33219.4]
  wire [10:0] buffer_13_774; // @[Modules.scala 78:156:@33220.4]
  wire [11:0] _T_78502; // @[Modules.scala 78:156:@33222.4]
  wire [10:0] _T_78503; // @[Modules.scala 78:156:@33223.4]
  wire [10:0] buffer_13_775; // @[Modules.scala 78:156:@33224.4]
  wire [11:0] _T_78505; // @[Modules.scala 78:156:@33226.4]
  wire [10:0] _T_78506; // @[Modules.scala 78:156:@33227.4]
  wire [10:0] buffer_13_776; // @[Modules.scala 78:156:@33228.4]
  wire [11:0] _T_78508; // @[Modules.scala 78:156:@33230.4]
  wire [10:0] _T_78509; // @[Modules.scala 78:156:@33231.4]
  wire [10:0] buffer_13_777; // @[Modules.scala 78:156:@33232.4]
  wire [11:0] _T_78511; // @[Modules.scala 78:156:@33234.4]
  wire [10:0] _T_78512; // @[Modules.scala 78:156:@33235.4]
  wire [10:0] buffer_13_778; // @[Modules.scala 78:156:@33236.4]
  wire [11:0] _T_78514; // @[Modules.scala 78:156:@33238.4]
  wire [10:0] _T_78515; // @[Modules.scala 78:156:@33239.4]
  wire [10:0] buffer_13_779; // @[Modules.scala 78:156:@33240.4]
  wire [11:0] _T_78517; // @[Modules.scala 78:156:@33242.4]
  wire [10:0] _T_78518; // @[Modules.scala 78:156:@33243.4]
  wire [10:0] buffer_13_780; // @[Modules.scala 78:156:@33244.4]
  wire [11:0] _T_78520; // @[Modules.scala 78:156:@33246.4]
  wire [10:0] _T_78521; // @[Modules.scala 78:156:@33247.4]
  wire [10:0] buffer_13_781; // @[Modules.scala 78:156:@33248.4]
  wire [11:0] _T_78523; // @[Modules.scala 78:156:@33250.4]
  wire [10:0] _T_78524; // @[Modules.scala 78:156:@33251.4]
  wire [10:0] buffer_13_782; // @[Modules.scala 78:156:@33252.4]
  wire [11:0] _T_78526; // @[Modules.scala 78:156:@33254.4]
  wire [10:0] _T_78527; // @[Modules.scala 78:156:@33255.4]
  wire [10:0] buffer_13_783; // @[Modules.scala 78:156:@33256.4]
  wire [11:0] _T_79137; // @[Modules.scala 65:57:@34137.4]
  wire [10:0] _T_79138; // @[Modules.scala 65:57:@34138.4]
  wire [10:0] buffer_14_392; // @[Modules.scala 65:57:@34139.4]
  wire [11:0] _T_79143; // @[Modules.scala 65:57:@34145.4]
  wire [10:0] _T_79144; // @[Modules.scala 65:57:@34146.4]
  wire [10:0] buffer_14_394; // @[Modules.scala 65:57:@34147.4]
  wire [11:0] _T_79158; // @[Modules.scala 65:57:@34165.4]
  wire [10:0] _T_79159; // @[Modules.scala 65:57:@34166.4]
  wire [10:0] buffer_14_399; // @[Modules.scala 65:57:@34167.4]
  wire [11:0] _T_79167; // @[Modules.scala 65:57:@34177.4]
  wire [10:0] _T_79168; // @[Modules.scala 65:57:@34178.4]
  wire [10:0] buffer_14_402; // @[Modules.scala 65:57:@34179.4]
  wire [11:0] _T_79176; // @[Modules.scala 65:57:@34189.4]
  wire [10:0] _T_79177; // @[Modules.scala 65:57:@34190.4]
  wire [10:0] buffer_14_405; // @[Modules.scala 65:57:@34191.4]
  wire [10:0] buffer_14_30; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79182; // @[Modules.scala 65:57:@34197.4]
  wire [10:0] _T_79183; // @[Modules.scala 65:57:@34198.4]
  wire [10:0] buffer_14_407; // @[Modules.scala 65:57:@34199.4]
  wire [11:0] _T_79200; // @[Modules.scala 65:57:@34221.4]
  wire [10:0] _T_79201; // @[Modules.scala 65:57:@34222.4]
  wire [10:0] buffer_14_413; // @[Modules.scala 65:57:@34223.4]
  wire [10:0] buffer_14_45; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79203; // @[Modules.scala 65:57:@34225.4]
  wire [10:0] _T_79204; // @[Modules.scala 65:57:@34226.4]
  wire [10:0] buffer_14_414; // @[Modules.scala 65:57:@34227.4]
  wire [10:0] buffer_14_48; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79209; // @[Modules.scala 65:57:@34233.4]
  wire [10:0] _T_79210; // @[Modules.scala 65:57:@34234.4]
  wire [10:0] buffer_14_416; // @[Modules.scala 65:57:@34235.4]
  wire [11:0] _T_79221; // @[Modules.scala 65:57:@34249.4]
  wire [10:0] _T_79222; // @[Modules.scala 65:57:@34250.4]
  wire [10:0] buffer_14_420; // @[Modules.scala 65:57:@34251.4]
  wire [11:0] _T_79230; // @[Modules.scala 65:57:@34261.4]
  wire [10:0] _T_79231; // @[Modules.scala 65:57:@34262.4]
  wire [10:0] buffer_14_423; // @[Modules.scala 65:57:@34263.4]
  wire [11:0] _T_79242; // @[Modules.scala 65:57:@34277.4]
  wire [10:0] _T_79243; // @[Modules.scala 65:57:@34278.4]
  wire [10:0] buffer_14_427; // @[Modules.scala 65:57:@34279.4]
  wire [10:0] buffer_14_88; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79269; // @[Modules.scala 65:57:@34313.4]
  wire [10:0] _T_79270; // @[Modules.scala 65:57:@34314.4]
  wire [10:0] buffer_14_436; // @[Modules.scala 65:57:@34315.4]
  wire [11:0] _T_79275; // @[Modules.scala 65:57:@34321.4]
  wire [10:0] _T_79276; // @[Modules.scala 65:57:@34322.4]
  wire [10:0] buffer_14_438; // @[Modules.scala 65:57:@34323.4]
  wire [11:0] _T_79278; // @[Modules.scala 65:57:@34325.4]
  wire [10:0] _T_79279; // @[Modules.scala 65:57:@34326.4]
  wire [10:0] buffer_14_439; // @[Modules.scala 65:57:@34327.4]
  wire [11:0] _T_79317; // @[Modules.scala 65:57:@34377.4]
  wire [10:0] _T_79318; // @[Modules.scala 65:57:@34378.4]
  wire [10:0] buffer_14_452; // @[Modules.scala 65:57:@34379.4]
  wire [10:0] buffer_14_134; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79338; // @[Modules.scala 65:57:@34405.4]
  wire [10:0] _T_79339; // @[Modules.scala 65:57:@34406.4]
  wire [10:0] buffer_14_459; // @[Modules.scala 65:57:@34407.4]
  wire [11:0] _T_79341; // @[Modules.scala 65:57:@34409.4]
  wire [10:0] _T_79342; // @[Modules.scala 65:57:@34410.4]
  wire [10:0] buffer_14_460; // @[Modules.scala 65:57:@34411.4]
  wire [11:0] _T_79344; // @[Modules.scala 65:57:@34413.4]
  wire [10:0] _T_79345; // @[Modules.scala 65:57:@34414.4]
  wire [10:0] buffer_14_461; // @[Modules.scala 65:57:@34415.4]
  wire [10:0] buffer_14_164; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79383; // @[Modules.scala 65:57:@34465.4]
  wire [10:0] _T_79384; // @[Modules.scala 65:57:@34466.4]
  wire [10:0] buffer_14_474; // @[Modules.scala 65:57:@34467.4]
  wire [11:0] _T_79392; // @[Modules.scala 65:57:@34477.4]
  wire [10:0] _T_79393; // @[Modules.scala 65:57:@34478.4]
  wire [10:0] buffer_14_477; // @[Modules.scala 65:57:@34479.4]
  wire [10:0] buffer_14_173; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79395; // @[Modules.scala 65:57:@34481.4]
  wire [10:0] _T_79396; // @[Modules.scala 65:57:@34482.4]
  wire [10:0] buffer_14_478; // @[Modules.scala 65:57:@34483.4]
  wire [10:0] buffer_14_180; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79407; // @[Modules.scala 65:57:@34497.4]
  wire [10:0] _T_79408; // @[Modules.scala 65:57:@34498.4]
  wire [10:0] buffer_14_482; // @[Modules.scala 65:57:@34499.4]
  wire [11:0] _T_79413; // @[Modules.scala 65:57:@34505.4]
  wire [10:0] _T_79414; // @[Modules.scala 65:57:@34506.4]
  wire [10:0] buffer_14_484; // @[Modules.scala 65:57:@34507.4]
  wire [11:0] _T_79416; // @[Modules.scala 65:57:@34509.4]
  wire [10:0] _T_79417; // @[Modules.scala 65:57:@34510.4]
  wire [10:0] buffer_14_485; // @[Modules.scala 65:57:@34511.4]
  wire [11:0] _T_79425; // @[Modules.scala 65:57:@34521.4]
  wire [10:0] _T_79426; // @[Modules.scala 65:57:@34522.4]
  wire [10:0] buffer_14_488; // @[Modules.scala 65:57:@34523.4]
  wire [11:0] _T_79449; // @[Modules.scala 65:57:@34553.4]
  wire [10:0] _T_79450; // @[Modules.scala 65:57:@34554.4]
  wire [10:0] buffer_14_496; // @[Modules.scala 65:57:@34555.4]
  wire [10:0] buffer_14_215; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79458; // @[Modules.scala 65:57:@34565.4]
  wire [10:0] _T_79459; // @[Modules.scala 65:57:@34566.4]
  wire [10:0] buffer_14_499; // @[Modules.scala 65:57:@34567.4]
  wire [10:0] buffer_14_216; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79461; // @[Modules.scala 65:57:@34569.4]
  wire [10:0] _T_79462; // @[Modules.scala 65:57:@34570.4]
  wire [10:0] buffer_14_500; // @[Modules.scala 65:57:@34571.4]
  wire [11:0] _T_79464; // @[Modules.scala 65:57:@34573.4]
  wire [10:0] _T_79465; // @[Modules.scala 65:57:@34574.4]
  wire [10:0] buffer_14_501; // @[Modules.scala 65:57:@34575.4]
  wire [11:0] _T_79485; // @[Modules.scala 65:57:@34601.4]
  wire [10:0] _T_79486; // @[Modules.scala 65:57:@34602.4]
  wire [10:0] buffer_14_508; // @[Modules.scala 65:57:@34603.4]
  wire [11:0] _T_79488; // @[Modules.scala 65:57:@34605.4]
  wire [10:0] _T_79489; // @[Modules.scala 65:57:@34606.4]
  wire [10:0] buffer_14_509; // @[Modules.scala 65:57:@34607.4]
  wire [11:0] _T_79491; // @[Modules.scala 65:57:@34609.4]
  wire [10:0] _T_79492; // @[Modules.scala 65:57:@34610.4]
  wire [10:0] buffer_14_510; // @[Modules.scala 65:57:@34611.4]
  wire [11:0] _T_79494; // @[Modules.scala 65:57:@34613.4]
  wire [10:0] _T_79495; // @[Modules.scala 65:57:@34614.4]
  wire [10:0] buffer_14_511; // @[Modules.scala 65:57:@34615.4]
  wire [11:0] _T_79503; // @[Modules.scala 65:57:@34625.4]
  wire [10:0] _T_79504; // @[Modules.scala 65:57:@34626.4]
  wire [10:0] buffer_14_514; // @[Modules.scala 65:57:@34627.4]
  wire [11:0] _T_79509; // @[Modules.scala 65:57:@34633.4]
  wire [10:0] _T_79510; // @[Modules.scala 65:57:@34634.4]
  wire [10:0] buffer_14_516; // @[Modules.scala 65:57:@34635.4]
  wire [11:0] _T_79515; // @[Modules.scala 65:57:@34641.4]
  wire [10:0] _T_79516; // @[Modules.scala 65:57:@34642.4]
  wire [10:0] buffer_14_518; // @[Modules.scala 65:57:@34643.4]
  wire [11:0] _T_79524; // @[Modules.scala 65:57:@34653.4]
  wire [10:0] _T_79525; // @[Modules.scala 65:57:@34654.4]
  wire [10:0] buffer_14_521; // @[Modules.scala 65:57:@34655.4]
  wire [11:0] _T_79536; // @[Modules.scala 65:57:@34669.4]
  wire [10:0] _T_79537; // @[Modules.scala 65:57:@34670.4]
  wire [10:0] buffer_14_525; // @[Modules.scala 65:57:@34671.4]
  wire [11:0] _T_79542; // @[Modules.scala 65:57:@34677.4]
  wire [10:0] _T_79543; // @[Modules.scala 65:57:@34678.4]
  wire [10:0] buffer_14_527; // @[Modules.scala 65:57:@34679.4]
  wire [11:0] _T_79557; // @[Modules.scala 65:57:@34697.4]
  wire [10:0] _T_79558; // @[Modules.scala 65:57:@34698.4]
  wire [10:0] buffer_14_532; // @[Modules.scala 65:57:@34699.4]
  wire [10:0] buffer_14_284; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79563; // @[Modules.scala 65:57:@34705.4]
  wire [10:0] _T_79564; // @[Modules.scala 65:57:@34706.4]
  wire [10:0] buffer_14_534; // @[Modules.scala 65:57:@34707.4]
  wire [11:0] _T_79569; // @[Modules.scala 65:57:@34713.4]
  wire [10:0] _T_79570; // @[Modules.scala 65:57:@34714.4]
  wire [10:0] buffer_14_536; // @[Modules.scala 65:57:@34715.4]
  wire [11:0] _T_79578; // @[Modules.scala 65:57:@34725.4]
  wire [10:0] _T_79579; // @[Modules.scala 65:57:@34726.4]
  wire [10:0] buffer_14_539; // @[Modules.scala 65:57:@34727.4]
  wire [11:0] _T_79590; // @[Modules.scala 65:57:@34741.4]
  wire [10:0] _T_79591; // @[Modules.scala 65:57:@34742.4]
  wire [10:0] buffer_14_543; // @[Modules.scala 65:57:@34743.4]
  wire [11:0] _T_79599; // @[Modules.scala 65:57:@34753.4]
  wire [10:0] _T_79600; // @[Modules.scala 65:57:@34754.4]
  wire [10:0] buffer_14_546; // @[Modules.scala 65:57:@34755.4]
  wire [11:0] _T_79602; // @[Modules.scala 65:57:@34757.4]
  wire [10:0] _T_79603; // @[Modules.scala 65:57:@34758.4]
  wire [10:0] buffer_14_547; // @[Modules.scala 65:57:@34759.4]
  wire [11:0] _T_79617; // @[Modules.scala 65:57:@34777.4]
  wire [10:0] _T_79618; // @[Modules.scala 65:57:@34778.4]
  wire [10:0] buffer_14_552; // @[Modules.scala 65:57:@34779.4]
  wire [11:0] _T_79626; // @[Modules.scala 65:57:@34789.4]
  wire [10:0] _T_79627; // @[Modules.scala 65:57:@34790.4]
  wire [10:0] buffer_14_555; // @[Modules.scala 65:57:@34791.4]
  wire [11:0] _T_79659; // @[Modules.scala 65:57:@34833.4]
  wire [10:0] _T_79660; // @[Modules.scala 65:57:@34834.4]
  wire [10:0] buffer_14_566; // @[Modules.scala 65:57:@34835.4]
  wire [11:0] _T_79665; // @[Modules.scala 65:57:@34841.4]
  wire [10:0] _T_79666; // @[Modules.scala 65:57:@34842.4]
  wire [10:0] buffer_14_568; // @[Modules.scala 65:57:@34843.4]
  wire [10:0] buffer_14_354; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79668; // @[Modules.scala 65:57:@34845.4]
  wire [10:0] _T_79669; // @[Modules.scala 65:57:@34846.4]
  wire [10:0] buffer_14_569; // @[Modules.scala 65:57:@34847.4]
  wire [11:0] _T_79671; // @[Modules.scala 65:57:@34849.4]
  wire [10:0] _T_79672; // @[Modules.scala 65:57:@34850.4]
  wire [10:0] buffer_14_570; // @[Modules.scala 65:57:@34851.4]
  wire [10:0] buffer_14_363; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79680; // @[Modules.scala 65:57:@34861.4]
  wire [10:0] _T_79681; // @[Modules.scala 65:57:@34862.4]
  wire [10:0] buffer_14_573; // @[Modules.scala 65:57:@34863.4]
  wire [11:0] _T_79683; // @[Modules.scala 65:57:@34865.4]
  wire [10:0] _T_79684; // @[Modules.scala 65:57:@34866.4]
  wire [10:0] buffer_14_574; // @[Modules.scala 65:57:@34867.4]
  wire [10:0] buffer_14_367; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79686; // @[Modules.scala 65:57:@34869.4]
  wire [10:0] _T_79687; // @[Modules.scala 65:57:@34870.4]
  wire [10:0] buffer_14_575; // @[Modules.scala 65:57:@34871.4]
  wire [10:0] buffer_14_368; // @[Modules.scala 32:22:@8.4]
  wire [10:0] buffer_14_369; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_79689; // @[Modules.scala 65:57:@34873.4]
  wire [10:0] _T_79690; // @[Modules.scala 65:57:@34874.4]
  wire [10:0] buffer_14_576; // @[Modules.scala 65:57:@34875.4]
  wire [11:0] _T_79692; // @[Modules.scala 65:57:@34877.4]
  wire [10:0] _T_79693; // @[Modules.scala 65:57:@34878.4]
  wire [10:0] buffer_14_577; // @[Modules.scala 65:57:@34879.4]
  wire [11:0] _T_79722; // @[Modules.scala 65:57:@34917.4]
  wire [10:0] _T_79723; // @[Modules.scala 65:57:@34918.4]
  wire [10:0] buffer_14_587; // @[Modules.scala 65:57:@34919.4]
  wire [11:0] _T_79725; // @[Modules.scala 68:83:@34921.4]
  wire [10:0] _T_79726; // @[Modules.scala 68:83:@34922.4]
  wire [10:0] buffer_14_588; // @[Modules.scala 68:83:@34923.4]
  wire [11:0] _T_79728; // @[Modules.scala 68:83:@34925.4]
  wire [10:0] _T_79729; // @[Modules.scala 68:83:@34926.4]
  wire [10:0] buffer_14_589; // @[Modules.scala 68:83:@34927.4]
  wire [11:0] _T_79731; // @[Modules.scala 68:83:@34929.4]
  wire [10:0] _T_79732; // @[Modules.scala 68:83:@34930.4]
  wire [10:0] buffer_14_590; // @[Modules.scala 68:83:@34931.4]
  wire [11:0] _T_79734; // @[Modules.scala 68:83:@34933.4]
  wire [10:0] _T_79735; // @[Modules.scala 68:83:@34934.4]
  wire [10:0] buffer_14_591; // @[Modules.scala 68:83:@34935.4]
  wire [11:0] _T_79737; // @[Modules.scala 68:83:@34937.4]
  wire [10:0] _T_79738; // @[Modules.scala 68:83:@34938.4]
  wire [10:0] buffer_14_592; // @[Modules.scala 68:83:@34939.4]
  wire [11:0] _T_79740; // @[Modules.scala 68:83:@34941.4]
  wire [10:0] _T_79741; // @[Modules.scala 68:83:@34942.4]
  wire [10:0] buffer_14_593; // @[Modules.scala 68:83:@34943.4]
  wire [11:0] _T_79743; // @[Modules.scala 68:83:@34945.4]
  wire [10:0] _T_79744; // @[Modules.scala 68:83:@34946.4]
  wire [10:0] buffer_14_594; // @[Modules.scala 68:83:@34947.4]
  wire [11:0] _T_79746; // @[Modules.scala 68:83:@34949.4]
  wire [10:0] _T_79747; // @[Modules.scala 68:83:@34950.4]
  wire [10:0] buffer_14_595; // @[Modules.scala 68:83:@34951.4]
  wire [11:0] _T_79755; // @[Modules.scala 68:83:@34961.4]
  wire [10:0] _T_79756; // @[Modules.scala 68:83:@34962.4]
  wire [10:0] buffer_14_598; // @[Modules.scala 68:83:@34963.4]
  wire [11:0] _T_79758; // @[Modules.scala 68:83:@34965.4]
  wire [10:0] _T_79759; // @[Modules.scala 68:83:@34966.4]
  wire [10:0] buffer_14_599; // @[Modules.scala 68:83:@34967.4]
  wire [11:0] _T_79761; // @[Modules.scala 68:83:@34969.4]
  wire [10:0] _T_79762; // @[Modules.scala 68:83:@34970.4]
  wire [10:0] buffer_14_600; // @[Modules.scala 68:83:@34971.4]
  wire [11:0] _T_79764; // @[Modules.scala 68:83:@34973.4]
  wire [10:0] _T_79765; // @[Modules.scala 68:83:@34974.4]
  wire [10:0] buffer_14_601; // @[Modules.scala 68:83:@34975.4]
  wire [11:0] _T_79767; // @[Modules.scala 68:83:@34977.4]
  wire [10:0] _T_79768; // @[Modules.scala 68:83:@34978.4]
  wire [10:0] buffer_14_602; // @[Modules.scala 68:83:@34979.4]
  wire [11:0] _T_79770; // @[Modules.scala 68:83:@34981.4]
  wire [10:0] _T_79771; // @[Modules.scala 68:83:@34982.4]
  wire [10:0] buffer_14_603; // @[Modules.scala 68:83:@34983.4]
  wire [11:0] _T_79773; // @[Modules.scala 68:83:@34985.4]
  wire [10:0] _T_79774; // @[Modules.scala 68:83:@34986.4]
  wire [10:0] buffer_14_604; // @[Modules.scala 68:83:@34987.4]
  wire [11:0] _T_79776; // @[Modules.scala 68:83:@34989.4]
  wire [10:0] _T_79777; // @[Modules.scala 68:83:@34990.4]
  wire [10:0] buffer_14_605; // @[Modules.scala 68:83:@34991.4]
  wire [11:0] _T_79779; // @[Modules.scala 68:83:@34993.4]
  wire [10:0] _T_79780; // @[Modules.scala 68:83:@34994.4]
  wire [10:0] buffer_14_606; // @[Modules.scala 68:83:@34995.4]
  wire [11:0] _T_79785; // @[Modules.scala 68:83:@35001.4]
  wire [10:0] _T_79786; // @[Modules.scala 68:83:@35002.4]
  wire [10:0] buffer_14_608; // @[Modules.scala 68:83:@35003.4]
  wire [11:0] _T_79788; // @[Modules.scala 68:83:@35005.4]
  wire [10:0] _T_79789; // @[Modules.scala 68:83:@35006.4]
  wire [10:0] buffer_14_609; // @[Modules.scala 68:83:@35007.4]
  wire [11:0] _T_79791; // @[Modules.scala 68:83:@35009.4]
  wire [10:0] _T_79792; // @[Modules.scala 68:83:@35010.4]
  wire [10:0] buffer_14_610; // @[Modules.scala 68:83:@35011.4]
  wire [11:0] _T_79794; // @[Modules.scala 68:83:@35013.4]
  wire [10:0] _T_79795; // @[Modules.scala 68:83:@35014.4]
  wire [10:0] buffer_14_611; // @[Modules.scala 68:83:@35015.4]
  wire [11:0] _T_79800; // @[Modules.scala 68:83:@35021.4]
  wire [10:0] _T_79801; // @[Modules.scala 68:83:@35022.4]
  wire [10:0] buffer_14_613; // @[Modules.scala 68:83:@35023.4]
  wire [11:0] _T_79803; // @[Modules.scala 68:83:@35025.4]
  wire [10:0] _T_79804; // @[Modules.scala 68:83:@35026.4]
  wire [10:0] buffer_14_614; // @[Modules.scala 68:83:@35027.4]
  wire [11:0] _T_79806; // @[Modules.scala 68:83:@35029.4]
  wire [10:0] _T_79807; // @[Modules.scala 68:83:@35030.4]
  wire [10:0] buffer_14_615; // @[Modules.scala 68:83:@35031.4]
  wire [11:0] _T_79812; // @[Modules.scala 68:83:@35037.4]
  wire [10:0] _T_79813; // @[Modules.scala 68:83:@35038.4]
  wire [10:0] buffer_14_617; // @[Modules.scala 68:83:@35039.4]
  wire [11:0] _T_79815; // @[Modules.scala 68:83:@35041.4]
  wire [10:0] _T_79816; // @[Modules.scala 68:83:@35042.4]
  wire [10:0] buffer_14_618; // @[Modules.scala 68:83:@35043.4]
  wire [11:0] _T_79824; // @[Modules.scala 68:83:@35053.4]
  wire [10:0] _T_79825; // @[Modules.scala 68:83:@35054.4]
  wire [10:0] buffer_14_621; // @[Modules.scala 68:83:@35055.4]
  wire [11:0] _T_79827; // @[Modules.scala 68:83:@35057.4]
  wire [10:0] _T_79828; // @[Modules.scala 68:83:@35058.4]
  wire [10:0] buffer_14_622; // @[Modules.scala 68:83:@35059.4]
  wire [11:0] _T_79833; // @[Modules.scala 68:83:@35065.4]
  wire [10:0] _T_79834; // @[Modules.scala 68:83:@35066.4]
  wire [10:0] buffer_14_624; // @[Modules.scala 68:83:@35067.4]
  wire [11:0] _T_79836; // @[Modules.scala 68:83:@35069.4]
  wire [10:0] _T_79837; // @[Modules.scala 68:83:@35070.4]
  wire [10:0] buffer_14_625; // @[Modules.scala 68:83:@35071.4]
  wire [11:0] _T_79845; // @[Modules.scala 68:83:@35081.4]
  wire [10:0] _T_79846; // @[Modules.scala 68:83:@35082.4]
  wire [10:0] buffer_14_628; // @[Modules.scala 68:83:@35083.4]
  wire [11:0] _T_79848; // @[Modules.scala 68:83:@35085.4]
  wire [10:0] _T_79849; // @[Modules.scala 68:83:@35086.4]
  wire [10:0] buffer_14_629; // @[Modules.scala 68:83:@35087.4]
  wire [11:0] _T_79851; // @[Modules.scala 68:83:@35089.4]
  wire [10:0] _T_79852; // @[Modules.scala 68:83:@35090.4]
  wire [10:0] buffer_14_630; // @[Modules.scala 68:83:@35091.4]
  wire [11:0] _T_79854; // @[Modules.scala 68:83:@35093.4]
  wire [10:0] _T_79855; // @[Modules.scala 68:83:@35094.4]
  wire [10:0] buffer_14_631; // @[Modules.scala 68:83:@35095.4]
  wire [11:0] _T_79860; // @[Modules.scala 68:83:@35101.4]
  wire [10:0] _T_79861; // @[Modules.scala 68:83:@35102.4]
  wire [10:0] buffer_14_633; // @[Modules.scala 68:83:@35103.4]
  wire [11:0] _T_79863; // @[Modules.scala 68:83:@35105.4]
  wire [10:0] _T_79864; // @[Modules.scala 68:83:@35106.4]
  wire [10:0] buffer_14_634; // @[Modules.scala 68:83:@35107.4]
  wire [11:0] _T_79866; // @[Modules.scala 68:83:@35109.4]
  wire [10:0] _T_79867; // @[Modules.scala 68:83:@35110.4]
  wire [10:0] buffer_14_635; // @[Modules.scala 68:83:@35111.4]
  wire [11:0] _T_79869; // @[Modules.scala 68:83:@35113.4]
  wire [10:0] _T_79870; // @[Modules.scala 68:83:@35114.4]
  wire [10:0] buffer_14_636; // @[Modules.scala 68:83:@35115.4]
  wire [11:0] _T_79875; // @[Modules.scala 68:83:@35121.4]
  wire [10:0] _T_79876; // @[Modules.scala 68:83:@35122.4]
  wire [10:0] buffer_14_638; // @[Modules.scala 68:83:@35123.4]
  wire [11:0] _T_79878; // @[Modules.scala 68:83:@35125.4]
  wire [10:0] _T_79879; // @[Modules.scala 68:83:@35126.4]
  wire [10:0] buffer_14_639; // @[Modules.scala 68:83:@35127.4]
  wire [11:0] _T_79881; // @[Modules.scala 68:83:@35129.4]
  wire [10:0] _T_79882; // @[Modules.scala 68:83:@35130.4]
  wire [10:0] buffer_14_640; // @[Modules.scala 68:83:@35131.4]
  wire [11:0] _T_79884; // @[Modules.scala 68:83:@35133.4]
  wire [10:0] _T_79885; // @[Modules.scala 68:83:@35134.4]
  wire [10:0] buffer_14_641; // @[Modules.scala 68:83:@35135.4]
  wire [11:0] _T_79887; // @[Modules.scala 68:83:@35137.4]
  wire [10:0] _T_79888; // @[Modules.scala 68:83:@35138.4]
  wire [10:0] buffer_14_642; // @[Modules.scala 68:83:@35139.4]
  wire [11:0] _T_79890; // @[Modules.scala 68:83:@35141.4]
  wire [10:0] _T_79891; // @[Modules.scala 68:83:@35142.4]
  wire [10:0] buffer_14_643; // @[Modules.scala 68:83:@35143.4]
  wire [11:0] _T_79893; // @[Modules.scala 68:83:@35145.4]
  wire [10:0] _T_79894; // @[Modules.scala 68:83:@35146.4]
  wire [10:0] buffer_14_644; // @[Modules.scala 68:83:@35147.4]
  wire [11:0] _T_79899; // @[Modules.scala 68:83:@35153.4]
  wire [10:0] _T_79900; // @[Modules.scala 68:83:@35154.4]
  wire [10:0] buffer_14_646; // @[Modules.scala 68:83:@35155.4]
  wire [11:0] _T_79902; // @[Modules.scala 68:83:@35157.4]
  wire [10:0] _T_79903; // @[Modules.scala 68:83:@35158.4]
  wire [10:0] buffer_14_647; // @[Modules.scala 68:83:@35159.4]
  wire [11:0] _T_79908; // @[Modules.scala 68:83:@35165.4]
  wire [10:0] _T_79909; // @[Modules.scala 68:83:@35166.4]
  wire [10:0] buffer_14_649; // @[Modules.scala 68:83:@35167.4]
  wire [11:0] _T_79911; // @[Modules.scala 68:83:@35169.4]
  wire [10:0] _T_79912; // @[Modules.scala 68:83:@35170.4]
  wire [10:0] buffer_14_650; // @[Modules.scala 68:83:@35171.4]
  wire [11:0] _T_79914; // @[Modules.scala 68:83:@35173.4]
  wire [10:0] _T_79915; // @[Modules.scala 68:83:@35174.4]
  wire [10:0] buffer_14_651; // @[Modules.scala 68:83:@35175.4]
  wire [11:0] _T_79917; // @[Modules.scala 68:83:@35177.4]
  wire [10:0] _T_79918; // @[Modules.scala 68:83:@35178.4]
  wire [10:0] buffer_14_652; // @[Modules.scala 68:83:@35179.4]
  wire [11:0] _T_79920; // @[Modules.scala 68:83:@35181.4]
  wire [10:0] _T_79921; // @[Modules.scala 68:83:@35182.4]
  wire [10:0] buffer_14_653; // @[Modules.scala 68:83:@35183.4]
  wire [11:0] _T_79923; // @[Modules.scala 68:83:@35185.4]
  wire [10:0] _T_79924; // @[Modules.scala 68:83:@35186.4]
  wire [10:0] buffer_14_654; // @[Modules.scala 68:83:@35187.4]
  wire [11:0] _T_79926; // @[Modules.scala 68:83:@35189.4]
  wire [10:0] _T_79927; // @[Modules.scala 68:83:@35190.4]
  wire [10:0] buffer_14_655; // @[Modules.scala 68:83:@35191.4]
  wire [11:0] _T_79929; // @[Modules.scala 68:83:@35193.4]
  wire [10:0] _T_79930; // @[Modules.scala 68:83:@35194.4]
  wire [10:0] buffer_14_656; // @[Modules.scala 68:83:@35195.4]
  wire [11:0] _T_79935; // @[Modules.scala 68:83:@35201.4]
  wire [10:0] _T_79936; // @[Modules.scala 68:83:@35202.4]
  wire [10:0] buffer_14_658; // @[Modules.scala 68:83:@35203.4]
  wire [11:0] _T_79938; // @[Modules.scala 68:83:@35205.4]
  wire [10:0] _T_79939; // @[Modules.scala 68:83:@35206.4]
  wire [10:0] buffer_14_659; // @[Modules.scala 68:83:@35207.4]
  wire [11:0] _T_79941; // @[Modules.scala 68:83:@35209.4]
  wire [10:0] _T_79942; // @[Modules.scala 68:83:@35210.4]
  wire [10:0] buffer_14_660; // @[Modules.scala 68:83:@35211.4]
  wire [11:0] _T_79944; // @[Modules.scala 68:83:@35213.4]
  wire [10:0] _T_79945; // @[Modules.scala 68:83:@35214.4]
  wire [10:0] buffer_14_661; // @[Modules.scala 68:83:@35215.4]
  wire [11:0] _T_79947; // @[Modules.scala 68:83:@35217.4]
  wire [10:0] _T_79948; // @[Modules.scala 68:83:@35218.4]
  wire [10:0] buffer_14_662; // @[Modules.scala 68:83:@35219.4]
  wire [11:0] _T_79950; // @[Modules.scala 68:83:@35221.4]
  wire [10:0] _T_79951; // @[Modules.scala 68:83:@35222.4]
  wire [10:0] buffer_14_663; // @[Modules.scala 68:83:@35223.4]
  wire [11:0] _T_79956; // @[Modules.scala 68:83:@35229.4]
  wire [10:0] _T_79957; // @[Modules.scala 68:83:@35230.4]
  wire [10:0] buffer_14_665; // @[Modules.scala 68:83:@35231.4]
  wire [11:0] _T_79965; // @[Modules.scala 68:83:@35241.4]
  wire [10:0] _T_79966; // @[Modules.scala 68:83:@35242.4]
  wire [10:0] buffer_14_668; // @[Modules.scala 68:83:@35243.4]
  wire [11:0] _T_79968; // @[Modules.scala 68:83:@35245.4]
  wire [10:0] _T_79969; // @[Modules.scala 68:83:@35246.4]
  wire [10:0] buffer_14_669; // @[Modules.scala 68:83:@35247.4]
  wire [11:0] _T_79977; // @[Modules.scala 68:83:@35257.4]
  wire [10:0] _T_79978; // @[Modules.scala 68:83:@35258.4]
  wire [10:0] buffer_14_672; // @[Modules.scala 68:83:@35259.4]
  wire [11:0] _T_79980; // @[Modules.scala 68:83:@35261.4]
  wire [10:0] _T_79981; // @[Modules.scala 68:83:@35262.4]
  wire [10:0] buffer_14_673; // @[Modules.scala 68:83:@35263.4]
  wire [11:0] _T_79986; // @[Modules.scala 68:83:@35269.4]
  wire [10:0] _T_79987; // @[Modules.scala 68:83:@35270.4]
  wire [10:0] buffer_14_675; // @[Modules.scala 68:83:@35271.4]
  wire [11:0] _T_79989; // @[Modules.scala 68:83:@35273.4]
  wire [10:0] _T_79990; // @[Modules.scala 68:83:@35274.4]
  wire [10:0] buffer_14_676; // @[Modules.scala 68:83:@35275.4]
  wire [11:0] _T_79992; // @[Modules.scala 68:83:@35277.4]
  wire [10:0] _T_79993; // @[Modules.scala 68:83:@35278.4]
  wire [10:0] buffer_14_677; // @[Modules.scala 68:83:@35279.4]
  wire [11:0] _T_79995; // @[Modules.scala 68:83:@35281.4]
  wire [10:0] _T_79996; // @[Modules.scala 68:83:@35282.4]
  wire [10:0] buffer_14_678; // @[Modules.scala 68:83:@35283.4]
  wire [11:0] _T_79998; // @[Modules.scala 68:83:@35285.4]
  wire [10:0] _T_79999; // @[Modules.scala 68:83:@35286.4]
  wire [10:0] buffer_14_679; // @[Modules.scala 68:83:@35287.4]
  wire [11:0] _T_80001; // @[Modules.scala 68:83:@35289.4]
  wire [10:0] _T_80002; // @[Modules.scala 68:83:@35290.4]
  wire [10:0] buffer_14_680; // @[Modules.scala 68:83:@35291.4]
  wire [11:0] _T_80004; // @[Modules.scala 68:83:@35293.4]
  wire [10:0] _T_80005; // @[Modules.scala 68:83:@35294.4]
  wire [10:0] buffer_14_681; // @[Modules.scala 68:83:@35295.4]
  wire [11:0] _T_80007; // @[Modules.scala 68:83:@35297.4]
  wire [10:0] _T_80008; // @[Modules.scala 68:83:@35298.4]
  wire [10:0] buffer_14_682; // @[Modules.scala 68:83:@35299.4]
  wire [11:0] _T_80010; // @[Modules.scala 68:83:@35301.4]
  wire [10:0] _T_80011; // @[Modules.scala 68:83:@35302.4]
  wire [10:0] buffer_14_683; // @[Modules.scala 68:83:@35303.4]
  wire [11:0] _T_80016; // @[Modules.scala 68:83:@35309.4]
  wire [10:0] _T_80017; // @[Modules.scala 68:83:@35310.4]
  wire [10:0] buffer_14_685; // @[Modules.scala 68:83:@35311.4]
  wire [11:0] _T_80019; // @[Modules.scala 71:109:@35313.4]
  wire [10:0] _T_80020; // @[Modules.scala 71:109:@35314.4]
  wire [10:0] buffer_14_686; // @[Modules.scala 71:109:@35315.4]
  wire [11:0] _T_80022; // @[Modules.scala 71:109:@35317.4]
  wire [10:0] _T_80023; // @[Modules.scala 71:109:@35318.4]
  wire [10:0] buffer_14_687; // @[Modules.scala 71:109:@35319.4]
  wire [11:0] _T_80025; // @[Modules.scala 71:109:@35321.4]
  wire [10:0] _T_80026; // @[Modules.scala 71:109:@35322.4]
  wire [10:0] buffer_14_688; // @[Modules.scala 71:109:@35323.4]
  wire [11:0] _T_80028; // @[Modules.scala 71:109:@35325.4]
  wire [10:0] _T_80029; // @[Modules.scala 71:109:@35326.4]
  wire [10:0] buffer_14_689; // @[Modules.scala 71:109:@35327.4]
  wire [11:0] _T_80034; // @[Modules.scala 71:109:@35333.4]
  wire [10:0] _T_80035; // @[Modules.scala 71:109:@35334.4]
  wire [10:0] buffer_14_691; // @[Modules.scala 71:109:@35335.4]
  wire [11:0] _T_80037; // @[Modules.scala 71:109:@35337.4]
  wire [10:0] _T_80038; // @[Modules.scala 71:109:@35338.4]
  wire [10:0] buffer_14_692; // @[Modules.scala 71:109:@35339.4]
  wire [11:0] _T_80040; // @[Modules.scala 71:109:@35341.4]
  wire [10:0] _T_80041; // @[Modules.scala 71:109:@35342.4]
  wire [10:0] buffer_14_693; // @[Modules.scala 71:109:@35343.4]
  wire [11:0] _T_80043; // @[Modules.scala 71:109:@35345.4]
  wire [10:0] _T_80044; // @[Modules.scala 71:109:@35346.4]
  wire [10:0] buffer_14_694; // @[Modules.scala 71:109:@35347.4]
  wire [11:0] _T_80046; // @[Modules.scala 71:109:@35349.4]
  wire [10:0] _T_80047; // @[Modules.scala 71:109:@35350.4]
  wire [10:0] buffer_14_695; // @[Modules.scala 71:109:@35351.4]
  wire [11:0] _T_80049; // @[Modules.scala 71:109:@35353.4]
  wire [10:0] _T_80050; // @[Modules.scala 71:109:@35354.4]
  wire [10:0] buffer_14_696; // @[Modules.scala 71:109:@35355.4]
  wire [11:0] _T_80052; // @[Modules.scala 71:109:@35357.4]
  wire [10:0] _T_80053; // @[Modules.scala 71:109:@35358.4]
  wire [10:0] buffer_14_697; // @[Modules.scala 71:109:@35359.4]
  wire [11:0] _T_80055; // @[Modules.scala 71:109:@35361.4]
  wire [10:0] _T_80056; // @[Modules.scala 71:109:@35362.4]
  wire [10:0] buffer_14_698; // @[Modules.scala 71:109:@35363.4]
  wire [11:0] _T_80058; // @[Modules.scala 71:109:@35365.4]
  wire [10:0] _T_80059; // @[Modules.scala 71:109:@35366.4]
  wire [10:0] buffer_14_699; // @[Modules.scala 71:109:@35367.4]
  wire [11:0] _T_80061; // @[Modules.scala 71:109:@35369.4]
  wire [10:0] _T_80062; // @[Modules.scala 71:109:@35370.4]
  wire [10:0] buffer_14_700; // @[Modules.scala 71:109:@35371.4]
  wire [11:0] _T_80064; // @[Modules.scala 71:109:@35373.4]
  wire [10:0] _T_80065; // @[Modules.scala 71:109:@35374.4]
  wire [10:0] buffer_14_701; // @[Modules.scala 71:109:@35375.4]
  wire [11:0] _T_80067; // @[Modules.scala 71:109:@35377.4]
  wire [10:0] _T_80068; // @[Modules.scala 71:109:@35378.4]
  wire [10:0] buffer_14_702; // @[Modules.scala 71:109:@35379.4]
  wire [11:0] _T_80070; // @[Modules.scala 71:109:@35381.4]
  wire [10:0] _T_80071; // @[Modules.scala 71:109:@35382.4]
  wire [10:0] buffer_14_703; // @[Modules.scala 71:109:@35383.4]
  wire [11:0] _T_80073; // @[Modules.scala 71:109:@35385.4]
  wire [10:0] _T_80074; // @[Modules.scala 71:109:@35386.4]
  wire [10:0] buffer_14_704; // @[Modules.scala 71:109:@35387.4]
  wire [11:0] _T_80076; // @[Modules.scala 71:109:@35389.4]
  wire [10:0] _T_80077; // @[Modules.scala 71:109:@35390.4]
  wire [10:0] buffer_14_705; // @[Modules.scala 71:109:@35391.4]
  wire [11:0] _T_80079; // @[Modules.scala 71:109:@35393.4]
  wire [10:0] _T_80080; // @[Modules.scala 71:109:@35394.4]
  wire [10:0] buffer_14_706; // @[Modules.scala 71:109:@35395.4]
  wire [11:0] _T_80082; // @[Modules.scala 71:109:@35397.4]
  wire [10:0] _T_80083; // @[Modules.scala 71:109:@35398.4]
  wire [10:0] buffer_14_707; // @[Modules.scala 71:109:@35399.4]
  wire [11:0] _T_80085; // @[Modules.scala 71:109:@35401.4]
  wire [10:0] _T_80086; // @[Modules.scala 71:109:@35402.4]
  wire [10:0] buffer_14_708; // @[Modules.scala 71:109:@35403.4]
  wire [11:0] _T_80088; // @[Modules.scala 71:109:@35405.4]
  wire [10:0] _T_80089; // @[Modules.scala 71:109:@35406.4]
  wire [10:0] buffer_14_709; // @[Modules.scala 71:109:@35407.4]
  wire [11:0] _T_80091; // @[Modules.scala 71:109:@35409.4]
  wire [10:0] _T_80092; // @[Modules.scala 71:109:@35410.4]
  wire [10:0] buffer_14_710; // @[Modules.scala 71:109:@35411.4]
  wire [11:0] _T_80094; // @[Modules.scala 71:109:@35413.4]
  wire [10:0] _T_80095; // @[Modules.scala 71:109:@35414.4]
  wire [10:0] buffer_14_711; // @[Modules.scala 71:109:@35415.4]
  wire [11:0] _T_80097; // @[Modules.scala 71:109:@35417.4]
  wire [10:0] _T_80098; // @[Modules.scala 71:109:@35418.4]
  wire [10:0] buffer_14_712; // @[Modules.scala 71:109:@35419.4]
  wire [11:0] _T_80100; // @[Modules.scala 71:109:@35421.4]
  wire [10:0] _T_80101; // @[Modules.scala 71:109:@35422.4]
  wire [10:0] buffer_14_713; // @[Modules.scala 71:109:@35423.4]
  wire [11:0] _T_80103; // @[Modules.scala 71:109:@35425.4]
  wire [10:0] _T_80104; // @[Modules.scala 71:109:@35426.4]
  wire [10:0] buffer_14_714; // @[Modules.scala 71:109:@35427.4]
  wire [11:0] _T_80106; // @[Modules.scala 71:109:@35429.4]
  wire [10:0] _T_80107; // @[Modules.scala 71:109:@35430.4]
  wire [10:0] buffer_14_715; // @[Modules.scala 71:109:@35431.4]
  wire [11:0] _T_80109; // @[Modules.scala 71:109:@35433.4]
  wire [10:0] _T_80110; // @[Modules.scala 71:109:@35434.4]
  wire [10:0] buffer_14_716; // @[Modules.scala 71:109:@35435.4]
  wire [11:0] _T_80112; // @[Modules.scala 71:109:@35437.4]
  wire [10:0] _T_80113; // @[Modules.scala 71:109:@35438.4]
  wire [10:0] buffer_14_717; // @[Modules.scala 71:109:@35439.4]
  wire [11:0] _T_80115; // @[Modules.scala 71:109:@35441.4]
  wire [10:0] _T_80116; // @[Modules.scala 71:109:@35442.4]
  wire [10:0] buffer_14_718; // @[Modules.scala 71:109:@35443.4]
  wire [11:0] _T_80118; // @[Modules.scala 71:109:@35445.4]
  wire [10:0] _T_80119; // @[Modules.scala 71:109:@35446.4]
  wire [10:0] buffer_14_719; // @[Modules.scala 71:109:@35447.4]
  wire [11:0] _T_80121; // @[Modules.scala 71:109:@35449.4]
  wire [10:0] _T_80122; // @[Modules.scala 71:109:@35450.4]
  wire [10:0] buffer_14_720; // @[Modules.scala 71:109:@35451.4]
  wire [11:0] _T_80124; // @[Modules.scala 71:109:@35453.4]
  wire [10:0] _T_80125; // @[Modules.scala 71:109:@35454.4]
  wire [10:0] buffer_14_721; // @[Modules.scala 71:109:@35455.4]
  wire [11:0] _T_80127; // @[Modules.scala 71:109:@35457.4]
  wire [10:0] _T_80128; // @[Modules.scala 71:109:@35458.4]
  wire [10:0] buffer_14_722; // @[Modules.scala 71:109:@35459.4]
  wire [11:0] _T_80130; // @[Modules.scala 71:109:@35461.4]
  wire [10:0] _T_80131; // @[Modules.scala 71:109:@35462.4]
  wire [10:0] buffer_14_723; // @[Modules.scala 71:109:@35463.4]
  wire [11:0] _T_80133; // @[Modules.scala 71:109:@35465.4]
  wire [10:0] _T_80134; // @[Modules.scala 71:109:@35466.4]
  wire [10:0] buffer_14_724; // @[Modules.scala 71:109:@35467.4]
  wire [11:0] _T_80136; // @[Modules.scala 71:109:@35469.4]
  wire [10:0] _T_80137; // @[Modules.scala 71:109:@35470.4]
  wire [10:0] buffer_14_725; // @[Modules.scala 71:109:@35471.4]
  wire [11:0] _T_80139; // @[Modules.scala 71:109:@35473.4]
  wire [10:0] _T_80140; // @[Modules.scala 71:109:@35474.4]
  wire [10:0] buffer_14_726; // @[Modules.scala 71:109:@35475.4]
  wire [11:0] _T_80142; // @[Modules.scala 71:109:@35477.4]
  wire [10:0] _T_80143; // @[Modules.scala 71:109:@35478.4]
  wire [10:0] buffer_14_727; // @[Modules.scala 71:109:@35479.4]
  wire [11:0] _T_80145; // @[Modules.scala 71:109:@35481.4]
  wire [10:0] _T_80146; // @[Modules.scala 71:109:@35482.4]
  wire [10:0] buffer_14_728; // @[Modules.scala 71:109:@35483.4]
  wire [11:0] _T_80148; // @[Modules.scala 71:109:@35485.4]
  wire [10:0] _T_80149; // @[Modules.scala 71:109:@35486.4]
  wire [10:0] buffer_14_729; // @[Modules.scala 71:109:@35487.4]
  wire [11:0] _T_80151; // @[Modules.scala 71:109:@35489.4]
  wire [10:0] _T_80152; // @[Modules.scala 71:109:@35490.4]
  wire [10:0] buffer_14_730; // @[Modules.scala 71:109:@35491.4]
  wire [11:0] _T_80154; // @[Modules.scala 71:109:@35493.4]
  wire [10:0] _T_80155; // @[Modules.scala 71:109:@35494.4]
  wire [10:0] buffer_14_731; // @[Modules.scala 71:109:@35495.4]
  wire [11:0] _T_80157; // @[Modules.scala 71:109:@35497.4]
  wire [10:0] _T_80158; // @[Modules.scala 71:109:@35498.4]
  wire [10:0] buffer_14_732; // @[Modules.scala 71:109:@35499.4]
  wire [11:0] _T_80160; // @[Modules.scala 71:109:@35501.4]
  wire [10:0] _T_80161; // @[Modules.scala 71:109:@35502.4]
  wire [10:0] buffer_14_733; // @[Modules.scala 71:109:@35503.4]
  wire [11:0] _T_80163; // @[Modules.scala 71:109:@35505.4]
  wire [10:0] _T_80164; // @[Modules.scala 71:109:@35506.4]
  wire [10:0] buffer_14_734; // @[Modules.scala 71:109:@35507.4]
  wire [11:0] _T_80166; // @[Modules.scala 78:156:@35510.4]
  wire [10:0] _T_80167; // @[Modules.scala 78:156:@35511.4]
  wire [10:0] buffer_14_736; // @[Modules.scala 78:156:@35512.4]
  wire [11:0] _T_80169; // @[Modules.scala 78:156:@35514.4]
  wire [10:0] _T_80170; // @[Modules.scala 78:156:@35515.4]
  wire [10:0] buffer_14_737; // @[Modules.scala 78:156:@35516.4]
  wire [11:0] _T_80172; // @[Modules.scala 78:156:@35518.4]
  wire [10:0] _T_80173; // @[Modules.scala 78:156:@35519.4]
  wire [10:0] buffer_14_738; // @[Modules.scala 78:156:@35520.4]
  wire [11:0] _T_80175; // @[Modules.scala 78:156:@35522.4]
  wire [10:0] _T_80176; // @[Modules.scala 78:156:@35523.4]
  wire [10:0] buffer_14_739; // @[Modules.scala 78:156:@35524.4]
  wire [11:0] _T_80178; // @[Modules.scala 78:156:@35526.4]
  wire [10:0] _T_80179; // @[Modules.scala 78:156:@35527.4]
  wire [10:0] buffer_14_740; // @[Modules.scala 78:156:@35528.4]
  wire [11:0] _T_80181; // @[Modules.scala 78:156:@35530.4]
  wire [10:0] _T_80182; // @[Modules.scala 78:156:@35531.4]
  wire [10:0] buffer_14_741; // @[Modules.scala 78:156:@35532.4]
  wire [11:0] _T_80184; // @[Modules.scala 78:156:@35534.4]
  wire [10:0] _T_80185; // @[Modules.scala 78:156:@35535.4]
  wire [10:0] buffer_14_742; // @[Modules.scala 78:156:@35536.4]
  wire [11:0] _T_80187; // @[Modules.scala 78:156:@35538.4]
  wire [10:0] _T_80188; // @[Modules.scala 78:156:@35539.4]
  wire [10:0] buffer_14_743; // @[Modules.scala 78:156:@35540.4]
  wire [11:0] _T_80190; // @[Modules.scala 78:156:@35542.4]
  wire [10:0] _T_80191; // @[Modules.scala 78:156:@35543.4]
  wire [10:0] buffer_14_744; // @[Modules.scala 78:156:@35544.4]
  wire [11:0] _T_80193; // @[Modules.scala 78:156:@35546.4]
  wire [10:0] _T_80194; // @[Modules.scala 78:156:@35547.4]
  wire [10:0] buffer_14_745; // @[Modules.scala 78:156:@35548.4]
  wire [11:0] _T_80196; // @[Modules.scala 78:156:@35550.4]
  wire [10:0] _T_80197; // @[Modules.scala 78:156:@35551.4]
  wire [10:0] buffer_14_746; // @[Modules.scala 78:156:@35552.4]
  wire [11:0] _T_80199; // @[Modules.scala 78:156:@35554.4]
  wire [10:0] _T_80200; // @[Modules.scala 78:156:@35555.4]
  wire [10:0] buffer_14_747; // @[Modules.scala 78:156:@35556.4]
  wire [11:0] _T_80202; // @[Modules.scala 78:156:@35558.4]
  wire [10:0] _T_80203; // @[Modules.scala 78:156:@35559.4]
  wire [10:0] buffer_14_748; // @[Modules.scala 78:156:@35560.4]
  wire [11:0] _T_80205; // @[Modules.scala 78:156:@35562.4]
  wire [10:0] _T_80206; // @[Modules.scala 78:156:@35563.4]
  wire [10:0] buffer_14_749; // @[Modules.scala 78:156:@35564.4]
  wire [11:0] _T_80208; // @[Modules.scala 78:156:@35566.4]
  wire [10:0] _T_80209; // @[Modules.scala 78:156:@35567.4]
  wire [10:0] buffer_14_750; // @[Modules.scala 78:156:@35568.4]
  wire [11:0] _T_80211; // @[Modules.scala 78:156:@35570.4]
  wire [10:0] _T_80212; // @[Modules.scala 78:156:@35571.4]
  wire [10:0] buffer_14_751; // @[Modules.scala 78:156:@35572.4]
  wire [11:0] _T_80214; // @[Modules.scala 78:156:@35574.4]
  wire [10:0] _T_80215; // @[Modules.scala 78:156:@35575.4]
  wire [10:0] buffer_14_752; // @[Modules.scala 78:156:@35576.4]
  wire [11:0] _T_80217; // @[Modules.scala 78:156:@35578.4]
  wire [10:0] _T_80218; // @[Modules.scala 78:156:@35579.4]
  wire [10:0] buffer_14_753; // @[Modules.scala 78:156:@35580.4]
  wire [11:0] _T_80220; // @[Modules.scala 78:156:@35582.4]
  wire [10:0] _T_80221; // @[Modules.scala 78:156:@35583.4]
  wire [10:0] buffer_14_754; // @[Modules.scala 78:156:@35584.4]
  wire [11:0] _T_80223; // @[Modules.scala 78:156:@35586.4]
  wire [10:0] _T_80224; // @[Modules.scala 78:156:@35587.4]
  wire [10:0] buffer_14_755; // @[Modules.scala 78:156:@35588.4]
  wire [11:0] _T_80226; // @[Modules.scala 78:156:@35590.4]
  wire [10:0] _T_80227; // @[Modules.scala 78:156:@35591.4]
  wire [10:0] buffer_14_756; // @[Modules.scala 78:156:@35592.4]
  wire [11:0] _T_80229; // @[Modules.scala 78:156:@35594.4]
  wire [10:0] _T_80230; // @[Modules.scala 78:156:@35595.4]
  wire [10:0] buffer_14_757; // @[Modules.scala 78:156:@35596.4]
  wire [11:0] _T_80232; // @[Modules.scala 78:156:@35598.4]
  wire [10:0] _T_80233; // @[Modules.scala 78:156:@35599.4]
  wire [10:0] buffer_14_758; // @[Modules.scala 78:156:@35600.4]
  wire [11:0] _T_80235; // @[Modules.scala 78:156:@35602.4]
  wire [10:0] _T_80236; // @[Modules.scala 78:156:@35603.4]
  wire [10:0] buffer_14_759; // @[Modules.scala 78:156:@35604.4]
  wire [11:0] _T_80238; // @[Modules.scala 78:156:@35606.4]
  wire [10:0] _T_80239; // @[Modules.scala 78:156:@35607.4]
  wire [10:0] buffer_14_760; // @[Modules.scala 78:156:@35608.4]
  wire [11:0] _T_80241; // @[Modules.scala 78:156:@35610.4]
  wire [10:0] _T_80242; // @[Modules.scala 78:156:@35611.4]
  wire [10:0] buffer_14_761; // @[Modules.scala 78:156:@35612.4]
  wire [11:0] _T_80244; // @[Modules.scala 78:156:@35614.4]
  wire [10:0] _T_80245; // @[Modules.scala 78:156:@35615.4]
  wire [10:0] buffer_14_762; // @[Modules.scala 78:156:@35616.4]
  wire [11:0] _T_80247; // @[Modules.scala 78:156:@35618.4]
  wire [10:0] _T_80248; // @[Modules.scala 78:156:@35619.4]
  wire [10:0] buffer_14_763; // @[Modules.scala 78:156:@35620.4]
  wire [11:0] _T_80250; // @[Modules.scala 78:156:@35622.4]
  wire [10:0] _T_80251; // @[Modules.scala 78:156:@35623.4]
  wire [10:0] buffer_14_764; // @[Modules.scala 78:156:@35624.4]
  wire [11:0] _T_80253; // @[Modules.scala 78:156:@35626.4]
  wire [10:0] _T_80254; // @[Modules.scala 78:156:@35627.4]
  wire [10:0] buffer_14_765; // @[Modules.scala 78:156:@35628.4]
  wire [11:0] _T_80256; // @[Modules.scala 78:156:@35630.4]
  wire [10:0] _T_80257; // @[Modules.scala 78:156:@35631.4]
  wire [10:0] buffer_14_766; // @[Modules.scala 78:156:@35632.4]
  wire [11:0] _T_80259; // @[Modules.scala 78:156:@35634.4]
  wire [10:0] _T_80260; // @[Modules.scala 78:156:@35635.4]
  wire [10:0] buffer_14_767; // @[Modules.scala 78:156:@35636.4]
  wire [11:0] _T_80262; // @[Modules.scala 78:156:@35638.4]
  wire [10:0] _T_80263; // @[Modules.scala 78:156:@35639.4]
  wire [10:0] buffer_14_768; // @[Modules.scala 78:156:@35640.4]
  wire [11:0] _T_80265; // @[Modules.scala 78:156:@35642.4]
  wire [10:0] _T_80266; // @[Modules.scala 78:156:@35643.4]
  wire [10:0] buffer_14_769; // @[Modules.scala 78:156:@35644.4]
  wire [11:0] _T_80268; // @[Modules.scala 78:156:@35646.4]
  wire [10:0] _T_80269; // @[Modules.scala 78:156:@35647.4]
  wire [10:0] buffer_14_770; // @[Modules.scala 78:156:@35648.4]
  wire [11:0] _T_80271; // @[Modules.scala 78:156:@35650.4]
  wire [10:0] _T_80272; // @[Modules.scala 78:156:@35651.4]
  wire [10:0] buffer_14_771; // @[Modules.scala 78:156:@35652.4]
  wire [11:0] _T_80274; // @[Modules.scala 78:156:@35654.4]
  wire [10:0] _T_80275; // @[Modules.scala 78:156:@35655.4]
  wire [10:0] buffer_14_772; // @[Modules.scala 78:156:@35656.4]
  wire [11:0] _T_80277; // @[Modules.scala 78:156:@35658.4]
  wire [10:0] _T_80278; // @[Modules.scala 78:156:@35659.4]
  wire [10:0] buffer_14_773; // @[Modules.scala 78:156:@35660.4]
  wire [11:0] _T_80280; // @[Modules.scala 78:156:@35662.4]
  wire [10:0] _T_80281; // @[Modules.scala 78:156:@35663.4]
  wire [10:0] buffer_14_774; // @[Modules.scala 78:156:@35664.4]
  wire [11:0] _T_80283; // @[Modules.scala 78:156:@35666.4]
  wire [10:0] _T_80284; // @[Modules.scala 78:156:@35667.4]
  wire [10:0] buffer_14_775; // @[Modules.scala 78:156:@35668.4]
  wire [11:0] _T_80286; // @[Modules.scala 78:156:@35670.4]
  wire [10:0] _T_80287; // @[Modules.scala 78:156:@35671.4]
  wire [10:0] buffer_14_776; // @[Modules.scala 78:156:@35672.4]
  wire [11:0] _T_80289; // @[Modules.scala 78:156:@35674.4]
  wire [10:0] _T_80290; // @[Modules.scala 78:156:@35675.4]
  wire [10:0] buffer_14_777; // @[Modules.scala 78:156:@35676.4]
  wire [11:0] _T_80292; // @[Modules.scala 78:156:@35678.4]
  wire [10:0] _T_80293; // @[Modules.scala 78:156:@35679.4]
  wire [10:0] buffer_14_778; // @[Modules.scala 78:156:@35680.4]
  wire [11:0] _T_80295; // @[Modules.scala 78:156:@35682.4]
  wire [10:0] _T_80296; // @[Modules.scala 78:156:@35683.4]
  wire [10:0] buffer_14_779; // @[Modules.scala 78:156:@35684.4]
  wire [11:0] _T_80298; // @[Modules.scala 78:156:@35686.4]
  wire [10:0] _T_80299; // @[Modules.scala 78:156:@35687.4]
  wire [10:0] buffer_14_780; // @[Modules.scala 78:156:@35688.4]
  wire [11:0] _T_80301; // @[Modules.scala 78:156:@35690.4]
  wire [10:0] _T_80302; // @[Modules.scala 78:156:@35691.4]
  wire [10:0] buffer_14_781; // @[Modules.scala 78:156:@35692.4]
  wire [11:0] _T_80304; // @[Modules.scala 78:156:@35694.4]
  wire [10:0] _T_80305; // @[Modules.scala 78:156:@35695.4]
  wire [10:0] buffer_14_782; // @[Modules.scala 78:156:@35696.4]
  wire [11:0] _T_80307; // @[Modules.scala 78:156:@35698.4]
  wire [10:0] _T_80308; // @[Modules.scala 78:156:@35699.4]
  wire [10:0] buffer_14_783; // @[Modules.scala 78:156:@35700.4]
  wire [5:0] _T_80589; // @[Modules.scala 37:46:@36108.4]
  wire [4:0] _T_80590; // @[Modules.scala 37:46:@36109.4]
  wire [4:0] _T_80591; // @[Modules.scala 37:46:@36110.4]
  wire [11:0] _T_80926; // @[Modules.scala 65:57:@36599.4]
  wire [10:0] _T_80927; // @[Modules.scala 65:57:@36600.4]
  wire [10:0] buffer_15_395; // @[Modules.scala 65:57:@36601.4]
  wire [11:0] _T_80929; // @[Modules.scala 65:57:@36603.4]
  wire [10:0] _T_80930; // @[Modules.scala 65:57:@36604.4]
  wire [10:0] buffer_15_396; // @[Modules.scala 65:57:@36605.4]
  wire [11:0] _T_80932; // @[Modules.scala 65:57:@36607.4]
  wire [10:0] _T_80933; // @[Modules.scala 65:57:@36608.4]
  wire [10:0] buffer_15_397; // @[Modules.scala 65:57:@36609.4]
  wire [11:0] _T_80935; // @[Modules.scala 65:57:@36611.4]
  wire [10:0] _T_80936; // @[Modules.scala 65:57:@36612.4]
  wire [10:0] buffer_15_398; // @[Modules.scala 65:57:@36613.4]
  wire [11:0] _T_80944; // @[Modules.scala 65:57:@36623.4]
  wire [10:0] _T_80945; // @[Modules.scala 65:57:@36624.4]
  wire [10:0] buffer_15_401; // @[Modules.scala 65:57:@36625.4]
  wire [11:0] _T_80950; // @[Modules.scala 65:57:@36631.4]
  wire [10:0] _T_80951; // @[Modules.scala 65:57:@36632.4]
  wire [10:0] buffer_15_403; // @[Modules.scala 65:57:@36633.4]
  wire [10:0] buffer_15_24; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_80953; // @[Modules.scala 65:57:@36635.4]
  wire [10:0] _T_80954; // @[Modules.scala 65:57:@36636.4]
  wire [10:0] buffer_15_404; // @[Modules.scala 65:57:@36637.4]
  wire [10:0] buffer_15_38; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_80974; // @[Modules.scala 65:57:@36663.4]
  wire [10:0] _T_80975; // @[Modules.scala 65:57:@36664.4]
  wire [10:0] buffer_15_411; // @[Modules.scala 65:57:@36665.4]
  wire [11:0] _T_80980; // @[Modules.scala 65:57:@36671.4]
  wire [10:0] _T_80981; // @[Modules.scala 65:57:@36672.4]
  wire [10:0] buffer_15_413; // @[Modules.scala 65:57:@36673.4]
  wire [11:0] _T_80983; // @[Modules.scala 65:57:@36675.4]
  wire [10:0] _T_80984; // @[Modules.scala 65:57:@36676.4]
  wire [10:0] buffer_15_414; // @[Modules.scala 65:57:@36677.4]
  wire [11:0] _T_81007; // @[Modules.scala 65:57:@36707.4]
  wire [10:0] _T_81008; // @[Modules.scala 65:57:@36708.4]
  wire [10:0] buffer_15_422; // @[Modules.scala 65:57:@36709.4]
  wire [11:0] _T_81013; // @[Modules.scala 65:57:@36715.4]
  wire [10:0] _T_81014; // @[Modules.scala 65:57:@36716.4]
  wire [10:0] buffer_15_424; // @[Modules.scala 65:57:@36717.4]
  wire [11:0] _T_81022; // @[Modules.scala 65:57:@36727.4]
  wire [10:0] _T_81023; // @[Modules.scala 65:57:@36728.4]
  wire [10:0] buffer_15_427; // @[Modules.scala 65:57:@36729.4]
  wire [11:0] _T_81031; // @[Modules.scala 65:57:@36739.4]
  wire [10:0] _T_81032; // @[Modules.scala 65:57:@36740.4]
  wire [10:0] buffer_15_430; // @[Modules.scala 65:57:@36741.4]
  wire [11:0] _T_81034; // @[Modules.scala 65:57:@36743.4]
  wire [10:0] _T_81035; // @[Modules.scala 65:57:@36744.4]
  wire [10:0] buffer_15_431; // @[Modules.scala 65:57:@36745.4]
  wire [11:0] _T_81043; // @[Modules.scala 65:57:@36755.4]
  wire [10:0] _T_81044; // @[Modules.scala 65:57:@36756.4]
  wire [10:0] buffer_15_434; // @[Modules.scala 65:57:@36757.4]
  wire [11:0] _T_81046; // @[Modules.scala 65:57:@36759.4]
  wire [10:0] _T_81047; // @[Modules.scala 65:57:@36760.4]
  wire [10:0] buffer_15_435; // @[Modules.scala 65:57:@36761.4]
  wire [11:0] _T_81049; // @[Modules.scala 65:57:@36763.4]
  wire [10:0] _T_81050; // @[Modules.scala 65:57:@36764.4]
  wire [10:0] buffer_15_436; // @[Modules.scala 65:57:@36765.4]
  wire [11:0] _T_81064; // @[Modules.scala 65:57:@36783.4]
  wire [10:0] _T_81065; // @[Modules.scala 65:57:@36784.4]
  wire [10:0] buffer_15_441; // @[Modules.scala 65:57:@36785.4]
  wire [11:0] _T_81067; // @[Modules.scala 65:57:@36787.4]
  wire [10:0] _T_81068; // @[Modules.scala 65:57:@36788.4]
  wire [10:0] buffer_15_442; // @[Modules.scala 65:57:@36789.4]
  wire [11:0] _T_81076; // @[Modules.scala 65:57:@36799.4]
  wire [10:0] _T_81077; // @[Modules.scala 65:57:@36800.4]
  wire [10:0] buffer_15_445; // @[Modules.scala 65:57:@36801.4]
  wire [11:0] _T_81091; // @[Modules.scala 65:57:@36819.4]
  wire [10:0] _T_81092; // @[Modules.scala 65:57:@36820.4]
  wire [10:0] buffer_15_450; // @[Modules.scala 65:57:@36821.4]
  wire [10:0] buffer_15_129; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81109; // @[Modules.scala 65:57:@36843.4]
  wire [10:0] _T_81110; // @[Modules.scala 65:57:@36844.4]
  wire [10:0] buffer_15_456; // @[Modules.scala 65:57:@36845.4]
  wire [11:0] _T_81130; // @[Modules.scala 65:57:@36871.4]
  wire [10:0] _T_81131; // @[Modules.scala 65:57:@36872.4]
  wire [10:0] buffer_15_463; // @[Modules.scala 65:57:@36873.4]
  wire [11:0] _T_81142; // @[Modules.scala 65:57:@36887.4]
  wire [10:0] _T_81143; // @[Modules.scala 65:57:@36888.4]
  wire [10:0] buffer_15_467; // @[Modules.scala 65:57:@36889.4]
  wire [11:0] _T_81151; // @[Modules.scala 65:57:@36899.4]
  wire [10:0] _T_81152; // @[Modules.scala 65:57:@36900.4]
  wire [10:0] buffer_15_470; // @[Modules.scala 65:57:@36901.4]
  wire [11:0] _T_81154; // @[Modules.scala 65:57:@36903.4]
  wire [10:0] _T_81155; // @[Modules.scala 65:57:@36904.4]
  wire [10:0] buffer_15_471; // @[Modules.scala 65:57:@36905.4]
  wire [11:0] _T_81160; // @[Modules.scala 65:57:@36911.4]
  wire [10:0] _T_81161; // @[Modules.scala 65:57:@36912.4]
  wire [10:0] buffer_15_473; // @[Modules.scala 65:57:@36913.4]
  wire [11:0] _T_81169; // @[Modules.scala 65:57:@36923.4]
  wire [10:0] _T_81170; // @[Modules.scala 65:57:@36924.4]
  wire [10:0] buffer_15_476; // @[Modules.scala 65:57:@36925.4]
  wire [11:0] _T_81187; // @[Modules.scala 65:57:@36947.4]
  wire [10:0] _T_81188; // @[Modules.scala 65:57:@36948.4]
  wire [10:0] buffer_15_482; // @[Modules.scala 65:57:@36949.4]
  wire [10:0] buffer_15_183; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81190; // @[Modules.scala 65:57:@36951.4]
  wire [10:0] _T_81191; // @[Modules.scala 65:57:@36952.4]
  wire [10:0] buffer_15_483; // @[Modules.scala 65:57:@36953.4]
  wire [11:0] _T_81193; // @[Modules.scala 65:57:@36955.4]
  wire [10:0] _T_81194; // @[Modules.scala 65:57:@36956.4]
  wire [10:0] buffer_15_484; // @[Modules.scala 65:57:@36957.4]
  wire [11:0] _T_81223; // @[Modules.scala 65:57:@36995.4]
  wire [10:0] _T_81224; // @[Modules.scala 65:57:@36996.4]
  wire [10:0] buffer_15_494; // @[Modules.scala 65:57:@36997.4]
  wire [11:0] _T_81244; // @[Modules.scala 65:57:@37023.4]
  wire [10:0] _T_81245; // @[Modules.scala 65:57:@37024.4]
  wire [10:0] buffer_15_501; // @[Modules.scala 65:57:@37025.4]
  wire [11:0] _T_81259; // @[Modules.scala 65:57:@37043.4]
  wire [10:0] _T_81260; // @[Modules.scala 65:57:@37044.4]
  wire [10:0] buffer_15_506; // @[Modules.scala 65:57:@37045.4]
  wire [11:0] _T_81262; // @[Modules.scala 65:57:@37047.4]
  wire [10:0] _T_81263; // @[Modules.scala 65:57:@37048.4]
  wire [10:0] buffer_15_507; // @[Modules.scala 65:57:@37049.4]
  wire [11:0] _T_81286; // @[Modules.scala 65:57:@37079.4]
  wire [10:0] _T_81287; // @[Modules.scala 65:57:@37080.4]
  wire [10:0] buffer_15_515; // @[Modules.scala 65:57:@37081.4]
  wire [10:0] buffer_15_249; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81289; // @[Modules.scala 65:57:@37083.4]
  wire [10:0] _T_81290; // @[Modules.scala 65:57:@37084.4]
  wire [10:0] buffer_15_516; // @[Modules.scala 65:57:@37085.4]
  wire [11:0] _T_81310; // @[Modules.scala 65:57:@37111.4]
  wire [10:0] _T_81311; // @[Modules.scala 65:57:@37112.4]
  wire [10:0] buffer_15_523; // @[Modules.scala 65:57:@37113.4]
  wire [11:0] _T_81325; // @[Modules.scala 65:57:@37131.4]
  wire [10:0] _T_81326; // @[Modules.scala 65:57:@37132.4]
  wire [10:0] buffer_15_528; // @[Modules.scala 65:57:@37133.4]
  wire [11:0] _T_81328; // @[Modules.scala 65:57:@37135.4]
  wire [10:0] _T_81329; // @[Modules.scala 65:57:@37136.4]
  wire [10:0] buffer_15_529; // @[Modules.scala 65:57:@37137.4]
  wire [11:0] _T_81343; // @[Modules.scala 65:57:@37155.4]
  wire [10:0] _T_81344; // @[Modules.scala 65:57:@37156.4]
  wire [10:0] buffer_15_534; // @[Modules.scala 65:57:@37157.4]
  wire [10:0] buffer_15_287; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81346; // @[Modules.scala 65:57:@37159.4]
  wire [10:0] _T_81347; // @[Modules.scala 65:57:@37160.4]
  wire [10:0] buffer_15_535; // @[Modules.scala 65:57:@37161.4]
  wire [11:0] _T_81349; // @[Modules.scala 65:57:@37163.4]
  wire [10:0] _T_81350; // @[Modules.scala 65:57:@37164.4]
  wire [10:0] buffer_15_536; // @[Modules.scala 65:57:@37165.4]
  wire [11:0] _T_81358; // @[Modules.scala 65:57:@37175.4]
  wire [10:0] _T_81359; // @[Modules.scala 65:57:@37176.4]
  wire [10:0] buffer_15_539; // @[Modules.scala 65:57:@37177.4]
  wire [11:0] _T_81364; // @[Modules.scala 65:57:@37183.4]
  wire [10:0] _T_81365; // @[Modules.scala 65:57:@37184.4]
  wire [10:0] buffer_15_541; // @[Modules.scala 65:57:@37185.4]
  wire [11:0] _T_81367; // @[Modules.scala 65:57:@37187.4]
  wire [10:0] _T_81368; // @[Modules.scala 65:57:@37188.4]
  wire [10:0] buffer_15_542; // @[Modules.scala 65:57:@37189.4]
  wire [11:0] _T_81370; // @[Modules.scala 65:57:@37191.4]
  wire [10:0] _T_81371; // @[Modules.scala 65:57:@37192.4]
  wire [10:0] buffer_15_543; // @[Modules.scala 65:57:@37193.4]
  wire [11:0] _T_81373; // @[Modules.scala 65:57:@37195.4]
  wire [10:0] _T_81374; // @[Modules.scala 65:57:@37196.4]
  wire [10:0] buffer_15_544; // @[Modules.scala 65:57:@37197.4]
  wire [10:0] buffer_15_308; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81379; // @[Modules.scala 65:57:@37203.4]
  wire [10:0] _T_81380; // @[Modules.scala 65:57:@37204.4]
  wire [10:0] buffer_15_546; // @[Modules.scala 65:57:@37205.4]
  wire [11:0] _T_81382; // @[Modules.scala 65:57:@37207.4]
  wire [10:0] _T_81383; // @[Modules.scala 65:57:@37208.4]
  wire [10:0] buffer_15_547; // @[Modules.scala 65:57:@37209.4]
  wire [11:0] _T_81388; // @[Modules.scala 65:57:@37215.4]
  wire [10:0] _T_81389; // @[Modules.scala 65:57:@37216.4]
  wire [10:0] buffer_15_549; // @[Modules.scala 65:57:@37217.4]
  wire [11:0] _T_81397; // @[Modules.scala 65:57:@37227.4]
  wire [10:0] _T_81398; // @[Modules.scala 65:57:@37228.4]
  wire [10:0] buffer_15_552; // @[Modules.scala 65:57:@37229.4]
  wire [11:0] _T_81400; // @[Modules.scala 65:57:@37231.4]
  wire [10:0] _T_81401; // @[Modules.scala 65:57:@37232.4]
  wire [10:0] buffer_15_553; // @[Modules.scala 65:57:@37233.4]
  wire [11:0] _T_81403; // @[Modules.scala 65:57:@37235.4]
  wire [10:0] _T_81404; // @[Modules.scala 65:57:@37236.4]
  wire [10:0] buffer_15_554; // @[Modules.scala 65:57:@37237.4]
  wire [10:0] buffer_15_338; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81424; // @[Modules.scala 65:57:@37263.4]
  wire [10:0] _T_81425; // @[Modules.scala 65:57:@37264.4]
  wire [10:0] buffer_15_561; // @[Modules.scala 65:57:@37265.4]
  wire [11:0] _T_81427; // @[Modules.scala 65:57:@37267.4]
  wire [10:0] _T_81428; // @[Modules.scala 65:57:@37268.4]
  wire [10:0] buffer_15_562; // @[Modules.scala 65:57:@37269.4]
  wire [11:0] _T_81442; // @[Modules.scala 65:57:@37287.4]
  wire [10:0] _T_81443; // @[Modules.scala 65:57:@37288.4]
  wire [10:0] buffer_15_567; // @[Modules.scala 65:57:@37289.4]
  wire [11:0] _T_81445; // @[Modules.scala 65:57:@37291.4]
  wire [10:0] _T_81446; // @[Modules.scala 65:57:@37292.4]
  wire [10:0] buffer_15_568; // @[Modules.scala 65:57:@37293.4]
  wire [10:0] buffer_15_356; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81451; // @[Modules.scala 65:57:@37299.4]
  wire [10:0] _T_81452; // @[Modules.scala 65:57:@37300.4]
  wire [10:0] buffer_15_570; // @[Modules.scala 65:57:@37301.4]
  wire [10:0] buffer_15_366; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81466; // @[Modules.scala 65:57:@37319.4]
  wire [10:0] _T_81467; // @[Modules.scala 65:57:@37320.4]
  wire [10:0] buffer_15_575; // @[Modules.scala 65:57:@37321.4]
  wire [10:0] buffer_15_389; // @[Modules.scala 32:22:@8.4]
  wire [11:0] _T_81499; // @[Modules.scala 65:57:@37363.4]
  wire [10:0] _T_81500; // @[Modules.scala 65:57:@37364.4]
  wire [10:0] buffer_15_586; // @[Modules.scala 65:57:@37365.4]
  wire [11:0] _T_81505; // @[Modules.scala 68:83:@37371.4]
  wire [10:0] _T_81506; // @[Modules.scala 68:83:@37372.4]
  wire [10:0] buffer_15_588; // @[Modules.scala 68:83:@37373.4]
  wire [11:0] _T_81508; // @[Modules.scala 68:83:@37375.4]
  wire [10:0] _T_81509; // @[Modules.scala 68:83:@37376.4]
  wire [10:0] buffer_15_589; // @[Modules.scala 68:83:@37377.4]
  wire [11:0] _T_81511; // @[Modules.scala 68:83:@37379.4]
  wire [10:0] _T_81512; // @[Modules.scala 68:83:@37380.4]
  wire [10:0] buffer_15_590; // @[Modules.scala 68:83:@37381.4]
  wire [11:0] _T_81514; // @[Modules.scala 68:83:@37383.4]
  wire [10:0] _T_81515; // @[Modules.scala 68:83:@37384.4]
  wire [10:0] buffer_15_591; // @[Modules.scala 68:83:@37385.4]
  wire [11:0] _T_81517; // @[Modules.scala 68:83:@37387.4]
  wire [10:0] _T_81518; // @[Modules.scala 68:83:@37388.4]
  wire [10:0] buffer_15_592; // @[Modules.scala 68:83:@37389.4]
  wire [11:0] _T_81520; // @[Modules.scala 68:83:@37391.4]
  wire [10:0] _T_81521; // @[Modules.scala 68:83:@37392.4]
  wire [10:0] buffer_15_593; // @[Modules.scala 68:83:@37393.4]
  wire [11:0] _T_81523; // @[Modules.scala 68:83:@37395.4]
  wire [10:0] _T_81524; // @[Modules.scala 68:83:@37396.4]
  wire [10:0] buffer_15_594; // @[Modules.scala 68:83:@37397.4]
  wire [11:0] _T_81526; // @[Modules.scala 68:83:@37399.4]
  wire [10:0] _T_81527; // @[Modules.scala 68:83:@37400.4]
  wire [10:0] buffer_15_595; // @[Modules.scala 68:83:@37401.4]
  wire [11:0] _T_81532; // @[Modules.scala 68:83:@37407.4]
  wire [10:0] _T_81533; // @[Modules.scala 68:83:@37408.4]
  wire [10:0] buffer_15_597; // @[Modules.scala 68:83:@37409.4]
  wire [11:0] _T_81535; // @[Modules.scala 68:83:@37411.4]
  wire [10:0] _T_81536; // @[Modules.scala 68:83:@37412.4]
  wire [10:0] buffer_15_598; // @[Modules.scala 68:83:@37413.4]
  wire [11:0] _T_81538; // @[Modules.scala 68:83:@37415.4]
  wire [10:0] _T_81539; // @[Modules.scala 68:83:@37416.4]
  wire [10:0] buffer_15_599; // @[Modules.scala 68:83:@37417.4]
  wire [11:0] _T_81547; // @[Modules.scala 68:83:@37427.4]
  wire [10:0] _T_81548; // @[Modules.scala 68:83:@37428.4]
  wire [10:0] buffer_15_602; // @[Modules.scala 68:83:@37429.4]
  wire [11:0] _T_81550; // @[Modules.scala 68:83:@37431.4]
  wire [10:0] _T_81551; // @[Modules.scala 68:83:@37432.4]
  wire [10:0] buffer_15_603; // @[Modules.scala 68:83:@37433.4]
  wire [11:0] _T_81553; // @[Modules.scala 68:83:@37435.4]
  wire [10:0] _T_81554; // @[Modules.scala 68:83:@37436.4]
  wire [10:0] buffer_15_604; // @[Modules.scala 68:83:@37437.4]
  wire [11:0] _T_81556; // @[Modules.scala 68:83:@37439.4]
  wire [10:0] _T_81557; // @[Modules.scala 68:83:@37440.4]
  wire [10:0] buffer_15_605; // @[Modules.scala 68:83:@37441.4]
  wire [11:0] _T_81559; // @[Modules.scala 68:83:@37443.4]
  wire [10:0] _T_81560; // @[Modules.scala 68:83:@37444.4]
  wire [10:0] buffer_15_606; // @[Modules.scala 68:83:@37445.4]
  wire [11:0] _T_81562; // @[Modules.scala 68:83:@37447.4]
  wire [10:0] _T_81563; // @[Modules.scala 68:83:@37448.4]
  wire [10:0] buffer_15_607; // @[Modules.scala 68:83:@37449.4]
  wire [11:0] _T_81565; // @[Modules.scala 68:83:@37451.4]
  wire [10:0] _T_81566; // @[Modules.scala 68:83:@37452.4]
  wire [10:0] buffer_15_608; // @[Modules.scala 68:83:@37453.4]
  wire [11:0] _T_81568; // @[Modules.scala 68:83:@37455.4]
  wire [10:0] _T_81569; // @[Modules.scala 68:83:@37456.4]
  wire [10:0] buffer_15_609; // @[Modules.scala 68:83:@37457.4]
  wire [11:0] _T_81571; // @[Modules.scala 68:83:@37459.4]
  wire [10:0] _T_81572; // @[Modules.scala 68:83:@37460.4]
  wire [10:0] buffer_15_610; // @[Modules.scala 68:83:@37461.4]
  wire [11:0] _T_81574; // @[Modules.scala 68:83:@37463.4]
  wire [10:0] _T_81575; // @[Modules.scala 68:83:@37464.4]
  wire [10:0] buffer_15_611; // @[Modules.scala 68:83:@37465.4]
  wire [11:0] _T_81577; // @[Modules.scala 68:83:@37467.4]
  wire [10:0] _T_81578; // @[Modules.scala 68:83:@37468.4]
  wire [10:0] buffer_15_612; // @[Modules.scala 68:83:@37469.4]
  wire [11:0] _T_81580; // @[Modules.scala 68:83:@37471.4]
  wire [10:0] _T_81581; // @[Modules.scala 68:83:@37472.4]
  wire [10:0] buffer_15_613; // @[Modules.scala 68:83:@37473.4]
  wire [11:0] _T_81583; // @[Modules.scala 68:83:@37475.4]
  wire [10:0] _T_81584; // @[Modules.scala 68:83:@37476.4]
  wire [10:0] buffer_15_614; // @[Modules.scala 68:83:@37477.4]
  wire [11:0] _T_81586; // @[Modules.scala 68:83:@37479.4]
  wire [10:0] _T_81587; // @[Modules.scala 68:83:@37480.4]
  wire [10:0] buffer_15_615; // @[Modules.scala 68:83:@37481.4]
  wire [11:0] _T_81589; // @[Modules.scala 68:83:@37483.4]
  wire [10:0] _T_81590; // @[Modules.scala 68:83:@37484.4]
  wire [10:0] buffer_15_616; // @[Modules.scala 68:83:@37485.4]
  wire [11:0] _T_81592; // @[Modules.scala 68:83:@37487.4]
  wire [10:0] _T_81593; // @[Modules.scala 68:83:@37488.4]
  wire [10:0] buffer_15_617; // @[Modules.scala 68:83:@37489.4]
  wire [11:0] _T_81595; // @[Modules.scala 68:83:@37491.4]
  wire [10:0] _T_81596; // @[Modules.scala 68:83:@37492.4]
  wire [10:0] buffer_15_618; // @[Modules.scala 68:83:@37493.4]
  wire [11:0] _T_81601; // @[Modules.scala 68:83:@37499.4]
  wire [10:0] _T_81602; // @[Modules.scala 68:83:@37500.4]
  wire [10:0] buffer_15_620; // @[Modules.scala 68:83:@37501.4]
  wire [11:0] _T_81604; // @[Modules.scala 68:83:@37503.4]
  wire [10:0] _T_81605; // @[Modules.scala 68:83:@37504.4]
  wire [10:0] buffer_15_621; // @[Modules.scala 68:83:@37505.4]
  wire [11:0] _T_81610; // @[Modules.scala 68:83:@37511.4]
  wire [10:0] _T_81611; // @[Modules.scala 68:83:@37512.4]
  wire [10:0] buffer_15_623; // @[Modules.scala 68:83:@37513.4]
  wire [11:0] _T_81616; // @[Modules.scala 68:83:@37519.4]
  wire [10:0] _T_81617; // @[Modules.scala 68:83:@37520.4]
  wire [10:0] buffer_15_625; // @[Modules.scala 68:83:@37521.4]
  wire [11:0] _T_81619; // @[Modules.scala 68:83:@37523.4]
  wire [10:0] _T_81620; // @[Modules.scala 68:83:@37524.4]
  wire [10:0] buffer_15_626; // @[Modules.scala 68:83:@37525.4]
  wire [11:0] _T_81622; // @[Modules.scala 68:83:@37527.4]
  wire [10:0] _T_81623; // @[Modules.scala 68:83:@37528.4]
  wire [10:0] buffer_15_627; // @[Modules.scala 68:83:@37529.4]
  wire [11:0] _T_81625; // @[Modules.scala 68:83:@37531.4]
  wire [10:0] _T_81626; // @[Modules.scala 68:83:@37532.4]
  wire [10:0] buffer_15_628; // @[Modules.scala 68:83:@37533.4]
  wire [11:0] _T_81628; // @[Modules.scala 68:83:@37535.4]
  wire [10:0] _T_81629; // @[Modules.scala 68:83:@37536.4]
  wire [10:0] buffer_15_629; // @[Modules.scala 68:83:@37537.4]
  wire [11:0] _T_81631; // @[Modules.scala 68:83:@37539.4]
  wire [10:0] _T_81632; // @[Modules.scala 68:83:@37540.4]
  wire [10:0] buffer_15_630; // @[Modules.scala 68:83:@37541.4]
  wire [11:0] _T_81637; // @[Modules.scala 68:83:@37547.4]
  wire [10:0] _T_81638; // @[Modules.scala 68:83:@37548.4]
  wire [10:0] buffer_15_632; // @[Modules.scala 68:83:@37549.4]
  wire [11:0] _T_81640; // @[Modules.scala 68:83:@37551.4]
  wire [10:0] _T_81641; // @[Modules.scala 68:83:@37552.4]
  wire [10:0] buffer_15_633; // @[Modules.scala 68:83:@37553.4]
  wire [11:0] _T_81643; // @[Modules.scala 68:83:@37555.4]
  wire [10:0] _T_81644; // @[Modules.scala 68:83:@37556.4]
  wire [10:0] buffer_15_634; // @[Modules.scala 68:83:@37557.4]
  wire [11:0] _T_81649; // @[Modules.scala 68:83:@37563.4]
  wire [10:0] _T_81650; // @[Modules.scala 68:83:@37564.4]
  wire [10:0] buffer_15_636; // @[Modules.scala 68:83:@37565.4]
  wire [11:0] _T_81658; // @[Modules.scala 68:83:@37575.4]
  wire [10:0] _T_81659; // @[Modules.scala 68:83:@37576.4]
  wire [10:0] buffer_15_639; // @[Modules.scala 68:83:@37577.4]
  wire [11:0] _T_81661; // @[Modules.scala 68:83:@37579.4]
  wire [10:0] _T_81662; // @[Modules.scala 68:83:@37580.4]
  wire [10:0] buffer_15_640; // @[Modules.scala 68:83:@37581.4]
  wire [11:0] _T_81667; // @[Modules.scala 68:83:@37587.4]
  wire [10:0] _T_81668; // @[Modules.scala 68:83:@37588.4]
  wire [10:0] buffer_15_642; // @[Modules.scala 68:83:@37589.4]
  wire [11:0] _T_81670; // @[Modules.scala 68:83:@37591.4]
  wire [10:0] _T_81671; // @[Modules.scala 68:83:@37592.4]
  wire [10:0] buffer_15_643; // @[Modules.scala 68:83:@37593.4]
  wire [11:0] _T_81676; // @[Modules.scala 68:83:@37599.4]
  wire [10:0] _T_81677; // @[Modules.scala 68:83:@37600.4]
  wire [10:0] buffer_15_645; // @[Modules.scala 68:83:@37601.4]
  wire [11:0] _T_81679; // @[Modules.scala 68:83:@37603.4]
  wire [10:0] _T_81680; // @[Modules.scala 68:83:@37604.4]
  wire [10:0] buffer_15_646; // @[Modules.scala 68:83:@37605.4]
  wire [11:0] _T_81688; // @[Modules.scala 68:83:@37615.4]
  wire [10:0] _T_81689; // @[Modules.scala 68:83:@37616.4]
  wire [10:0] buffer_15_649; // @[Modules.scala 68:83:@37617.4]
  wire [11:0] _T_81691; // @[Modules.scala 68:83:@37619.4]
  wire [10:0] _T_81692; // @[Modules.scala 68:83:@37620.4]
  wire [10:0] buffer_15_650; // @[Modules.scala 68:83:@37621.4]
  wire [11:0] _T_81694; // @[Modules.scala 68:83:@37623.4]
  wire [10:0] _T_81695; // @[Modules.scala 68:83:@37624.4]
  wire [10:0] buffer_15_651; // @[Modules.scala 68:83:@37625.4]
  wire [11:0] _T_81697; // @[Modules.scala 68:83:@37627.4]
  wire [10:0] _T_81698; // @[Modules.scala 68:83:@37628.4]
  wire [10:0] buffer_15_652; // @[Modules.scala 68:83:@37629.4]
  wire [11:0] _T_81700; // @[Modules.scala 68:83:@37631.4]
  wire [10:0] _T_81701; // @[Modules.scala 68:83:@37632.4]
  wire [10:0] buffer_15_653; // @[Modules.scala 68:83:@37633.4]
  wire [11:0] _T_81706; // @[Modules.scala 68:83:@37639.4]
  wire [10:0] _T_81707; // @[Modules.scala 68:83:@37640.4]
  wire [10:0] buffer_15_655; // @[Modules.scala 68:83:@37641.4]
  wire [11:0] _T_81709; // @[Modules.scala 68:83:@37643.4]
  wire [10:0] _T_81710; // @[Modules.scala 68:83:@37644.4]
  wire [10:0] buffer_15_656; // @[Modules.scala 68:83:@37645.4]
  wire [11:0] _T_81718; // @[Modules.scala 68:83:@37655.4]
  wire [10:0] _T_81719; // @[Modules.scala 68:83:@37656.4]
  wire [10:0] buffer_15_659; // @[Modules.scala 68:83:@37657.4]
  wire [11:0] _T_81721; // @[Modules.scala 68:83:@37659.4]
  wire [10:0] _T_81722; // @[Modules.scala 68:83:@37660.4]
  wire [10:0] buffer_15_660; // @[Modules.scala 68:83:@37661.4]
  wire [11:0] _T_81724; // @[Modules.scala 68:83:@37663.4]
  wire [10:0] _T_81725; // @[Modules.scala 68:83:@37664.4]
  wire [10:0] buffer_15_661; // @[Modules.scala 68:83:@37665.4]
  wire [11:0] _T_81727; // @[Modules.scala 68:83:@37667.4]
  wire [10:0] _T_81728; // @[Modules.scala 68:83:@37668.4]
  wire [10:0] buffer_15_662; // @[Modules.scala 68:83:@37669.4]
  wire [11:0] _T_81730; // @[Modules.scala 68:83:@37671.4]
  wire [10:0] _T_81731; // @[Modules.scala 68:83:@37672.4]
  wire [10:0] buffer_15_663; // @[Modules.scala 68:83:@37673.4]
  wire [11:0] _T_81733; // @[Modules.scala 68:83:@37675.4]
  wire [10:0] _T_81734; // @[Modules.scala 68:83:@37676.4]
  wire [10:0] buffer_15_664; // @[Modules.scala 68:83:@37677.4]
  wire [11:0] _T_81736; // @[Modules.scala 68:83:@37679.4]
  wire [10:0] _T_81737; // @[Modules.scala 68:83:@37680.4]
  wire [10:0] buffer_15_665; // @[Modules.scala 68:83:@37681.4]
  wire [11:0] _T_81739; // @[Modules.scala 68:83:@37683.4]
  wire [10:0] _T_81740; // @[Modules.scala 68:83:@37684.4]
  wire [10:0] buffer_15_666; // @[Modules.scala 68:83:@37685.4]
  wire [11:0] _T_81745; // @[Modules.scala 68:83:@37691.4]
  wire [10:0] _T_81746; // @[Modules.scala 68:83:@37692.4]
  wire [10:0] buffer_15_668; // @[Modules.scala 68:83:@37693.4]
  wire [11:0] _T_81748; // @[Modules.scala 68:83:@37695.4]
  wire [10:0] _T_81749; // @[Modules.scala 68:83:@37696.4]
  wire [10:0] buffer_15_669; // @[Modules.scala 68:83:@37697.4]
  wire [11:0] _T_81754; // @[Modules.scala 68:83:@37703.4]
  wire [10:0] _T_81755; // @[Modules.scala 68:83:@37704.4]
  wire [10:0] buffer_15_671; // @[Modules.scala 68:83:@37705.4]
  wire [11:0] _T_81757; // @[Modules.scala 68:83:@37707.4]
  wire [10:0] _T_81758; // @[Modules.scala 68:83:@37708.4]
  wire [10:0] buffer_15_672; // @[Modules.scala 68:83:@37709.4]
  wire [11:0] _T_81760; // @[Modules.scala 68:83:@37711.4]
  wire [10:0] _T_81761; // @[Modules.scala 68:83:@37712.4]
  wire [10:0] buffer_15_673; // @[Modules.scala 68:83:@37713.4]
  wire [11:0] _T_81766; // @[Modules.scala 68:83:@37719.4]
  wire [10:0] _T_81767; // @[Modules.scala 68:83:@37720.4]
  wire [10:0] buffer_15_675; // @[Modules.scala 68:83:@37721.4]
  wire [11:0] _T_81769; // @[Modules.scala 68:83:@37723.4]
  wire [10:0] _T_81770; // @[Modules.scala 68:83:@37724.4]
  wire [10:0] buffer_15_676; // @[Modules.scala 68:83:@37725.4]
  wire [11:0] _T_81772; // @[Modules.scala 68:83:@37727.4]
  wire [10:0] _T_81773; // @[Modules.scala 68:83:@37728.4]
  wire [10:0] buffer_15_677; // @[Modules.scala 68:83:@37729.4]
  wire [11:0] _T_81778; // @[Modules.scala 68:83:@37735.4]
  wire [10:0] _T_81779; // @[Modules.scala 68:83:@37736.4]
  wire [10:0] buffer_15_679; // @[Modules.scala 68:83:@37737.4]
  wire [11:0] _T_81796; // @[Modules.scala 68:83:@37759.4]
  wire [10:0] _T_81797; // @[Modules.scala 68:83:@37760.4]
  wire [10:0] buffer_15_685; // @[Modules.scala 68:83:@37761.4]
  wire [11:0] _T_81799; // @[Modules.scala 71:109:@37763.4]
  wire [10:0] _T_81800; // @[Modules.scala 71:109:@37764.4]
  wire [10:0] buffer_15_686; // @[Modules.scala 71:109:@37765.4]
  wire [11:0] _T_81802; // @[Modules.scala 71:109:@37767.4]
  wire [10:0] _T_81803; // @[Modules.scala 71:109:@37768.4]
  wire [10:0] buffer_15_687; // @[Modules.scala 71:109:@37769.4]
  wire [11:0] _T_81805; // @[Modules.scala 71:109:@37771.4]
  wire [10:0] _T_81806; // @[Modules.scala 71:109:@37772.4]
  wire [10:0] buffer_15_688; // @[Modules.scala 71:109:@37773.4]
  wire [11:0] _T_81808; // @[Modules.scala 71:109:@37775.4]
  wire [10:0] _T_81809; // @[Modules.scala 71:109:@37776.4]
  wire [10:0] buffer_15_689; // @[Modules.scala 71:109:@37777.4]
  wire [11:0] _T_81811; // @[Modules.scala 71:109:@37779.4]
  wire [10:0] _T_81812; // @[Modules.scala 71:109:@37780.4]
  wire [10:0] buffer_15_690; // @[Modules.scala 71:109:@37781.4]
  wire [11:0] _T_81814; // @[Modules.scala 71:109:@37783.4]
  wire [10:0] _T_81815; // @[Modules.scala 71:109:@37784.4]
  wire [10:0] buffer_15_691; // @[Modules.scala 71:109:@37785.4]
  wire [11:0] _T_81820; // @[Modules.scala 71:109:@37791.4]
  wire [10:0] _T_81821; // @[Modules.scala 71:109:@37792.4]
  wire [10:0] buffer_15_693; // @[Modules.scala 71:109:@37793.4]
  wire [11:0] _T_81823; // @[Modules.scala 71:109:@37795.4]
  wire [10:0] _T_81824; // @[Modules.scala 71:109:@37796.4]
  wire [10:0] buffer_15_694; // @[Modules.scala 71:109:@37797.4]
  wire [11:0] _T_81826; // @[Modules.scala 71:109:@37799.4]
  wire [10:0] _T_81827; // @[Modules.scala 71:109:@37800.4]
  wire [10:0] buffer_15_695; // @[Modules.scala 71:109:@37801.4]
  wire [11:0] _T_81829; // @[Modules.scala 71:109:@37803.4]
  wire [10:0] _T_81830; // @[Modules.scala 71:109:@37804.4]
  wire [10:0] buffer_15_696; // @[Modules.scala 71:109:@37805.4]
  wire [11:0] _T_81832; // @[Modules.scala 71:109:@37807.4]
  wire [10:0] _T_81833; // @[Modules.scala 71:109:@37808.4]
  wire [10:0] buffer_15_697; // @[Modules.scala 71:109:@37809.4]
  wire [11:0] _T_81835; // @[Modules.scala 71:109:@37811.4]
  wire [10:0] _T_81836; // @[Modules.scala 71:109:@37812.4]
  wire [10:0] buffer_15_698; // @[Modules.scala 71:109:@37813.4]
  wire [11:0] _T_81838; // @[Modules.scala 71:109:@37815.4]
  wire [10:0] _T_81839; // @[Modules.scala 71:109:@37816.4]
  wire [10:0] buffer_15_699; // @[Modules.scala 71:109:@37817.4]
  wire [11:0] _T_81841; // @[Modules.scala 71:109:@37819.4]
  wire [10:0] _T_81842; // @[Modules.scala 71:109:@37820.4]
  wire [10:0] buffer_15_700; // @[Modules.scala 71:109:@37821.4]
  wire [11:0] _T_81844; // @[Modules.scala 71:109:@37823.4]
  wire [10:0] _T_81845; // @[Modules.scala 71:109:@37824.4]
  wire [10:0] buffer_15_701; // @[Modules.scala 71:109:@37825.4]
  wire [11:0] _T_81847; // @[Modules.scala 71:109:@37827.4]
  wire [10:0] _T_81848; // @[Modules.scala 71:109:@37828.4]
  wire [10:0] buffer_15_702; // @[Modules.scala 71:109:@37829.4]
  wire [11:0] _T_81850; // @[Modules.scala 71:109:@37831.4]
  wire [10:0] _T_81851; // @[Modules.scala 71:109:@37832.4]
  wire [10:0] buffer_15_703; // @[Modules.scala 71:109:@37833.4]
  wire [11:0] _T_81853; // @[Modules.scala 71:109:@37835.4]
  wire [10:0] _T_81854; // @[Modules.scala 71:109:@37836.4]
  wire [10:0] buffer_15_704; // @[Modules.scala 71:109:@37837.4]
  wire [11:0] _T_81856; // @[Modules.scala 71:109:@37839.4]
  wire [10:0] _T_81857; // @[Modules.scala 71:109:@37840.4]
  wire [10:0] buffer_15_705; // @[Modules.scala 71:109:@37841.4]
  wire [11:0] _T_81859; // @[Modules.scala 71:109:@37843.4]
  wire [10:0] _T_81860; // @[Modules.scala 71:109:@37844.4]
  wire [10:0] buffer_15_706; // @[Modules.scala 71:109:@37845.4]
  wire [11:0] _T_81862; // @[Modules.scala 71:109:@37847.4]
  wire [10:0] _T_81863; // @[Modules.scala 71:109:@37848.4]
  wire [10:0] buffer_15_707; // @[Modules.scala 71:109:@37849.4]
  wire [11:0] _T_81865; // @[Modules.scala 71:109:@37851.4]
  wire [10:0] _T_81866; // @[Modules.scala 71:109:@37852.4]
  wire [10:0] buffer_15_708; // @[Modules.scala 71:109:@37853.4]
  wire [11:0] _T_81868; // @[Modules.scala 71:109:@37855.4]
  wire [10:0] _T_81869; // @[Modules.scala 71:109:@37856.4]
  wire [10:0] buffer_15_709; // @[Modules.scala 71:109:@37857.4]
  wire [11:0] _T_81871; // @[Modules.scala 71:109:@37859.4]
  wire [10:0] _T_81872; // @[Modules.scala 71:109:@37860.4]
  wire [10:0] buffer_15_710; // @[Modules.scala 71:109:@37861.4]
  wire [11:0] _T_81874; // @[Modules.scala 71:109:@37863.4]
  wire [10:0] _T_81875; // @[Modules.scala 71:109:@37864.4]
  wire [10:0] buffer_15_711; // @[Modules.scala 71:109:@37865.4]
  wire [11:0] _T_81877; // @[Modules.scala 71:109:@37867.4]
  wire [10:0] _T_81878; // @[Modules.scala 71:109:@37868.4]
  wire [10:0] buffer_15_712; // @[Modules.scala 71:109:@37869.4]
  wire [11:0] _T_81880; // @[Modules.scala 71:109:@37871.4]
  wire [10:0] _T_81881; // @[Modules.scala 71:109:@37872.4]
  wire [10:0] buffer_15_713; // @[Modules.scala 71:109:@37873.4]
  wire [11:0] _T_81883; // @[Modules.scala 71:109:@37875.4]
  wire [10:0] _T_81884; // @[Modules.scala 71:109:@37876.4]
  wire [10:0] buffer_15_714; // @[Modules.scala 71:109:@37877.4]
  wire [11:0] _T_81886; // @[Modules.scala 71:109:@37879.4]
  wire [10:0] _T_81887; // @[Modules.scala 71:109:@37880.4]
  wire [10:0] buffer_15_715; // @[Modules.scala 71:109:@37881.4]
  wire [11:0] _T_81889; // @[Modules.scala 71:109:@37883.4]
  wire [10:0] _T_81890; // @[Modules.scala 71:109:@37884.4]
  wire [10:0] buffer_15_716; // @[Modules.scala 71:109:@37885.4]
  wire [11:0] _T_81892; // @[Modules.scala 71:109:@37887.4]
  wire [10:0] _T_81893; // @[Modules.scala 71:109:@37888.4]
  wire [10:0] buffer_15_717; // @[Modules.scala 71:109:@37889.4]
  wire [11:0] _T_81895; // @[Modules.scala 71:109:@37891.4]
  wire [10:0] _T_81896; // @[Modules.scala 71:109:@37892.4]
  wire [10:0] buffer_15_718; // @[Modules.scala 71:109:@37893.4]
  wire [11:0] _T_81898; // @[Modules.scala 71:109:@37895.4]
  wire [10:0] _T_81899; // @[Modules.scala 71:109:@37896.4]
  wire [10:0] buffer_15_719; // @[Modules.scala 71:109:@37897.4]
  wire [11:0] _T_81901; // @[Modules.scala 71:109:@37899.4]
  wire [10:0] _T_81902; // @[Modules.scala 71:109:@37900.4]
  wire [10:0] buffer_15_720; // @[Modules.scala 71:109:@37901.4]
  wire [11:0] _T_81904; // @[Modules.scala 71:109:@37903.4]
  wire [10:0] _T_81905; // @[Modules.scala 71:109:@37904.4]
  wire [10:0] buffer_15_721; // @[Modules.scala 71:109:@37905.4]
  wire [11:0] _T_81907; // @[Modules.scala 71:109:@37907.4]
  wire [10:0] _T_81908; // @[Modules.scala 71:109:@37908.4]
  wire [10:0] buffer_15_722; // @[Modules.scala 71:109:@37909.4]
  wire [11:0] _T_81910; // @[Modules.scala 71:109:@37911.4]
  wire [10:0] _T_81911; // @[Modules.scala 71:109:@37912.4]
  wire [10:0] buffer_15_723; // @[Modules.scala 71:109:@37913.4]
  wire [11:0] _T_81913; // @[Modules.scala 71:109:@37915.4]
  wire [10:0] _T_81914; // @[Modules.scala 71:109:@37916.4]
  wire [10:0] buffer_15_724; // @[Modules.scala 71:109:@37917.4]
  wire [11:0] _T_81916; // @[Modules.scala 71:109:@37919.4]
  wire [10:0] _T_81917; // @[Modules.scala 71:109:@37920.4]
  wire [10:0] buffer_15_725; // @[Modules.scala 71:109:@37921.4]
  wire [11:0] _T_81919; // @[Modules.scala 71:109:@37923.4]
  wire [10:0] _T_81920; // @[Modules.scala 71:109:@37924.4]
  wire [10:0] buffer_15_726; // @[Modules.scala 71:109:@37925.4]
  wire [11:0] _T_81922; // @[Modules.scala 71:109:@37927.4]
  wire [10:0] _T_81923; // @[Modules.scala 71:109:@37928.4]
  wire [10:0] buffer_15_727; // @[Modules.scala 71:109:@37929.4]
  wire [11:0] _T_81925; // @[Modules.scala 71:109:@37931.4]
  wire [10:0] _T_81926; // @[Modules.scala 71:109:@37932.4]
  wire [10:0] buffer_15_728; // @[Modules.scala 71:109:@37933.4]
  wire [11:0] _T_81928; // @[Modules.scala 71:109:@37935.4]
  wire [10:0] _T_81929; // @[Modules.scala 71:109:@37936.4]
  wire [10:0] buffer_15_729; // @[Modules.scala 71:109:@37937.4]
  wire [11:0] _T_81931; // @[Modules.scala 71:109:@37939.4]
  wire [10:0] _T_81932; // @[Modules.scala 71:109:@37940.4]
  wire [10:0] buffer_15_730; // @[Modules.scala 71:109:@37941.4]
  wire [11:0] _T_81934; // @[Modules.scala 71:109:@37943.4]
  wire [10:0] _T_81935; // @[Modules.scala 71:109:@37944.4]
  wire [10:0] buffer_15_731; // @[Modules.scala 71:109:@37945.4]
  wire [11:0] _T_81937; // @[Modules.scala 71:109:@37947.4]
  wire [10:0] _T_81938; // @[Modules.scala 71:109:@37948.4]
  wire [10:0] buffer_15_732; // @[Modules.scala 71:109:@37949.4]
  wire [11:0] _T_81940; // @[Modules.scala 71:109:@37951.4]
  wire [10:0] _T_81941; // @[Modules.scala 71:109:@37952.4]
  wire [10:0] buffer_15_733; // @[Modules.scala 71:109:@37953.4]
  wire [11:0] _T_81943; // @[Modules.scala 71:109:@37955.4]
  wire [10:0] _T_81944; // @[Modules.scala 71:109:@37956.4]
  wire [10:0] buffer_15_734; // @[Modules.scala 71:109:@37957.4]
  wire [11:0] _T_81946; // @[Modules.scala 78:156:@37960.4]
  wire [10:0] _T_81947; // @[Modules.scala 78:156:@37961.4]
  wire [10:0] buffer_15_736; // @[Modules.scala 78:156:@37962.4]
  wire [11:0] _T_81949; // @[Modules.scala 78:156:@37964.4]
  wire [10:0] _T_81950; // @[Modules.scala 78:156:@37965.4]
  wire [10:0] buffer_15_737; // @[Modules.scala 78:156:@37966.4]
  wire [11:0] _T_81952; // @[Modules.scala 78:156:@37968.4]
  wire [10:0] _T_81953; // @[Modules.scala 78:156:@37969.4]
  wire [10:0] buffer_15_738; // @[Modules.scala 78:156:@37970.4]
  wire [11:0] _T_81955; // @[Modules.scala 78:156:@37972.4]
  wire [10:0] _T_81956; // @[Modules.scala 78:156:@37973.4]
  wire [10:0] buffer_15_739; // @[Modules.scala 78:156:@37974.4]
  wire [11:0] _T_81958; // @[Modules.scala 78:156:@37976.4]
  wire [10:0] _T_81959; // @[Modules.scala 78:156:@37977.4]
  wire [10:0] buffer_15_740; // @[Modules.scala 78:156:@37978.4]
  wire [11:0] _T_81961; // @[Modules.scala 78:156:@37980.4]
  wire [10:0] _T_81962; // @[Modules.scala 78:156:@37981.4]
  wire [10:0] buffer_15_741; // @[Modules.scala 78:156:@37982.4]
  wire [11:0] _T_81964; // @[Modules.scala 78:156:@37984.4]
  wire [10:0] _T_81965; // @[Modules.scala 78:156:@37985.4]
  wire [10:0] buffer_15_742; // @[Modules.scala 78:156:@37986.4]
  wire [11:0] _T_81967; // @[Modules.scala 78:156:@37988.4]
  wire [10:0] _T_81968; // @[Modules.scala 78:156:@37989.4]
  wire [10:0] buffer_15_743; // @[Modules.scala 78:156:@37990.4]
  wire [11:0] _T_81970; // @[Modules.scala 78:156:@37992.4]
  wire [10:0] _T_81971; // @[Modules.scala 78:156:@37993.4]
  wire [10:0] buffer_15_744; // @[Modules.scala 78:156:@37994.4]
  wire [11:0] _T_81973; // @[Modules.scala 78:156:@37996.4]
  wire [10:0] _T_81974; // @[Modules.scala 78:156:@37997.4]
  wire [10:0] buffer_15_745; // @[Modules.scala 78:156:@37998.4]
  wire [11:0] _T_81976; // @[Modules.scala 78:156:@38000.4]
  wire [10:0] _T_81977; // @[Modules.scala 78:156:@38001.4]
  wire [10:0] buffer_15_746; // @[Modules.scala 78:156:@38002.4]
  wire [11:0] _T_81979; // @[Modules.scala 78:156:@38004.4]
  wire [10:0] _T_81980; // @[Modules.scala 78:156:@38005.4]
  wire [10:0] buffer_15_747; // @[Modules.scala 78:156:@38006.4]
  wire [11:0] _T_81982; // @[Modules.scala 78:156:@38008.4]
  wire [10:0] _T_81983; // @[Modules.scala 78:156:@38009.4]
  wire [10:0] buffer_15_748; // @[Modules.scala 78:156:@38010.4]
  wire [11:0] _T_81985; // @[Modules.scala 78:156:@38012.4]
  wire [10:0] _T_81986; // @[Modules.scala 78:156:@38013.4]
  wire [10:0] buffer_15_749; // @[Modules.scala 78:156:@38014.4]
  wire [11:0] _T_81988; // @[Modules.scala 78:156:@38016.4]
  wire [10:0] _T_81989; // @[Modules.scala 78:156:@38017.4]
  wire [10:0] buffer_15_750; // @[Modules.scala 78:156:@38018.4]
  wire [11:0] _T_81991; // @[Modules.scala 78:156:@38020.4]
  wire [10:0] _T_81992; // @[Modules.scala 78:156:@38021.4]
  wire [10:0] buffer_15_751; // @[Modules.scala 78:156:@38022.4]
  wire [11:0] _T_81994; // @[Modules.scala 78:156:@38024.4]
  wire [10:0] _T_81995; // @[Modules.scala 78:156:@38025.4]
  wire [10:0] buffer_15_752; // @[Modules.scala 78:156:@38026.4]
  wire [11:0] _T_81997; // @[Modules.scala 78:156:@38028.4]
  wire [10:0] _T_81998; // @[Modules.scala 78:156:@38029.4]
  wire [10:0] buffer_15_753; // @[Modules.scala 78:156:@38030.4]
  wire [11:0] _T_82000; // @[Modules.scala 78:156:@38032.4]
  wire [10:0] _T_82001; // @[Modules.scala 78:156:@38033.4]
  wire [10:0] buffer_15_754; // @[Modules.scala 78:156:@38034.4]
  wire [11:0] _T_82003; // @[Modules.scala 78:156:@38036.4]
  wire [10:0] _T_82004; // @[Modules.scala 78:156:@38037.4]
  wire [10:0] buffer_15_755; // @[Modules.scala 78:156:@38038.4]
  wire [11:0] _T_82006; // @[Modules.scala 78:156:@38040.4]
  wire [10:0] _T_82007; // @[Modules.scala 78:156:@38041.4]
  wire [10:0] buffer_15_756; // @[Modules.scala 78:156:@38042.4]
  wire [11:0] _T_82009; // @[Modules.scala 78:156:@38044.4]
  wire [10:0] _T_82010; // @[Modules.scala 78:156:@38045.4]
  wire [10:0] buffer_15_757; // @[Modules.scala 78:156:@38046.4]
  wire [11:0] _T_82012; // @[Modules.scala 78:156:@38048.4]
  wire [10:0] _T_82013; // @[Modules.scala 78:156:@38049.4]
  wire [10:0] buffer_15_758; // @[Modules.scala 78:156:@38050.4]
  wire [11:0] _T_82015; // @[Modules.scala 78:156:@38052.4]
  wire [10:0] _T_82016; // @[Modules.scala 78:156:@38053.4]
  wire [10:0] buffer_15_759; // @[Modules.scala 78:156:@38054.4]
  wire [11:0] _T_82018; // @[Modules.scala 78:156:@38056.4]
  wire [10:0] _T_82019; // @[Modules.scala 78:156:@38057.4]
  wire [10:0] buffer_15_760; // @[Modules.scala 78:156:@38058.4]
  wire [11:0] _T_82021; // @[Modules.scala 78:156:@38060.4]
  wire [10:0] _T_82022; // @[Modules.scala 78:156:@38061.4]
  wire [10:0] buffer_15_761; // @[Modules.scala 78:156:@38062.4]
  wire [11:0] _T_82024; // @[Modules.scala 78:156:@38064.4]
  wire [10:0] _T_82025; // @[Modules.scala 78:156:@38065.4]
  wire [10:0] buffer_15_762; // @[Modules.scala 78:156:@38066.4]
  wire [11:0] _T_82027; // @[Modules.scala 78:156:@38068.4]
  wire [10:0] _T_82028; // @[Modules.scala 78:156:@38069.4]
  wire [10:0] buffer_15_763; // @[Modules.scala 78:156:@38070.4]
  wire [11:0] _T_82030; // @[Modules.scala 78:156:@38072.4]
  wire [10:0] _T_82031; // @[Modules.scala 78:156:@38073.4]
  wire [10:0] buffer_15_764; // @[Modules.scala 78:156:@38074.4]
  wire [11:0] _T_82033; // @[Modules.scala 78:156:@38076.4]
  wire [10:0] _T_82034; // @[Modules.scala 78:156:@38077.4]
  wire [10:0] buffer_15_765; // @[Modules.scala 78:156:@38078.4]
  wire [11:0] _T_82036; // @[Modules.scala 78:156:@38080.4]
  wire [10:0] _T_82037; // @[Modules.scala 78:156:@38081.4]
  wire [10:0] buffer_15_766; // @[Modules.scala 78:156:@38082.4]
  wire [11:0] _T_82039; // @[Modules.scala 78:156:@38084.4]
  wire [10:0] _T_82040; // @[Modules.scala 78:156:@38085.4]
  wire [10:0] buffer_15_767; // @[Modules.scala 78:156:@38086.4]
  wire [11:0] _T_82042; // @[Modules.scala 78:156:@38088.4]
  wire [10:0] _T_82043; // @[Modules.scala 78:156:@38089.4]
  wire [10:0] buffer_15_768; // @[Modules.scala 78:156:@38090.4]
  wire [11:0] _T_82045; // @[Modules.scala 78:156:@38092.4]
  wire [10:0] _T_82046; // @[Modules.scala 78:156:@38093.4]
  wire [10:0] buffer_15_769; // @[Modules.scala 78:156:@38094.4]
  wire [11:0] _T_82048; // @[Modules.scala 78:156:@38096.4]
  wire [10:0] _T_82049; // @[Modules.scala 78:156:@38097.4]
  wire [10:0] buffer_15_770; // @[Modules.scala 78:156:@38098.4]
  wire [11:0] _T_82051; // @[Modules.scala 78:156:@38100.4]
  wire [10:0] _T_82052; // @[Modules.scala 78:156:@38101.4]
  wire [10:0] buffer_15_771; // @[Modules.scala 78:156:@38102.4]
  wire [11:0] _T_82054; // @[Modules.scala 78:156:@38104.4]
  wire [10:0] _T_82055; // @[Modules.scala 78:156:@38105.4]
  wire [10:0] buffer_15_772; // @[Modules.scala 78:156:@38106.4]
  wire [11:0] _T_82057; // @[Modules.scala 78:156:@38108.4]
  wire [10:0] _T_82058; // @[Modules.scala 78:156:@38109.4]
  wire [10:0] buffer_15_773; // @[Modules.scala 78:156:@38110.4]
  wire [11:0] _T_82060; // @[Modules.scala 78:156:@38112.4]
  wire [10:0] _T_82061; // @[Modules.scala 78:156:@38113.4]
  wire [10:0] buffer_15_774; // @[Modules.scala 78:156:@38114.4]
  wire [11:0] _T_82063; // @[Modules.scala 78:156:@38116.4]
  wire [10:0] _T_82064; // @[Modules.scala 78:156:@38117.4]
  wire [10:0] buffer_15_775; // @[Modules.scala 78:156:@38118.4]
  wire [11:0] _T_82066; // @[Modules.scala 78:156:@38120.4]
  wire [10:0] _T_82067; // @[Modules.scala 78:156:@38121.4]
  wire [10:0] buffer_15_776; // @[Modules.scala 78:156:@38122.4]
  wire [11:0] _T_82069; // @[Modules.scala 78:156:@38124.4]
  wire [10:0] _T_82070; // @[Modules.scala 78:156:@38125.4]
  wire [10:0] buffer_15_777; // @[Modules.scala 78:156:@38126.4]
  wire [11:0] _T_82072; // @[Modules.scala 78:156:@38128.4]
  wire [10:0] _T_82073; // @[Modules.scala 78:156:@38129.4]
  wire [10:0] buffer_15_778; // @[Modules.scala 78:156:@38130.4]
  wire [11:0] _T_82075; // @[Modules.scala 78:156:@38132.4]
  wire [10:0] _T_82076; // @[Modules.scala 78:156:@38133.4]
  wire [10:0] buffer_15_779; // @[Modules.scala 78:156:@38134.4]
  wire [11:0] _T_82078; // @[Modules.scala 78:156:@38136.4]
  wire [10:0] _T_82079; // @[Modules.scala 78:156:@38137.4]
  wire [10:0] buffer_15_780; // @[Modules.scala 78:156:@38138.4]
  wire [11:0] _T_82081; // @[Modules.scala 78:156:@38140.4]
  wire [10:0] _T_82082; // @[Modules.scala 78:156:@38141.4]
  wire [10:0] buffer_15_781; // @[Modules.scala 78:156:@38142.4]
  wire [11:0] _T_82084; // @[Modules.scala 78:156:@38144.4]
  wire [10:0] _T_82085; // @[Modules.scala 78:156:@38145.4]
  wire [10:0] buffer_15_782; // @[Modules.scala 78:156:@38146.4]
  wire [11:0] _T_82087; // @[Modules.scala 78:156:@38148.4]
  wire [10:0] _T_82088; // @[Modules.scala 78:156:@38149.4]
  wire [10:0] buffer_15_783; // @[Modules.scala 78:156:@38150.4]
  assign _T_54270 = $signed(io_in_16) + $signed(io_in_17); // @[Modules.scala 37:46:@17.4]
  assign _T_54271 = _T_54270[4:0]; // @[Modules.scala 37:46:@18.4]
  assign _T_54272 = $signed(_T_54271); // @[Modules.scala 37:46:@19.4]
  assign _T_54274 = $signed(io_in_20) + $signed(io_in_21); // @[Modules.scala 37:46:@22.4]
  assign _T_54275 = _T_54274[4:0]; // @[Modules.scala 37:46:@23.4]
  assign _T_54276 = $signed(_T_54275); // @[Modules.scala 37:46:@24.4]
  assign _T_54278 = $signed(io_in_32) + $signed(io_in_33); // @[Modules.scala 37:46:@31.4]
  assign _T_54279 = _T_54278[4:0]; // @[Modules.scala 37:46:@32.4]
  assign _T_54280 = $signed(_T_54279); // @[Modules.scala 37:46:@33.4]
  assign _T_54290 = $signed(io_in_52) + $signed(io_in_53); // @[Modules.scala 37:46:@44.4]
  assign _T_54291 = _T_54290[4:0]; // @[Modules.scala 37:46:@45.4]
  assign _T_54292 = $signed(_T_54291); // @[Modules.scala 37:46:@46.4]
  assign _T_54300 = $signed(io_in_78) + $signed(io_in_79); // @[Modules.scala 37:46:@60.4]
  assign _T_54301 = _T_54300[4:0]; // @[Modules.scala 37:46:@61.4]
  assign _T_54302 = $signed(_T_54301); // @[Modules.scala 37:46:@62.4]
  assign _T_54305 = $signed(io_in_88) + $signed(io_in_89); // @[Modules.scala 37:46:@68.4]
  assign _T_54306 = _T_54305[4:0]; // @[Modules.scala 37:46:@69.4]
  assign _T_54307 = $signed(_T_54306); // @[Modules.scala 37:46:@70.4]
  assign _T_54308 = $signed(io_in_90) + $signed(io_in_91); // @[Modules.scala 37:46:@72.4]
  assign _T_54309 = _T_54308[4:0]; // @[Modules.scala 37:46:@73.4]
  assign _T_54310 = $signed(_T_54309); // @[Modules.scala 37:46:@74.4]
  assign _T_54311 = $signed(io_in_94) + $signed(io_in_95); // @[Modules.scala 37:46:@77.4]
  assign _T_54312 = _T_54311[4:0]; // @[Modules.scala 37:46:@78.4]
  assign _T_54313 = $signed(_T_54312); // @[Modules.scala 37:46:@79.4]
  assign _T_54314 = $signed(io_in_98) + $signed(io_in_99); // @[Modules.scala 37:46:@82.4]
  assign _T_54315 = _T_54314[4:0]; // @[Modules.scala 37:46:@83.4]
  assign _T_54316 = $signed(_T_54315); // @[Modules.scala 37:46:@84.4]
  assign _T_54317 = $signed(io_in_100) + $signed(io_in_101); // @[Modules.scala 37:46:@86.4]
  assign _T_54318 = _T_54317[4:0]; // @[Modules.scala 37:46:@87.4]
  assign _T_54319 = $signed(_T_54318); // @[Modules.scala 37:46:@88.4]
  assign _T_54320 = $signed(io_in_102) + $signed(io_in_103); // @[Modules.scala 37:46:@90.4]
  assign _T_54321 = _T_54320[4:0]; // @[Modules.scala 37:46:@91.4]
  assign _T_54322 = $signed(_T_54321); // @[Modules.scala 37:46:@92.4]
  assign _T_54323 = $signed(io_in_104) + $signed(io_in_105); // @[Modules.scala 37:46:@94.4]
  assign _T_54324 = _T_54323[4:0]; // @[Modules.scala 37:46:@95.4]
  assign _T_54325 = $signed(_T_54324); // @[Modules.scala 37:46:@96.4]
  assign _T_54326 = $signed(io_in_106) + $signed(io_in_107); // @[Modules.scala 37:46:@98.4]
  assign _T_54327 = _T_54326[4:0]; // @[Modules.scala 37:46:@99.4]
  assign _T_54328 = $signed(_T_54327); // @[Modules.scala 37:46:@100.4]
  assign _T_54329 = $signed(io_in_110) + $signed(io_in_111); // @[Modules.scala 37:46:@103.4]
  assign _T_54330 = _T_54329[4:0]; // @[Modules.scala 37:46:@104.4]
  assign _T_54331 = $signed(_T_54330); // @[Modules.scala 37:46:@105.4]
  assign _T_54333 = $signed(io_in_118) + $signed(io_in_119); // @[Modules.scala 37:46:@110.4]
  assign _T_54334 = _T_54333[4:0]; // @[Modules.scala 37:46:@111.4]
  assign _T_54335 = $signed(_T_54334); // @[Modules.scala 37:46:@112.4]
  assign _T_54340 = $signed(io_in_132) + $signed(io_in_133); // @[Modules.scala 37:46:@120.4]
  assign _T_54341 = _T_54340[4:0]; // @[Modules.scala 37:46:@121.4]
  assign _T_54342 = $signed(_T_54341); // @[Modules.scala 37:46:@122.4]
  assign _T_54343 = $signed(io_in_134) + $signed(io_in_135); // @[Modules.scala 37:46:@124.4]
  assign _T_54344 = _T_54343[4:0]; // @[Modules.scala 37:46:@125.4]
  assign _T_54345 = $signed(_T_54344); // @[Modules.scala 37:46:@126.4]
  assign _T_54347 = $signed(io_in_140) + $signed(io_in_141); // @[Modules.scala 37:46:@130.4]
  assign _T_54348 = _T_54347[4:0]; // @[Modules.scala 37:46:@131.4]
  assign _T_54349 = $signed(_T_54348); // @[Modules.scala 37:46:@132.4]
  assign _T_54351 = $signed(io_in_146) + $signed(io_in_147); // @[Modules.scala 37:46:@136.4]
  assign _T_54352 = _T_54351[4:0]; // @[Modules.scala 37:46:@137.4]
  assign _T_54353 = $signed(_T_54352); // @[Modules.scala 37:46:@138.4]
  assign _T_54354 = $signed(io_in_148) + $signed(io_in_149); // @[Modules.scala 37:46:@140.4]
  assign _T_54355 = _T_54354[4:0]; // @[Modules.scala 37:46:@141.4]
  assign _T_54356 = $signed(_T_54355); // @[Modules.scala 37:46:@142.4]
  assign _T_54363 = $signed(io_in_162) + $signed(io_in_163); // @[Modules.scala 37:46:@150.4]
  assign _T_54364 = _T_54363[4:0]; // @[Modules.scala 37:46:@151.4]
  assign _T_54365 = $signed(_T_54364); // @[Modules.scala 37:46:@152.4]
  assign _T_54374 = $signed(io_in_186) + $signed(io_in_187); // @[Modules.scala 37:46:@165.4]
  assign _T_54375 = _T_54374[4:0]; // @[Modules.scala 37:46:@166.4]
  assign _T_54376 = $signed(_T_54375); // @[Modules.scala 37:46:@167.4]
  assign _T_54383 = $signed(io_in_210) + $signed(io_in_211); // @[Modules.scala 37:46:@180.4]
  assign _T_54384 = _T_54383[4:0]; // @[Modules.scala 37:46:@181.4]
  assign _T_54385 = $signed(_T_54384); // @[Modules.scala 37:46:@182.4]
  assign _T_54433 = $signed(io_in_316) + $signed(io_in_317); // @[Modules.scala 37:46:@236.4]
  assign _T_54434 = _T_54433[4:0]; // @[Modules.scala 37:46:@237.4]
  assign _T_54435 = $signed(_T_54434); // @[Modules.scala 37:46:@238.4]
  assign _T_54436 = $signed(io_in_318) + $signed(io_in_319); // @[Modules.scala 37:46:@240.4]
  assign _T_54437 = _T_54436[4:0]; // @[Modules.scala 37:46:@241.4]
  assign _T_54438 = $signed(_T_54437); // @[Modules.scala 37:46:@242.4]
  assign _T_54442 = $signed(io_in_328) + $signed(io_in_329); // @[Modules.scala 37:46:@248.4]
  assign _T_54443 = _T_54442[4:0]; // @[Modules.scala 37:46:@249.4]
  assign _T_54444 = $signed(_T_54443); // @[Modules.scala 37:46:@250.4]
  assign _T_54448 = $signed(io_in_342) + $signed(io_in_343); // @[Modules.scala 37:46:@258.4]
  assign _T_54449 = _T_54448[4:0]; // @[Modules.scala 37:46:@259.4]
  assign _T_54450 = $signed(_T_54449); // @[Modules.scala 37:46:@260.4]
  assign _T_54451 = $signed(io_in_344) + $signed(io_in_345); // @[Modules.scala 37:46:@262.4]
  assign _T_54452 = _T_54451[4:0]; // @[Modules.scala 37:46:@263.4]
  assign _T_54453 = $signed(_T_54452); // @[Modules.scala 37:46:@264.4]
  assign _T_54454 = $signed(io_in_346) + $signed(io_in_347); // @[Modules.scala 37:46:@266.4]
  assign _T_54455 = _T_54454[4:0]; // @[Modules.scala 37:46:@267.4]
  assign _T_54456 = $signed(_T_54455); // @[Modules.scala 37:46:@268.4]
  assign _T_54457 = $signed(io_in_348) + $signed(io_in_349); // @[Modules.scala 37:46:@270.4]
  assign _T_54458 = _T_54457[4:0]; // @[Modules.scala 37:46:@271.4]
  assign _T_54459 = $signed(_T_54458); // @[Modules.scala 37:46:@272.4]
  assign _T_54460 = $signed(io_in_350) + $signed(io_in_351); // @[Modules.scala 37:46:@274.4]
  assign _T_54461 = _T_54460[4:0]; // @[Modules.scala 37:46:@275.4]
  assign _T_54462 = $signed(_T_54461); // @[Modules.scala 37:46:@276.4]
  assign _T_54463 = $signed(io_in_352) + $signed(io_in_353); // @[Modules.scala 37:46:@278.4]
  assign _T_54464 = _T_54463[4:0]; // @[Modules.scala 37:46:@279.4]
  assign _T_54465 = $signed(_T_54464); // @[Modules.scala 37:46:@280.4]
  assign _T_54466 = $signed(io_in_354) + $signed(io_in_355); // @[Modules.scala 37:46:@282.4]
  assign _T_54467 = _T_54466[4:0]; // @[Modules.scala 37:46:@283.4]
  assign _T_54468 = $signed(_T_54467); // @[Modules.scala 37:46:@284.4]
  assign _T_54469 = $signed(io_in_356) + $signed(io_in_357); // @[Modules.scala 37:46:@286.4]
  assign _T_54470 = _T_54469[4:0]; // @[Modules.scala 37:46:@287.4]
  assign _T_54471 = $signed(_T_54470); // @[Modules.scala 37:46:@288.4]
  assign _T_54472 = $signed(io_in_358) + $signed(io_in_359); // @[Modules.scala 37:46:@290.4]
  assign _T_54473 = _T_54472[4:0]; // @[Modules.scala 37:46:@291.4]
  assign _T_54474 = $signed(_T_54473); // @[Modules.scala 37:46:@292.4]
  assign _T_54478 = $signed(io_in_368) + $signed(io_in_369); // @[Modules.scala 37:46:@298.4]
  assign _T_54479 = _T_54478[4:0]; // @[Modules.scala 37:46:@299.4]
  assign _T_54480 = $signed(_T_54479); // @[Modules.scala 37:46:@300.4]
  assign _T_54481 = $signed(io_in_370) + $signed(io_in_371); // @[Modules.scala 37:46:@302.4]
  assign _T_54482 = _T_54481[4:0]; // @[Modules.scala 37:46:@303.4]
  assign _T_54483 = $signed(_T_54482); // @[Modules.scala 37:46:@304.4]
  assign _T_54484 = $signed(io_in_372) + $signed(io_in_373); // @[Modules.scala 37:46:@306.4]
  assign _T_54485 = _T_54484[4:0]; // @[Modules.scala 37:46:@307.4]
  assign _T_54486 = $signed(_T_54485); // @[Modules.scala 37:46:@308.4]
  assign _T_54487 = $signed(io_in_374) + $signed(io_in_375); // @[Modules.scala 37:46:@310.4]
  assign _T_54488 = _T_54487[4:0]; // @[Modules.scala 37:46:@311.4]
  assign _T_54489 = $signed(_T_54488); // @[Modules.scala 37:46:@312.4]
  assign _T_54490 = $signed(io_in_376) + $signed(io_in_377); // @[Modules.scala 37:46:@314.4]
  assign _T_54491 = _T_54490[4:0]; // @[Modules.scala 37:46:@315.4]
  assign _T_54492 = $signed(_T_54491); // @[Modules.scala 37:46:@316.4]
  assign _T_54493 = $signed(io_in_378) + $signed(io_in_379); // @[Modules.scala 37:46:@318.4]
  assign _T_54494 = _T_54493[4:0]; // @[Modules.scala 37:46:@319.4]
  assign _T_54495 = $signed(_T_54494); // @[Modules.scala 37:46:@320.4]
  assign _T_54496 = $signed(io_in_380) + $signed(io_in_381); // @[Modules.scala 37:46:@322.4]
  assign _T_54497 = _T_54496[4:0]; // @[Modules.scala 37:46:@323.4]
  assign _T_54498 = $signed(_T_54497); // @[Modules.scala 37:46:@324.4]
  assign _T_54499 = $signed(io_in_382) + $signed(io_in_383); // @[Modules.scala 37:46:@326.4]
  assign _T_54500 = _T_54499[4:0]; // @[Modules.scala 37:46:@327.4]
  assign _T_54501 = $signed(_T_54500); // @[Modules.scala 37:46:@328.4]
  assign _T_54502 = $signed(io_in_386) + $signed(io_in_387); // @[Modules.scala 37:46:@331.4]
  assign _T_54503 = _T_54502[4:0]; // @[Modules.scala 37:46:@332.4]
  assign _T_54504 = $signed(_T_54503); // @[Modules.scala 37:46:@333.4]
  assign _T_54507 = $signed(io_in_396) + $signed(io_in_397); // @[Modules.scala 37:46:@339.4]
  assign _T_54508 = _T_54507[4:0]; // @[Modules.scala 37:46:@340.4]
  assign _T_54509 = $signed(_T_54508); // @[Modules.scala 37:46:@341.4]
  assign _T_54510 = $signed(io_in_398) + $signed(io_in_399); // @[Modules.scala 37:46:@343.4]
  assign _T_54511 = _T_54510[4:0]; // @[Modules.scala 37:46:@344.4]
  assign _T_54512 = $signed(_T_54511); // @[Modules.scala 37:46:@345.4]
  assign _T_54513 = $signed(io_in_400) + $signed(io_in_401); // @[Modules.scala 37:46:@347.4]
  assign _T_54514 = _T_54513[4:0]; // @[Modules.scala 37:46:@348.4]
  assign _T_54515 = $signed(_T_54514); // @[Modules.scala 37:46:@349.4]
  assign _T_54516 = $signed(io_in_402) + $signed(io_in_403); // @[Modules.scala 37:46:@351.4]
  assign _T_54517 = _T_54516[4:0]; // @[Modules.scala 37:46:@352.4]
  assign _T_54518 = $signed(_T_54517); // @[Modules.scala 37:46:@353.4]
  assign _T_54519 = $signed(io_in_404) + $signed(io_in_405); // @[Modules.scala 37:46:@355.4]
  assign _T_54520 = _T_54519[4:0]; // @[Modules.scala 37:46:@356.4]
  assign _T_54521 = $signed(_T_54520); // @[Modules.scala 37:46:@357.4]
  assign _T_54522 = $signed(io_in_406) + $signed(io_in_407); // @[Modules.scala 37:46:@359.4]
  assign _T_54523 = _T_54522[4:0]; // @[Modules.scala 37:46:@360.4]
  assign _T_54524 = $signed(_T_54523); // @[Modules.scala 37:46:@361.4]
  assign _T_54525 = $signed(io_in_408) + $signed(io_in_409); // @[Modules.scala 37:46:@363.4]
  assign _T_54526 = _T_54525[4:0]; // @[Modules.scala 37:46:@364.4]
  assign _T_54527 = $signed(_T_54526); // @[Modules.scala 37:46:@365.4]
  assign _T_54528 = $signed(io_in_410) + $signed(io_in_411); // @[Modules.scala 37:46:@367.4]
  assign _T_54529 = _T_54528[4:0]; // @[Modules.scala 37:46:@368.4]
  assign _T_54530 = $signed(_T_54529); // @[Modules.scala 37:46:@369.4]
  assign _T_54531 = $signed(io_in_412) + $signed(io_in_413); // @[Modules.scala 37:46:@371.4]
  assign _T_54532 = _T_54531[4:0]; // @[Modules.scala 37:46:@372.4]
  assign _T_54533 = $signed(_T_54532); // @[Modules.scala 37:46:@373.4]
  assign _T_54534 = $signed(io_in_414) + $signed(io_in_415); // @[Modules.scala 37:46:@375.4]
  assign _T_54535 = _T_54534[4:0]; // @[Modules.scala 37:46:@376.4]
  assign _T_54536 = $signed(_T_54535); // @[Modules.scala 37:46:@377.4]
  assign _T_54538 = $signed(io_in_426) + $signed(io_in_427); // @[Modules.scala 37:46:@384.4]
  assign _T_54539 = _T_54538[4:0]; // @[Modules.scala 37:46:@385.4]
  assign _T_54540 = $signed(_T_54539); // @[Modules.scala 37:46:@386.4]
  assign _T_54541 = $signed(io_in_428) + $signed(io_in_429); // @[Modules.scala 37:46:@388.4]
  assign _T_54542 = _T_54541[4:0]; // @[Modules.scala 37:46:@389.4]
  assign _T_54543 = $signed(_T_54542); // @[Modules.scala 37:46:@390.4]
  assign _T_54544 = $signed(io_in_430) + $signed(io_in_431); // @[Modules.scala 37:46:@392.4]
  assign _T_54545 = _T_54544[4:0]; // @[Modules.scala 37:46:@393.4]
  assign _T_54546 = $signed(_T_54545); // @[Modules.scala 37:46:@394.4]
  assign _T_54547 = $signed(io_in_432) + $signed(io_in_433); // @[Modules.scala 37:46:@396.4]
  assign _T_54548 = _T_54547[4:0]; // @[Modules.scala 37:46:@397.4]
  assign _T_54549 = $signed(_T_54548); // @[Modules.scala 37:46:@398.4]
  assign _T_54550 = $signed(io_in_434) + $signed(io_in_435); // @[Modules.scala 37:46:@400.4]
  assign _T_54551 = _T_54550[4:0]; // @[Modules.scala 37:46:@401.4]
  assign _T_54552 = $signed(_T_54551); // @[Modules.scala 37:46:@402.4]
  assign _T_54553 = $signed(io_in_436) + $signed(io_in_437); // @[Modules.scala 37:46:@404.4]
  assign _T_54554 = _T_54553[4:0]; // @[Modules.scala 37:46:@405.4]
  assign _T_54555 = $signed(_T_54554); // @[Modules.scala 37:46:@406.4]
  assign _T_54558 = $signed(io_in_448) + $signed(io_in_449); // @[Modules.scala 37:46:@413.4]
  assign _T_54559 = _T_54558[4:0]; // @[Modules.scala 37:46:@414.4]
  assign _T_54560 = $signed(_T_54559); // @[Modules.scala 37:46:@415.4]
  assign _T_54562 = $signed(io_in_454) + $signed(io_in_455); // @[Modules.scala 37:46:@419.4]
  assign _T_54563 = _T_54562[4:0]; // @[Modules.scala 37:46:@420.4]
  assign _T_54564 = $signed(_T_54563); // @[Modules.scala 37:46:@421.4]
  assign _T_54565 = $signed(io_in_456) + $signed(io_in_457); // @[Modules.scala 37:46:@423.4]
  assign _T_54566 = _T_54565[4:0]; // @[Modules.scala 37:46:@424.4]
  assign _T_54567 = $signed(_T_54566); // @[Modules.scala 37:46:@425.4]
  assign _T_54568 = $signed(io_in_458) + $signed(io_in_459); // @[Modules.scala 37:46:@427.4]
  assign _T_54569 = _T_54568[4:0]; // @[Modules.scala 37:46:@428.4]
  assign _T_54570 = $signed(_T_54569); // @[Modules.scala 37:46:@429.4]
  assign _T_54571 = $signed(io_in_462) + $signed(io_in_463); // @[Modules.scala 37:46:@432.4]
  assign _T_54572 = _T_54571[4:0]; // @[Modules.scala 37:46:@433.4]
  assign _T_54573 = $signed(_T_54572); // @[Modules.scala 37:46:@434.4]
  assign _T_54574 = $signed(io_in_464) + $signed(io_in_465); // @[Modules.scala 37:46:@436.4]
  assign _T_54575 = _T_54574[4:0]; // @[Modules.scala 37:46:@437.4]
  assign _T_54576 = $signed(_T_54575); // @[Modules.scala 37:46:@438.4]
  assign _T_54577 = $signed(io_in_466) + $signed(io_in_467); // @[Modules.scala 37:46:@440.4]
  assign _T_54578 = _T_54577[4:0]; // @[Modules.scala 37:46:@441.4]
  assign _T_54579 = $signed(_T_54578); // @[Modules.scala 37:46:@442.4]
  assign _T_54585 = $signed(io_in_482) + $signed(io_in_483); // @[Modules.scala 37:46:@451.4]
  assign _T_54586 = _T_54585[4:0]; // @[Modules.scala 37:46:@452.4]
  assign _T_54587 = $signed(_T_54586); // @[Modules.scala 37:46:@453.4]
  assign _T_54588 = $signed(io_in_484) + $signed(io_in_485); // @[Modules.scala 37:46:@455.4]
  assign _T_54589 = _T_54588[4:0]; // @[Modules.scala 37:46:@456.4]
  assign _T_54590 = $signed(_T_54589); // @[Modules.scala 37:46:@457.4]
  assign _T_54591 = $signed(io_in_486) + $signed(io_in_487); // @[Modules.scala 37:46:@459.4]
  assign _T_54592 = _T_54591[4:0]; // @[Modules.scala 37:46:@460.4]
  assign _T_54593 = $signed(_T_54592); // @[Modules.scala 37:46:@461.4]
  assign _T_54594 = $signed(io_in_490) + $signed(io_in_491); // @[Modules.scala 37:46:@464.4]
  assign _T_54595 = _T_54594[4:0]; // @[Modules.scala 37:46:@465.4]
  assign _T_54596 = $signed(_T_54595); // @[Modules.scala 37:46:@466.4]
  assign _T_54598 = $signed(io_in_498) + $signed(io_in_499); // @[Modules.scala 37:46:@471.4]
  assign _T_54599 = _T_54598[4:0]; // @[Modules.scala 37:46:@472.4]
  assign _T_54600 = $signed(_T_54599); // @[Modules.scala 37:46:@473.4]
  assign _T_54606 = $signed(io_in_512) + $signed(io_in_513); // @[Modules.scala 37:46:@481.4]
  assign _T_54607 = _T_54606[4:0]; // @[Modules.scala 37:46:@482.4]
  assign _T_54608 = $signed(_T_54607); // @[Modules.scala 37:46:@483.4]
  assign _T_54609 = $signed(io_in_514) + $signed(io_in_515); // @[Modules.scala 37:46:@485.4]
  assign _T_54610 = _T_54609[4:0]; // @[Modules.scala 37:46:@486.4]
  assign _T_54611 = $signed(_T_54610); // @[Modules.scala 37:46:@487.4]
  assign _T_54612 = $signed(io_in_518) + $signed(io_in_519); // @[Modules.scala 37:46:@490.4]
  assign _T_54613 = _T_54612[4:0]; // @[Modules.scala 37:46:@491.4]
  assign _T_54614 = $signed(_T_54613); // @[Modules.scala 37:46:@492.4]
  assign _T_54615 = $signed(io_in_526) + $signed(io_in_527); // @[Modules.scala 37:46:@497.4]
  assign _T_54616 = _T_54615[4:0]; // @[Modules.scala 37:46:@498.4]
  assign _T_54617 = $signed(_T_54616); // @[Modules.scala 37:46:@499.4]
  assign _T_54618 = $signed(io_in_528) + $signed(io_in_529); // @[Modules.scala 37:46:@501.4]
  assign _T_54619 = _T_54618[4:0]; // @[Modules.scala 37:46:@502.4]
  assign _T_54620 = $signed(_T_54619); // @[Modules.scala 37:46:@503.4]
  assign _T_54634 = $signed(io_in_576) + $signed(io_in_577); // @[Modules.scala 37:46:@528.4]
  assign _T_54635 = _T_54634[4:0]; // @[Modules.scala 37:46:@529.4]
  assign _T_54636 = $signed(_T_54635); // @[Modules.scala 37:46:@530.4]
  assign _T_54638 = $signed(io_in_584) + $signed(io_in_585); // @[Modules.scala 37:46:@535.4]
  assign _T_54639 = _T_54638[4:0]; // @[Modules.scala 37:46:@536.4]
  assign _T_54640 = $signed(_T_54639); // @[Modules.scala 37:46:@537.4]
  assign _T_54646 = $signed(io_in_600) + $signed(io_in_601); // @[Modules.scala 37:46:@546.4]
  assign _T_54647 = _T_54646[4:0]; // @[Modules.scala 37:46:@547.4]
  assign _T_54648 = $signed(_T_54647); // @[Modules.scala 37:46:@548.4]
  assign _T_54649 = $signed(io_in_604) + $signed(io_in_605); // @[Modules.scala 37:46:@551.4]
  assign _T_54650 = _T_54649[4:0]; // @[Modules.scala 37:46:@552.4]
  assign _T_54651 = $signed(_T_54650); // @[Modules.scala 37:46:@553.4]
  assign _T_54652 = $signed(io_in_606) + $signed(io_in_607); // @[Modules.scala 37:46:@555.4]
  assign _T_54653 = _T_54652[4:0]; // @[Modules.scala 37:46:@556.4]
  assign _T_54654 = $signed(_T_54653); // @[Modules.scala 37:46:@557.4]
  assign _T_54657 = $signed(io_in_612) + $signed(io_in_613); // @[Modules.scala 37:46:@561.4]
  assign _T_54658 = _T_54657[4:0]; // @[Modules.scala 37:46:@562.4]
  assign _T_54659 = $signed(_T_54658); // @[Modules.scala 37:46:@563.4]
  assign _T_54660 = $signed(io_in_618) + $signed(io_in_619); // @[Modules.scala 37:46:@567.4]
  assign _T_54661 = _T_54660[4:0]; // @[Modules.scala 37:46:@568.4]
  assign _T_54662 = $signed(_T_54661); // @[Modules.scala 37:46:@569.4]
  assign _T_54672 = $signed(io_in_640) + $signed(io_in_641); // @[Modules.scala 37:46:@581.4]
  assign _T_54673 = _T_54672[4:0]; // @[Modules.scala 37:46:@582.4]
  assign _T_54674 = $signed(_T_54673); // @[Modules.scala 37:46:@583.4]
  assign _T_54675 = $signed(io_in_646) + $signed(io_in_647); // @[Modules.scala 37:46:@587.4]
  assign _T_54676 = _T_54675[4:0]; // @[Modules.scala 37:46:@588.4]
  assign _T_54677 = $signed(_T_54676); // @[Modules.scala 37:46:@589.4]
  assign _T_54685 = $signed(io_in_664) + $signed(io_in_665); // @[Modules.scala 37:46:@599.4]
  assign _T_54686 = _T_54685[4:0]; // @[Modules.scala 37:46:@600.4]
  assign _T_54687 = $signed(_T_54686); // @[Modules.scala 37:46:@601.4]
  assign _T_54688 = $signed(io_in_666) + $signed(io_in_667); // @[Modules.scala 37:46:@603.4]
  assign _T_54689 = _T_54688[4:0]; // @[Modules.scala 37:46:@604.4]
  assign _T_54690 = $signed(_T_54689); // @[Modules.scala 37:46:@605.4]
  assign _T_54691 = $signed(io_in_668) + $signed(io_in_669); // @[Modules.scala 37:46:@607.4]
  assign _T_54692 = _T_54691[4:0]; // @[Modules.scala 37:46:@608.4]
  assign _T_54693 = $signed(_T_54692); // @[Modules.scala 37:46:@609.4]
  assign _T_54695 = $signed(io_in_676) + $signed(io_in_677); // @[Modules.scala 37:46:@614.4]
  assign _T_54696 = _T_54695[4:0]; // @[Modules.scala 37:46:@615.4]
  assign _T_54697 = $signed(_T_54696); // @[Modules.scala 37:46:@616.4]
  assign _T_54698 = $signed(io_in_678) + $signed(io_in_679); // @[Modules.scala 37:46:@618.4]
  assign _T_54699 = _T_54698[4:0]; // @[Modules.scala 37:46:@619.4]
  assign _T_54700 = $signed(_T_54699); // @[Modules.scala 37:46:@620.4]
  assign _T_54701 = $signed(io_in_680) + $signed(io_in_681); // @[Modules.scala 37:46:@622.4]
  assign _T_54702 = _T_54701[4:0]; // @[Modules.scala 37:46:@623.4]
  assign _T_54703 = $signed(_T_54702); // @[Modules.scala 37:46:@624.4]
  assign _T_54706 = $signed(io_in_688) + $signed(io_in_689); // @[Modules.scala 37:46:@629.4]
  assign _T_54707 = _T_54706[4:0]; // @[Modules.scala 37:46:@630.4]
  assign _T_54708 = $signed(_T_54707); // @[Modules.scala 37:46:@631.4]
  assign _T_54709 = $signed(io_in_690) + $signed(io_in_691); // @[Modules.scala 37:46:@633.4]
  assign _T_54710 = _T_54709[4:0]; // @[Modules.scala 37:46:@634.4]
  assign _T_54711 = $signed(_T_54710); // @[Modules.scala 37:46:@635.4]
  assign _T_54712 = $signed(io_in_692) + $signed(io_in_693); // @[Modules.scala 37:46:@637.4]
  assign _T_54713 = _T_54712[4:0]; // @[Modules.scala 37:46:@638.4]
  assign _T_54714 = $signed(_T_54713); // @[Modules.scala 37:46:@639.4]
  assign _T_54715 = $signed(io_in_694) + $signed(io_in_695); // @[Modules.scala 37:46:@641.4]
  assign _T_54716 = _T_54715[4:0]; // @[Modules.scala 37:46:@642.4]
  assign _T_54717 = $signed(_T_54716); // @[Modules.scala 37:46:@643.4]
  assign _T_54718 = $signed(io_in_696) + $signed(io_in_697); // @[Modules.scala 37:46:@645.4]
  assign _T_54719 = _T_54718[4:0]; // @[Modules.scala 37:46:@646.4]
  assign _T_54720 = $signed(_T_54719); // @[Modules.scala 37:46:@647.4]
  assign _T_54721 = $signed(io_in_704) + $signed(io_in_705); // @[Modules.scala 37:46:@652.4]
  assign _T_54722 = _T_54721[4:0]; // @[Modules.scala 37:46:@653.4]
  assign _T_54723 = $signed(_T_54722); // @[Modules.scala 37:46:@654.4]
  assign _T_54724 = $signed(io_in_706) + $signed(io_in_707); // @[Modules.scala 37:46:@656.4]
  assign _T_54725 = _T_54724[4:0]; // @[Modules.scala 37:46:@657.4]
  assign _T_54726 = $signed(_T_54725); // @[Modules.scala 37:46:@658.4]
  assign _T_54727 = $signed(io_in_708) + $signed(io_in_709); // @[Modules.scala 37:46:@660.4]
  assign _T_54728 = _T_54727[4:0]; // @[Modules.scala 37:46:@661.4]
  assign _T_54729 = $signed(_T_54728); // @[Modules.scala 37:46:@662.4]
  assign _T_54730 = $signed(io_in_712) + $signed(io_in_713); // @[Modules.scala 37:46:@665.4]
  assign _T_54731 = _T_54730[4:0]; // @[Modules.scala 37:46:@666.4]
  assign _T_54732 = $signed(_T_54731); // @[Modules.scala 37:46:@667.4]
  assign _T_54733 = $signed(io_in_714) + $signed(io_in_715); // @[Modules.scala 37:46:@669.4]
  assign _T_54734 = _T_54733[4:0]; // @[Modules.scala 37:46:@670.4]
  assign _T_54735 = $signed(_T_54734); // @[Modules.scala 37:46:@671.4]
  assign _T_54736 = $signed(io_in_716) + $signed(io_in_717); // @[Modules.scala 37:46:@673.4]
  assign _T_54737 = _T_54736[4:0]; // @[Modules.scala 37:46:@674.4]
  assign _T_54738 = $signed(_T_54737); // @[Modules.scala 37:46:@675.4]
  assign _T_54739 = $signed(io_in_718) + $signed(io_in_719); // @[Modules.scala 37:46:@677.4]
  assign _T_54740 = _T_54739[4:0]; // @[Modules.scala 37:46:@678.4]
  assign _T_54741 = $signed(_T_54740); // @[Modules.scala 37:46:@679.4]
  assign _T_54742 = $signed(io_in_720) + $signed(io_in_721); // @[Modules.scala 37:46:@681.4]
  assign _T_54743 = _T_54742[4:0]; // @[Modules.scala 37:46:@682.4]
  assign _T_54744 = $signed(_T_54743); // @[Modules.scala 37:46:@683.4]
  assign _T_54745 = $signed(io_in_722) + $signed(io_in_723); // @[Modules.scala 37:46:@685.4]
  assign _T_54746 = _T_54745[4:0]; // @[Modules.scala 37:46:@686.4]
  assign _T_54747 = $signed(_T_54746); // @[Modules.scala 37:46:@687.4]
  assign _T_54749 = $signed(io_in_732) + $signed(io_in_733); // @[Modules.scala 37:46:@693.4]
  assign _T_54750 = _T_54749[4:0]; // @[Modules.scala 37:46:@694.4]
  assign _T_54751 = $signed(_T_54750); // @[Modules.scala 37:46:@695.4]
  assign _T_54752 = $signed(io_in_734) + $signed(io_in_735); // @[Modules.scala 37:46:@697.4]
  assign _T_54753 = _T_54752[4:0]; // @[Modules.scala 37:46:@698.4]
  assign _T_54754 = $signed(_T_54753); // @[Modules.scala 37:46:@699.4]
  assign _T_54759 = $signed(io_in_748) + $signed(io_in_749); // @[Modules.scala 37:46:@707.4]
  assign _T_54760 = _T_54759[4:0]; // @[Modules.scala 37:46:@708.4]
  assign _T_54761 = $signed(_T_54760); // @[Modules.scala 37:46:@709.4]
  assign _T_54762 = $signed(io_in_752) + $signed(io_in_753); // @[Modules.scala 37:46:@712.4]
  assign _T_54763 = _T_54762[4:0]; // @[Modules.scala 37:46:@713.4]
  assign _T_54764 = $signed(_T_54763); // @[Modules.scala 37:46:@714.4]
  assign _T_54765 = $signed(io_in_754) + $signed(io_in_755); // @[Modules.scala 37:46:@716.4]
  assign _T_54766 = _T_54765[4:0]; // @[Modules.scala 37:46:@717.4]
  assign _T_54767 = $signed(_T_54766); // @[Modules.scala 37:46:@718.4]
  assign _T_54774 = $signed(io_in_776) + $signed(io_in_777); // @[Modules.scala 37:46:@730.4]
  assign _T_54775 = _T_54774[4:0]; // @[Modules.scala 37:46:@731.4]
  assign _T_54776 = $signed(_T_54775); // @[Modules.scala 37:46:@732.4]
  assign _T_54778 = $signed(io_in_782) + $signed(io_in_783); // @[Modules.scala 37:46:@736.4]
  assign _T_54779 = _T_54778[4:0]; // @[Modules.scala 37:46:@737.4]
  assign _T_54780 = $signed(_T_54779); // @[Modules.scala 37:46:@738.4]
  assign buffer_0_0 = {{6{io_in_1[4]}},io_in_1}; // @[Modules.scala 32:22:@8.4]
  assign _T_54781 = $signed(buffer_0_0) + $signed(11'sh0); // @[Modules.scala 65:57:@740.4]
  assign _T_54782 = _T_54781[10:0]; // @[Modules.scala 65:57:@741.4]
  assign buffer_0_392 = $signed(_T_54782); // @[Modules.scala 65:57:@742.4]
  assign buffer_0_2 = {{6{io_in_5[4]}},io_in_5}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_3 = {{6{io_in_7[4]}},io_in_7}; // @[Modules.scala 32:22:@8.4]
  assign _T_54784 = $signed(buffer_0_2) + $signed(buffer_0_3); // @[Modules.scala 65:57:@744.4]
  assign _T_54785 = _T_54784[10:0]; // @[Modules.scala 65:57:@745.4]
  assign buffer_0_393 = $signed(_T_54785); // @[Modules.scala 65:57:@746.4]
  assign buffer_0_4 = {{6{io_in_9[4]}},io_in_9}; // @[Modules.scala 32:22:@8.4]
  assign _T_54787 = $signed(buffer_0_4) + $signed(11'sh0); // @[Modules.scala 65:57:@748.4]
  assign _T_54788 = _T_54787[10:0]; // @[Modules.scala 65:57:@749.4]
  assign buffer_0_394 = $signed(_T_54788); // @[Modules.scala 65:57:@750.4]
  assign _T_54790 = $signed(11'sh0) + $signed(11'sh0); // @[Modules.scala 65:57:@752.4]
  assign _T_54791 = _T_54790[10:0]; // @[Modules.scala 65:57:@753.4]
  assign buffer_0_395 = $signed(_T_54791); // @[Modules.scala 65:57:@754.4]
  assign buffer_0_8 = {{6{_T_54272[4]}},_T_54272}; // @[Modules.scala 32:22:@8.4]
  assign _T_54793 = $signed(buffer_0_8) + $signed(11'sh0); // @[Modules.scala 65:57:@756.4]
  assign _T_54794 = _T_54793[10:0]; // @[Modules.scala 65:57:@757.4]
  assign buffer_0_396 = $signed(_T_54794); // @[Modules.scala 65:57:@758.4]
  assign buffer_0_10 = {{6{_T_54276[4]}},_T_54276}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_11 = {{6{io_in_23[4]}},io_in_23}; // @[Modules.scala 32:22:@8.4]
  assign _T_54796 = $signed(buffer_0_10) + $signed(buffer_0_11); // @[Modules.scala 65:57:@760.4]
  assign _T_54797 = _T_54796[10:0]; // @[Modules.scala 65:57:@761.4]
  assign buffer_0_397 = $signed(_T_54797); // @[Modules.scala 65:57:@762.4]
  assign buffer_0_12 = {{6{io_in_25[4]}},io_in_25}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_13 = {{6{io_in_26[4]}},io_in_26}; // @[Modules.scala 32:22:@8.4]
  assign _T_54799 = $signed(buffer_0_12) + $signed(buffer_0_13); // @[Modules.scala 65:57:@764.4]
  assign _T_54800 = _T_54799[10:0]; // @[Modules.scala 65:57:@765.4]
  assign buffer_0_398 = $signed(_T_54800); // @[Modules.scala 65:57:@766.4]
  assign buffer_0_15 = {{6{io_in_31[4]}},io_in_31}; // @[Modules.scala 32:22:@8.4]
  assign _T_54802 = $signed(11'sh0) + $signed(buffer_0_15); // @[Modules.scala 65:57:@768.4]
  assign _T_54803 = _T_54802[10:0]; // @[Modules.scala 65:57:@769.4]
  assign buffer_0_399 = $signed(_T_54803); // @[Modules.scala 65:57:@770.4]
  assign buffer_0_16 = {{6{_T_54280[4]}},_T_54280}; // @[Modules.scala 32:22:@8.4]
  assign _T_54805 = $signed(buffer_0_16) + $signed(11'sh0); // @[Modules.scala 65:57:@772.4]
  assign _T_54806 = _T_54805[10:0]; // @[Modules.scala 65:57:@773.4]
  assign buffer_0_400 = $signed(_T_54806); // @[Modules.scala 65:57:@774.4]
  assign buffer_0_26 = {{6{_T_54292[4]}},_T_54292}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_27 = {{6{io_in_54[4]}},io_in_54}; // @[Modules.scala 32:22:@8.4]
  assign _T_54820 = $signed(buffer_0_26) + $signed(buffer_0_27); // @[Modules.scala 65:57:@792.4]
  assign _T_54821 = _T_54820[10:0]; // @[Modules.scala 65:57:@793.4]
  assign buffer_0_405 = $signed(_T_54821); // @[Modules.scala 65:57:@794.4]
  assign buffer_0_28 = {{6{io_in_56[4]}},io_in_56}; // @[Modules.scala 32:22:@8.4]
  assign _T_54823 = $signed(buffer_0_28) + $signed(11'sh0); // @[Modules.scala 65:57:@796.4]
  assign _T_54824 = _T_54823[10:0]; // @[Modules.scala 65:57:@797.4]
  assign buffer_0_406 = $signed(_T_54824); // @[Modules.scala 65:57:@798.4]
  assign buffer_0_32 = {{6{io_in_65[4]}},io_in_65}; // @[Modules.scala 32:22:@8.4]
  assign _T_54829 = $signed(buffer_0_32) + $signed(11'sh0); // @[Modules.scala 65:57:@804.4]
  assign _T_54830 = _T_54829[10:0]; // @[Modules.scala 65:57:@805.4]
  assign buffer_0_408 = $signed(_T_54830); // @[Modules.scala 65:57:@806.4]
  assign buffer_0_37 = {{6{io_in_75[4]}},io_in_75}; // @[Modules.scala 32:22:@8.4]
  assign _T_54835 = $signed(11'sh0) + $signed(buffer_0_37); // @[Modules.scala 65:57:@812.4]
  assign _T_54836 = _T_54835[10:0]; // @[Modules.scala 65:57:@813.4]
  assign buffer_0_410 = $signed(_T_54836); // @[Modules.scala 65:57:@814.4]
  assign buffer_0_38 = {{6{io_in_76[4]}},io_in_76}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_39 = {{6{_T_54302[4]}},_T_54302}; // @[Modules.scala 32:22:@8.4]
  assign _T_54838 = $signed(buffer_0_38) + $signed(buffer_0_39); // @[Modules.scala 65:57:@816.4]
  assign _T_54839 = _T_54838[10:0]; // @[Modules.scala 65:57:@817.4]
  assign buffer_0_411 = $signed(_T_54839); // @[Modules.scala 65:57:@818.4]
  assign buffer_0_41 = {{6{io_in_82[4]}},io_in_82}; // @[Modules.scala 32:22:@8.4]
  assign _T_54841 = $signed(11'sh0) + $signed(buffer_0_41); // @[Modules.scala 65:57:@820.4]
  assign _T_54842 = _T_54841[10:0]; // @[Modules.scala 65:57:@821.4]
  assign buffer_0_412 = $signed(_T_54842); // @[Modules.scala 65:57:@822.4]
  assign buffer_0_42 = {{6{io_in_84[4]}},io_in_84}; // @[Modules.scala 32:22:@8.4]
  assign _T_54844 = $signed(buffer_0_42) + $signed(11'sh0); // @[Modules.scala 65:57:@824.4]
  assign _T_54845 = _T_54844[10:0]; // @[Modules.scala 65:57:@825.4]
  assign buffer_0_413 = $signed(_T_54845); // @[Modules.scala 65:57:@826.4]
  assign buffer_0_44 = {{6{_T_54307[4]}},_T_54307}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_45 = {{6{_T_54310[4]}},_T_54310}; // @[Modules.scala 32:22:@8.4]
  assign _T_54847 = $signed(buffer_0_44) + $signed(buffer_0_45); // @[Modules.scala 65:57:@828.4]
  assign _T_54848 = _T_54847[10:0]; // @[Modules.scala 65:57:@829.4]
  assign buffer_0_414 = $signed(_T_54848); // @[Modules.scala 65:57:@830.4]
  assign buffer_0_46 = {{6{io_in_93[4]}},io_in_93}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_47 = {{6{_T_54313[4]}},_T_54313}; // @[Modules.scala 32:22:@8.4]
  assign _T_54850 = $signed(buffer_0_46) + $signed(buffer_0_47); // @[Modules.scala 65:57:@832.4]
  assign _T_54851 = _T_54850[10:0]; // @[Modules.scala 65:57:@833.4]
  assign buffer_0_415 = $signed(_T_54851); // @[Modules.scala 65:57:@834.4]
  assign buffer_0_48 = {{6{io_in_97[4]}},io_in_97}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_49 = {{6{_T_54316[4]}},_T_54316}; // @[Modules.scala 32:22:@8.4]
  assign _T_54853 = $signed(buffer_0_48) + $signed(buffer_0_49); // @[Modules.scala 65:57:@836.4]
  assign _T_54854 = _T_54853[10:0]; // @[Modules.scala 65:57:@837.4]
  assign buffer_0_416 = $signed(_T_54854); // @[Modules.scala 65:57:@838.4]
  assign buffer_0_50 = {{6{_T_54319[4]}},_T_54319}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_51 = {{6{_T_54322[4]}},_T_54322}; // @[Modules.scala 32:22:@8.4]
  assign _T_54856 = $signed(buffer_0_50) + $signed(buffer_0_51); // @[Modules.scala 65:57:@840.4]
  assign _T_54857 = _T_54856[10:0]; // @[Modules.scala 65:57:@841.4]
  assign buffer_0_417 = $signed(_T_54857); // @[Modules.scala 65:57:@842.4]
  assign buffer_0_52 = {{6{_T_54325[4]}},_T_54325}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_53 = {{6{_T_54328[4]}},_T_54328}; // @[Modules.scala 32:22:@8.4]
  assign _T_54859 = $signed(buffer_0_52) + $signed(buffer_0_53); // @[Modules.scala 65:57:@844.4]
  assign _T_54860 = _T_54859[10:0]; // @[Modules.scala 65:57:@845.4]
  assign buffer_0_418 = $signed(_T_54860); // @[Modules.scala 65:57:@846.4]
  assign buffer_0_54 = {{6{io_in_108[4]}},io_in_108}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_55 = {{6{_T_54331[4]}},_T_54331}; // @[Modules.scala 32:22:@8.4]
  assign _T_54862 = $signed(buffer_0_54) + $signed(buffer_0_55); // @[Modules.scala 65:57:@848.4]
  assign _T_54863 = _T_54862[10:0]; // @[Modules.scala 65:57:@849.4]
  assign buffer_0_419 = $signed(_T_54863); // @[Modules.scala 65:57:@850.4]
  assign buffer_0_56 = {{6{io_in_113[4]}},io_in_113}; // @[Modules.scala 32:22:@8.4]
  assign _T_54865 = $signed(buffer_0_56) + $signed(11'sh0); // @[Modules.scala 65:57:@852.4]
  assign _T_54866 = _T_54865[10:0]; // @[Modules.scala 65:57:@853.4]
  assign buffer_0_420 = $signed(_T_54866); // @[Modules.scala 65:57:@854.4]
  assign buffer_0_58 = {{6{io_in_116[4]}},io_in_116}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_59 = {{6{_T_54335[4]}},_T_54335}; // @[Modules.scala 32:22:@8.4]
  assign _T_54868 = $signed(buffer_0_58) + $signed(buffer_0_59); // @[Modules.scala 65:57:@856.4]
  assign _T_54869 = _T_54868[10:0]; // @[Modules.scala 65:57:@857.4]
  assign buffer_0_421 = $signed(_T_54869); // @[Modules.scala 65:57:@858.4]
  assign buffer_0_64 = {{6{io_in_129[4]}},io_in_129}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_65 = {{6{io_in_131[4]}},io_in_131}; // @[Modules.scala 32:22:@8.4]
  assign _T_54877 = $signed(buffer_0_64) + $signed(buffer_0_65); // @[Modules.scala 65:57:@868.4]
  assign _T_54878 = _T_54877[10:0]; // @[Modules.scala 65:57:@869.4]
  assign buffer_0_424 = $signed(_T_54878); // @[Modules.scala 65:57:@870.4]
  assign buffer_0_66 = {{6{_T_54342[4]}},_T_54342}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_67 = {{6{_T_54345[4]}},_T_54345}; // @[Modules.scala 32:22:@8.4]
  assign _T_54880 = $signed(buffer_0_66) + $signed(buffer_0_67); // @[Modules.scala 65:57:@872.4]
  assign _T_54881 = _T_54880[10:0]; // @[Modules.scala 65:57:@873.4]
  assign buffer_0_425 = $signed(_T_54881); // @[Modules.scala 65:57:@874.4]
  assign buffer_0_68 = {{6{io_in_136[4]}},io_in_136}; // @[Modules.scala 32:22:@8.4]
  assign _T_54883 = $signed(buffer_0_68) + $signed(11'sh0); // @[Modules.scala 65:57:@876.4]
  assign _T_54884 = _T_54883[10:0]; // @[Modules.scala 65:57:@877.4]
  assign buffer_0_426 = $signed(_T_54884); // @[Modules.scala 65:57:@878.4]
  assign buffer_0_70 = {{6{_T_54349[4]}},_T_54349}; // @[Modules.scala 32:22:@8.4]
  assign _T_54886 = $signed(buffer_0_70) + $signed(11'sh0); // @[Modules.scala 65:57:@880.4]
  assign _T_54887 = _T_54886[10:0]; // @[Modules.scala 65:57:@881.4]
  assign buffer_0_427 = $signed(_T_54887); // @[Modules.scala 65:57:@882.4]
  assign buffer_0_72 = {{6{io_in_144[4]}},io_in_144}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_73 = {{6{_T_54353[4]}},_T_54353}; // @[Modules.scala 32:22:@8.4]
  assign _T_54889 = $signed(buffer_0_72) + $signed(buffer_0_73); // @[Modules.scala 65:57:@884.4]
  assign _T_54890 = _T_54889[10:0]; // @[Modules.scala 65:57:@885.4]
  assign buffer_0_428 = $signed(_T_54890); // @[Modules.scala 65:57:@886.4]
  assign buffer_0_74 = {{6{_T_54356[4]}},_T_54356}; // @[Modules.scala 32:22:@8.4]
  assign _T_54892 = $signed(buffer_0_74) + $signed(11'sh0); // @[Modules.scala 65:57:@888.4]
  assign _T_54893 = _T_54892[10:0]; // @[Modules.scala 65:57:@889.4]
  assign buffer_0_429 = $signed(_T_54893); // @[Modules.scala 65:57:@890.4]
  assign buffer_0_81 = {{6{_T_54365[4]}},_T_54365}; // @[Modules.scala 32:22:@8.4]
  assign _T_54901 = $signed(11'sh0) + $signed(buffer_0_81); // @[Modules.scala 65:57:@900.4]
  assign _T_54902 = _T_54901[10:0]; // @[Modules.scala 65:57:@901.4]
  assign buffer_0_432 = $signed(_T_54902); // @[Modules.scala 65:57:@902.4]
  assign buffer_0_82 = {{6{io_in_164[4]}},io_in_164}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_83 = {{6{io_in_167[4]}},io_in_167}; // @[Modules.scala 32:22:@8.4]
  assign _T_54904 = $signed(buffer_0_82) + $signed(buffer_0_83); // @[Modules.scala 65:57:@904.4]
  assign _T_54905 = _T_54904[10:0]; // @[Modules.scala 65:57:@905.4]
  assign buffer_0_433 = $signed(_T_54905); // @[Modules.scala 65:57:@906.4]
  assign buffer_0_86 = {{6{io_in_172[4]}},io_in_172}; // @[Modules.scala 32:22:@8.4]
  assign _T_54910 = $signed(buffer_0_86) + $signed(11'sh0); // @[Modules.scala 65:57:@912.4]
  assign _T_54911 = _T_54910[10:0]; // @[Modules.scala 65:57:@913.4]
  assign buffer_0_435 = $signed(_T_54911); // @[Modules.scala 65:57:@914.4]
  assign buffer_0_93 = {{6{_T_54376[4]}},_T_54376}; // @[Modules.scala 32:22:@8.4]
  assign _T_54919 = $signed(11'sh0) + $signed(buffer_0_93); // @[Modules.scala 65:57:@924.4]
  assign _T_54920 = _T_54919[10:0]; // @[Modules.scala 65:57:@925.4]
  assign buffer_0_438 = $signed(_T_54920); // @[Modules.scala 65:57:@926.4]
  assign buffer_0_95 = {{6{io_in_190[4]}},io_in_190}; // @[Modules.scala 32:22:@8.4]
  assign _T_54922 = $signed(11'sh0) + $signed(buffer_0_95); // @[Modules.scala 65:57:@928.4]
  assign _T_54923 = _T_54922[10:0]; // @[Modules.scala 65:57:@929.4]
  assign buffer_0_439 = $signed(_T_54923); // @[Modules.scala 65:57:@930.4]
  assign buffer_0_98 = {{6{io_in_196[4]}},io_in_196}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_99 = {{6{io_in_198[4]}},io_in_198}; // @[Modules.scala 32:22:@8.4]
  assign _T_54928 = $signed(buffer_0_98) + $signed(buffer_0_99); // @[Modules.scala 65:57:@936.4]
  assign _T_54929 = _T_54928[10:0]; // @[Modules.scala 65:57:@937.4]
  assign buffer_0_441 = $signed(_T_54929); // @[Modules.scala 65:57:@938.4]
  assign buffer_0_103 = {{6{io_in_207[4]}},io_in_207}; // @[Modules.scala 32:22:@8.4]
  assign _T_54934 = $signed(11'sh0) + $signed(buffer_0_103); // @[Modules.scala 65:57:@944.4]
  assign _T_54935 = _T_54934[10:0]; // @[Modules.scala 65:57:@945.4]
  assign buffer_0_443 = $signed(_T_54935); // @[Modules.scala 65:57:@946.4]
  assign buffer_0_104 = {{6{io_in_209[4]}},io_in_209}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_105 = {{6{_T_54385[4]}},_T_54385}; // @[Modules.scala 32:22:@8.4]
  assign _T_54937 = $signed(buffer_0_104) + $signed(buffer_0_105); // @[Modules.scala 65:57:@948.4]
  assign _T_54938 = _T_54937[10:0]; // @[Modules.scala 65:57:@949.4]
  assign buffer_0_444 = $signed(_T_54938); // @[Modules.scala 65:57:@950.4]
  assign buffer_0_106 = {{6{io_in_212[4]}},io_in_212}; // @[Modules.scala 32:22:@8.4]
  assign _T_54940 = $signed(buffer_0_106) + $signed(11'sh0); // @[Modules.scala 65:57:@952.4]
  assign _T_54941 = _T_54940[10:0]; // @[Modules.scala 65:57:@953.4]
  assign buffer_0_445 = $signed(_T_54941); // @[Modules.scala 65:57:@954.4]
  assign buffer_0_118 = {{6{io_in_237[4]}},io_in_237}; // @[Modules.scala 32:22:@8.4]
  assign _T_54958 = $signed(buffer_0_118) + $signed(11'sh0); // @[Modules.scala 65:57:@976.4]
  assign _T_54959 = _T_54958[10:0]; // @[Modules.scala 65:57:@977.4]
  assign buffer_0_451 = $signed(_T_54959); // @[Modules.scala 65:57:@978.4]
  assign buffer_0_131 = {{6{io_in_262[4]}},io_in_262}; // @[Modules.scala 32:22:@8.4]
  assign _T_54976 = $signed(11'sh0) + $signed(buffer_0_131); // @[Modules.scala 65:57:@1000.4]
  assign _T_54977 = _T_54976[10:0]; // @[Modules.scala 65:57:@1001.4]
  assign buffer_0_457 = $signed(_T_54977); // @[Modules.scala 65:57:@1002.4]
  assign buffer_0_144 = {{6{io_in_289[4]}},io_in_289}; // @[Modules.scala 32:22:@8.4]
  assign _T_54997 = $signed(buffer_0_144) + $signed(11'sh0); // @[Modules.scala 65:57:@1028.4]
  assign _T_54998 = _T_54997[10:0]; // @[Modules.scala 65:57:@1029.4]
  assign buffer_0_464 = $signed(_T_54998); // @[Modules.scala 65:57:@1030.4]
  assign buffer_0_157 = {{6{io_in_315[4]}},io_in_315}; // @[Modules.scala 32:22:@8.4]
  assign _T_55015 = $signed(11'sh0) + $signed(buffer_0_157); // @[Modules.scala 65:57:@1052.4]
  assign _T_55016 = _T_55015[10:0]; // @[Modules.scala 65:57:@1053.4]
  assign buffer_0_470 = $signed(_T_55016); // @[Modules.scala 65:57:@1054.4]
  assign buffer_0_158 = {{6{_T_54435[4]}},_T_54435}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_159 = {{6{_T_54438[4]}},_T_54438}; // @[Modules.scala 32:22:@8.4]
  assign _T_55018 = $signed(buffer_0_158) + $signed(buffer_0_159); // @[Modules.scala 65:57:@1056.4]
  assign _T_55019 = _T_55018[10:0]; // @[Modules.scala 65:57:@1057.4]
  assign buffer_0_471 = $signed(_T_55019); // @[Modules.scala 65:57:@1058.4]
  assign buffer_0_162 = {{6{io_in_325[4]}},io_in_325}; // @[Modules.scala 32:22:@8.4]
  assign _T_55024 = $signed(buffer_0_162) + $signed(11'sh0); // @[Modules.scala 65:57:@1064.4]
  assign _T_55025 = _T_55024[10:0]; // @[Modules.scala 65:57:@1065.4]
  assign buffer_0_473 = $signed(_T_55025); // @[Modules.scala 65:57:@1066.4]
  assign buffer_0_164 = {{6{_T_54444[4]}},_T_54444}; // @[Modules.scala 32:22:@8.4]
  assign _T_55027 = $signed(buffer_0_164) + $signed(11'sh0); // @[Modules.scala 65:57:@1068.4]
  assign _T_55028 = _T_55027[10:0]; // @[Modules.scala 65:57:@1069.4]
  assign buffer_0_474 = $signed(_T_55028); // @[Modules.scala 65:57:@1070.4]
  assign buffer_0_167 = {{6{io_in_335[4]}},io_in_335}; // @[Modules.scala 32:22:@8.4]
  assign _T_55030 = $signed(11'sh0) + $signed(buffer_0_167); // @[Modules.scala 65:57:@1072.4]
  assign _T_55031 = _T_55030[10:0]; // @[Modules.scala 65:57:@1073.4]
  assign buffer_0_475 = $signed(_T_55031); // @[Modules.scala 65:57:@1074.4]
  assign buffer_0_168 = {{6{io_in_336[4]}},io_in_336}; // @[Modules.scala 32:22:@8.4]
  assign _T_55033 = $signed(buffer_0_168) + $signed(11'sh0); // @[Modules.scala 65:57:@1076.4]
  assign _T_55034 = _T_55033[10:0]; // @[Modules.scala 65:57:@1077.4]
  assign buffer_0_476 = $signed(_T_55034); // @[Modules.scala 65:57:@1078.4]
  assign buffer_0_170 = {{6{io_in_341[4]}},io_in_341}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_171 = {{6{_T_54450[4]}},_T_54450}; // @[Modules.scala 32:22:@8.4]
  assign _T_55036 = $signed(buffer_0_170) + $signed(buffer_0_171); // @[Modules.scala 65:57:@1080.4]
  assign _T_55037 = _T_55036[10:0]; // @[Modules.scala 65:57:@1081.4]
  assign buffer_0_477 = $signed(_T_55037); // @[Modules.scala 65:57:@1082.4]
  assign buffer_0_172 = {{6{_T_54453[4]}},_T_54453}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_173 = {{6{_T_54456[4]}},_T_54456}; // @[Modules.scala 32:22:@8.4]
  assign _T_55039 = $signed(buffer_0_172) + $signed(buffer_0_173); // @[Modules.scala 65:57:@1084.4]
  assign _T_55040 = _T_55039[10:0]; // @[Modules.scala 65:57:@1085.4]
  assign buffer_0_478 = $signed(_T_55040); // @[Modules.scala 65:57:@1086.4]
  assign buffer_0_174 = {{6{_T_54459[4]}},_T_54459}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_175 = {{6{_T_54462[4]}},_T_54462}; // @[Modules.scala 32:22:@8.4]
  assign _T_55042 = $signed(buffer_0_174) + $signed(buffer_0_175); // @[Modules.scala 65:57:@1088.4]
  assign _T_55043 = _T_55042[10:0]; // @[Modules.scala 65:57:@1089.4]
  assign buffer_0_479 = $signed(_T_55043); // @[Modules.scala 65:57:@1090.4]
  assign buffer_0_176 = {{6{_T_54465[4]}},_T_54465}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_177 = {{6{_T_54468[4]}},_T_54468}; // @[Modules.scala 32:22:@8.4]
  assign _T_55045 = $signed(buffer_0_176) + $signed(buffer_0_177); // @[Modules.scala 65:57:@1092.4]
  assign _T_55046 = _T_55045[10:0]; // @[Modules.scala 65:57:@1093.4]
  assign buffer_0_480 = $signed(_T_55046); // @[Modules.scala 65:57:@1094.4]
  assign buffer_0_178 = {{6{_T_54471[4]}},_T_54471}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_179 = {{6{_T_54474[4]}},_T_54474}; // @[Modules.scala 32:22:@8.4]
  assign _T_55048 = $signed(buffer_0_178) + $signed(buffer_0_179); // @[Modules.scala 65:57:@1096.4]
  assign _T_55049 = _T_55048[10:0]; // @[Modules.scala 65:57:@1097.4]
  assign buffer_0_481 = $signed(_T_55049); // @[Modules.scala 65:57:@1098.4]
  assign buffer_0_181 = {{6{io_in_363[4]}},io_in_363}; // @[Modules.scala 32:22:@8.4]
  assign _T_55051 = $signed(11'sh0) + $signed(buffer_0_181); // @[Modules.scala 65:57:@1100.4]
  assign _T_55052 = _T_55051[10:0]; // @[Modules.scala 65:57:@1101.4]
  assign buffer_0_482 = $signed(_T_55052); // @[Modules.scala 65:57:@1102.4]
  assign buffer_0_184 = {{6{_T_54480[4]}},_T_54480}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_185 = {{6{_T_54483[4]}},_T_54483}; // @[Modules.scala 32:22:@8.4]
  assign _T_55057 = $signed(buffer_0_184) + $signed(buffer_0_185); // @[Modules.scala 65:57:@1108.4]
  assign _T_55058 = _T_55057[10:0]; // @[Modules.scala 65:57:@1109.4]
  assign buffer_0_484 = $signed(_T_55058); // @[Modules.scala 65:57:@1110.4]
  assign buffer_0_186 = {{6{_T_54486[4]}},_T_54486}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_187 = {{6{_T_54489[4]}},_T_54489}; // @[Modules.scala 32:22:@8.4]
  assign _T_55060 = $signed(buffer_0_186) + $signed(buffer_0_187); // @[Modules.scala 65:57:@1112.4]
  assign _T_55061 = _T_55060[10:0]; // @[Modules.scala 65:57:@1113.4]
  assign buffer_0_485 = $signed(_T_55061); // @[Modules.scala 65:57:@1114.4]
  assign buffer_0_188 = {{6{_T_54492[4]}},_T_54492}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_189 = {{6{_T_54495[4]}},_T_54495}; // @[Modules.scala 32:22:@8.4]
  assign _T_55063 = $signed(buffer_0_188) + $signed(buffer_0_189); // @[Modules.scala 65:57:@1116.4]
  assign _T_55064 = _T_55063[10:0]; // @[Modules.scala 65:57:@1117.4]
  assign buffer_0_486 = $signed(_T_55064); // @[Modules.scala 65:57:@1118.4]
  assign buffer_0_190 = {{6{_T_54498[4]}},_T_54498}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_191 = {{6{_T_54501[4]}},_T_54501}; // @[Modules.scala 32:22:@8.4]
  assign _T_55066 = $signed(buffer_0_190) + $signed(buffer_0_191); // @[Modules.scala 65:57:@1120.4]
  assign _T_55067 = _T_55066[10:0]; // @[Modules.scala 65:57:@1121.4]
  assign buffer_0_487 = $signed(_T_55067); // @[Modules.scala 65:57:@1122.4]
  assign buffer_0_192 = {{6{io_in_385[4]}},io_in_385}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_193 = {{6{_T_54504[4]}},_T_54504}; // @[Modules.scala 32:22:@8.4]
  assign _T_55069 = $signed(buffer_0_192) + $signed(buffer_0_193); // @[Modules.scala 65:57:@1124.4]
  assign _T_55070 = _T_55069[10:0]; // @[Modules.scala 65:57:@1125.4]
  assign buffer_0_488 = $signed(_T_55070); // @[Modules.scala 65:57:@1126.4]
  assign buffer_0_194 = {{6{io_in_388[4]}},io_in_388}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_195 = {{6{io_in_391[4]}},io_in_391}; // @[Modules.scala 32:22:@8.4]
  assign _T_55072 = $signed(buffer_0_194) + $signed(buffer_0_195); // @[Modules.scala 65:57:@1128.4]
  assign _T_55073 = _T_55072[10:0]; // @[Modules.scala 65:57:@1129.4]
  assign buffer_0_489 = $signed(_T_55073); // @[Modules.scala 65:57:@1130.4]
  assign buffer_0_198 = {{6{_T_54509[4]}},_T_54509}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_199 = {{6{_T_54512[4]}},_T_54512}; // @[Modules.scala 32:22:@8.4]
  assign _T_55078 = $signed(buffer_0_198) + $signed(buffer_0_199); // @[Modules.scala 65:57:@1136.4]
  assign _T_55079 = _T_55078[10:0]; // @[Modules.scala 65:57:@1137.4]
  assign buffer_0_491 = $signed(_T_55079); // @[Modules.scala 65:57:@1138.4]
  assign buffer_0_200 = {{6{_T_54515[4]}},_T_54515}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_201 = {{6{_T_54518[4]}},_T_54518}; // @[Modules.scala 32:22:@8.4]
  assign _T_55081 = $signed(buffer_0_200) + $signed(buffer_0_201); // @[Modules.scala 65:57:@1140.4]
  assign _T_55082 = _T_55081[10:0]; // @[Modules.scala 65:57:@1141.4]
  assign buffer_0_492 = $signed(_T_55082); // @[Modules.scala 65:57:@1142.4]
  assign buffer_0_202 = {{6{_T_54521[4]}},_T_54521}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_203 = {{6{_T_54524[4]}},_T_54524}; // @[Modules.scala 32:22:@8.4]
  assign _T_55084 = $signed(buffer_0_202) + $signed(buffer_0_203); // @[Modules.scala 65:57:@1144.4]
  assign _T_55085 = _T_55084[10:0]; // @[Modules.scala 65:57:@1145.4]
  assign buffer_0_493 = $signed(_T_55085); // @[Modules.scala 65:57:@1146.4]
  assign buffer_0_204 = {{6{_T_54527[4]}},_T_54527}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_205 = {{6{_T_54530[4]}},_T_54530}; // @[Modules.scala 32:22:@8.4]
  assign _T_55087 = $signed(buffer_0_204) + $signed(buffer_0_205); // @[Modules.scala 65:57:@1148.4]
  assign _T_55088 = _T_55087[10:0]; // @[Modules.scala 65:57:@1149.4]
  assign buffer_0_494 = $signed(_T_55088); // @[Modules.scala 65:57:@1150.4]
  assign buffer_0_206 = {{6{_T_54533[4]}},_T_54533}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_207 = {{6{_T_54536[4]}},_T_54536}; // @[Modules.scala 32:22:@8.4]
  assign _T_55090 = $signed(buffer_0_206) + $signed(buffer_0_207); // @[Modules.scala 65:57:@1152.4]
  assign _T_55091 = _T_55090[10:0]; // @[Modules.scala 65:57:@1153.4]
  assign buffer_0_495 = $signed(_T_55091); // @[Modules.scala 65:57:@1154.4]
  assign buffer_0_208 = {{6{io_in_416[4]}},io_in_416}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_209 = {{6{io_in_419[4]}},io_in_419}; // @[Modules.scala 32:22:@8.4]
  assign _T_55093 = $signed(buffer_0_208) + $signed(buffer_0_209); // @[Modules.scala 65:57:@1156.4]
  assign _T_55094 = _T_55093[10:0]; // @[Modules.scala 65:57:@1157.4]
  assign buffer_0_496 = $signed(_T_55094); // @[Modules.scala 65:57:@1158.4]
  assign buffer_0_210 = {{6{io_in_421[4]}},io_in_421}; // @[Modules.scala 32:22:@8.4]
  assign _T_55096 = $signed(buffer_0_210) + $signed(11'sh0); // @[Modules.scala 65:57:@1160.4]
  assign _T_55097 = _T_55096[10:0]; // @[Modules.scala 65:57:@1161.4]
  assign buffer_0_497 = $signed(_T_55097); // @[Modules.scala 65:57:@1162.4]
  assign buffer_0_212 = {{6{io_in_425[4]}},io_in_425}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_213 = {{6{_T_54540[4]}},_T_54540}; // @[Modules.scala 32:22:@8.4]
  assign _T_55099 = $signed(buffer_0_212) + $signed(buffer_0_213); // @[Modules.scala 65:57:@1164.4]
  assign _T_55100 = _T_55099[10:0]; // @[Modules.scala 65:57:@1165.4]
  assign buffer_0_498 = $signed(_T_55100); // @[Modules.scala 65:57:@1166.4]
  assign buffer_0_214 = {{6{_T_54543[4]}},_T_54543}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_215 = {{6{_T_54546[4]}},_T_54546}; // @[Modules.scala 32:22:@8.4]
  assign _T_55102 = $signed(buffer_0_214) + $signed(buffer_0_215); // @[Modules.scala 65:57:@1168.4]
  assign _T_55103 = _T_55102[10:0]; // @[Modules.scala 65:57:@1169.4]
  assign buffer_0_499 = $signed(_T_55103); // @[Modules.scala 65:57:@1170.4]
  assign buffer_0_216 = {{6{_T_54549[4]}},_T_54549}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_217 = {{6{_T_54552[4]}},_T_54552}; // @[Modules.scala 32:22:@8.4]
  assign _T_55105 = $signed(buffer_0_216) + $signed(buffer_0_217); // @[Modules.scala 65:57:@1172.4]
  assign _T_55106 = _T_55105[10:0]; // @[Modules.scala 65:57:@1173.4]
  assign buffer_0_500 = $signed(_T_55106); // @[Modules.scala 65:57:@1174.4]
  assign buffer_0_218 = {{6{_T_54555[4]}},_T_54555}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_219 = {{6{io_in_438[4]}},io_in_438}; // @[Modules.scala 32:22:@8.4]
  assign _T_55108 = $signed(buffer_0_218) + $signed(buffer_0_219); // @[Modules.scala 65:57:@1176.4]
  assign _T_55109 = _T_55108[10:0]; // @[Modules.scala 65:57:@1177.4]
  assign buffer_0_501 = $signed(_T_55109); // @[Modules.scala 65:57:@1178.4]
  assign buffer_0_220 = {{6{io_in_440[4]}},io_in_440}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_221 = {{6{io_in_443[4]}},io_in_443}; // @[Modules.scala 32:22:@8.4]
  assign _T_55111 = $signed(buffer_0_220) + $signed(buffer_0_221); // @[Modules.scala 65:57:@1180.4]
  assign _T_55112 = _T_55111[10:0]; // @[Modules.scala 65:57:@1181.4]
  assign buffer_0_502 = $signed(_T_55112); // @[Modules.scala 65:57:@1182.4]
  assign buffer_0_224 = {{6{_T_54560[4]}},_T_54560}; // @[Modules.scala 32:22:@8.4]
  assign _T_55117 = $signed(buffer_0_224) + $signed(11'sh0); // @[Modules.scala 65:57:@1188.4]
  assign _T_55118 = _T_55117[10:0]; // @[Modules.scala 65:57:@1189.4]
  assign buffer_0_504 = $signed(_T_55118); // @[Modules.scala 65:57:@1190.4]
  assign buffer_0_226 = {{6{io_in_453[4]}},io_in_453}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_227 = {{6{_T_54564[4]}},_T_54564}; // @[Modules.scala 32:22:@8.4]
  assign _T_55120 = $signed(buffer_0_226) + $signed(buffer_0_227); // @[Modules.scala 65:57:@1192.4]
  assign _T_55121 = _T_55120[10:0]; // @[Modules.scala 65:57:@1193.4]
  assign buffer_0_505 = $signed(_T_55121); // @[Modules.scala 65:57:@1194.4]
  assign buffer_0_228 = {{6{_T_54567[4]}},_T_54567}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_229 = {{6{_T_54570[4]}},_T_54570}; // @[Modules.scala 32:22:@8.4]
  assign _T_55123 = $signed(buffer_0_228) + $signed(buffer_0_229); // @[Modules.scala 65:57:@1196.4]
  assign _T_55124 = _T_55123[10:0]; // @[Modules.scala 65:57:@1197.4]
  assign buffer_0_506 = $signed(_T_55124); // @[Modules.scala 65:57:@1198.4]
  assign buffer_0_230 = {{6{io_in_460[4]}},io_in_460}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_231 = {{6{_T_54573[4]}},_T_54573}; // @[Modules.scala 32:22:@8.4]
  assign _T_55126 = $signed(buffer_0_230) + $signed(buffer_0_231); // @[Modules.scala 65:57:@1200.4]
  assign _T_55127 = _T_55126[10:0]; // @[Modules.scala 65:57:@1201.4]
  assign buffer_0_507 = $signed(_T_55127); // @[Modules.scala 65:57:@1202.4]
  assign buffer_0_232 = {{6{_T_54576[4]}},_T_54576}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_233 = {{6{_T_54579[4]}},_T_54579}; // @[Modules.scala 32:22:@8.4]
  assign _T_55129 = $signed(buffer_0_232) + $signed(buffer_0_233); // @[Modules.scala 65:57:@1204.4]
  assign _T_55130 = _T_55129[10:0]; // @[Modules.scala 65:57:@1205.4]
  assign buffer_0_508 = $signed(_T_55130); // @[Modules.scala 65:57:@1206.4]
  assign buffer_0_234 = {{6{io_in_468[4]}},io_in_468}; // @[Modules.scala 32:22:@8.4]
  assign _T_55132 = $signed(buffer_0_234) + $signed(11'sh0); // @[Modules.scala 65:57:@1208.4]
  assign _T_55133 = _T_55132[10:0]; // @[Modules.scala 65:57:@1209.4]
  assign buffer_0_509 = $signed(_T_55133); // @[Modules.scala 65:57:@1210.4]
  assign buffer_0_239 = {{6{io_in_478[4]}},io_in_478}; // @[Modules.scala 32:22:@8.4]
  assign _T_55138 = $signed(11'sh0) + $signed(buffer_0_239); // @[Modules.scala 65:57:@1216.4]
  assign _T_55139 = _T_55138[10:0]; // @[Modules.scala 65:57:@1217.4]
  assign buffer_0_511 = $signed(_T_55139); // @[Modules.scala 65:57:@1218.4]
  assign buffer_0_241 = {{6{_T_54587[4]}},_T_54587}; // @[Modules.scala 32:22:@8.4]
  assign _T_55141 = $signed(11'sh0) + $signed(buffer_0_241); // @[Modules.scala 65:57:@1220.4]
  assign _T_55142 = _T_55141[10:0]; // @[Modules.scala 65:57:@1221.4]
  assign buffer_0_512 = $signed(_T_55142); // @[Modules.scala 65:57:@1222.4]
  assign buffer_0_242 = {{6{_T_54590[4]}},_T_54590}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_243 = {{6{_T_54593[4]}},_T_54593}; // @[Modules.scala 32:22:@8.4]
  assign _T_55144 = $signed(buffer_0_242) + $signed(buffer_0_243); // @[Modules.scala 65:57:@1224.4]
  assign _T_55145 = _T_55144[10:0]; // @[Modules.scala 65:57:@1225.4]
  assign buffer_0_513 = $signed(_T_55145); // @[Modules.scala 65:57:@1226.4]
  assign buffer_0_244 = {{6{io_in_489[4]}},io_in_489}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_245 = {{6{_T_54596[4]}},_T_54596}; // @[Modules.scala 32:22:@8.4]
  assign _T_55147 = $signed(buffer_0_244) + $signed(buffer_0_245); // @[Modules.scala 65:57:@1228.4]
  assign _T_55148 = _T_55147[10:0]; // @[Modules.scala 65:57:@1229.4]
  assign buffer_0_514 = $signed(_T_55148); // @[Modules.scala 65:57:@1230.4]
  assign buffer_0_246 = {{6{io_in_492[4]}},io_in_492}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_247 = {{6{io_in_494[4]}},io_in_494}; // @[Modules.scala 32:22:@8.4]
  assign _T_55150 = $signed(buffer_0_246) + $signed(buffer_0_247); // @[Modules.scala 65:57:@1232.4]
  assign _T_55151 = _T_55150[10:0]; // @[Modules.scala 65:57:@1233.4]
  assign buffer_0_515 = $signed(_T_55151); // @[Modules.scala 65:57:@1234.4]
  assign buffer_0_249 = {{6{_T_54600[4]}},_T_54600}; // @[Modules.scala 32:22:@8.4]
  assign _T_55153 = $signed(11'sh0) + $signed(buffer_0_249); // @[Modules.scala 65:57:@1236.4]
  assign _T_55154 = _T_55153[10:0]; // @[Modules.scala 65:57:@1237.4]
  assign buffer_0_516 = $signed(_T_55154); // @[Modules.scala 65:57:@1238.4]
  assign buffer_0_253 = {{6{io_in_507[4]}},io_in_507}; // @[Modules.scala 32:22:@8.4]
  assign _T_55159 = $signed(11'sh0) + $signed(buffer_0_253); // @[Modules.scala 65:57:@1244.4]
  assign _T_55160 = _T_55159[10:0]; // @[Modules.scala 65:57:@1245.4]
  assign buffer_0_518 = $signed(_T_55160); // @[Modules.scala 65:57:@1246.4]
  assign buffer_0_256 = {{6{_T_54608[4]}},_T_54608}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_257 = {{6{_T_54611[4]}},_T_54611}; // @[Modules.scala 32:22:@8.4]
  assign _T_55165 = $signed(buffer_0_256) + $signed(buffer_0_257); // @[Modules.scala 65:57:@1252.4]
  assign _T_55166 = _T_55165[10:0]; // @[Modules.scala 65:57:@1253.4]
  assign buffer_0_520 = $signed(_T_55166); // @[Modules.scala 65:57:@1254.4]
  assign buffer_0_258 = {{6{io_in_516[4]}},io_in_516}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_259 = {{6{_T_54614[4]}},_T_54614}; // @[Modules.scala 32:22:@8.4]
  assign _T_55168 = $signed(buffer_0_258) + $signed(buffer_0_259); // @[Modules.scala 65:57:@1256.4]
  assign _T_55169 = _T_55168[10:0]; // @[Modules.scala 65:57:@1257.4]
  assign buffer_0_521 = $signed(_T_55169); // @[Modules.scala 65:57:@1258.4]
  assign buffer_0_260 = {{6{io_in_521[4]}},io_in_521}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_261 = {{6{io_in_523[4]}},io_in_523}; // @[Modules.scala 32:22:@8.4]
  assign _T_55171 = $signed(buffer_0_260) + $signed(buffer_0_261); // @[Modules.scala 65:57:@1260.4]
  assign _T_55172 = _T_55171[10:0]; // @[Modules.scala 65:57:@1261.4]
  assign buffer_0_522 = $signed(_T_55172); // @[Modules.scala 65:57:@1262.4]
  assign buffer_0_262 = {{6{io_in_525[4]}},io_in_525}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_263 = {{6{_T_54617[4]}},_T_54617}; // @[Modules.scala 32:22:@8.4]
  assign _T_55174 = $signed(buffer_0_262) + $signed(buffer_0_263); // @[Modules.scala 65:57:@1264.4]
  assign _T_55175 = _T_55174[10:0]; // @[Modules.scala 65:57:@1265.4]
  assign buffer_0_523 = $signed(_T_55175); // @[Modules.scala 65:57:@1266.4]
  assign buffer_0_264 = {{6{_T_54620[4]}},_T_54620}; // @[Modules.scala 32:22:@8.4]
  assign _T_55177 = $signed(buffer_0_264) + $signed(11'sh0); // @[Modules.scala 65:57:@1268.4]
  assign _T_55178 = _T_55177[10:0]; // @[Modules.scala 65:57:@1269.4]
  assign buffer_0_524 = $signed(_T_55178); // @[Modules.scala 65:57:@1270.4]
  assign buffer_0_266 = {{6{io_in_532[4]}},io_in_532}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_267 = {{6{io_in_535[4]}},io_in_535}; // @[Modules.scala 32:22:@8.4]
  assign _T_55180 = $signed(buffer_0_266) + $signed(buffer_0_267); // @[Modules.scala 65:57:@1272.4]
  assign _T_55181 = _T_55180[10:0]; // @[Modules.scala 65:57:@1273.4]
  assign buffer_0_525 = $signed(_T_55181); // @[Modules.scala 65:57:@1274.4]
  assign buffer_0_271 = {{6{io_in_543[4]}},io_in_543}; // @[Modules.scala 32:22:@8.4]
  assign _T_55186 = $signed(11'sh0) + $signed(buffer_0_271); // @[Modules.scala 65:57:@1280.4]
  assign _T_55187 = _T_55186[10:0]; // @[Modules.scala 65:57:@1281.4]
  assign buffer_0_527 = $signed(_T_55187); // @[Modules.scala 65:57:@1282.4]
  assign buffer_0_275 = {{6{io_in_550[4]}},io_in_550}; // @[Modules.scala 32:22:@8.4]
  assign _T_55192 = $signed(11'sh0) + $signed(buffer_0_275); // @[Modules.scala 65:57:@1288.4]
  assign _T_55193 = _T_55192[10:0]; // @[Modules.scala 65:57:@1289.4]
  assign buffer_0_529 = $signed(_T_55193); // @[Modules.scala 65:57:@1290.4]
  assign buffer_0_276 = {{6{io_in_552[4]}},io_in_552}; // @[Modules.scala 32:22:@8.4]
  assign _T_55195 = $signed(buffer_0_276) + $signed(11'sh0); // @[Modules.scala 65:57:@1292.4]
  assign _T_55196 = _T_55195[10:0]; // @[Modules.scala 65:57:@1293.4]
  assign buffer_0_530 = $signed(_T_55196); // @[Modules.scala 65:57:@1294.4]
  assign buffer_0_278 = {{6{io_in_556[4]}},io_in_556}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_279 = {{6{io_in_559[4]}},io_in_559}; // @[Modules.scala 32:22:@8.4]
  assign _T_55198 = $signed(buffer_0_278) + $signed(buffer_0_279); // @[Modules.scala 65:57:@1296.4]
  assign _T_55199 = _T_55198[10:0]; // @[Modules.scala 65:57:@1297.4]
  assign buffer_0_531 = $signed(_T_55199); // @[Modules.scala 65:57:@1298.4]
  assign buffer_0_285 = {{6{io_in_571[4]}},io_in_571}; // @[Modules.scala 32:22:@8.4]
  assign _T_55207 = $signed(11'sh0) + $signed(buffer_0_285); // @[Modules.scala 65:57:@1308.4]
  assign _T_55208 = _T_55207[10:0]; // @[Modules.scala 65:57:@1309.4]
  assign buffer_0_534 = $signed(_T_55208); // @[Modules.scala 65:57:@1310.4]
  assign buffer_0_286 = {{6{io_in_573[4]}},io_in_573}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_287 = {{6{io_in_575[4]}},io_in_575}; // @[Modules.scala 32:22:@8.4]
  assign _T_55210 = $signed(buffer_0_286) + $signed(buffer_0_287); // @[Modules.scala 65:57:@1312.4]
  assign _T_55211 = _T_55210[10:0]; // @[Modules.scala 65:57:@1313.4]
  assign buffer_0_535 = $signed(_T_55211); // @[Modules.scala 65:57:@1314.4]
  assign buffer_0_288 = {{6{_T_54636[4]}},_T_54636}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_289 = {{6{io_in_578[4]}},io_in_578}; // @[Modules.scala 32:22:@8.4]
  assign _T_55213 = $signed(buffer_0_288) + $signed(buffer_0_289); // @[Modules.scala 65:57:@1316.4]
  assign _T_55214 = _T_55213[10:0]; // @[Modules.scala 65:57:@1317.4]
  assign buffer_0_536 = $signed(_T_55214); // @[Modules.scala 65:57:@1318.4]
  assign buffer_0_290 = {{6{io_in_580[4]}},io_in_580}; // @[Modules.scala 32:22:@8.4]
  assign _T_55216 = $signed(buffer_0_290) + $signed(11'sh0); // @[Modules.scala 65:57:@1320.4]
  assign _T_55217 = _T_55216[10:0]; // @[Modules.scala 65:57:@1321.4]
  assign buffer_0_537 = $signed(_T_55217); // @[Modules.scala 65:57:@1322.4]
  assign buffer_0_292 = {{6{_T_54640[4]}},_T_54640}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_293 = {{6{io_in_587[4]}},io_in_587}; // @[Modules.scala 32:22:@8.4]
  assign _T_55219 = $signed(buffer_0_292) + $signed(buffer_0_293); // @[Modules.scala 65:57:@1324.4]
  assign _T_55220 = _T_55219[10:0]; // @[Modules.scala 65:57:@1325.4]
  assign buffer_0_538 = $signed(_T_55220); // @[Modules.scala 65:57:@1326.4]
  assign buffer_0_294 = {{6{io_in_589[4]}},io_in_589}; // @[Modules.scala 32:22:@8.4]
  assign _T_55222 = $signed(buffer_0_294) + $signed(11'sh0); // @[Modules.scala 65:57:@1328.4]
  assign _T_55223 = _T_55222[10:0]; // @[Modules.scala 65:57:@1329.4]
  assign buffer_0_539 = $signed(_T_55223); // @[Modules.scala 65:57:@1330.4]
  assign buffer_0_300 = {{6{_T_54648[4]}},_T_54648}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_301 = {{6{io_in_602[4]}},io_in_602}; // @[Modules.scala 32:22:@8.4]
  assign _T_55231 = $signed(buffer_0_300) + $signed(buffer_0_301); // @[Modules.scala 65:57:@1340.4]
  assign _T_55232 = _T_55231[10:0]; // @[Modules.scala 65:57:@1341.4]
  assign buffer_0_542 = $signed(_T_55232); // @[Modules.scala 65:57:@1342.4]
  assign buffer_0_302 = {{6{_T_54651[4]}},_T_54651}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_303 = {{6{_T_54654[4]}},_T_54654}; // @[Modules.scala 32:22:@8.4]
  assign _T_55234 = $signed(buffer_0_302) + $signed(buffer_0_303); // @[Modules.scala 65:57:@1344.4]
  assign _T_55235 = _T_55234[10:0]; // @[Modules.scala 65:57:@1345.4]
  assign buffer_0_543 = $signed(_T_55235); // @[Modules.scala 65:57:@1346.4]
  assign buffer_0_306 = {{6{_T_54659[4]}},_T_54659}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_307 = {{6{io_in_615[4]}},io_in_615}; // @[Modules.scala 32:22:@8.4]
  assign _T_55240 = $signed(buffer_0_306) + $signed(buffer_0_307); // @[Modules.scala 65:57:@1352.4]
  assign _T_55241 = _T_55240[10:0]; // @[Modules.scala 65:57:@1353.4]
  assign buffer_0_545 = $signed(_T_55241); // @[Modules.scala 65:57:@1354.4]
  assign buffer_0_308 = {{6{io_in_617[4]}},io_in_617}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_309 = {{6{_T_54662[4]}},_T_54662}; // @[Modules.scala 32:22:@8.4]
  assign _T_55243 = $signed(buffer_0_308) + $signed(buffer_0_309); // @[Modules.scala 65:57:@1356.4]
  assign _T_55244 = _T_55243[10:0]; // @[Modules.scala 65:57:@1357.4]
  assign buffer_0_546 = $signed(_T_55244); // @[Modules.scala 65:57:@1358.4]
  assign buffer_0_319 = {{6{io_in_639[4]}},io_in_639}; // @[Modules.scala 32:22:@8.4]
  assign _T_55258 = $signed(11'sh0) + $signed(buffer_0_319); // @[Modules.scala 65:57:@1376.4]
  assign _T_55259 = _T_55258[10:0]; // @[Modules.scala 65:57:@1377.4]
  assign buffer_0_551 = $signed(_T_55259); // @[Modules.scala 65:57:@1378.4]
  assign buffer_0_320 = {{6{_T_54674[4]}},_T_54674}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_321 = {{6{io_in_643[4]}},io_in_643}; // @[Modules.scala 32:22:@8.4]
  assign _T_55261 = $signed(buffer_0_320) + $signed(buffer_0_321); // @[Modules.scala 65:57:@1380.4]
  assign _T_55262 = _T_55261[10:0]; // @[Modules.scala 65:57:@1381.4]
  assign buffer_0_552 = $signed(_T_55262); // @[Modules.scala 65:57:@1382.4]
  assign buffer_0_322 = {{6{io_in_645[4]}},io_in_645}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_323 = {{6{_T_54677[4]}},_T_54677}; // @[Modules.scala 32:22:@8.4]
  assign _T_55264 = $signed(buffer_0_322) + $signed(buffer_0_323); // @[Modules.scala 65:57:@1384.4]
  assign _T_55265 = _T_55264[10:0]; // @[Modules.scala 65:57:@1385.4]
  assign buffer_0_553 = $signed(_T_55265); // @[Modules.scala 65:57:@1386.4]
  assign buffer_0_331 = {{6{io_in_663[4]}},io_in_663}; // @[Modules.scala 32:22:@8.4]
  assign _T_55276 = $signed(11'sh0) + $signed(buffer_0_331); // @[Modules.scala 65:57:@1400.4]
  assign _T_55277 = _T_55276[10:0]; // @[Modules.scala 65:57:@1401.4]
  assign buffer_0_557 = $signed(_T_55277); // @[Modules.scala 65:57:@1402.4]
  assign buffer_0_332 = {{6{_T_54687[4]}},_T_54687}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_333 = {{6{_T_54690[4]}},_T_54690}; // @[Modules.scala 32:22:@8.4]
  assign _T_55279 = $signed(buffer_0_332) + $signed(buffer_0_333); // @[Modules.scala 65:57:@1404.4]
  assign _T_55280 = _T_55279[10:0]; // @[Modules.scala 65:57:@1405.4]
  assign buffer_0_558 = $signed(_T_55280); // @[Modules.scala 65:57:@1406.4]
  assign buffer_0_334 = {{6{_T_54693[4]}},_T_54693}; // @[Modules.scala 32:22:@8.4]
  assign _T_55282 = $signed(buffer_0_334) + $signed(11'sh0); // @[Modules.scala 65:57:@1408.4]
  assign _T_55283 = _T_55282[10:0]; // @[Modules.scala 65:57:@1409.4]
  assign buffer_0_559 = $signed(_T_55283); // @[Modules.scala 65:57:@1410.4]
  assign buffer_0_336 = {{6{io_in_673[4]}},io_in_673}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_337 = {{6{io_in_674[4]}},io_in_674}; // @[Modules.scala 32:22:@8.4]
  assign _T_55285 = $signed(buffer_0_336) + $signed(buffer_0_337); // @[Modules.scala 65:57:@1412.4]
  assign _T_55286 = _T_55285[10:0]; // @[Modules.scala 65:57:@1413.4]
  assign buffer_0_560 = $signed(_T_55286); // @[Modules.scala 65:57:@1414.4]
  assign buffer_0_338 = {{6{_T_54697[4]}},_T_54697}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_339 = {{6{_T_54700[4]}},_T_54700}; // @[Modules.scala 32:22:@8.4]
  assign _T_55288 = $signed(buffer_0_338) + $signed(buffer_0_339); // @[Modules.scala 65:57:@1416.4]
  assign _T_55289 = _T_55288[10:0]; // @[Modules.scala 65:57:@1417.4]
  assign buffer_0_561 = $signed(_T_55289); // @[Modules.scala 65:57:@1418.4]
  assign buffer_0_340 = {{6{_T_54703[4]}},_T_54703}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_341 = {{6{io_in_682[4]}},io_in_682}; // @[Modules.scala 32:22:@8.4]
  assign _T_55291 = $signed(buffer_0_340) + $signed(buffer_0_341); // @[Modules.scala 65:57:@1420.4]
  assign _T_55292 = _T_55291[10:0]; // @[Modules.scala 65:57:@1421.4]
  assign buffer_0_562 = $signed(_T_55292); // @[Modules.scala 65:57:@1422.4]
  assign buffer_0_344 = {{6{_T_54708[4]}},_T_54708}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_345 = {{6{_T_54711[4]}},_T_54711}; // @[Modules.scala 32:22:@8.4]
  assign _T_55297 = $signed(buffer_0_344) + $signed(buffer_0_345); // @[Modules.scala 65:57:@1428.4]
  assign _T_55298 = _T_55297[10:0]; // @[Modules.scala 65:57:@1429.4]
  assign buffer_0_564 = $signed(_T_55298); // @[Modules.scala 65:57:@1430.4]
  assign buffer_0_346 = {{6{_T_54714[4]}},_T_54714}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_347 = {{6{_T_54717[4]}},_T_54717}; // @[Modules.scala 32:22:@8.4]
  assign _T_55300 = $signed(buffer_0_346) + $signed(buffer_0_347); // @[Modules.scala 65:57:@1432.4]
  assign _T_55301 = _T_55300[10:0]; // @[Modules.scala 65:57:@1433.4]
  assign buffer_0_565 = $signed(_T_55301); // @[Modules.scala 65:57:@1434.4]
  assign buffer_0_348 = {{6{_T_54720[4]}},_T_54720}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_349 = {{6{io_in_699[4]}},io_in_699}; // @[Modules.scala 32:22:@8.4]
  assign _T_55303 = $signed(buffer_0_348) + $signed(buffer_0_349); // @[Modules.scala 65:57:@1436.4]
  assign _T_55304 = _T_55303[10:0]; // @[Modules.scala 65:57:@1437.4]
  assign buffer_0_566 = $signed(_T_55304); // @[Modules.scala 65:57:@1438.4]
  assign buffer_0_350 = {{6{io_in_701[4]}},io_in_701}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_351 = {{6{io_in_702[4]}},io_in_702}; // @[Modules.scala 32:22:@8.4]
  assign _T_55306 = $signed(buffer_0_350) + $signed(buffer_0_351); // @[Modules.scala 65:57:@1440.4]
  assign _T_55307 = _T_55306[10:0]; // @[Modules.scala 65:57:@1441.4]
  assign buffer_0_567 = $signed(_T_55307); // @[Modules.scala 65:57:@1442.4]
  assign buffer_0_352 = {{6{_T_54723[4]}},_T_54723}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_353 = {{6{_T_54726[4]}},_T_54726}; // @[Modules.scala 32:22:@8.4]
  assign _T_55309 = $signed(buffer_0_352) + $signed(buffer_0_353); // @[Modules.scala 65:57:@1444.4]
  assign _T_55310 = _T_55309[10:0]; // @[Modules.scala 65:57:@1445.4]
  assign buffer_0_568 = $signed(_T_55310); // @[Modules.scala 65:57:@1446.4]
  assign buffer_0_354 = {{6{_T_54729[4]}},_T_54729}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_355 = {{6{io_in_710[4]}},io_in_710}; // @[Modules.scala 32:22:@8.4]
  assign _T_55312 = $signed(buffer_0_354) + $signed(buffer_0_355); // @[Modules.scala 65:57:@1448.4]
  assign _T_55313 = _T_55312[10:0]; // @[Modules.scala 65:57:@1449.4]
  assign buffer_0_569 = $signed(_T_55313); // @[Modules.scala 65:57:@1450.4]
  assign buffer_0_356 = {{6{_T_54732[4]}},_T_54732}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_357 = {{6{_T_54735[4]}},_T_54735}; // @[Modules.scala 32:22:@8.4]
  assign _T_55315 = $signed(buffer_0_356) + $signed(buffer_0_357); // @[Modules.scala 65:57:@1452.4]
  assign _T_55316 = _T_55315[10:0]; // @[Modules.scala 65:57:@1453.4]
  assign buffer_0_570 = $signed(_T_55316); // @[Modules.scala 65:57:@1454.4]
  assign buffer_0_358 = {{6{_T_54738[4]}},_T_54738}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_359 = {{6{_T_54741[4]}},_T_54741}; // @[Modules.scala 32:22:@8.4]
  assign _T_55318 = $signed(buffer_0_358) + $signed(buffer_0_359); // @[Modules.scala 65:57:@1456.4]
  assign _T_55319 = _T_55318[10:0]; // @[Modules.scala 65:57:@1457.4]
  assign buffer_0_571 = $signed(_T_55319); // @[Modules.scala 65:57:@1458.4]
  assign buffer_0_360 = {{6{_T_54744[4]}},_T_54744}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_361 = {{6{_T_54747[4]}},_T_54747}; // @[Modules.scala 32:22:@8.4]
  assign _T_55321 = $signed(buffer_0_360) + $signed(buffer_0_361); // @[Modules.scala 65:57:@1460.4]
  assign _T_55322 = _T_55321[10:0]; // @[Modules.scala 65:57:@1461.4]
  assign buffer_0_572 = $signed(_T_55322); // @[Modules.scala 65:57:@1462.4]
  assign buffer_0_362 = {{6{io_in_724[4]}},io_in_724}; // @[Modules.scala 32:22:@8.4]
  assign _T_55324 = $signed(buffer_0_362) + $signed(11'sh0); // @[Modules.scala 65:57:@1464.4]
  assign _T_55325 = _T_55324[10:0]; // @[Modules.scala 65:57:@1465.4]
  assign buffer_0_573 = $signed(_T_55325); // @[Modules.scala 65:57:@1466.4]
  assign buffer_0_364 = {{6{io_in_728[4]}},io_in_728}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_365 = {{6{io_in_731[4]}},io_in_731}; // @[Modules.scala 32:22:@8.4]
  assign _T_55327 = $signed(buffer_0_364) + $signed(buffer_0_365); // @[Modules.scala 65:57:@1468.4]
  assign _T_55328 = _T_55327[10:0]; // @[Modules.scala 65:57:@1469.4]
  assign buffer_0_574 = $signed(_T_55328); // @[Modules.scala 65:57:@1470.4]
  assign buffer_0_366 = {{6{_T_54751[4]}},_T_54751}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_367 = {{6{_T_54754[4]}},_T_54754}; // @[Modules.scala 32:22:@8.4]
  assign _T_55330 = $signed(buffer_0_366) + $signed(buffer_0_367); // @[Modules.scala 65:57:@1472.4]
  assign _T_55331 = _T_55330[10:0]; // @[Modules.scala 65:57:@1473.4]
  assign buffer_0_575 = $signed(_T_55331); // @[Modules.scala 65:57:@1474.4]
  assign buffer_0_370 = {{6{io_in_740[4]}},io_in_740}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_371 = {{6{io_in_742[4]}},io_in_742}; // @[Modules.scala 32:22:@8.4]
  assign _T_55336 = $signed(buffer_0_370) + $signed(buffer_0_371); // @[Modules.scala 65:57:@1480.4]
  assign _T_55337 = _T_55336[10:0]; // @[Modules.scala 65:57:@1481.4]
  assign buffer_0_577 = $signed(_T_55337); // @[Modules.scala 65:57:@1482.4]
  assign buffer_0_374 = {{6{_T_54761[4]}},_T_54761}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_375 = {{6{io_in_750[4]}},io_in_750}; // @[Modules.scala 32:22:@8.4]
  assign _T_55342 = $signed(buffer_0_374) + $signed(buffer_0_375); // @[Modules.scala 65:57:@1488.4]
  assign _T_55343 = _T_55342[10:0]; // @[Modules.scala 65:57:@1489.4]
  assign buffer_0_579 = $signed(_T_55343); // @[Modules.scala 65:57:@1490.4]
  assign buffer_0_376 = {{6{_T_54764[4]}},_T_54764}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_377 = {{6{_T_54767[4]}},_T_54767}; // @[Modules.scala 32:22:@8.4]
  assign _T_55345 = $signed(buffer_0_376) + $signed(buffer_0_377); // @[Modules.scala 65:57:@1492.4]
  assign _T_55346 = _T_55345[10:0]; // @[Modules.scala 65:57:@1493.4]
  assign buffer_0_580 = $signed(_T_55346); // @[Modules.scala 65:57:@1494.4]
  assign buffer_0_378 = {{6{io_in_757[4]}},io_in_757}; // @[Modules.scala 32:22:@8.4]
  assign _T_55348 = $signed(buffer_0_378) + $signed(11'sh0); // @[Modules.scala 65:57:@1496.4]
  assign _T_55349 = _T_55348[10:0]; // @[Modules.scala 65:57:@1497.4]
  assign buffer_0_581 = $signed(_T_55349); // @[Modules.scala 65:57:@1498.4]
  assign buffer_0_380 = {{6{io_in_760[4]}},io_in_760}; // @[Modules.scala 32:22:@8.4]
  assign _T_55351 = $signed(buffer_0_380) + $signed(11'sh0); // @[Modules.scala 65:57:@1500.4]
  assign _T_55352 = _T_55351[10:0]; // @[Modules.scala 65:57:@1501.4]
  assign buffer_0_582 = $signed(_T_55352); // @[Modules.scala 65:57:@1502.4]
  assign buffer_0_384 = {{6{io_in_768[4]}},io_in_768}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_385 = {{6{io_in_771[4]}},io_in_771}; // @[Modules.scala 32:22:@8.4]
  assign _T_55357 = $signed(buffer_0_384) + $signed(buffer_0_385); // @[Modules.scala 65:57:@1508.4]
  assign _T_55358 = _T_55357[10:0]; // @[Modules.scala 65:57:@1509.4]
  assign buffer_0_584 = $signed(_T_55358); // @[Modules.scala 65:57:@1510.4]
  assign buffer_0_388 = {{6{_T_54776[4]}},_T_54776}; // @[Modules.scala 32:22:@8.4]
  assign _T_55363 = $signed(buffer_0_388) + $signed(11'sh0); // @[Modules.scala 65:57:@1516.4]
  assign _T_55364 = _T_55363[10:0]; // @[Modules.scala 65:57:@1517.4]
  assign buffer_0_586 = $signed(_T_55364); // @[Modules.scala 65:57:@1518.4]
  assign buffer_0_390 = {{6{io_in_781[4]}},io_in_781}; // @[Modules.scala 32:22:@8.4]
  assign buffer_0_391 = {{6{_T_54780[4]}},_T_54780}; // @[Modules.scala 32:22:@8.4]
  assign _T_55366 = $signed(buffer_0_390) + $signed(buffer_0_391); // @[Modules.scala 65:57:@1520.4]
  assign _T_55367 = _T_55366[10:0]; // @[Modules.scala 65:57:@1521.4]
  assign buffer_0_587 = $signed(_T_55367); // @[Modules.scala 65:57:@1522.4]
  assign _T_55369 = $signed(buffer_0_392) + $signed(buffer_0_393); // @[Modules.scala 68:83:@1524.4]
  assign _T_55370 = _T_55369[10:0]; // @[Modules.scala 68:83:@1525.4]
  assign buffer_0_588 = $signed(_T_55370); // @[Modules.scala 68:83:@1526.4]
  assign _T_55372 = $signed(buffer_0_394) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1528.4]
  assign _T_55373 = _T_55372[10:0]; // @[Modules.scala 68:83:@1529.4]
  assign buffer_0_589 = $signed(_T_55373); // @[Modules.scala 68:83:@1530.4]
  assign _T_55375 = $signed(buffer_0_396) + $signed(buffer_0_397); // @[Modules.scala 68:83:@1532.4]
  assign _T_55376 = _T_55375[10:0]; // @[Modules.scala 68:83:@1533.4]
  assign buffer_0_590 = $signed(_T_55376); // @[Modules.scala 68:83:@1534.4]
  assign _T_55378 = $signed(buffer_0_398) + $signed(buffer_0_399); // @[Modules.scala 68:83:@1536.4]
  assign _T_55379 = _T_55378[10:0]; // @[Modules.scala 68:83:@1537.4]
  assign buffer_0_591 = $signed(_T_55379); // @[Modules.scala 68:83:@1538.4]
  assign _T_55381 = $signed(buffer_0_400) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1540.4]
  assign _T_55382 = _T_55381[10:0]; // @[Modules.scala 68:83:@1541.4]
  assign buffer_0_592 = $signed(_T_55382); // @[Modules.scala 68:83:@1542.4]
  assign _T_55384 = $signed(buffer_0_395) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1544.4]
  assign _T_55385 = _T_55384[10:0]; // @[Modules.scala 68:83:@1545.4]
  assign buffer_0_593 = $signed(_T_55385); // @[Modules.scala 68:83:@1546.4]
  assign _T_55387 = $signed(buffer_0_395) + $signed(buffer_0_405); // @[Modules.scala 68:83:@1548.4]
  assign _T_55388 = _T_55387[10:0]; // @[Modules.scala 68:83:@1549.4]
  assign buffer_0_594 = $signed(_T_55388); // @[Modules.scala 68:83:@1550.4]
  assign _T_55390 = $signed(buffer_0_406) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1552.4]
  assign _T_55391 = _T_55390[10:0]; // @[Modules.scala 68:83:@1553.4]
  assign buffer_0_595 = $signed(_T_55391); // @[Modules.scala 68:83:@1554.4]
  assign _T_55393 = $signed(buffer_0_408) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1556.4]
  assign _T_55394 = _T_55393[10:0]; // @[Modules.scala 68:83:@1557.4]
  assign buffer_0_596 = $signed(_T_55394); // @[Modules.scala 68:83:@1558.4]
  assign _T_55396 = $signed(buffer_0_410) + $signed(buffer_0_411); // @[Modules.scala 68:83:@1560.4]
  assign _T_55397 = _T_55396[10:0]; // @[Modules.scala 68:83:@1561.4]
  assign buffer_0_597 = $signed(_T_55397); // @[Modules.scala 68:83:@1562.4]
  assign _T_55399 = $signed(buffer_0_412) + $signed(buffer_0_413); // @[Modules.scala 68:83:@1564.4]
  assign _T_55400 = _T_55399[10:0]; // @[Modules.scala 68:83:@1565.4]
  assign buffer_0_598 = $signed(_T_55400); // @[Modules.scala 68:83:@1566.4]
  assign _T_55402 = $signed(buffer_0_414) + $signed(buffer_0_415); // @[Modules.scala 68:83:@1568.4]
  assign _T_55403 = _T_55402[10:0]; // @[Modules.scala 68:83:@1569.4]
  assign buffer_0_599 = $signed(_T_55403); // @[Modules.scala 68:83:@1570.4]
  assign _T_55405 = $signed(buffer_0_416) + $signed(buffer_0_417); // @[Modules.scala 68:83:@1572.4]
  assign _T_55406 = _T_55405[10:0]; // @[Modules.scala 68:83:@1573.4]
  assign buffer_0_600 = $signed(_T_55406); // @[Modules.scala 68:83:@1574.4]
  assign _T_55408 = $signed(buffer_0_418) + $signed(buffer_0_419); // @[Modules.scala 68:83:@1576.4]
  assign _T_55409 = _T_55408[10:0]; // @[Modules.scala 68:83:@1577.4]
  assign buffer_0_601 = $signed(_T_55409); // @[Modules.scala 68:83:@1578.4]
  assign _T_55411 = $signed(buffer_0_420) + $signed(buffer_0_421); // @[Modules.scala 68:83:@1580.4]
  assign _T_55412 = _T_55411[10:0]; // @[Modules.scala 68:83:@1581.4]
  assign buffer_0_602 = $signed(_T_55412); // @[Modules.scala 68:83:@1582.4]
  assign _T_55417 = $signed(buffer_0_424) + $signed(buffer_0_425); // @[Modules.scala 68:83:@1588.4]
  assign _T_55418 = _T_55417[10:0]; // @[Modules.scala 68:83:@1589.4]
  assign buffer_0_604 = $signed(_T_55418); // @[Modules.scala 68:83:@1590.4]
  assign _T_55420 = $signed(buffer_0_426) + $signed(buffer_0_427); // @[Modules.scala 68:83:@1592.4]
  assign _T_55421 = _T_55420[10:0]; // @[Modules.scala 68:83:@1593.4]
  assign buffer_0_605 = $signed(_T_55421); // @[Modules.scala 68:83:@1594.4]
  assign _T_55423 = $signed(buffer_0_428) + $signed(buffer_0_429); // @[Modules.scala 68:83:@1596.4]
  assign _T_55424 = _T_55423[10:0]; // @[Modules.scala 68:83:@1597.4]
  assign buffer_0_606 = $signed(_T_55424); // @[Modules.scala 68:83:@1598.4]
  assign _T_55429 = $signed(buffer_0_432) + $signed(buffer_0_433); // @[Modules.scala 68:83:@1604.4]
  assign _T_55430 = _T_55429[10:0]; // @[Modules.scala 68:83:@1605.4]
  assign buffer_0_608 = $signed(_T_55430); // @[Modules.scala 68:83:@1606.4]
  assign _T_55432 = $signed(buffer_0_395) + $signed(buffer_0_435); // @[Modules.scala 68:83:@1608.4]
  assign _T_55433 = _T_55432[10:0]; // @[Modules.scala 68:83:@1609.4]
  assign buffer_0_609 = $signed(_T_55433); // @[Modules.scala 68:83:@1610.4]
  assign _T_55438 = $signed(buffer_0_438) + $signed(buffer_0_439); // @[Modules.scala 68:83:@1616.4]
  assign _T_55439 = _T_55438[10:0]; // @[Modules.scala 68:83:@1617.4]
  assign buffer_0_611 = $signed(_T_55439); // @[Modules.scala 68:83:@1618.4]
  assign _T_55441 = $signed(buffer_0_395) + $signed(buffer_0_441); // @[Modules.scala 68:83:@1620.4]
  assign _T_55442 = _T_55441[10:0]; // @[Modules.scala 68:83:@1621.4]
  assign buffer_0_612 = $signed(_T_55442); // @[Modules.scala 68:83:@1622.4]
  assign _T_55444 = $signed(buffer_0_395) + $signed(buffer_0_443); // @[Modules.scala 68:83:@1624.4]
  assign _T_55445 = _T_55444[10:0]; // @[Modules.scala 68:83:@1625.4]
  assign buffer_0_613 = $signed(_T_55445); // @[Modules.scala 68:83:@1626.4]
  assign _T_55447 = $signed(buffer_0_444) + $signed(buffer_0_445); // @[Modules.scala 68:83:@1628.4]
  assign _T_55448 = _T_55447[10:0]; // @[Modules.scala 68:83:@1629.4]
  assign buffer_0_614 = $signed(_T_55448); // @[Modules.scala 68:83:@1630.4]
  assign _T_55456 = $signed(buffer_0_395) + $signed(buffer_0_451); // @[Modules.scala 68:83:@1640.4]
  assign _T_55457 = _T_55456[10:0]; // @[Modules.scala 68:83:@1641.4]
  assign buffer_0_617 = $signed(_T_55457); // @[Modules.scala 68:83:@1642.4]
  assign _T_55465 = $signed(buffer_0_395) + $signed(buffer_0_457); // @[Modules.scala 68:83:@1652.4]
  assign _T_55466 = _T_55465[10:0]; // @[Modules.scala 68:83:@1653.4]
  assign buffer_0_620 = $signed(_T_55466); // @[Modules.scala 68:83:@1654.4]
  assign _T_55477 = $signed(buffer_0_464) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1668.4]
  assign _T_55478 = _T_55477[10:0]; // @[Modules.scala 68:83:@1669.4]
  assign buffer_0_624 = $signed(_T_55478); // @[Modules.scala 68:83:@1670.4]
  assign _T_55486 = $signed(buffer_0_470) + $signed(buffer_0_471); // @[Modules.scala 68:83:@1680.4]
  assign _T_55487 = _T_55486[10:0]; // @[Modules.scala 68:83:@1681.4]
  assign buffer_0_627 = $signed(_T_55487); // @[Modules.scala 68:83:@1682.4]
  assign _T_55489 = $signed(buffer_0_395) + $signed(buffer_0_473); // @[Modules.scala 68:83:@1684.4]
  assign _T_55490 = _T_55489[10:0]; // @[Modules.scala 68:83:@1685.4]
  assign buffer_0_628 = $signed(_T_55490); // @[Modules.scala 68:83:@1686.4]
  assign _T_55492 = $signed(buffer_0_474) + $signed(buffer_0_475); // @[Modules.scala 68:83:@1688.4]
  assign _T_55493 = _T_55492[10:0]; // @[Modules.scala 68:83:@1689.4]
  assign buffer_0_629 = $signed(_T_55493); // @[Modules.scala 68:83:@1690.4]
  assign _T_55495 = $signed(buffer_0_476) + $signed(buffer_0_477); // @[Modules.scala 68:83:@1692.4]
  assign _T_55496 = _T_55495[10:0]; // @[Modules.scala 68:83:@1693.4]
  assign buffer_0_630 = $signed(_T_55496); // @[Modules.scala 68:83:@1694.4]
  assign _T_55498 = $signed(buffer_0_478) + $signed(buffer_0_479); // @[Modules.scala 68:83:@1696.4]
  assign _T_55499 = _T_55498[10:0]; // @[Modules.scala 68:83:@1697.4]
  assign buffer_0_631 = $signed(_T_55499); // @[Modules.scala 68:83:@1698.4]
  assign _T_55501 = $signed(buffer_0_480) + $signed(buffer_0_481); // @[Modules.scala 68:83:@1700.4]
  assign _T_55502 = _T_55501[10:0]; // @[Modules.scala 68:83:@1701.4]
  assign buffer_0_632 = $signed(_T_55502); // @[Modules.scala 68:83:@1702.4]
  assign _T_55504 = $signed(buffer_0_482) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1704.4]
  assign _T_55505 = _T_55504[10:0]; // @[Modules.scala 68:83:@1705.4]
  assign buffer_0_633 = $signed(_T_55505); // @[Modules.scala 68:83:@1706.4]
  assign _T_55507 = $signed(buffer_0_484) + $signed(buffer_0_485); // @[Modules.scala 68:83:@1708.4]
  assign _T_55508 = _T_55507[10:0]; // @[Modules.scala 68:83:@1709.4]
  assign buffer_0_634 = $signed(_T_55508); // @[Modules.scala 68:83:@1710.4]
  assign _T_55510 = $signed(buffer_0_486) + $signed(buffer_0_487); // @[Modules.scala 68:83:@1712.4]
  assign _T_55511 = _T_55510[10:0]; // @[Modules.scala 68:83:@1713.4]
  assign buffer_0_635 = $signed(_T_55511); // @[Modules.scala 68:83:@1714.4]
  assign _T_55513 = $signed(buffer_0_488) + $signed(buffer_0_489); // @[Modules.scala 68:83:@1716.4]
  assign _T_55514 = _T_55513[10:0]; // @[Modules.scala 68:83:@1717.4]
  assign buffer_0_636 = $signed(_T_55514); // @[Modules.scala 68:83:@1718.4]
  assign _T_55516 = $signed(buffer_0_395) + $signed(buffer_0_491); // @[Modules.scala 68:83:@1720.4]
  assign _T_55517 = _T_55516[10:0]; // @[Modules.scala 68:83:@1721.4]
  assign buffer_0_637 = $signed(_T_55517); // @[Modules.scala 68:83:@1722.4]
  assign _T_55519 = $signed(buffer_0_492) + $signed(buffer_0_493); // @[Modules.scala 68:83:@1724.4]
  assign _T_55520 = _T_55519[10:0]; // @[Modules.scala 68:83:@1725.4]
  assign buffer_0_638 = $signed(_T_55520); // @[Modules.scala 68:83:@1726.4]
  assign _T_55522 = $signed(buffer_0_494) + $signed(buffer_0_495); // @[Modules.scala 68:83:@1728.4]
  assign _T_55523 = _T_55522[10:0]; // @[Modules.scala 68:83:@1729.4]
  assign buffer_0_639 = $signed(_T_55523); // @[Modules.scala 68:83:@1730.4]
  assign _T_55525 = $signed(buffer_0_496) + $signed(buffer_0_497); // @[Modules.scala 68:83:@1732.4]
  assign _T_55526 = _T_55525[10:0]; // @[Modules.scala 68:83:@1733.4]
  assign buffer_0_640 = $signed(_T_55526); // @[Modules.scala 68:83:@1734.4]
  assign _T_55528 = $signed(buffer_0_498) + $signed(buffer_0_499); // @[Modules.scala 68:83:@1736.4]
  assign _T_55529 = _T_55528[10:0]; // @[Modules.scala 68:83:@1737.4]
  assign buffer_0_641 = $signed(_T_55529); // @[Modules.scala 68:83:@1738.4]
  assign _T_55531 = $signed(buffer_0_500) + $signed(buffer_0_501); // @[Modules.scala 68:83:@1740.4]
  assign _T_55532 = _T_55531[10:0]; // @[Modules.scala 68:83:@1741.4]
  assign buffer_0_642 = $signed(_T_55532); // @[Modules.scala 68:83:@1742.4]
  assign _T_55534 = $signed(buffer_0_502) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1744.4]
  assign _T_55535 = _T_55534[10:0]; // @[Modules.scala 68:83:@1745.4]
  assign buffer_0_643 = $signed(_T_55535); // @[Modules.scala 68:83:@1746.4]
  assign _T_55537 = $signed(buffer_0_504) + $signed(buffer_0_505); // @[Modules.scala 68:83:@1748.4]
  assign _T_55538 = _T_55537[10:0]; // @[Modules.scala 68:83:@1749.4]
  assign buffer_0_644 = $signed(_T_55538); // @[Modules.scala 68:83:@1750.4]
  assign _T_55540 = $signed(buffer_0_506) + $signed(buffer_0_507); // @[Modules.scala 68:83:@1752.4]
  assign _T_55541 = _T_55540[10:0]; // @[Modules.scala 68:83:@1753.4]
  assign buffer_0_645 = $signed(_T_55541); // @[Modules.scala 68:83:@1754.4]
  assign _T_55543 = $signed(buffer_0_508) + $signed(buffer_0_509); // @[Modules.scala 68:83:@1756.4]
  assign _T_55544 = _T_55543[10:0]; // @[Modules.scala 68:83:@1757.4]
  assign buffer_0_646 = $signed(_T_55544); // @[Modules.scala 68:83:@1758.4]
  assign _T_55546 = $signed(buffer_0_395) + $signed(buffer_0_511); // @[Modules.scala 68:83:@1760.4]
  assign _T_55547 = _T_55546[10:0]; // @[Modules.scala 68:83:@1761.4]
  assign buffer_0_647 = $signed(_T_55547); // @[Modules.scala 68:83:@1762.4]
  assign _T_55549 = $signed(buffer_0_512) + $signed(buffer_0_513); // @[Modules.scala 68:83:@1764.4]
  assign _T_55550 = _T_55549[10:0]; // @[Modules.scala 68:83:@1765.4]
  assign buffer_0_648 = $signed(_T_55550); // @[Modules.scala 68:83:@1766.4]
  assign _T_55552 = $signed(buffer_0_514) + $signed(buffer_0_515); // @[Modules.scala 68:83:@1768.4]
  assign _T_55553 = _T_55552[10:0]; // @[Modules.scala 68:83:@1769.4]
  assign buffer_0_649 = $signed(_T_55553); // @[Modules.scala 68:83:@1770.4]
  assign _T_55555 = $signed(buffer_0_516) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1772.4]
  assign _T_55556 = _T_55555[10:0]; // @[Modules.scala 68:83:@1773.4]
  assign buffer_0_650 = $signed(_T_55556); // @[Modules.scala 68:83:@1774.4]
  assign _T_55558 = $signed(buffer_0_518) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1776.4]
  assign _T_55559 = _T_55558[10:0]; // @[Modules.scala 68:83:@1777.4]
  assign buffer_0_651 = $signed(_T_55559); // @[Modules.scala 68:83:@1778.4]
  assign _T_55561 = $signed(buffer_0_520) + $signed(buffer_0_521); // @[Modules.scala 68:83:@1780.4]
  assign _T_55562 = _T_55561[10:0]; // @[Modules.scala 68:83:@1781.4]
  assign buffer_0_652 = $signed(_T_55562); // @[Modules.scala 68:83:@1782.4]
  assign _T_55564 = $signed(buffer_0_522) + $signed(buffer_0_523); // @[Modules.scala 68:83:@1784.4]
  assign _T_55565 = _T_55564[10:0]; // @[Modules.scala 68:83:@1785.4]
  assign buffer_0_653 = $signed(_T_55565); // @[Modules.scala 68:83:@1786.4]
  assign _T_55567 = $signed(buffer_0_524) + $signed(buffer_0_525); // @[Modules.scala 68:83:@1788.4]
  assign _T_55568 = _T_55567[10:0]; // @[Modules.scala 68:83:@1789.4]
  assign buffer_0_654 = $signed(_T_55568); // @[Modules.scala 68:83:@1790.4]
  assign _T_55570 = $signed(buffer_0_395) + $signed(buffer_0_527); // @[Modules.scala 68:83:@1792.4]
  assign _T_55571 = _T_55570[10:0]; // @[Modules.scala 68:83:@1793.4]
  assign buffer_0_655 = $signed(_T_55571); // @[Modules.scala 68:83:@1794.4]
  assign _T_55573 = $signed(buffer_0_395) + $signed(buffer_0_529); // @[Modules.scala 68:83:@1796.4]
  assign _T_55574 = _T_55573[10:0]; // @[Modules.scala 68:83:@1797.4]
  assign buffer_0_656 = $signed(_T_55574); // @[Modules.scala 68:83:@1798.4]
  assign _T_55576 = $signed(buffer_0_530) + $signed(buffer_0_531); // @[Modules.scala 68:83:@1800.4]
  assign _T_55577 = _T_55576[10:0]; // @[Modules.scala 68:83:@1801.4]
  assign buffer_0_657 = $signed(_T_55577); // @[Modules.scala 68:83:@1802.4]
  assign _T_55582 = $signed(buffer_0_534) + $signed(buffer_0_535); // @[Modules.scala 68:83:@1808.4]
  assign _T_55583 = _T_55582[10:0]; // @[Modules.scala 68:83:@1809.4]
  assign buffer_0_659 = $signed(_T_55583); // @[Modules.scala 68:83:@1810.4]
  assign _T_55585 = $signed(buffer_0_536) + $signed(buffer_0_537); // @[Modules.scala 68:83:@1812.4]
  assign _T_55586 = _T_55585[10:0]; // @[Modules.scala 68:83:@1813.4]
  assign buffer_0_660 = $signed(_T_55586); // @[Modules.scala 68:83:@1814.4]
  assign _T_55588 = $signed(buffer_0_538) + $signed(buffer_0_539); // @[Modules.scala 68:83:@1816.4]
  assign _T_55589 = _T_55588[10:0]; // @[Modules.scala 68:83:@1817.4]
  assign buffer_0_661 = $signed(_T_55589); // @[Modules.scala 68:83:@1818.4]
  assign _T_55594 = $signed(buffer_0_542) + $signed(buffer_0_543); // @[Modules.scala 68:83:@1824.4]
  assign _T_55595 = _T_55594[10:0]; // @[Modules.scala 68:83:@1825.4]
  assign buffer_0_663 = $signed(_T_55595); // @[Modules.scala 68:83:@1826.4]
  assign _T_55597 = $signed(buffer_0_395) + $signed(buffer_0_545); // @[Modules.scala 68:83:@1828.4]
  assign _T_55598 = _T_55597[10:0]; // @[Modules.scala 68:83:@1829.4]
  assign buffer_0_664 = $signed(_T_55598); // @[Modules.scala 68:83:@1830.4]
  assign _T_55600 = $signed(buffer_0_546) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1832.4]
  assign _T_55601 = _T_55600[10:0]; // @[Modules.scala 68:83:@1833.4]
  assign buffer_0_665 = $signed(_T_55601); // @[Modules.scala 68:83:@1834.4]
  assign _T_55606 = $signed(buffer_0_395) + $signed(buffer_0_551); // @[Modules.scala 68:83:@1840.4]
  assign _T_55607 = _T_55606[10:0]; // @[Modules.scala 68:83:@1841.4]
  assign buffer_0_667 = $signed(_T_55607); // @[Modules.scala 68:83:@1842.4]
  assign _T_55609 = $signed(buffer_0_552) + $signed(buffer_0_553); // @[Modules.scala 68:83:@1844.4]
  assign _T_55610 = _T_55609[10:0]; // @[Modules.scala 68:83:@1845.4]
  assign buffer_0_668 = $signed(_T_55610); // @[Modules.scala 68:83:@1846.4]
  assign _T_55615 = $signed(buffer_0_395) + $signed(buffer_0_557); // @[Modules.scala 68:83:@1852.4]
  assign _T_55616 = _T_55615[10:0]; // @[Modules.scala 68:83:@1853.4]
  assign buffer_0_670 = $signed(_T_55616); // @[Modules.scala 68:83:@1854.4]
  assign _T_55618 = $signed(buffer_0_558) + $signed(buffer_0_559); // @[Modules.scala 68:83:@1856.4]
  assign _T_55619 = _T_55618[10:0]; // @[Modules.scala 68:83:@1857.4]
  assign buffer_0_671 = $signed(_T_55619); // @[Modules.scala 68:83:@1858.4]
  assign _T_55621 = $signed(buffer_0_560) + $signed(buffer_0_561); // @[Modules.scala 68:83:@1860.4]
  assign _T_55622 = _T_55621[10:0]; // @[Modules.scala 68:83:@1861.4]
  assign buffer_0_672 = $signed(_T_55622); // @[Modules.scala 68:83:@1862.4]
  assign _T_55624 = $signed(buffer_0_562) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1864.4]
  assign _T_55625 = _T_55624[10:0]; // @[Modules.scala 68:83:@1865.4]
  assign buffer_0_673 = $signed(_T_55625); // @[Modules.scala 68:83:@1866.4]
  assign _T_55627 = $signed(buffer_0_564) + $signed(buffer_0_565); // @[Modules.scala 68:83:@1868.4]
  assign _T_55628 = _T_55627[10:0]; // @[Modules.scala 68:83:@1869.4]
  assign buffer_0_674 = $signed(_T_55628); // @[Modules.scala 68:83:@1870.4]
  assign _T_55630 = $signed(buffer_0_566) + $signed(buffer_0_567); // @[Modules.scala 68:83:@1872.4]
  assign _T_55631 = _T_55630[10:0]; // @[Modules.scala 68:83:@1873.4]
  assign buffer_0_675 = $signed(_T_55631); // @[Modules.scala 68:83:@1874.4]
  assign _T_55633 = $signed(buffer_0_568) + $signed(buffer_0_569); // @[Modules.scala 68:83:@1876.4]
  assign _T_55634 = _T_55633[10:0]; // @[Modules.scala 68:83:@1877.4]
  assign buffer_0_676 = $signed(_T_55634); // @[Modules.scala 68:83:@1878.4]
  assign _T_55636 = $signed(buffer_0_570) + $signed(buffer_0_571); // @[Modules.scala 68:83:@1880.4]
  assign _T_55637 = _T_55636[10:0]; // @[Modules.scala 68:83:@1881.4]
  assign buffer_0_677 = $signed(_T_55637); // @[Modules.scala 68:83:@1882.4]
  assign _T_55639 = $signed(buffer_0_572) + $signed(buffer_0_573); // @[Modules.scala 68:83:@1884.4]
  assign _T_55640 = _T_55639[10:0]; // @[Modules.scala 68:83:@1885.4]
  assign buffer_0_678 = $signed(_T_55640); // @[Modules.scala 68:83:@1886.4]
  assign _T_55642 = $signed(buffer_0_574) + $signed(buffer_0_575); // @[Modules.scala 68:83:@1888.4]
  assign _T_55643 = _T_55642[10:0]; // @[Modules.scala 68:83:@1889.4]
  assign buffer_0_679 = $signed(_T_55643); // @[Modules.scala 68:83:@1890.4]
  assign _T_55645 = $signed(buffer_0_395) + $signed(buffer_0_577); // @[Modules.scala 68:83:@1892.4]
  assign _T_55646 = _T_55645[10:0]; // @[Modules.scala 68:83:@1893.4]
  assign buffer_0_680 = $signed(_T_55646); // @[Modules.scala 68:83:@1894.4]
  assign _T_55648 = $signed(buffer_0_395) + $signed(buffer_0_579); // @[Modules.scala 68:83:@1896.4]
  assign _T_55649 = _T_55648[10:0]; // @[Modules.scala 68:83:@1897.4]
  assign buffer_0_681 = $signed(_T_55649); // @[Modules.scala 68:83:@1898.4]
  assign _T_55651 = $signed(buffer_0_580) + $signed(buffer_0_581); // @[Modules.scala 68:83:@1900.4]
  assign _T_55652 = _T_55651[10:0]; // @[Modules.scala 68:83:@1901.4]
  assign buffer_0_682 = $signed(_T_55652); // @[Modules.scala 68:83:@1902.4]
  assign _T_55654 = $signed(buffer_0_582) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1904.4]
  assign _T_55655 = _T_55654[10:0]; // @[Modules.scala 68:83:@1905.4]
  assign buffer_0_683 = $signed(_T_55655); // @[Modules.scala 68:83:@1906.4]
  assign _T_55657 = $signed(buffer_0_584) + $signed(buffer_0_395); // @[Modules.scala 68:83:@1908.4]
  assign _T_55658 = _T_55657[10:0]; // @[Modules.scala 68:83:@1909.4]
  assign buffer_0_684 = $signed(_T_55658); // @[Modules.scala 68:83:@1910.4]
  assign _T_55660 = $signed(buffer_0_586) + $signed(buffer_0_587); // @[Modules.scala 68:83:@1912.4]
  assign _T_55661 = _T_55660[10:0]; // @[Modules.scala 68:83:@1913.4]
  assign buffer_0_685 = $signed(_T_55661); // @[Modules.scala 68:83:@1914.4]
  assign _T_55663 = $signed(buffer_0_588) + $signed(buffer_0_589); // @[Modules.scala 71:109:@1916.4]
  assign _T_55664 = _T_55663[10:0]; // @[Modules.scala 71:109:@1917.4]
  assign buffer_0_686 = $signed(_T_55664); // @[Modules.scala 71:109:@1918.4]
  assign _T_55666 = $signed(buffer_0_590) + $signed(buffer_0_591); // @[Modules.scala 71:109:@1920.4]
  assign _T_55667 = _T_55666[10:0]; // @[Modules.scala 71:109:@1921.4]
  assign buffer_0_687 = $signed(_T_55667); // @[Modules.scala 71:109:@1922.4]
  assign _T_55669 = $signed(buffer_0_592) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1924.4]
  assign _T_55670 = _T_55669[10:0]; // @[Modules.scala 71:109:@1925.4]
  assign buffer_0_688 = $signed(_T_55670); // @[Modules.scala 71:109:@1926.4]
  assign _T_55672 = $signed(buffer_0_594) + $signed(buffer_0_595); // @[Modules.scala 71:109:@1928.4]
  assign _T_55673 = _T_55672[10:0]; // @[Modules.scala 71:109:@1929.4]
  assign buffer_0_689 = $signed(_T_55673); // @[Modules.scala 71:109:@1930.4]
  assign _T_55675 = $signed(buffer_0_596) + $signed(buffer_0_597); // @[Modules.scala 71:109:@1932.4]
  assign _T_55676 = _T_55675[10:0]; // @[Modules.scala 71:109:@1933.4]
  assign buffer_0_690 = $signed(_T_55676); // @[Modules.scala 71:109:@1934.4]
  assign _T_55678 = $signed(buffer_0_598) + $signed(buffer_0_599); // @[Modules.scala 71:109:@1936.4]
  assign _T_55679 = _T_55678[10:0]; // @[Modules.scala 71:109:@1937.4]
  assign buffer_0_691 = $signed(_T_55679); // @[Modules.scala 71:109:@1938.4]
  assign _T_55681 = $signed(buffer_0_600) + $signed(buffer_0_601); // @[Modules.scala 71:109:@1940.4]
  assign _T_55682 = _T_55681[10:0]; // @[Modules.scala 71:109:@1941.4]
  assign buffer_0_692 = $signed(_T_55682); // @[Modules.scala 71:109:@1942.4]
  assign _T_55684 = $signed(buffer_0_602) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1944.4]
  assign _T_55685 = _T_55684[10:0]; // @[Modules.scala 71:109:@1945.4]
  assign buffer_0_693 = $signed(_T_55685); // @[Modules.scala 71:109:@1946.4]
  assign _T_55687 = $signed(buffer_0_604) + $signed(buffer_0_605); // @[Modules.scala 71:109:@1948.4]
  assign _T_55688 = _T_55687[10:0]; // @[Modules.scala 71:109:@1949.4]
  assign buffer_0_694 = $signed(_T_55688); // @[Modules.scala 71:109:@1950.4]
  assign _T_55690 = $signed(buffer_0_606) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1952.4]
  assign _T_55691 = _T_55690[10:0]; // @[Modules.scala 71:109:@1953.4]
  assign buffer_0_695 = $signed(_T_55691); // @[Modules.scala 71:109:@1954.4]
  assign _T_55693 = $signed(buffer_0_608) + $signed(buffer_0_609); // @[Modules.scala 71:109:@1956.4]
  assign _T_55694 = _T_55693[10:0]; // @[Modules.scala 71:109:@1957.4]
  assign buffer_0_696 = $signed(_T_55694); // @[Modules.scala 71:109:@1958.4]
  assign _T_55696 = $signed(buffer_0_593) + $signed(buffer_0_611); // @[Modules.scala 71:109:@1960.4]
  assign _T_55697 = _T_55696[10:0]; // @[Modules.scala 71:109:@1961.4]
  assign buffer_0_697 = $signed(_T_55697); // @[Modules.scala 71:109:@1962.4]
  assign _T_55699 = $signed(buffer_0_612) + $signed(buffer_0_613); // @[Modules.scala 71:109:@1964.4]
  assign _T_55700 = _T_55699[10:0]; // @[Modules.scala 71:109:@1965.4]
  assign buffer_0_698 = $signed(_T_55700); // @[Modules.scala 71:109:@1966.4]
  assign _T_55702 = $signed(buffer_0_614) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1968.4]
  assign _T_55703 = _T_55702[10:0]; // @[Modules.scala 71:109:@1969.4]
  assign buffer_0_699 = $signed(_T_55703); // @[Modules.scala 71:109:@1970.4]
  assign _T_55705 = $signed(buffer_0_593) + $signed(buffer_0_617); // @[Modules.scala 71:109:@1972.4]
  assign _T_55706 = _T_55705[10:0]; // @[Modules.scala 71:109:@1973.4]
  assign buffer_0_700 = $signed(_T_55706); // @[Modules.scala 71:109:@1974.4]
  assign _T_55708 = $signed(buffer_0_593) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1976.4]
  assign _T_55709 = _T_55708[10:0]; // @[Modules.scala 71:109:@1977.4]
  assign buffer_0_701 = $signed(_T_55709); // @[Modules.scala 71:109:@1978.4]
  assign _T_55711 = $signed(buffer_0_620) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1980.4]
  assign _T_55712 = _T_55711[10:0]; // @[Modules.scala 71:109:@1981.4]
  assign buffer_0_702 = $signed(_T_55712); // @[Modules.scala 71:109:@1982.4]
  assign _T_55717 = $signed(buffer_0_624) + $signed(buffer_0_593); // @[Modules.scala 71:109:@1988.4]
  assign _T_55718 = _T_55717[10:0]; // @[Modules.scala 71:109:@1989.4]
  assign buffer_0_704 = $signed(_T_55718); // @[Modules.scala 71:109:@1990.4]
  assign _T_55720 = $signed(buffer_0_593) + $signed(buffer_0_627); // @[Modules.scala 71:109:@1992.4]
  assign _T_55721 = _T_55720[10:0]; // @[Modules.scala 71:109:@1993.4]
  assign buffer_0_705 = $signed(_T_55721); // @[Modules.scala 71:109:@1994.4]
  assign _T_55723 = $signed(buffer_0_628) + $signed(buffer_0_629); // @[Modules.scala 71:109:@1996.4]
  assign _T_55724 = _T_55723[10:0]; // @[Modules.scala 71:109:@1997.4]
  assign buffer_0_706 = $signed(_T_55724); // @[Modules.scala 71:109:@1998.4]
  assign _T_55726 = $signed(buffer_0_630) + $signed(buffer_0_631); // @[Modules.scala 71:109:@2000.4]
  assign _T_55727 = _T_55726[10:0]; // @[Modules.scala 71:109:@2001.4]
  assign buffer_0_707 = $signed(_T_55727); // @[Modules.scala 71:109:@2002.4]
  assign _T_55729 = $signed(buffer_0_632) + $signed(buffer_0_633); // @[Modules.scala 71:109:@2004.4]
  assign _T_55730 = _T_55729[10:0]; // @[Modules.scala 71:109:@2005.4]
  assign buffer_0_708 = $signed(_T_55730); // @[Modules.scala 71:109:@2006.4]
  assign _T_55732 = $signed(buffer_0_634) + $signed(buffer_0_635); // @[Modules.scala 71:109:@2008.4]
  assign _T_55733 = _T_55732[10:0]; // @[Modules.scala 71:109:@2009.4]
  assign buffer_0_709 = $signed(_T_55733); // @[Modules.scala 71:109:@2010.4]
  assign _T_55735 = $signed(buffer_0_636) + $signed(buffer_0_637); // @[Modules.scala 71:109:@2012.4]
  assign _T_55736 = _T_55735[10:0]; // @[Modules.scala 71:109:@2013.4]
  assign buffer_0_710 = $signed(_T_55736); // @[Modules.scala 71:109:@2014.4]
  assign _T_55738 = $signed(buffer_0_638) + $signed(buffer_0_639); // @[Modules.scala 71:109:@2016.4]
  assign _T_55739 = _T_55738[10:0]; // @[Modules.scala 71:109:@2017.4]
  assign buffer_0_711 = $signed(_T_55739); // @[Modules.scala 71:109:@2018.4]
  assign _T_55741 = $signed(buffer_0_640) + $signed(buffer_0_641); // @[Modules.scala 71:109:@2020.4]
  assign _T_55742 = _T_55741[10:0]; // @[Modules.scala 71:109:@2021.4]
  assign buffer_0_712 = $signed(_T_55742); // @[Modules.scala 71:109:@2022.4]
  assign _T_55744 = $signed(buffer_0_642) + $signed(buffer_0_643); // @[Modules.scala 71:109:@2024.4]
  assign _T_55745 = _T_55744[10:0]; // @[Modules.scala 71:109:@2025.4]
  assign buffer_0_713 = $signed(_T_55745); // @[Modules.scala 71:109:@2026.4]
  assign _T_55747 = $signed(buffer_0_644) + $signed(buffer_0_645); // @[Modules.scala 71:109:@2028.4]
  assign _T_55748 = _T_55747[10:0]; // @[Modules.scala 71:109:@2029.4]
  assign buffer_0_714 = $signed(_T_55748); // @[Modules.scala 71:109:@2030.4]
  assign _T_55750 = $signed(buffer_0_646) + $signed(buffer_0_647); // @[Modules.scala 71:109:@2032.4]
  assign _T_55751 = _T_55750[10:0]; // @[Modules.scala 71:109:@2033.4]
  assign buffer_0_715 = $signed(_T_55751); // @[Modules.scala 71:109:@2034.4]
  assign _T_55753 = $signed(buffer_0_648) + $signed(buffer_0_649); // @[Modules.scala 71:109:@2036.4]
  assign _T_55754 = _T_55753[10:0]; // @[Modules.scala 71:109:@2037.4]
  assign buffer_0_716 = $signed(_T_55754); // @[Modules.scala 71:109:@2038.4]
  assign _T_55756 = $signed(buffer_0_650) + $signed(buffer_0_651); // @[Modules.scala 71:109:@2040.4]
  assign _T_55757 = _T_55756[10:0]; // @[Modules.scala 71:109:@2041.4]
  assign buffer_0_717 = $signed(_T_55757); // @[Modules.scala 71:109:@2042.4]
  assign _T_55759 = $signed(buffer_0_652) + $signed(buffer_0_653); // @[Modules.scala 71:109:@2044.4]
  assign _T_55760 = _T_55759[10:0]; // @[Modules.scala 71:109:@2045.4]
  assign buffer_0_718 = $signed(_T_55760); // @[Modules.scala 71:109:@2046.4]
  assign _T_55762 = $signed(buffer_0_654) + $signed(buffer_0_655); // @[Modules.scala 71:109:@2048.4]
  assign _T_55763 = _T_55762[10:0]; // @[Modules.scala 71:109:@2049.4]
  assign buffer_0_719 = $signed(_T_55763); // @[Modules.scala 71:109:@2050.4]
  assign _T_55765 = $signed(buffer_0_656) + $signed(buffer_0_657); // @[Modules.scala 71:109:@2052.4]
  assign _T_55766 = _T_55765[10:0]; // @[Modules.scala 71:109:@2053.4]
  assign buffer_0_720 = $signed(_T_55766); // @[Modules.scala 71:109:@2054.4]
  assign _T_55768 = $signed(buffer_0_593) + $signed(buffer_0_659); // @[Modules.scala 71:109:@2056.4]
  assign _T_55769 = _T_55768[10:0]; // @[Modules.scala 71:109:@2057.4]
  assign buffer_0_721 = $signed(_T_55769); // @[Modules.scala 71:109:@2058.4]
  assign _T_55771 = $signed(buffer_0_660) + $signed(buffer_0_661); // @[Modules.scala 71:109:@2060.4]
  assign _T_55772 = _T_55771[10:0]; // @[Modules.scala 71:109:@2061.4]
  assign buffer_0_722 = $signed(_T_55772); // @[Modules.scala 71:109:@2062.4]
  assign _T_55774 = $signed(buffer_0_593) + $signed(buffer_0_663); // @[Modules.scala 71:109:@2064.4]
  assign _T_55775 = _T_55774[10:0]; // @[Modules.scala 71:109:@2065.4]
  assign buffer_0_723 = $signed(_T_55775); // @[Modules.scala 71:109:@2066.4]
  assign _T_55777 = $signed(buffer_0_664) + $signed(buffer_0_665); // @[Modules.scala 71:109:@2068.4]
  assign _T_55778 = _T_55777[10:0]; // @[Modules.scala 71:109:@2069.4]
  assign buffer_0_724 = $signed(_T_55778); // @[Modules.scala 71:109:@2070.4]
  assign _T_55780 = $signed(buffer_0_593) + $signed(buffer_0_667); // @[Modules.scala 71:109:@2072.4]
  assign _T_55781 = _T_55780[10:0]; // @[Modules.scala 71:109:@2073.4]
  assign buffer_0_725 = $signed(_T_55781); // @[Modules.scala 71:109:@2074.4]
  assign _T_55783 = $signed(buffer_0_668) + $signed(buffer_0_593); // @[Modules.scala 71:109:@2076.4]
  assign _T_55784 = _T_55783[10:0]; // @[Modules.scala 71:109:@2077.4]
  assign buffer_0_726 = $signed(_T_55784); // @[Modules.scala 71:109:@2078.4]
  assign _T_55786 = $signed(buffer_0_670) + $signed(buffer_0_671); // @[Modules.scala 71:109:@2080.4]
  assign _T_55787 = _T_55786[10:0]; // @[Modules.scala 71:109:@2081.4]
  assign buffer_0_727 = $signed(_T_55787); // @[Modules.scala 71:109:@2082.4]
  assign _T_55789 = $signed(buffer_0_672) + $signed(buffer_0_673); // @[Modules.scala 71:109:@2084.4]
  assign _T_55790 = _T_55789[10:0]; // @[Modules.scala 71:109:@2085.4]
  assign buffer_0_728 = $signed(_T_55790); // @[Modules.scala 71:109:@2086.4]
  assign _T_55792 = $signed(buffer_0_674) + $signed(buffer_0_675); // @[Modules.scala 71:109:@2088.4]
  assign _T_55793 = _T_55792[10:0]; // @[Modules.scala 71:109:@2089.4]
  assign buffer_0_729 = $signed(_T_55793); // @[Modules.scala 71:109:@2090.4]
  assign _T_55795 = $signed(buffer_0_676) + $signed(buffer_0_677); // @[Modules.scala 71:109:@2092.4]
  assign _T_55796 = _T_55795[10:0]; // @[Modules.scala 71:109:@2093.4]
  assign buffer_0_730 = $signed(_T_55796); // @[Modules.scala 71:109:@2094.4]
  assign _T_55798 = $signed(buffer_0_678) + $signed(buffer_0_679); // @[Modules.scala 71:109:@2096.4]
  assign _T_55799 = _T_55798[10:0]; // @[Modules.scala 71:109:@2097.4]
  assign buffer_0_731 = $signed(_T_55799); // @[Modules.scala 71:109:@2098.4]
  assign _T_55801 = $signed(buffer_0_680) + $signed(buffer_0_681); // @[Modules.scala 71:109:@2100.4]
  assign _T_55802 = _T_55801[10:0]; // @[Modules.scala 71:109:@2101.4]
  assign buffer_0_732 = $signed(_T_55802); // @[Modules.scala 71:109:@2102.4]
  assign _T_55804 = $signed(buffer_0_682) + $signed(buffer_0_683); // @[Modules.scala 71:109:@2104.4]
  assign _T_55805 = _T_55804[10:0]; // @[Modules.scala 71:109:@2105.4]
  assign buffer_0_733 = $signed(_T_55805); // @[Modules.scala 71:109:@2106.4]
  assign _T_55807 = $signed(buffer_0_684) + $signed(buffer_0_685); // @[Modules.scala 71:109:@2108.4]
  assign _T_55808 = _T_55807[10:0]; // @[Modules.scala 71:109:@2109.4]
  assign buffer_0_734 = $signed(_T_55808); // @[Modules.scala 71:109:@2110.4]
  assign _T_55810 = $signed(buffer_0_686) + $signed(buffer_0_687); // @[Modules.scala 78:156:@2113.4]
  assign _T_55811 = _T_55810[10:0]; // @[Modules.scala 78:156:@2114.4]
  assign buffer_0_736 = $signed(_T_55811); // @[Modules.scala 78:156:@2115.4]
  assign _T_55813 = $signed(buffer_0_736) + $signed(buffer_0_688); // @[Modules.scala 78:156:@2117.4]
  assign _T_55814 = _T_55813[10:0]; // @[Modules.scala 78:156:@2118.4]
  assign buffer_0_737 = $signed(_T_55814); // @[Modules.scala 78:156:@2119.4]
  assign _T_55816 = $signed(buffer_0_737) + $signed(buffer_0_689); // @[Modules.scala 78:156:@2121.4]
  assign _T_55817 = _T_55816[10:0]; // @[Modules.scala 78:156:@2122.4]
  assign buffer_0_738 = $signed(_T_55817); // @[Modules.scala 78:156:@2123.4]
  assign _T_55819 = $signed(buffer_0_738) + $signed(buffer_0_690); // @[Modules.scala 78:156:@2125.4]
  assign _T_55820 = _T_55819[10:0]; // @[Modules.scala 78:156:@2126.4]
  assign buffer_0_739 = $signed(_T_55820); // @[Modules.scala 78:156:@2127.4]
  assign _T_55822 = $signed(buffer_0_739) + $signed(buffer_0_691); // @[Modules.scala 78:156:@2129.4]
  assign _T_55823 = _T_55822[10:0]; // @[Modules.scala 78:156:@2130.4]
  assign buffer_0_740 = $signed(_T_55823); // @[Modules.scala 78:156:@2131.4]
  assign _T_55825 = $signed(buffer_0_740) + $signed(buffer_0_692); // @[Modules.scala 78:156:@2133.4]
  assign _T_55826 = _T_55825[10:0]; // @[Modules.scala 78:156:@2134.4]
  assign buffer_0_741 = $signed(_T_55826); // @[Modules.scala 78:156:@2135.4]
  assign _T_55828 = $signed(buffer_0_741) + $signed(buffer_0_693); // @[Modules.scala 78:156:@2137.4]
  assign _T_55829 = _T_55828[10:0]; // @[Modules.scala 78:156:@2138.4]
  assign buffer_0_742 = $signed(_T_55829); // @[Modules.scala 78:156:@2139.4]
  assign _T_55831 = $signed(buffer_0_742) + $signed(buffer_0_694); // @[Modules.scala 78:156:@2141.4]
  assign _T_55832 = _T_55831[10:0]; // @[Modules.scala 78:156:@2142.4]
  assign buffer_0_743 = $signed(_T_55832); // @[Modules.scala 78:156:@2143.4]
  assign _T_55834 = $signed(buffer_0_743) + $signed(buffer_0_695); // @[Modules.scala 78:156:@2145.4]
  assign _T_55835 = _T_55834[10:0]; // @[Modules.scala 78:156:@2146.4]
  assign buffer_0_744 = $signed(_T_55835); // @[Modules.scala 78:156:@2147.4]
  assign _T_55837 = $signed(buffer_0_744) + $signed(buffer_0_696); // @[Modules.scala 78:156:@2149.4]
  assign _T_55838 = _T_55837[10:0]; // @[Modules.scala 78:156:@2150.4]
  assign buffer_0_745 = $signed(_T_55838); // @[Modules.scala 78:156:@2151.4]
  assign _T_55840 = $signed(buffer_0_745) + $signed(buffer_0_697); // @[Modules.scala 78:156:@2153.4]
  assign _T_55841 = _T_55840[10:0]; // @[Modules.scala 78:156:@2154.4]
  assign buffer_0_746 = $signed(_T_55841); // @[Modules.scala 78:156:@2155.4]
  assign _T_55843 = $signed(buffer_0_746) + $signed(buffer_0_698); // @[Modules.scala 78:156:@2157.4]
  assign _T_55844 = _T_55843[10:0]; // @[Modules.scala 78:156:@2158.4]
  assign buffer_0_747 = $signed(_T_55844); // @[Modules.scala 78:156:@2159.4]
  assign _T_55846 = $signed(buffer_0_747) + $signed(buffer_0_699); // @[Modules.scala 78:156:@2161.4]
  assign _T_55847 = _T_55846[10:0]; // @[Modules.scala 78:156:@2162.4]
  assign buffer_0_748 = $signed(_T_55847); // @[Modules.scala 78:156:@2163.4]
  assign _T_55849 = $signed(buffer_0_748) + $signed(buffer_0_700); // @[Modules.scala 78:156:@2165.4]
  assign _T_55850 = _T_55849[10:0]; // @[Modules.scala 78:156:@2166.4]
  assign buffer_0_749 = $signed(_T_55850); // @[Modules.scala 78:156:@2167.4]
  assign _T_55852 = $signed(buffer_0_749) + $signed(buffer_0_701); // @[Modules.scala 78:156:@2169.4]
  assign _T_55853 = _T_55852[10:0]; // @[Modules.scala 78:156:@2170.4]
  assign buffer_0_750 = $signed(_T_55853); // @[Modules.scala 78:156:@2171.4]
  assign _T_55855 = $signed(buffer_0_750) + $signed(buffer_0_702); // @[Modules.scala 78:156:@2173.4]
  assign _T_55856 = _T_55855[10:0]; // @[Modules.scala 78:156:@2174.4]
  assign buffer_0_751 = $signed(_T_55856); // @[Modules.scala 78:156:@2175.4]
  assign _T_55858 = $signed(buffer_0_751) + $signed(buffer_0_701); // @[Modules.scala 78:156:@2177.4]
  assign _T_55859 = _T_55858[10:0]; // @[Modules.scala 78:156:@2178.4]
  assign buffer_0_752 = $signed(_T_55859); // @[Modules.scala 78:156:@2179.4]
  assign _T_55861 = $signed(buffer_0_752) + $signed(buffer_0_704); // @[Modules.scala 78:156:@2181.4]
  assign _T_55862 = _T_55861[10:0]; // @[Modules.scala 78:156:@2182.4]
  assign buffer_0_753 = $signed(_T_55862); // @[Modules.scala 78:156:@2183.4]
  assign _T_55864 = $signed(buffer_0_753) + $signed(buffer_0_705); // @[Modules.scala 78:156:@2185.4]
  assign _T_55865 = _T_55864[10:0]; // @[Modules.scala 78:156:@2186.4]
  assign buffer_0_754 = $signed(_T_55865); // @[Modules.scala 78:156:@2187.4]
  assign _T_55867 = $signed(buffer_0_754) + $signed(buffer_0_706); // @[Modules.scala 78:156:@2189.4]
  assign _T_55868 = _T_55867[10:0]; // @[Modules.scala 78:156:@2190.4]
  assign buffer_0_755 = $signed(_T_55868); // @[Modules.scala 78:156:@2191.4]
  assign _T_55870 = $signed(buffer_0_755) + $signed(buffer_0_707); // @[Modules.scala 78:156:@2193.4]
  assign _T_55871 = _T_55870[10:0]; // @[Modules.scala 78:156:@2194.4]
  assign buffer_0_756 = $signed(_T_55871); // @[Modules.scala 78:156:@2195.4]
  assign _T_55873 = $signed(buffer_0_756) + $signed(buffer_0_708); // @[Modules.scala 78:156:@2197.4]
  assign _T_55874 = _T_55873[10:0]; // @[Modules.scala 78:156:@2198.4]
  assign buffer_0_757 = $signed(_T_55874); // @[Modules.scala 78:156:@2199.4]
  assign _T_55876 = $signed(buffer_0_757) + $signed(buffer_0_709); // @[Modules.scala 78:156:@2201.4]
  assign _T_55877 = _T_55876[10:0]; // @[Modules.scala 78:156:@2202.4]
  assign buffer_0_758 = $signed(_T_55877); // @[Modules.scala 78:156:@2203.4]
  assign _T_55879 = $signed(buffer_0_758) + $signed(buffer_0_710); // @[Modules.scala 78:156:@2205.4]
  assign _T_55880 = _T_55879[10:0]; // @[Modules.scala 78:156:@2206.4]
  assign buffer_0_759 = $signed(_T_55880); // @[Modules.scala 78:156:@2207.4]
  assign _T_55882 = $signed(buffer_0_759) + $signed(buffer_0_711); // @[Modules.scala 78:156:@2209.4]
  assign _T_55883 = _T_55882[10:0]; // @[Modules.scala 78:156:@2210.4]
  assign buffer_0_760 = $signed(_T_55883); // @[Modules.scala 78:156:@2211.4]
  assign _T_55885 = $signed(buffer_0_760) + $signed(buffer_0_712); // @[Modules.scala 78:156:@2213.4]
  assign _T_55886 = _T_55885[10:0]; // @[Modules.scala 78:156:@2214.4]
  assign buffer_0_761 = $signed(_T_55886); // @[Modules.scala 78:156:@2215.4]
  assign _T_55888 = $signed(buffer_0_761) + $signed(buffer_0_713); // @[Modules.scala 78:156:@2217.4]
  assign _T_55889 = _T_55888[10:0]; // @[Modules.scala 78:156:@2218.4]
  assign buffer_0_762 = $signed(_T_55889); // @[Modules.scala 78:156:@2219.4]
  assign _T_55891 = $signed(buffer_0_762) + $signed(buffer_0_714); // @[Modules.scala 78:156:@2221.4]
  assign _T_55892 = _T_55891[10:0]; // @[Modules.scala 78:156:@2222.4]
  assign buffer_0_763 = $signed(_T_55892); // @[Modules.scala 78:156:@2223.4]
  assign _T_55894 = $signed(buffer_0_763) + $signed(buffer_0_715); // @[Modules.scala 78:156:@2225.4]
  assign _T_55895 = _T_55894[10:0]; // @[Modules.scala 78:156:@2226.4]
  assign buffer_0_764 = $signed(_T_55895); // @[Modules.scala 78:156:@2227.4]
  assign _T_55897 = $signed(buffer_0_764) + $signed(buffer_0_716); // @[Modules.scala 78:156:@2229.4]
  assign _T_55898 = _T_55897[10:0]; // @[Modules.scala 78:156:@2230.4]
  assign buffer_0_765 = $signed(_T_55898); // @[Modules.scala 78:156:@2231.4]
  assign _T_55900 = $signed(buffer_0_765) + $signed(buffer_0_717); // @[Modules.scala 78:156:@2233.4]
  assign _T_55901 = _T_55900[10:0]; // @[Modules.scala 78:156:@2234.4]
  assign buffer_0_766 = $signed(_T_55901); // @[Modules.scala 78:156:@2235.4]
  assign _T_55903 = $signed(buffer_0_766) + $signed(buffer_0_718); // @[Modules.scala 78:156:@2237.4]
  assign _T_55904 = _T_55903[10:0]; // @[Modules.scala 78:156:@2238.4]
  assign buffer_0_767 = $signed(_T_55904); // @[Modules.scala 78:156:@2239.4]
  assign _T_55906 = $signed(buffer_0_767) + $signed(buffer_0_719); // @[Modules.scala 78:156:@2241.4]
  assign _T_55907 = _T_55906[10:0]; // @[Modules.scala 78:156:@2242.4]
  assign buffer_0_768 = $signed(_T_55907); // @[Modules.scala 78:156:@2243.4]
  assign _T_55909 = $signed(buffer_0_768) + $signed(buffer_0_720); // @[Modules.scala 78:156:@2245.4]
  assign _T_55910 = _T_55909[10:0]; // @[Modules.scala 78:156:@2246.4]
  assign buffer_0_769 = $signed(_T_55910); // @[Modules.scala 78:156:@2247.4]
  assign _T_55912 = $signed(buffer_0_769) + $signed(buffer_0_721); // @[Modules.scala 78:156:@2249.4]
  assign _T_55913 = _T_55912[10:0]; // @[Modules.scala 78:156:@2250.4]
  assign buffer_0_770 = $signed(_T_55913); // @[Modules.scala 78:156:@2251.4]
  assign _T_55915 = $signed(buffer_0_770) + $signed(buffer_0_722); // @[Modules.scala 78:156:@2253.4]
  assign _T_55916 = _T_55915[10:0]; // @[Modules.scala 78:156:@2254.4]
  assign buffer_0_771 = $signed(_T_55916); // @[Modules.scala 78:156:@2255.4]
  assign _T_55918 = $signed(buffer_0_771) + $signed(buffer_0_723); // @[Modules.scala 78:156:@2257.4]
  assign _T_55919 = _T_55918[10:0]; // @[Modules.scala 78:156:@2258.4]
  assign buffer_0_772 = $signed(_T_55919); // @[Modules.scala 78:156:@2259.4]
  assign _T_55921 = $signed(buffer_0_772) + $signed(buffer_0_724); // @[Modules.scala 78:156:@2261.4]
  assign _T_55922 = _T_55921[10:0]; // @[Modules.scala 78:156:@2262.4]
  assign buffer_0_773 = $signed(_T_55922); // @[Modules.scala 78:156:@2263.4]
  assign _T_55924 = $signed(buffer_0_773) + $signed(buffer_0_725); // @[Modules.scala 78:156:@2265.4]
  assign _T_55925 = _T_55924[10:0]; // @[Modules.scala 78:156:@2266.4]
  assign buffer_0_774 = $signed(_T_55925); // @[Modules.scala 78:156:@2267.4]
  assign _T_55927 = $signed(buffer_0_774) + $signed(buffer_0_726); // @[Modules.scala 78:156:@2269.4]
  assign _T_55928 = _T_55927[10:0]; // @[Modules.scala 78:156:@2270.4]
  assign buffer_0_775 = $signed(_T_55928); // @[Modules.scala 78:156:@2271.4]
  assign _T_55930 = $signed(buffer_0_775) + $signed(buffer_0_727); // @[Modules.scala 78:156:@2273.4]
  assign _T_55931 = _T_55930[10:0]; // @[Modules.scala 78:156:@2274.4]
  assign buffer_0_776 = $signed(_T_55931); // @[Modules.scala 78:156:@2275.4]
  assign _T_55933 = $signed(buffer_0_776) + $signed(buffer_0_728); // @[Modules.scala 78:156:@2277.4]
  assign _T_55934 = _T_55933[10:0]; // @[Modules.scala 78:156:@2278.4]
  assign buffer_0_777 = $signed(_T_55934); // @[Modules.scala 78:156:@2279.4]
  assign _T_55936 = $signed(buffer_0_777) + $signed(buffer_0_729); // @[Modules.scala 78:156:@2281.4]
  assign _T_55937 = _T_55936[10:0]; // @[Modules.scala 78:156:@2282.4]
  assign buffer_0_778 = $signed(_T_55937); // @[Modules.scala 78:156:@2283.4]
  assign _T_55939 = $signed(buffer_0_778) + $signed(buffer_0_730); // @[Modules.scala 78:156:@2285.4]
  assign _T_55940 = _T_55939[10:0]; // @[Modules.scala 78:156:@2286.4]
  assign buffer_0_779 = $signed(_T_55940); // @[Modules.scala 78:156:@2287.4]
  assign _T_55942 = $signed(buffer_0_779) + $signed(buffer_0_731); // @[Modules.scala 78:156:@2289.4]
  assign _T_55943 = _T_55942[10:0]; // @[Modules.scala 78:156:@2290.4]
  assign buffer_0_780 = $signed(_T_55943); // @[Modules.scala 78:156:@2291.4]
  assign _T_55945 = $signed(buffer_0_780) + $signed(buffer_0_732); // @[Modules.scala 78:156:@2293.4]
  assign _T_55946 = _T_55945[10:0]; // @[Modules.scala 78:156:@2294.4]
  assign buffer_0_781 = $signed(_T_55946); // @[Modules.scala 78:156:@2295.4]
  assign _T_55948 = $signed(buffer_0_781) + $signed(buffer_0_733); // @[Modules.scala 78:156:@2297.4]
  assign _T_55949 = _T_55948[10:0]; // @[Modules.scala 78:156:@2298.4]
  assign buffer_0_782 = $signed(_T_55949); // @[Modules.scala 78:156:@2299.4]
  assign _T_55951 = $signed(buffer_0_782) + $signed(buffer_0_734); // @[Modules.scala 78:156:@2301.4]
  assign _T_55952 = _T_55951[10:0]; // @[Modules.scala 78:156:@2302.4]
  assign buffer_0_783 = $signed(_T_55952); // @[Modules.scala 78:156:@2303.4]
  assign _T_55956 = $signed(io_in_4) + $signed(io_in_5); // @[Modules.scala 37:46:@2308.4]
  assign _T_55957 = _T_55956[4:0]; // @[Modules.scala 37:46:@2309.4]
  assign _T_55958 = $signed(_T_55957); // @[Modules.scala 37:46:@2310.4]
  assign _T_55959 = $signed(io_in_6) + $signed(io_in_7); // @[Modules.scala 37:46:@2312.4]
  assign _T_55960 = _T_55959[4:0]; // @[Modules.scala 37:46:@2313.4]
  assign _T_55961 = $signed(_T_55960); // @[Modules.scala 37:46:@2314.4]
  assign _T_55962 = $signed(io_in_8) + $signed(io_in_9); // @[Modules.scala 37:46:@2316.4]
  assign _T_55963 = _T_55962[4:0]; // @[Modules.scala 37:46:@2317.4]
  assign _T_55964 = $signed(_T_55963); // @[Modules.scala 37:46:@2318.4]
  assign _T_55966 = $signed(io_in_12) + $signed(io_in_13); // @[Modules.scala 37:46:@2321.4]
  assign _T_55967 = _T_55966[4:0]; // @[Modules.scala 37:46:@2322.4]
  assign _T_55968 = $signed(_T_55967); // @[Modules.scala 37:46:@2323.4]
  assign _T_55969 = $signed(io_in_14) + $signed(io_in_15); // @[Modules.scala 37:46:@2325.4]
  assign _T_55970 = _T_55969[4:0]; // @[Modules.scala 37:46:@2326.4]
  assign _T_55971 = $signed(_T_55970); // @[Modules.scala 37:46:@2327.4]
  assign _T_55975 = $signed(io_in_24) + $signed(io_in_25); // @[Modules.scala 37:46:@2336.4]
  assign _T_55976 = _T_55975[4:0]; // @[Modules.scala 37:46:@2337.4]
  assign _T_55977 = $signed(_T_55976); // @[Modules.scala 37:46:@2338.4]
  assign _T_55979 = $signed(io_in_30) + $signed(io_in_31); // @[Modules.scala 37:46:@2342.4]
  assign _T_55980 = _T_55979[4:0]; // @[Modules.scala 37:46:@2343.4]
  assign _T_55981 = $signed(_T_55980); // @[Modules.scala 37:46:@2344.4]
  assign _T_55985 = $signed(io_in_34) + $signed(io_in_35); // @[Modules.scala 37:46:@2350.4]
  assign _T_55986 = _T_55985[4:0]; // @[Modules.scala 37:46:@2351.4]
  assign _T_55987 = $signed(_T_55986); // @[Modules.scala 37:46:@2352.4]
  assign _T_55988 = $signed(io_in_36) + $signed(io_in_37); // @[Modules.scala 37:46:@2354.4]
  assign _T_55989 = _T_55988[4:0]; // @[Modules.scala 37:46:@2355.4]
  assign _T_55990 = $signed(_T_55989); // @[Modules.scala 37:46:@2356.4]
  assign _T_55991 = $signed(io_in_38) + $signed(io_in_39); // @[Modules.scala 37:46:@2358.4]
  assign _T_55992 = _T_55991[4:0]; // @[Modules.scala 37:46:@2359.4]
  assign _T_55993 = $signed(_T_55992); // @[Modules.scala 37:46:@2360.4]
  assign _T_55994 = $signed(io_in_40) + $signed(io_in_41); // @[Modules.scala 37:46:@2362.4]
  assign _T_55995 = _T_55994[4:0]; // @[Modules.scala 37:46:@2363.4]
  assign _T_55996 = $signed(_T_55995); // @[Modules.scala 37:46:@2364.4]
  assign _T_55997 = $signed(io_in_42) + $signed(io_in_43); // @[Modules.scala 37:46:@2366.4]
  assign _T_55998 = _T_55997[4:0]; // @[Modules.scala 37:46:@2367.4]
  assign _T_55999 = $signed(_T_55998); // @[Modules.scala 37:46:@2368.4]
  assign _T_56000 = $signed(io_in_46) + $signed(io_in_47); // @[Modules.scala 37:46:@2371.4]
  assign _T_56001 = _T_56000[4:0]; // @[Modules.scala 37:46:@2372.4]
  assign _T_56002 = $signed(_T_56001); // @[Modules.scala 37:46:@2373.4]
  assign _T_56003 = $signed(io_in_48) + $signed(io_in_49); // @[Modules.scala 37:46:@2375.4]
  assign _T_56004 = _T_56003[4:0]; // @[Modules.scala 37:46:@2376.4]
  assign _T_56005 = $signed(_T_56004); // @[Modules.scala 37:46:@2377.4]
  assign _T_56006 = $signed(io_in_50) + $signed(io_in_51); // @[Modules.scala 37:46:@2379.4]
  assign _T_56007 = _T_56006[4:0]; // @[Modules.scala 37:46:@2380.4]
  assign _T_56008 = $signed(_T_56007); // @[Modules.scala 37:46:@2381.4]
  assign _T_56009 = $signed(io_in_58) + $signed(io_in_59); // @[Modules.scala 37:46:@2386.4]
  assign _T_56010 = _T_56009[4:0]; // @[Modules.scala 37:46:@2387.4]
  assign _T_56011 = $signed(_T_56010); // @[Modules.scala 37:46:@2388.4]
  assign _T_56012 = $signed(io_in_60) + $signed(io_in_61); // @[Modules.scala 37:46:@2390.4]
  assign _T_56013 = _T_56012[4:0]; // @[Modules.scala 37:46:@2391.4]
  assign _T_56014 = $signed(_T_56013); // @[Modules.scala 37:46:@2392.4]
  assign _T_56015 = $signed(io_in_62) + $signed(io_in_63); // @[Modules.scala 37:46:@2394.4]
  assign _T_56016 = _T_56015[4:0]; // @[Modules.scala 37:46:@2395.4]
  assign _T_56017 = $signed(_T_56016); // @[Modules.scala 37:46:@2396.4]
  assign _T_56018 = $signed(io_in_64) + $signed(io_in_65); // @[Modules.scala 37:46:@2398.4]
  assign _T_56019 = _T_56018[4:0]; // @[Modules.scala 37:46:@2399.4]
  assign _T_56020 = $signed(_T_56019); // @[Modules.scala 37:46:@2400.4]
  assign _T_56021 = $signed(io_in_66) + $signed(io_in_67); // @[Modules.scala 37:46:@2402.4]
  assign _T_56022 = _T_56021[4:0]; // @[Modules.scala 37:46:@2403.4]
  assign _T_56023 = $signed(_T_56022); // @[Modules.scala 37:46:@2404.4]
  assign _T_56024 = $signed(io_in_68) + $signed(io_in_69); // @[Modules.scala 37:46:@2406.4]
  assign _T_56025 = _T_56024[4:0]; // @[Modules.scala 37:46:@2407.4]
  assign _T_56026 = $signed(_T_56025); // @[Modules.scala 37:46:@2408.4]
  assign _T_56027 = $signed(io_in_70) + $signed(io_in_71); // @[Modules.scala 37:46:@2410.4]
  assign _T_56028 = _T_56027[4:0]; // @[Modules.scala 37:46:@2411.4]
  assign _T_56029 = $signed(_T_56028); // @[Modules.scala 37:46:@2412.4]
  assign _T_56030 = $signed(io_in_72) + $signed(io_in_73); // @[Modules.scala 37:46:@2414.4]
  assign _T_56031 = _T_56030[4:0]; // @[Modules.scala 37:46:@2415.4]
  assign _T_56032 = $signed(_T_56031); // @[Modules.scala 37:46:@2416.4]
  assign _T_56033 = $signed(io_in_74) + $signed(io_in_75); // @[Modules.scala 37:46:@2418.4]
  assign _T_56034 = _T_56033[4:0]; // @[Modules.scala 37:46:@2419.4]
  assign _T_56035 = $signed(_T_56034); // @[Modules.scala 37:46:@2420.4]
  assign _T_56036 = $signed(io_in_76) + $signed(io_in_77); // @[Modules.scala 37:46:@2422.4]
  assign _T_56037 = _T_56036[4:0]; // @[Modules.scala 37:46:@2423.4]
  assign _T_56038 = $signed(_T_56037); // @[Modules.scala 37:46:@2424.4]
  assign _T_56042 = $signed(io_in_80) + $signed(io_in_81); // @[Modules.scala 37:46:@2430.4]
  assign _T_56043 = _T_56042[4:0]; // @[Modules.scala 37:46:@2431.4]
  assign _T_56044 = $signed(_T_56043); // @[Modules.scala 37:46:@2432.4]
  assign _T_56052 = $signed(io_in_92) + $signed(io_in_93); // @[Modules.scala 37:46:@2445.4]
  assign _T_56053 = _T_56052[4:0]; // @[Modules.scala 37:46:@2446.4]
  assign _T_56054 = $signed(_T_56053); // @[Modules.scala 37:46:@2447.4]
  assign _T_56058 = $signed(io_in_96) + $signed(io_in_97); // @[Modules.scala 37:46:@2453.4]
  assign _T_56059 = _T_56058[4:0]; // @[Modules.scala 37:46:@2454.4]
  assign _T_56060 = $signed(_T_56059); // @[Modules.scala 37:46:@2455.4]
  assign _T_56076 = $signed(io_in_108) + $signed(io_in_109); // @[Modules.scala 37:46:@2477.4]
  assign _T_56077 = _T_56076[4:0]; // @[Modules.scala 37:46:@2478.4]
  assign _T_56078 = $signed(_T_56077); // @[Modules.scala 37:46:@2479.4]
  assign _T_56087 = $signed(io_in_128) + $signed(io_in_129); // @[Modules.scala 37:46:@2493.4]
  assign _T_56088 = _T_56087[4:0]; // @[Modules.scala 37:46:@2494.4]
  assign _T_56089 = $signed(_T_56088); // @[Modules.scala 37:46:@2495.4]
  assign _T_56090 = $signed(io_in_130) + $signed(io_in_131); // @[Modules.scala 37:46:@2497.4]
  assign _T_56091 = _T_56090[4:0]; // @[Modules.scala 37:46:@2498.4]
  assign _T_56092 = $signed(_T_56091); // @[Modules.scala 37:46:@2499.4]
  assign _T_56096 = $signed(io_in_136) + $signed(io_in_137); // @[Modules.scala 37:46:@2506.4]
  assign _T_56097 = _T_56096[4:0]; // @[Modules.scala 37:46:@2507.4]
  assign _T_56098 = $signed(_T_56097); // @[Modules.scala 37:46:@2508.4]
  assign _T_56106 = $signed(io_in_166) + $signed(io_in_167); // @[Modules.scala 37:46:@2524.4]
  assign _T_56107 = _T_56106[4:0]; // @[Modules.scala 37:46:@2525.4]
  assign _T_56108 = $signed(_T_56107); // @[Modules.scala 37:46:@2526.4]
  assign _T_56109 = $signed(io_in_170) + $signed(io_in_171); // @[Modules.scala 37:46:@2529.4]
  assign _T_56110 = _T_56109[4:0]; // @[Modules.scala 37:46:@2530.4]
  assign _T_56111 = $signed(_T_56110); // @[Modules.scala 37:46:@2531.4]
  assign _T_56112 = $signed(io_in_174) + $signed(io_in_175); // @[Modules.scala 37:46:@2534.4]
  assign _T_56113 = _T_56112[4:0]; // @[Modules.scala 37:46:@2535.4]
  assign _T_56114 = $signed(_T_56113); // @[Modules.scala 37:46:@2536.4]
  assign _T_56115 = $signed(io_in_176) + $signed(io_in_177); // @[Modules.scala 37:46:@2538.4]
  assign _T_56116 = _T_56115[4:0]; // @[Modules.scala 37:46:@2539.4]
  assign _T_56117 = $signed(_T_56116); // @[Modules.scala 37:46:@2540.4]
  assign _T_56123 = $signed(io_in_196) + $signed(io_in_197); // @[Modules.scala 37:46:@2554.4]
  assign _T_56124 = _T_56123[4:0]; // @[Modules.scala 37:46:@2555.4]
  assign _T_56125 = $signed(_T_56124); // @[Modules.scala 37:46:@2556.4]
  assign _T_56126 = $signed(io_in_202) + $signed(io_in_203); // @[Modules.scala 37:46:@2560.4]
  assign _T_56127 = _T_56126[4:0]; // @[Modules.scala 37:46:@2561.4]
  assign _T_56128 = $signed(_T_56127); // @[Modules.scala 37:46:@2562.4]
  assign _T_56132 = $signed(io_in_220) + $signed(io_in_221); // @[Modules.scala 37:46:@2575.4]
  assign _T_56133 = _T_56132[4:0]; // @[Modules.scala 37:46:@2576.4]
  assign _T_56134 = $signed(_T_56133); // @[Modules.scala 37:46:@2577.4]
  assign _T_56135 = $signed(io_in_224) + $signed(io_in_225); // @[Modules.scala 37:46:@2580.4]
  assign _T_56136 = _T_56135[4:0]; // @[Modules.scala 37:46:@2581.4]
  assign _T_56137 = $signed(_T_56136); // @[Modules.scala 37:46:@2582.4]
  assign _T_56145 = $signed(io_in_240) + $signed(io_in_241); // @[Modules.scala 37:46:@2591.4]
  assign _T_56146 = _T_56145[4:0]; // @[Modules.scala 37:46:@2592.4]
  assign _T_56147 = $signed(_T_56146); // @[Modules.scala 37:46:@2593.4]
  assign _T_56150 = $signed(io_in_248) + $signed(io_in_249); // @[Modules.scala 37:46:@2598.4]
  assign _T_56151 = _T_56150[4:0]; // @[Modules.scala 37:46:@2599.4]
  assign _T_56152 = $signed(_T_56151); // @[Modules.scala 37:46:@2600.4]
  assign _T_56153 = $signed(io_in_250) + $signed(io_in_251); // @[Modules.scala 37:46:@2602.4]
  assign _T_56154 = _T_56153[4:0]; // @[Modules.scala 37:46:@2603.4]
  assign _T_56155 = $signed(_T_56154); // @[Modules.scala 37:46:@2604.4]
  assign _T_56161 = $signed(io_in_266) + $signed(io_in_267); // @[Modules.scala 37:46:@2613.4]
  assign _T_56162 = _T_56161[4:0]; // @[Modules.scala 37:46:@2614.4]
  assign _T_56163 = $signed(_T_56162); // @[Modules.scala 37:46:@2615.4]
  assign _T_56167 = $signed(io_in_276) + $signed(io_in_277); // @[Modules.scala 37:46:@2621.4]
  assign _T_56168 = _T_56167[4:0]; // @[Modules.scala 37:46:@2622.4]
  assign _T_56169 = $signed(_T_56168); // @[Modules.scala 37:46:@2623.4]
  assign _T_56170 = $signed(io_in_278) + $signed(io_in_279); // @[Modules.scala 37:46:@2625.4]
  assign _T_56171 = _T_56170[4:0]; // @[Modules.scala 37:46:@2626.4]
  assign _T_56172 = $signed(_T_56171); // @[Modules.scala 37:46:@2627.4]
  assign _T_56176 = $signed(io_in_292) + $signed(io_in_293); // @[Modules.scala 37:46:@2635.4]
  assign _T_56177 = _T_56176[4:0]; // @[Modules.scala 37:46:@2636.4]
  assign _T_56178 = $signed(_T_56177); // @[Modules.scala 37:46:@2637.4]
  assign _T_56182 = $signed(io_in_304) + $signed(io_in_305); // @[Modules.scala 37:46:@2644.4]
  assign _T_56183 = _T_56182[4:0]; // @[Modules.scala 37:46:@2645.4]
  assign _T_56184 = $signed(_T_56183); // @[Modules.scala 37:46:@2646.4]
  assign _T_56185 = $signed(io_in_306) + $signed(io_in_307); // @[Modules.scala 37:46:@2648.4]
  assign _T_56186 = _T_56185[4:0]; // @[Modules.scala 37:46:@2649.4]
  assign _T_56187 = $signed(_T_56186); // @[Modules.scala 37:46:@2650.4]
  assign _T_56195 = $signed(io_in_320) + $signed(io_in_321); // @[Modules.scala 37:46:@2661.4]
  assign _T_56196 = _T_56195[4:0]; // @[Modules.scala 37:46:@2662.4]
  assign _T_56197 = $signed(_T_56196); // @[Modules.scala 37:46:@2663.4]
  assign _T_56201 = $signed(io_in_332) + $signed(io_in_333); // @[Modules.scala 37:46:@2670.4]
  assign _T_56202 = _T_56201[4:0]; // @[Modules.scala 37:46:@2671.4]
  assign _T_56203 = $signed(_T_56202); // @[Modules.scala 37:46:@2672.4]
  assign _T_56204 = $signed(io_in_334) + $signed(io_in_335); // @[Modules.scala 37:46:@2674.4]
  assign _T_56205 = _T_56204[4:0]; // @[Modules.scala 37:46:@2675.4]
  assign _T_56206 = $signed(_T_56205); // @[Modules.scala 37:46:@2676.4]
  assign _T_56224 = $signed(io_in_360) + $signed(io_in_361); // @[Modules.scala 37:46:@2702.4]
  assign _T_56225 = _T_56224[4:0]; // @[Modules.scala 37:46:@2703.4]
  assign _T_56226 = $signed(_T_56225); // @[Modules.scala 37:46:@2704.4]
  assign _T_56249 = $signed(io_in_392) + $signed(io_in_393); // @[Modules.scala 37:46:@2736.4]
  assign _T_56250 = _T_56249[4:0]; // @[Modules.scala 37:46:@2737.4]
  assign _T_56251 = $signed(_T_56250); // @[Modules.scala 37:46:@2738.4]
  assign _T_56281 = $signed(io_in_440) + $signed(io_in_441); // @[Modules.scala 37:46:@2784.4]
  assign _T_56282 = _T_56281[4:0]; // @[Modules.scala 37:46:@2785.4]
  assign _T_56283 = $signed(_T_56282); // @[Modules.scala 37:46:@2786.4]
  assign _T_56284 = $signed(io_in_442) + $signed(io_in_443); // @[Modules.scala 37:46:@2788.4]
  assign _T_56285 = _T_56284[4:0]; // @[Modules.scala 37:46:@2789.4]
  assign _T_56286 = $signed(_T_56285); // @[Modules.scala 37:46:@2790.4]
  assign _T_56288 = $signed(io_in_450) + $signed(io_in_451); // @[Modules.scala 37:46:@2795.4]
  assign _T_56289 = _T_56288[4:0]; // @[Modules.scala 37:46:@2796.4]
  assign _T_56290 = $signed(_T_56289); // @[Modules.scala 37:46:@2797.4]
  assign _T_56296 = $signed(io_in_468) + $signed(io_in_469); // @[Modules.scala 37:46:@2807.4]
  assign _T_56297 = _T_56296[4:0]; // @[Modules.scala 37:46:@2808.4]
  assign _T_56298 = $signed(_T_56297); // @[Modules.scala 37:46:@2809.4]
  assign _T_56299 = $signed(io_in_470) + $signed(io_in_471); // @[Modules.scala 37:46:@2811.4]
  assign _T_56300 = _T_56299[4:0]; // @[Modules.scala 37:46:@2812.4]
  assign _T_56301 = $signed(_T_56300); // @[Modules.scala 37:46:@2813.4]
  assign _T_56303 = $signed(io_in_478) + $signed(io_in_479); // @[Modules.scala 37:46:@2818.4]
  assign _T_56304 = _T_56303[4:0]; // @[Modules.scala 37:46:@2819.4]
  assign _T_56305 = $signed(_T_56304); // @[Modules.scala 37:46:@2820.4]
  assign _T_56315 = $signed(io_in_494) + $signed(io_in_495); // @[Modules.scala 37:46:@2832.4]
  assign _T_56316 = _T_56315[4:0]; // @[Modules.scala 37:46:@2833.4]
  assign _T_56317 = $signed(_T_56316); // @[Modules.scala 37:46:@2834.4]
  assign _T_56318 = $signed(io_in_496) + $signed(io_in_497); // @[Modules.scala 37:46:@2836.4]
  assign _T_56319 = _T_56318[4:0]; // @[Modules.scala 37:46:@2837.4]
  assign _T_56320 = $signed(_T_56319); // @[Modules.scala 37:46:@2838.4]
  assign _T_56326 = $signed(io_in_506) + $signed(io_in_507); // @[Modules.scala 37:46:@2847.4]
  assign _T_56327 = _T_56326[4:0]; // @[Modules.scala 37:46:@2848.4]
  assign _T_56328 = $signed(_T_56327); // @[Modules.scala 37:46:@2849.4]
  assign _T_56329 = $signed(io_in_510) + $signed(io_in_511); // @[Modules.scala 37:46:@2852.4]
  assign _T_56330 = _T_56329[4:0]; // @[Modules.scala 37:46:@2853.4]
  assign _T_56331 = $signed(_T_56330); // @[Modules.scala 37:46:@2854.4]
  assign _T_56338 = $signed(io_in_520) + $signed(io_in_521); // @[Modules.scala 37:46:@2863.4]
  assign _T_56339 = _T_56338[4:0]; // @[Modules.scala 37:46:@2864.4]
  assign _T_56340 = $signed(_T_56339); // @[Modules.scala 37:46:@2865.4]
  assign _T_56341 = $signed(io_in_522) + $signed(io_in_523); // @[Modules.scala 37:46:@2867.4]
  assign _T_56342 = _T_56341[4:0]; // @[Modules.scala 37:46:@2868.4]
  assign _T_56343 = $signed(_T_56342); // @[Modules.scala 37:46:@2869.4]
  assign _T_56344 = $signed(io_in_524) + $signed(io_in_525); // @[Modules.scala 37:46:@2871.4]
  assign _T_56345 = _T_56344[4:0]; // @[Modules.scala 37:46:@2872.4]
  assign _T_56346 = $signed(_T_56345); // @[Modules.scala 37:46:@2873.4]
  assign _T_56349 = $signed(io_in_532) + $signed(io_in_533); // @[Modules.scala 37:46:@2878.4]
  assign _T_56350 = _T_56349[4:0]; // @[Modules.scala 37:46:@2879.4]
  assign _T_56351 = $signed(_T_56350); // @[Modules.scala 37:46:@2880.4]
  assign _T_56352 = $signed(io_in_534) + $signed(io_in_535); // @[Modules.scala 37:46:@2882.4]
  assign _T_56353 = _T_56352[4:0]; // @[Modules.scala 37:46:@2883.4]
  assign _T_56354 = $signed(_T_56353); // @[Modules.scala 37:46:@2884.4]
  assign _T_56355 = $signed(io_in_536) + $signed(io_in_537); // @[Modules.scala 37:46:@2886.4]
  assign _T_56356 = _T_56355[4:0]; // @[Modules.scala 37:46:@2887.4]
  assign _T_56357 = $signed(_T_56356); // @[Modules.scala 37:46:@2888.4]
  assign _T_56358 = $signed(io_in_538) + $signed(io_in_539); // @[Modules.scala 37:46:@2890.4]
  assign _T_56359 = _T_56358[4:0]; // @[Modules.scala 37:46:@2891.4]
  assign _T_56360 = $signed(_T_56359); // @[Modules.scala 37:46:@2892.4]
  assign _T_56361 = $signed(io_in_540) + $signed(io_in_541); // @[Modules.scala 37:46:@2894.4]
  assign _T_56362 = _T_56361[4:0]; // @[Modules.scala 37:46:@2895.4]
  assign _T_56363 = $signed(_T_56362); // @[Modules.scala 37:46:@2896.4]
  assign _T_56364 = $signed(io_in_542) + $signed(io_in_543); // @[Modules.scala 37:46:@2898.4]
  assign _T_56365 = _T_56364[4:0]; // @[Modules.scala 37:46:@2899.4]
  assign _T_56366 = $signed(_T_56365); // @[Modules.scala 37:46:@2900.4]
  assign _T_56367 = $signed(io_in_544) + $signed(io_in_545); // @[Modules.scala 37:46:@2902.4]
  assign _T_56368 = _T_56367[4:0]; // @[Modules.scala 37:46:@2903.4]
  assign _T_56369 = $signed(_T_56368); // @[Modules.scala 37:46:@2904.4]
  assign _T_56370 = $signed(io_in_548) + $signed(io_in_549); // @[Modules.scala 37:46:@2907.4]
  assign _T_56371 = _T_56370[4:0]; // @[Modules.scala 37:46:@2908.4]
  assign _T_56372 = $signed(_T_56371); // @[Modules.scala 37:46:@2909.4]
  assign _T_56373 = $signed(io_in_550) + $signed(io_in_551); // @[Modules.scala 37:46:@2911.4]
  assign _T_56374 = _T_56373[4:0]; // @[Modules.scala 37:46:@2912.4]
  assign _T_56375 = $signed(_T_56374); // @[Modules.scala 37:46:@2913.4]
  assign _T_56378 = $signed(io_in_562) + $signed(io_in_563); // @[Modules.scala 37:46:@2920.4]
  assign _T_56379 = _T_56378[4:0]; // @[Modules.scala 37:46:@2921.4]
  assign _T_56380 = $signed(_T_56379); // @[Modules.scala 37:46:@2922.4]
  assign _T_56381 = $signed(io_in_564) + $signed(io_in_565); // @[Modules.scala 37:46:@2924.4]
  assign _T_56382 = _T_56381[4:0]; // @[Modules.scala 37:46:@2925.4]
  assign _T_56383 = $signed(_T_56382); // @[Modules.scala 37:46:@2926.4]
  assign _T_56384 = $signed(io_in_568) + $signed(io_in_569); // @[Modules.scala 37:46:@2929.4]
  assign _T_56385 = _T_56384[4:0]; // @[Modules.scala 37:46:@2930.4]
  assign _T_56386 = $signed(_T_56385); // @[Modules.scala 37:46:@2931.4]
  assign _T_56387 = $signed(io_in_570) + $signed(io_in_571); // @[Modules.scala 37:46:@2933.4]
  assign _T_56388 = _T_56387[4:0]; // @[Modules.scala 37:46:@2934.4]
  assign _T_56389 = $signed(_T_56388); // @[Modules.scala 37:46:@2935.4]
  assign _T_56390 = $signed(io_in_572) + $signed(io_in_573); // @[Modules.scala 37:46:@2937.4]
  assign _T_56391 = _T_56390[4:0]; // @[Modules.scala 37:46:@2938.4]
  assign _T_56392 = $signed(_T_56391); // @[Modules.scala 37:46:@2939.4]
  assign _T_56393 = $signed(io_in_574) + $signed(io_in_575); // @[Modules.scala 37:46:@2941.4]
  assign _T_56394 = _T_56393[4:0]; // @[Modules.scala 37:46:@2942.4]
  assign _T_56395 = $signed(_T_56394); // @[Modules.scala 37:46:@2943.4]
  assign _T_56396 = $signed(io_in_578) + $signed(io_in_579); // @[Modules.scala 37:46:@2946.4]
  assign _T_56397 = _T_56396[4:0]; // @[Modules.scala 37:46:@2947.4]
  assign _T_56398 = $signed(_T_56397); // @[Modules.scala 37:46:@2948.4]
  assign _T_56401 = $signed(io_in_590) + $signed(io_in_591); // @[Modules.scala 37:46:@2955.4]
  assign _T_56402 = _T_56401[4:0]; // @[Modules.scala 37:46:@2956.4]
  assign _T_56403 = $signed(_T_56402); // @[Modules.scala 37:46:@2957.4]
  assign _T_56404 = $signed(io_in_592) + $signed(io_in_593); // @[Modules.scala 37:46:@2959.4]
  assign _T_56405 = _T_56404[4:0]; // @[Modules.scala 37:46:@2960.4]
  assign _T_56406 = $signed(_T_56405); // @[Modules.scala 37:46:@2961.4]
  assign _T_56407 = $signed(io_in_598) + $signed(io_in_599); // @[Modules.scala 37:46:@2965.4]
  assign _T_56408 = _T_56407[4:0]; // @[Modules.scala 37:46:@2966.4]
  assign _T_56409 = $signed(_T_56408); // @[Modules.scala 37:46:@2967.4]
  assign _T_56413 = $signed(io_in_602) + $signed(io_in_603); // @[Modules.scala 37:46:@2973.4]
  assign _T_56414 = _T_56413[4:0]; // @[Modules.scala 37:46:@2974.4]
  assign _T_56415 = $signed(_T_56414); // @[Modules.scala 37:46:@2975.4]
  assign _T_56430 = $signed(io_in_624) + $signed(io_in_625); // @[Modules.scala 37:46:@2996.4]
  assign _T_56431 = _T_56430[4:0]; // @[Modules.scala 37:46:@2997.4]
  assign _T_56432 = $signed(_T_56431); // @[Modules.scala 37:46:@2998.4]
  assign _T_56433 = $signed(io_in_626) + $signed(io_in_627); // @[Modules.scala 37:46:@3000.4]
  assign _T_56434 = _T_56433[4:0]; // @[Modules.scala 37:46:@3001.4]
  assign _T_56435 = $signed(_T_56434); // @[Modules.scala 37:46:@3002.4]
  assign _T_56436 = $signed(io_in_628) + $signed(io_in_629); // @[Modules.scala 37:46:@3004.4]
  assign _T_56437 = _T_56436[4:0]; // @[Modules.scala 37:46:@3005.4]
  assign _T_56438 = $signed(_T_56437); // @[Modules.scala 37:46:@3006.4]
  assign _T_56439 = $signed(io_in_630) + $signed(io_in_631); // @[Modules.scala 37:46:@3008.4]
  assign _T_56440 = _T_56439[4:0]; // @[Modules.scala 37:46:@3009.4]
  assign _T_56441 = $signed(_T_56440); // @[Modules.scala 37:46:@3010.4]
  assign _T_56442 = $signed(io_in_632) + $signed(io_in_633); // @[Modules.scala 37:46:@3012.4]
  assign _T_56443 = _T_56442[4:0]; // @[Modules.scala 37:46:@3013.4]
  assign _T_56444 = $signed(_T_56443); // @[Modules.scala 37:46:@3014.4]
  assign _T_56445 = $signed(io_in_636) + $signed(io_in_637); // @[Modules.scala 37:46:@3017.4]
  assign _T_56446 = _T_56445[4:0]; // @[Modules.scala 37:46:@3018.4]
  assign _T_56447 = $signed(_T_56446); // @[Modules.scala 37:46:@3019.4]
  assign _T_56449 = $signed(io_in_642) + $signed(io_in_643); // @[Modules.scala 37:46:@3023.4]
  assign _T_56450 = _T_56449[4:0]; // @[Modules.scala 37:46:@3024.4]
  assign _T_56451 = $signed(_T_56450); // @[Modules.scala 37:46:@3025.4]
  assign _T_56456 = $signed(io_in_648) + $signed(io_in_649); // @[Modules.scala 37:46:@3032.4]
  assign _T_56457 = _T_56456[4:0]; // @[Modules.scala 37:46:@3033.4]
  assign _T_56458 = $signed(_T_56457); // @[Modules.scala 37:46:@3034.4]
  assign _T_56459 = $signed(io_in_650) + $signed(io_in_651); // @[Modules.scala 37:46:@3036.4]
  assign _T_56460 = _T_56459[4:0]; // @[Modules.scala 37:46:@3037.4]
  assign _T_56461 = $signed(_T_56460); // @[Modules.scala 37:46:@3038.4]
  assign _T_56462 = $signed(io_in_652) + $signed(io_in_653); // @[Modules.scala 37:46:@3040.4]
  assign _T_56463 = _T_56462[4:0]; // @[Modules.scala 37:46:@3041.4]
  assign _T_56464 = $signed(_T_56463); // @[Modules.scala 37:46:@3042.4]
  assign _T_56465 = $signed(io_in_654) + $signed(io_in_655); // @[Modules.scala 37:46:@3044.4]
  assign _T_56466 = _T_56465[4:0]; // @[Modules.scala 37:46:@3045.4]
  assign _T_56467 = $signed(_T_56466); // @[Modules.scala 37:46:@3046.4]
  assign _T_56468 = $signed(io_in_656) + $signed(io_in_657); // @[Modules.scala 37:46:@3048.4]
  assign _T_56469 = _T_56468[4:0]; // @[Modules.scala 37:46:@3049.4]
  assign _T_56470 = $signed(_T_56469); // @[Modules.scala 37:46:@3050.4]
  assign _T_56471 = $signed(io_in_658) + $signed(io_in_659); // @[Modules.scala 37:46:@3052.4]
  assign _T_56472 = _T_56471[4:0]; // @[Modules.scala 37:46:@3053.4]
  assign _T_56473 = $signed(_T_56472); // @[Modules.scala 37:46:@3054.4]
  assign _T_56475 = $signed(io_in_662) + $signed(io_in_663); // @[Modules.scala 37:46:@3057.4]
  assign _T_56476 = _T_56475[4:0]; // @[Modules.scala 37:46:@3058.4]
  assign _T_56477 = $signed(_T_56476); // @[Modules.scala 37:46:@3059.4]
  assign _T_56483 = $signed(io_in_674) + $signed(io_in_675); // @[Modules.scala 37:46:@3066.4]
  assign _T_56484 = _T_56483[4:0]; // @[Modules.scala 37:46:@3067.4]
  assign _T_56485 = $signed(_T_56484); // @[Modules.scala 37:46:@3068.4]
  assign _T_56492 = $signed(io_in_682) + $signed(io_in_683); // @[Modules.scala 37:46:@3079.4]
  assign _T_56493 = _T_56492[4:0]; // @[Modules.scala 37:46:@3080.4]
  assign _T_56494 = $signed(_T_56493); // @[Modules.scala 37:46:@3081.4]
  assign _T_56495 = $signed(io_in_684) + $signed(io_in_685); // @[Modules.scala 37:46:@3083.4]
  assign _T_56496 = _T_56495[4:0]; // @[Modules.scala 37:46:@3084.4]
  assign _T_56497 = $signed(_T_56496); // @[Modules.scala 37:46:@3085.4]
  assign _T_56500 = $signed(io_in_700) + $signed(io_in_701); // @[Modules.scala 37:46:@3094.4]
  assign _T_56501 = _T_56500[4:0]; // @[Modules.scala 37:46:@3095.4]
  assign _T_56502 = $signed(_T_56501); // @[Modules.scala 37:46:@3096.4]
  assign _T_56503 = $signed(io_in_702) + $signed(io_in_703); // @[Modules.scala 37:46:@3098.4]
  assign _T_56504 = _T_56503[4:0]; // @[Modules.scala 37:46:@3099.4]
  assign _T_56505 = $signed(_T_56504); // @[Modules.scala 37:46:@3100.4]
  assign _T_56519 = $signed(io_in_724) + $signed(io_in_725); // @[Modules.scala 37:46:@3121.4]
  assign _T_56520 = _T_56519[4:0]; // @[Modules.scala 37:46:@3122.4]
  assign _T_56521 = $signed(_T_56520); // @[Modules.scala 37:46:@3123.4]
  assign _T_56541 = $signed(io_in_758) + $signed(io_in_759); // @[Modules.scala 37:46:@3150.4]
  assign _T_56542 = _T_56541[4:0]; // @[Modules.scala 37:46:@3151.4]
  assign _T_56543 = $signed(_T_56542); // @[Modules.scala 37:46:@3152.4]
  assign _T_56544 = $signed(io_in_760) + $signed(io_in_761); // @[Modules.scala 37:46:@3154.4]
  assign _T_56545 = _T_56544[4:0]; // @[Modules.scala 37:46:@3155.4]
  assign _T_56546 = $signed(_T_56545); // @[Modules.scala 37:46:@3156.4]
  assign _T_56547 = $signed(io_in_762) + $signed(io_in_763); // @[Modules.scala 37:46:@3158.4]
  assign _T_56548 = _T_56547[4:0]; // @[Modules.scala 37:46:@3159.4]
  assign _T_56549 = $signed(_T_56548); // @[Modules.scala 37:46:@3160.4]
  assign _T_56551 = $signed(io_in_766) + $signed(io_in_767); // @[Modules.scala 37:46:@3163.4]
  assign _T_56552 = _T_56551[4:0]; // @[Modules.scala 37:46:@3164.4]
  assign _T_56553 = $signed(_T_56552); // @[Modules.scala 37:46:@3165.4]
  assign buffer_1_2 = {{6{_T_55958[4]}},_T_55958}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_3 = {{6{_T_55961[4]}},_T_55961}; // @[Modules.scala 32:22:@8.4]
  assign _T_56564 = $signed(buffer_1_2) + $signed(buffer_1_3); // @[Modules.scala 65:57:@3179.4]
  assign _T_56565 = _T_56564[10:0]; // @[Modules.scala 65:57:@3180.4]
  assign buffer_1_393 = $signed(_T_56565); // @[Modules.scala 65:57:@3181.4]
  assign buffer_1_4 = {{6{_T_55964[4]}},_T_55964}; // @[Modules.scala 32:22:@8.4]
  assign _T_56567 = $signed(buffer_1_4) + $signed(11'sh0); // @[Modules.scala 65:57:@3183.4]
  assign _T_56568 = _T_56567[10:0]; // @[Modules.scala 65:57:@3184.4]
  assign buffer_1_394 = $signed(_T_56568); // @[Modules.scala 65:57:@3185.4]
  assign buffer_1_6 = {{6{_T_55968[4]}},_T_55968}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_7 = {{6{_T_55971[4]}},_T_55971}; // @[Modules.scala 32:22:@8.4]
  assign _T_56570 = $signed(buffer_1_6) + $signed(buffer_1_7); // @[Modules.scala 65:57:@3187.4]
  assign _T_56571 = _T_56570[10:0]; // @[Modules.scala 65:57:@3188.4]
  assign buffer_1_395 = $signed(_T_56571); // @[Modules.scala 65:57:@3189.4]
  assign buffer_1_8 = {{6{io_in_16[4]}},io_in_16}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_9 = {{6{io_in_18[4]}},io_in_18}; // @[Modules.scala 32:22:@8.4]
  assign _T_56573 = $signed(buffer_1_8) + $signed(buffer_1_9); // @[Modules.scala 65:57:@3191.4]
  assign _T_56574 = _T_56573[10:0]; // @[Modules.scala 65:57:@3192.4]
  assign buffer_1_396 = $signed(_T_56574); // @[Modules.scala 65:57:@3193.4]
  assign buffer_1_11 = {{6{io_in_22[4]}},io_in_22}; // @[Modules.scala 32:22:@8.4]
  assign _T_56576 = $signed(buffer_0_10) + $signed(buffer_1_11); // @[Modules.scala 65:57:@3195.4]
  assign _T_56577 = _T_56576[10:0]; // @[Modules.scala 65:57:@3196.4]
  assign buffer_1_397 = $signed(_T_56577); // @[Modules.scala 65:57:@3197.4]
  assign buffer_1_12 = {{6{_T_55977[4]}},_T_55977}; // @[Modules.scala 32:22:@8.4]
  assign _T_56579 = $signed(buffer_1_12) + $signed(11'sh0); // @[Modules.scala 65:57:@3199.4]
  assign _T_56580 = _T_56579[10:0]; // @[Modules.scala 65:57:@3200.4]
  assign buffer_1_398 = $signed(_T_56580); // @[Modules.scala 65:57:@3201.4]
  assign buffer_1_14 = {{6{io_in_28[4]}},io_in_28}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_15 = {{6{_T_55981[4]}},_T_55981}; // @[Modules.scala 32:22:@8.4]
  assign _T_56582 = $signed(buffer_1_14) + $signed(buffer_1_15); // @[Modules.scala 65:57:@3203.4]
  assign _T_56583 = _T_56582[10:0]; // @[Modules.scala 65:57:@3204.4]
  assign buffer_1_399 = $signed(_T_56583); // @[Modules.scala 65:57:@3205.4]
  assign buffer_1_17 = {{6{_T_55987[4]}},_T_55987}; // @[Modules.scala 32:22:@8.4]
  assign _T_56585 = $signed(buffer_0_16) + $signed(buffer_1_17); // @[Modules.scala 65:57:@3207.4]
  assign _T_56586 = _T_56585[10:0]; // @[Modules.scala 65:57:@3208.4]
  assign buffer_1_400 = $signed(_T_56586); // @[Modules.scala 65:57:@3209.4]
  assign buffer_1_18 = {{6{_T_55990[4]}},_T_55990}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_19 = {{6{_T_55993[4]}},_T_55993}; // @[Modules.scala 32:22:@8.4]
  assign _T_56588 = $signed(buffer_1_18) + $signed(buffer_1_19); // @[Modules.scala 65:57:@3211.4]
  assign _T_56589 = _T_56588[10:0]; // @[Modules.scala 65:57:@3212.4]
  assign buffer_1_401 = $signed(_T_56589); // @[Modules.scala 65:57:@3213.4]
  assign buffer_1_20 = {{6{_T_55996[4]}},_T_55996}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_21 = {{6{_T_55999[4]}},_T_55999}; // @[Modules.scala 32:22:@8.4]
  assign _T_56591 = $signed(buffer_1_20) + $signed(buffer_1_21); // @[Modules.scala 65:57:@3215.4]
  assign _T_56592 = _T_56591[10:0]; // @[Modules.scala 65:57:@3216.4]
  assign buffer_1_402 = $signed(_T_56592); // @[Modules.scala 65:57:@3217.4]
  assign buffer_1_22 = {{6{io_in_45[4]}},io_in_45}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_23 = {{6{_T_56002[4]}},_T_56002}; // @[Modules.scala 32:22:@8.4]
  assign _T_56594 = $signed(buffer_1_22) + $signed(buffer_1_23); // @[Modules.scala 65:57:@3219.4]
  assign _T_56595 = _T_56594[10:0]; // @[Modules.scala 65:57:@3220.4]
  assign buffer_1_403 = $signed(_T_56595); // @[Modules.scala 65:57:@3221.4]
  assign buffer_1_24 = {{6{_T_56005[4]}},_T_56005}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_25 = {{6{_T_56008[4]}},_T_56008}; // @[Modules.scala 32:22:@8.4]
  assign _T_56597 = $signed(buffer_1_24) + $signed(buffer_1_25); // @[Modules.scala 65:57:@3223.4]
  assign _T_56598 = _T_56597[10:0]; // @[Modules.scala 65:57:@3224.4]
  assign buffer_1_404 = $signed(_T_56598); // @[Modules.scala 65:57:@3225.4]
  assign buffer_1_26 = {{6{io_in_52[4]}},io_in_52}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_27 = {{6{io_in_55[4]}},io_in_55}; // @[Modules.scala 32:22:@8.4]
  assign _T_56600 = $signed(buffer_1_26) + $signed(buffer_1_27); // @[Modules.scala 65:57:@3227.4]
  assign _T_56601 = _T_56600[10:0]; // @[Modules.scala 65:57:@3228.4]
  assign buffer_1_405 = $signed(_T_56601); // @[Modules.scala 65:57:@3229.4]
  assign buffer_1_28 = {{6{io_in_57[4]}},io_in_57}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_29 = {{6{_T_56011[4]}},_T_56011}; // @[Modules.scala 32:22:@8.4]
  assign _T_56603 = $signed(buffer_1_28) + $signed(buffer_1_29); // @[Modules.scala 65:57:@3231.4]
  assign _T_56604 = _T_56603[10:0]; // @[Modules.scala 65:57:@3232.4]
  assign buffer_1_406 = $signed(_T_56604); // @[Modules.scala 65:57:@3233.4]
  assign buffer_1_30 = {{6{_T_56014[4]}},_T_56014}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_31 = {{6{_T_56017[4]}},_T_56017}; // @[Modules.scala 32:22:@8.4]
  assign _T_56606 = $signed(buffer_1_30) + $signed(buffer_1_31); // @[Modules.scala 65:57:@3235.4]
  assign _T_56607 = _T_56606[10:0]; // @[Modules.scala 65:57:@3236.4]
  assign buffer_1_407 = $signed(_T_56607); // @[Modules.scala 65:57:@3237.4]
  assign buffer_1_32 = {{6{_T_56020[4]}},_T_56020}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_33 = {{6{_T_56023[4]}},_T_56023}; // @[Modules.scala 32:22:@8.4]
  assign _T_56609 = $signed(buffer_1_32) + $signed(buffer_1_33); // @[Modules.scala 65:57:@3239.4]
  assign _T_56610 = _T_56609[10:0]; // @[Modules.scala 65:57:@3240.4]
  assign buffer_1_408 = $signed(_T_56610); // @[Modules.scala 65:57:@3241.4]
  assign buffer_1_34 = {{6{_T_56026[4]}},_T_56026}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_35 = {{6{_T_56029[4]}},_T_56029}; // @[Modules.scala 32:22:@8.4]
  assign _T_56612 = $signed(buffer_1_34) + $signed(buffer_1_35); // @[Modules.scala 65:57:@3243.4]
  assign _T_56613 = _T_56612[10:0]; // @[Modules.scala 65:57:@3244.4]
  assign buffer_1_409 = $signed(_T_56613); // @[Modules.scala 65:57:@3245.4]
  assign buffer_1_36 = {{6{_T_56032[4]}},_T_56032}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_37 = {{6{_T_56035[4]}},_T_56035}; // @[Modules.scala 32:22:@8.4]
  assign _T_56615 = $signed(buffer_1_36) + $signed(buffer_1_37); // @[Modules.scala 65:57:@3247.4]
  assign _T_56616 = _T_56615[10:0]; // @[Modules.scala 65:57:@3248.4]
  assign buffer_1_410 = $signed(_T_56616); // @[Modules.scala 65:57:@3249.4]
  assign buffer_1_38 = {{6{_T_56038[4]}},_T_56038}; // @[Modules.scala 32:22:@8.4]
  assign _T_56618 = $signed(buffer_1_38) + $signed(buffer_0_39); // @[Modules.scala 65:57:@3251.4]
  assign _T_56619 = _T_56618[10:0]; // @[Modules.scala 65:57:@3252.4]
  assign buffer_1_411 = $signed(_T_56619); // @[Modules.scala 65:57:@3253.4]
  assign buffer_1_40 = {{6{_T_56044[4]}},_T_56044}; // @[Modules.scala 32:22:@8.4]
  assign _T_56621 = $signed(buffer_1_40) + $signed(11'sh0); // @[Modules.scala 65:57:@3255.4]
  assign _T_56622 = _T_56621[10:0]; // @[Modules.scala 65:57:@3256.4]
  assign buffer_1_412 = $signed(_T_56622); // @[Modules.scala 65:57:@3257.4]
  assign buffer_1_42 = {{6{io_in_85[4]}},io_in_85}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_43 = {{6{io_in_87[4]}},io_in_87}; // @[Modules.scala 32:22:@8.4]
  assign _T_56624 = $signed(buffer_1_42) + $signed(buffer_1_43); // @[Modules.scala 65:57:@3259.4]
  assign _T_56625 = _T_56624[10:0]; // @[Modules.scala 65:57:@3260.4]
  assign buffer_1_413 = $signed(_T_56625); // @[Modules.scala 65:57:@3261.4]
  assign buffer_1_46 = {{6{_T_56054[4]}},_T_56054}; // @[Modules.scala 32:22:@8.4]
  assign _T_56630 = $signed(buffer_1_46) + $signed(buffer_0_47); // @[Modules.scala 65:57:@3267.4]
  assign _T_56631 = _T_56630[10:0]; // @[Modules.scala 65:57:@3268.4]
  assign buffer_1_415 = $signed(_T_56631); // @[Modules.scala 65:57:@3269.4]
  assign buffer_1_48 = {{6{_T_56060[4]}},_T_56060}; // @[Modules.scala 32:22:@8.4]
  assign _T_56633 = $signed(buffer_1_48) + $signed(buffer_0_49); // @[Modules.scala 65:57:@3271.4]
  assign _T_56634 = _T_56633[10:0]; // @[Modules.scala 65:57:@3272.4]
  assign buffer_1_416 = $signed(_T_56634); // @[Modules.scala 65:57:@3273.4]
  assign buffer_1_54 = {{6{_T_56078[4]}},_T_56078}; // @[Modules.scala 32:22:@8.4]
  assign _T_56642 = $signed(buffer_1_54) + $signed(buffer_0_55); // @[Modules.scala 65:57:@3283.4]
  assign _T_56643 = _T_56642[10:0]; // @[Modules.scala 65:57:@3284.4]
  assign buffer_1_419 = $signed(_T_56643); // @[Modules.scala 65:57:@3285.4]
  assign buffer_1_57 = {{6{io_in_115[4]}},io_in_115}; // @[Modules.scala 32:22:@8.4]
  assign _T_56645 = $signed(11'sh0) + $signed(buffer_1_57); // @[Modules.scala 65:57:@3287.4]
  assign _T_56646 = _T_56645[10:0]; // @[Modules.scala 65:57:@3288.4]
  assign buffer_1_420 = $signed(_T_56646); // @[Modules.scala 65:57:@3289.4]
  assign _T_56648 = $signed(buffer_0_58) + $signed(11'sh0); // @[Modules.scala 65:57:@3291.4]
  assign _T_56649 = _T_56648[10:0]; // @[Modules.scala 65:57:@3292.4]
  assign buffer_1_421 = $signed(_T_56649); // @[Modules.scala 65:57:@3293.4]
  assign buffer_1_63 = {{6{io_in_127[4]}},io_in_127}; // @[Modules.scala 32:22:@8.4]
  assign _T_56654 = $signed(11'sh0) + $signed(buffer_1_63); // @[Modules.scala 65:57:@3299.4]
  assign _T_56655 = _T_56654[10:0]; // @[Modules.scala 65:57:@3300.4]
  assign buffer_1_423 = $signed(_T_56655); // @[Modules.scala 65:57:@3301.4]
  assign buffer_1_64 = {{6{_T_56089[4]}},_T_56089}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_65 = {{6{_T_56092[4]}},_T_56092}; // @[Modules.scala 32:22:@8.4]
  assign _T_56657 = $signed(buffer_1_64) + $signed(buffer_1_65); // @[Modules.scala 65:57:@3303.4]
  assign _T_56658 = _T_56657[10:0]; // @[Modules.scala 65:57:@3304.4]
  assign buffer_1_424 = $signed(_T_56658); // @[Modules.scala 65:57:@3305.4]
  assign buffer_1_66 = {{6{io_in_133[4]}},io_in_133}; // @[Modules.scala 32:22:@8.4]
  assign _T_56660 = $signed(buffer_1_66) + $signed(buffer_0_67); // @[Modules.scala 65:57:@3307.4]
  assign _T_56661 = _T_56660[10:0]; // @[Modules.scala 65:57:@3308.4]
  assign buffer_1_425 = $signed(_T_56661); // @[Modules.scala 65:57:@3309.4]
  assign buffer_1_68 = {{6{_T_56098[4]}},_T_56098}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_69 = {{6{io_in_139[4]}},io_in_139}; // @[Modules.scala 32:22:@8.4]
  assign _T_56663 = $signed(buffer_1_68) + $signed(buffer_1_69); // @[Modules.scala 65:57:@3311.4]
  assign _T_56664 = _T_56663[10:0]; // @[Modules.scala 65:57:@3312.4]
  assign buffer_1_426 = $signed(_T_56664); // @[Modules.scala 65:57:@3313.4]
  assign buffer_1_70 = {{6{io_in_140[4]}},io_in_140}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_71 = {{6{io_in_143[4]}},io_in_143}; // @[Modules.scala 32:22:@8.4]
  assign _T_56666 = $signed(buffer_1_70) + $signed(buffer_1_71); // @[Modules.scala 65:57:@3315.4]
  assign _T_56667 = _T_56666[10:0]; // @[Modules.scala 65:57:@3316.4]
  assign buffer_1_427 = $signed(_T_56667); // @[Modules.scala 65:57:@3317.4]
  assign buffer_1_74 = {{6{io_in_148[4]}},io_in_148}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_75 = {{6{io_in_150[4]}},io_in_150}; // @[Modules.scala 32:22:@8.4]
  assign _T_56672 = $signed(buffer_1_74) + $signed(buffer_1_75); // @[Modules.scala 65:57:@3323.4]
  assign _T_56673 = _T_56672[10:0]; // @[Modules.scala 65:57:@3324.4]
  assign buffer_1_429 = $signed(_T_56673); // @[Modules.scala 65:57:@3325.4]
  assign buffer_1_78 = {{6{io_in_156[4]}},io_in_156}; // @[Modules.scala 32:22:@8.4]
  assign _T_56678 = $signed(buffer_1_78) + $signed(11'sh0); // @[Modules.scala 65:57:@3331.4]
  assign _T_56679 = _T_56678[10:0]; // @[Modules.scala 65:57:@3332.4]
  assign buffer_1_431 = $signed(_T_56679); // @[Modules.scala 65:57:@3333.4]
  assign buffer_1_81 = {{6{io_in_163[4]}},io_in_163}; // @[Modules.scala 32:22:@8.4]
  assign _T_56681 = $signed(11'sh0) + $signed(buffer_1_81); // @[Modules.scala 65:57:@3335.4]
  assign _T_56682 = _T_56681[10:0]; // @[Modules.scala 65:57:@3336.4]
  assign buffer_1_432 = $signed(_T_56682); // @[Modules.scala 65:57:@3337.4]
  assign buffer_1_83 = {{6{_T_56108[4]}},_T_56108}; // @[Modules.scala 32:22:@8.4]
  assign _T_56684 = $signed(11'sh0) + $signed(buffer_1_83); // @[Modules.scala 65:57:@3339.4]
  assign _T_56685 = _T_56684[10:0]; // @[Modules.scala 65:57:@3340.4]
  assign buffer_1_433 = $signed(_T_56685); // @[Modules.scala 65:57:@3341.4]
  assign buffer_1_84 = {{6{io_in_169[4]}},io_in_169}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_85 = {{6{_T_56111[4]}},_T_56111}; // @[Modules.scala 32:22:@8.4]
  assign _T_56687 = $signed(buffer_1_84) + $signed(buffer_1_85); // @[Modules.scala 65:57:@3343.4]
  assign _T_56688 = _T_56687[10:0]; // @[Modules.scala 65:57:@3344.4]
  assign buffer_1_434 = $signed(_T_56688); // @[Modules.scala 65:57:@3345.4]
  assign buffer_1_87 = {{6{_T_56114[4]}},_T_56114}; // @[Modules.scala 32:22:@8.4]
  assign _T_56690 = $signed(buffer_0_86) + $signed(buffer_1_87); // @[Modules.scala 65:57:@3347.4]
  assign _T_56691 = _T_56690[10:0]; // @[Modules.scala 65:57:@3348.4]
  assign buffer_1_435 = $signed(_T_56691); // @[Modules.scala 65:57:@3349.4]
  assign buffer_1_88 = {{6{_T_56117[4]}},_T_56117}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_89 = {{6{io_in_178[4]}},io_in_178}; // @[Modules.scala 32:22:@8.4]
  assign _T_56693 = $signed(buffer_1_88) + $signed(buffer_1_89); // @[Modules.scala 65:57:@3351.4]
  assign _T_56694 = _T_56693[10:0]; // @[Modules.scala 65:57:@3352.4]
  assign buffer_1_436 = $signed(_T_56694); // @[Modules.scala 65:57:@3353.4]
  assign buffer_1_91 = {{6{io_in_182[4]}},io_in_182}; // @[Modules.scala 32:22:@8.4]
  assign _T_56696 = $signed(11'sh0) + $signed(buffer_1_91); // @[Modules.scala 65:57:@3355.4]
  assign _T_56697 = _T_56696[10:0]; // @[Modules.scala 65:57:@3356.4]
  assign buffer_1_437 = $signed(_T_56697); // @[Modules.scala 65:57:@3357.4]
  assign buffer_1_94 = {{6{io_in_188[4]}},io_in_188}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_95 = {{6{io_in_191[4]}},io_in_191}; // @[Modules.scala 32:22:@8.4]
  assign _T_56702 = $signed(buffer_1_94) + $signed(buffer_1_95); // @[Modules.scala 65:57:@3363.4]
  assign _T_56703 = _T_56702[10:0]; // @[Modules.scala 65:57:@3364.4]
  assign buffer_1_439 = $signed(_T_56703); // @[Modules.scala 65:57:@3365.4]
  assign buffer_1_96 = {{6{io_in_193[4]}},io_in_193}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_97 = {{6{io_in_195[4]}},io_in_195}; // @[Modules.scala 32:22:@8.4]
  assign _T_56705 = $signed(buffer_1_96) + $signed(buffer_1_97); // @[Modules.scala 65:57:@3367.4]
  assign _T_56706 = _T_56705[10:0]; // @[Modules.scala 65:57:@3368.4]
  assign buffer_1_440 = $signed(_T_56706); // @[Modules.scala 65:57:@3369.4]
  assign buffer_1_98 = {{6{_T_56125[4]}},_T_56125}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_99 = {{6{io_in_199[4]}},io_in_199}; // @[Modules.scala 32:22:@8.4]
  assign _T_56708 = $signed(buffer_1_98) + $signed(buffer_1_99); // @[Modules.scala 65:57:@3371.4]
  assign _T_56709 = _T_56708[10:0]; // @[Modules.scala 65:57:@3372.4]
  assign buffer_1_441 = $signed(_T_56709); // @[Modules.scala 65:57:@3373.4]
  assign buffer_1_100 = {{6{io_in_201[4]}},io_in_201}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_101 = {{6{_T_56128[4]}},_T_56128}; // @[Modules.scala 32:22:@8.4]
  assign _T_56711 = $signed(buffer_1_100) + $signed(buffer_1_101); // @[Modules.scala 65:57:@3375.4]
  assign _T_56712 = _T_56711[10:0]; // @[Modules.scala 65:57:@3376.4]
  assign buffer_1_442 = $signed(_T_56712); // @[Modules.scala 65:57:@3377.4]
  assign buffer_1_102 = {{6{io_in_205[4]}},io_in_205}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_103 = {{6{io_in_206[4]}},io_in_206}; // @[Modules.scala 32:22:@8.4]
  assign _T_56714 = $signed(buffer_1_102) + $signed(buffer_1_103); // @[Modules.scala 65:57:@3379.4]
  assign _T_56715 = _T_56714[10:0]; // @[Modules.scala 65:57:@3380.4]
  assign buffer_1_443 = $signed(_T_56715); // @[Modules.scala 65:57:@3381.4]
  assign buffer_1_104 = {{6{io_in_208[4]}},io_in_208}; // @[Modules.scala 32:22:@8.4]
  assign _T_56717 = $signed(buffer_1_104) + $signed(buffer_0_105); // @[Modules.scala 65:57:@3383.4]
  assign _T_56718 = _T_56717[10:0]; // @[Modules.scala 65:57:@3384.4]
  assign buffer_1_444 = $signed(_T_56718); // @[Modules.scala 65:57:@3385.4]
  assign buffer_1_106 = {{6{io_in_213[4]}},io_in_213}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_107 = {{6{io_in_215[4]}},io_in_215}; // @[Modules.scala 32:22:@8.4]
  assign _T_56720 = $signed(buffer_1_106) + $signed(buffer_1_107); // @[Modules.scala 65:57:@3387.4]
  assign _T_56721 = _T_56720[10:0]; // @[Modules.scala 65:57:@3388.4]
  assign buffer_1_445 = $signed(_T_56721); // @[Modules.scala 65:57:@3389.4]
  assign buffer_1_108 = {{6{io_in_217[4]}},io_in_217}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_109 = {{6{io_in_219[4]}},io_in_219}; // @[Modules.scala 32:22:@8.4]
  assign _T_56723 = $signed(buffer_1_108) + $signed(buffer_1_109); // @[Modules.scala 65:57:@3391.4]
  assign _T_56724 = _T_56723[10:0]; // @[Modules.scala 65:57:@3392.4]
  assign buffer_1_446 = $signed(_T_56724); // @[Modules.scala 65:57:@3393.4]
  assign buffer_1_110 = {{6{_T_56134[4]}},_T_56134}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_111 = {{6{io_in_223[4]}},io_in_223}; // @[Modules.scala 32:22:@8.4]
  assign _T_56726 = $signed(buffer_1_110) + $signed(buffer_1_111); // @[Modules.scala 65:57:@3395.4]
  assign _T_56727 = _T_56726[10:0]; // @[Modules.scala 65:57:@3396.4]
  assign buffer_1_447 = $signed(_T_56727); // @[Modules.scala 65:57:@3397.4]
  assign buffer_1_112 = {{6{_T_56137[4]}},_T_56137}; // @[Modules.scala 32:22:@8.4]
  assign _T_56729 = $signed(buffer_1_112) + $signed(11'sh0); // @[Modules.scala 65:57:@3399.4]
  assign _T_56730 = _T_56729[10:0]; // @[Modules.scala 65:57:@3400.4]
  assign buffer_1_448 = $signed(_T_56730); // @[Modules.scala 65:57:@3401.4]
  assign buffer_1_120 = {{6{_T_56147[4]}},_T_56147}; // @[Modules.scala 32:22:@8.4]
  assign _T_56741 = $signed(buffer_1_120) + $signed(11'sh0); // @[Modules.scala 65:57:@3415.4]
  assign _T_56742 = _T_56741[10:0]; // @[Modules.scala 65:57:@3416.4]
  assign buffer_1_452 = $signed(_T_56742); // @[Modules.scala 65:57:@3417.4]
  assign buffer_1_123 = {{6{io_in_247[4]}},io_in_247}; // @[Modules.scala 32:22:@8.4]
  assign _T_56744 = $signed(11'sh0) + $signed(buffer_1_123); // @[Modules.scala 65:57:@3419.4]
  assign _T_56745 = _T_56744[10:0]; // @[Modules.scala 65:57:@3420.4]
  assign buffer_1_453 = $signed(_T_56745); // @[Modules.scala 65:57:@3421.4]
  assign buffer_1_124 = {{6{_T_56152[4]}},_T_56152}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_125 = {{6{_T_56155[4]}},_T_56155}; // @[Modules.scala 32:22:@8.4]
  assign _T_56747 = $signed(buffer_1_124) + $signed(buffer_1_125); // @[Modules.scala 65:57:@3423.4]
  assign _T_56748 = _T_56747[10:0]; // @[Modules.scala 65:57:@3424.4]
  assign buffer_1_454 = $signed(_T_56748); // @[Modules.scala 65:57:@3425.4]
  assign buffer_1_126 = {{6{io_in_253[4]}},io_in_253}; // @[Modules.scala 32:22:@8.4]
  assign _T_56750 = $signed(buffer_1_126) + $signed(11'sh0); // @[Modules.scala 65:57:@3427.4]
  assign _T_56751 = _T_56750[10:0]; // @[Modules.scala 65:57:@3428.4]
  assign buffer_1_455 = $signed(_T_56751); // @[Modules.scala 65:57:@3429.4]
  assign buffer_1_130 = {{6{io_in_260[4]}},io_in_260}; // @[Modules.scala 32:22:@8.4]
  assign _T_56756 = $signed(buffer_1_130) + $signed(11'sh0); // @[Modules.scala 65:57:@3435.4]
  assign _T_56757 = _T_56756[10:0]; // @[Modules.scala 65:57:@3436.4]
  assign buffer_1_457 = $signed(_T_56757); // @[Modules.scala 65:57:@3437.4]
  assign buffer_1_133 = {{6{_T_56163[4]}},_T_56163}; // @[Modules.scala 32:22:@8.4]
  assign _T_56759 = $signed(11'sh0) + $signed(buffer_1_133); // @[Modules.scala 65:57:@3439.4]
  assign _T_56760 = _T_56759[10:0]; // @[Modules.scala 65:57:@3440.4]
  assign buffer_1_458 = $signed(_T_56760); // @[Modules.scala 65:57:@3441.4]
  assign buffer_1_137 = {{6{io_in_275[4]}},io_in_275}; // @[Modules.scala 32:22:@8.4]
  assign _T_56765 = $signed(11'sh0) + $signed(buffer_1_137); // @[Modules.scala 65:57:@3447.4]
  assign _T_56766 = _T_56765[10:0]; // @[Modules.scala 65:57:@3448.4]
  assign buffer_1_460 = $signed(_T_56766); // @[Modules.scala 65:57:@3449.4]
  assign buffer_1_138 = {{6{_T_56169[4]}},_T_56169}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_139 = {{6{_T_56172[4]}},_T_56172}; // @[Modules.scala 32:22:@8.4]
  assign _T_56768 = $signed(buffer_1_138) + $signed(buffer_1_139); // @[Modules.scala 65:57:@3451.4]
  assign _T_56769 = _T_56768[10:0]; // @[Modules.scala 65:57:@3452.4]
  assign buffer_1_461 = $signed(_T_56769); // @[Modules.scala 65:57:@3453.4]
  assign buffer_1_140 = {{6{io_in_281[4]}},io_in_281}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_141 = {{6{io_in_283[4]}},io_in_283}; // @[Modules.scala 32:22:@8.4]
  assign _T_56771 = $signed(buffer_1_140) + $signed(buffer_1_141); // @[Modules.scala 65:57:@3455.4]
  assign _T_56772 = _T_56771[10:0]; // @[Modules.scala 65:57:@3456.4]
  assign buffer_1_462 = $signed(_T_56772); // @[Modules.scala 65:57:@3457.4]
  assign buffer_1_146 = {{6{_T_56178[4]}},_T_56178}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_147 = {{6{io_in_294[4]}},io_in_294}; // @[Modules.scala 32:22:@8.4]
  assign _T_56780 = $signed(buffer_1_146) + $signed(buffer_1_147); // @[Modules.scala 65:57:@3467.4]
  assign _T_56781 = _T_56780[10:0]; // @[Modules.scala 65:57:@3468.4]
  assign buffer_1_465 = $signed(_T_56781); // @[Modules.scala 65:57:@3469.4]
  assign buffer_1_151 = {{6{io_in_303[4]}},io_in_303}; // @[Modules.scala 32:22:@8.4]
  assign _T_56786 = $signed(11'sh0) + $signed(buffer_1_151); // @[Modules.scala 65:57:@3475.4]
  assign _T_56787 = _T_56786[10:0]; // @[Modules.scala 65:57:@3476.4]
  assign buffer_1_467 = $signed(_T_56787); // @[Modules.scala 65:57:@3477.4]
  assign buffer_1_152 = {{6{_T_56184[4]}},_T_56184}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_153 = {{6{_T_56187[4]}},_T_56187}; // @[Modules.scala 32:22:@8.4]
  assign _T_56789 = $signed(buffer_1_152) + $signed(buffer_1_153); // @[Modules.scala 65:57:@3479.4]
  assign _T_56790 = _T_56789[10:0]; // @[Modules.scala 65:57:@3480.4]
  assign buffer_1_468 = $signed(_T_56790); // @[Modules.scala 65:57:@3481.4]
  assign buffer_1_157 = {{6{io_in_314[4]}},io_in_314}; // @[Modules.scala 32:22:@8.4]
  assign _T_56795 = $signed(11'sh0) + $signed(buffer_1_157); // @[Modules.scala 65:57:@3487.4]
  assign _T_56796 = _T_56795[10:0]; // @[Modules.scala 65:57:@3488.4]
  assign buffer_1_470 = $signed(_T_56796); // @[Modules.scala 65:57:@3489.4]
  assign _T_56798 = $signed(11'sh0) + $signed(buffer_0_159); // @[Modules.scala 65:57:@3491.4]
  assign _T_56799 = _T_56798[10:0]; // @[Modules.scala 65:57:@3492.4]
  assign buffer_1_471 = $signed(_T_56799); // @[Modules.scala 65:57:@3493.4]
  assign buffer_1_160 = {{6{_T_56197[4]}},_T_56197}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_161 = {{6{io_in_322[4]}},io_in_322}; // @[Modules.scala 32:22:@8.4]
  assign _T_56801 = $signed(buffer_1_160) + $signed(buffer_1_161); // @[Modules.scala 65:57:@3495.4]
  assign _T_56802 = _T_56801[10:0]; // @[Modules.scala 65:57:@3496.4]
  assign buffer_1_472 = $signed(_T_56802); // @[Modules.scala 65:57:@3497.4]
  assign buffer_1_165 = {{6{io_in_331[4]}},io_in_331}; // @[Modules.scala 32:22:@8.4]
  assign _T_56807 = $signed(11'sh0) + $signed(buffer_1_165); // @[Modules.scala 65:57:@3503.4]
  assign _T_56808 = _T_56807[10:0]; // @[Modules.scala 65:57:@3504.4]
  assign buffer_1_474 = $signed(_T_56808); // @[Modules.scala 65:57:@3505.4]
  assign buffer_1_166 = {{6{_T_56203[4]}},_T_56203}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_167 = {{6{_T_56206[4]}},_T_56206}; // @[Modules.scala 32:22:@8.4]
  assign _T_56810 = $signed(buffer_1_166) + $signed(buffer_1_167); // @[Modules.scala 65:57:@3507.4]
  assign _T_56811 = _T_56810[10:0]; // @[Modules.scala 65:57:@3508.4]
  assign buffer_1_475 = $signed(_T_56811); // @[Modules.scala 65:57:@3509.4]
  assign _T_56822 = $signed(buffer_0_174) + $signed(11'sh0); // @[Modules.scala 65:57:@3523.4]
  assign _T_56823 = _T_56822[10:0]; // @[Modules.scala 65:57:@3524.4]
  assign buffer_1_479 = $signed(_T_56823); // @[Modules.scala 65:57:@3525.4]
  assign buffer_1_179 = {{6{io_in_359[4]}},io_in_359}; // @[Modules.scala 32:22:@8.4]
  assign _T_56828 = $signed(11'sh0) + $signed(buffer_1_179); // @[Modules.scala 65:57:@3531.4]
  assign _T_56829 = _T_56828[10:0]; // @[Modules.scala 65:57:@3532.4]
  assign buffer_1_481 = $signed(_T_56829); // @[Modules.scala 65:57:@3533.4]
  assign buffer_1_180 = {{6{_T_56226[4]}},_T_56226}; // @[Modules.scala 32:22:@8.4]
  assign _T_56831 = $signed(buffer_1_180) + $signed(11'sh0); // @[Modules.scala 65:57:@3535.4]
  assign _T_56832 = _T_56831[10:0]; // @[Modules.scala 65:57:@3536.4]
  assign buffer_1_482 = $signed(_T_56832); // @[Modules.scala 65:57:@3537.4]
  assign buffer_1_184 = {{6{io_in_369[4]}},io_in_369}; // @[Modules.scala 32:22:@8.4]
  assign _T_56837 = $signed(buffer_1_184) + $signed(buffer_0_185); // @[Modules.scala 65:57:@3543.4]
  assign _T_56838 = _T_56837[10:0]; // @[Modules.scala 65:57:@3544.4]
  assign buffer_1_484 = $signed(_T_56838); // @[Modules.scala 65:57:@3545.4]
  assign _T_56843 = $signed(buffer_0_188) + $signed(11'sh0); // @[Modules.scala 65:57:@3551.4]
  assign _T_56844 = _T_56843[10:0]; // @[Modules.scala 65:57:@3552.4]
  assign buffer_1_486 = $signed(_T_56844); // @[Modules.scala 65:57:@3553.4]
  assign _T_56852 = $signed(buffer_0_194) + $signed(11'sh0); // @[Modules.scala 65:57:@3563.4]
  assign _T_56853 = _T_56852[10:0]; // @[Modules.scala 65:57:@3564.4]
  assign buffer_1_489 = $signed(_T_56853); // @[Modules.scala 65:57:@3565.4]
  assign buffer_1_196 = {{6{_T_56251[4]}},_T_56251}; // @[Modules.scala 32:22:@8.4]
  assign _T_56855 = $signed(buffer_1_196) + $signed(11'sh0); // @[Modules.scala 65:57:@3567.4]
  assign _T_56856 = _T_56855[10:0]; // @[Modules.scala 65:57:@3568.4]
  assign buffer_1_490 = $signed(_T_56856); // @[Modules.scala 65:57:@3569.4]
  assign buffer_1_198 = {{6{io_in_397[4]}},io_in_397}; // @[Modules.scala 32:22:@8.4]
  assign _T_56858 = $signed(buffer_1_198) + $signed(buffer_0_199); // @[Modules.scala 65:57:@3571.4]
  assign _T_56859 = _T_56858[10:0]; // @[Modules.scala 65:57:@3572.4]
  assign buffer_1_491 = $signed(_T_56859); // @[Modules.scala 65:57:@3573.4]
  assign buffer_1_202 = {{6{io_in_404[4]}},io_in_404}; // @[Modules.scala 32:22:@8.4]
  assign _T_56864 = $signed(buffer_1_202) + $signed(11'sh0); // @[Modules.scala 65:57:@3579.4]
  assign _T_56865 = _T_56864[10:0]; // @[Modules.scala 65:57:@3580.4]
  assign buffer_1_493 = $signed(_T_56865); // @[Modules.scala 65:57:@3581.4]
  assign buffer_1_204 = {{6{io_in_408[4]}},io_in_408}; // @[Modules.scala 32:22:@8.4]
  assign _T_56867 = $signed(buffer_1_204) + $signed(11'sh0); // @[Modules.scala 65:57:@3583.4]
  assign _T_56868 = _T_56867[10:0]; // @[Modules.scala 65:57:@3584.4]
  assign buffer_1_494 = $signed(_T_56868); // @[Modules.scala 65:57:@3585.4]
  assign _T_56873 = $signed(buffer_0_208) + $signed(11'sh0); // @[Modules.scala 65:57:@3591.4]
  assign _T_56874 = _T_56873[10:0]; // @[Modules.scala 65:57:@3592.4]
  assign buffer_1_496 = $signed(_T_56874); // @[Modules.scala 65:57:@3593.4]
  assign buffer_1_211 = {{6{io_in_422[4]}},io_in_422}; // @[Modules.scala 32:22:@8.4]
  assign _T_56876 = $signed(buffer_0_210) + $signed(buffer_1_211); // @[Modules.scala 65:57:@3595.4]
  assign _T_56877 = _T_56876[10:0]; // @[Modules.scala 65:57:@3596.4]
  assign buffer_1_497 = $signed(_T_56877); // @[Modules.scala 65:57:@3597.4]
  assign _T_56879 = $signed(buffer_0_212) + $signed(11'sh0); // @[Modules.scala 65:57:@3599.4]
  assign _T_56880 = _T_56879[10:0]; // @[Modules.scala 65:57:@3600.4]
  assign buffer_1_498 = $signed(_T_56880); // @[Modules.scala 65:57:@3601.4]
  assign buffer_1_219 = {{6{io_in_439[4]}},io_in_439}; // @[Modules.scala 32:22:@8.4]
  assign _T_56888 = $signed(11'sh0) + $signed(buffer_1_219); // @[Modules.scala 65:57:@3611.4]
  assign _T_56889 = _T_56888[10:0]; // @[Modules.scala 65:57:@3612.4]
  assign buffer_1_501 = $signed(_T_56889); // @[Modules.scala 65:57:@3613.4]
  assign buffer_1_220 = {{6{_T_56283[4]}},_T_56283}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_221 = {{6{_T_56286[4]}},_T_56286}; // @[Modules.scala 32:22:@8.4]
  assign _T_56891 = $signed(buffer_1_220) + $signed(buffer_1_221); // @[Modules.scala 65:57:@3615.4]
  assign _T_56892 = _T_56891[10:0]; // @[Modules.scala 65:57:@3616.4]
  assign buffer_1_502 = $signed(_T_56892); // @[Modules.scala 65:57:@3617.4]
  assign buffer_1_222 = {{6{io_in_444[4]}},io_in_444}; // @[Modules.scala 32:22:@8.4]
  assign _T_56894 = $signed(buffer_1_222) + $signed(11'sh0); // @[Modules.scala 65:57:@3619.4]
  assign _T_56895 = _T_56894[10:0]; // @[Modules.scala 65:57:@3620.4]
  assign buffer_1_503 = $signed(_T_56895); // @[Modules.scala 65:57:@3621.4]
  assign buffer_1_224 = {{6{io_in_449[4]}},io_in_449}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_225 = {{6{_T_56290[4]}},_T_56290}; // @[Modules.scala 32:22:@8.4]
  assign _T_56897 = $signed(buffer_1_224) + $signed(buffer_1_225); // @[Modules.scala 65:57:@3623.4]
  assign _T_56898 = _T_56897[10:0]; // @[Modules.scala 65:57:@3624.4]
  assign buffer_1_504 = $signed(_T_56898); // @[Modules.scala 65:57:@3625.4]
  assign buffer_1_228 = {{6{io_in_457[4]}},io_in_457}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_229 = {{6{io_in_458[4]}},io_in_458}; // @[Modules.scala 32:22:@8.4]
  assign _T_56903 = $signed(buffer_1_228) + $signed(buffer_1_229); // @[Modules.scala 65:57:@3631.4]
  assign _T_56904 = _T_56903[10:0]; // @[Modules.scala 65:57:@3632.4]
  assign buffer_1_506 = $signed(_T_56904); // @[Modules.scala 65:57:@3633.4]
  assign buffer_1_233 = {{6{io_in_467[4]}},io_in_467}; // @[Modules.scala 32:22:@8.4]
  assign _T_56909 = $signed(11'sh0) + $signed(buffer_1_233); // @[Modules.scala 65:57:@3639.4]
  assign _T_56910 = _T_56909[10:0]; // @[Modules.scala 65:57:@3640.4]
  assign buffer_1_508 = $signed(_T_56910); // @[Modules.scala 65:57:@3641.4]
  assign buffer_1_234 = {{6{_T_56298[4]}},_T_56298}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_235 = {{6{_T_56301[4]}},_T_56301}; // @[Modules.scala 32:22:@8.4]
  assign _T_56912 = $signed(buffer_1_234) + $signed(buffer_1_235); // @[Modules.scala 65:57:@3643.4]
  assign _T_56913 = _T_56912[10:0]; // @[Modules.scala 65:57:@3644.4]
  assign buffer_1_509 = $signed(_T_56913); // @[Modules.scala 65:57:@3645.4]
  assign buffer_1_236 = {{6{io_in_472[4]}},io_in_472}; // @[Modules.scala 32:22:@8.4]
  assign _T_56915 = $signed(buffer_1_236) + $signed(11'sh0); // @[Modules.scala 65:57:@3647.4]
  assign _T_56916 = _T_56915[10:0]; // @[Modules.scala 65:57:@3648.4]
  assign buffer_1_510 = $signed(_T_56916); // @[Modules.scala 65:57:@3649.4]
  assign buffer_1_238 = {{6{io_in_477[4]}},io_in_477}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_239 = {{6{_T_56305[4]}},_T_56305}; // @[Modules.scala 32:22:@8.4]
  assign _T_56918 = $signed(buffer_1_238) + $signed(buffer_1_239); // @[Modules.scala 65:57:@3651.4]
  assign _T_56919 = _T_56918[10:0]; // @[Modules.scala 65:57:@3652.4]
  assign buffer_1_511 = $signed(_T_56919); // @[Modules.scala 65:57:@3653.4]
  assign buffer_1_247 = {{6{_T_56317[4]}},_T_56317}; // @[Modules.scala 32:22:@8.4]
  assign _T_56930 = $signed(11'sh0) + $signed(buffer_1_247); // @[Modules.scala 65:57:@3667.4]
  assign _T_56931 = _T_56930[10:0]; // @[Modules.scala 65:57:@3668.4]
  assign buffer_1_515 = $signed(_T_56931); // @[Modules.scala 65:57:@3669.4]
  assign buffer_1_248 = {{6{_T_56320[4]}},_T_56320}; // @[Modules.scala 32:22:@8.4]
  assign _T_56933 = $signed(buffer_1_248) + $signed(buffer_0_249); // @[Modules.scala 65:57:@3671.4]
  assign _T_56934 = _T_56933[10:0]; // @[Modules.scala 65:57:@3672.4]
  assign buffer_1_516 = $signed(_T_56934); // @[Modules.scala 65:57:@3673.4]
  assign buffer_1_252 = {{6{io_in_505[4]}},io_in_505}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_253 = {{6{_T_56328[4]}},_T_56328}; // @[Modules.scala 32:22:@8.4]
  assign _T_56939 = $signed(buffer_1_252) + $signed(buffer_1_253); // @[Modules.scala 65:57:@3679.4]
  assign _T_56940 = _T_56939[10:0]; // @[Modules.scala 65:57:@3680.4]
  assign buffer_1_518 = $signed(_T_56940); // @[Modules.scala 65:57:@3681.4]
  assign buffer_1_254 = {{6{io_in_508[4]}},io_in_508}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_255 = {{6{_T_56331[4]}},_T_56331}; // @[Modules.scala 32:22:@8.4]
  assign _T_56942 = $signed(buffer_1_254) + $signed(buffer_1_255); // @[Modules.scala 65:57:@3683.4]
  assign _T_56943 = _T_56942[10:0]; // @[Modules.scala 65:57:@3684.4]
  assign buffer_1_519 = $signed(_T_56943); // @[Modules.scala 65:57:@3685.4]
  assign _T_56945 = $signed(11'sh0) + $signed(buffer_0_257); // @[Modules.scala 65:57:@3687.4]
  assign _T_56946 = _T_56945[10:0]; // @[Modules.scala 65:57:@3688.4]
  assign buffer_1_520 = $signed(_T_56946); // @[Modules.scala 65:57:@3689.4]
  assign buffer_1_260 = {{6{_T_56340[4]}},_T_56340}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_261 = {{6{_T_56343[4]}},_T_56343}; // @[Modules.scala 32:22:@8.4]
  assign _T_56951 = $signed(buffer_1_260) + $signed(buffer_1_261); // @[Modules.scala 65:57:@3695.4]
  assign _T_56952 = _T_56951[10:0]; // @[Modules.scala 65:57:@3696.4]
  assign buffer_1_522 = $signed(_T_56952); // @[Modules.scala 65:57:@3697.4]
  assign buffer_1_262 = {{6{_T_56346[4]}},_T_56346}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_263 = {{6{io_in_526[4]}},io_in_526}; // @[Modules.scala 32:22:@8.4]
  assign _T_56954 = $signed(buffer_1_262) + $signed(buffer_1_263); // @[Modules.scala 65:57:@3699.4]
  assign _T_56955 = _T_56954[10:0]; // @[Modules.scala 65:57:@3700.4]
  assign buffer_1_523 = $signed(_T_56955); // @[Modules.scala 65:57:@3701.4]
  assign buffer_1_266 = {{6{_T_56351[4]}},_T_56351}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_267 = {{6{_T_56354[4]}},_T_56354}; // @[Modules.scala 32:22:@8.4]
  assign _T_56960 = $signed(buffer_1_266) + $signed(buffer_1_267); // @[Modules.scala 65:57:@3707.4]
  assign _T_56961 = _T_56960[10:0]; // @[Modules.scala 65:57:@3708.4]
  assign buffer_1_525 = $signed(_T_56961); // @[Modules.scala 65:57:@3709.4]
  assign buffer_1_268 = {{6{_T_56357[4]}},_T_56357}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_269 = {{6{_T_56360[4]}},_T_56360}; // @[Modules.scala 32:22:@8.4]
  assign _T_56963 = $signed(buffer_1_268) + $signed(buffer_1_269); // @[Modules.scala 65:57:@3711.4]
  assign _T_56964 = _T_56963[10:0]; // @[Modules.scala 65:57:@3712.4]
  assign buffer_1_526 = $signed(_T_56964); // @[Modules.scala 65:57:@3713.4]
  assign buffer_1_270 = {{6{_T_56363[4]}},_T_56363}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_271 = {{6{_T_56366[4]}},_T_56366}; // @[Modules.scala 32:22:@8.4]
  assign _T_56966 = $signed(buffer_1_270) + $signed(buffer_1_271); // @[Modules.scala 65:57:@3715.4]
  assign _T_56967 = _T_56966[10:0]; // @[Modules.scala 65:57:@3716.4]
  assign buffer_1_527 = $signed(_T_56967); // @[Modules.scala 65:57:@3717.4]
  assign buffer_1_272 = {{6{_T_56369[4]}},_T_56369}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_273 = {{6{io_in_547[4]}},io_in_547}; // @[Modules.scala 32:22:@8.4]
  assign _T_56969 = $signed(buffer_1_272) + $signed(buffer_1_273); // @[Modules.scala 65:57:@3719.4]
  assign _T_56970 = _T_56969[10:0]; // @[Modules.scala 65:57:@3720.4]
  assign buffer_1_528 = $signed(_T_56970); // @[Modules.scala 65:57:@3721.4]
  assign buffer_1_274 = {{6{_T_56372[4]}},_T_56372}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_275 = {{6{_T_56375[4]}},_T_56375}; // @[Modules.scala 32:22:@8.4]
  assign _T_56972 = $signed(buffer_1_274) + $signed(buffer_1_275); // @[Modules.scala 65:57:@3723.4]
  assign _T_56973 = _T_56972[10:0]; // @[Modules.scala 65:57:@3724.4]
  assign buffer_1_529 = $signed(_T_56973); // @[Modules.scala 65:57:@3725.4]
  assign buffer_1_277 = {{6{io_in_554[4]}},io_in_554}; // @[Modules.scala 32:22:@8.4]
  assign _T_56975 = $signed(buffer_0_276) + $signed(buffer_1_277); // @[Modules.scala 65:57:@3727.4]
  assign _T_56976 = _T_56975[10:0]; // @[Modules.scala 65:57:@3728.4]
  assign buffer_1_530 = $signed(_T_56976); // @[Modules.scala 65:57:@3729.4]
  assign buffer_1_280 = {{6{io_in_561[4]}},io_in_561}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_281 = {{6{_T_56380[4]}},_T_56380}; // @[Modules.scala 32:22:@8.4]
  assign _T_56981 = $signed(buffer_1_280) + $signed(buffer_1_281); // @[Modules.scala 65:57:@3735.4]
  assign _T_56982 = _T_56981[10:0]; // @[Modules.scala 65:57:@3736.4]
  assign buffer_1_532 = $signed(_T_56982); // @[Modules.scala 65:57:@3737.4]
  assign buffer_1_282 = {{6{_T_56383[4]}},_T_56383}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_283 = {{6{io_in_566[4]}},io_in_566}; // @[Modules.scala 32:22:@8.4]
  assign _T_56984 = $signed(buffer_1_282) + $signed(buffer_1_283); // @[Modules.scala 65:57:@3739.4]
  assign _T_56985 = _T_56984[10:0]; // @[Modules.scala 65:57:@3740.4]
  assign buffer_1_533 = $signed(_T_56985); // @[Modules.scala 65:57:@3741.4]
  assign buffer_1_284 = {{6{_T_56386[4]}},_T_56386}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_285 = {{6{_T_56389[4]}},_T_56389}; // @[Modules.scala 32:22:@8.4]
  assign _T_56987 = $signed(buffer_1_284) + $signed(buffer_1_285); // @[Modules.scala 65:57:@3743.4]
  assign _T_56988 = _T_56987[10:0]; // @[Modules.scala 65:57:@3744.4]
  assign buffer_1_534 = $signed(_T_56988); // @[Modules.scala 65:57:@3745.4]
  assign buffer_1_286 = {{6{_T_56392[4]}},_T_56392}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_287 = {{6{_T_56395[4]}},_T_56395}; // @[Modules.scala 32:22:@8.4]
  assign _T_56990 = $signed(buffer_1_286) + $signed(buffer_1_287); // @[Modules.scala 65:57:@3747.4]
  assign _T_56991 = _T_56990[10:0]; // @[Modules.scala 65:57:@3748.4]
  assign buffer_1_535 = $signed(_T_56991); // @[Modules.scala 65:57:@3749.4]
  assign buffer_1_288 = {{6{io_in_576[4]}},io_in_576}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_289 = {{6{_T_56398[4]}},_T_56398}; // @[Modules.scala 32:22:@8.4]
  assign _T_56993 = $signed(buffer_1_288) + $signed(buffer_1_289); // @[Modules.scala 65:57:@3751.4]
  assign _T_56994 = _T_56993[10:0]; // @[Modules.scala 65:57:@3752.4]
  assign buffer_1_536 = $signed(_T_56994); // @[Modules.scala 65:57:@3753.4]
  assign buffer_1_291 = {{6{io_in_582[4]}},io_in_582}; // @[Modules.scala 32:22:@8.4]
  assign _T_56996 = $signed(buffer_0_290) + $signed(buffer_1_291); // @[Modules.scala 65:57:@3755.4]
  assign _T_56997 = _T_56996[10:0]; // @[Modules.scala 65:57:@3756.4]
  assign buffer_1_537 = $signed(_T_56997); // @[Modules.scala 65:57:@3757.4]
  assign _T_56999 = $signed(11'sh0) + $signed(buffer_0_293); // @[Modules.scala 65:57:@3759.4]
  assign _T_57000 = _T_56999[10:0]; // @[Modules.scala 65:57:@3760.4]
  assign buffer_1_538 = $signed(_T_57000); // @[Modules.scala 65:57:@3761.4]
  assign buffer_1_295 = {{6{_T_56403[4]}},_T_56403}; // @[Modules.scala 32:22:@8.4]
  assign _T_57002 = $signed(11'sh0) + $signed(buffer_1_295); // @[Modules.scala 65:57:@3763.4]
  assign _T_57003 = _T_57002[10:0]; // @[Modules.scala 65:57:@3764.4]
  assign buffer_1_539 = $signed(_T_57003); // @[Modules.scala 65:57:@3765.4]
  assign buffer_1_296 = {{6{_T_56406[4]}},_T_56406}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_297 = {{6{io_in_594[4]}},io_in_594}; // @[Modules.scala 32:22:@8.4]
  assign _T_57005 = $signed(buffer_1_296) + $signed(buffer_1_297); // @[Modules.scala 65:57:@3767.4]
  assign _T_57006 = _T_57005[10:0]; // @[Modules.scala 65:57:@3768.4]
  assign buffer_1_540 = $signed(_T_57006); // @[Modules.scala 65:57:@3769.4]
  assign buffer_1_298 = {{6{io_in_596[4]}},io_in_596}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_299 = {{6{_T_56409[4]}},_T_56409}; // @[Modules.scala 32:22:@8.4]
  assign _T_57008 = $signed(buffer_1_298) + $signed(buffer_1_299); // @[Modules.scala 65:57:@3771.4]
  assign _T_57009 = _T_57008[10:0]; // @[Modules.scala 65:57:@3772.4]
  assign buffer_1_541 = $signed(_T_57009); // @[Modules.scala 65:57:@3773.4]
  assign buffer_1_301 = {{6{_T_56415[4]}},_T_56415}; // @[Modules.scala 32:22:@8.4]
  assign _T_57011 = $signed(buffer_0_300) + $signed(buffer_1_301); // @[Modules.scala 65:57:@3775.4]
  assign _T_57012 = _T_57011[10:0]; // @[Modules.scala 65:57:@3776.4]
  assign buffer_1_542 = $signed(_T_57012); // @[Modules.scala 65:57:@3777.4]
  assign _T_57020 = $signed(11'sh0) + $signed(buffer_0_307); // @[Modules.scala 65:57:@3787.4]
  assign _T_57021 = _T_57020[10:0]; // @[Modules.scala 65:57:@3788.4]
  assign buffer_1_545 = $signed(_T_57021); // @[Modules.scala 65:57:@3789.4]
  assign _T_57023 = $signed(11'sh0) + $signed(buffer_0_309); // @[Modules.scala 65:57:@3791.4]
  assign _T_57024 = _T_57023[10:0]; // @[Modules.scala 65:57:@3792.4]
  assign buffer_1_546 = $signed(_T_57024); // @[Modules.scala 65:57:@3793.4]
  assign buffer_1_310 = {{6{io_in_620[4]}},io_in_620}; // @[Modules.scala 32:22:@8.4]
  assign _T_57026 = $signed(buffer_1_310) + $signed(11'sh0); // @[Modules.scala 65:57:@3795.4]
  assign _T_57027 = _T_57026[10:0]; // @[Modules.scala 65:57:@3796.4]
  assign buffer_1_547 = $signed(_T_57027); // @[Modules.scala 65:57:@3797.4]
  assign buffer_1_312 = {{6{_T_56432[4]}},_T_56432}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_313 = {{6{_T_56435[4]}},_T_56435}; // @[Modules.scala 32:22:@8.4]
  assign _T_57029 = $signed(buffer_1_312) + $signed(buffer_1_313); // @[Modules.scala 65:57:@3799.4]
  assign _T_57030 = _T_57029[10:0]; // @[Modules.scala 65:57:@3800.4]
  assign buffer_1_548 = $signed(_T_57030); // @[Modules.scala 65:57:@3801.4]
  assign buffer_1_314 = {{6{_T_56438[4]}},_T_56438}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_315 = {{6{_T_56441[4]}},_T_56441}; // @[Modules.scala 32:22:@8.4]
  assign _T_57032 = $signed(buffer_1_314) + $signed(buffer_1_315); // @[Modules.scala 65:57:@3803.4]
  assign _T_57033 = _T_57032[10:0]; // @[Modules.scala 65:57:@3804.4]
  assign buffer_1_549 = $signed(_T_57033); // @[Modules.scala 65:57:@3805.4]
  assign buffer_1_316 = {{6{_T_56444[4]}},_T_56444}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_317 = {{6{io_in_634[4]}},io_in_634}; // @[Modules.scala 32:22:@8.4]
  assign _T_57035 = $signed(buffer_1_316) + $signed(buffer_1_317); // @[Modules.scala 65:57:@3807.4]
  assign _T_57036 = _T_57035[10:0]; // @[Modules.scala 65:57:@3808.4]
  assign buffer_1_550 = $signed(_T_57036); // @[Modules.scala 65:57:@3809.4]
  assign buffer_1_318 = {{6{_T_56447[4]}},_T_56447}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_319 = {{6{io_in_638[4]}},io_in_638}; // @[Modules.scala 32:22:@8.4]
  assign _T_57038 = $signed(buffer_1_318) + $signed(buffer_1_319); // @[Modules.scala 65:57:@3811.4]
  assign _T_57039 = _T_57038[10:0]; // @[Modules.scala 65:57:@3812.4]
  assign buffer_1_551 = $signed(_T_57039); // @[Modules.scala 65:57:@3813.4]
  assign buffer_1_321 = {{6{_T_56451[4]}},_T_56451}; // @[Modules.scala 32:22:@8.4]
  assign _T_57041 = $signed(11'sh0) + $signed(buffer_1_321); // @[Modules.scala 65:57:@3815.4]
  assign _T_57042 = _T_57041[10:0]; // @[Modules.scala 65:57:@3816.4]
  assign buffer_1_552 = $signed(_T_57042); // @[Modules.scala 65:57:@3817.4]
  assign _T_57044 = $signed(11'sh0) + $signed(buffer_0_323); // @[Modules.scala 65:57:@3819.4]
  assign _T_57045 = _T_57044[10:0]; // @[Modules.scala 65:57:@3820.4]
  assign buffer_1_553 = $signed(_T_57045); // @[Modules.scala 65:57:@3821.4]
  assign buffer_1_324 = {{6{_T_56458[4]}},_T_56458}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_325 = {{6{_T_56461[4]}},_T_56461}; // @[Modules.scala 32:22:@8.4]
  assign _T_57047 = $signed(buffer_1_324) + $signed(buffer_1_325); // @[Modules.scala 65:57:@3823.4]
  assign _T_57048 = _T_57047[10:0]; // @[Modules.scala 65:57:@3824.4]
  assign buffer_1_554 = $signed(_T_57048); // @[Modules.scala 65:57:@3825.4]
  assign buffer_1_326 = {{6{_T_56464[4]}},_T_56464}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_327 = {{6{_T_56467[4]}},_T_56467}; // @[Modules.scala 32:22:@8.4]
  assign _T_57050 = $signed(buffer_1_326) + $signed(buffer_1_327); // @[Modules.scala 65:57:@3827.4]
  assign _T_57051 = _T_57050[10:0]; // @[Modules.scala 65:57:@3828.4]
  assign buffer_1_555 = $signed(_T_57051); // @[Modules.scala 65:57:@3829.4]
  assign buffer_1_328 = {{6{_T_56470[4]}},_T_56470}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_329 = {{6{_T_56473[4]}},_T_56473}; // @[Modules.scala 32:22:@8.4]
  assign _T_57053 = $signed(buffer_1_328) + $signed(buffer_1_329); // @[Modules.scala 65:57:@3831.4]
  assign _T_57054 = _T_57053[10:0]; // @[Modules.scala 65:57:@3832.4]
  assign buffer_1_556 = $signed(_T_57054); // @[Modules.scala 65:57:@3833.4]
  assign buffer_1_331 = {{6{_T_56477[4]}},_T_56477}; // @[Modules.scala 32:22:@8.4]
  assign _T_57056 = $signed(11'sh0) + $signed(buffer_1_331); // @[Modules.scala 65:57:@3835.4]
  assign _T_57057 = _T_57056[10:0]; // @[Modules.scala 65:57:@3836.4]
  assign buffer_1_557 = $signed(_T_57057); // @[Modules.scala 65:57:@3837.4]
  assign buffer_1_337 = {{6{_T_56485[4]}},_T_56485}; // @[Modules.scala 32:22:@8.4]
  assign _T_57065 = $signed(11'sh0) + $signed(buffer_1_337); // @[Modules.scala 65:57:@3847.4]
  assign _T_57066 = _T_57065[10:0]; // @[Modules.scala 65:57:@3848.4]
  assign buffer_1_560 = $signed(_T_57066); // @[Modules.scala 65:57:@3849.4]
  assign buffer_1_340 = {{6{io_in_681[4]}},io_in_681}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_341 = {{6{_T_56494[4]}},_T_56494}; // @[Modules.scala 32:22:@8.4]
  assign _T_57071 = $signed(buffer_1_340) + $signed(buffer_1_341); // @[Modules.scala 65:57:@3855.4]
  assign _T_57072 = _T_57071[10:0]; // @[Modules.scala 65:57:@3856.4]
  assign buffer_1_562 = $signed(_T_57072); // @[Modules.scala 65:57:@3857.4]
  assign buffer_1_342 = {{6{_T_56497[4]}},_T_56497}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_343 = {{6{io_in_686[4]}},io_in_686}; // @[Modules.scala 32:22:@8.4]
  assign _T_57074 = $signed(buffer_1_342) + $signed(buffer_1_343); // @[Modules.scala 65:57:@3859.4]
  assign _T_57075 = _T_57074[10:0]; // @[Modules.scala 65:57:@3860.4]
  assign buffer_1_563 = $signed(_T_57075); // @[Modules.scala 65:57:@3861.4]
  assign buffer_1_344 = {{6{io_in_688[4]}},io_in_688}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_345 = {{6{io_in_690[4]}},io_in_690}; // @[Modules.scala 32:22:@8.4]
  assign _T_57077 = $signed(buffer_1_344) + $signed(buffer_1_345); // @[Modules.scala 65:57:@3863.4]
  assign _T_57078 = _T_57077[10:0]; // @[Modules.scala 65:57:@3864.4]
  assign buffer_1_564 = $signed(_T_57078); // @[Modules.scala 65:57:@3865.4]
  assign buffer_1_347 = {{6{io_in_695[4]}},io_in_695}; // @[Modules.scala 32:22:@8.4]
  assign _T_57080 = $signed(11'sh0) + $signed(buffer_1_347); // @[Modules.scala 65:57:@3867.4]
  assign _T_57081 = _T_57080[10:0]; // @[Modules.scala 65:57:@3868.4]
  assign buffer_1_565 = $signed(_T_57081); // @[Modules.scala 65:57:@3869.4]
  assign buffer_1_348 = {{6{io_in_696[4]}},io_in_696}; // @[Modules.scala 32:22:@8.4]
  assign _T_57083 = $signed(buffer_1_348) + $signed(11'sh0); // @[Modules.scala 65:57:@3871.4]
  assign _T_57084 = _T_57083[10:0]; // @[Modules.scala 65:57:@3872.4]
  assign buffer_1_566 = $signed(_T_57084); // @[Modules.scala 65:57:@3873.4]
  assign buffer_1_350 = {{6{_T_56502[4]}},_T_56502}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_351 = {{6{_T_56505[4]}},_T_56505}; // @[Modules.scala 32:22:@8.4]
  assign _T_57086 = $signed(buffer_1_350) + $signed(buffer_1_351); // @[Modules.scala 65:57:@3875.4]
  assign _T_57087 = _T_57086[10:0]; // @[Modules.scala 65:57:@3876.4]
  assign buffer_1_567 = $signed(_T_57087); // @[Modules.scala 65:57:@3877.4]
  assign buffer_1_355 = {{6{io_in_711[4]}},io_in_711}; // @[Modules.scala 32:22:@8.4]
  assign _T_57092 = $signed(11'sh0) + $signed(buffer_1_355); // @[Modules.scala 65:57:@3883.4]
  assign _T_57093 = _T_57092[10:0]; // @[Modules.scala 65:57:@3884.4]
  assign buffer_1_569 = $signed(_T_57093); // @[Modules.scala 65:57:@3885.4]
  assign buffer_1_357 = {{6{io_in_715[4]}},io_in_715}; // @[Modules.scala 32:22:@8.4]
  assign _T_57095 = $signed(11'sh0) + $signed(buffer_1_357); // @[Modules.scala 65:57:@3887.4]
  assign _T_57096 = _T_57095[10:0]; // @[Modules.scala 65:57:@3888.4]
  assign buffer_1_570 = $signed(_T_57096); // @[Modules.scala 65:57:@3889.4]
  assign buffer_1_358 = {{6{io_in_716[4]}},io_in_716}; // @[Modules.scala 32:22:@8.4]
  assign _T_57098 = $signed(buffer_1_358) + $signed(11'sh0); // @[Modules.scala 65:57:@3891.4]
  assign _T_57099 = _T_57098[10:0]; // @[Modules.scala 65:57:@3892.4]
  assign buffer_1_571 = $signed(_T_57099); // @[Modules.scala 65:57:@3893.4]
  assign _T_57101 = $signed(11'sh0) + $signed(buffer_0_361); // @[Modules.scala 65:57:@3895.4]
  assign _T_57102 = _T_57101[10:0]; // @[Modules.scala 65:57:@3896.4]
  assign buffer_1_572 = $signed(_T_57102); // @[Modules.scala 65:57:@3897.4]
  assign buffer_1_362 = {{6{_T_56521[4]}},_T_56521}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_363 = {{6{io_in_726[4]}},io_in_726}; // @[Modules.scala 32:22:@8.4]
  assign _T_57104 = $signed(buffer_1_362) + $signed(buffer_1_363); // @[Modules.scala 65:57:@3899.4]
  assign _T_57105 = _T_57104[10:0]; // @[Modules.scala 65:57:@3900.4]
  assign buffer_1_573 = $signed(_T_57105); // @[Modules.scala 65:57:@3901.4]
  assign buffer_1_378 = {{6{io_in_756[4]}},io_in_756}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_379 = {{6{_T_56543[4]}},_T_56543}; // @[Modules.scala 32:22:@8.4]
  assign _T_57128 = $signed(buffer_1_378) + $signed(buffer_1_379); // @[Modules.scala 65:57:@3931.4]
  assign _T_57129 = _T_57128[10:0]; // @[Modules.scala 65:57:@3932.4]
  assign buffer_1_581 = $signed(_T_57129); // @[Modules.scala 65:57:@3933.4]
  assign buffer_1_380 = {{6{_T_56546[4]}},_T_56546}; // @[Modules.scala 32:22:@8.4]
  assign buffer_1_381 = {{6{_T_56549[4]}},_T_56549}; // @[Modules.scala 32:22:@8.4]
  assign _T_57131 = $signed(buffer_1_380) + $signed(buffer_1_381); // @[Modules.scala 65:57:@3935.4]
  assign _T_57132 = _T_57131[10:0]; // @[Modules.scala 65:57:@3936.4]
  assign buffer_1_582 = $signed(_T_57132); // @[Modules.scala 65:57:@3937.4]
  assign buffer_1_383 = {{6{_T_56553[4]}},_T_56553}; // @[Modules.scala 32:22:@8.4]
  assign _T_57134 = $signed(11'sh0) + $signed(buffer_1_383); // @[Modules.scala 65:57:@3939.4]
  assign _T_57135 = _T_57134[10:0]; // @[Modules.scala 65:57:@3940.4]
  assign buffer_1_583 = $signed(_T_57135); // @[Modules.scala 65:57:@3941.4]
  assign buffer_1_390 = {{6{io_in_780[4]}},io_in_780}; // @[Modules.scala 32:22:@8.4]
  assign _T_57146 = $signed(buffer_1_390) + $signed(11'sh0); // @[Modules.scala 65:57:@3955.4]
  assign _T_57147 = _T_57146[10:0]; // @[Modules.scala 65:57:@3956.4]
  assign buffer_1_587 = $signed(_T_57147); // @[Modules.scala 65:57:@3957.4]
  assign _T_57149 = $signed(buffer_0_395) + $signed(buffer_1_393); // @[Modules.scala 68:83:@3959.4]
  assign _T_57150 = _T_57149[10:0]; // @[Modules.scala 68:83:@3960.4]
  assign buffer_1_588 = $signed(_T_57150); // @[Modules.scala 68:83:@3961.4]
  assign _T_57152 = $signed(buffer_1_394) + $signed(buffer_1_395); // @[Modules.scala 68:83:@3963.4]
  assign _T_57153 = _T_57152[10:0]; // @[Modules.scala 68:83:@3964.4]
  assign buffer_1_589 = $signed(_T_57153); // @[Modules.scala 68:83:@3965.4]
  assign _T_57155 = $signed(buffer_1_396) + $signed(buffer_1_397); // @[Modules.scala 68:83:@3967.4]
  assign _T_57156 = _T_57155[10:0]; // @[Modules.scala 68:83:@3968.4]
  assign buffer_1_590 = $signed(_T_57156); // @[Modules.scala 68:83:@3969.4]
  assign _T_57158 = $signed(buffer_1_398) + $signed(buffer_1_399); // @[Modules.scala 68:83:@3971.4]
  assign _T_57159 = _T_57158[10:0]; // @[Modules.scala 68:83:@3972.4]
  assign buffer_1_591 = $signed(_T_57159); // @[Modules.scala 68:83:@3973.4]
  assign _T_57161 = $signed(buffer_1_400) + $signed(buffer_1_401); // @[Modules.scala 68:83:@3975.4]
  assign _T_57162 = _T_57161[10:0]; // @[Modules.scala 68:83:@3976.4]
  assign buffer_1_592 = $signed(_T_57162); // @[Modules.scala 68:83:@3977.4]
  assign _T_57164 = $signed(buffer_1_402) + $signed(buffer_1_403); // @[Modules.scala 68:83:@3979.4]
  assign _T_57165 = _T_57164[10:0]; // @[Modules.scala 68:83:@3980.4]
  assign buffer_1_593 = $signed(_T_57165); // @[Modules.scala 68:83:@3981.4]
  assign _T_57167 = $signed(buffer_1_404) + $signed(buffer_1_405); // @[Modules.scala 68:83:@3983.4]
  assign _T_57168 = _T_57167[10:0]; // @[Modules.scala 68:83:@3984.4]
  assign buffer_1_594 = $signed(_T_57168); // @[Modules.scala 68:83:@3985.4]
  assign _T_57170 = $signed(buffer_1_406) + $signed(buffer_1_407); // @[Modules.scala 68:83:@3987.4]
  assign _T_57171 = _T_57170[10:0]; // @[Modules.scala 68:83:@3988.4]
  assign buffer_1_595 = $signed(_T_57171); // @[Modules.scala 68:83:@3989.4]
  assign _T_57173 = $signed(buffer_1_408) + $signed(buffer_1_409); // @[Modules.scala 68:83:@3991.4]
  assign _T_57174 = _T_57173[10:0]; // @[Modules.scala 68:83:@3992.4]
  assign buffer_1_596 = $signed(_T_57174); // @[Modules.scala 68:83:@3993.4]
  assign _T_57176 = $signed(buffer_1_410) + $signed(buffer_1_411); // @[Modules.scala 68:83:@3995.4]
  assign _T_57177 = _T_57176[10:0]; // @[Modules.scala 68:83:@3996.4]
  assign buffer_1_597 = $signed(_T_57177); // @[Modules.scala 68:83:@3997.4]
  assign _T_57179 = $signed(buffer_1_412) + $signed(buffer_1_413); // @[Modules.scala 68:83:@3999.4]
  assign _T_57180 = _T_57179[10:0]; // @[Modules.scala 68:83:@4000.4]
  assign buffer_1_598 = $signed(_T_57180); // @[Modules.scala 68:83:@4001.4]
  assign _T_57182 = $signed(buffer_0_414) + $signed(buffer_1_415); // @[Modules.scala 68:83:@4003.4]
  assign _T_57183 = _T_57182[10:0]; // @[Modules.scala 68:83:@4004.4]
  assign buffer_1_599 = $signed(_T_57183); // @[Modules.scala 68:83:@4005.4]
  assign _T_57185 = $signed(buffer_1_416) + $signed(buffer_0_417); // @[Modules.scala 68:83:@4007.4]
  assign _T_57186 = _T_57185[10:0]; // @[Modules.scala 68:83:@4008.4]
  assign buffer_1_600 = $signed(_T_57186); // @[Modules.scala 68:83:@4009.4]
  assign _T_57188 = $signed(buffer_0_418) + $signed(buffer_1_419); // @[Modules.scala 68:83:@4011.4]
  assign _T_57189 = _T_57188[10:0]; // @[Modules.scala 68:83:@4012.4]
  assign buffer_1_601 = $signed(_T_57189); // @[Modules.scala 68:83:@4013.4]
  assign _T_57191 = $signed(buffer_1_420) + $signed(buffer_1_421); // @[Modules.scala 68:83:@4015.4]
  assign _T_57192 = _T_57191[10:0]; // @[Modules.scala 68:83:@4016.4]
  assign buffer_1_602 = $signed(_T_57192); // @[Modules.scala 68:83:@4017.4]
  assign _T_57194 = $signed(buffer_0_395) + $signed(buffer_1_423); // @[Modules.scala 68:83:@4019.4]
  assign _T_57195 = _T_57194[10:0]; // @[Modules.scala 68:83:@4020.4]
  assign buffer_1_603 = $signed(_T_57195); // @[Modules.scala 68:83:@4021.4]
  assign _T_57197 = $signed(buffer_1_424) + $signed(buffer_1_425); // @[Modules.scala 68:83:@4023.4]
  assign _T_57198 = _T_57197[10:0]; // @[Modules.scala 68:83:@4024.4]
  assign buffer_1_604 = $signed(_T_57198); // @[Modules.scala 68:83:@4025.4]
  assign _T_57200 = $signed(buffer_1_426) + $signed(buffer_1_427); // @[Modules.scala 68:83:@4027.4]
  assign _T_57201 = _T_57200[10:0]; // @[Modules.scala 68:83:@4028.4]
  assign buffer_1_605 = $signed(_T_57201); // @[Modules.scala 68:83:@4029.4]
  assign _T_57203 = $signed(buffer_0_395) + $signed(buffer_1_429); // @[Modules.scala 68:83:@4031.4]
  assign _T_57204 = _T_57203[10:0]; // @[Modules.scala 68:83:@4032.4]
  assign buffer_1_606 = $signed(_T_57204); // @[Modules.scala 68:83:@4033.4]
  assign _T_57206 = $signed(buffer_0_395) + $signed(buffer_1_431); // @[Modules.scala 68:83:@4035.4]
  assign _T_57207 = _T_57206[10:0]; // @[Modules.scala 68:83:@4036.4]
  assign buffer_1_607 = $signed(_T_57207); // @[Modules.scala 68:83:@4037.4]
  assign _T_57209 = $signed(buffer_1_432) + $signed(buffer_1_433); // @[Modules.scala 68:83:@4039.4]
  assign _T_57210 = _T_57209[10:0]; // @[Modules.scala 68:83:@4040.4]
  assign buffer_1_608 = $signed(_T_57210); // @[Modules.scala 68:83:@4041.4]
  assign _T_57212 = $signed(buffer_1_434) + $signed(buffer_1_435); // @[Modules.scala 68:83:@4043.4]
  assign _T_57213 = _T_57212[10:0]; // @[Modules.scala 68:83:@4044.4]
  assign buffer_1_609 = $signed(_T_57213); // @[Modules.scala 68:83:@4045.4]
  assign _T_57215 = $signed(buffer_1_436) + $signed(buffer_1_437); // @[Modules.scala 68:83:@4047.4]
  assign _T_57216 = _T_57215[10:0]; // @[Modules.scala 68:83:@4048.4]
  assign buffer_1_610 = $signed(_T_57216); // @[Modules.scala 68:83:@4049.4]
  assign _T_57218 = $signed(buffer_0_438) + $signed(buffer_1_439); // @[Modules.scala 68:83:@4051.4]
  assign _T_57219 = _T_57218[10:0]; // @[Modules.scala 68:83:@4052.4]
  assign buffer_1_611 = $signed(_T_57219); // @[Modules.scala 68:83:@4053.4]
  assign _T_57221 = $signed(buffer_1_440) + $signed(buffer_1_441); // @[Modules.scala 68:83:@4055.4]
  assign _T_57222 = _T_57221[10:0]; // @[Modules.scala 68:83:@4056.4]
  assign buffer_1_612 = $signed(_T_57222); // @[Modules.scala 68:83:@4057.4]
  assign _T_57224 = $signed(buffer_1_442) + $signed(buffer_1_443); // @[Modules.scala 68:83:@4059.4]
  assign _T_57225 = _T_57224[10:0]; // @[Modules.scala 68:83:@4060.4]
  assign buffer_1_613 = $signed(_T_57225); // @[Modules.scala 68:83:@4061.4]
  assign _T_57227 = $signed(buffer_1_444) + $signed(buffer_1_445); // @[Modules.scala 68:83:@4063.4]
  assign _T_57228 = _T_57227[10:0]; // @[Modules.scala 68:83:@4064.4]
  assign buffer_1_614 = $signed(_T_57228); // @[Modules.scala 68:83:@4065.4]
  assign _T_57230 = $signed(buffer_1_446) + $signed(buffer_1_447); // @[Modules.scala 68:83:@4067.4]
  assign _T_57231 = _T_57230[10:0]; // @[Modules.scala 68:83:@4068.4]
  assign buffer_1_615 = $signed(_T_57231); // @[Modules.scala 68:83:@4069.4]
  assign _T_57233 = $signed(buffer_1_448) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4071.4]
  assign _T_57234 = _T_57233[10:0]; // @[Modules.scala 68:83:@4072.4]
  assign buffer_1_616 = $signed(_T_57234); // @[Modules.scala 68:83:@4073.4]
  assign _T_57239 = $signed(buffer_1_452) + $signed(buffer_1_453); // @[Modules.scala 68:83:@4079.4]
  assign _T_57240 = _T_57239[10:0]; // @[Modules.scala 68:83:@4080.4]
  assign buffer_1_618 = $signed(_T_57240); // @[Modules.scala 68:83:@4081.4]
  assign _T_57242 = $signed(buffer_1_454) + $signed(buffer_1_455); // @[Modules.scala 68:83:@4083.4]
  assign _T_57243 = _T_57242[10:0]; // @[Modules.scala 68:83:@4084.4]
  assign buffer_1_619 = $signed(_T_57243); // @[Modules.scala 68:83:@4085.4]
  assign _T_57245 = $signed(buffer_0_395) + $signed(buffer_1_457); // @[Modules.scala 68:83:@4087.4]
  assign _T_57246 = _T_57245[10:0]; // @[Modules.scala 68:83:@4088.4]
  assign buffer_1_620 = $signed(_T_57246); // @[Modules.scala 68:83:@4089.4]
  assign _T_57248 = $signed(buffer_1_458) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4091.4]
  assign _T_57249 = _T_57248[10:0]; // @[Modules.scala 68:83:@4092.4]
  assign buffer_1_621 = $signed(_T_57249); // @[Modules.scala 68:83:@4093.4]
  assign _T_57251 = $signed(buffer_1_460) + $signed(buffer_1_461); // @[Modules.scala 68:83:@4095.4]
  assign _T_57252 = _T_57251[10:0]; // @[Modules.scala 68:83:@4096.4]
  assign buffer_1_622 = $signed(_T_57252); // @[Modules.scala 68:83:@4097.4]
  assign _T_57254 = $signed(buffer_1_462) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4099.4]
  assign _T_57255 = _T_57254[10:0]; // @[Modules.scala 68:83:@4100.4]
  assign buffer_1_623 = $signed(_T_57255); // @[Modules.scala 68:83:@4101.4]
  assign _T_57257 = $signed(buffer_0_464) + $signed(buffer_1_465); // @[Modules.scala 68:83:@4103.4]
  assign _T_57258 = _T_57257[10:0]; // @[Modules.scala 68:83:@4104.4]
  assign buffer_1_624 = $signed(_T_57258); // @[Modules.scala 68:83:@4105.4]
  assign _T_57260 = $signed(buffer_0_395) + $signed(buffer_1_467); // @[Modules.scala 68:83:@4107.4]
  assign _T_57261 = _T_57260[10:0]; // @[Modules.scala 68:83:@4108.4]
  assign buffer_1_625 = $signed(_T_57261); // @[Modules.scala 68:83:@4109.4]
  assign _T_57263 = $signed(buffer_1_468) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4111.4]
  assign _T_57264 = _T_57263[10:0]; // @[Modules.scala 68:83:@4112.4]
  assign buffer_1_626 = $signed(_T_57264); // @[Modules.scala 68:83:@4113.4]
  assign _T_57266 = $signed(buffer_1_470) + $signed(buffer_1_471); // @[Modules.scala 68:83:@4115.4]
  assign _T_57267 = _T_57266[10:0]; // @[Modules.scala 68:83:@4116.4]
  assign buffer_1_627 = $signed(_T_57267); // @[Modules.scala 68:83:@4117.4]
  assign _T_57269 = $signed(buffer_1_472) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4119.4]
  assign _T_57270 = _T_57269[10:0]; // @[Modules.scala 68:83:@4120.4]
  assign buffer_1_628 = $signed(_T_57270); // @[Modules.scala 68:83:@4121.4]
  assign _T_57272 = $signed(buffer_1_474) + $signed(buffer_1_475); // @[Modules.scala 68:83:@4123.4]
  assign _T_57273 = _T_57272[10:0]; // @[Modules.scala 68:83:@4124.4]
  assign buffer_1_629 = $signed(_T_57273); // @[Modules.scala 68:83:@4125.4]
  assign _T_57278 = $signed(buffer_0_478) + $signed(buffer_1_479); // @[Modules.scala 68:83:@4131.4]
  assign _T_57279 = _T_57278[10:0]; // @[Modules.scala 68:83:@4132.4]
  assign buffer_1_631 = $signed(_T_57279); // @[Modules.scala 68:83:@4133.4]
  assign _T_57281 = $signed(buffer_0_395) + $signed(buffer_1_481); // @[Modules.scala 68:83:@4135.4]
  assign _T_57282 = _T_57281[10:0]; // @[Modules.scala 68:83:@4136.4]
  assign buffer_1_632 = $signed(_T_57282); // @[Modules.scala 68:83:@4137.4]
  assign _T_57284 = $signed(buffer_1_482) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4139.4]
  assign _T_57285 = _T_57284[10:0]; // @[Modules.scala 68:83:@4140.4]
  assign buffer_1_633 = $signed(_T_57285); // @[Modules.scala 68:83:@4141.4]
  assign _T_57287 = $signed(buffer_1_484) + $signed(buffer_0_485); // @[Modules.scala 68:83:@4143.4]
  assign _T_57288 = _T_57287[10:0]; // @[Modules.scala 68:83:@4144.4]
  assign buffer_1_634 = $signed(_T_57288); // @[Modules.scala 68:83:@4145.4]
  assign _T_57290 = $signed(buffer_1_486) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4147.4]
  assign _T_57291 = _T_57290[10:0]; // @[Modules.scala 68:83:@4148.4]
  assign buffer_1_635 = $signed(_T_57291); // @[Modules.scala 68:83:@4149.4]
  assign _T_57293 = $signed(buffer_0_488) + $signed(buffer_1_489); // @[Modules.scala 68:83:@4151.4]
  assign _T_57294 = _T_57293[10:0]; // @[Modules.scala 68:83:@4152.4]
  assign buffer_1_636 = $signed(_T_57294); // @[Modules.scala 68:83:@4153.4]
  assign _T_57296 = $signed(buffer_1_490) + $signed(buffer_1_491); // @[Modules.scala 68:83:@4155.4]
  assign _T_57297 = _T_57296[10:0]; // @[Modules.scala 68:83:@4156.4]
  assign buffer_1_637 = $signed(_T_57297); // @[Modules.scala 68:83:@4157.4]
  assign _T_57299 = $signed(buffer_0_492) + $signed(buffer_1_493); // @[Modules.scala 68:83:@4159.4]
  assign _T_57300 = _T_57299[10:0]; // @[Modules.scala 68:83:@4160.4]
  assign buffer_1_638 = $signed(_T_57300); // @[Modules.scala 68:83:@4161.4]
  assign _T_57302 = $signed(buffer_1_494) + $signed(buffer_0_495); // @[Modules.scala 68:83:@4163.4]
  assign _T_57303 = _T_57302[10:0]; // @[Modules.scala 68:83:@4164.4]
  assign buffer_1_639 = $signed(_T_57303); // @[Modules.scala 68:83:@4165.4]
  assign _T_57305 = $signed(buffer_1_496) + $signed(buffer_1_497); // @[Modules.scala 68:83:@4167.4]
  assign _T_57306 = _T_57305[10:0]; // @[Modules.scala 68:83:@4168.4]
  assign buffer_1_640 = $signed(_T_57306); // @[Modules.scala 68:83:@4169.4]
  assign _T_57308 = $signed(buffer_1_498) + $signed(buffer_0_499); // @[Modules.scala 68:83:@4171.4]
  assign _T_57309 = _T_57308[10:0]; // @[Modules.scala 68:83:@4172.4]
  assign buffer_1_641 = $signed(_T_57309); // @[Modules.scala 68:83:@4173.4]
  assign _T_57311 = $signed(buffer_0_395) + $signed(buffer_1_501); // @[Modules.scala 68:83:@4175.4]
  assign _T_57312 = _T_57311[10:0]; // @[Modules.scala 68:83:@4176.4]
  assign buffer_1_642 = $signed(_T_57312); // @[Modules.scala 68:83:@4177.4]
  assign _T_57314 = $signed(buffer_1_502) + $signed(buffer_1_503); // @[Modules.scala 68:83:@4179.4]
  assign _T_57315 = _T_57314[10:0]; // @[Modules.scala 68:83:@4180.4]
  assign buffer_1_643 = $signed(_T_57315); // @[Modules.scala 68:83:@4181.4]
  assign _T_57317 = $signed(buffer_1_504) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4183.4]
  assign _T_57318 = _T_57317[10:0]; // @[Modules.scala 68:83:@4184.4]
  assign buffer_1_644 = $signed(_T_57318); // @[Modules.scala 68:83:@4185.4]
  assign _T_57320 = $signed(buffer_1_506) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4187.4]
  assign _T_57321 = _T_57320[10:0]; // @[Modules.scala 68:83:@4188.4]
  assign buffer_1_645 = $signed(_T_57321); // @[Modules.scala 68:83:@4189.4]
  assign _T_57323 = $signed(buffer_1_508) + $signed(buffer_1_509); // @[Modules.scala 68:83:@4191.4]
  assign _T_57324 = _T_57323[10:0]; // @[Modules.scala 68:83:@4192.4]
  assign buffer_1_646 = $signed(_T_57324); // @[Modules.scala 68:83:@4193.4]
  assign _T_57326 = $signed(buffer_1_510) + $signed(buffer_1_511); // @[Modules.scala 68:83:@4195.4]
  assign _T_57327 = _T_57326[10:0]; // @[Modules.scala 68:83:@4196.4]
  assign buffer_1_647 = $signed(_T_57327); // @[Modules.scala 68:83:@4197.4]
  assign _T_57329 = $signed(buffer_0_512) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4199.4]
  assign _T_57330 = _T_57329[10:0]; // @[Modules.scala 68:83:@4200.4]
  assign buffer_1_648 = $signed(_T_57330); // @[Modules.scala 68:83:@4201.4]
  assign _T_57332 = $signed(buffer_0_395) + $signed(buffer_1_515); // @[Modules.scala 68:83:@4203.4]
  assign _T_57333 = _T_57332[10:0]; // @[Modules.scala 68:83:@4204.4]
  assign buffer_1_649 = $signed(_T_57333); // @[Modules.scala 68:83:@4205.4]
  assign _T_57335 = $signed(buffer_1_516) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4207.4]
  assign _T_57336 = _T_57335[10:0]; // @[Modules.scala 68:83:@4208.4]
  assign buffer_1_650 = $signed(_T_57336); // @[Modules.scala 68:83:@4209.4]
  assign _T_57338 = $signed(buffer_1_518) + $signed(buffer_1_519); // @[Modules.scala 68:83:@4211.4]
  assign _T_57339 = _T_57338[10:0]; // @[Modules.scala 68:83:@4212.4]
  assign buffer_1_651 = $signed(_T_57339); // @[Modules.scala 68:83:@4213.4]
  assign _T_57341 = $signed(buffer_1_520) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4215.4]
  assign _T_57342 = _T_57341[10:0]; // @[Modules.scala 68:83:@4216.4]
  assign buffer_1_652 = $signed(_T_57342); // @[Modules.scala 68:83:@4217.4]
  assign _T_57344 = $signed(buffer_1_522) + $signed(buffer_1_523); // @[Modules.scala 68:83:@4219.4]
  assign _T_57345 = _T_57344[10:0]; // @[Modules.scala 68:83:@4220.4]
  assign buffer_1_653 = $signed(_T_57345); // @[Modules.scala 68:83:@4221.4]
  assign _T_57347 = $signed(buffer_0_395) + $signed(buffer_1_525); // @[Modules.scala 68:83:@4223.4]
  assign _T_57348 = _T_57347[10:0]; // @[Modules.scala 68:83:@4224.4]
  assign buffer_1_654 = $signed(_T_57348); // @[Modules.scala 68:83:@4225.4]
  assign _T_57350 = $signed(buffer_1_526) + $signed(buffer_1_527); // @[Modules.scala 68:83:@4227.4]
  assign _T_57351 = _T_57350[10:0]; // @[Modules.scala 68:83:@4228.4]
  assign buffer_1_655 = $signed(_T_57351); // @[Modules.scala 68:83:@4229.4]
  assign _T_57353 = $signed(buffer_1_528) + $signed(buffer_1_529); // @[Modules.scala 68:83:@4231.4]
  assign _T_57354 = _T_57353[10:0]; // @[Modules.scala 68:83:@4232.4]
  assign buffer_1_656 = $signed(_T_57354); // @[Modules.scala 68:83:@4233.4]
  assign _T_57356 = $signed(buffer_1_530) + $signed(buffer_0_395); // @[Modules.scala 68:83:@4235.4]
  assign _T_57357 = _T_57356[10:0]; // @[Modules.scala 68:83:@4236.4]
  assign buffer_1_657 = $signed(_T_57357); // @[Modules.scala 68:83:@4237.4]
  assign _T_57359 = $signed(buffer_1_532) + $signed(buffer_1_533); // @[Modules.scala 68:83:@4239.4]
  assign _T_57360 = _T_57359[10:0]; // @[Modules.scala 68:83:@4240.4]
  assign buffer_1_658 = $signed(_T_57360); // @[Modules.scala 68:83:@4241.4]
  assign _T_57362 = $signed(buffer_1_534) + $signed(buffer_1_535); // @[Modules.scala 68:83:@4243.4]
  assign _T_57363 = _T_57362[10:0]; // @[Modules.scala 68:83:@4244.4]
  assign buffer_1_659 = $signed(_T_57363); // @[Modules.scala 68:83:@4245.4]
  assign _T_57365 = $signed(buffer_1_536) + $signed(buffer_1_537); // @[Modules.scala 68:83:@4247.4]
  assign _T_57366 = _T_57365[10:0]; // @[Modules.scala 68:83:@4248.4]
  assign buffer_1_660 = $signed(_T_57366); // @[Modules.scala 68:83:@4249.4]
  assign _T_57368 = $signed(buffer_1_538) + $signed(buffer_1_539); // @[Modules.scala 68:83:@4251.4]
  assign _T_57369 = _T_57368[10:0]; // @[Modules.scala 68:83:@4252.4]
  assign buffer_1_661 = $signed(_T_57369); // @[Modules.scala 68:83:@4253.4]
  assign _T_57371 = $signed(buffer_1_540) + $signed(buffer_1_541); // @[Modules.scala 68:83:@4255.4]
  assign _T_57372 = _T_57371[10:0]; // @[Modules.scala 68:83:@4256.4]
  assign buffer_1_662 = $signed(_T_57372); // @[Modules.scala 68:83:@4257.4]
  assign _T_57374 = $signed(buffer_1_542) + $signed(buffer_0_543); // @[Modules.scala 68:83:@4259.4]
  assign _T_57375 = _T_57374[10:0]; // @[Modules.scala 68:83:@4260.4]
  assign buffer_1_663 = $signed(_T_57375); // @[Modules.scala 68:83:@4261.4]
  assign _T_57377 = $signed(buffer_0_395) + $signed(buffer_1_545); // @[Modules.scala 68:83:@4263.4]
  assign _T_57378 = _T_57377[10:0]; // @[Modules.scala 68:83:@4264.4]
  assign buffer_1_664 = $signed(_T_57378); // @[Modules.scala 68:83:@4265.4]
  assign _T_57380 = $signed(buffer_1_546) + $signed(buffer_1_547); // @[Modules.scala 68:83:@4267.4]
  assign _T_57381 = _T_57380[10:0]; // @[Modules.scala 68:83:@4268.4]
  assign buffer_1_665 = $signed(_T_57381); // @[Modules.scala 68:83:@4269.4]
  assign _T_57383 = $signed(buffer_1_548) + $signed(buffer_1_549); // @[Modules.scala 68:83:@4271.4]
  assign _T_57384 = _T_57383[10:0]; // @[Modules.scala 68:83:@4272.4]
  assign buffer_1_666 = $signed(_T_57384); // @[Modules.scala 68:83:@4273.4]
  assign _T_57386 = $signed(buffer_1_550) + $signed(buffer_1_551); // @[Modules.scala 68:83:@4275.4]
  assign _T_57387 = _T_57386[10:0]; // @[Modules.scala 68:83:@4276.4]
  assign buffer_1_667 = $signed(_T_57387); // @[Modules.scala 68:83:@4277.4]
  assign _T_57389 = $signed(buffer_1_552) + $signed(buffer_1_553); // @[Modules.scala 68:83:@4279.4]
  assign _T_57390 = _T_57389[10:0]; // @[Modules.scala 68:83:@4280.4]
  assign buffer_1_668 = $signed(_T_57390); // @[Modules.scala 68:83:@4281.4]
  assign _T_57392 = $signed(buffer_1_554) + $signed(buffer_1_555); // @[Modules.scala 68:83:@4283.4]
  assign _T_57393 = _T_57392[10:0]; // @[Modules.scala 68:83:@4284.4]
  assign buffer_1_669 = $signed(_T_57393); // @[Modules.scala 68:83:@4285.4]
  assign _T_57395 = $signed(buffer_1_556) + $signed(buffer_1_557); // @[Modules.scala 68:83:@4287.4]
  assign _T_57396 = _T_57395[10:0]; // @[Modules.scala 68:83:@4288.4]
  assign buffer_1_670 = $signed(_T_57396); // @[Modules.scala 68:83:@4289.4]
  assign _T_57401 = $signed(buffer_1_560) + $signed(buffer_0_561); // @[Modules.scala 68:83:@4295.4]
  assign _T_57402 = _T_57401[10:0]; // @[Modules.scala 68:83:@4296.4]
  assign buffer_1_672 = $signed(_T_57402); // @[Modules.scala 68:83:@4297.4]
  assign _T_57404 = $signed(buffer_1_562) + $signed(buffer_1_563); // @[Modules.scala 68:83:@4299.4]
  assign _T_57405 = _T_57404[10:0]; // @[Modules.scala 68:83:@4300.4]
  assign buffer_1_673 = $signed(_T_57405); // @[Modules.scala 68:83:@4301.4]
  assign _T_57407 = $signed(buffer_1_564) + $signed(buffer_1_565); // @[Modules.scala 68:83:@4303.4]
  assign _T_57408 = _T_57407[10:0]; // @[Modules.scala 68:83:@4304.4]
  assign buffer_1_674 = $signed(_T_57408); // @[Modules.scala 68:83:@4305.4]
  assign _T_57410 = $signed(buffer_1_566) + $signed(buffer_1_567); // @[Modules.scala 68:83:@4307.4]
  assign _T_57411 = _T_57410[10:0]; // @[Modules.scala 68:83:@4308.4]
  assign buffer_1_675 = $signed(_T_57411); // @[Modules.scala 68:83:@4309.4]
  assign _T_57413 = $signed(buffer_0_568) + $signed(buffer_1_569); // @[Modules.scala 68:83:@4311.4]
  assign _T_57414 = _T_57413[10:0]; // @[Modules.scala 68:83:@4312.4]
  assign buffer_1_676 = $signed(_T_57414); // @[Modules.scala 68:83:@4313.4]
  assign _T_57416 = $signed(buffer_1_570) + $signed(buffer_1_571); // @[Modules.scala 68:83:@4315.4]
  assign _T_57417 = _T_57416[10:0]; // @[Modules.scala 68:83:@4316.4]
  assign buffer_1_677 = $signed(_T_57417); // @[Modules.scala 68:83:@4317.4]
  assign _T_57419 = $signed(buffer_1_572) + $signed(buffer_1_573); // @[Modules.scala 68:83:@4319.4]
  assign _T_57420 = _T_57419[10:0]; // @[Modules.scala 68:83:@4320.4]
  assign buffer_1_678 = $signed(_T_57420); // @[Modules.scala 68:83:@4321.4]
  assign _T_57431 = $signed(buffer_0_580) + $signed(buffer_1_581); // @[Modules.scala 68:83:@4335.4]
  assign _T_57432 = _T_57431[10:0]; // @[Modules.scala 68:83:@4336.4]
  assign buffer_1_682 = $signed(_T_57432); // @[Modules.scala 68:83:@4337.4]
  assign _T_57434 = $signed(buffer_1_582) + $signed(buffer_1_583); // @[Modules.scala 68:83:@4339.4]
  assign _T_57435 = _T_57434[10:0]; // @[Modules.scala 68:83:@4340.4]
  assign buffer_1_683 = $signed(_T_57435); // @[Modules.scala 68:83:@4341.4]
  assign _T_57440 = $signed(buffer_0_395) + $signed(buffer_1_587); // @[Modules.scala 68:83:@4347.4]
  assign _T_57441 = _T_57440[10:0]; // @[Modules.scala 68:83:@4348.4]
  assign buffer_1_685 = $signed(_T_57441); // @[Modules.scala 68:83:@4349.4]
  assign _T_57443 = $signed(buffer_1_588) + $signed(buffer_1_589); // @[Modules.scala 71:109:@4351.4]
  assign _T_57444 = _T_57443[10:0]; // @[Modules.scala 71:109:@4352.4]
  assign buffer_1_686 = $signed(_T_57444); // @[Modules.scala 71:109:@4353.4]
  assign _T_57446 = $signed(buffer_1_590) + $signed(buffer_1_591); // @[Modules.scala 71:109:@4355.4]
  assign _T_57447 = _T_57446[10:0]; // @[Modules.scala 71:109:@4356.4]
  assign buffer_1_687 = $signed(_T_57447); // @[Modules.scala 71:109:@4357.4]
  assign _T_57449 = $signed(buffer_1_592) + $signed(buffer_1_593); // @[Modules.scala 71:109:@4359.4]
  assign _T_57450 = _T_57449[10:0]; // @[Modules.scala 71:109:@4360.4]
  assign buffer_1_688 = $signed(_T_57450); // @[Modules.scala 71:109:@4361.4]
  assign _T_57452 = $signed(buffer_1_594) + $signed(buffer_1_595); // @[Modules.scala 71:109:@4363.4]
  assign _T_57453 = _T_57452[10:0]; // @[Modules.scala 71:109:@4364.4]
  assign buffer_1_689 = $signed(_T_57453); // @[Modules.scala 71:109:@4365.4]
  assign _T_57455 = $signed(buffer_1_596) + $signed(buffer_1_597); // @[Modules.scala 71:109:@4367.4]
  assign _T_57456 = _T_57455[10:0]; // @[Modules.scala 71:109:@4368.4]
  assign buffer_1_690 = $signed(_T_57456); // @[Modules.scala 71:109:@4369.4]
  assign _T_57458 = $signed(buffer_1_598) + $signed(buffer_1_599); // @[Modules.scala 71:109:@4371.4]
  assign _T_57459 = _T_57458[10:0]; // @[Modules.scala 71:109:@4372.4]
  assign buffer_1_691 = $signed(_T_57459); // @[Modules.scala 71:109:@4373.4]
  assign _T_57461 = $signed(buffer_1_600) + $signed(buffer_1_601); // @[Modules.scala 71:109:@4375.4]
  assign _T_57462 = _T_57461[10:0]; // @[Modules.scala 71:109:@4376.4]
  assign buffer_1_692 = $signed(_T_57462); // @[Modules.scala 71:109:@4377.4]
  assign _T_57464 = $signed(buffer_1_602) + $signed(buffer_1_603); // @[Modules.scala 71:109:@4379.4]
  assign _T_57465 = _T_57464[10:0]; // @[Modules.scala 71:109:@4380.4]
  assign buffer_1_693 = $signed(_T_57465); // @[Modules.scala 71:109:@4381.4]
  assign _T_57467 = $signed(buffer_1_604) + $signed(buffer_1_605); // @[Modules.scala 71:109:@4383.4]
  assign _T_57468 = _T_57467[10:0]; // @[Modules.scala 71:109:@4384.4]
  assign buffer_1_694 = $signed(_T_57468); // @[Modules.scala 71:109:@4385.4]
  assign _T_57470 = $signed(buffer_1_606) + $signed(buffer_1_607); // @[Modules.scala 71:109:@4387.4]
  assign _T_57471 = _T_57470[10:0]; // @[Modules.scala 71:109:@4388.4]
  assign buffer_1_695 = $signed(_T_57471); // @[Modules.scala 71:109:@4389.4]
  assign _T_57473 = $signed(buffer_1_608) + $signed(buffer_1_609); // @[Modules.scala 71:109:@4391.4]
  assign _T_57474 = _T_57473[10:0]; // @[Modules.scala 71:109:@4392.4]
  assign buffer_1_696 = $signed(_T_57474); // @[Modules.scala 71:109:@4393.4]
  assign _T_57476 = $signed(buffer_1_610) + $signed(buffer_1_611); // @[Modules.scala 71:109:@4395.4]
  assign _T_57477 = _T_57476[10:0]; // @[Modules.scala 71:109:@4396.4]
  assign buffer_1_697 = $signed(_T_57477); // @[Modules.scala 71:109:@4397.4]
  assign _T_57479 = $signed(buffer_1_612) + $signed(buffer_1_613); // @[Modules.scala 71:109:@4399.4]
  assign _T_57480 = _T_57479[10:0]; // @[Modules.scala 71:109:@4400.4]
  assign buffer_1_698 = $signed(_T_57480); // @[Modules.scala 71:109:@4401.4]
  assign _T_57482 = $signed(buffer_1_614) + $signed(buffer_1_615); // @[Modules.scala 71:109:@4403.4]
  assign _T_57483 = _T_57482[10:0]; // @[Modules.scala 71:109:@4404.4]
  assign buffer_1_699 = $signed(_T_57483); // @[Modules.scala 71:109:@4405.4]
  assign _T_57485 = $signed(buffer_1_616) + $signed(buffer_0_593); // @[Modules.scala 71:109:@4407.4]
  assign _T_57486 = _T_57485[10:0]; // @[Modules.scala 71:109:@4408.4]
  assign buffer_1_700 = $signed(_T_57486); // @[Modules.scala 71:109:@4409.4]
  assign _T_57488 = $signed(buffer_1_618) + $signed(buffer_1_619); // @[Modules.scala 71:109:@4411.4]
  assign _T_57489 = _T_57488[10:0]; // @[Modules.scala 71:109:@4412.4]
  assign buffer_1_701 = $signed(_T_57489); // @[Modules.scala 71:109:@4413.4]
  assign _T_57491 = $signed(buffer_1_620) + $signed(buffer_1_621); // @[Modules.scala 71:109:@4415.4]
  assign _T_57492 = _T_57491[10:0]; // @[Modules.scala 71:109:@4416.4]
  assign buffer_1_702 = $signed(_T_57492); // @[Modules.scala 71:109:@4417.4]
  assign _T_57494 = $signed(buffer_1_622) + $signed(buffer_1_623); // @[Modules.scala 71:109:@4419.4]
  assign _T_57495 = _T_57494[10:0]; // @[Modules.scala 71:109:@4420.4]
  assign buffer_1_703 = $signed(_T_57495); // @[Modules.scala 71:109:@4421.4]
  assign _T_57497 = $signed(buffer_1_624) + $signed(buffer_1_625); // @[Modules.scala 71:109:@4423.4]
  assign _T_57498 = _T_57497[10:0]; // @[Modules.scala 71:109:@4424.4]
  assign buffer_1_704 = $signed(_T_57498); // @[Modules.scala 71:109:@4425.4]
  assign _T_57500 = $signed(buffer_1_626) + $signed(buffer_1_627); // @[Modules.scala 71:109:@4427.4]
  assign _T_57501 = _T_57500[10:0]; // @[Modules.scala 71:109:@4428.4]
  assign buffer_1_705 = $signed(_T_57501); // @[Modules.scala 71:109:@4429.4]
  assign _T_57503 = $signed(buffer_1_628) + $signed(buffer_1_629); // @[Modules.scala 71:109:@4431.4]
  assign _T_57504 = _T_57503[10:0]; // @[Modules.scala 71:109:@4432.4]
  assign buffer_1_706 = $signed(_T_57504); // @[Modules.scala 71:109:@4433.4]
  assign _T_57506 = $signed(buffer_0_630) + $signed(buffer_1_631); // @[Modules.scala 71:109:@4435.4]
  assign _T_57507 = _T_57506[10:0]; // @[Modules.scala 71:109:@4436.4]
  assign buffer_1_707 = $signed(_T_57507); // @[Modules.scala 71:109:@4437.4]
  assign _T_57509 = $signed(buffer_1_632) + $signed(buffer_1_633); // @[Modules.scala 71:109:@4439.4]
  assign _T_57510 = _T_57509[10:0]; // @[Modules.scala 71:109:@4440.4]
  assign buffer_1_708 = $signed(_T_57510); // @[Modules.scala 71:109:@4441.4]
  assign _T_57512 = $signed(buffer_1_634) + $signed(buffer_1_635); // @[Modules.scala 71:109:@4443.4]
  assign _T_57513 = _T_57512[10:0]; // @[Modules.scala 71:109:@4444.4]
  assign buffer_1_709 = $signed(_T_57513); // @[Modules.scala 71:109:@4445.4]
  assign _T_57515 = $signed(buffer_1_636) + $signed(buffer_1_637); // @[Modules.scala 71:109:@4447.4]
  assign _T_57516 = _T_57515[10:0]; // @[Modules.scala 71:109:@4448.4]
  assign buffer_1_710 = $signed(_T_57516); // @[Modules.scala 71:109:@4449.4]
  assign _T_57518 = $signed(buffer_1_638) + $signed(buffer_1_639); // @[Modules.scala 71:109:@4451.4]
  assign _T_57519 = _T_57518[10:0]; // @[Modules.scala 71:109:@4452.4]
  assign buffer_1_711 = $signed(_T_57519); // @[Modules.scala 71:109:@4453.4]
  assign _T_57521 = $signed(buffer_1_640) + $signed(buffer_1_641); // @[Modules.scala 71:109:@4455.4]
  assign _T_57522 = _T_57521[10:0]; // @[Modules.scala 71:109:@4456.4]
  assign buffer_1_712 = $signed(_T_57522); // @[Modules.scala 71:109:@4457.4]
  assign _T_57524 = $signed(buffer_1_642) + $signed(buffer_1_643); // @[Modules.scala 71:109:@4459.4]
  assign _T_57525 = _T_57524[10:0]; // @[Modules.scala 71:109:@4460.4]
  assign buffer_1_713 = $signed(_T_57525); // @[Modules.scala 71:109:@4461.4]
  assign _T_57527 = $signed(buffer_1_644) + $signed(buffer_1_645); // @[Modules.scala 71:109:@4463.4]
  assign _T_57528 = _T_57527[10:0]; // @[Modules.scala 71:109:@4464.4]
  assign buffer_1_714 = $signed(_T_57528); // @[Modules.scala 71:109:@4465.4]
  assign _T_57530 = $signed(buffer_1_646) + $signed(buffer_1_647); // @[Modules.scala 71:109:@4467.4]
  assign _T_57531 = _T_57530[10:0]; // @[Modules.scala 71:109:@4468.4]
  assign buffer_1_715 = $signed(_T_57531); // @[Modules.scala 71:109:@4469.4]
  assign _T_57533 = $signed(buffer_1_648) + $signed(buffer_1_649); // @[Modules.scala 71:109:@4471.4]
  assign _T_57534 = _T_57533[10:0]; // @[Modules.scala 71:109:@4472.4]
  assign buffer_1_716 = $signed(_T_57534); // @[Modules.scala 71:109:@4473.4]
  assign _T_57536 = $signed(buffer_1_650) + $signed(buffer_1_651); // @[Modules.scala 71:109:@4475.4]
  assign _T_57537 = _T_57536[10:0]; // @[Modules.scala 71:109:@4476.4]
  assign buffer_1_717 = $signed(_T_57537); // @[Modules.scala 71:109:@4477.4]
  assign _T_57539 = $signed(buffer_1_652) + $signed(buffer_1_653); // @[Modules.scala 71:109:@4479.4]
  assign _T_57540 = _T_57539[10:0]; // @[Modules.scala 71:109:@4480.4]
  assign buffer_1_718 = $signed(_T_57540); // @[Modules.scala 71:109:@4481.4]
  assign _T_57542 = $signed(buffer_1_654) + $signed(buffer_1_655); // @[Modules.scala 71:109:@4483.4]
  assign _T_57543 = _T_57542[10:0]; // @[Modules.scala 71:109:@4484.4]
  assign buffer_1_719 = $signed(_T_57543); // @[Modules.scala 71:109:@4485.4]
  assign _T_57545 = $signed(buffer_1_656) + $signed(buffer_1_657); // @[Modules.scala 71:109:@4487.4]
  assign _T_57546 = _T_57545[10:0]; // @[Modules.scala 71:109:@4488.4]
  assign buffer_1_720 = $signed(_T_57546); // @[Modules.scala 71:109:@4489.4]
  assign _T_57548 = $signed(buffer_1_658) + $signed(buffer_1_659); // @[Modules.scala 71:109:@4491.4]
  assign _T_57549 = _T_57548[10:0]; // @[Modules.scala 71:109:@4492.4]
  assign buffer_1_721 = $signed(_T_57549); // @[Modules.scala 71:109:@4493.4]
  assign _T_57551 = $signed(buffer_1_660) + $signed(buffer_1_661); // @[Modules.scala 71:109:@4495.4]
  assign _T_57552 = _T_57551[10:0]; // @[Modules.scala 71:109:@4496.4]
  assign buffer_1_722 = $signed(_T_57552); // @[Modules.scala 71:109:@4497.4]
  assign _T_57554 = $signed(buffer_1_662) + $signed(buffer_1_663); // @[Modules.scala 71:109:@4499.4]
  assign _T_57555 = _T_57554[10:0]; // @[Modules.scala 71:109:@4500.4]
  assign buffer_1_723 = $signed(_T_57555); // @[Modules.scala 71:109:@4501.4]
  assign _T_57557 = $signed(buffer_1_664) + $signed(buffer_1_665); // @[Modules.scala 71:109:@4503.4]
  assign _T_57558 = _T_57557[10:0]; // @[Modules.scala 71:109:@4504.4]
  assign buffer_1_724 = $signed(_T_57558); // @[Modules.scala 71:109:@4505.4]
  assign _T_57560 = $signed(buffer_1_666) + $signed(buffer_1_667); // @[Modules.scala 71:109:@4507.4]
  assign _T_57561 = _T_57560[10:0]; // @[Modules.scala 71:109:@4508.4]
  assign buffer_1_725 = $signed(_T_57561); // @[Modules.scala 71:109:@4509.4]
  assign _T_57563 = $signed(buffer_1_668) + $signed(buffer_1_669); // @[Modules.scala 71:109:@4511.4]
  assign _T_57564 = _T_57563[10:0]; // @[Modules.scala 71:109:@4512.4]
  assign buffer_1_726 = $signed(_T_57564); // @[Modules.scala 71:109:@4513.4]
  assign _T_57566 = $signed(buffer_1_670) + $signed(buffer_0_593); // @[Modules.scala 71:109:@4515.4]
  assign _T_57567 = _T_57566[10:0]; // @[Modules.scala 71:109:@4516.4]
  assign buffer_1_727 = $signed(_T_57567); // @[Modules.scala 71:109:@4517.4]
  assign _T_57569 = $signed(buffer_1_672) + $signed(buffer_1_673); // @[Modules.scala 71:109:@4519.4]
  assign _T_57570 = _T_57569[10:0]; // @[Modules.scala 71:109:@4520.4]
  assign buffer_1_728 = $signed(_T_57570); // @[Modules.scala 71:109:@4521.4]
  assign _T_57572 = $signed(buffer_1_674) + $signed(buffer_1_675); // @[Modules.scala 71:109:@4523.4]
  assign _T_57573 = _T_57572[10:0]; // @[Modules.scala 71:109:@4524.4]
  assign buffer_1_729 = $signed(_T_57573); // @[Modules.scala 71:109:@4525.4]
  assign _T_57575 = $signed(buffer_1_676) + $signed(buffer_1_677); // @[Modules.scala 71:109:@4527.4]
  assign _T_57576 = _T_57575[10:0]; // @[Modules.scala 71:109:@4528.4]
  assign buffer_1_730 = $signed(_T_57576); // @[Modules.scala 71:109:@4529.4]
  assign _T_57578 = $signed(buffer_1_678) + $signed(buffer_0_593); // @[Modules.scala 71:109:@4531.4]
  assign _T_57579 = _T_57578[10:0]; // @[Modules.scala 71:109:@4532.4]
  assign buffer_1_731 = $signed(_T_57579); // @[Modules.scala 71:109:@4533.4]
  assign _T_57581 = $signed(buffer_0_593) + $signed(buffer_0_681); // @[Modules.scala 71:109:@4535.4]
  assign _T_57582 = _T_57581[10:0]; // @[Modules.scala 71:109:@4536.4]
  assign buffer_1_732 = $signed(_T_57582); // @[Modules.scala 71:109:@4537.4]
  assign _T_57584 = $signed(buffer_1_682) + $signed(buffer_1_683); // @[Modules.scala 71:109:@4539.4]
  assign _T_57585 = _T_57584[10:0]; // @[Modules.scala 71:109:@4540.4]
  assign buffer_1_733 = $signed(_T_57585); // @[Modules.scala 71:109:@4541.4]
  assign _T_57587 = $signed(buffer_0_593) + $signed(buffer_1_685); // @[Modules.scala 71:109:@4543.4]
  assign _T_57588 = _T_57587[10:0]; // @[Modules.scala 71:109:@4544.4]
  assign buffer_1_734 = $signed(_T_57588); // @[Modules.scala 71:109:@4545.4]
  assign _T_57590 = $signed(buffer_1_686) + $signed(buffer_1_687); // @[Modules.scala 78:156:@4548.4]
  assign _T_57591 = _T_57590[10:0]; // @[Modules.scala 78:156:@4549.4]
  assign buffer_1_736 = $signed(_T_57591); // @[Modules.scala 78:156:@4550.4]
  assign _T_57593 = $signed(buffer_1_736) + $signed(buffer_1_688); // @[Modules.scala 78:156:@4552.4]
  assign _T_57594 = _T_57593[10:0]; // @[Modules.scala 78:156:@4553.4]
  assign buffer_1_737 = $signed(_T_57594); // @[Modules.scala 78:156:@4554.4]
  assign _T_57596 = $signed(buffer_1_737) + $signed(buffer_1_689); // @[Modules.scala 78:156:@4556.4]
  assign _T_57597 = _T_57596[10:0]; // @[Modules.scala 78:156:@4557.4]
  assign buffer_1_738 = $signed(_T_57597); // @[Modules.scala 78:156:@4558.4]
  assign _T_57599 = $signed(buffer_1_738) + $signed(buffer_1_690); // @[Modules.scala 78:156:@4560.4]
  assign _T_57600 = _T_57599[10:0]; // @[Modules.scala 78:156:@4561.4]
  assign buffer_1_739 = $signed(_T_57600); // @[Modules.scala 78:156:@4562.4]
  assign _T_57602 = $signed(buffer_1_739) + $signed(buffer_1_691); // @[Modules.scala 78:156:@4564.4]
  assign _T_57603 = _T_57602[10:0]; // @[Modules.scala 78:156:@4565.4]
  assign buffer_1_740 = $signed(_T_57603); // @[Modules.scala 78:156:@4566.4]
  assign _T_57605 = $signed(buffer_1_740) + $signed(buffer_1_692); // @[Modules.scala 78:156:@4568.4]
  assign _T_57606 = _T_57605[10:0]; // @[Modules.scala 78:156:@4569.4]
  assign buffer_1_741 = $signed(_T_57606); // @[Modules.scala 78:156:@4570.4]
  assign _T_57608 = $signed(buffer_1_741) + $signed(buffer_1_693); // @[Modules.scala 78:156:@4572.4]
  assign _T_57609 = _T_57608[10:0]; // @[Modules.scala 78:156:@4573.4]
  assign buffer_1_742 = $signed(_T_57609); // @[Modules.scala 78:156:@4574.4]
  assign _T_57611 = $signed(buffer_1_742) + $signed(buffer_1_694); // @[Modules.scala 78:156:@4576.4]
  assign _T_57612 = _T_57611[10:0]; // @[Modules.scala 78:156:@4577.4]
  assign buffer_1_743 = $signed(_T_57612); // @[Modules.scala 78:156:@4578.4]
  assign _T_57614 = $signed(buffer_1_743) + $signed(buffer_1_695); // @[Modules.scala 78:156:@4580.4]
  assign _T_57615 = _T_57614[10:0]; // @[Modules.scala 78:156:@4581.4]
  assign buffer_1_744 = $signed(_T_57615); // @[Modules.scala 78:156:@4582.4]
  assign _T_57617 = $signed(buffer_1_744) + $signed(buffer_1_696); // @[Modules.scala 78:156:@4584.4]
  assign _T_57618 = _T_57617[10:0]; // @[Modules.scala 78:156:@4585.4]
  assign buffer_1_745 = $signed(_T_57618); // @[Modules.scala 78:156:@4586.4]
  assign _T_57620 = $signed(buffer_1_745) + $signed(buffer_1_697); // @[Modules.scala 78:156:@4588.4]
  assign _T_57621 = _T_57620[10:0]; // @[Modules.scala 78:156:@4589.4]
  assign buffer_1_746 = $signed(_T_57621); // @[Modules.scala 78:156:@4590.4]
  assign _T_57623 = $signed(buffer_1_746) + $signed(buffer_1_698); // @[Modules.scala 78:156:@4592.4]
  assign _T_57624 = _T_57623[10:0]; // @[Modules.scala 78:156:@4593.4]
  assign buffer_1_747 = $signed(_T_57624); // @[Modules.scala 78:156:@4594.4]
  assign _T_57626 = $signed(buffer_1_747) + $signed(buffer_1_699); // @[Modules.scala 78:156:@4596.4]
  assign _T_57627 = _T_57626[10:0]; // @[Modules.scala 78:156:@4597.4]
  assign buffer_1_748 = $signed(_T_57627); // @[Modules.scala 78:156:@4598.4]
  assign _T_57629 = $signed(buffer_1_748) + $signed(buffer_1_700); // @[Modules.scala 78:156:@4600.4]
  assign _T_57630 = _T_57629[10:0]; // @[Modules.scala 78:156:@4601.4]
  assign buffer_1_749 = $signed(_T_57630); // @[Modules.scala 78:156:@4602.4]
  assign _T_57632 = $signed(buffer_1_749) + $signed(buffer_1_701); // @[Modules.scala 78:156:@4604.4]
  assign _T_57633 = _T_57632[10:0]; // @[Modules.scala 78:156:@4605.4]
  assign buffer_1_750 = $signed(_T_57633); // @[Modules.scala 78:156:@4606.4]
  assign _T_57635 = $signed(buffer_1_750) + $signed(buffer_1_702); // @[Modules.scala 78:156:@4608.4]
  assign _T_57636 = _T_57635[10:0]; // @[Modules.scala 78:156:@4609.4]
  assign buffer_1_751 = $signed(_T_57636); // @[Modules.scala 78:156:@4610.4]
  assign _T_57638 = $signed(buffer_1_751) + $signed(buffer_1_703); // @[Modules.scala 78:156:@4612.4]
  assign _T_57639 = _T_57638[10:0]; // @[Modules.scala 78:156:@4613.4]
  assign buffer_1_752 = $signed(_T_57639); // @[Modules.scala 78:156:@4614.4]
  assign _T_57641 = $signed(buffer_1_752) + $signed(buffer_1_704); // @[Modules.scala 78:156:@4616.4]
  assign _T_57642 = _T_57641[10:0]; // @[Modules.scala 78:156:@4617.4]
  assign buffer_1_753 = $signed(_T_57642); // @[Modules.scala 78:156:@4618.4]
  assign _T_57644 = $signed(buffer_1_753) + $signed(buffer_1_705); // @[Modules.scala 78:156:@4620.4]
  assign _T_57645 = _T_57644[10:0]; // @[Modules.scala 78:156:@4621.4]
  assign buffer_1_754 = $signed(_T_57645); // @[Modules.scala 78:156:@4622.4]
  assign _T_57647 = $signed(buffer_1_754) + $signed(buffer_1_706); // @[Modules.scala 78:156:@4624.4]
  assign _T_57648 = _T_57647[10:0]; // @[Modules.scala 78:156:@4625.4]
  assign buffer_1_755 = $signed(_T_57648); // @[Modules.scala 78:156:@4626.4]
  assign _T_57650 = $signed(buffer_1_755) + $signed(buffer_1_707); // @[Modules.scala 78:156:@4628.4]
  assign _T_57651 = _T_57650[10:0]; // @[Modules.scala 78:156:@4629.4]
  assign buffer_1_756 = $signed(_T_57651); // @[Modules.scala 78:156:@4630.4]
  assign _T_57653 = $signed(buffer_1_756) + $signed(buffer_1_708); // @[Modules.scala 78:156:@4632.4]
  assign _T_57654 = _T_57653[10:0]; // @[Modules.scala 78:156:@4633.4]
  assign buffer_1_757 = $signed(_T_57654); // @[Modules.scala 78:156:@4634.4]
  assign _T_57656 = $signed(buffer_1_757) + $signed(buffer_1_709); // @[Modules.scala 78:156:@4636.4]
  assign _T_57657 = _T_57656[10:0]; // @[Modules.scala 78:156:@4637.4]
  assign buffer_1_758 = $signed(_T_57657); // @[Modules.scala 78:156:@4638.4]
  assign _T_57659 = $signed(buffer_1_758) + $signed(buffer_1_710); // @[Modules.scala 78:156:@4640.4]
  assign _T_57660 = _T_57659[10:0]; // @[Modules.scala 78:156:@4641.4]
  assign buffer_1_759 = $signed(_T_57660); // @[Modules.scala 78:156:@4642.4]
  assign _T_57662 = $signed(buffer_1_759) + $signed(buffer_1_711); // @[Modules.scala 78:156:@4644.4]
  assign _T_57663 = _T_57662[10:0]; // @[Modules.scala 78:156:@4645.4]
  assign buffer_1_760 = $signed(_T_57663); // @[Modules.scala 78:156:@4646.4]
  assign _T_57665 = $signed(buffer_1_760) + $signed(buffer_1_712); // @[Modules.scala 78:156:@4648.4]
  assign _T_57666 = _T_57665[10:0]; // @[Modules.scala 78:156:@4649.4]
  assign buffer_1_761 = $signed(_T_57666); // @[Modules.scala 78:156:@4650.4]
  assign _T_57668 = $signed(buffer_1_761) + $signed(buffer_1_713); // @[Modules.scala 78:156:@4652.4]
  assign _T_57669 = _T_57668[10:0]; // @[Modules.scala 78:156:@4653.4]
  assign buffer_1_762 = $signed(_T_57669); // @[Modules.scala 78:156:@4654.4]
  assign _T_57671 = $signed(buffer_1_762) + $signed(buffer_1_714); // @[Modules.scala 78:156:@4656.4]
  assign _T_57672 = _T_57671[10:0]; // @[Modules.scala 78:156:@4657.4]
  assign buffer_1_763 = $signed(_T_57672); // @[Modules.scala 78:156:@4658.4]
  assign _T_57674 = $signed(buffer_1_763) + $signed(buffer_1_715); // @[Modules.scala 78:156:@4660.4]
  assign _T_57675 = _T_57674[10:0]; // @[Modules.scala 78:156:@4661.4]
  assign buffer_1_764 = $signed(_T_57675); // @[Modules.scala 78:156:@4662.4]
  assign _T_57677 = $signed(buffer_1_764) + $signed(buffer_1_716); // @[Modules.scala 78:156:@4664.4]
  assign _T_57678 = _T_57677[10:0]; // @[Modules.scala 78:156:@4665.4]
  assign buffer_1_765 = $signed(_T_57678); // @[Modules.scala 78:156:@4666.4]
  assign _T_57680 = $signed(buffer_1_765) + $signed(buffer_1_717); // @[Modules.scala 78:156:@4668.4]
  assign _T_57681 = _T_57680[10:0]; // @[Modules.scala 78:156:@4669.4]
  assign buffer_1_766 = $signed(_T_57681); // @[Modules.scala 78:156:@4670.4]
  assign _T_57683 = $signed(buffer_1_766) + $signed(buffer_1_718); // @[Modules.scala 78:156:@4672.4]
  assign _T_57684 = _T_57683[10:0]; // @[Modules.scala 78:156:@4673.4]
  assign buffer_1_767 = $signed(_T_57684); // @[Modules.scala 78:156:@4674.4]
  assign _T_57686 = $signed(buffer_1_767) + $signed(buffer_1_719); // @[Modules.scala 78:156:@4676.4]
  assign _T_57687 = _T_57686[10:0]; // @[Modules.scala 78:156:@4677.4]
  assign buffer_1_768 = $signed(_T_57687); // @[Modules.scala 78:156:@4678.4]
  assign _T_57689 = $signed(buffer_1_768) + $signed(buffer_1_720); // @[Modules.scala 78:156:@4680.4]
  assign _T_57690 = _T_57689[10:0]; // @[Modules.scala 78:156:@4681.4]
  assign buffer_1_769 = $signed(_T_57690); // @[Modules.scala 78:156:@4682.4]
  assign _T_57692 = $signed(buffer_1_769) + $signed(buffer_1_721); // @[Modules.scala 78:156:@4684.4]
  assign _T_57693 = _T_57692[10:0]; // @[Modules.scala 78:156:@4685.4]
  assign buffer_1_770 = $signed(_T_57693); // @[Modules.scala 78:156:@4686.4]
  assign _T_57695 = $signed(buffer_1_770) + $signed(buffer_1_722); // @[Modules.scala 78:156:@4688.4]
  assign _T_57696 = _T_57695[10:0]; // @[Modules.scala 78:156:@4689.4]
  assign buffer_1_771 = $signed(_T_57696); // @[Modules.scala 78:156:@4690.4]
  assign _T_57698 = $signed(buffer_1_771) + $signed(buffer_1_723); // @[Modules.scala 78:156:@4692.4]
  assign _T_57699 = _T_57698[10:0]; // @[Modules.scala 78:156:@4693.4]
  assign buffer_1_772 = $signed(_T_57699); // @[Modules.scala 78:156:@4694.4]
  assign _T_57701 = $signed(buffer_1_772) + $signed(buffer_1_724); // @[Modules.scala 78:156:@4696.4]
  assign _T_57702 = _T_57701[10:0]; // @[Modules.scala 78:156:@4697.4]
  assign buffer_1_773 = $signed(_T_57702); // @[Modules.scala 78:156:@4698.4]
  assign _T_57704 = $signed(buffer_1_773) + $signed(buffer_1_725); // @[Modules.scala 78:156:@4700.4]
  assign _T_57705 = _T_57704[10:0]; // @[Modules.scala 78:156:@4701.4]
  assign buffer_1_774 = $signed(_T_57705); // @[Modules.scala 78:156:@4702.4]
  assign _T_57707 = $signed(buffer_1_774) + $signed(buffer_1_726); // @[Modules.scala 78:156:@4704.4]
  assign _T_57708 = _T_57707[10:0]; // @[Modules.scala 78:156:@4705.4]
  assign buffer_1_775 = $signed(_T_57708); // @[Modules.scala 78:156:@4706.4]
  assign _T_57710 = $signed(buffer_1_775) + $signed(buffer_1_727); // @[Modules.scala 78:156:@4708.4]
  assign _T_57711 = _T_57710[10:0]; // @[Modules.scala 78:156:@4709.4]
  assign buffer_1_776 = $signed(_T_57711); // @[Modules.scala 78:156:@4710.4]
  assign _T_57713 = $signed(buffer_1_776) + $signed(buffer_1_728); // @[Modules.scala 78:156:@4712.4]
  assign _T_57714 = _T_57713[10:0]; // @[Modules.scala 78:156:@4713.4]
  assign buffer_1_777 = $signed(_T_57714); // @[Modules.scala 78:156:@4714.4]
  assign _T_57716 = $signed(buffer_1_777) + $signed(buffer_1_729); // @[Modules.scala 78:156:@4716.4]
  assign _T_57717 = _T_57716[10:0]; // @[Modules.scala 78:156:@4717.4]
  assign buffer_1_778 = $signed(_T_57717); // @[Modules.scala 78:156:@4718.4]
  assign _T_57719 = $signed(buffer_1_778) + $signed(buffer_1_730); // @[Modules.scala 78:156:@4720.4]
  assign _T_57720 = _T_57719[10:0]; // @[Modules.scala 78:156:@4721.4]
  assign buffer_1_779 = $signed(_T_57720); // @[Modules.scala 78:156:@4722.4]
  assign _T_57722 = $signed(buffer_1_779) + $signed(buffer_1_731); // @[Modules.scala 78:156:@4724.4]
  assign _T_57723 = _T_57722[10:0]; // @[Modules.scala 78:156:@4725.4]
  assign buffer_1_780 = $signed(_T_57723); // @[Modules.scala 78:156:@4726.4]
  assign _T_57725 = $signed(buffer_1_780) + $signed(buffer_1_732); // @[Modules.scala 78:156:@4728.4]
  assign _T_57726 = _T_57725[10:0]; // @[Modules.scala 78:156:@4729.4]
  assign buffer_1_781 = $signed(_T_57726); // @[Modules.scala 78:156:@4730.4]
  assign _T_57728 = $signed(buffer_1_781) + $signed(buffer_1_733); // @[Modules.scala 78:156:@4732.4]
  assign _T_57729 = _T_57728[10:0]; // @[Modules.scala 78:156:@4733.4]
  assign buffer_1_782 = $signed(_T_57729); // @[Modules.scala 78:156:@4734.4]
  assign _T_57731 = $signed(buffer_1_782) + $signed(buffer_1_734); // @[Modules.scala 78:156:@4736.4]
  assign _T_57732 = _T_57731[10:0]; // @[Modules.scala 78:156:@4737.4]
  assign buffer_1_783 = $signed(_T_57732); // @[Modules.scala 78:156:@4738.4]
  assign _T_57736 = $signed(io_in_10) + $signed(io_in_11); // @[Modules.scala 37:46:@4746.4]
  assign _T_57737 = _T_57736[4:0]; // @[Modules.scala 37:46:@4747.4]
  assign _T_57738 = $signed(_T_57737); // @[Modules.scala 37:46:@4748.4]
  assign _T_57741 = $signed(io_in_22) + $signed(io_in_23); // @[Modules.scala 37:46:@4755.4]
  assign _T_57742 = _T_57741[4:0]; // @[Modules.scala 37:46:@4756.4]
  assign _T_57743 = $signed(_T_57742); // @[Modules.scala 37:46:@4757.4]
  assign _T_57770 = $signed(io_in_56) + $signed(io_in_57); // @[Modules.scala 37:46:@4796.4]
  assign _T_57771 = _T_57770[4:0]; // @[Modules.scala 37:46:@4797.4]
  assign _T_57772 = $signed(_T_57771); // @[Modules.scala 37:46:@4798.4]
  assign _T_57793 = $signed(io_in_82) + $signed(io_in_83); // @[Modules.scala 37:46:@4830.4]
  assign _T_57794 = _T_57793[4:0]; // @[Modules.scala 37:46:@4831.4]
  assign _T_57795 = $signed(_T_57794); // @[Modules.scala 37:46:@4832.4]
  assign _T_57836 = $signed(io_in_160) + $signed(io_in_161); // @[Modules.scala 37:46:@4890.4]
  assign _T_57837 = _T_57836[4:0]; // @[Modules.scala 37:46:@4891.4]
  assign _T_57838 = $signed(_T_57837); // @[Modules.scala 37:46:@4892.4]
  assign _T_57842 = $signed(io_in_164) + $signed(io_in_165); // @[Modules.scala 37:46:@4898.4]
  assign _T_57843 = _T_57842[4:0]; // @[Modules.scala 37:46:@4899.4]
  assign _T_57844 = $signed(_T_57843); // @[Modules.scala 37:46:@4900.4]
  assign _T_57858 = $signed(io_in_190) + $signed(io_in_191); // @[Modules.scala 37:46:@4917.4]
  assign _T_57859 = _T_57858[4:0]; // @[Modules.scala 37:46:@4918.4]
  assign _T_57860 = $signed(_T_57859); // @[Modules.scala 37:46:@4919.4]
  assign _T_57861 = $signed(io_in_192) + $signed(io_in_193); // @[Modules.scala 37:46:@4921.4]
  assign _T_57862 = _T_57861[4:0]; // @[Modules.scala 37:46:@4922.4]
  assign _T_57863 = $signed(_T_57862); // @[Modules.scala 37:46:@4923.4]
  assign _T_57864 = $signed(io_in_194) + $signed(io_in_195); // @[Modules.scala 37:46:@4925.4]
  assign _T_57865 = _T_57864[4:0]; // @[Modules.scala 37:46:@4926.4]
  assign _T_57866 = $signed(_T_57865); // @[Modules.scala 37:46:@4927.4]
  assign _T_57876 = $signed(io_in_214) + $signed(io_in_215); // @[Modules.scala 37:46:@4941.4]
  assign _T_57877 = _T_57876[4:0]; // @[Modules.scala 37:46:@4942.4]
  assign _T_57878 = $signed(_T_57877); // @[Modules.scala 37:46:@4943.4]
  assign _T_57879 = $signed(io_in_218) + $signed(io_in_219); // @[Modules.scala 37:46:@4946.4]
  assign _T_57880 = _T_57879[4:0]; // @[Modules.scala 37:46:@4947.4]
  assign _T_57881 = $signed(_T_57880); // @[Modules.scala 37:46:@4948.4]
  assign _T_57885 = $signed(io_in_222) + $signed(io_in_223); // @[Modules.scala 37:46:@4954.4]
  assign _T_57886 = _T_57885[4:0]; // @[Modules.scala 37:46:@4955.4]
  assign _T_57887 = $signed(_T_57886); // @[Modules.scala 37:46:@4956.4]
  assign _T_57923 = $signed(io_in_288) + $signed(io_in_289); // @[Modules.scala 37:46:@5002.4]
  assign _T_57924 = _T_57923[4:0]; // @[Modules.scala 37:46:@5003.4]
  assign _T_57925 = $signed(_T_57924); // @[Modules.scala 37:46:@5004.4]
  assign _T_57926 = $signed(io_in_290) + $signed(io_in_291); // @[Modules.scala 37:46:@5006.4]
  assign _T_57927 = _T_57926[4:0]; // @[Modules.scala 37:46:@5007.4]
  assign _T_57928 = $signed(_T_57927); // @[Modules.scala 37:46:@5008.4]
  assign _T_57941 = $signed(io_in_314) + $signed(io_in_315); // @[Modules.scala 37:46:@5024.4]
  assign _T_57942 = _T_57941[4:0]; // @[Modules.scala 37:46:@5025.4]
  assign _T_57943 = $signed(_T_57942); // @[Modules.scala 37:46:@5026.4]
  assign _T_57999 = $signed(io_in_384) + $signed(io_in_385); // @[Modules.scala 37:46:@5107.4]
  assign _T_58000 = _T_57999[4:0]; // @[Modules.scala 37:46:@5108.4]
  assign _T_58001 = $signed(_T_58000); // @[Modules.scala 37:46:@5109.4]
  assign _T_58038 = $signed(io_in_422) + $signed(io_in_423); // @[Modules.scala 37:46:@5159.4]
  assign _T_58039 = _T_58038[4:0]; // @[Modules.scala 37:46:@5160.4]
  assign _T_58040 = $signed(_T_58039); // @[Modules.scala 37:46:@5161.4]
  assign _T_58066 = $signed(io_in_460) + $signed(io_in_461); // @[Modules.scala 37:46:@5196.4]
  assign _T_58067 = _T_58066[4:0]; // @[Modules.scala 37:46:@5197.4]
  assign _T_58068 = $signed(_T_58067); // @[Modules.scala 37:46:@5198.4]
  assign _T_58081 = $signed(io_in_476) + $signed(io_in_477); // @[Modules.scala 37:46:@5216.4]
  assign _T_58082 = _T_58081[4:0]; // @[Modules.scala 37:46:@5217.4]
  assign _T_58083 = $signed(_T_58082); // @[Modules.scala 37:46:@5218.4]
  assign _T_58089 = $signed(io_in_488) + $signed(io_in_489); // @[Modules.scala 37:46:@5228.4]
  assign _T_58090 = _T_58089[4:0]; // @[Modules.scala 37:46:@5229.4]
  assign _T_58091 = $signed(_T_58090); // @[Modules.scala 37:46:@5230.4]
  assign _T_58113 = $signed(io_in_516) + $signed(io_in_517); // @[Modules.scala 37:46:@5257.4]
  assign _T_58114 = _T_58113[4:0]; // @[Modules.scala 37:46:@5258.4]
  assign _T_58115 = $signed(_T_58114); // @[Modules.scala 37:46:@5259.4]
  assign _T_58126 = $signed(io_in_552) + $signed(io_in_553); // @[Modules.scala 37:46:@5278.4]
  assign _T_58127 = _T_58126[4:0]; // @[Modules.scala 37:46:@5279.4]
  assign _T_58128 = $signed(_T_58127); // @[Modules.scala 37:46:@5280.4]
  assign _T_58149 = $signed(io_in_596) + $signed(io_in_597); // @[Modules.scala 37:46:@5312.4]
  assign _T_58150 = _T_58149[4:0]; // @[Modules.scala 37:46:@5313.4]
  assign _T_58151 = $signed(_T_58150); // @[Modules.scala 37:46:@5314.4]
  assign _T_58156 = $signed(io_in_608) + $signed(io_in_609); // @[Modules.scala 37:46:@5324.4]
  assign _T_58157 = _T_58156[4:0]; // @[Modules.scala 37:46:@5325.4]
  assign _T_58158 = $signed(_T_58157); // @[Modules.scala 37:46:@5326.4]
  assign _T_58160 = $signed(io_in_616) + $signed(io_in_617); // @[Modules.scala 37:46:@5331.4]
  assign _T_58161 = _T_58160[4:0]; // @[Modules.scala 37:46:@5332.4]
  assign _T_58162 = $signed(_T_58161); // @[Modules.scala 37:46:@5333.4]
  assign _T_58172 = $signed(io_in_634) + $signed(io_in_635); // @[Modules.scala 37:46:@5346.4]
  assign _T_58173 = _T_58172[4:0]; // @[Modules.scala 37:46:@5347.4]
  assign _T_58174 = $signed(_T_58173); // @[Modules.scala 37:46:@5348.4]
  assign _T_58189 = $signed(io_in_660) + $signed(io_in_661); // @[Modules.scala 37:46:@5374.4]
  assign _T_58190 = _T_58189[4:0]; // @[Modules.scala 37:46:@5375.4]
  assign _T_58191 = $signed(_T_58190); // @[Modules.scala 37:46:@5376.4]
  assign _T_58202 = $signed(io_in_670) + $signed(io_in_671); // @[Modules.scala 37:46:@5391.4]
  assign _T_58203 = _T_58202[4:0]; // @[Modules.scala 37:46:@5392.4]
  assign _T_58204 = $signed(_T_58203); // @[Modules.scala 37:46:@5393.4]
  assign _T_58237 = $signed(io_in_728) + $signed(io_in_729); // @[Modules.scala 37:46:@5438.4]
  assign _T_58238 = _T_58237[4:0]; // @[Modules.scala 37:46:@5439.4]
  assign _T_58239 = $signed(_T_58238); // @[Modules.scala 37:46:@5440.4]
  assign _T_58240 = $signed(io_in_730) + $signed(io_in_731); // @[Modules.scala 37:46:@5442.4]
  assign _T_58241 = _T_58240[4:0]; // @[Modules.scala 37:46:@5443.4]
  assign _T_58242 = $signed(_T_58241); // @[Modules.scala 37:46:@5444.4]
  assign buffer_2_2 = {{6{io_in_4[4]}},io_in_4}; // @[Modules.scala 32:22:@8.4]
  assign _T_58269 = $signed(buffer_2_2) + $signed(11'sh0); // @[Modules.scala 65:57:@5482.4]
  assign _T_58270 = _T_58269[10:0]; // @[Modules.scala 65:57:@5483.4]
  assign buffer_2_393 = $signed(_T_58270); // @[Modules.scala 65:57:@5484.4]
  assign buffer_2_4 = {{6{io_in_8[4]}},io_in_8}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_5 = {{6{_T_57738[4]}},_T_57738}; // @[Modules.scala 32:22:@8.4]
  assign _T_58272 = $signed(buffer_2_4) + $signed(buffer_2_5); // @[Modules.scala 65:57:@5486.4]
  assign _T_58273 = _T_58272[10:0]; // @[Modules.scala 65:57:@5487.4]
  assign buffer_2_394 = $signed(_T_58273); // @[Modules.scala 65:57:@5488.4]
  assign buffer_2_9 = {{6{io_in_19[4]}},io_in_19}; // @[Modules.scala 32:22:@8.4]
  assign _T_58278 = $signed(buffer_1_8) + $signed(buffer_2_9); // @[Modules.scala 65:57:@5494.4]
  assign _T_58279 = _T_58278[10:0]; // @[Modules.scala 65:57:@5495.4]
  assign buffer_2_396 = $signed(_T_58279); // @[Modules.scala 65:57:@5496.4]
  assign buffer_2_10 = {{6{io_in_20[4]}},io_in_20}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_11 = {{6{_T_57743[4]}},_T_57743}; // @[Modules.scala 32:22:@8.4]
  assign _T_58281 = $signed(buffer_2_10) + $signed(buffer_2_11); // @[Modules.scala 65:57:@5498.4]
  assign _T_58282 = _T_58281[10:0]; // @[Modules.scala 65:57:@5499.4]
  assign buffer_2_397 = $signed(_T_58282); // @[Modules.scala 65:57:@5500.4]
  assign _T_58284 = $signed(11'sh0) + $signed(buffer_0_13); // @[Modules.scala 65:57:@5502.4]
  assign _T_58285 = _T_58284[10:0]; // @[Modules.scala 65:57:@5503.4]
  assign buffer_2_398 = $signed(_T_58285); // @[Modules.scala 65:57:@5504.4]
  assign buffer_2_15 = {{6{io_in_30[4]}},io_in_30}; // @[Modules.scala 32:22:@8.4]
  assign _T_58287 = $signed(11'sh0) + $signed(buffer_2_15); // @[Modules.scala 65:57:@5506.4]
  assign _T_58288 = _T_58287[10:0]; // @[Modules.scala 65:57:@5507.4]
  assign buffer_2_399 = $signed(_T_58288); // @[Modules.scala 65:57:@5508.4]
  assign _T_58290 = $signed(11'sh0) + $signed(buffer_1_17); // @[Modules.scala 65:57:@5510.4]
  assign _T_58291 = _T_58290[10:0]; // @[Modules.scala 65:57:@5511.4]
  assign buffer_2_400 = $signed(_T_58291); // @[Modules.scala 65:57:@5512.4]
  assign buffer_2_20 = {{6{io_in_40[4]}},io_in_40}; // @[Modules.scala 32:22:@8.4]
  assign _T_58296 = $signed(buffer_2_20) + $signed(buffer_1_21); // @[Modules.scala 65:57:@5518.4]
  assign _T_58297 = _T_58296[10:0]; // @[Modules.scala 65:57:@5519.4]
  assign buffer_2_402 = $signed(_T_58297); // @[Modules.scala 65:57:@5520.4]
  assign _T_58299 = $signed(11'sh0) + $signed(buffer_1_23); // @[Modules.scala 65:57:@5522.4]
  assign _T_58300 = _T_58299[10:0]; // @[Modules.scala 65:57:@5523.4]
  assign buffer_2_403 = $signed(_T_58300); // @[Modules.scala 65:57:@5524.4]
  assign _T_58305 = $signed(11'sh0) + $signed(buffer_1_27); // @[Modules.scala 65:57:@5530.4]
  assign _T_58306 = _T_58305[10:0]; // @[Modules.scala 65:57:@5531.4]
  assign buffer_2_405 = $signed(_T_58306); // @[Modules.scala 65:57:@5532.4]
  assign buffer_2_28 = {{6{_T_57772[4]}},_T_57772}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_29 = {{6{io_in_59[4]}},io_in_59}; // @[Modules.scala 32:22:@8.4]
  assign _T_58308 = $signed(buffer_2_28) + $signed(buffer_2_29); // @[Modules.scala 65:57:@5534.4]
  assign _T_58309 = _T_58308[10:0]; // @[Modules.scala 65:57:@5535.4]
  assign buffer_2_406 = $signed(_T_58309); // @[Modules.scala 65:57:@5536.4]
  assign buffer_2_31 = {{6{io_in_63[4]}},io_in_63}; // @[Modules.scala 32:22:@8.4]
  assign _T_58311 = $signed(11'sh0) + $signed(buffer_2_31); // @[Modules.scala 65:57:@5538.4]
  assign _T_58312 = _T_58311[10:0]; // @[Modules.scala 65:57:@5539.4]
  assign buffer_2_407 = $signed(_T_58312); // @[Modules.scala 65:57:@5540.4]
  assign buffer_2_35 = {{6{io_in_71[4]}},io_in_71}; // @[Modules.scala 32:22:@8.4]
  assign _T_58317 = $signed(buffer_1_34) + $signed(buffer_2_35); // @[Modules.scala 65:57:@5546.4]
  assign _T_58318 = _T_58317[10:0]; // @[Modules.scala 65:57:@5547.4]
  assign buffer_2_409 = $signed(_T_58318); // @[Modules.scala 65:57:@5548.4]
  assign buffer_2_39 = {{6{io_in_78[4]}},io_in_78}; // @[Modules.scala 32:22:@8.4]
  assign _T_58323 = $signed(buffer_1_38) + $signed(buffer_2_39); // @[Modules.scala 65:57:@5554.4]
  assign _T_58324 = _T_58323[10:0]; // @[Modules.scala 65:57:@5555.4]
  assign buffer_2_411 = $signed(_T_58324); // @[Modules.scala 65:57:@5556.4]
  assign buffer_2_41 = {{6{_T_57795[4]}},_T_57795}; // @[Modules.scala 32:22:@8.4]
  assign _T_58326 = $signed(11'sh0) + $signed(buffer_2_41); // @[Modules.scala 65:57:@5558.4]
  assign _T_58327 = _T_58326[10:0]; // @[Modules.scala 65:57:@5559.4]
  assign buffer_2_412 = $signed(_T_58327); // @[Modules.scala 65:57:@5560.4]
  assign _T_58329 = $signed(11'sh0) + $signed(buffer_1_43); // @[Modules.scala 65:57:@5562.4]
  assign _T_58330 = _T_58329[10:0]; // @[Modules.scala 65:57:@5563.4]
  assign buffer_2_413 = $signed(_T_58330); // @[Modules.scala 65:57:@5564.4]
  assign buffer_2_44 = {{6{io_in_88[4]}},io_in_88}; // @[Modules.scala 32:22:@8.4]
  assign _T_58332 = $signed(buffer_2_44) + $signed(buffer_0_45); // @[Modules.scala 65:57:@5566.4]
  assign _T_58333 = _T_58332[10:0]; // @[Modules.scala 65:57:@5567.4]
  assign buffer_2_414 = $signed(_T_58333); // @[Modules.scala 65:57:@5568.4]
  assign _T_58335 = $signed(buffer_1_46) + $signed(11'sh0); // @[Modules.scala 65:57:@5570.4]
  assign _T_58336 = _T_58335[10:0]; // @[Modules.scala 65:57:@5571.4]
  assign buffer_2_415 = $signed(_T_58336); // @[Modules.scala 65:57:@5572.4]
  assign buffer_2_50 = {{6{io_in_100[4]}},io_in_100}; // @[Modules.scala 32:22:@8.4]
  assign _T_58341 = $signed(buffer_2_50) + $signed(buffer_0_51); // @[Modules.scala 65:57:@5578.4]
  assign _T_58342 = _T_58341[10:0]; // @[Modules.scala 65:57:@5579.4]
  assign buffer_2_417 = $signed(_T_58342); // @[Modules.scala 65:57:@5580.4]
  assign _T_58362 = $signed(buffer_0_64) + $signed(11'sh0); // @[Modules.scala 65:57:@5606.4]
  assign _T_58363 = _T_58362[10:0]; // @[Modules.scala 65:57:@5607.4]
  assign buffer_2_424 = $signed(_T_58363); // @[Modules.scala 65:57:@5608.4]
  assign buffer_2_70 = {{6{io_in_141[4]}},io_in_141}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_71 = {{6{io_in_142[4]}},io_in_142}; // @[Modules.scala 32:22:@8.4]
  assign _T_58371 = $signed(buffer_2_70) + $signed(buffer_2_71); // @[Modules.scala 65:57:@5618.4]
  assign _T_58372 = _T_58371[10:0]; // @[Modules.scala 65:57:@5619.4]
  assign buffer_2_427 = $signed(_T_58372); // @[Modules.scala 65:57:@5620.4]
  assign buffer_2_79 = {{6{io_in_159[4]}},io_in_159}; // @[Modules.scala 32:22:@8.4]
  assign _T_58383 = $signed(11'sh0) + $signed(buffer_2_79); // @[Modules.scala 65:57:@5634.4]
  assign _T_58384 = _T_58383[10:0]; // @[Modules.scala 65:57:@5635.4]
  assign buffer_2_431 = $signed(_T_58384); // @[Modules.scala 65:57:@5636.4]
  assign buffer_2_80 = {{6{_T_57838[4]}},_T_57838}; // @[Modules.scala 32:22:@8.4]
  assign _T_58386 = $signed(buffer_2_80) + $signed(buffer_0_81); // @[Modules.scala 65:57:@5638.4]
  assign _T_58387 = _T_58386[10:0]; // @[Modules.scala 65:57:@5639.4]
  assign buffer_2_432 = $signed(_T_58387); // @[Modules.scala 65:57:@5640.4]
  assign buffer_2_82 = {{6{_T_57844[4]}},_T_57844}; // @[Modules.scala 32:22:@8.4]
  assign _T_58389 = $signed(buffer_2_82) + $signed(buffer_1_83); // @[Modules.scala 65:57:@5642.4]
  assign _T_58390 = _T_58389[10:0]; // @[Modules.scala 65:57:@5643.4]
  assign buffer_2_433 = $signed(_T_58390); // @[Modules.scala 65:57:@5644.4]
  assign buffer_2_84 = {{6{io_in_168[4]}},io_in_168}; // @[Modules.scala 32:22:@8.4]
  assign _T_58392 = $signed(buffer_2_84) + $signed(11'sh0); // @[Modules.scala 65:57:@5646.4]
  assign _T_58393 = _T_58392[10:0]; // @[Modules.scala 65:57:@5647.4]
  assign buffer_2_434 = $signed(_T_58393); // @[Modules.scala 65:57:@5648.4]
  assign buffer_2_95 = {{6{_T_57860[4]}},_T_57860}; // @[Modules.scala 32:22:@8.4]
  assign _T_58407 = $signed(11'sh0) + $signed(buffer_2_95); // @[Modules.scala 65:57:@5666.4]
  assign _T_58408 = _T_58407[10:0]; // @[Modules.scala 65:57:@5667.4]
  assign buffer_2_439 = $signed(_T_58408); // @[Modules.scala 65:57:@5668.4]
  assign buffer_2_96 = {{6{_T_57863[4]}},_T_57863}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_97 = {{6{_T_57866[4]}},_T_57866}; // @[Modules.scala 32:22:@8.4]
  assign _T_58410 = $signed(buffer_2_96) + $signed(buffer_2_97); // @[Modules.scala 65:57:@5670.4]
  assign _T_58411 = _T_58410[10:0]; // @[Modules.scala 65:57:@5671.4]
  assign buffer_2_440 = $signed(_T_58411); // @[Modules.scala 65:57:@5672.4]
  assign _T_58413 = $signed(buffer_0_98) + $signed(11'sh0); // @[Modules.scala 65:57:@5674.4]
  assign _T_58414 = _T_58413[10:0]; // @[Modules.scala 65:57:@5675.4]
  assign buffer_2_441 = $signed(_T_58414); // @[Modules.scala 65:57:@5676.4]
  assign _T_58422 = $signed(11'sh0) + $signed(buffer_0_105); // @[Modules.scala 65:57:@5686.4]
  assign _T_58423 = _T_58422[10:0]; // @[Modules.scala 65:57:@5687.4]
  assign buffer_2_444 = $signed(_T_58423); // @[Modules.scala 65:57:@5688.4]
  assign buffer_2_107 = {{6{_T_57878[4]}},_T_57878}; // @[Modules.scala 32:22:@8.4]
  assign _T_58425 = $signed(buffer_0_106) + $signed(buffer_2_107); // @[Modules.scala 65:57:@5690.4]
  assign _T_58426 = _T_58425[10:0]; // @[Modules.scala 65:57:@5691.4]
  assign buffer_2_445 = $signed(_T_58426); // @[Modules.scala 65:57:@5692.4]
  assign buffer_2_109 = {{6{_T_57881[4]}},_T_57881}; // @[Modules.scala 32:22:@8.4]
  assign _T_58428 = $signed(buffer_1_108) + $signed(buffer_2_109); // @[Modules.scala 65:57:@5694.4]
  assign _T_58429 = _T_58428[10:0]; // @[Modules.scala 65:57:@5695.4]
  assign buffer_2_446 = $signed(_T_58429); // @[Modules.scala 65:57:@5696.4]
  assign buffer_2_111 = {{6{_T_57887[4]}},_T_57887}; // @[Modules.scala 32:22:@8.4]
  assign _T_58431 = $signed(buffer_1_110) + $signed(buffer_2_111); // @[Modules.scala 65:57:@5698.4]
  assign _T_58432 = _T_58431[10:0]; // @[Modules.scala 65:57:@5699.4]
  assign buffer_2_447 = $signed(_T_58432); // @[Modules.scala 65:57:@5700.4]
  assign buffer_2_117 = {{6{io_in_235[4]}},io_in_235}; // @[Modules.scala 32:22:@8.4]
  assign _T_58440 = $signed(11'sh0) + $signed(buffer_2_117); // @[Modules.scala 65:57:@5710.4]
  assign _T_58441 = _T_58440[10:0]; // @[Modules.scala 65:57:@5711.4]
  assign buffer_2_450 = $signed(_T_58441); // @[Modules.scala 65:57:@5712.4]
  assign buffer_2_130 = {{6{io_in_261[4]}},io_in_261}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_131 = {{6{io_in_263[4]}},io_in_263}; // @[Modules.scala 32:22:@8.4]
  assign _T_58461 = $signed(buffer_2_130) + $signed(buffer_2_131); // @[Modules.scala 65:57:@5738.4]
  assign _T_58462 = _T_58461[10:0]; // @[Modules.scala 65:57:@5739.4]
  assign buffer_2_457 = $signed(_T_58462); // @[Modules.scala 65:57:@5740.4]
  assign buffer_2_143 = {{6{io_in_287[4]}},io_in_287}; // @[Modules.scala 32:22:@8.4]
  assign _T_58479 = $signed(11'sh0) + $signed(buffer_2_143); // @[Modules.scala 65:57:@5762.4]
  assign _T_58480 = _T_58479[10:0]; // @[Modules.scala 65:57:@5763.4]
  assign buffer_2_463 = $signed(_T_58480); // @[Modules.scala 65:57:@5764.4]
  assign buffer_2_144 = {{6{_T_57925[4]}},_T_57925}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_145 = {{6{_T_57928[4]}},_T_57928}; // @[Modules.scala 32:22:@8.4]
  assign _T_58482 = $signed(buffer_2_144) + $signed(buffer_2_145); // @[Modules.scala 65:57:@5766.4]
  assign _T_58483 = _T_58482[10:0]; // @[Modules.scala 65:57:@5767.4]
  assign buffer_2_464 = $signed(_T_58483); // @[Modules.scala 65:57:@5768.4]
  assign buffer_2_152 = {{6{io_in_305[4]}},io_in_305}; // @[Modules.scala 32:22:@8.4]
  assign _T_58494 = $signed(buffer_2_152) + $signed(buffer_1_153); // @[Modules.scala 65:57:@5782.4]
  assign _T_58495 = _T_58494[10:0]; // @[Modules.scala 65:57:@5783.4]
  assign buffer_2_468 = $signed(_T_58495); // @[Modules.scala 65:57:@5784.4]
  assign buffer_2_157 = {{6{_T_57943[4]}},_T_57943}; // @[Modules.scala 32:22:@8.4]
  assign _T_58500 = $signed(11'sh0) + $signed(buffer_2_157); // @[Modules.scala 65:57:@5790.4]
  assign _T_58501 = _T_58500[10:0]; // @[Modules.scala 65:57:@5791.4]
  assign buffer_2_470 = $signed(_T_58501); // @[Modules.scala 65:57:@5792.4]
  assign buffer_2_160 = {{6{io_in_320[4]}},io_in_320}; // @[Modules.scala 32:22:@8.4]
  assign _T_58506 = $signed(buffer_2_160) + $signed(buffer_1_161); // @[Modules.scala 65:57:@5798.4]
  assign _T_58507 = _T_58506[10:0]; // @[Modules.scala 65:57:@5799.4]
  assign buffer_2_472 = $signed(_T_58507); // @[Modules.scala 65:57:@5800.4]
  assign buffer_2_166 = {{6{io_in_333[4]}},io_in_333}; // @[Modules.scala 32:22:@8.4]
  assign _T_58515 = $signed(buffer_2_166) + $signed(buffer_1_167); // @[Modules.scala 65:57:@5810.4]
  assign _T_58516 = _T_58515[10:0]; // @[Modules.scala 65:57:@5811.4]
  assign buffer_2_475 = $signed(_T_58516); // @[Modules.scala 65:57:@5812.4]
  assign buffer_2_177 = {{6{io_in_354[4]}},io_in_354}; // @[Modules.scala 32:22:@8.4]
  assign _T_58530 = $signed(11'sh0) + $signed(buffer_2_177); // @[Modules.scala 65:57:@5830.4]
  assign _T_58531 = _T_58530[10:0]; // @[Modules.scala 65:57:@5831.4]
  assign buffer_2_480 = $signed(_T_58531); // @[Modules.scala 65:57:@5832.4]
  assign buffer_2_180 = {{6{io_in_361[4]}},io_in_361}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_181 = {{6{io_in_362[4]}},io_in_362}; // @[Modules.scala 32:22:@8.4]
  assign _T_58536 = $signed(buffer_2_180) + $signed(buffer_2_181); // @[Modules.scala 65:57:@5838.4]
  assign _T_58537 = _T_58536[10:0]; // @[Modules.scala 65:57:@5839.4]
  assign buffer_2_482 = $signed(_T_58537); // @[Modules.scala 65:57:@5840.4]
  assign buffer_2_192 = {{6{_T_58001[4]}},_T_58001}; // @[Modules.scala 32:22:@8.4]
  assign _T_58554 = $signed(buffer_2_192) + $signed(11'sh0); // @[Modules.scala 65:57:@5862.4]
  assign _T_58555 = _T_58554[10:0]; // @[Modules.scala 65:57:@5863.4]
  assign buffer_2_488 = $signed(_T_58555); // @[Modules.scala 65:57:@5864.4]
  assign buffer_2_205 = {{6{io_in_411[4]}},io_in_411}; // @[Modules.scala 32:22:@8.4]
  assign _T_58572 = $signed(buffer_0_204) + $signed(buffer_2_205); // @[Modules.scala 65:57:@5886.4]
  assign _T_58573 = _T_58572[10:0]; // @[Modules.scala 65:57:@5887.4]
  assign buffer_2_494 = $signed(_T_58573); // @[Modules.scala 65:57:@5888.4]
  assign buffer_2_211 = {{6{_T_58040[4]}},_T_58040}; // @[Modules.scala 32:22:@8.4]
  assign _T_58581 = $signed(buffer_0_210) + $signed(buffer_2_211); // @[Modules.scala 65:57:@5898.4]
  assign _T_58582 = _T_58581[10:0]; // @[Modules.scala 65:57:@5899.4]
  assign buffer_2_497 = $signed(_T_58582); // @[Modules.scala 65:57:@5900.4]
  assign _T_58584 = $signed(11'sh0) + $signed(buffer_0_213); // @[Modules.scala 65:57:@5902.4]
  assign _T_58585 = _T_58584[10:0]; // @[Modules.scala 65:57:@5903.4]
  assign buffer_2_498 = $signed(_T_58585); // @[Modules.scala 65:57:@5904.4]
  assign _T_58587 = $signed(buffer_0_214) + $signed(11'sh0); // @[Modules.scala 65:57:@5906.4]
  assign _T_58588 = _T_58587[10:0]; // @[Modules.scala 65:57:@5907.4]
  assign buffer_2_499 = $signed(_T_58588); // @[Modules.scala 65:57:@5908.4]
  assign _T_58596 = $signed(11'sh0) + $signed(buffer_1_221); // @[Modules.scala 65:57:@5918.4]
  assign _T_58597 = _T_58596[10:0]; // @[Modules.scala 65:57:@5919.4]
  assign buffer_2_502 = $signed(_T_58597); // @[Modules.scala 65:57:@5920.4]
  assign _T_58602 = $signed(buffer_1_224) + $signed(11'sh0); // @[Modules.scala 65:57:@5926.4]
  assign _T_58603 = _T_58602[10:0]; // @[Modules.scala 65:57:@5927.4]
  assign buffer_2_504 = $signed(_T_58603); // @[Modules.scala 65:57:@5928.4]
  assign buffer_2_227 = {{6{io_in_455[4]}},io_in_455}; // @[Modules.scala 32:22:@8.4]
  assign _T_58605 = $signed(11'sh0) + $signed(buffer_2_227); // @[Modules.scala 65:57:@5930.4]
  assign _T_58606 = _T_58605[10:0]; // @[Modules.scala 65:57:@5931.4]
  assign buffer_2_505 = $signed(_T_58606); // @[Modules.scala 65:57:@5932.4]
  assign buffer_2_228 = {{6{io_in_456[4]}},io_in_456}; // @[Modules.scala 32:22:@8.4]
  assign _T_58608 = $signed(buffer_2_228) + $signed(11'sh0); // @[Modules.scala 65:57:@5934.4]
  assign _T_58609 = _T_58608[10:0]; // @[Modules.scala 65:57:@5935.4]
  assign buffer_2_506 = $signed(_T_58609); // @[Modules.scala 65:57:@5936.4]
  assign buffer_2_230 = {{6{_T_58068[4]}},_T_58068}; // @[Modules.scala 32:22:@8.4]
  assign _T_58611 = $signed(buffer_2_230) + $signed(buffer_0_231); // @[Modules.scala 65:57:@5938.4]
  assign _T_58612 = _T_58611[10:0]; // @[Modules.scala 65:57:@5939.4]
  assign buffer_2_507 = $signed(_T_58612); // @[Modules.scala 65:57:@5940.4]
  assign buffer_2_232 = {{6{io_in_465[4]}},io_in_465}; // @[Modules.scala 32:22:@8.4]
  assign _T_58614 = $signed(buffer_2_232) + $signed(buffer_0_233); // @[Modules.scala 65:57:@5942.4]
  assign _T_58615 = _T_58614[10:0]; // @[Modules.scala 65:57:@5943.4]
  assign buffer_2_508 = $signed(_T_58615); // @[Modules.scala 65:57:@5944.4]
  assign _T_58617 = $signed(11'sh0) + $signed(buffer_1_235); // @[Modules.scala 65:57:@5946.4]
  assign _T_58618 = _T_58617[10:0]; // @[Modules.scala 65:57:@5947.4]
  assign buffer_2_509 = $signed(_T_58618); // @[Modules.scala 65:57:@5948.4]
  assign buffer_2_238 = {{6{_T_58083[4]}},_T_58083}; // @[Modules.scala 32:22:@8.4]
  assign _T_58623 = $signed(buffer_2_238) + $signed(buffer_0_239); // @[Modules.scala 65:57:@5954.4]
  assign _T_58624 = _T_58623[10:0]; // @[Modules.scala 65:57:@5955.4]
  assign buffer_2_511 = $signed(_T_58624); // @[Modules.scala 65:57:@5956.4]
  assign buffer_2_242 = {{6{io_in_485[4]}},io_in_485}; // @[Modules.scala 32:22:@8.4]
  assign _T_58629 = $signed(buffer_2_242) + $signed(buffer_0_243); // @[Modules.scala 65:57:@5962.4]
  assign _T_58630 = _T_58629[10:0]; // @[Modules.scala 65:57:@5963.4]
  assign buffer_2_513 = $signed(_T_58630); // @[Modules.scala 65:57:@5964.4]
  assign buffer_2_244 = {{6{_T_58091[4]}},_T_58091}; // @[Modules.scala 32:22:@8.4]
  assign _T_58632 = $signed(buffer_2_244) + $signed(buffer_0_245); // @[Modules.scala 65:57:@5966.4]
  assign _T_58633 = _T_58632[10:0]; // @[Modules.scala 65:57:@5967.4]
  assign buffer_2_514 = $signed(_T_58633); // @[Modules.scala 65:57:@5968.4]
  assign _T_58638 = $signed(buffer_1_248) + $signed(11'sh0); // @[Modules.scala 65:57:@5974.4]
  assign _T_58639 = _T_58638[10:0]; // @[Modules.scala 65:57:@5975.4]
  assign buffer_2_516 = $signed(_T_58639); // @[Modules.scala 65:57:@5976.4]
  assign buffer_2_258 = {{6{_T_58115[4]}},_T_58115}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_259 = {{6{io_in_518[4]}},io_in_518}; // @[Modules.scala 32:22:@8.4]
  assign _T_58653 = $signed(buffer_2_258) + $signed(buffer_2_259); // @[Modules.scala 65:57:@5994.4]
  assign _T_58654 = _T_58653[10:0]; // @[Modules.scala 65:57:@5995.4]
  assign buffer_2_521 = $signed(_T_58654); // @[Modules.scala 65:57:@5996.4]
  assign _T_58656 = $signed(11'sh0) + $signed(buffer_0_261); // @[Modules.scala 65:57:@5998.4]
  assign _T_58657 = _T_58656[10:0]; // @[Modules.scala 65:57:@5999.4]
  assign buffer_2_522 = $signed(_T_58657); // @[Modules.scala 65:57:@6000.4]
  assign buffer_2_272 = {{6{io_in_545[4]}},io_in_545}; // @[Modules.scala 32:22:@8.4]
  assign _T_58674 = $signed(buffer_2_272) + $signed(buffer_1_273); // @[Modules.scala 65:57:@6022.4]
  assign _T_58675 = _T_58674[10:0]; // @[Modules.scala 65:57:@6023.4]
  assign buffer_2_528 = $signed(_T_58675); // @[Modules.scala 65:57:@6024.4]
  assign buffer_2_274 = {{6{io_in_549[4]}},io_in_549}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_275 = {{6{io_in_551[4]}},io_in_551}; // @[Modules.scala 32:22:@8.4]
  assign _T_58677 = $signed(buffer_2_274) + $signed(buffer_2_275); // @[Modules.scala 65:57:@6026.4]
  assign _T_58678 = _T_58677[10:0]; // @[Modules.scala 65:57:@6027.4]
  assign buffer_2_529 = $signed(_T_58678); // @[Modules.scala 65:57:@6028.4]
  assign buffer_2_276 = {{6{_T_58128[4]}},_T_58128}; // @[Modules.scala 32:22:@8.4]
  assign _T_58680 = $signed(buffer_2_276) + $signed(11'sh0); // @[Modules.scala 65:57:@6030.4]
  assign _T_58681 = _T_58680[10:0]; // @[Modules.scala 65:57:@6031.4]
  assign buffer_2_530 = $signed(_T_58681); // @[Modules.scala 65:57:@6032.4]
  assign _T_58683 = $signed(11'sh0) + $signed(buffer_0_279); // @[Modules.scala 65:57:@6034.4]
  assign _T_58684 = _T_58683[10:0]; // @[Modules.scala 65:57:@6035.4]
  assign buffer_2_531 = $signed(_T_58684); // @[Modules.scala 65:57:@6036.4]
  assign buffer_2_280 = {{6{io_in_560[4]}},io_in_560}; // @[Modules.scala 32:22:@8.4]
  assign _T_58686 = $signed(buffer_2_280) + $signed(11'sh0); // @[Modules.scala 65:57:@6038.4]
  assign _T_58687 = _T_58686[10:0]; // @[Modules.scala 65:57:@6039.4]
  assign buffer_2_532 = $signed(_T_58687); // @[Modules.scala 65:57:@6040.4]
  assign _T_58695 = $signed(11'sh0) + $signed(buffer_1_287); // @[Modules.scala 65:57:@6050.4]
  assign _T_58696 = _T_58695[10:0]; // @[Modules.scala 65:57:@6051.4]
  assign buffer_2_535 = $signed(_T_58696); // @[Modules.scala 65:57:@6052.4]
  assign _T_58698 = $signed(buffer_0_288) + $signed(buffer_1_289); // @[Modules.scala 65:57:@6054.4]
  assign _T_58699 = _T_58698[10:0]; // @[Modules.scala 65:57:@6055.4]
  assign buffer_2_536 = $signed(_T_58699); // @[Modules.scala 65:57:@6056.4]
  assign buffer_2_294 = {{6{io_in_588[4]}},io_in_588}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_295 = {{6{io_in_590[4]}},io_in_590}; // @[Modules.scala 32:22:@8.4]
  assign _T_58707 = $signed(buffer_2_294) + $signed(buffer_2_295); // @[Modules.scala 65:57:@6066.4]
  assign _T_58708 = _T_58707[10:0]; // @[Modules.scala 65:57:@6067.4]
  assign buffer_2_539 = $signed(_T_58708); // @[Modules.scala 65:57:@6068.4]
  assign buffer_2_297 = {{6{io_in_595[4]}},io_in_595}; // @[Modules.scala 32:22:@8.4]
  assign _T_58710 = $signed(11'sh0) + $signed(buffer_2_297); // @[Modules.scala 65:57:@6070.4]
  assign _T_58711 = _T_58710[10:0]; // @[Modules.scala 65:57:@6071.4]
  assign buffer_2_540 = $signed(_T_58711); // @[Modules.scala 65:57:@6072.4]
  assign buffer_2_298 = {{6{_T_58151[4]}},_T_58151}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_299 = {{6{io_in_598[4]}},io_in_598}; // @[Modules.scala 32:22:@8.4]
  assign _T_58713 = $signed(buffer_2_298) + $signed(buffer_2_299); // @[Modules.scala 65:57:@6074.4]
  assign _T_58714 = _T_58713[10:0]; // @[Modules.scala 65:57:@6075.4]
  assign buffer_2_541 = $signed(_T_58714); // @[Modules.scala 65:57:@6076.4]
  assign buffer_2_300 = {{6{io_in_601[4]}},io_in_601}; // @[Modules.scala 32:22:@8.4]
  assign _T_58716 = $signed(buffer_2_300) + $signed(buffer_1_301); // @[Modules.scala 65:57:@6078.4]
  assign _T_58717 = _T_58716[10:0]; // @[Modules.scala 65:57:@6079.4]
  assign buffer_2_542 = $signed(_T_58717); // @[Modules.scala 65:57:@6080.4]
  assign buffer_2_302 = {{6{io_in_605[4]}},io_in_605}; // @[Modules.scala 32:22:@8.4]
  assign _T_58719 = $signed(buffer_2_302) + $signed(11'sh0); // @[Modules.scala 65:57:@6082.4]
  assign _T_58720 = _T_58719[10:0]; // @[Modules.scala 65:57:@6083.4]
  assign buffer_2_543 = $signed(_T_58720); // @[Modules.scala 65:57:@6084.4]
  assign buffer_2_304 = {{6{_T_58158[4]}},_T_58158}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_305 = {{6{io_in_610[4]}},io_in_610}; // @[Modules.scala 32:22:@8.4]
  assign _T_58722 = $signed(buffer_2_304) + $signed(buffer_2_305); // @[Modules.scala 65:57:@6086.4]
  assign _T_58723 = _T_58722[10:0]; // @[Modules.scala 65:57:@6087.4]
  assign buffer_2_544 = $signed(_T_58723); // @[Modules.scala 65:57:@6088.4]
  assign buffer_2_308 = {{6{_T_58162[4]}},_T_58162}; // @[Modules.scala 32:22:@8.4]
  assign _T_58728 = $signed(buffer_2_308) + $signed(11'sh0); // @[Modules.scala 65:57:@6094.4]
  assign _T_58729 = _T_58728[10:0]; // @[Modules.scala 65:57:@6095.4]
  assign buffer_2_546 = $signed(_T_58729); // @[Modules.scala 65:57:@6096.4]
  assign buffer_2_312 = {{6{io_in_624[4]}},io_in_624}; // @[Modules.scala 32:22:@8.4]
  assign _T_58734 = $signed(buffer_2_312) + $signed(11'sh0); // @[Modules.scala 65:57:@6102.4]
  assign _T_58735 = _T_58734[10:0]; // @[Modules.scala 65:57:@6103.4]
  assign buffer_2_548 = $signed(_T_58735); // @[Modules.scala 65:57:@6104.4]
  assign buffer_2_317 = {{6{_T_58174[4]}},_T_58174}; // @[Modules.scala 32:22:@8.4]
  assign _T_58740 = $signed(buffer_1_316) + $signed(buffer_2_317); // @[Modules.scala 65:57:@6110.4]
  assign _T_58741 = _T_58740[10:0]; // @[Modules.scala 65:57:@6111.4]
  assign buffer_2_550 = $signed(_T_58741); // @[Modules.scala 65:57:@6112.4]
  assign buffer_2_322 = {{6{io_in_644[4]}},io_in_644}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_323 = {{6{io_in_646[4]}},io_in_646}; // @[Modules.scala 32:22:@8.4]
  assign _T_58749 = $signed(buffer_2_322) + $signed(buffer_2_323); // @[Modules.scala 65:57:@6122.4]
  assign _T_58750 = _T_58749[10:0]; // @[Modules.scala 65:57:@6123.4]
  assign buffer_2_553 = $signed(_T_58750); // @[Modules.scala 65:57:@6124.4]
  assign buffer_2_324 = {{6{io_in_649[4]}},io_in_649}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_325 = {{6{io_in_650[4]}},io_in_650}; // @[Modules.scala 32:22:@8.4]
  assign _T_58752 = $signed(buffer_2_324) + $signed(buffer_2_325); // @[Modules.scala 65:57:@6126.4]
  assign _T_58753 = _T_58752[10:0]; // @[Modules.scala 65:57:@6127.4]
  assign buffer_2_554 = $signed(_T_58753); // @[Modules.scala 65:57:@6128.4]
  assign _T_58755 = $signed(buffer_1_326) + $signed(11'sh0); // @[Modules.scala 65:57:@6130.4]
  assign _T_58756 = _T_58755[10:0]; // @[Modules.scala 65:57:@6131.4]
  assign buffer_2_555 = $signed(_T_58756); // @[Modules.scala 65:57:@6132.4]
  assign buffer_2_328 = {{6{io_in_656[4]}},io_in_656}; // @[Modules.scala 32:22:@8.4]
  assign _T_58758 = $signed(buffer_2_328) + $signed(buffer_1_329); // @[Modules.scala 65:57:@6134.4]
  assign _T_58759 = _T_58758[10:0]; // @[Modules.scala 65:57:@6135.4]
  assign buffer_2_556 = $signed(_T_58759); // @[Modules.scala 65:57:@6136.4]
  assign buffer_2_330 = {{6{_T_58191[4]}},_T_58191}; // @[Modules.scala 32:22:@8.4]
  assign _T_58761 = $signed(buffer_2_330) + $signed(buffer_1_331); // @[Modules.scala 65:57:@6138.4]
  assign _T_58762 = _T_58761[10:0]; // @[Modules.scala 65:57:@6139.4]
  assign buffer_2_557 = $signed(_T_58762); // @[Modules.scala 65:57:@6140.4]
  assign buffer_2_335 = {{6{_T_58204[4]}},_T_58204}; // @[Modules.scala 32:22:@8.4]
  assign _T_58767 = $signed(11'sh0) + $signed(buffer_2_335); // @[Modules.scala 65:57:@6146.4]
  assign _T_58768 = _T_58767[10:0]; // @[Modules.scala 65:57:@6147.4]
  assign buffer_2_559 = $signed(_T_58768); // @[Modules.scala 65:57:@6148.4]
  assign _T_58770 = $signed(11'sh0) + $signed(buffer_0_337); // @[Modules.scala 65:57:@6150.4]
  assign _T_58771 = _T_58770[10:0]; // @[Modules.scala 65:57:@6151.4]
  assign buffer_2_560 = $signed(_T_58771); // @[Modules.scala 65:57:@6152.4]
  assign buffer_2_342 = {{6{io_in_684[4]}},io_in_684}; // @[Modules.scala 32:22:@8.4]
  assign _T_58779 = $signed(buffer_2_342) + $signed(11'sh0); // @[Modules.scala 65:57:@6162.4]
  assign _T_58780 = _T_58779[10:0]; // @[Modules.scala 65:57:@6163.4]
  assign buffer_2_563 = $signed(_T_58780); // @[Modules.scala 65:57:@6164.4]
  assign buffer_2_344 = {{6{io_in_689[4]}},io_in_689}; // @[Modules.scala 32:22:@8.4]
  assign _T_58782 = $signed(buffer_2_344) + $signed(buffer_0_345); // @[Modules.scala 65:57:@6166.4]
  assign _T_58783 = _T_58782[10:0]; // @[Modules.scala 65:57:@6167.4]
  assign buffer_2_564 = $signed(_T_58783); // @[Modules.scala 65:57:@6168.4]
  assign _T_58788 = $signed(11'sh0) + $signed(buffer_0_349); // @[Modules.scala 65:57:@6174.4]
  assign _T_58789 = _T_58788[10:0]; // @[Modules.scala 65:57:@6175.4]
  assign buffer_2_566 = $signed(_T_58789); // @[Modules.scala 65:57:@6176.4]
  assign _T_58791 = $signed(11'sh0) + $signed(buffer_0_351); // @[Modules.scala 65:57:@6178.4]
  assign _T_58792 = _T_58791[10:0]; // @[Modules.scala 65:57:@6179.4]
  assign buffer_2_567 = $signed(_T_58792); // @[Modules.scala 65:57:@6180.4]
  assign buffer_2_364 = {{6{_T_58239[4]}},_T_58239}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_365 = {{6{_T_58242[4]}},_T_58242}; // @[Modules.scala 32:22:@8.4]
  assign _T_58812 = $signed(buffer_2_364) + $signed(buffer_2_365); // @[Modules.scala 65:57:@6206.4]
  assign _T_58813 = _T_58812[10:0]; // @[Modules.scala 65:57:@6207.4]
  assign buffer_2_574 = $signed(_T_58813); // @[Modules.scala 65:57:@6208.4]
  assign buffer_2_366 = {{6{io_in_732[4]}},io_in_732}; // @[Modules.scala 32:22:@8.4]
  assign _T_58815 = $signed(buffer_2_366) + $signed(11'sh0); // @[Modules.scala 65:57:@6210.4]
  assign _T_58816 = _T_58815[10:0]; // @[Modules.scala 65:57:@6211.4]
  assign buffer_2_575 = $signed(_T_58816); // @[Modules.scala 65:57:@6212.4]
  assign buffer_2_374 = {{6{io_in_748[4]}},io_in_748}; // @[Modules.scala 32:22:@8.4]
  assign buffer_2_375 = {{6{io_in_751[4]}},io_in_751}; // @[Modules.scala 32:22:@8.4]
  assign _T_58827 = $signed(buffer_2_374) + $signed(buffer_2_375); // @[Modules.scala 65:57:@6226.4]
  assign _T_58828 = _T_58827[10:0]; // @[Modules.scala 65:57:@6227.4]
  assign buffer_2_579 = $signed(_T_58828); // @[Modules.scala 65:57:@6228.4]
  assign buffer_2_377 = {{6{io_in_754[4]}},io_in_754}; // @[Modules.scala 32:22:@8.4]
  assign _T_58830 = $signed(buffer_0_376) + $signed(buffer_2_377); // @[Modules.scala 65:57:@6230.4]
  assign _T_58831 = _T_58830[10:0]; // @[Modules.scala 65:57:@6231.4]
  assign buffer_2_580 = $signed(_T_58831); // @[Modules.scala 65:57:@6232.4]
  assign _T_58833 = $signed(11'sh0) + $signed(buffer_1_379); // @[Modules.scala 65:57:@6234.4]
  assign _T_58834 = _T_58833[10:0]; // @[Modules.scala 65:57:@6235.4]
  assign buffer_2_581 = $signed(_T_58834); // @[Modules.scala 65:57:@6236.4]
  assign buffer_2_391 = {{6{io_in_783[4]}},io_in_783}; // @[Modules.scala 32:22:@8.4]
  assign _T_58851 = $signed(buffer_1_390) + $signed(buffer_2_391); // @[Modules.scala 65:57:@6258.4]
  assign _T_58852 = _T_58851[10:0]; // @[Modules.scala 65:57:@6259.4]
  assign buffer_2_587 = $signed(_T_58852); // @[Modules.scala 65:57:@6260.4]
  assign _T_58854 = $signed(buffer_0_392) + $signed(buffer_2_393); // @[Modules.scala 68:83:@6262.4]
  assign _T_58855 = _T_58854[10:0]; // @[Modules.scala 68:83:@6263.4]
  assign buffer_2_588 = $signed(_T_58855); // @[Modules.scala 68:83:@6264.4]
  assign _T_58857 = $signed(buffer_2_394) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6266.4]
  assign _T_58858 = _T_58857[10:0]; // @[Modules.scala 68:83:@6267.4]
  assign buffer_2_589 = $signed(_T_58858); // @[Modules.scala 68:83:@6268.4]
  assign _T_58860 = $signed(buffer_2_396) + $signed(buffer_2_397); // @[Modules.scala 68:83:@6270.4]
  assign _T_58861 = _T_58860[10:0]; // @[Modules.scala 68:83:@6271.4]
  assign buffer_2_590 = $signed(_T_58861); // @[Modules.scala 68:83:@6272.4]
  assign _T_58863 = $signed(buffer_2_398) + $signed(buffer_2_399); // @[Modules.scala 68:83:@6274.4]
  assign _T_58864 = _T_58863[10:0]; // @[Modules.scala 68:83:@6275.4]
  assign buffer_2_591 = $signed(_T_58864); // @[Modules.scala 68:83:@6276.4]
  assign _T_58866 = $signed(buffer_2_400) + $signed(buffer_1_401); // @[Modules.scala 68:83:@6278.4]
  assign _T_58867 = _T_58866[10:0]; // @[Modules.scala 68:83:@6279.4]
  assign buffer_2_592 = $signed(_T_58867); // @[Modules.scala 68:83:@6280.4]
  assign _T_58869 = $signed(buffer_2_402) + $signed(buffer_2_403); // @[Modules.scala 68:83:@6282.4]
  assign _T_58870 = _T_58869[10:0]; // @[Modules.scala 68:83:@6283.4]
  assign buffer_2_593 = $signed(_T_58870); // @[Modules.scala 68:83:@6284.4]
  assign _T_58872 = $signed(buffer_1_404) + $signed(buffer_2_405); // @[Modules.scala 68:83:@6286.4]
  assign _T_58873 = _T_58872[10:0]; // @[Modules.scala 68:83:@6287.4]
  assign buffer_2_594 = $signed(_T_58873); // @[Modules.scala 68:83:@6288.4]
  assign _T_58875 = $signed(buffer_2_406) + $signed(buffer_2_407); // @[Modules.scala 68:83:@6290.4]
  assign _T_58876 = _T_58875[10:0]; // @[Modules.scala 68:83:@6291.4]
  assign buffer_2_595 = $signed(_T_58876); // @[Modules.scala 68:83:@6292.4]
  assign _T_58878 = $signed(buffer_1_408) + $signed(buffer_2_409); // @[Modules.scala 68:83:@6294.4]
  assign _T_58879 = _T_58878[10:0]; // @[Modules.scala 68:83:@6295.4]
  assign buffer_2_596 = $signed(_T_58879); // @[Modules.scala 68:83:@6296.4]
  assign _T_58881 = $signed(buffer_1_410) + $signed(buffer_2_411); // @[Modules.scala 68:83:@6298.4]
  assign _T_58882 = _T_58881[10:0]; // @[Modules.scala 68:83:@6299.4]
  assign buffer_2_597 = $signed(_T_58882); // @[Modules.scala 68:83:@6300.4]
  assign _T_58884 = $signed(buffer_2_412) + $signed(buffer_2_413); // @[Modules.scala 68:83:@6302.4]
  assign _T_58885 = _T_58884[10:0]; // @[Modules.scala 68:83:@6303.4]
  assign buffer_2_598 = $signed(_T_58885); // @[Modules.scala 68:83:@6304.4]
  assign _T_58887 = $signed(buffer_2_414) + $signed(buffer_2_415); // @[Modules.scala 68:83:@6306.4]
  assign _T_58888 = _T_58887[10:0]; // @[Modules.scala 68:83:@6307.4]
  assign buffer_2_599 = $signed(_T_58888); // @[Modules.scala 68:83:@6308.4]
  assign _T_58890 = $signed(buffer_0_395) + $signed(buffer_2_417); // @[Modules.scala 68:83:@6310.4]
  assign _T_58891 = _T_58890[10:0]; // @[Modules.scala 68:83:@6311.4]
  assign buffer_2_600 = $signed(_T_58891); // @[Modules.scala 68:83:@6312.4]
  assign _T_58893 = $signed(buffer_0_418) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6314.4]
  assign _T_58894 = _T_58893[10:0]; // @[Modules.scala 68:83:@6315.4]
  assign buffer_2_601 = $signed(_T_58894); // @[Modules.scala 68:83:@6316.4]
  assign _T_58896 = $signed(buffer_0_420) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6318.4]
  assign _T_58897 = _T_58896[10:0]; // @[Modules.scala 68:83:@6319.4]
  assign buffer_2_602 = $signed(_T_58897); // @[Modules.scala 68:83:@6320.4]
  assign _T_58902 = $signed(buffer_2_424) + $signed(buffer_1_425); // @[Modules.scala 68:83:@6326.4]
  assign _T_58903 = _T_58902[10:0]; // @[Modules.scala 68:83:@6327.4]
  assign buffer_2_604 = $signed(_T_58903); // @[Modules.scala 68:83:@6328.4]
  assign _T_58905 = $signed(buffer_0_426) + $signed(buffer_2_427); // @[Modules.scala 68:83:@6330.4]
  assign _T_58906 = _T_58905[10:0]; // @[Modules.scala 68:83:@6331.4]
  assign buffer_2_605 = $signed(_T_58906); // @[Modules.scala 68:83:@6332.4]
  assign _T_58911 = $signed(buffer_0_395) + $signed(buffer_2_431); // @[Modules.scala 68:83:@6338.4]
  assign _T_58912 = _T_58911[10:0]; // @[Modules.scala 68:83:@6339.4]
  assign buffer_2_607 = $signed(_T_58912); // @[Modules.scala 68:83:@6340.4]
  assign _T_58914 = $signed(buffer_2_432) + $signed(buffer_2_433); // @[Modules.scala 68:83:@6342.4]
  assign _T_58915 = _T_58914[10:0]; // @[Modules.scala 68:83:@6343.4]
  assign buffer_2_608 = $signed(_T_58915); // @[Modules.scala 68:83:@6344.4]
  assign _T_58917 = $signed(buffer_2_434) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6346.4]
  assign _T_58918 = _T_58917[10:0]; // @[Modules.scala 68:83:@6347.4]
  assign buffer_2_609 = $signed(_T_58918); // @[Modules.scala 68:83:@6348.4]
  assign _T_58923 = $signed(buffer_0_395) + $signed(buffer_2_439); // @[Modules.scala 68:83:@6354.4]
  assign _T_58924 = _T_58923[10:0]; // @[Modules.scala 68:83:@6355.4]
  assign buffer_2_611 = $signed(_T_58924); // @[Modules.scala 68:83:@6356.4]
  assign _T_58926 = $signed(buffer_2_440) + $signed(buffer_2_441); // @[Modules.scala 68:83:@6358.4]
  assign _T_58927 = _T_58926[10:0]; // @[Modules.scala 68:83:@6359.4]
  assign buffer_2_612 = $signed(_T_58927); // @[Modules.scala 68:83:@6360.4]
  assign _T_58932 = $signed(buffer_2_444) + $signed(buffer_2_445); // @[Modules.scala 68:83:@6366.4]
  assign _T_58933 = _T_58932[10:0]; // @[Modules.scala 68:83:@6367.4]
  assign buffer_2_614 = $signed(_T_58933); // @[Modules.scala 68:83:@6368.4]
  assign _T_58935 = $signed(buffer_2_446) + $signed(buffer_2_447); // @[Modules.scala 68:83:@6370.4]
  assign _T_58936 = _T_58935[10:0]; // @[Modules.scala 68:83:@6371.4]
  assign buffer_2_615 = $signed(_T_58936); // @[Modules.scala 68:83:@6372.4]
  assign _T_58941 = $signed(buffer_2_450) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6378.4]
  assign _T_58942 = _T_58941[10:0]; // @[Modules.scala 68:83:@6379.4]
  assign buffer_2_617 = $signed(_T_58942); // @[Modules.scala 68:83:@6380.4]
  assign _T_58944 = $signed(buffer_0_395) + $signed(buffer_1_453); // @[Modules.scala 68:83:@6382.4]
  assign _T_58945 = _T_58944[10:0]; // @[Modules.scala 68:83:@6383.4]
  assign buffer_2_618 = $signed(_T_58945); // @[Modules.scala 68:83:@6384.4]
  assign _T_58947 = $signed(buffer_1_454) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6386.4]
  assign _T_58948 = _T_58947[10:0]; // @[Modules.scala 68:83:@6387.4]
  assign buffer_2_619 = $signed(_T_58948); // @[Modules.scala 68:83:@6388.4]
  assign _T_58950 = $signed(buffer_0_395) + $signed(buffer_2_457); // @[Modules.scala 68:83:@6390.4]
  assign _T_58951 = _T_58950[10:0]; // @[Modules.scala 68:83:@6391.4]
  assign buffer_2_620 = $signed(_T_58951); // @[Modules.scala 68:83:@6392.4]
  assign _T_58956 = $signed(buffer_0_395) + $signed(buffer_1_461); // @[Modules.scala 68:83:@6398.4]
  assign _T_58957 = _T_58956[10:0]; // @[Modules.scala 68:83:@6399.4]
  assign buffer_2_622 = $signed(_T_58957); // @[Modules.scala 68:83:@6400.4]
  assign _T_58959 = $signed(buffer_0_395) + $signed(buffer_2_463); // @[Modules.scala 68:83:@6402.4]
  assign _T_58960 = _T_58959[10:0]; // @[Modules.scala 68:83:@6403.4]
  assign buffer_2_623 = $signed(_T_58960); // @[Modules.scala 68:83:@6404.4]
  assign _T_58962 = $signed(buffer_2_464) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6406.4]
  assign _T_58963 = _T_58962[10:0]; // @[Modules.scala 68:83:@6407.4]
  assign buffer_2_624 = $signed(_T_58963); // @[Modules.scala 68:83:@6408.4]
  assign _T_58968 = $signed(buffer_2_468) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6414.4]
  assign _T_58969 = _T_58968[10:0]; // @[Modules.scala 68:83:@6415.4]
  assign buffer_2_626 = $signed(_T_58969); // @[Modules.scala 68:83:@6416.4]
  assign _T_58971 = $signed(buffer_2_470) + $signed(buffer_0_471); // @[Modules.scala 68:83:@6418.4]
  assign _T_58972 = _T_58971[10:0]; // @[Modules.scala 68:83:@6419.4]
  assign buffer_2_627 = $signed(_T_58972); // @[Modules.scala 68:83:@6420.4]
  assign _T_58974 = $signed(buffer_2_472) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6422.4]
  assign _T_58975 = _T_58974[10:0]; // @[Modules.scala 68:83:@6423.4]
  assign buffer_2_628 = $signed(_T_58975); // @[Modules.scala 68:83:@6424.4]
  assign _T_58977 = $signed(buffer_0_395) + $signed(buffer_2_475); // @[Modules.scala 68:83:@6426.4]
  assign _T_58978 = _T_58977[10:0]; // @[Modules.scala 68:83:@6427.4]
  assign buffer_2_629 = $signed(_T_58978); // @[Modules.scala 68:83:@6428.4]
  assign _T_58986 = $signed(buffer_2_480) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6438.4]
  assign _T_58987 = _T_58986[10:0]; // @[Modules.scala 68:83:@6439.4]
  assign buffer_2_632 = $signed(_T_58987); // @[Modules.scala 68:83:@6440.4]
  assign _T_58989 = $signed(buffer_2_482) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6442.4]
  assign _T_58990 = _T_58989[10:0]; // @[Modules.scala 68:83:@6443.4]
  assign buffer_2_633 = $signed(_T_58990); // @[Modules.scala 68:83:@6444.4]
  assign _T_58998 = $signed(buffer_2_488) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6454.4]
  assign _T_58999 = _T_58998[10:0]; // @[Modules.scala 68:83:@6455.4]
  assign buffer_2_636 = $signed(_T_58999); // @[Modules.scala 68:83:@6456.4]
  assign _T_59001 = $signed(buffer_1_490) + $signed(buffer_0_491); // @[Modules.scala 68:83:@6458.4]
  assign _T_59002 = _T_59001[10:0]; // @[Modules.scala 68:83:@6459.4]
  assign buffer_2_637 = $signed(_T_59002); // @[Modules.scala 68:83:@6460.4]
  assign _T_59007 = $signed(buffer_2_494) + $signed(buffer_0_495); // @[Modules.scala 68:83:@6466.4]
  assign _T_59008 = _T_59007[10:0]; // @[Modules.scala 68:83:@6467.4]
  assign buffer_2_639 = $signed(_T_59008); // @[Modules.scala 68:83:@6468.4]
  assign _T_59010 = $signed(buffer_0_395) + $signed(buffer_2_497); // @[Modules.scala 68:83:@6470.4]
  assign _T_59011 = _T_59010[10:0]; // @[Modules.scala 68:83:@6471.4]
  assign buffer_2_640 = $signed(_T_59011); // @[Modules.scala 68:83:@6472.4]
  assign _T_59013 = $signed(buffer_2_498) + $signed(buffer_2_499); // @[Modules.scala 68:83:@6474.4]
  assign _T_59014 = _T_59013[10:0]; // @[Modules.scala 68:83:@6475.4]
  assign buffer_2_641 = $signed(_T_59014); // @[Modules.scala 68:83:@6476.4]
  assign _T_59016 = $signed(buffer_0_500) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6478.4]
  assign _T_59017 = _T_59016[10:0]; // @[Modules.scala 68:83:@6479.4]
  assign buffer_2_642 = $signed(_T_59017); // @[Modules.scala 68:83:@6480.4]
  assign _T_59019 = $signed(buffer_2_502) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6482.4]
  assign _T_59020 = _T_59019[10:0]; // @[Modules.scala 68:83:@6483.4]
  assign buffer_2_643 = $signed(_T_59020); // @[Modules.scala 68:83:@6484.4]
  assign _T_59022 = $signed(buffer_2_504) + $signed(buffer_2_505); // @[Modules.scala 68:83:@6486.4]
  assign _T_59023 = _T_59022[10:0]; // @[Modules.scala 68:83:@6487.4]
  assign buffer_2_644 = $signed(_T_59023); // @[Modules.scala 68:83:@6488.4]
  assign _T_59025 = $signed(buffer_2_506) + $signed(buffer_2_507); // @[Modules.scala 68:83:@6490.4]
  assign _T_59026 = _T_59025[10:0]; // @[Modules.scala 68:83:@6491.4]
  assign buffer_2_645 = $signed(_T_59026); // @[Modules.scala 68:83:@6492.4]
  assign _T_59028 = $signed(buffer_2_508) + $signed(buffer_2_509); // @[Modules.scala 68:83:@6494.4]
  assign _T_59029 = _T_59028[10:0]; // @[Modules.scala 68:83:@6495.4]
  assign buffer_2_646 = $signed(_T_59029); // @[Modules.scala 68:83:@6496.4]
  assign _T_59031 = $signed(buffer_0_395) + $signed(buffer_2_511); // @[Modules.scala 68:83:@6498.4]
  assign _T_59032 = _T_59031[10:0]; // @[Modules.scala 68:83:@6499.4]
  assign buffer_2_647 = $signed(_T_59032); // @[Modules.scala 68:83:@6500.4]
  assign _T_59034 = $signed(buffer_0_395) + $signed(buffer_2_513); // @[Modules.scala 68:83:@6502.4]
  assign _T_59035 = _T_59034[10:0]; // @[Modules.scala 68:83:@6503.4]
  assign buffer_2_648 = $signed(_T_59035); // @[Modules.scala 68:83:@6504.4]
  assign _T_59037 = $signed(buffer_2_514) + $signed(buffer_1_515); // @[Modules.scala 68:83:@6506.4]
  assign _T_59038 = _T_59037[10:0]; // @[Modules.scala 68:83:@6507.4]
  assign buffer_2_649 = $signed(_T_59038); // @[Modules.scala 68:83:@6508.4]
  assign _T_59040 = $signed(buffer_2_516) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6510.4]
  assign _T_59041 = _T_59040[10:0]; // @[Modules.scala 68:83:@6511.4]
  assign buffer_2_650 = $signed(_T_59041); // @[Modules.scala 68:83:@6512.4]
  assign _T_59046 = $signed(buffer_1_520) + $signed(buffer_2_521); // @[Modules.scala 68:83:@6518.4]
  assign _T_59047 = _T_59046[10:0]; // @[Modules.scala 68:83:@6519.4]
  assign buffer_2_652 = $signed(_T_59047); // @[Modules.scala 68:83:@6520.4]
  assign _T_59049 = $signed(buffer_2_522) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6522.4]
  assign _T_59050 = _T_59049[10:0]; // @[Modules.scala 68:83:@6523.4]
  assign buffer_2_653 = $signed(_T_59050); // @[Modules.scala 68:83:@6524.4]
  assign _T_59058 = $signed(buffer_2_528) + $signed(buffer_2_529); // @[Modules.scala 68:83:@6534.4]
  assign _T_59059 = _T_59058[10:0]; // @[Modules.scala 68:83:@6535.4]
  assign buffer_2_656 = $signed(_T_59059); // @[Modules.scala 68:83:@6536.4]
  assign _T_59061 = $signed(buffer_2_530) + $signed(buffer_2_531); // @[Modules.scala 68:83:@6538.4]
  assign _T_59062 = _T_59061[10:0]; // @[Modules.scala 68:83:@6539.4]
  assign buffer_2_657 = $signed(_T_59062); // @[Modules.scala 68:83:@6540.4]
  assign _T_59064 = $signed(buffer_2_532) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6542.4]
  assign _T_59065 = _T_59064[10:0]; // @[Modules.scala 68:83:@6543.4]
  assign buffer_2_658 = $signed(_T_59065); // @[Modules.scala 68:83:@6544.4]
  assign _T_59067 = $signed(buffer_0_534) + $signed(buffer_2_535); // @[Modules.scala 68:83:@6546.4]
  assign _T_59068 = _T_59067[10:0]; // @[Modules.scala 68:83:@6547.4]
  assign buffer_2_659 = $signed(_T_59068); // @[Modules.scala 68:83:@6548.4]
  assign _T_59070 = $signed(buffer_2_536) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6550.4]
  assign _T_59071 = _T_59070[10:0]; // @[Modules.scala 68:83:@6551.4]
  assign buffer_2_660 = $signed(_T_59071); // @[Modules.scala 68:83:@6552.4]
  assign _T_59073 = $signed(buffer_1_538) + $signed(buffer_2_539); // @[Modules.scala 68:83:@6554.4]
  assign _T_59074 = _T_59073[10:0]; // @[Modules.scala 68:83:@6555.4]
  assign buffer_2_661 = $signed(_T_59074); // @[Modules.scala 68:83:@6556.4]
  assign _T_59076 = $signed(buffer_2_540) + $signed(buffer_2_541); // @[Modules.scala 68:83:@6558.4]
  assign _T_59077 = _T_59076[10:0]; // @[Modules.scala 68:83:@6559.4]
  assign buffer_2_662 = $signed(_T_59077); // @[Modules.scala 68:83:@6560.4]
  assign _T_59079 = $signed(buffer_2_542) + $signed(buffer_2_543); // @[Modules.scala 68:83:@6562.4]
  assign _T_59080 = _T_59079[10:0]; // @[Modules.scala 68:83:@6563.4]
  assign buffer_2_663 = $signed(_T_59080); // @[Modules.scala 68:83:@6564.4]
  assign _T_59082 = $signed(buffer_2_544) + $signed(buffer_1_545); // @[Modules.scala 68:83:@6566.4]
  assign _T_59083 = _T_59082[10:0]; // @[Modules.scala 68:83:@6567.4]
  assign buffer_2_664 = $signed(_T_59083); // @[Modules.scala 68:83:@6568.4]
  assign _T_59085 = $signed(buffer_2_546) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6570.4]
  assign _T_59086 = _T_59085[10:0]; // @[Modules.scala 68:83:@6571.4]
  assign buffer_2_665 = $signed(_T_59086); // @[Modules.scala 68:83:@6572.4]
  assign _T_59088 = $signed(buffer_2_548) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6574.4]
  assign _T_59089 = _T_59088[10:0]; // @[Modules.scala 68:83:@6575.4]
  assign buffer_2_666 = $signed(_T_59089); // @[Modules.scala 68:83:@6576.4]
  assign _T_59091 = $signed(buffer_2_550) + $signed(buffer_1_551); // @[Modules.scala 68:83:@6578.4]
  assign _T_59092 = _T_59091[10:0]; // @[Modules.scala 68:83:@6579.4]
  assign buffer_2_667 = $signed(_T_59092); // @[Modules.scala 68:83:@6580.4]
  assign _T_59094 = $signed(buffer_1_552) + $signed(buffer_2_553); // @[Modules.scala 68:83:@6582.4]
  assign _T_59095 = _T_59094[10:0]; // @[Modules.scala 68:83:@6583.4]
  assign buffer_2_668 = $signed(_T_59095); // @[Modules.scala 68:83:@6584.4]
  assign _T_59097 = $signed(buffer_2_554) + $signed(buffer_2_555); // @[Modules.scala 68:83:@6586.4]
  assign _T_59098 = _T_59097[10:0]; // @[Modules.scala 68:83:@6587.4]
  assign buffer_2_669 = $signed(_T_59098); // @[Modules.scala 68:83:@6588.4]
  assign _T_59100 = $signed(buffer_2_556) + $signed(buffer_2_557); // @[Modules.scala 68:83:@6590.4]
  assign _T_59101 = _T_59100[10:0]; // @[Modules.scala 68:83:@6591.4]
  assign buffer_2_670 = $signed(_T_59101); // @[Modules.scala 68:83:@6592.4]
  assign _T_59103 = $signed(buffer_0_558) + $signed(buffer_2_559); // @[Modules.scala 68:83:@6594.4]
  assign _T_59104 = _T_59103[10:0]; // @[Modules.scala 68:83:@6595.4]
  assign buffer_2_671 = $signed(_T_59104); // @[Modules.scala 68:83:@6596.4]
  assign _T_59106 = $signed(buffer_2_560) + $signed(buffer_0_395); // @[Modules.scala 68:83:@6598.4]
  assign _T_59107 = _T_59106[10:0]; // @[Modules.scala 68:83:@6599.4]
  assign buffer_2_672 = $signed(_T_59107); // @[Modules.scala 68:83:@6600.4]
  assign _T_59109 = $signed(buffer_0_395) + $signed(buffer_2_563); // @[Modules.scala 68:83:@6602.4]
  assign _T_59110 = _T_59109[10:0]; // @[Modules.scala 68:83:@6603.4]
  assign buffer_2_673 = $signed(_T_59110); // @[Modules.scala 68:83:@6604.4]
  assign _T_59112 = $signed(buffer_2_564) + $signed(buffer_0_565); // @[Modules.scala 68:83:@6606.4]
  assign _T_59113 = _T_59112[10:0]; // @[Modules.scala 68:83:@6607.4]
  assign buffer_2_674 = $signed(_T_59113); // @[Modules.scala 68:83:@6608.4]
  assign _T_59115 = $signed(buffer_2_566) + $signed(buffer_2_567); // @[Modules.scala 68:83:@6610.4]
  assign _T_59116 = _T_59115[10:0]; // @[Modules.scala 68:83:@6611.4]
  assign buffer_2_675 = $signed(_T_59116); // @[Modules.scala 68:83:@6612.4]
  assign _T_59127 = $signed(buffer_2_574) + $signed(buffer_2_575); // @[Modules.scala 68:83:@6626.4]
  assign _T_59128 = _T_59127[10:0]; // @[Modules.scala 68:83:@6627.4]
  assign buffer_2_679 = $signed(_T_59128); // @[Modules.scala 68:83:@6628.4]
  assign _T_59133 = $signed(buffer_0_395) + $signed(buffer_2_579); // @[Modules.scala 68:83:@6634.4]
  assign _T_59134 = _T_59133[10:0]; // @[Modules.scala 68:83:@6635.4]
  assign buffer_2_681 = $signed(_T_59134); // @[Modules.scala 68:83:@6636.4]
  assign _T_59136 = $signed(buffer_2_580) + $signed(buffer_2_581); // @[Modules.scala 68:83:@6638.4]
  assign _T_59137 = _T_59136[10:0]; // @[Modules.scala 68:83:@6639.4]
  assign buffer_2_682 = $signed(_T_59137); // @[Modules.scala 68:83:@6640.4]
  assign _T_59145 = $signed(buffer_0_395) + $signed(buffer_2_587); // @[Modules.scala 68:83:@6650.4]
  assign _T_59146 = _T_59145[10:0]; // @[Modules.scala 68:83:@6651.4]
  assign buffer_2_685 = $signed(_T_59146); // @[Modules.scala 68:83:@6652.4]
  assign _T_59148 = $signed(buffer_2_588) + $signed(buffer_2_589); // @[Modules.scala 71:109:@6654.4]
  assign _T_59149 = _T_59148[10:0]; // @[Modules.scala 71:109:@6655.4]
  assign buffer_2_686 = $signed(_T_59149); // @[Modules.scala 71:109:@6656.4]
  assign _T_59151 = $signed(buffer_2_590) + $signed(buffer_2_591); // @[Modules.scala 71:109:@6658.4]
  assign _T_59152 = _T_59151[10:0]; // @[Modules.scala 71:109:@6659.4]
  assign buffer_2_687 = $signed(_T_59152); // @[Modules.scala 71:109:@6660.4]
  assign _T_59154 = $signed(buffer_2_592) + $signed(buffer_2_593); // @[Modules.scala 71:109:@6662.4]
  assign _T_59155 = _T_59154[10:0]; // @[Modules.scala 71:109:@6663.4]
  assign buffer_2_688 = $signed(_T_59155); // @[Modules.scala 71:109:@6664.4]
  assign _T_59157 = $signed(buffer_2_594) + $signed(buffer_2_595); // @[Modules.scala 71:109:@6666.4]
  assign _T_59158 = _T_59157[10:0]; // @[Modules.scala 71:109:@6667.4]
  assign buffer_2_689 = $signed(_T_59158); // @[Modules.scala 71:109:@6668.4]
  assign _T_59160 = $signed(buffer_2_596) + $signed(buffer_2_597); // @[Modules.scala 71:109:@6670.4]
  assign _T_59161 = _T_59160[10:0]; // @[Modules.scala 71:109:@6671.4]
  assign buffer_2_690 = $signed(_T_59161); // @[Modules.scala 71:109:@6672.4]
  assign _T_59163 = $signed(buffer_2_598) + $signed(buffer_2_599); // @[Modules.scala 71:109:@6674.4]
  assign _T_59164 = _T_59163[10:0]; // @[Modules.scala 71:109:@6675.4]
  assign buffer_2_691 = $signed(_T_59164); // @[Modules.scala 71:109:@6676.4]
  assign _T_59166 = $signed(buffer_2_600) + $signed(buffer_2_601); // @[Modules.scala 71:109:@6678.4]
  assign _T_59167 = _T_59166[10:0]; // @[Modules.scala 71:109:@6679.4]
  assign buffer_2_692 = $signed(_T_59167); // @[Modules.scala 71:109:@6680.4]
  assign _T_59169 = $signed(buffer_2_602) + $signed(buffer_0_593); // @[Modules.scala 71:109:@6682.4]
  assign _T_59170 = _T_59169[10:0]; // @[Modules.scala 71:109:@6683.4]
  assign buffer_2_693 = $signed(_T_59170); // @[Modules.scala 71:109:@6684.4]
  assign _T_59172 = $signed(buffer_2_604) + $signed(buffer_2_605); // @[Modules.scala 71:109:@6686.4]
  assign _T_59173 = _T_59172[10:0]; // @[Modules.scala 71:109:@6687.4]
  assign buffer_2_694 = $signed(_T_59173); // @[Modules.scala 71:109:@6688.4]
  assign _T_59175 = $signed(buffer_0_593) + $signed(buffer_2_607); // @[Modules.scala 71:109:@6690.4]
  assign _T_59176 = _T_59175[10:0]; // @[Modules.scala 71:109:@6691.4]
  assign buffer_2_695 = $signed(_T_59176); // @[Modules.scala 71:109:@6692.4]
  assign _T_59178 = $signed(buffer_2_608) + $signed(buffer_2_609); // @[Modules.scala 71:109:@6694.4]
  assign _T_59179 = _T_59178[10:0]; // @[Modules.scala 71:109:@6695.4]
  assign buffer_2_696 = $signed(_T_59179); // @[Modules.scala 71:109:@6696.4]
  assign _T_59181 = $signed(buffer_0_593) + $signed(buffer_2_611); // @[Modules.scala 71:109:@6698.4]
  assign _T_59182 = _T_59181[10:0]; // @[Modules.scala 71:109:@6699.4]
  assign buffer_2_697 = $signed(_T_59182); // @[Modules.scala 71:109:@6700.4]
  assign _T_59184 = $signed(buffer_2_612) + $signed(buffer_0_593); // @[Modules.scala 71:109:@6702.4]
  assign _T_59185 = _T_59184[10:0]; // @[Modules.scala 71:109:@6703.4]
  assign buffer_2_698 = $signed(_T_59185); // @[Modules.scala 71:109:@6704.4]
  assign _T_59187 = $signed(buffer_2_614) + $signed(buffer_2_615); // @[Modules.scala 71:109:@6706.4]
  assign _T_59188 = _T_59187[10:0]; // @[Modules.scala 71:109:@6707.4]
  assign buffer_2_699 = $signed(_T_59188); // @[Modules.scala 71:109:@6708.4]
  assign _T_59190 = $signed(buffer_0_593) + $signed(buffer_2_617); // @[Modules.scala 71:109:@6710.4]
  assign _T_59191 = _T_59190[10:0]; // @[Modules.scala 71:109:@6711.4]
  assign buffer_2_700 = $signed(_T_59191); // @[Modules.scala 71:109:@6712.4]
  assign _T_59193 = $signed(buffer_2_618) + $signed(buffer_2_619); // @[Modules.scala 71:109:@6714.4]
  assign _T_59194 = _T_59193[10:0]; // @[Modules.scala 71:109:@6715.4]
  assign buffer_2_701 = $signed(_T_59194); // @[Modules.scala 71:109:@6716.4]
  assign _T_59196 = $signed(buffer_2_620) + $signed(buffer_0_593); // @[Modules.scala 71:109:@6718.4]
  assign _T_59197 = _T_59196[10:0]; // @[Modules.scala 71:109:@6719.4]
  assign buffer_2_702 = $signed(_T_59197); // @[Modules.scala 71:109:@6720.4]
  assign _T_59199 = $signed(buffer_2_622) + $signed(buffer_2_623); // @[Modules.scala 71:109:@6722.4]
  assign _T_59200 = _T_59199[10:0]; // @[Modules.scala 71:109:@6723.4]
  assign buffer_2_703 = $signed(_T_59200); // @[Modules.scala 71:109:@6724.4]
  assign _T_59202 = $signed(buffer_2_624) + $signed(buffer_0_593); // @[Modules.scala 71:109:@6726.4]
  assign _T_59203 = _T_59202[10:0]; // @[Modules.scala 71:109:@6727.4]
  assign buffer_2_704 = $signed(_T_59203); // @[Modules.scala 71:109:@6728.4]
  assign _T_59205 = $signed(buffer_2_626) + $signed(buffer_2_627); // @[Modules.scala 71:109:@6730.4]
  assign _T_59206 = _T_59205[10:0]; // @[Modules.scala 71:109:@6731.4]
  assign buffer_2_705 = $signed(_T_59206); // @[Modules.scala 71:109:@6732.4]
  assign _T_59208 = $signed(buffer_2_628) + $signed(buffer_2_629); // @[Modules.scala 71:109:@6734.4]
  assign _T_59209 = _T_59208[10:0]; // @[Modules.scala 71:109:@6735.4]
  assign buffer_2_706 = $signed(_T_59209); // @[Modules.scala 71:109:@6736.4]
  assign _T_59214 = $signed(buffer_2_632) + $signed(buffer_2_633); // @[Modules.scala 71:109:@6742.4]
  assign _T_59215 = _T_59214[10:0]; // @[Modules.scala 71:109:@6743.4]
  assign buffer_2_708 = $signed(_T_59215); // @[Modules.scala 71:109:@6744.4]
  assign _T_59217 = $signed(buffer_1_634) + $signed(buffer_0_635); // @[Modules.scala 71:109:@6746.4]
  assign _T_59218 = _T_59217[10:0]; // @[Modules.scala 71:109:@6747.4]
  assign buffer_2_709 = $signed(_T_59218); // @[Modules.scala 71:109:@6748.4]
  assign _T_59220 = $signed(buffer_2_636) + $signed(buffer_2_637); // @[Modules.scala 71:109:@6750.4]
  assign _T_59221 = _T_59220[10:0]; // @[Modules.scala 71:109:@6751.4]
  assign buffer_2_710 = $signed(_T_59221); // @[Modules.scala 71:109:@6752.4]
  assign _T_59223 = $signed(buffer_0_638) + $signed(buffer_2_639); // @[Modules.scala 71:109:@6754.4]
  assign _T_59224 = _T_59223[10:0]; // @[Modules.scala 71:109:@6755.4]
  assign buffer_2_711 = $signed(_T_59224); // @[Modules.scala 71:109:@6756.4]
  assign _T_59226 = $signed(buffer_2_640) + $signed(buffer_2_641); // @[Modules.scala 71:109:@6758.4]
  assign _T_59227 = _T_59226[10:0]; // @[Modules.scala 71:109:@6759.4]
  assign buffer_2_712 = $signed(_T_59227); // @[Modules.scala 71:109:@6760.4]
  assign _T_59229 = $signed(buffer_2_642) + $signed(buffer_2_643); // @[Modules.scala 71:109:@6762.4]
  assign _T_59230 = _T_59229[10:0]; // @[Modules.scala 71:109:@6763.4]
  assign buffer_2_713 = $signed(_T_59230); // @[Modules.scala 71:109:@6764.4]
  assign _T_59232 = $signed(buffer_2_644) + $signed(buffer_2_645); // @[Modules.scala 71:109:@6766.4]
  assign _T_59233 = _T_59232[10:0]; // @[Modules.scala 71:109:@6767.4]
  assign buffer_2_714 = $signed(_T_59233); // @[Modules.scala 71:109:@6768.4]
  assign _T_59235 = $signed(buffer_2_646) + $signed(buffer_2_647); // @[Modules.scala 71:109:@6770.4]
  assign _T_59236 = _T_59235[10:0]; // @[Modules.scala 71:109:@6771.4]
  assign buffer_2_715 = $signed(_T_59236); // @[Modules.scala 71:109:@6772.4]
  assign _T_59238 = $signed(buffer_2_648) + $signed(buffer_2_649); // @[Modules.scala 71:109:@6774.4]
  assign _T_59239 = _T_59238[10:0]; // @[Modules.scala 71:109:@6775.4]
  assign buffer_2_716 = $signed(_T_59239); // @[Modules.scala 71:109:@6776.4]
  assign _T_59241 = $signed(buffer_2_650) + $signed(buffer_0_593); // @[Modules.scala 71:109:@6778.4]
  assign _T_59242 = _T_59241[10:0]; // @[Modules.scala 71:109:@6779.4]
  assign buffer_2_717 = $signed(_T_59242); // @[Modules.scala 71:109:@6780.4]
  assign _T_59244 = $signed(buffer_2_652) + $signed(buffer_2_653); // @[Modules.scala 71:109:@6782.4]
  assign _T_59245 = _T_59244[10:0]; // @[Modules.scala 71:109:@6783.4]
  assign buffer_2_718 = $signed(_T_59245); // @[Modules.scala 71:109:@6784.4]
  assign _T_59247 = $signed(buffer_0_593) + $signed(buffer_0_655); // @[Modules.scala 71:109:@6786.4]
  assign _T_59248 = _T_59247[10:0]; // @[Modules.scala 71:109:@6787.4]
  assign buffer_2_719 = $signed(_T_59248); // @[Modules.scala 71:109:@6788.4]
  assign _T_59250 = $signed(buffer_2_656) + $signed(buffer_2_657); // @[Modules.scala 71:109:@6790.4]
  assign _T_59251 = _T_59250[10:0]; // @[Modules.scala 71:109:@6791.4]
  assign buffer_2_720 = $signed(_T_59251); // @[Modules.scala 71:109:@6792.4]
  assign _T_59253 = $signed(buffer_2_658) + $signed(buffer_2_659); // @[Modules.scala 71:109:@6794.4]
  assign _T_59254 = _T_59253[10:0]; // @[Modules.scala 71:109:@6795.4]
  assign buffer_2_721 = $signed(_T_59254); // @[Modules.scala 71:109:@6796.4]
  assign _T_59256 = $signed(buffer_2_660) + $signed(buffer_2_661); // @[Modules.scala 71:109:@6798.4]
  assign _T_59257 = _T_59256[10:0]; // @[Modules.scala 71:109:@6799.4]
  assign buffer_2_722 = $signed(_T_59257); // @[Modules.scala 71:109:@6800.4]
  assign _T_59259 = $signed(buffer_2_662) + $signed(buffer_2_663); // @[Modules.scala 71:109:@6802.4]
  assign _T_59260 = _T_59259[10:0]; // @[Modules.scala 71:109:@6803.4]
  assign buffer_2_723 = $signed(_T_59260); // @[Modules.scala 71:109:@6804.4]
  assign _T_59262 = $signed(buffer_2_664) + $signed(buffer_2_665); // @[Modules.scala 71:109:@6806.4]
  assign _T_59263 = _T_59262[10:0]; // @[Modules.scala 71:109:@6807.4]
  assign buffer_2_724 = $signed(_T_59263); // @[Modules.scala 71:109:@6808.4]
  assign _T_59265 = $signed(buffer_2_666) + $signed(buffer_2_667); // @[Modules.scala 71:109:@6810.4]
  assign _T_59266 = _T_59265[10:0]; // @[Modules.scala 71:109:@6811.4]
  assign buffer_2_725 = $signed(_T_59266); // @[Modules.scala 71:109:@6812.4]
  assign _T_59268 = $signed(buffer_2_668) + $signed(buffer_2_669); // @[Modules.scala 71:109:@6814.4]
  assign _T_59269 = _T_59268[10:0]; // @[Modules.scala 71:109:@6815.4]
  assign buffer_2_726 = $signed(_T_59269); // @[Modules.scala 71:109:@6816.4]
  assign _T_59271 = $signed(buffer_2_670) + $signed(buffer_2_671); // @[Modules.scala 71:109:@6818.4]
  assign _T_59272 = _T_59271[10:0]; // @[Modules.scala 71:109:@6819.4]
  assign buffer_2_727 = $signed(_T_59272); // @[Modules.scala 71:109:@6820.4]
  assign _T_59274 = $signed(buffer_2_672) + $signed(buffer_2_673); // @[Modules.scala 71:109:@6822.4]
  assign _T_59275 = _T_59274[10:0]; // @[Modules.scala 71:109:@6823.4]
  assign buffer_2_728 = $signed(_T_59275); // @[Modules.scala 71:109:@6824.4]
  assign _T_59277 = $signed(buffer_2_674) + $signed(buffer_2_675); // @[Modules.scala 71:109:@6826.4]
  assign _T_59278 = _T_59277[10:0]; // @[Modules.scala 71:109:@6827.4]
  assign buffer_2_729 = $signed(_T_59278); // @[Modules.scala 71:109:@6828.4]
  assign _T_59283 = $signed(buffer_0_678) + $signed(buffer_2_679); // @[Modules.scala 71:109:@6834.4]
  assign _T_59284 = _T_59283[10:0]; // @[Modules.scala 71:109:@6835.4]
  assign buffer_2_731 = $signed(_T_59284); // @[Modules.scala 71:109:@6836.4]
  assign _T_59286 = $signed(buffer_0_593) + $signed(buffer_2_681); // @[Modules.scala 71:109:@6838.4]
  assign _T_59287 = _T_59286[10:0]; // @[Modules.scala 71:109:@6839.4]
  assign buffer_2_732 = $signed(_T_59287); // @[Modules.scala 71:109:@6840.4]
  assign _T_59289 = $signed(buffer_2_682) + $signed(buffer_0_683); // @[Modules.scala 71:109:@6842.4]
  assign _T_59290 = _T_59289[10:0]; // @[Modules.scala 71:109:@6843.4]
  assign buffer_2_733 = $signed(_T_59290); // @[Modules.scala 71:109:@6844.4]
  assign _T_59292 = $signed(buffer_0_593) + $signed(buffer_2_685); // @[Modules.scala 71:109:@6846.4]
  assign _T_59293 = _T_59292[10:0]; // @[Modules.scala 71:109:@6847.4]
  assign buffer_2_734 = $signed(_T_59293); // @[Modules.scala 71:109:@6848.4]
  assign _T_59295 = $signed(buffer_2_686) + $signed(buffer_2_687); // @[Modules.scala 78:156:@6851.4]
  assign _T_59296 = _T_59295[10:0]; // @[Modules.scala 78:156:@6852.4]
  assign buffer_2_736 = $signed(_T_59296); // @[Modules.scala 78:156:@6853.4]
  assign _T_59298 = $signed(buffer_2_736) + $signed(buffer_2_688); // @[Modules.scala 78:156:@6855.4]
  assign _T_59299 = _T_59298[10:0]; // @[Modules.scala 78:156:@6856.4]
  assign buffer_2_737 = $signed(_T_59299); // @[Modules.scala 78:156:@6857.4]
  assign _T_59301 = $signed(buffer_2_737) + $signed(buffer_2_689); // @[Modules.scala 78:156:@6859.4]
  assign _T_59302 = _T_59301[10:0]; // @[Modules.scala 78:156:@6860.4]
  assign buffer_2_738 = $signed(_T_59302); // @[Modules.scala 78:156:@6861.4]
  assign _T_59304 = $signed(buffer_2_738) + $signed(buffer_2_690); // @[Modules.scala 78:156:@6863.4]
  assign _T_59305 = _T_59304[10:0]; // @[Modules.scala 78:156:@6864.4]
  assign buffer_2_739 = $signed(_T_59305); // @[Modules.scala 78:156:@6865.4]
  assign _T_59307 = $signed(buffer_2_739) + $signed(buffer_2_691); // @[Modules.scala 78:156:@6867.4]
  assign _T_59308 = _T_59307[10:0]; // @[Modules.scala 78:156:@6868.4]
  assign buffer_2_740 = $signed(_T_59308); // @[Modules.scala 78:156:@6869.4]
  assign _T_59310 = $signed(buffer_2_740) + $signed(buffer_2_692); // @[Modules.scala 78:156:@6871.4]
  assign _T_59311 = _T_59310[10:0]; // @[Modules.scala 78:156:@6872.4]
  assign buffer_2_741 = $signed(_T_59311); // @[Modules.scala 78:156:@6873.4]
  assign _T_59313 = $signed(buffer_2_741) + $signed(buffer_2_693); // @[Modules.scala 78:156:@6875.4]
  assign _T_59314 = _T_59313[10:0]; // @[Modules.scala 78:156:@6876.4]
  assign buffer_2_742 = $signed(_T_59314); // @[Modules.scala 78:156:@6877.4]
  assign _T_59316 = $signed(buffer_2_742) + $signed(buffer_2_694); // @[Modules.scala 78:156:@6879.4]
  assign _T_59317 = _T_59316[10:0]; // @[Modules.scala 78:156:@6880.4]
  assign buffer_2_743 = $signed(_T_59317); // @[Modules.scala 78:156:@6881.4]
  assign _T_59319 = $signed(buffer_2_743) + $signed(buffer_2_695); // @[Modules.scala 78:156:@6883.4]
  assign _T_59320 = _T_59319[10:0]; // @[Modules.scala 78:156:@6884.4]
  assign buffer_2_744 = $signed(_T_59320); // @[Modules.scala 78:156:@6885.4]
  assign _T_59322 = $signed(buffer_2_744) + $signed(buffer_2_696); // @[Modules.scala 78:156:@6887.4]
  assign _T_59323 = _T_59322[10:0]; // @[Modules.scala 78:156:@6888.4]
  assign buffer_2_745 = $signed(_T_59323); // @[Modules.scala 78:156:@6889.4]
  assign _T_59325 = $signed(buffer_2_745) + $signed(buffer_2_697); // @[Modules.scala 78:156:@6891.4]
  assign _T_59326 = _T_59325[10:0]; // @[Modules.scala 78:156:@6892.4]
  assign buffer_2_746 = $signed(_T_59326); // @[Modules.scala 78:156:@6893.4]
  assign _T_59328 = $signed(buffer_2_746) + $signed(buffer_2_698); // @[Modules.scala 78:156:@6895.4]
  assign _T_59329 = _T_59328[10:0]; // @[Modules.scala 78:156:@6896.4]
  assign buffer_2_747 = $signed(_T_59329); // @[Modules.scala 78:156:@6897.4]
  assign _T_59331 = $signed(buffer_2_747) + $signed(buffer_2_699); // @[Modules.scala 78:156:@6899.4]
  assign _T_59332 = _T_59331[10:0]; // @[Modules.scala 78:156:@6900.4]
  assign buffer_2_748 = $signed(_T_59332); // @[Modules.scala 78:156:@6901.4]
  assign _T_59334 = $signed(buffer_2_748) + $signed(buffer_2_700); // @[Modules.scala 78:156:@6903.4]
  assign _T_59335 = _T_59334[10:0]; // @[Modules.scala 78:156:@6904.4]
  assign buffer_2_749 = $signed(_T_59335); // @[Modules.scala 78:156:@6905.4]
  assign _T_59337 = $signed(buffer_2_749) + $signed(buffer_2_701); // @[Modules.scala 78:156:@6907.4]
  assign _T_59338 = _T_59337[10:0]; // @[Modules.scala 78:156:@6908.4]
  assign buffer_2_750 = $signed(_T_59338); // @[Modules.scala 78:156:@6909.4]
  assign _T_59340 = $signed(buffer_2_750) + $signed(buffer_2_702); // @[Modules.scala 78:156:@6911.4]
  assign _T_59341 = _T_59340[10:0]; // @[Modules.scala 78:156:@6912.4]
  assign buffer_2_751 = $signed(_T_59341); // @[Modules.scala 78:156:@6913.4]
  assign _T_59343 = $signed(buffer_2_751) + $signed(buffer_2_703); // @[Modules.scala 78:156:@6915.4]
  assign _T_59344 = _T_59343[10:0]; // @[Modules.scala 78:156:@6916.4]
  assign buffer_2_752 = $signed(_T_59344); // @[Modules.scala 78:156:@6917.4]
  assign _T_59346 = $signed(buffer_2_752) + $signed(buffer_2_704); // @[Modules.scala 78:156:@6919.4]
  assign _T_59347 = _T_59346[10:0]; // @[Modules.scala 78:156:@6920.4]
  assign buffer_2_753 = $signed(_T_59347); // @[Modules.scala 78:156:@6921.4]
  assign _T_59349 = $signed(buffer_2_753) + $signed(buffer_2_705); // @[Modules.scala 78:156:@6923.4]
  assign _T_59350 = _T_59349[10:0]; // @[Modules.scala 78:156:@6924.4]
  assign buffer_2_754 = $signed(_T_59350); // @[Modules.scala 78:156:@6925.4]
  assign _T_59352 = $signed(buffer_2_754) + $signed(buffer_2_706); // @[Modules.scala 78:156:@6927.4]
  assign _T_59353 = _T_59352[10:0]; // @[Modules.scala 78:156:@6928.4]
  assign buffer_2_755 = $signed(_T_59353); // @[Modules.scala 78:156:@6929.4]
  assign _T_59355 = $signed(buffer_2_755) + $signed(buffer_0_707); // @[Modules.scala 78:156:@6931.4]
  assign _T_59356 = _T_59355[10:0]; // @[Modules.scala 78:156:@6932.4]
  assign buffer_2_756 = $signed(_T_59356); // @[Modules.scala 78:156:@6933.4]
  assign _T_59358 = $signed(buffer_2_756) + $signed(buffer_2_708); // @[Modules.scala 78:156:@6935.4]
  assign _T_59359 = _T_59358[10:0]; // @[Modules.scala 78:156:@6936.4]
  assign buffer_2_757 = $signed(_T_59359); // @[Modules.scala 78:156:@6937.4]
  assign _T_59361 = $signed(buffer_2_757) + $signed(buffer_2_709); // @[Modules.scala 78:156:@6939.4]
  assign _T_59362 = _T_59361[10:0]; // @[Modules.scala 78:156:@6940.4]
  assign buffer_2_758 = $signed(_T_59362); // @[Modules.scala 78:156:@6941.4]
  assign _T_59364 = $signed(buffer_2_758) + $signed(buffer_2_710); // @[Modules.scala 78:156:@6943.4]
  assign _T_59365 = _T_59364[10:0]; // @[Modules.scala 78:156:@6944.4]
  assign buffer_2_759 = $signed(_T_59365); // @[Modules.scala 78:156:@6945.4]
  assign _T_59367 = $signed(buffer_2_759) + $signed(buffer_2_711); // @[Modules.scala 78:156:@6947.4]
  assign _T_59368 = _T_59367[10:0]; // @[Modules.scala 78:156:@6948.4]
  assign buffer_2_760 = $signed(_T_59368); // @[Modules.scala 78:156:@6949.4]
  assign _T_59370 = $signed(buffer_2_760) + $signed(buffer_2_712); // @[Modules.scala 78:156:@6951.4]
  assign _T_59371 = _T_59370[10:0]; // @[Modules.scala 78:156:@6952.4]
  assign buffer_2_761 = $signed(_T_59371); // @[Modules.scala 78:156:@6953.4]
  assign _T_59373 = $signed(buffer_2_761) + $signed(buffer_2_713); // @[Modules.scala 78:156:@6955.4]
  assign _T_59374 = _T_59373[10:0]; // @[Modules.scala 78:156:@6956.4]
  assign buffer_2_762 = $signed(_T_59374); // @[Modules.scala 78:156:@6957.4]
  assign _T_59376 = $signed(buffer_2_762) + $signed(buffer_2_714); // @[Modules.scala 78:156:@6959.4]
  assign _T_59377 = _T_59376[10:0]; // @[Modules.scala 78:156:@6960.4]
  assign buffer_2_763 = $signed(_T_59377); // @[Modules.scala 78:156:@6961.4]
  assign _T_59379 = $signed(buffer_2_763) + $signed(buffer_2_715); // @[Modules.scala 78:156:@6963.4]
  assign _T_59380 = _T_59379[10:0]; // @[Modules.scala 78:156:@6964.4]
  assign buffer_2_764 = $signed(_T_59380); // @[Modules.scala 78:156:@6965.4]
  assign _T_59382 = $signed(buffer_2_764) + $signed(buffer_2_716); // @[Modules.scala 78:156:@6967.4]
  assign _T_59383 = _T_59382[10:0]; // @[Modules.scala 78:156:@6968.4]
  assign buffer_2_765 = $signed(_T_59383); // @[Modules.scala 78:156:@6969.4]
  assign _T_59385 = $signed(buffer_2_765) + $signed(buffer_2_717); // @[Modules.scala 78:156:@6971.4]
  assign _T_59386 = _T_59385[10:0]; // @[Modules.scala 78:156:@6972.4]
  assign buffer_2_766 = $signed(_T_59386); // @[Modules.scala 78:156:@6973.4]
  assign _T_59388 = $signed(buffer_2_766) + $signed(buffer_2_718); // @[Modules.scala 78:156:@6975.4]
  assign _T_59389 = _T_59388[10:0]; // @[Modules.scala 78:156:@6976.4]
  assign buffer_2_767 = $signed(_T_59389); // @[Modules.scala 78:156:@6977.4]
  assign _T_59391 = $signed(buffer_2_767) + $signed(buffer_2_719); // @[Modules.scala 78:156:@6979.4]
  assign _T_59392 = _T_59391[10:0]; // @[Modules.scala 78:156:@6980.4]
  assign buffer_2_768 = $signed(_T_59392); // @[Modules.scala 78:156:@6981.4]
  assign _T_59394 = $signed(buffer_2_768) + $signed(buffer_2_720); // @[Modules.scala 78:156:@6983.4]
  assign _T_59395 = _T_59394[10:0]; // @[Modules.scala 78:156:@6984.4]
  assign buffer_2_769 = $signed(_T_59395); // @[Modules.scala 78:156:@6985.4]
  assign _T_59397 = $signed(buffer_2_769) + $signed(buffer_2_721); // @[Modules.scala 78:156:@6987.4]
  assign _T_59398 = _T_59397[10:0]; // @[Modules.scala 78:156:@6988.4]
  assign buffer_2_770 = $signed(_T_59398); // @[Modules.scala 78:156:@6989.4]
  assign _T_59400 = $signed(buffer_2_770) + $signed(buffer_2_722); // @[Modules.scala 78:156:@6991.4]
  assign _T_59401 = _T_59400[10:0]; // @[Modules.scala 78:156:@6992.4]
  assign buffer_2_771 = $signed(_T_59401); // @[Modules.scala 78:156:@6993.4]
  assign _T_59403 = $signed(buffer_2_771) + $signed(buffer_2_723); // @[Modules.scala 78:156:@6995.4]
  assign _T_59404 = _T_59403[10:0]; // @[Modules.scala 78:156:@6996.4]
  assign buffer_2_772 = $signed(_T_59404); // @[Modules.scala 78:156:@6997.4]
  assign _T_59406 = $signed(buffer_2_772) + $signed(buffer_2_724); // @[Modules.scala 78:156:@6999.4]
  assign _T_59407 = _T_59406[10:0]; // @[Modules.scala 78:156:@7000.4]
  assign buffer_2_773 = $signed(_T_59407); // @[Modules.scala 78:156:@7001.4]
  assign _T_59409 = $signed(buffer_2_773) + $signed(buffer_2_725); // @[Modules.scala 78:156:@7003.4]
  assign _T_59410 = _T_59409[10:0]; // @[Modules.scala 78:156:@7004.4]
  assign buffer_2_774 = $signed(_T_59410); // @[Modules.scala 78:156:@7005.4]
  assign _T_59412 = $signed(buffer_2_774) + $signed(buffer_2_726); // @[Modules.scala 78:156:@7007.4]
  assign _T_59413 = _T_59412[10:0]; // @[Modules.scala 78:156:@7008.4]
  assign buffer_2_775 = $signed(_T_59413); // @[Modules.scala 78:156:@7009.4]
  assign _T_59415 = $signed(buffer_2_775) + $signed(buffer_2_727); // @[Modules.scala 78:156:@7011.4]
  assign _T_59416 = _T_59415[10:0]; // @[Modules.scala 78:156:@7012.4]
  assign buffer_2_776 = $signed(_T_59416); // @[Modules.scala 78:156:@7013.4]
  assign _T_59418 = $signed(buffer_2_776) + $signed(buffer_2_728); // @[Modules.scala 78:156:@7015.4]
  assign _T_59419 = _T_59418[10:0]; // @[Modules.scala 78:156:@7016.4]
  assign buffer_2_777 = $signed(_T_59419); // @[Modules.scala 78:156:@7017.4]
  assign _T_59421 = $signed(buffer_2_777) + $signed(buffer_2_729); // @[Modules.scala 78:156:@7019.4]
  assign _T_59422 = _T_59421[10:0]; // @[Modules.scala 78:156:@7020.4]
  assign buffer_2_778 = $signed(_T_59422); // @[Modules.scala 78:156:@7021.4]
  assign _T_59424 = $signed(buffer_2_778) + $signed(buffer_0_701); // @[Modules.scala 78:156:@7023.4]
  assign _T_59425 = _T_59424[10:0]; // @[Modules.scala 78:156:@7024.4]
  assign buffer_2_779 = $signed(_T_59425); // @[Modules.scala 78:156:@7025.4]
  assign _T_59427 = $signed(buffer_2_779) + $signed(buffer_2_731); // @[Modules.scala 78:156:@7027.4]
  assign _T_59428 = _T_59427[10:0]; // @[Modules.scala 78:156:@7028.4]
  assign buffer_2_780 = $signed(_T_59428); // @[Modules.scala 78:156:@7029.4]
  assign _T_59430 = $signed(buffer_2_780) + $signed(buffer_2_732); // @[Modules.scala 78:156:@7031.4]
  assign _T_59431 = _T_59430[10:0]; // @[Modules.scala 78:156:@7032.4]
  assign buffer_2_781 = $signed(_T_59431); // @[Modules.scala 78:156:@7033.4]
  assign _T_59433 = $signed(buffer_2_781) + $signed(buffer_2_733); // @[Modules.scala 78:156:@7035.4]
  assign _T_59434 = _T_59433[10:0]; // @[Modules.scala 78:156:@7036.4]
  assign buffer_2_782 = $signed(_T_59434); // @[Modules.scala 78:156:@7037.4]
  assign _T_59436 = $signed(buffer_2_782) + $signed(buffer_2_734); // @[Modules.scala 78:156:@7039.4]
  assign _T_59437 = _T_59436[10:0]; // @[Modules.scala 78:156:@7040.4]
  assign buffer_2_783 = $signed(_T_59437); // @[Modules.scala 78:156:@7041.4]
  assign _T_59453 = $signed(io_in_26) + $signed(io_in_27); // @[Modules.scala 37:46:@7069.4]
  assign _T_59454 = _T_59453[4:0]; // @[Modules.scala 37:46:@7070.4]
  assign _T_59455 = $signed(_T_59454); // @[Modules.scala 37:46:@7071.4]
  assign _T_59456 = $signed(io_in_28) + $signed(io_in_29); // @[Modules.scala 37:46:@7073.4]
  assign _T_59457 = _T_59456[4:0]; // @[Modules.scala 37:46:@7074.4]
  assign _T_59458 = $signed(_T_59457); // @[Modules.scala 37:46:@7075.4]
  assign _T_59506 = $signed(io_in_114) + $signed(io_in_115); // @[Modules.scala 37:46:@7143.4]
  assign _T_59507 = _T_59506[4:0]; // @[Modules.scala 37:46:@7144.4]
  assign _T_59508 = $signed(_T_59507); // @[Modules.scala 37:46:@7145.4]
  assign _T_59513 = $signed(io_in_120) + $signed(io_in_121); // @[Modules.scala 37:46:@7152.4]
  assign _T_59514 = _T_59513[4:0]; // @[Modules.scala 37:46:@7153.4]
  assign _T_59515 = $signed(_T_59514); // @[Modules.scala 37:46:@7154.4]
  assign _T_59516 = $signed(io_in_122) + $signed(io_in_123); // @[Modules.scala 37:46:@7156.4]
  assign _T_59517 = _T_59516[4:0]; // @[Modules.scala 37:46:@7157.4]
  assign _T_59518 = $signed(_T_59517); // @[Modules.scala 37:46:@7158.4]
  assign _T_59519 = $signed(io_in_124) + $signed(io_in_125); // @[Modules.scala 37:46:@7160.4]
  assign _T_59520 = _T_59519[4:0]; // @[Modules.scala 37:46:@7161.4]
  assign _T_59521 = $signed(_T_59520); // @[Modules.scala 37:46:@7162.4]
  assign _T_59522 = $signed(io_in_126) + $signed(io_in_127); // @[Modules.scala 37:46:@7164.4]
  assign _T_59523 = _T_59522[4:0]; // @[Modules.scala 37:46:@7165.4]
  assign _T_59524 = $signed(_T_59523); // @[Modules.scala 37:46:@7166.4]
  assign _T_59544 = $signed(io_in_150) + $signed(io_in_151); // @[Modules.scala 37:46:@7197.4]
  assign _T_59545 = _T_59544[4:0]; // @[Modules.scala 37:46:@7198.4]
  assign _T_59546 = $signed(_T_59545); // @[Modules.scala 37:46:@7199.4]
  assign _T_59547 = $signed(io_in_154) + $signed(io_in_155); // @[Modules.scala 37:46:@7202.4]
  assign _T_59548 = _T_59547[4:0]; // @[Modules.scala 37:46:@7203.4]
  assign _T_59549 = $signed(_T_59548); // @[Modules.scala 37:46:@7204.4]
  assign _T_59550 = $signed(io_in_158) + $signed(io_in_159); // @[Modules.scala 37:46:@7207.4]
  assign _T_59551 = _T_59550[4:0]; // @[Modules.scala 37:46:@7208.4]
  assign _T_59552 = $signed(_T_59551); // @[Modules.scala 37:46:@7209.4]
  assign _T_59568 = $signed(io_in_172) + $signed(io_in_173); // @[Modules.scala 37:46:@7232.4]
  assign _T_59569 = _T_59568[4:0]; // @[Modules.scala 37:46:@7233.4]
  assign _T_59570 = $signed(_T_59569); // @[Modules.scala 37:46:@7234.4]
  assign _T_59577 = $signed(io_in_178) + $signed(io_in_179); // @[Modules.scala 37:46:@7244.4]
  assign _T_59578 = _T_59577[4:0]; // @[Modules.scala 37:46:@7245.4]
  assign _T_59579 = $signed(_T_59578); // @[Modules.scala 37:46:@7246.4]
  assign _T_59580 = $signed(io_in_180) + $signed(io_in_181); // @[Modules.scala 37:46:@7248.4]
  assign _T_59581 = _T_59580[4:0]; // @[Modules.scala 37:46:@7249.4]
  assign _T_59582 = $signed(_T_59581); // @[Modules.scala 37:46:@7250.4]
  assign _T_59590 = $signed(io_in_198) + $signed(io_in_199); // @[Modules.scala 37:46:@7266.4]
  assign _T_59591 = _T_59590[4:0]; // @[Modules.scala 37:46:@7267.4]
  assign _T_59592 = $signed(_T_59591); // @[Modules.scala 37:46:@7268.4]
  assign _T_59593 = $signed(io_in_200) + $signed(io_in_201); // @[Modules.scala 37:46:@7270.4]
  assign _T_59594 = _T_59593[4:0]; // @[Modules.scala 37:46:@7271.4]
  assign _T_59595 = $signed(_T_59594); // @[Modules.scala 37:46:@7272.4]
  assign _T_59599 = $signed(io_in_206) + $signed(io_in_207); // @[Modules.scala 37:46:@7279.4]
  assign _T_59600 = _T_59599[4:0]; // @[Modules.scala 37:46:@7280.4]
  assign _T_59601 = $signed(_T_59600); // @[Modules.scala 37:46:@7281.4]
  assign _T_59602 = $signed(io_in_208) + $signed(io_in_209); // @[Modules.scala 37:46:@7283.4]
  assign _T_59603 = _T_59602[4:0]; // @[Modules.scala 37:46:@7284.4]
  assign _T_59604 = $signed(_T_59603); // @[Modules.scala 37:46:@7285.4]
  assign _T_59605 = $signed(io_in_212) + $signed(io_in_213); // @[Modules.scala 37:46:@7288.4]
  assign _T_59606 = _T_59605[4:0]; // @[Modules.scala 37:46:@7289.4]
  assign _T_59607 = $signed(_T_59606); // @[Modules.scala 37:46:@7290.4]
  assign _T_59620 = $signed(io_in_226) + $signed(io_in_227); // @[Modules.scala 37:46:@7310.4]
  assign _T_59621 = _T_59620[4:0]; // @[Modules.scala 37:46:@7311.4]
  assign _T_59622 = $signed(_T_59621); // @[Modules.scala 37:46:@7312.4]
  assign _T_59623 = $signed(io_in_228) + $signed(io_in_229); // @[Modules.scala 37:46:@7314.4]
  assign _T_59624 = _T_59623[4:0]; // @[Modules.scala 37:46:@7315.4]
  assign _T_59625 = $signed(_T_59624); // @[Modules.scala 37:46:@7316.4]
  assign _T_59626 = $signed(io_in_234) + $signed(io_in_235); // @[Modules.scala 37:46:@7320.4]
  assign _T_59627 = _T_59626[4:0]; // @[Modules.scala 37:46:@7321.4]
  assign _T_59628 = $signed(_T_59627); // @[Modules.scala 37:46:@7322.4]
  assign _T_59629 = $signed(io_in_236) + $signed(io_in_237); // @[Modules.scala 37:46:@7324.4]
  assign _T_59630 = _T_59629[4:0]; // @[Modules.scala 37:46:@7325.4]
  assign _T_59631 = $signed(_T_59630); // @[Modules.scala 37:46:@7326.4]
  assign _T_59632 = $signed(io_in_238) + $signed(io_in_239); // @[Modules.scala 37:46:@7328.4]
  assign _T_59633 = _T_59632[4:0]; // @[Modules.scala 37:46:@7329.4]
  assign _T_59634 = $signed(_T_59633); // @[Modules.scala 37:46:@7330.4]
  assign _T_59638 = $signed(io_in_242) + $signed(io_in_243); // @[Modules.scala 37:46:@7336.4]
  assign _T_59639 = _T_59638[4:0]; // @[Modules.scala 37:46:@7337.4]
  assign _T_59640 = $signed(_T_59639); // @[Modules.scala 37:46:@7338.4]
  assign _T_59641 = $signed(io_in_246) + $signed(io_in_247); // @[Modules.scala 37:46:@7341.4]
  assign _T_59642 = _T_59641[4:0]; // @[Modules.scala 37:46:@7342.4]
  assign _T_59643 = $signed(_T_59642); // @[Modules.scala 37:46:@7343.4]
  assign _T_59650 = $signed(io_in_252) + $signed(io_in_253); // @[Modules.scala 37:46:@7353.4]
  assign _T_59651 = _T_59650[4:0]; // @[Modules.scala 37:46:@7354.4]
  assign _T_59652 = $signed(_T_59651); // @[Modules.scala 37:46:@7355.4]
  assign _T_59653 = $signed(io_in_254) + $signed(io_in_255); // @[Modules.scala 37:46:@7357.4]
  assign _T_59654 = _T_59653[4:0]; // @[Modules.scala 37:46:@7358.4]
  assign _T_59655 = $signed(_T_59654); // @[Modules.scala 37:46:@7359.4]
  assign _T_59656 = $signed(io_in_256) + $signed(io_in_257); // @[Modules.scala 37:46:@7361.4]
  assign _T_59657 = _T_59656[4:0]; // @[Modules.scala 37:46:@7362.4]
  assign _T_59658 = $signed(_T_59657); // @[Modules.scala 37:46:@7363.4]
  assign _T_59660 = $signed(io_in_264) + $signed(io_in_265); // @[Modules.scala 37:46:@7368.4]
  assign _T_59661 = _T_59660[4:0]; // @[Modules.scala 37:46:@7369.4]
  assign _T_59662 = $signed(_T_59661); // @[Modules.scala 37:46:@7370.4]
  assign _T_59666 = $signed(io_in_268) + $signed(io_in_269); // @[Modules.scala 37:46:@7376.4]
  assign _T_59667 = _T_59666[4:0]; // @[Modules.scala 37:46:@7377.4]
  assign _T_59668 = $signed(_T_59667); // @[Modules.scala 37:46:@7378.4]
  assign _T_59669 = $signed(io_in_270) + $signed(io_in_271); // @[Modules.scala 37:46:@7380.4]
  assign _T_59670 = _T_59669[4:0]; // @[Modules.scala 37:46:@7381.4]
  assign _T_59671 = $signed(_T_59670); // @[Modules.scala 37:46:@7382.4]
  assign _T_59672 = $signed(io_in_272) + $signed(io_in_273); // @[Modules.scala 37:46:@7384.4]
  assign _T_59673 = _T_59672[4:0]; // @[Modules.scala 37:46:@7385.4]
  assign _T_59674 = $signed(_T_59673); // @[Modules.scala 37:46:@7386.4]
  assign _T_59675 = $signed(io_in_274) + $signed(io_in_275); // @[Modules.scala 37:46:@7388.4]
  assign _T_59676 = _T_59675[4:0]; // @[Modules.scala 37:46:@7389.4]
  assign _T_59677 = $signed(_T_59676); // @[Modules.scala 37:46:@7390.4]
  assign _T_59684 = $signed(io_in_280) + $signed(io_in_281); // @[Modules.scala 37:46:@7400.4]
  assign _T_59685 = _T_59684[4:0]; // @[Modules.scala 37:46:@7401.4]
  assign _T_59686 = $signed(_T_59685); // @[Modules.scala 37:46:@7402.4]
  assign _T_59687 = $signed(io_in_282) + $signed(io_in_283); // @[Modules.scala 37:46:@7404.4]
  assign _T_59688 = _T_59687[4:0]; // @[Modules.scala 37:46:@7405.4]
  assign _T_59689 = $signed(_T_59688); // @[Modules.scala 37:46:@7406.4]
  assign _T_59694 = $signed(io_in_296) + $signed(io_in_297); // @[Modules.scala 37:46:@7414.4]
  assign _T_59695 = _T_59694[4:0]; // @[Modules.scala 37:46:@7415.4]
  assign _T_59696 = $signed(_T_59695); // @[Modules.scala 37:46:@7416.4]
  assign _T_59704 = $signed(io_in_310) + $signed(io_in_311); // @[Modules.scala 37:46:@7430.4]
  assign _T_59705 = _T_59704[4:0]; // @[Modules.scala 37:46:@7431.4]
  assign _T_59706 = $signed(_T_59705); // @[Modules.scala 37:46:@7432.4]
  assign _T_59738 = $signed(io_in_390) + $signed(io_in_391); // @[Modules.scala 37:46:@7473.4]
  assign _T_59739 = _T_59738[4:0]; // @[Modules.scala 37:46:@7474.4]
  assign _T_59740 = $signed(_T_59739); // @[Modules.scala 37:46:@7475.4]
  assign _T_59751 = $signed(io_in_418) + $signed(io_in_419); // @[Modules.scala 37:46:@7493.4]
  assign _T_59752 = _T_59751[4:0]; // @[Modules.scala 37:46:@7494.4]
  assign _T_59753 = $signed(_T_59752); // @[Modules.scala 37:46:@7495.4]
  assign _T_59757 = $signed(io_in_424) + $signed(io_in_425); // @[Modules.scala 37:46:@7502.4]
  assign _T_59758 = _T_59757[4:0]; // @[Modules.scala 37:46:@7503.4]
  assign _T_59759 = $signed(_T_59758); // @[Modules.scala 37:46:@7504.4]
  assign _T_59769 = $signed(io_in_444) + $signed(io_in_445); // @[Modules.scala 37:46:@7518.4]
  assign _T_59770 = _T_59769[4:0]; // @[Modules.scala 37:46:@7519.4]
  assign _T_59771 = $signed(_T_59770); // @[Modules.scala 37:46:@7520.4]
  assign _T_59772 = $signed(io_in_446) + $signed(io_in_447); // @[Modules.scala 37:46:@7522.4]
  assign _T_59773 = _T_59772[4:0]; // @[Modules.scala 37:46:@7523.4]
  assign _T_59774 = $signed(_T_59773); // @[Modules.scala 37:46:@7524.4]
  assign _T_59778 = $signed(io_in_452) + $signed(io_in_453); // @[Modules.scala 37:46:@7531.4]
  assign _T_59779 = _T_59778[4:0]; // @[Modules.scala 37:46:@7532.4]
  assign _T_59780 = $signed(_T_59779); // @[Modules.scala 37:46:@7533.4]
  assign _T_59798 = $signed(io_in_472) + $signed(io_in_473); // @[Modules.scala 37:46:@7556.4]
  assign _T_59799 = _T_59798[4:0]; // @[Modules.scala 37:46:@7557.4]
  assign _T_59800 = $signed(_T_59799); // @[Modules.scala 37:46:@7558.4]
  assign _T_59801 = $signed(io_in_474) + $signed(io_in_475); // @[Modules.scala 37:46:@7560.4]
  assign _T_59802 = _T_59801[4:0]; // @[Modules.scala 37:46:@7561.4]
  assign _T_59803 = $signed(_T_59802); // @[Modules.scala 37:46:@7562.4]
  assign _T_59808 = $signed(io_in_480) + $signed(io_in_481); // @[Modules.scala 37:46:@7569.4]
  assign _T_59809 = _T_59808[4:0]; // @[Modules.scala 37:46:@7570.4]
  assign _T_59810 = $signed(_T_59809); // @[Modules.scala 37:46:@7571.4]
  assign _T_59824 = $signed(io_in_500) + $signed(io_in_501); // @[Modules.scala 37:46:@7591.4]
  assign _T_59825 = _T_59824[4:0]; // @[Modules.scala 37:46:@7592.4]
  assign _T_59826 = $signed(_T_59825); // @[Modules.scala 37:46:@7593.4]
  assign _T_59827 = $signed(io_in_502) + $signed(io_in_503); // @[Modules.scala 37:46:@7595.4]
  assign _T_59828 = _T_59827[4:0]; // @[Modules.scala 37:46:@7596.4]
  assign _T_59829 = $signed(_T_59828); // @[Modules.scala 37:46:@7597.4]
  assign _T_59833 = $signed(io_in_508) + $signed(io_in_509); // @[Modules.scala 37:46:@7604.4]
  assign _T_59834 = _T_59833[4:0]; // @[Modules.scala 37:46:@7605.4]
  assign _T_59835 = $signed(_T_59834); // @[Modules.scala 37:46:@7606.4]
  assign _T_59855 = $signed(io_in_530) + $signed(io_in_531); // @[Modules.scala 37:46:@7633.4]
  assign _T_59856 = _T_59855[4:0]; // @[Modules.scala 37:46:@7634.4]
  assign _T_59857 = $signed(_T_59856); // @[Modules.scala 37:46:@7635.4]
  assign _T_59877 = $signed(io_in_554) + $signed(io_in_555); // @[Modules.scala 37:46:@7663.4]
  assign _T_59878 = _T_59877[4:0]; // @[Modules.scala 37:46:@7664.4]
  assign _T_59879 = $signed(_T_59878); // @[Modules.scala 37:46:@7665.4]
  assign _T_59880 = $signed(io_in_556) + $signed(io_in_557); // @[Modules.scala 37:46:@7667.4]
  assign _T_59881 = _T_59880[4:0]; // @[Modules.scala 37:46:@7668.4]
  assign _T_59882 = $signed(_T_59881); // @[Modules.scala 37:46:@7669.4]
  assign _T_59889 = $signed(io_in_566) + $signed(io_in_567); // @[Modules.scala 37:46:@7681.4]
  assign _T_59890 = _T_59889[4:0]; // @[Modules.scala 37:46:@7682.4]
  assign _T_59891 = $signed(_T_59890); // @[Modules.scala 37:46:@7683.4]
  assign _T_59898 = $signed(io_in_582) + $signed(io_in_583); // @[Modules.scala 37:46:@7698.4]
  assign _T_59899 = _T_59898[4:0]; // @[Modules.scala 37:46:@7699.4]
  assign _T_59900 = $signed(_T_59899); // @[Modules.scala 37:46:@7700.4]
  assign _T_59904 = $signed(io_in_586) + $signed(io_in_587); // @[Modules.scala 37:46:@7706.4]
  assign _T_59905 = _T_59904[4:0]; // @[Modules.scala 37:46:@7707.4]
  assign _T_59906 = $signed(_T_59905); // @[Modules.scala 37:46:@7708.4]
  assign _T_59914 = $signed(io_in_594) + $signed(io_in_595); // @[Modules.scala 37:46:@7719.4]
  assign _T_59915 = _T_59914[4:0]; // @[Modules.scala 37:46:@7720.4]
  assign _T_59916 = $signed(_T_59915); // @[Modules.scala 37:46:@7721.4]
  assign _T_59922 = $signed(io_in_610) + $signed(io_in_611); // @[Modules.scala 37:46:@7733.4]
  assign _T_59923 = _T_59922[4:0]; // @[Modules.scala 37:46:@7734.4]
  assign _T_59924 = $signed(_T_59923); // @[Modules.scala 37:46:@7735.4]
  assign _T_59932 = $signed(io_in_620) + $signed(io_in_621); // @[Modules.scala 37:46:@7747.4]
  assign _T_59933 = _T_59932[4:0]; // @[Modules.scala 37:46:@7748.4]
  assign _T_59934 = $signed(_T_59933); // @[Modules.scala 37:46:@7749.4]
  assign _T_59945 = $signed(io_in_638) + $signed(io_in_639); // @[Modules.scala 37:46:@7768.4]
  assign _T_59946 = _T_59945[4:0]; // @[Modules.scala 37:46:@7769.4]
  assign _T_59947 = $signed(_T_59946); // @[Modules.scala 37:46:@7770.4]
  assign _T_59979 = $signed(io_in_686) + $signed(io_in_687); // @[Modules.scala 37:46:@7822.4]
  assign _T_59980 = _T_59979[4:0]; // @[Modules.scala 37:46:@7823.4]
  assign _T_59981 = $signed(_T_59980); // @[Modules.scala 37:46:@7824.4]
  assign _T_59987 = $signed(io_in_698) + $signed(io_in_699); // @[Modules.scala 37:46:@7831.4]
  assign _T_59988 = _T_59987[4:0]; // @[Modules.scala 37:46:@7832.4]
  assign _T_59989 = $signed(_T_59988); // @[Modules.scala 37:46:@7833.4]
  assign _T_59999 = $signed(io_in_710) + $signed(io_in_711); // @[Modules.scala 37:46:@7849.4]
  assign _T_60000 = _T_59999[4:0]; // @[Modules.scala 37:46:@7850.4]
  assign _T_60001 = $signed(_T_60000); // @[Modules.scala 37:46:@7851.4]
  assign _T_60020 = $signed(io_in_736) + $signed(io_in_737); // @[Modules.scala 37:46:@7880.4]
  assign _T_60021 = _T_60020[4:0]; // @[Modules.scala 37:46:@7881.4]
  assign _T_60022 = $signed(_T_60021); // @[Modules.scala 37:46:@7882.4]
  assign _T_60023 = $signed(io_in_738) + $signed(io_in_739); // @[Modules.scala 37:46:@7884.4]
  assign _T_60024 = _T_60023[4:0]; // @[Modules.scala 37:46:@7885.4]
  assign _T_60025 = $signed(_T_60024); // @[Modules.scala 37:46:@7886.4]
  assign _T_60026 = $signed(io_in_740) + $signed(io_in_741); // @[Modules.scala 37:46:@7888.4]
  assign _T_60027 = _T_60026[4:0]; // @[Modules.scala 37:46:@7889.4]
  assign _T_60028 = $signed(_T_60027); // @[Modules.scala 37:46:@7890.4]
  assign _T_60029 = $signed(io_in_744) + $signed(io_in_745); // @[Modules.scala 37:46:@7893.4]
  assign _T_60030 = _T_60029[4:0]; // @[Modules.scala 37:46:@7894.4]
  assign _T_60031 = $signed(_T_60030); // @[Modules.scala 37:46:@7895.4]
  assign _T_60032 = $signed(io_in_746) + $signed(io_in_747); // @[Modules.scala 37:46:@7897.4]
  assign _T_60033 = _T_60032[4:0]; // @[Modules.scala 37:46:@7898.4]
  assign _T_60034 = $signed(_T_60033); // @[Modules.scala 37:46:@7899.4]
  assign _T_60036 = $signed(io_in_756) + $signed(io_in_757); // @[Modules.scala 37:46:@7905.4]
  assign _T_60037 = _T_60036[4:0]; // @[Modules.scala 37:46:@7906.4]
  assign _T_60038 = $signed(_T_60037); // @[Modules.scala 37:46:@7907.4]
  assign _T_60046 = $signed(io_in_764) + $signed(io_in_765); // @[Modules.scala 37:46:@7918.4]
  assign _T_60047 = _T_60046[4:0]; // @[Modules.scala 37:46:@7919.4]
  assign _T_60048 = $signed(_T_60047); // @[Modules.scala 37:46:@7920.4]
  assign _T_60052 = $signed(io_in_768) + $signed(io_in_769); // @[Modules.scala 37:46:@7926.4]
  assign _T_60053 = _T_60052[4:0]; // @[Modules.scala 37:46:@7927.4]
  assign _T_60054 = $signed(_T_60053); // @[Modules.scala 37:46:@7928.4]
  assign _T_60055 = $signed(io_in_770) + $signed(io_in_771); // @[Modules.scala 37:46:@7930.4]
  assign _T_60056 = _T_60055[4:0]; // @[Modules.scala 37:46:@7931.4]
  assign _T_60057 = $signed(_T_60056); // @[Modules.scala 37:46:@7932.4]
  assign _T_60058 = $signed(io_in_772) + $signed(io_in_773); // @[Modules.scala 37:46:@7934.4]
  assign _T_60059 = _T_60058[4:0]; // @[Modules.scala 37:46:@7935.4]
  assign _T_60060 = $signed(_T_60059); // @[Modules.scala 37:46:@7936.4]
  assign _T_60061 = $signed(io_in_774) + $signed(io_in_775); // @[Modules.scala 37:46:@7938.4]
  assign _T_60062 = _T_60061[4:0]; // @[Modules.scala 37:46:@7939.4]
  assign _T_60063 = $signed(_T_60062); // @[Modules.scala 37:46:@7940.4]
  assign buffer_3_0 = {{6{io_in_0[4]}},io_in_0}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_1 = {{6{io_in_2[4]}},io_in_2}; // @[Modules.scala 32:22:@8.4]
  assign _T_60068 = $signed(buffer_3_0) + $signed(buffer_3_1); // @[Modules.scala 65:57:@7949.4]
  assign _T_60069 = _T_60068[10:0]; // @[Modules.scala 65:57:@7950.4]
  assign buffer_3_392 = $signed(_T_60069); // @[Modules.scala 65:57:@7951.4]
  assign buffer_3_5 = {{6{io_in_10[4]}},io_in_10}; // @[Modules.scala 32:22:@8.4]
  assign _T_60074 = $signed(11'sh0) + $signed(buffer_3_5); // @[Modules.scala 65:57:@7957.4]
  assign _T_60075 = _T_60074[10:0]; // @[Modules.scala 65:57:@7958.4]
  assign buffer_3_394 = $signed(_T_60075); // @[Modules.scala 65:57:@7959.4]
  assign _T_60080 = $signed(buffer_1_8) + $signed(11'sh0); // @[Modules.scala 65:57:@7965.4]
  assign _T_60081 = _T_60080[10:0]; // @[Modules.scala 65:57:@7966.4]
  assign buffer_3_396 = $signed(_T_60081); // @[Modules.scala 65:57:@7967.4]
  assign _T_60083 = $signed(buffer_2_10) + $signed(buffer_0_11); // @[Modules.scala 65:57:@7969.4]
  assign _T_60084 = _T_60083[10:0]; // @[Modules.scala 65:57:@7970.4]
  assign buffer_3_397 = $signed(_T_60084); // @[Modules.scala 65:57:@7971.4]
  assign buffer_3_12 = {{6{io_in_24[4]}},io_in_24}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_13 = {{6{_T_59455[4]}},_T_59455}; // @[Modules.scala 32:22:@8.4]
  assign _T_60086 = $signed(buffer_3_12) + $signed(buffer_3_13); // @[Modules.scala 65:57:@7973.4]
  assign _T_60087 = _T_60086[10:0]; // @[Modules.scala 65:57:@7974.4]
  assign buffer_3_398 = $signed(_T_60087); // @[Modules.scala 65:57:@7975.4]
  assign buffer_3_14 = {{6{_T_59458[4]}},_T_59458}; // @[Modules.scala 32:22:@8.4]
  assign _T_60089 = $signed(buffer_3_14) + $signed(11'sh0); // @[Modules.scala 65:57:@7977.4]
  assign _T_60090 = _T_60089[10:0]; // @[Modules.scala 65:57:@7978.4]
  assign buffer_3_399 = $signed(_T_60090); // @[Modules.scala 65:57:@7979.4]
  assign buffer_3_16 = {{6{io_in_32[4]}},io_in_32}; // @[Modules.scala 32:22:@8.4]
  assign _T_60092 = $signed(buffer_3_16) + $signed(11'sh0); // @[Modules.scala 65:57:@7981.4]
  assign _T_60093 = _T_60092[10:0]; // @[Modules.scala 65:57:@7982.4]
  assign buffer_3_400 = $signed(_T_60093); // @[Modules.scala 65:57:@7983.4]
  assign _T_60101 = $signed(buffer_1_22) + $signed(11'sh0); // @[Modules.scala 65:57:@7993.4]
  assign _T_60102 = _T_60101[10:0]; // @[Modules.scala 65:57:@7994.4]
  assign buffer_3_403 = $signed(_T_60102); // @[Modules.scala 65:57:@7995.4]
  assign _T_60104 = $signed(11'sh0) + $signed(buffer_1_25); // @[Modules.scala 65:57:@7997.4]
  assign _T_60105 = _T_60104[10:0]; // @[Modules.scala 65:57:@7998.4]
  assign buffer_3_404 = $signed(_T_60105); // @[Modules.scala 65:57:@7999.4]
  assign buffer_3_26 = {{6{io_in_53[4]}},io_in_53}; // @[Modules.scala 32:22:@8.4]
  assign _T_60107 = $signed(buffer_3_26) + $signed(11'sh0); // @[Modules.scala 65:57:@8001.4]
  assign _T_60108 = _T_60107[10:0]; // @[Modules.scala 65:57:@8002.4]
  assign buffer_3_405 = $signed(_T_60108); // @[Modules.scala 65:57:@8003.4]
  assign buffer_3_29 = {{6{io_in_58[4]}},io_in_58}; // @[Modules.scala 32:22:@8.4]
  assign _T_60110 = $signed(11'sh0) + $signed(buffer_3_29); // @[Modules.scala 65:57:@8005.4]
  assign _T_60111 = _T_60110[10:0]; // @[Modules.scala 65:57:@8006.4]
  assign buffer_3_406 = $signed(_T_60111); // @[Modules.scala 65:57:@8007.4]
  assign buffer_3_30 = {{6{io_in_61[4]}},io_in_61}; // @[Modules.scala 32:22:@8.4]
  assign _T_60113 = $signed(buffer_3_30) + $signed(11'sh0); // @[Modules.scala 65:57:@8009.4]
  assign _T_60114 = _T_60113[10:0]; // @[Modules.scala 65:57:@8010.4]
  assign buffer_3_407 = $signed(_T_60114); // @[Modules.scala 65:57:@8011.4]
  assign _T_60128 = $signed(buffer_1_40) + $signed(buffer_2_41); // @[Modules.scala 65:57:@8029.4]
  assign _T_60129 = _T_60128[10:0]; // @[Modules.scala 65:57:@8030.4]
  assign buffer_3_412 = $signed(_T_60129); // @[Modules.scala 65:57:@8031.4]
  assign buffer_3_43 = {{6{io_in_86[4]}},io_in_86}; // @[Modules.scala 32:22:@8.4]
  assign _T_60131 = $signed(buffer_0_42) + $signed(buffer_3_43); // @[Modules.scala 65:57:@8033.4]
  assign _T_60132 = _T_60131[10:0]; // @[Modules.scala 65:57:@8034.4]
  assign buffer_3_413 = $signed(_T_60132); // @[Modules.scala 65:57:@8035.4]
  assign _T_60137 = $signed(11'sh0) + $signed(buffer_0_47); // @[Modules.scala 65:57:@8041.4]
  assign _T_60138 = _T_60137[10:0]; // @[Modules.scala 65:57:@8042.4]
  assign buffer_3_415 = $signed(_T_60138); // @[Modules.scala 65:57:@8043.4]
  assign buffer_3_49 = {{6{io_in_98[4]}},io_in_98}; // @[Modules.scala 32:22:@8.4]
  assign _T_60140 = $signed(buffer_1_48) + $signed(buffer_3_49); // @[Modules.scala 65:57:@8045.4]
  assign _T_60141 = _T_60140[10:0]; // @[Modules.scala 65:57:@8046.4]
  assign buffer_3_416 = $signed(_T_60141); // @[Modules.scala 65:57:@8047.4]
  assign _T_60143 = $signed(buffer_0_50) + $signed(11'sh0); // @[Modules.scala 65:57:@8049.4]
  assign _T_60144 = _T_60143[10:0]; // @[Modules.scala 65:57:@8050.4]
  assign buffer_3_417 = $signed(_T_60144); // @[Modules.scala 65:57:@8051.4]
  assign buffer_3_54 = {{6{io_in_109[4]}},io_in_109}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_55 = {{6{io_in_110[4]}},io_in_110}; // @[Modules.scala 32:22:@8.4]
  assign _T_60149 = $signed(buffer_3_54) + $signed(buffer_3_55); // @[Modules.scala 65:57:@8057.4]
  assign _T_60150 = _T_60149[10:0]; // @[Modules.scala 65:57:@8058.4]
  assign buffer_3_419 = $signed(_T_60150); // @[Modules.scala 65:57:@8059.4]
  assign buffer_3_56 = {{6{io_in_112[4]}},io_in_112}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_57 = {{6{_T_59508[4]}},_T_59508}; // @[Modules.scala 32:22:@8.4]
  assign _T_60152 = $signed(buffer_3_56) + $signed(buffer_3_57); // @[Modules.scala 65:57:@8061.4]
  assign _T_60153 = _T_60152[10:0]; // @[Modules.scala 65:57:@8062.4]
  assign buffer_3_420 = $signed(_T_60153); // @[Modules.scala 65:57:@8063.4]
  assign _T_60155 = $signed(11'sh0) + $signed(buffer_0_59); // @[Modules.scala 65:57:@8065.4]
  assign _T_60156 = _T_60155[10:0]; // @[Modules.scala 65:57:@8066.4]
  assign buffer_3_421 = $signed(_T_60156); // @[Modules.scala 65:57:@8067.4]
  assign buffer_3_60 = {{6{_T_59515[4]}},_T_59515}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_61 = {{6{_T_59518[4]}},_T_59518}; // @[Modules.scala 32:22:@8.4]
  assign _T_60158 = $signed(buffer_3_60) + $signed(buffer_3_61); // @[Modules.scala 65:57:@8069.4]
  assign _T_60159 = _T_60158[10:0]; // @[Modules.scala 65:57:@8070.4]
  assign buffer_3_422 = $signed(_T_60159); // @[Modules.scala 65:57:@8071.4]
  assign buffer_3_62 = {{6{_T_59521[4]}},_T_59521}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_63 = {{6{_T_59524[4]}},_T_59524}; // @[Modules.scala 32:22:@8.4]
  assign _T_60161 = $signed(buffer_3_62) + $signed(buffer_3_63); // @[Modules.scala 65:57:@8073.4]
  assign _T_60162 = _T_60161[10:0]; // @[Modules.scala 65:57:@8074.4]
  assign buffer_3_423 = $signed(_T_60162); // @[Modules.scala 65:57:@8075.4]
  assign buffer_3_67 = {{6{io_in_134[4]}},io_in_134}; // @[Modules.scala 32:22:@8.4]
  assign _T_60167 = $signed(11'sh0) + $signed(buffer_3_67); // @[Modules.scala 65:57:@8081.4]
  assign _T_60168 = _T_60167[10:0]; // @[Modules.scala 65:57:@8082.4]
  assign buffer_3_425 = $signed(_T_60168); // @[Modules.scala 65:57:@8083.4]
  assign buffer_3_69 = {{6{io_in_138[4]}},io_in_138}; // @[Modules.scala 32:22:@8.4]
  assign _T_60170 = $signed(buffer_1_68) + $signed(buffer_3_69); // @[Modules.scala 65:57:@8085.4]
  assign _T_60171 = _T_60170[10:0]; // @[Modules.scala 65:57:@8086.4]
  assign buffer_3_426 = $signed(_T_60171); // @[Modules.scala 65:57:@8087.4]
  assign _T_60173 = $signed(buffer_0_70) + $signed(buffer_1_71); // @[Modules.scala 65:57:@8089.4]
  assign _T_60174 = _T_60173[10:0]; // @[Modules.scala 65:57:@8090.4]
  assign buffer_3_427 = $signed(_T_60174); // @[Modules.scala 65:57:@8091.4]
  assign buffer_3_72 = {{6{io_in_145[4]}},io_in_145}; // @[Modules.scala 32:22:@8.4]
  assign _T_60176 = $signed(buffer_3_72) + $signed(buffer_0_73); // @[Modules.scala 65:57:@8093.4]
  assign _T_60177 = _T_60176[10:0]; // @[Modules.scala 65:57:@8094.4]
  assign buffer_3_428 = $signed(_T_60177); // @[Modules.scala 65:57:@8095.4]
  assign buffer_3_75 = {{6{_T_59546[4]}},_T_59546}; // @[Modules.scala 32:22:@8.4]
  assign _T_60179 = $signed(buffer_0_74) + $signed(buffer_3_75); // @[Modules.scala 65:57:@8097.4]
  assign _T_60180 = _T_60179[10:0]; // @[Modules.scala 65:57:@8098.4]
  assign buffer_3_429 = $signed(_T_60180); // @[Modules.scala 65:57:@8099.4]
  assign buffer_3_76 = {{6{io_in_153[4]}},io_in_153}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_77 = {{6{_T_59549[4]}},_T_59549}; // @[Modules.scala 32:22:@8.4]
  assign _T_60182 = $signed(buffer_3_76) + $signed(buffer_3_77); // @[Modules.scala 65:57:@8101.4]
  assign _T_60183 = _T_60182[10:0]; // @[Modules.scala 65:57:@8102.4]
  assign buffer_3_430 = $signed(_T_60183); // @[Modules.scala 65:57:@8103.4]
  assign buffer_3_79 = {{6{_T_59552[4]}},_T_59552}; // @[Modules.scala 32:22:@8.4]
  assign _T_60185 = $signed(buffer_1_78) + $signed(buffer_3_79); // @[Modules.scala 65:57:@8105.4]
  assign _T_60186 = _T_60185[10:0]; // @[Modules.scala 65:57:@8106.4]
  assign buffer_3_431 = $signed(_T_60186); // @[Modules.scala 65:57:@8107.4]
  assign buffer_3_86 = {{6{_T_59570[4]}},_T_59570}; // @[Modules.scala 32:22:@8.4]
  assign _T_60197 = $signed(buffer_3_86) + $signed(buffer_1_87); // @[Modules.scala 65:57:@8121.4]
  assign _T_60198 = _T_60197[10:0]; // @[Modules.scala 65:57:@8122.4]
  assign buffer_3_435 = $signed(_T_60198); // @[Modules.scala 65:57:@8123.4]
  assign buffer_3_89 = {{6{_T_59579[4]}},_T_59579}; // @[Modules.scala 32:22:@8.4]
  assign _T_60200 = $signed(buffer_1_88) + $signed(buffer_3_89); // @[Modules.scala 65:57:@8125.4]
  assign _T_60201 = _T_60200[10:0]; // @[Modules.scala 65:57:@8126.4]
  assign buffer_3_436 = $signed(_T_60201); // @[Modules.scala 65:57:@8127.4]
  assign buffer_3_90 = {{6{_T_59582[4]}},_T_59582}; // @[Modules.scala 32:22:@8.4]
  assign _T_60203 = $signed(buffer_3_90) + $signed(11'sh0); // @[Modules.scala 65:57:@8129.4]
  assign _T_60204 = _T_60203[10:0]; // @[Modules.scala 65:57:@8130.4]
  assign buffer_3_437 = $signed(_T_60204); // @[Modules.scala 65:57:@8131.4]
  assign buffer_3_92 = {{6{io_in_184[4]}},io_in_184}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_93 = {{6{io_in_186[4]}},io_in_186}; // @[Modules.scala 32:22:@8.4]
  assign _T_60206 = $signed(buffer_3_92) + $signed(buffer_3_93); // @[Modules.scala 65:57:@8133.4]
  assign _T_60207 = _T_60206[10:0]; // @[Modules.scala 65:57:@8134.4]
  assign buffer_3_438 = $signed(_T_60207); // @[Modules.scala 65:57:@8135.4]
  assign _T_60209 = $signed(buffer_1_94) + $signed(buffer_0_95); // @[Modules.scala 65:57:@8137.4]
  assign _T_60210 = _T_60209[10:0]; // @[Modules.scala 65:57:@8138.4]
  assign buffer_3_439 = $signed(_T_60210); // @[Modules.scala 65:57:@8139.4]
  assign buffer_3_98 = {{6{io_in_197[4]}},io_in_197}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_99 = {{6{_T_59592[4]}},_T_59592}; // @[Modules.scala 32:22:@8.4]
  assign _T_60215 = $signed(buffer_3_98) + $signed(buffer_3_99); // @[Modules.scala 65:57:@8145.4]
  assign _T_60216 = _T_60215[10:0]; // @[Modules.scala 65:57:@8146.4]
  assign buffer_3_441 = $signed(_T_60216); // @[Modules.scala 65:57:@8147.4]
  assign buffer_3_100 = {{6{_T_59595[4]}},_T_59595}; // @[Modules.scala 32:22:@8.4]
  assign _T_60218 = $signed(buffer_3_100) + $signed(buffer_1_101); // @[Modules.scala 65:57:@8149.4]
  assign _T_60219 = _T_60218[10:0]; // @[Modules.scala 65:57:@8150.4]
  assign buffer_3_442 = $signed(_T_60219); // @[Modules.scala 65:57:@8151.4]
  assign buffer_3_103 = {{6{_T_59601[4]}},_T_59601}; // @[Modules.scala 32:22:@8.4]
  assign _T_60221 = $signed(buffer_1_102) + $signed(buffer_3_103); // @[Modules.scala 65:57:@8153.4]
  assign _T_60222 = _T_60221[10:0]; // @[Modules.scala 65:57:@8154.4]
  assign buffer_3_443 = $signed(_T_60222); // @[Modules.scala 65:57:@8155.4]
  assign buffer_3_104 = {{6{_T_59604[4]}},_T_59604}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_105 = {{6{io_in_210[4]}},io_in_210}; // @[Modules.scala 32:22:@8.4]
  assign _T_60224 = $signed(buffer_3_104) + $signed(buffer_3_105); // @[Modules.scala 65:57:@8157.4]
  assign _T_60225 = _T_60224[10:0]; // @[Modules.scala 65:57:@8158.4]
  assign buffer_3_444 = $signed(_T_60225); // @[Modules.scala 65:57:@8159.4]
  assign buffer_3_106 = {{6{_T_59607[4]}},_T_59607}; // @[Modules.scala 32:22:@8.4]
  assign _T_60227 = $signed(buffer_3_106) + $signed(buffer_2_107); // @[Modules.scala 65:57:@8161.4]
  assign _T_60228 = _T_60227[10:0]; // @[Modules.scala 65:57:@8162.4]
  assign buffer_3_445 = $signed(_T_60228); // @[Modules.scala 65:57:@8163.4]
  assign buffer_3_109 = {{6{io_in_218[4]}},io_in_218}; // @[Modules.scala 32:22:@8.4]
  assign _T_60230 = $signed(buffer_1_108) + $signed(buffer_3_109); // @[Modules.scala 65:57:@8165.4]
  assign _T_60231 = _T_60230[10:0]; // @[Modules.scala 65:57:@8166.4]
  assign buffer_3_446 = $signed(_T_60231); // @[Modules.scala 65:57:@8167.4]
  assign buffer_3_113 = {{6{_T_59622[4]}},_T_59622}; // @[Modules.scala 32:22:@8.4]
  assign _T_60236 = $signed(buffer_1_112) + $signed(buffer_3_113); // @[Modules.scala 65:57:@8173.4]
  assign _T_60237 = _T_60236[10:0]; // @[Modules.scala 65:57:@8174.4]
  assign buffer_3_448 = $signed(_T_60237); // @[Modules.scala 65:57:@8175.4]
  assign buffer_3_114 = {{6{_T_59625[4]}},_T_59625}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_115 = {{6{io_in_231[4]}},io_in_231}; // @[Modules.scala 32:22:@8.4]
  assign _T_60239 = $signed(buffer_3_114) + $signed(buffer_3_115); // @[Modules.scala 65:57:@8177.4]
  assign _T_60240 = _T_60239[10:0]; // @[Modules.scala 65:57:@8178.4]
  assign buffer_3_449 = $signed(_T_60240); // @[Modules.scala 65:57:@8179.4]
  assign buffer_3_116 = {{6{io_in_232[4]}},io_in_232}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_117 = {{6{_T_59628[4]}},_T_59628}; // @[Modules.scala 32:22:@8.4]
  assign _T_60242 = $signed(buffer_3_116) + $signed(buffer_3_117); // @[Modules.scala 65:57:@8181.4]
  assign _T_60243 = _T_60242[10:0]; // @[Modules.scala 65:57:@8182.4]
  assign buffer_3_450 = $signed(_T_60243); // @[Modules.scala 65:57:@8183.4]
  assign buffer_3_118 = {{6{_T_59631[4]}},_T_59631}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_119 = {{6{_T_59634[4]}},_T_59634}; // @[Modules.scala 32:22:@8.4]
  assign _T_60245 = $signed(buffer_3_118) + $signed(buffer_3_119); // @[Modules.scala 65:57:@8185.4]
  assign _T_60246 = _T_60245[10:0]; // @[Modules.scala 65:57:@8186.4]
  assign buffer_3_451 = $signed(_T_60246); // @[Modules.scala 65:57:@8187.4]
  assign buffer_3_121 = {{6{_T_59640[4]}},_T_59640}; // @[Modules.scala 32:22:@8.4]
  assign _T_60248 = $signed(buffer_1_120) + $signed(buffer_3_121); // @[Modules.scala 65:57:@8189.4]
  assign _T_60249 = _T_60248[10:0]; // @[Modules.scala 65:57:@8190.4]
  assign buffer_3_452 = $signed(_T_60249); // @[Modules.scala 65:57:@8191.4]
  assign buffer_3_122 = {{6{io_in_244[4]}},io_in_244}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_123 = {{6{_T_59643[4]}},_T_59643}; // @[Modules.scala 32:22:@8.4]
  assign _T_60251 = $signed(buffer_3_122) + $signed(buffer_3_123); // @[Modules.scala 65:57:@8193.4]
  assign _T_60252 = _T_60251[10:0]; // @[Modules.scala 65:57:@8194.4]
  assign buffer_3_453 = $signed(_T_60252); // @[Modules.scala 65:57:@8195.4]
  assign buffer_3_126 = {{6{_T_59652[4]}},_T_59652}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_127 = {{6{_T_59655[4]}},_T_59655}; // @[Modules.scala 32:22:@8.4]
  assign _T_60257 = $signed(buffer_3_126) + $signed(buffer_3_127); // @[Modules.scala 65:57:@8201.4]
  assign _T_60258 = _T_60257[10:0]; // @[Modules.scala 65:57:@8202.4]
  assign buffer_3_455 = $signed(_T_60258); // @[Modules.scala 65:57:@8203.4]
  assign buffer_3_128 = {{6{_T_59658[4]}},_T_59658}; // @[Modules.scala 32:22:@8.4]
  assign _T_60260 = $signed(buffer_3_128) + $signed(11'sh0); // @[Modules.scala 65:57:@8205.4]
  assign _T_60261 = _T_60260[10:0]; // @[Modules.scala 65:57:@8206.4]
  assign buffer_3_456 = $signed(_T_60261); // @[Modules.scala 65:57:@8207.4]
  assign buffer_3_132 = {{6{_T_59662[4]}},_T_59662}; // @[Modules.scala 32:22:@8.4]
  assign _T_60266 = $signed(buffer_3_132) + $signed(buffer_1_133); // @[Modules.scala 65:57:@8213.4]
  assign _T_60267 = _T_60266[10:0]; // @[Modules.scala 65:57:@8214.4]
  assign buffer_3_458 = $signed(_T_60267); // @[Modules.scala 65:57:@8215.4]
  assign buffer_3_134 = {{6{_T_59668[4]}},_T_59668}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_135 = {{6{_T_59671[4]}},_T_59671}; // @[Modules.scala 32:22:@8.4]
  assign _T_60269 = $signed(buffer_3_134) + $signed(buffer_3_135); // @[Modules.scala 65:57:@8217.4]
  assign _T_60270 = _T_60269[10:0]; // @[Modules.scala 65:57:@8218.4]
  assign buffer_3_459 = $signed(_T_60270); // @[Modules.scala 65:57:@8219.4]
  assign buffer_3_136 = {{6{_T_59674[4]}},_T_59674}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_137 = {{6{_T_59677[4]}},_T_59677}; // @[Modules.scala 32:22:@8.4]
  assign _T_60272 = $signed(buffer_3_136) + $signed(buffer_3_137); // @[Modules.scala 65:57:@8221.4]
  assign _T_60273 = _T_60272[10:0]; // @[Modules.scala 65:57:@8222.4]
  assign buffer_3_460 = $signed(_T_60273); // @[Modules.scala 65:57:@8223.4]
  assign buffer_3_140 = {{6{_T_59686[4]}},_T_59686}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_141 = {{6{_T_59689[4]}},_T_59689}; // @[Modules.scala 32:22:@8.4]
  assign _T_60278 = $signed(buffer_3_140) + $signed(buffer_3_141); // @[Modules.scala 65:57:@8229.4]
  assign _T_60279 = _T_60278[10:0]; // @[Modules.scala 65:57:@8230.4]
  assign buffer_3_462 = $signed(_T_60279); // @[Modules.scala 65:57:@8231.4]
  assign buffer_3_142 = {{6{io_in_284[4]}},io_in_284}; // @[Modules.scala 32:22:@8.4]
  assign _T_60281 = $signed(buffer_3_142) + $signed(11'sh0); // @[Modules.scala 65:57:@8233.4]
  assign _T_60282 = _T_60281[10:0]; // @[Modules.scala 65:57:@8234.4]
  assign buffer_3_463 = $signed(_T_60282); // @[Modules.scala 65:57:@8235.4]
  assign buffer_3_147 = {{6{io_in_295[4]}},io_in_295}; // @[Modules.scala 32:22:@8.4]
  assign _T_60287 = $signed(11'sh0) + $signed(buffer_3_147); // @[Modules.scala 65:57:@8241.4]
  assign _T_60288 = _T_60287[10:0]; // @[Modules.scala 65:57:@8242.4]
  assign buffer_3_465 = $signed(_T_60288); // @[Modules.scala 65:57:@8243.4]
  assign buffer_3_148 = {{6{_T_59696[4]}},_T_59696}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_149 = {{6{io_in_298[4]}},io_in_298}; // @[Modules.scala 32:22:@8.4]
  assign _T_60290 = $signed(buffer_3_148) + $signed(buffer_3_149); // @[Modules.scala 65:57:@8245.4]
  assign _T_60291 = _T_60290[10:0]; // @[Modules.scala 65:57:@8246.4]
  assign buffer_3_466 = $signed(_T_60291); // @[Modules.scala 65:57:@8247.4]
  assign buffer_3_150 = {{6{io_in_300[4]}},io_in_300}; // @[Modules.scala 32:22:@8.4]
  assign _T_60293 = $signed(buffer_3_150) + $signed(11'sh0); // @[Modules.scala 65:57:@8249.4]
  assign _T_60294 = _T_60293[10:0]; // @[Modules.scala 65:57:@8250.4]
  assign buffer_3_467 = $signed(_T_60294); // @[Modules.scala 65:57:@8251.4]
  assign buffer_3_154 = {{6{io_in_309[4]}},io_in_309}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_155 = {{6{_T_59706[4]}},_T_59706}; // @[Modules.scala 32:22:@8.4]
  assign _T_60299 = $signed(buffer_3_154) + $signed(buffer_3_155); // @[Modules.scala 65:57:@8257.4]
  assign _T_60300 = _T_60299[10:0]; // @[Modules.scala 65:57:@8258.4]
  assign buffer_3_469 = $signed(_T_60300); // @[Modules.scala 65:57:@8259.4]
  assign buffer_3_167 = {{6{io_in_334[4]}},io_in_334}; // @[Modules.scala 32:22:@8.4]
  assign _T_60317 = $signed(11'sh0) + $signed(buffer_3_167); // @[Modules.scala 65:57:@8281.4]
  assign _T_60318 = _T_60317[10:0]; // @[Modules.scala 65:57:@8282.4]
  assign buffer_3_475 = $signed(_T_60318); // @[Modules.scala 65:57:@8283.4]
  assign buffer_3_168 = {{6{io_in_337[4]}},io_in_337}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_169 = {{6{io_in_338[4]}},io_in_338}; // @[Modules.scala 32:22:@8.4]
  assign _T_60320 = $signed(buffer_3_168) + $signed(buffer_3_169); // @[Modules.scala 65:57:@8285.4]
  assign _T_60321 = _T_60320[10:0]; // @[Modules.scala 65:57:@8286.4]
  assign buffer_3_476 = $signed(_T_60321); // @[Modules.scala 65:57:@8287.4]
  assign buffer_3_182 = {{6{io_in_365[4]}},io_in_365}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_183 = {{6{io_in_366[4]}},io_in_366}; // @[Modules.scala 32:22:@8.4]
  assign _T_60341 = $signed(buffer_3_182) + $signed(buffer_3_183); // @[Modules.scala 65:57:@8313.4]
  assign _T_60342 = _T_60341[10:0]; // @[Modules.scala 65:57:@8314.4]
  assign buffer_3_483 = $signed(_T_60342); // @[Modules.scala 65:57:@8315.4]
  assign buffer_3_187 = {{6{io_in_375[4]}},io_in_375}; // @[Modules.scala 32:22:@8.4]
  assign _T_60347 = $signed(11'sh0) + $signed(buffer_3_187); // @[Modules.scala 65:57:@8321.4]
  assign _T_60348 = _T_60347[10:0]; // @[Modules.scala 65:57:@8322.4]
  assign buffer_3_485 = $signed(_T_60348); // @[Modules.scala 65:57:@8323.4]
  assign buffer_3_190 = {{6{io_in_381[4]}},io_in_381}; // @[Modules.scala 32:22:@8.4]
  assign _T_60353 = $signed(buffer_3_190) + $signed(11'sh0); // @[Modules.scala 65:57:@8329.4]
  assign _T_60354 = _T_60353[10:0]; // @[Modules.scala 65:57:@8330.4]
  assign buffer_3_487 = $signed(_T_60354); // @[Modules.scala 65:57:@8331.4]
  assign buffer_3_195 = {{6{_T_59740[4]}},_T_59740}; // @[Modules.scala 32:22:@8.4]
  assign _T_60359 = $signed(11'sh0) + $signed(buffer_3_195); // @[Modules.scala 65:57:@8337.4]
  assign _T_60360 = _T_60359[10:0]; // @[Modules.scala 65:57:@8338.4]
  assign buffer_3_489 = $signed(_T_60360); // @[Modules.scala 65:57:@8339.4]
  assign buffer_3_197 = {{6{io_in_394[4]}},io_in_394}; // @[Modules.scala 32:22:@8.4]
  assign _T_60362 = $signed(buffer_1_196) + $signed(buffer_3_197); // @[Modules.scala 65:57:@8341.4]
  assign _T_60363 = _T_60362[10:0]; // @[Modules.scala 65:57:@8342.4]
  assign buffer_3_490 = $signed(_T_60363); // @[Modules.scala 65:57:@8343.4]
  assign buffer_3_200 = {{6{io_in_401[4]}},io_in_401}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_201 = {{6{io_in_402[4]}},io_in_402}; // @[Modules.scala 32:22:@8.4]
  assign _T_60368 = $signed(buffer_3_200) + $signed(buffer_3_201); // @[Modules.scala 65:57:@8349.4]
  assign _T_60369 = _T_60368[10:0]; // @[Modules.scala 65:57:@8350.4]
  assign buffer_3_492 = $signed(_T_60369); // @[Modules.scala 65:57:@8351.4]
  assign buffer_3_205 = {{6{io_in_410[4]}},io_in_410}; // @[Modules.scala 32:22:@8.4]
  assign _T_60374 = $signed(11'sh0) + $signed(buffer_3_205); // @[Modules.scala 65:57:@8357.4]
  assign _T_60375 = _T_60374[10:0]; // @[Modules.scala 65:57:@8358.4]
  assign buffer_3_494 = $signed(_T_60375); // @[Modules.scala 65:57:@8359.4]
  assign buffer_3_208 = {{6{io_in_417[4]}},io_in_417}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_209 = {{6{_T_59753[4]}},_T_59753}; // @[Modules.scala 32:22:@8.4]
  assign _T_60380 = $signed(buffer_3_208) + $signed(buffer_3_209); // @[Modules.scala 65:57:@8365.4]
  assign _T_60381 = _T_60380[10:0]; // @[Modules.scala 65:57:@8366.4]
  assign buffer_3_496 = $signed(_T_60381); // @[Modules.scala 65:57:@8367.4]
  assign buffer_3_210 = {{6{io_in_420[4]}},io_in_420}; // @[Modules.scala 32:22:@8.4]
  assign _T_60383 = $signed(buffer_3_210) + $signed(buffer_2_211); // @[Modules.scala 65:57:@8369.4]
  assign _T_60384 = _T_60383[10:0]; // @[Modules.scala 65:57:@8370.4]
  assign buffer_3_497 = $signed(_T_60384); // @[Modules.scala 65:57:@8371.4]
  assign buffer_3_212 = {{6{_T_59759[4]}},_T_59759}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_213 = {{6{io_in_427[4]}},io_in_427}; // @[Modules.scala 32:22:@8.4]
  assign _T_60386 = $signed(buffer_3_212) + $signed(buffer_3_213); // @[Modules.scala 65:57:@8373.4]
  assign _T_60387 = _T_60386[10:0]; // @[Modules.scala 65:57:@8374.4]
  assign buffer_3_498 = $signed(_T_60387); // @[Modules.scala 65:57:@8375.4]
  assign buffer_3_220 = {{6{io_in_441[4]}},io_in_441}; // @[Modules.scala 32:22:@8.4]
  assign _T_60398 = $signed(buffer_3_220) + $signed(11'sh0); // @[Modules.scala 65:57:@8389.4]
  assign _T_60399 = _T_60398[10:0]; // @[Modules.scala 65:57:@8390.4]
  assign buffer_3_502 = $signed(_T_60399); // @[Modules.scala 65:57:@8391.4]
  assign buffer_3_222 = {{6{_T_59771[4]}},_T_59771}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_223 = {{6{_T_59774[4]}},_T_59774}; // @[Modules.scala 32:22:@8.4]
  assign _T_60401 = $signed(buffer_3_222) + $signed(buffer_3_223); // @[Modules.scala 65:57:@8393.4]
  assign _T_60402 = _T_60401[10:0]; // @[Modules.scala 65:57:@8394.4]
  assign buffer_3_503 = $signed(_T_60402); // @[Modules.scala 65:57:@8395.4]
  assign buffer_3_224 = {{6{io_in_448[4]}},io_in_448}; // @[Modules.scala 32:22:@8.4]
  assign _T_60404 = $signed(buffer_3_224) + $signed(buffer_1_225); // @[Modules.scala 65:57:@8397.4]
  assign _T_60405 = _T_60404[10:0]; // @[Modules.scala 65:57:@8398.4]
  assign buffer_3_504 = $signed(_T_60405); // @[Modules.scala 65:57:@8399.4]
  assign buffer_3_226 = {{6{_T_59780[4]}},_T_59780}; // @[Modules.scala 32:22:@8.4]
  assign _T_60407 = $signed(buffer_3_226) + $signed(buffer_0_227); // @[Modules.scala 65:57:@8401.4]
  assign _T_60408 = _T_60407[10:0]; // @[Modules.scala 65:57:@8402.4]
  assign buffer_3_505 = $signed(_T_60408); // @[Modules.scala 65:57:@8403.4]
  assign _T_60416 = $signed(11'sh0) + $signed(buffer_0_233); // @[Modules.scala 65:57:@8413.4]
  assign _T_60417 = _T_60416[10:0]; // @[Modules.scala 65:57:@8414.4]
  assign buffer_3_508 = $signed(_T_60417); // @[Modules.scala 65:57:@8415.4]
  assign buffer_3_236 = {{6{_T_59800[4]}},_T_59800}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_237 = {{6{_T_59803[4]}},_T_59803}; // @[Modules.scala 32:22:@8.4]
  assign _T_60422 = $signed(buffer_3_236) + $signed(buffer_3_237); // @[Modules.scala 65:57:@8421.4]
  assign _T_60423 = _T_60422[10:0]; // @[Modules.scala 65:57:@8422.4]
  assign buffer_3_510 = $signed(_T_60423); // @[Modules.scala 65:57:@8423.4]
  assign _T_60425 = $signed(11'sh0) + $signed(buffer_1_239); // @[Modules.scala 65:57:@8425.4]
  assign _T_60426 = _T_60425[10:0]; // @[Modules.scala 65:57:@8426.4]
  assign buffer_3_511 = $signed(_T_60426); // @[Modules.scala 65:57:@8427.4]
  assign buffer_3_240 = {{6{_T_59810[4]}},_T_59810}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_241 = {{6{io_in_482[4]}},io_in_482}; // @[Modules.scala 32:22:@8.4]
  assign _T_60428 = $signed(buffer_3_240) + $signed(buffer_3_241); // @[Modules.scala 65:57:@8429.4]
  assign _T_60429 = _T_60428[10:0]; // @[Modules.scala 65:57:@8430.4]
  assign buffer_3_512 = $signed(_T_60429); // @[Modules.scala 65:57:@8431.4]
  assign buffer_3_246 = {{6{io_in_493[4]}},io_in_493}; // @[Modules.scala 32:22:@8.4]
  assign _T_60437 = $signed(buffer_3_246) + $signed(buffer_1_247); // @[Modules.scala 65:57:@8441.4]
  assign _T_60438 = _T_60437[10:0]; // @[Modules.scala 65:57:@8442.4]
  assign buffer_3_515 = $signed(_T_60438); // @[Modules.scala 65:57:@8443.4]
  assign buffer_3_250 = {{6{_T_59826[4]}},_T_59826}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_251 = {{6{_T_59829[4]}},_T_59829}; // @[Modules.scala 32:22:@8.4]
  assign _T_60443 = $signed(buffer_3_250) + $signed(buffer_3_251); // @[Modules.scala 65:57:@8449.4]
  assign _T_60444 = _T_60443[10:0]; // @[Modules.scala 65:57:@8450.4]
  assign buffer_3_517 = $signed(_T_60444); // @[Modules.scala 65:57:@8451.4]
  assign buffer_3_252 = {{6{io_in_504[4]}},io_in_504}; // @[Modules.scala 32:22:@8.4]
  assign _T_60446 = $signed(buffer_3_252) + $signed(buffer_1_253); // @[Modules.scala 65:57:@8453.4]
  assign _T_60447 = _T_60446[10:0]; // @[Modules.scala 65:57:@8454.4]
  assign buffer_3_518 = $signed(_T_60447); // @[Modules.scala 65:57:@8455.4]
  assign buffer_3_254 = {{6{_T_59835[4]}},_T_59835}; // @[Modules.scala 32:22:@8.4]
  assign _T_60449 = $signed(buffer_3_254) + $signed(buffer_1_255); // @[Modules.scala 65:57:@8457.4]
  assign _T_60450 = _T_60449[10:0]; // @[Modules.scala 65:57:@8458.4]
  assign buffer_3_519 = $signed(_T_60450); // @[Modules.scala 65:57:@8459.4]
  assign buffer_3_265 = {{6{_T_59857[4]}},_T_59857}; // @[Modules.scala 32:22:@8.4]
  assign _T_60464 = $signed(buffer_0_264) + $signed(buffer_3_265); // @[Modules.scala 65:57:@8477.4]
  assign _T_60465 = _T_60464[10:0]; // @[Modules.scala 65:57:@8478.4]
  assign buffer_3_524 = $signed(_T_60465); // @[Modules.scala 65:57:@8479.4]
  assign buffer_3_270 = {{6{io_in_540[4]}},io_in_540}; // @[Modules.scala 32:22:@8.4]
  assign _T_60473 = $signed(buffer_3_270) + $signed(11'sh0); // @[Modules.scala 65:57:@8489.4]
  assign _T_60474 = _T_60473[10:0]; // @[Modules.scala 65:57:@8490.4]
  assign buffer_3_527 = $signed(_T_60474); // @[Modules.scala 65:57:@8491.4]
  assign buffer_3_273 = {{6{io_in_546[4]}},io_in_546}; // @[Modules.scala 32:22:@8.4]
  assign _T_60476 = $signed(11'sh0) + $signed(buffer_3_273); // @[Modules.scala 65:57:@8493.4]
  assign _T_60477 = _T_60476[10:0]; // @[Modules.scala 65:57:@8494.4]
  assign buffer_3_528 = $signed(_T_60477); // @[Modules.scala 65:57:@8495.4]
  assign buffer_3_277 = {{6{_T_59879[4]}},_T_59879}; // @[Modules.scala 32:22:@8.4]
  assign _T_60482 = $signed(buffer_2_276) + $signed(buffer_3_277); // @[Modules.scala 65:57:@8501.4]
  assign _T_60483 = _T_60482[10:0]; // @[Modules.scala 65:57:@8502.4]
  assign buffer_3_530 = $signed(_T_60483); // @[Modules.scala 65:57:@8503.4]
  assign buffer_3_278 = {{6{_T_59882[4]}},_T_59882}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_279 = {{6{io_in_558[4]}},io_in_558}; // @[Modules.scala 32:22:@8.4]
  assign _T_60485 = $signed(buffer_3_278) + $signed(buffer_3_279); // @[Modules.scala 65:57:@8505.4]
  assign _T_60486 = _T_60485[10:0]; // @[Modules.scala 65:57:@8506.4]
  assign buffer_3_531 = $signed(_T_60486); // @[Modules.scala 65:57:@8507.4]
  assign _T_60488 = $signed(buffer_2_280) + $signed(buffer_1_281); // @[Modules.scala 65:57:@8509.4]
  assign _T_60489 = _T_60488[10:0]; // @[Modules.scala 65:57:@8510.4]
  assign buffer_3_532 = $signed(_T_60489); // @[Modules.scala 65:57:@8511.4]
  assign buffer_3_283 = {{6{_T_59891[4]}},_T_59891}; // @[Modules.scala 32:22:@8.4]
  assign _T_60491 = $signed(buffer_1_282) + $signed(buffer_3_283); // @[Modules.scala 65:57:@8513.4]
  assign _T_60492 = _T_60491[10:0]; // @[Modules.scala 65:57:@8514.4]
  assign buffer_3_533 = $signed(_T_60492); // @[Modules.scala 65:57:@8515.4]
  assign buffer_3_286 = {{6{io_in_572[4]}},io_in_572}; // @[Modules.scala 32:22:@8.4]
  assign _T_60497 = $signed(buffer_3_286) + $signed(buffer_0_287); // @[Modules.scala 65:57:@8521.4]
  assign _T_60498 = _T_60497[10:0]; // @[Modules.scala 65:57:@8522.4]
  assign buffer_3_535 = $signed(_T_60498); // @[Modules.scala 65:57:@8523.4]
  assign _T_60500 = $signed(buffer_1_288) + $signed(buffer_0_289); // @[Modules.scala 65:57:@8525.4]
  assign _T_60501 = _T_60500[10:0]; // @[Modules.scala 65:57:@8526.4]
  assign buffer_3_536 = $signed(_T_60501); // @[Modules.scala 65:57:@8527.4]
  assign buffer_3_291 = {{6{_T_59900[4]}},_T_59900}; // @[Modules.scala 32:22:@8.4]
  assign _T_60503 = $signed(buffer_0_290) + $signed(buffer_3_291); // @[Modules.scala 65:57:@8529.4]
  assign _T_60504 = _T_60503[10:0]; // @[Modules.scala 65:57:@8530.4]
  assign buffer_3_537 = $signed(_T_60504); // @[Modules.scala 65:57:@8531.4]
  assign buffer_3_293 = {{6{_T_59906[4]}},_T_59906}; // @[Modules.scala 32:22:@8.4]
  assign _T_60506 = $signed(buffer_0_292) + $signed(buffer_3_293); // @[Modules.scala 65:57:@8533.4]
  assign _T_60507 = _T_60506[10:0]; // @[Modules.scala 65:57:@8534.4]
  assign buffer_3_538 = $signed(_T_60507); // @[Modules.scala 65:57:@8535.4]
  assign buffer_3_297 = {{6{_T_59916[4]}},_T_59916}; // @[Modules.scala 32:22:@8.4]
  assign _T_60512 = $signed(buffer_1_296) + $signed(buffer_3_297); // @[Modules.scala 65:57:@8541.4]
  assign _T_60513 = _T_60512[10:0]; // @[Modules.scala 65:57:@8542.4]
  assign buffer_3_540 = $signed(_T_60513); // @[Modules.scala 65:57:@8543.4]
  assign _T_60515 = $signed(buffer_1_298) + $signed(11'sh0); // @[Modules.scala 65:57:@8545.4]
  assign _T_60516 = _T_60515[10:0]; // @[Modules.scala 65:57:@8546.4]
  assign buffer_3_541 = $signed(_T_60516); // @[Modules.scala 65:57:@8547.4]
  assign _T_60518 = $signed(buffer_2_300) + $signed(11'sh0); // @[Modules.scala 65:57:@8549.4]
  assign _T_60519 = _T_60518[10:0]; // @[Modules.scala 65:57:@8550.4]
  assign buffer_3_542 = $signed(_T_60519); // @[Modules.scala 65:57:@8551.4]
  assign _T_60521 = $signed(buffer_2_302) + $signed(buffer_0_303); // @[Modules.scala 65:57:@8553.4]
  assign _T_60522 = _T_60521[10:0]; // @[Modules.scala 65:57:@8554.4]
  assign buffer_3_543 = $signed(_T_60522); // @[Modules.scala 65:57:@8555.4]
  assign buffer_3_304 = {{6{io_in_609[4]}},io_in_609}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_305 = {{6{_T_59924[4]}},_T_59924}; // @[Modules.scala 32:22:@8.4]
  assign _T_60524 = $signed(buffer_3_304) + $signed(buffer_3_305); // @[Modules.scala 65:57:@8557.4]
  assign _T_60525 = _T_60524[10:0]; // @[Modules.scala 65:57:@8558.4]
  assign buffer_3_544 = $signed(_T_60525); // @[Modules.scala 65:57:@8559.4]
  assign buffer_3_307 = {{6{io_in_614[4]}},io_in_614}; // @[Modules.scala 32:22:@8.4]
  assign _T_60527 = $signed(buffer_0_306) + $signed(buffer_3_307); // @[Modules.scala 65:57:@8561.4]
  assign _T_60528 = _T_60527[10:0]; // @[Modules.scala 65:57:@8562.4]
  assign buffer_3_545 = $signed(_T_60528); // @[Modules.scala 65:57:@8563.4]
  assign buffer_3_310 = {{6{_T_59934[4]}},_T_59934}; // @[Modules.scala 32:22:@8.4]
  assign _T_60533 = $signed(buffer_3_310) + $signed(11'sh0); // @[Modules.scala 65:57:@8569.4]
  assign _T_60534 = _T_60533[10:0]; // @[Modules.scala 65:57:@8570.4]
  assign buffer_3_547 = $signed(_T_60534); // @[Modules.scala 65:57:@8571.4]
  assign buffer_3_313 = {{6{io_in_627[4]}},io_in_627}; // @[Modules.scala 32:22:@8.4]
  assign _T_60536 = $signed(buffer_1_312) + $signed(buffer_3_313); // @[Modules.scala 65:57:@8573.4]
  assign _T_60537 = _T_60536[10:0]; // @[Modules.scala 65:57:@8574.4]
  assign buffer_3_548 = $signed(_T_60537); // @[Modules.scala 65:57:@8575.4]
  assign buffer_3_315 = {{6{io_in_630[4]}},io_in_630}; // @[Modules.scala 32:22:@8.4]
  assign _T_60539 = $signed(buffer_1_314) + $signed(buffer_3_315); // @[Modules.scala 65:57:@8577.4]
  assign _T_60540 = _T_60539[10:0]; // @[Modules.scala 65:57:@8578.4]
  assign buffer_3_549 = $signed(_T_60540); // @[Modules.scala 65:57:@8579.4]
  assign buffer_3_316 = {{6{io_in_632[4]}},io_in_632}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_317 = {{6{io_in_635[4]}},io_in_635}; // @[Modules.scala 32:22:@8.4]
  assign _T_60542 = $signed(buffer_3_316) + $signed(buffer_3_317); // @[Modules.scala 65:57:@8581.4]
  assign _T_60543 = _T_60542[10:0]; // @[Modules.scala 65:57:@8582.4]
  assign buffer_3_550 = $signed(_T_60543); // @[Modules.scala 65:57:@8583.4]
  assign buffer_3_319 = {{6{_T_59947[4]}},_T_59947}; // @[Modules.scala 32:22:@8.4]
  assign _T_60545 = $signed(buffer_1_318) + $signed(buffer_3_319); // @[Modules.scala 65:57:@8585.4]
  assign _T_60546 = _T_60545[10:0]; // @[Modules.scala 65:57:@8586.4]
  assign buffer_3_551 = $signed(_T_60546); // @[Modules.scala 65:57:@8587.4]
  assign buffer_3_321 = {{6{io_in_642[4]}},io_in_642}; // @[Modules.scala 32:22:@8.4]
  assign _T_60548 = $signed(buffer_0_320) + $signed(buffer_3_321); // @[Modules.scala 65:57:@8589.4]
  assign _T_60549 = _T_60548[10:0]; // @[Modules.scala 65:57:@8590.4]
  assign buffer_3_552 = $signed(_T_60549); // @[Modules.scala 65:57:@8591.4]
  assign _T_60551 = $signed(buffer_2_322) + $signed(buffer_0_323); // @[Modules.scala 65:57:@8593.4]
  assign _T_60552 = _T_60551[10:0]; // @[Modules.scala 65:57:@8594.4]
  assign buffer_3_553 = $signed(_T_60552); // @[Modules.scala 65:57:@8595.4]
  assign buffer_3_325 = {{6{io_in_651[4]}},io_in_651}; // @[Modules.scala 32:22:@8.4]
  assign _T_60554 = $signed(buffer_1_324) + $signed(buffer_3_325); // @[Modules.scala 65:57:@8597.4]
  assign _T_60555 = _T_60554[10:0]; // @[Modules.scala 65:57:@8598.4]
  assign buffer_3_554 = $signed(_T_60555); // @[Modules.scala 65:57:@8599.4]
  assign buffer_3_326 = {{6{io_in_653[4]}},io_in_653}; // @[Modules.scala 32:22:@8.4]
  assign _T_60557 = $signed(buffer_3_326) + $signed(buffer_1_327); // @[Modules.scala 65:57:@8601.4]
  assign _T_60558 = _T_60557[10:0]; // @[Modules.scala 65:57:@8602.4]
  assign buffer_3_555 = $signed(_T_60558); // @[Modules.scala 65:57:@8603.4]
  assign _T_60560 = $signed(buffer_2_328) + $signed(11'sh0); // @[Modules.scala 65:57:@8605.4]
  assign _T_60561 = _T_60560[10:0]; // @[Modules.scala 65:57:@8606.4]
  assign buffer_3_556 = $signed(_T_60561); // @[Modules.scala 65:57:@8607.4]
  assign buffer_3_333 = {{6{io_in_666[4]}},io_in_666}; // @[Modules.scala 32:22:@8.4]
  assign _T_60566 = $signed(11'sh0) + $signed(buffer_3_333); // @[Modules.scala 65:57:@8613.4]
  assign _T_60567 = _T_60566[10:0]; // @[Modules.scala 65:57:@8614.4]
  assign buffer_3_558 = $signed(_T_60567); // @[Modules.scala 65:57:@8615.4]
  assign buffer_3_335 = {{6{io_in_670[4]}},io_in_670}; // @[Modules.scala 32:22:@8.4]
  assign _T_60569 = $signed(buffer_0_334) + $signed(buffer_3_335); // @[Modules.scala 65:57:@8617.4]
  assign _T_60570 = _T_60569[10:0]; // @[Modules.scala 65:57:@8618.4]
  assign buffer_3_559 = $signed(_T_60570); // @[Modules.scala 65:57:@8619.4]
  assign buffer_3_336 = {{6{io_in_672[4]}},io_in_672}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_337 = {{6{io_in_675[4]}},io_in_675}; // @[Modules.scala 32:22:@8.4]
  assign _T_60572 = $signed(buffer_3_336) + $signed(buffer_3_337); // @[Modules.scala 65:57:@8621.4]
  assign _T_60573 = _T_60572[10:0]; // @[Modules.scala 65:57:@8622.4]
  assign buffer_3_560 = $signed(_T_60573); // @[Modules.scala 65:57:@8623.4]
  assign _T_60578 = $signed(buffer_0_340) + $signed(buffer_1_341); // @[Modules.scala 65:57:@8629.4]
  assign _T_60579 = _T_60578[10:0]; // @[Modules.scala 65:57:@8630.4]
  assign buffer_3_562 = $signed(_T_60579); // @[Modules.scala 65:57:@8631.4]
  assign buffer_3_342 = {{6{io_in_685[4]}},io_in_685}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_343 = {{6{_T_59981[4]}},_T_59981}; // @[Modules.scala 32:22:@8.4]
  assign _T_60581 = $signed(buffer_3_342) + $signed(buffer_3_343); // @[Modules.scala 65:57:@8633.4]
  assign _T_60582 = _T_60581[10:0]; // @[Modules.scala 65:57:@8634.4]
  assign buffer_3_563 = $signed(_T_60582); // @[Modules.scala 65:57:@8635.4]
  assign buffer_3_349 = {{6{_T_59989[4]}},_T_59989}; // @[Modules.scala 32:22:@8.4]
  assign _T_60590 = $signed(11'sh0) + $signed(buffer_3_349); // @[Modules.scala 65:57:@8645.4]
  assign _T_60591 = _T_60590[10:0]; // @[Modules.scala 65:57:@8646.4]
  assign buffer_3_566 = $signed(_T_60591); // @[Modules.scala 65:57:@8647.4]
  assign buffer_3_351 = {{6{io_in_703[4]}},io_in_703}; // @[Modules.scala 32:22:@8.4]
  assign _T_60593 = $signed(buffer_0_350) + $signed(buffer_3_351); // @[Modules.scala 65:57:@8649.4]
  assign _T_60594 = _T_60593[10:0]; // @[Modules.scala 65:57:@8650.4]
  assign buffer_3_567 = $signed(_T_60594); // @[Modules.scala 65:57:@8651.4]
  assign buffer_3_355 = {{6{_T_60001[4]}},_T_60001}; // @[Modules.scala 32:22:@8.4]
  assign _T_60599 = $signed(buffer_0_354) + $signed(buffer_3_355); // @[Modules.scala 65:57:@8657.4]
  assign _T_60600 = _T_60599[10:0]; // @[Modules.scala 65:57:@8658.4]
  assign buffer_3_569 = $signed(_T_60600); // @[Modules.scala 65:57:@8659.4]
  assign _T_60611 = $signed(buffer_0_362) + $signed(buffer_1_363); // @[Modules.scala 65:57:@8673.4]
  assign _T_60612 = _T_60611[10:0]; // @[Modules.scala 65:57:@8674.4]
  assign buffer_3_573 = $signed(_T_60612); // @[Modules.scala 65:57:@8675.4]
  assign buffer_3_365 = {{6{io_in_730[4]}},io_in_730}; // @[Modules.scala 32:22:@8.4]
  assign _T_60614 = $signed(buffer_2_364) + $signed(buffer_3_365); // @[Modules.scala 65:57:@8677.4]
  assign _T_60615 = _T_60614[10:0]; // @[Modules.scala 65:57:@8678.4]
  assign buffer_3_574 = $signed(_T_60615); // @[Modules.scala 65:57:@8679.4]
  assign buffer_3_368 = {{6{_T_60022[4]}},_T_60022}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_369 = {{6{_T_60025[4]}},_T_60025}; // @[Modules.scala 32:22:@8.4]
  assign _T_60620 = $signed(buffer_3_368) + $signed(buffer_3_369); // @[Modules.scala 65:57:@8685.4]
  assign _T_60621 = _T_60620[10:0]; // @[Modules.scala 65:57:@8686.4]
  assign buffer_3_576 = $signed(_T_60621); // @[Modules.scala 65:57:@8687.4]
  assign buffer_3_370 = {{6{_T_60028[4]}},_T_60028}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_371 = {{6{io_in_743[4]}},io_in_743}; // @[Modules.scala 32:22:@8.4]
  assign _T_60623 = $signed(buffer_3_370) + $signed(buffer_3_371); // @[Modules.scala 65:57:@8689.4]
  assign _T_60624 = _T_60623[10:0]; // @[Modules.scala 65:57:@8690.4]
  assign buffer_3_577 = $signed(_T_60624); // @[Modules.scala 65:57:@8691.4]
  assign buffer_3_372 = {{6{_T_60031[4]}},_T_60031}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_373 = {{6{_T_60034[4]}},_T_60034}; // @[Modules.scala 32:22:@8.4]
  assign _T_60626 = $signed(buffer_3_372) + $signed(buffer_3_373); // @[Modules.scala 65:57:@8693.4]
  assign _T_60627 = _T_60626[10:0]; // @[Modules.scala 65:57:@8694.4]
  assign buffer_3_578 = $signed(_T_60627); // @[Modules.scala 65:57:@8695.4]
  assign _T_60629 = $signed(11'sh0) + $signed(buffer_0_375); // @[Modules.scala 65:57:@8697.4]
  assign _T_60630 = _T_60629[10:0]; // @[Modules.scala 65:57:@8698.4]
  assign buffer_3_579 = $signed(_T_60630); // @[Modules.scala 65:57:@8699.4]
  assign buffer_3_376 = {{6{io_in_752[4]}},io_in_752}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_377 = {{6{io_in_755[4]}},io_in_755}; // @[Modules.scala 32:22:@8.4]
  assign _T_60632 = $signed(buffer_3_376) + $signed(buffer_3_377); // @[Modules.scala 65:57:@8701.4]
  assign _T_60633 = _T_60632[10:0]; // @[Modules.scala 65:57:@8702.4]
  assign buffer_3_580 = $signed(_T_60633); // @[Modules.scala 65:57:@8703.4]
  assign buffer_3_378 = {{6{_T_60038[4]}},_T_60038}; // @[Modules.scala 32:22:@8.4]
  assign _T_60635 = $signed(buffer_3_378) + $signed(11'sh0); // @[Modules.scala 65:57:@8705.4]
  assign _T_60636 = _T_60635[10:0]; // @[Modules.scala 65:57:@8706.4]
  assign buffer_3_581 = $signed(_T_60636); // @[Modules.scala 65:57:@8707.4]
  assign buffer_3_382 = {{6{_T_60048[4]}},_T_60048}; // @[Modules.scala 32:22:@8.4]
  assign _T_60641 = $signed(buffer_3_382) + $signed(buffer_1_383); // @[Modules.scala 65:57:@8713.4]
  assign _T_60642 = _T_60641[10:0]; // @[Modules.scala 65:57:@8714.4]
  assign buffer_3_583 = $signed(_T_60642); // @[Modules.scala 65:57:@8715.4]
  assign buffer_3_384 = {{6{_T_60054[4]}},_T_60054}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_385 = {{6{_T_60057[4]}},_T_60057}; // @[Modules.scala 32:22:@8.4]
  assign _T_60644 = $signed(buffer_3_384) + $signed(buffer_3_385); // @[Modules.scala 65:57:@8717.4]
  assign _T_60645 = _T_60644[10:0]; // @[Modules.scala 65:57:@8718.4]
  assign buffer_3_584 = $signed(_T_60645); // @[Modules.scala 65:57:@8719.4]
  assign buffer_3_386 = {{6{_T_60060[4]}},_T_60060}; // @[Modules.scala 32:22:@8.4]
  assign buffer_3_387 = {{6{_T_60063[4]}},_T_60063}; // @[Modules.scala 32:22:@8.4]
  assign _T_60647 = $signed(buffer_3_386) + $signed(buffer_3_387); // @[Modules.scala 65:57:@8721.4]
  assign _T_60648 = _T_60647[10:0]; // @[Modules.scala 65:57:@8722.4]
  assign buffer_3_585 = $signed(_T_60648); // @[Modules.scala 65:57:@8723.4]
  assign buffer_3_389 = {{6{io_in_779[4]}},io_in_779}; // @[Modules.scala 32:22:@8.4]
  assign _T_60650 = $signed(11'sh0) + $signed(buffer_3_389); // @[Modules.scala 65:57:@8725.4]
  assign _T_60651 = _T_60650[10:0]; // @[Modules.scala 65:57:@8726.4]
  assign buffer_3_586 = $signed(_T_60651); // @[Modules.scala 65:57:@8727.4]
  assign _T_60653 = $signed(buffer_1_390) + $signed(buffer_0_391); // @[Modules.scala 65:57:@8729.4]
  assign _T_60654 = _T_60653[10:0]; // @[Modules.scala 65:57:@8730.4]
  assign buffer_3_587 = $signed(_T_60654); // @[Modules.scala 65:57:@8731.4]
  assign _T_60656 = $signed(buffer_3_392) + $signed(buffer_1_393); // @[Modules.scala 68:83:@8733.4]
  assign _T_60657 = _T_60656[10:0]; // @[Modules.scala 68:83:@8734.4]
  assign buffer_3_588 = $signed(_T_60657); // @[Modules.scala 68:83:@8735.4]
  assign _T_60659 = $signed(buffer_3_394) + $signed(buffer_1_395); // @[Modules.scala 68:83:@8737.4]
  assign _T_60660 = _T_60659[10:0]; // @[Modules.scala 68:83:@8738.4]
  assign buffer_3_589 = $signed(_T_60660); // @[Modules.scala 68:83:@8739.4]
  assign _T_60662 = $signed(buffer_3_396) + $signed(buffer_3_397); // @[Modules.scala 68:83:@8741.4]
  assign _T_60663 = _T_60662[10:0]; // @[Modules.scala 68:83:@8742.4]
  assign buffer_3_590 = $signed(_T_60663); // @[Modules.scala 68:83:@8743.4]
  assign _T_60665 = $signed(buffer_3_398) + $signed(buffer_3_399); // @[Modules.scala 68:83:@8745.4]
  assign _T_60666 = _T_60665[10:0]; // @[Modules.scala 68:83:@8746.4]
  assign buffer_3_591 = $signed(_T_60666); // @[Modules.scala 68:83:@8747.4]
  assign _T_60668 = $signed(buffer_3_400) + $signed(buffer_1_401); // @[Modules.scala 68:83:@8749.4]
  assign _T_60669 = _T_60668[10:0]; // @[Modules.scala 68:83:@8750.4]
  assign buffer_3_592 = $signed(_T_60669); // @[Modules.scala 68:83:@8751.4]
  assign _T_60671 = $signed(buffer_0_395) + $signed(buffer_3_403); // @[Modules.scala 68:83:@8753.4]
  assign _T_60672 = _T_60671[10:0]; // @[Modules.scala 68:83:@8754.4]
  assign buffer_3_593 = $signed(_T_60672); // @[Modules.scala 68:83:@8755.4]
  assign _T_60674 = $signed(buffer_3_404) + $signed(buffer_3_405); // @[Modules.scala 68:83:@8757.4]
  assign _T_60675 = _T_60674[10:0]; // @[Modules.scala 68:83:@8758.4]
  assign buffer_3_594 = $signed(_T_60675); // @[Modules.scala 68:83:@8759.4]
  assign _T_60677 = $signed(buffer_3_406) + $signed(buffer_3_407); // @[Modules.scala 68:83:@8761.4]
  assign _T_60678 = _T_60677[10:0]; // @[Modules.scala 68:83:@8762.4]
  assign buffer_3_595 = $signed(_T_60678); // @[Modules.scala 68:83:@8763.4]
  assign _T_60686 = $signed(buffer_3_412) + $signed(buffer_3_413); // @[Modules.scala 68:83:@8773.4]
  assign _T_60687 = _T_60686[10:0]; // @[Modules.scala 68:83:@8774.4]
  assign buffer_3_598 = $signed(_T_60687); // @[Modules.scala 68:83:@8775.4]
  assign _T_60689 = $signed(buffer_0_395) + $signed(buffer_3_415); // @[Modules.scala 68:83:@8777.4]
  assign _T_60690 = _T_60689[10:0]; // @[Modules.scala 68:83:@8778.4]
  assign buffer_3_599 = $signed(_T_60690); // @[Modules.scala 68:83:@8779.4]
  assign _T_60692 = $signed(buffer_3_416) + $signed(buffer_3_417); // @[Modules.scala 68:83:@8781.4]
  assign _T_60693 = _T_60692[10:0]; // @[Modules.scala 68:83:@8782.4]
  assign buffer_3_600 = $signed(_T_60693); // @[Modules.scala 68:83:@8783.4]
  assign _T_60695 = $signed(buffer_0_395) + $signed(buffer_3_419); // @[Modules.scala 68:83:@8785.4]
  assign _T_60696 = _T_60695[10:0]; // @[Modules.scala 68:83:@8786.4]
  assign buffer_3_601 = $signed(_T_60696); // @[Modules.scala 68:83:@8787.4]
  assign _T_60698 = $signed(buffer_3_420) + $signed(buffer_3_421); // @[Modules.scala 68:83:@8789.4]
  assign _T_60699 = _T_60698[10:0]; // @[Modules.scala 68:83:@8790.4]
  assign buffer_3_602 = $signed(_T_60699); // @[Modules.scala 68:83:@8791.4]
  assign _T_60701 = $signed(buffer_3_422) + $signed(buffer_3_423); // @[Modules.scala 68:83:@8793.4]
  assign _T_60702 = _T_60701[10:0]; // @[Modules.scala 68:83:@8794.4]
  assign buffer_3_603 = $signed(_T_60702); // @[Modules.scala 68:83:@8795.4]
  assign _T_60704 = $signed(buffer_1_424) + $signed(buffer_3_425); // @[Modules.scala 68:83:@8797.4]
  assign _T_60705 = _T_60704[10:0]; // @[Modules.scala 68:83:@8798.4]
  assign buffer_3_604 = $signed(_T_60705); // @[Modules.scala 68:83:@8799.4]
  assign _T_60707 = $signed(buffer_3_426) + $signed(buffer_3_427); // @[Modules.scala 68:83:@8801.4]
  assign _T_60708 = _T_60707[10:0]; // @[Modules.scala 68:83:@8802.4]
  assign buffer_3_605 = $signed(_T_60708); // @[Modules.scala 68:83:@8803.4]
  assign _T_60710 = $signed(buffer_3_428) + $signed(buffer_3_429); // @[Modules.scala 68:83:@8805.4]
  assign _T_60711 = _T_60710[10:0]; // @[Modules.scala 68:83:@8806.4]
  assign buffer_3_606 = $signed(_T_60711); // @[Modules.scala 68:83:@8807.4]
  assign _T_60713 = $signed(buffer_3_430) + $signed(buffer_3_431); // @[Modules.scala 68:83:@8809.4]
  assign _T_60714 = _T_60713[10:0]; // @[Modules.scala 68:83:@8810.4]
  assign buffer_3_607 = $signed(_T_60714); // @[Modules.scala 68:83:@8811.4]
  assign _T_60719 = $signed(buffer_1_434) + $signed(buffer_3_435); // @[Modules.scala 68:83:@8817.4]
  assign _T_60720 = _T_60719[10:0]; // @[Modules.scala 68:83:@8818.4]
  assign buffer_3_609 = $signed(_T_60720); // @[Modules.scala 68:83:@8819.4]
  assign _T_60722 = $signed(buffer_3_436) + $signed(buffer_3_437); // @[Modules.scala 68:83:@8821.4]
  assign _T_60723 = _T_60722[10:0]; // @[Modules.scala 68:83:@8822.4]
  assign buffer_3_610 = $signed(_T_60723); // @[Modules.scala 68:83:@8823.4]
  assign _T_60725 = $signed(buffer_3_438) + $signed(buffer_3_439); // @[Modules.scala 68:83:@8825.4]
  assign _T_60726 = _T_60725[10:0]; // @[Modules.scala 68:83:@8826.4]
  assign buffer_3_611 = $signed(_T_60726); // @[Modules.scala 68:83:@8827.4]
  assign _T_60728 = $signed(buffer_2_440) + $signed(buffer_3_441); // @[Modules.scala 68:83:@8829.4]
  assign _T_60729 = _T_60728[10:0]; // @[Modules.scala 68:83:@8830.4]
  assign buffer_3_612 = $signed(_T_60729); // @[Modules.scala 68:83:@8831.4]
  assign _T_60731 = $signed(buffer_3_442) + $signed(buffer_3_443); // @[Modules.scala 68:83:@8833.4]
  assign _T_60732 = _T_60731[10:0]; // @[Modules.scala 68:83:@8834.4]
  assign buffer_3_613 = $signed(_T_60732); // @[Modules.scala 68:83:@8835.4]
  assign _T_60734 = $signed(buffer_3_444) + $signed(buffer_3_445); // @[Modules.scala 68:83:@8837.4]
  assign _T_60735 = _T_60734[10:0]; // @[Modules.scala 68:83:@8838.4]
  assign buffer_3_614 = $signed(_T_60735); // @[Modules.scala 68:83:@8839.4]
  assign _T_60737 = $signed(buffer_3_446) + $signed(buffer_2_447); // @[Modules.scala 68:83:@8841.4]
  assign _T_60738 = _T_60737[10:0]; // @[Modules.scala 68:83:@8842.4]
  assign buffer_3_615 = $signed(_T_60738); // @[Modules.scala 68:83:@8843.4]
  assign _T_60740 = $signed(buffer_3_448) + $signed(buffer_3_449); // @[Modules.scala 68:83:@8845.4]
  assign _T_60741 = _T_60740[10:0]; // @[Modules.scala 68:83:@8846.4]
  assign buffer_3_616 = $signed(_T_60741); // @[Modules.scala 68:83:@8847.4]
  assign _T_60743 = $signed(buffer_3_450) + $signed(buffer_3_451); // @[Modules.scala 68:83:@8849.4]
  assign _T_60744 = _T_60743[10:0]; // @[Modules.scala 68:83:@8850.4]
  assign buffer_3_617 = $signed(_T_60744); // @[Modules.scala 68:83:@8851.4]
  assign _T_60746 = $signed(buffer_3_452) + $signed(buffer_3_453); // @[Modules.scala 68:83:@8853.4]
  assign _T_60747 = _T_60746[10:0]; // @[Modules.scala 68:83:@8854.4]
  assign buffer_3_618 = $signed(_T_60747); // @[Modules.scala 68:83:@8855.4]
  assign _T_60749 = $signed(buffer_1_454) + $signed(buffer_3_455); // @[Modules.scala 68:83:@8857.4]
  assign _T_60750 = _T_60749[10:0]; // @[Modules.scala 68:83:@8858.4]
  assign buffer_3_619 = $signed(_T_60750); // @[Modules.scala 68:83:@8859.4]
  assign _T_60752 = $signed(buffer_3_456) + $signed(buffer_2_457); // @[Modules.scala 68:83:@8861.4]
  assign _T_60753 = _T_60752[10:0]; // @[Modules.scala 68:83:@8862.4]
  assign buffer_3_620 = $signed(_T_60753); // @[Modules.scala 68:83:@8863.4]
  assign _T_60755 = $signed(buffer_3_458) + $signed(buffer_3_459); // @[Modules.scala 68:83:@8865.4]
  assign _T_60756 = _T_60755[10:0]; // @[Modules.scala 68:83:@8866.4]
  assign buffer_3_621 = $signed(_T_60756); // @[Modules.scala 68:83:@8867.4]
  assign _T_60758 = $signed(buffer_3_460) + $signed(buffer_1_461); // @[Modules.scala 68:83:@8869.4]
  assign _T_60759 = _T_60758[10:0]; // @[Modules.scala 68:83:@8870.4]
  assign buffer_3_622 = $signed(_T_60759); // @[Modules.scala 68:83:@8871.4]
  assign _T_60761 = $signed(buffer_3_462) + $signed(buffer_3_463); // @[Modules.scala 68:83:@8873.4]
  assign _T_60762 = _T_60761[10:0]; // @[Modules.scala 68:83:@8874.4]
  assign buffer_3_623 = $signed(_T_60762); // @[Modules.scala 68:83:@8875.4]
  assign _T_60764 = $signed(buffer_0_395) + $signed(buffer_3_465); // @[Modules.scala 68:83:@8877.4]
  assign _T_60765 = _T_60764[10:0]; // @[Modules.scala 68:83:@8878.4]
  assign buffer_3_624 = $signed(_T_60765); // @[Modules.scala 68:83:@8879.4]
  assign _T_60767 = $signed(buffer_3_466) + $signed(buffer_3_467); // @[Modules.scala 68:83:@8881.4]
  assign _T_60768 = _T_60767[10:0]; // @[Modules.scala 68:83:@8882.4]
  assign buffer_3_625 = $signed(_T_60768); // @[Modules.scala 68:83:@8883.4]
  assign _T_60770 = $signed(buffer_1_468) + $signed(buffer_3_469); // @[Modules.scala 68:83:@8885.4]
  assign _T_60771 = _T_60770[10:0]; // @[Modules.scala 68:83:@8886.4]
  assign buffer_3_626 = $signed(_T_60771); // @[Modules.scala 68:83:@8887.4]
  assign _T_60779 = $signed(buffer_0_395) + $signed(buffer_3_475); // @[Modules.scala 68:83:@8897.4]
  assign _T_60780 = _T_60779[10:0]; // @[Modules.scala 68:83:@8898.4]
  assign buffer_3_629 = $signed(_T_60780); // @[Modules.scala 68:83:@8899.4]
  assign _T_60782 = $signed(buffer_3_476) + $signed(buffer_0_395); // @[Modules.scala 68:83:@8901.4]
  assign _T_60783 = _T_60782[10:0]; // @[Modules.scala 68:83:@8902.4]
  assign buffer_3_630 = $signed(_T_60783); // @[Modules.scala 68:83:@8903.4]
  assign _T_60791 = $signed(buffer_0_395) + $signed(buffer_3_483); // @[Modules.scala 68:83:@8913.4]
  assign _T_60792 = _T_60791[10:0]; // @[Modules.scala 68:83:@8914.4]
  assign buffer_3_633 = $signed(_T_60792); // @[Modules.scala 68:83:@8915.4]
  assign _T_60794 = $signed(buffer_0_395) + $signed(buffer_3_485); // @[Modules.scala 68:83:@8917.4]
  assign _T_60795 = _T_60794[10:0]; // @[Modules.scala 68:83:@8918.4]
  assign buffer_3_634 = $signed(_T_60795); // @[Modules.scala 68:83:@8919.4]
  assign _T_60797 = $signed(buffer_0_395) + $signed(buffer_3_487); // @[Modules.scala 68:83:@8921.4]
  assign _T_60798 = _T_60797[10:0]; // @[Modules.scala 68:83:@8922.4]
  assign buffer_3_635 = $signed(_T_60798); // @[Modules.scala 68:83:@8923.4]
  assign _T_60800 = $signed(buffer_0_395) + $signed(buffer_3_489); // @[Modules.scala 68:83:@8925.4]
  assign _T_60801 = _T_60800[10:0]; // @[Modules.scala 68:83:@8926.4]
  assign buffer_3_636 = $signed(_T_60801); // @[Modules.scala 68:83:@8927.4]
  assign _T_60803 = $signed(buffer_3_490) + $signed(buffer_0_395); // @[Modules.scala 68:83:@8929.4]
  assign _T_60804 = _T_60803[10:0]; // @[Modules.scala 68:83:@8930.4]
  assign buffer_3_637 = $signed(_T_60804); // @[Modules.scala 68:83:@8931.4]
  assign _T_60806 = $signed(buffer_3_492) + $signed(buffer_0_395); // @[Modules.scala 68:83:@8933.4]
  assign _T_60807 = _T_60806[10:0]; // @[Modules.scala 68:83:@8934.4]
  assign buffer_3_638 = $signed(_T_60807); // @[Modules.scala 68:83:@8935.4]
  assign _T_60809 = $signed(buffer_3_494) + $signed(buffer_0_395); // @[Modules.scala 68:83:@8937.4]
  assign _T_60810 = _T_60809[10:0]; // @[Modules.scala 68:83:@8938.4]
  assign buffer_3_639 = $signed(_T_60810); // @[Modules.scala 68:83:@8939.4]
  assign _T_60812 = $signed(buffer_3_496) + $signed(buffer_3_497); // @[Modules.scala 68:83:@8941.4]
  assign _T_60813 = _T_60812[10:0]; // @[Modules.scala 68:83:@8942.4]
  assign buffer_3_640 = $signed(_T_60813); // @[Modules.scala 68:83:@8943.4]
  assign _T_60815 = $signed(buffer_3_498) + $signed(buffer_2_499); // @[Modules.scala 68:83:@8945.4]
  assign _T_60816 = _T_60815[10:0]; // @[Modules.scala 68:83:@8946.4]
  assign buffer_3_641 = $signed(_T_60816); // @[Modules.scala 68:83:@8947.4]
  assign _T_60821 = $signed(buffer_3_502) + $signed(buffer_3_503); // @[Modules.scala 68:83:@8953.4]
  assign _T_60822 = _T_60821[10:0]; // @[Modules.scala 68:83:@8954.4]
  assign buffer_3_643 = $signed(_T_60822); // @[Modules.scala 68:83:@8955.4]
  assign _T_60824 = $signed(buffer_3_504) + $signed(buffer_3_505); // @[Modules.scala 68:83:@8957.4]
  assign _T_60825 = _T_60824[10:0]; // @[Modules.scala 68:83:@8958.4]
  assign buffer_3_644 = $signed(_T_60825); // @[Modules.scala 68:83:@8959.4]
  assign _T_60830 = $signed(buffer_3_508) + $signed(buffer_1_509); // @[Modules.scala 68:83:@8965.4]
  assign _T_60831 = _T_60830[10:0]; // @[Modules.scala 68:83:@8966.4]
  assign buffer_3_646 = $signed(_T_60831); // @[Modules.scala 68:83:@8967.4]
  assign _T_60833 = $signed(buffer_3_510) + $signed(buffer_3_511); // @[Modules.scala 68:83:@8969.4]
  assign _T_60834 = _T_60833[10:0]; // @[Modules.scala 68:83:@8970.4]
  assign buffer_3_647 = $signed(_T_60834); // @[Modules.scala 68:83:@8971.4]
  assign _T_60836 = $signed(buffer_3_512) + $signed(buffer_0_395); // @[Modules.scala 68:83:@8973.4]
  assign _T_60837 = _T_60836[10:0]; // @[Modules.scala 68:83:@8974.4]
  assign buffer_3_648 = $signed(_T_60837); // @[Modules.scala 68:83:@8975.4]
  assign _T_60839 = $signed(buffer_0_395) + $signed(buffer_3_515); // @[Modules.scala 68:83:@8977.4]
  assign _T_60840 = _T_60839[10:0]; // @[Modules.scala 68:83:@8978.4]
  assign buffer_3_649 = $signed(_T_60840); // @[Modules.scala 68:83:@8979.4]
  assign _T_60842 = $signed(buffer_1_516) + $signed(buffer_3_517); // @[Modules.scala 68:83:@8981.4]
  assign _T_60843 = _T_60842[10:0]; // @[Modules.scala 68:83:@8982.4]
  assign buffer_3_650 = $signed(_T_60843); // @[Modules.scala 68:83:@8983.4]
  assign _T_60845 = $signed(buffer_3_518) + $signed(buffer_3_519); // @[Modules.scala 68:83:@8985.4]
  assign _T_60846 = _T_60845[10:0]; // @[Modules.scala 68:83:@8986.4]
  assign buffer_3_651 = $signed(_T_60846); // @[Modules.scala 68:83:@8987.4]
  assign _T_60851 = $signed(buffer_1_522) + $signed(buffer_0_523); // @[Modules.scala 68:83:@8993.4]
  assign _T_60852 = _T_60851[10:0]; // @[Modules.scala 68:83:@8994.4]
  assign buffer_3_653 = $signed(_T_60852); // @[Modules.scala 68:83:@8995.4]
  assign _T_60854 = $signed(buffer_3_524) + $signed(buffer_1_525); // @[Modules.scala 68:83:@8997.4]
  assign _T_60855 = _T_60854[10:0]; // @[Modules.scala 68:83:@8998.4]
  assign buffer_3_654 = $signed(_T_60855); // @[Modules.scala 68:83:@8999.4]
  assign _T_60857 = $signed(buffer_1_526) + $signed(buffer_3_527); // @[Modules.scala 68:83:@9001.4]
  assign _T_60858 = _T_60857[10:0]; // @[Modules.scala 68:83:@9002.4]
  assign buffer_3_655 = $signed(_T_60858); // @[Modules.scala 68:83:@9003.4]
  assign _T_60860 = $signed(buffer_3_528) + $signed(buffer_0_395); // @[Modules.scala 68:83:@9005.4]
  assign _T_60861 = _T_60860[10:0]; // @[Modules.scala 68:83:@9006.4]
  assign buffer_3_656 = $signed(_T_60861); // @[Modules.scala 68:83:@9007.4]
  assign _T_60863 = $signed(buffer_3_530) + $signed(buffer_3_531); // @[Modules.scala 68:83:@9009.4]
  assign _T_60864 = _T_60863[10:0]; // @[Modules.scala 68:83:@9010.4]
  assign buffer_3_657 = $signed(_T_60864); // @[Modules.scala 68:83:@9011.4]
  assign _T_60866 = $signed(buffer_3_532) + $signed(buffer_3_533); // @[Modules.scala 68:83:@9013.4]
  assign _T_60867 = _T_60866[10:0]; // @[Modules.scala 68:83:@9014.4]
  assign buffer_3_658 = $signed(_T_60867); // @[Modules.scala 68:83:@9015.4]
  assign _T_60869 = $signed(buffer_1_534) + $signed(buffer_3_535); // @[Modules.scala 68:83:@9017.4]
  assign _T_60870 = _T_60869[10:0]; // @[Modules.scala 68:83:@9018.4]
  assign buffer_3_659 = $signed(_T_60870); // @[Modules.scala 68:83:@9019.4]
  assign _T_60872 = $signed(buffer_3_536) + $signed(buffer_3_537); // @[Modules.scala 68:83:@9021.4]
  assign _T_60873 = _T_60872[10:0]; // @[Modules.scala 68:83:@9022.4]
  assign buffer_3_660 = $signed(_T_60873); // @[Modules.scala 68:83:@9023.4]
  assign _T_60875 = $signed(buffer_3_538) + $signed(buffer_1_539); // @[Modules.scala 68:83:@9025.4]
  assign _T_60876 = _T_60875[10:0]; // @[Modules.scala 68:83:@9026.4]
  assign buffer_3_661 = $signed(_T_60876); // @[Modules.scala 68:83:@9027.4]
  assign _T_60878 = $signed(buffer_3_540) + $signed(buffer_3_541); // @[Modules.scala 68:83:@9029.4]
  assign _T_60879 = _T_60878[10:0]; // @[Modules.scala 68:83:@9030.4]
  assign buffer_3_662 = $signed(_T_60879); // @[Modules.scala 68:83:@9031.4]
  assign _T_60881 = $signed(buffer_3_542) + $signed(buffer_3_543); // @[Modules.scala 68:83:@9033.4]
  assign _T_60882 = _T_60881[10:0]; // @[Modules.scala 68:83:@9034.4]
  assign buffer_3_663 = $signed(_T_60882); // @[Modules.scala 68:83:@9035.4]
  assign _T_60884 = $signed(buffer_3_544) + $signed(buffer_3_545); // @[Modules.scala 68:83:@9037.4]
  assign _T_60885 = _T_60884[10:0]; // @[Modules.scala 68:83:@9038.4]
  assign buffer_3_664 = $signed(_T_60885); // @[Modules.scala 68:83:@9039.4]
  assign _T_60887 = $signed(buffer_1_546) + $signed(buffer_3_547); // @[Modules.scala 68:83:@9041.4]
  assign _T_60888 = _T_60887[10:0]; // @[Modules.scala 68:83:@9042.4]
  assign buffer_3_665 = $signed(_T_60888); // @[Modules.scala 68:83:@9043.4]
  assign _T_60890 = $signed(buffer_3_548) + $signed(buffer_3_549); // @[Modules.scala 68:83:@9045.4]
  assign _T_60891 = _T_60890[10:0]; // @[Modules.scala 68:83:@9046.4]
  assign buffer_3_666 = $signed(_T_60891); // @[Modules.scala 68:83:@9047.4]
  assign _T_60893 = $signed(buffer_3_550) + $signed(buffer_3_551); // @[Modules.scala 68:83:@9049.4]
  assign _T_60894 = _T_60893[10:0]; // @[Modules.scala 68:83:@9050.4]
  assign buffer_3_667 = $signed(_T_60894); // @[Modules.scala 68:83:@9051.4]
  assign _T_60896 = $signed(buffer_3_552) + $signed(buffer_3_553); // @[Modules.scala 68:83:@9053.4]
  assign _T_60897 = _T_60896[10:0]; // @[Modules.scala 68:83:@9054.4]
  assign buffer_3_668 = $signed(_T_60897); // @[Modules.scala 68:83:@9055.4]
  assign _T_60899 = $signed(buffer_3_554) + $signed(buffer_3_555); // @[Modules.scala 68:83:@9057.4]
  assign _T_60900 = _T_60899[10:0]; // @[Modules.scala 68:83:@9058.4]
  assign buffer_3_669 = $signed(_T_60900); // @[Modules.scala 68:83:@9059.4]
  assign _T_60902 = $signed(buffer_3_556) + $signed(buffer_0_395); // @[Modules.scala 68:83:@9061.4]
  assign _T_60903 = _T_60902[10:0]; // @[Modules.scala 68:83:@9062.4]
  assign buffer_3_670 = $signed(_T_60903); // @[Modules.scala 68:83:@9063.4]
  assign _T_60905 = $signed(buffer_3_558) + $signed(buffer_3_559); // @[Modules.scala 68:83:@9065.4]
  assign _T_60906 = _T_60905[10:0]; // @[Modules.scala 68:83:@9066.4]
  assign buffer_3_671 = $signed(_T_60906); // @[Modules.scala 68:83:@9067.4]
  assign _T_60908 = $signed(buffer_3_560) + $signed(buffer_0_561); // @[Modules.scala 68:83:@9069.4]
  assign _T_60909 = _T_60908[10:0]; // @[Modules.scala 68:83:@9070.4]
  assign buffer_3_672 = $signed(_T_60909); // @[Modules.scala 68:83:@9071.4]
  assign _T_60911 = $signed(buffer_3_562) + $signed(buffer_3_563); // @[Modules.scala 68:83:@9073.4]
  assign _T_60912 = _T_60911[10:0]; // @[Modules.scala 68:83:@9074.4]
  assign buffer_3_673 = $signed(_T_60912); // @[Modules.scala 68:83:@9075.4]
  assign _T_60917 = $signed(buffer_3_566) + $signed(buffer_3_567); // @[Modules.scala 68:83:@9081.4]
  assign _T_60918 = _T_60917[10:0]; // @[Modules.scala 68:83:@9082.4]
  assign buffer_3_675 = $signed(_T_60918); // @[Modules.scala 68:83:@9083.4]
  assign _T_60920 = $signed(buffer_0_568) + $signed(buffer_3_569); // @[Modules.scala 68:83:@9085.4]
  assign _T_60921 = _T_60920[10:0]; // @[Modules.scala 68:83:@9086.4]
  assign buffer_3_676 = $signed(_T_60921); // @[Modules.scala 68:83:@9087.4]
  assign _T_60923 = $signed(buffer_0_570) + $signed(buffer_1_571); // @[Modules.scala 68:83:@9089.4]
  assign _T_60924 = _T_60923[10:0]; // @[Modules.scala 68:83:@9090.4]
  assign buffer_3_677 = $signed(_T_60924); // @[Modules.scala 68:83:@9091.4]
  assign _T_60926 = $signed(buffer_0_395) + $signed(buffer_3_573); // @[Modules.scala 68:83:@9093.4]
  assign _T_60927 = _T_60926[10:0]; // @[Modules.scala 68:83:@9094.4]
  assign buffer_3_678 = $signed(_T_60927); // @[Modules.scala 68:83:@9095.4]
  assign _T_60929 = $signed(buffer_3_574) + $signed(buffer_0_575); // @[Modules.scala 68:83:@9097.4]
  assign _T_60930 = _T_60929[10:0]; // @[Modules.scala 68:83:@9098.4]
  assign buffer_3_679 = $signed(_T_60930); // @[Modules.scala 68:83:@9099.4]
  assign _T_60932 = $signed(buffer_3_576) + $signed(buffer_3_577); // @[Modules.scala 68:83:@9101.4]
  assign _T_60933 = _T_60932[10:0]; // @[Modules.scala 68:83:@9102.4]
  assign buffer_3_680 = $signed(_T_60933); // @[Modules.scala 68:83:@9103.4]
  assign _T_60935 = $signed(buffer_3_578) + $signed(buffer_3_579); // @[Modules.scala 68:83:@9105.4]
  assign _T_60936 = _T_60935[10:0]; // @[Modules.scala 68:83:@9106.4]
  assign buffer_3_681 = $signed(_T_60936); // @[Modules.scala 68:83:@9107.4]
  assign _T_60938 = $signed(buffer_3_580) + $signed(buffer_3_581); // @[Modules.scala 68:83:@9109.4]
  assign _T_60939 = _T_60938[10:0]; // @[Modules.scala 68:83:@9110.4]
  assign buffer_3_682 = $signed(_T_60939); // @[Modules.scala 68:83:@9111.4]
  assign _T_60941 = $signed(buffer_1_582) + $signed(buffer_3_583); // @[Modules.scala 68:83:@9113.4]
  assign _T_60942 = _T_60941[10:0]; // @[Modules.scala 68:83:@9114.4]
  assign buffer_3_683 = $signed(_T_60942); // @[Modules.scala 68:83:@9115.4]
  assign _T_60944 = $signed(buffer_3_584) + $signed(buffer_3_585); // @[Modules.scala 68:83:@9117.4]
  assign _T_60945 = _T_60944[10:0]; // @[Modules.scala 68:83:@9118.4]
  assign buffer_3_684 = $signed(_T_60945); // @[Modules.scala 68:83:@9119.4]
  assign _T_60947 = $signed(buffer_3_586) + $signed(buffer_3_587); // @[Modules.scala 68:83:@9121.4]
  assign _T_60948 = _T_60947[10:0]; // @[Modules.scala 68:83:@9122.4]
  assign buffer_3_685 = $signed(_T_60948); // @[Modules.scala 68:83:@9123.4]
  assign _T_60950 = $signed(buffer_3_588) + $signed(buffer_3_589); // @[Modules.scala 71:109:@9125.4]
  assign _T_60951 = _T_60950[10:0]; // @[Modules.scala 71:109:@9126.4]
  assign buffer_3_686 = $signed(_T_60951); // @[Modules.scala 71:109:@9127.4]
  assign _T_60953 = $signed(buffer_3_590) + $signed(buffer_3_591); // @[Modules.scala 71:109:@9129.4]
  assign _T_60954 = _T_60953[10:0]; // @[Modules.scala 71:109:@9130.4]
  assign buffer_3_687 = $signed(_T_60954); // @[Modules.scala 71:109:@9131.4]
  assign _T_60956 = $signed(buffer_3_592) + $signed(buffer_3_593); // @[Modules.scala 71:109:@9133.4]
  assign _T_60957 = _T_60956[10:0]; // @[Modules.scala 71:109:@9134.4]
  assign buffer_3_688 = $signed(_T_60957); // @[Modules.scala 71:109:@9135.4]
  assign _T_60959 = $signed(buffer_3_594) + $signed(buffer_3_595); // @[Modules.scala 71:109:@9137.4]
  assign _T_60960 = _T_60959[10:0]; // @[Modules.scala 71:109:@9138.4]
  assign buffer_3_689 = $signed(_T_60960); // @[Modules.scala 71:109:@9139.4]
  assign _T_60965 = $signed(buffer_3_598) + $signed(buffer_3_599); // @[Modules.scala 71:109:@9145.4]
  assign _T_60966 = _T_60965[10:0]; // @[Modules.scala 71:109:@9146.4]
  assign buffer_3_691 = $signed(_T_60966); // @[Modules.scala 71:109:@9147.4]
  assign _T_60968 = $signed(buffer_3_600) + $signed(buffer_3_601); // @[Modules.scala 71:109:@9149.4]
  assign _T_60969 = _T_60968[10:0]; // @[Modules.scala 71:109:@9150.4]
  assign buffer_3_692 = $signed(_T_60969); // @[Modules.scala 71:109:@9151.4]
  assign _T_60971 = $signed(buffer_3_602) + $signed(buffer_3_603); // @[Modules.scala 71:109:@9153.4]
  assign _T_60972 = _T_60971[10:0]; // @[Modules.scala 71:109:@9154.4]
  assign buffer_3_693 = $signed(_T_60972); // @[Modules.scala 71:109:@9155.4]
  assign _T_60974 = $signed(buffer_3_604) + $signed(buffer_3_605); // @[Modules.scala 71:109:@9157.4]
  assign _T_60975 = _T_60974[10:0]; // @[Modules.scala 71:109:@9158.4]
  assign buffer_3_694 = $signed(_T_60975); // @[Modules.scala 71:109:@9159.4]
  assign _T_60977 = $signed(buffer_3_606) + $signed(buffer_3_607); // @[Modules.scala 71:109:@9161.4]
  assign _T_60978 = _T_60977[10:0]; // @[Modules.scala 71:109:@9162.4]
  assign buffer_3_695 = $signed(_T_60978); // @[Modules.scala 71:109:@9163.4]
  assign _T_60980 = $signed(buffer_2_608) + $signed(buffer_3_609); // @[Modules.scala 71:109:@9165.4]
  assign _T_60981 = _T_60980[10:0]; // @[Modules.scala 71:109:@9166.4]
  assign buffer_3_696 = $signed(_T_60981); // @[Modules.scala 71:109:@9167.4]
  assign _T_60983 = $signed(buffer_3_610) + $signed(buffer_3_611); // @[Modules.scala 71:109:@9169.4]
  assign _T_60984 = _T_60983[10:0]; // @[Modules.scala 71:109:@9170.4]
  assign buffer_3_697 = $signed(_T_60984); // @[Modules.scala 71:109:@9171.4]
  assign _T_60986 = $signed(buffer_3_612) + $signed(buffer_3_613); // @[Modules.scala 71:109:@9173.4]
  assign _T_60987 = _T_60986[10:0]; // @[Modules.scala 71:109:@9174.4]
  assign buffer_3_698 = $signed(_T_60987); // @[Modules.scala 71:109:@9175.4]
  assign _T_60989 = $signed(buffer_3_614) + $signed(buffer_3_615); // @[Modules.scala 71:109:@9177.4]
  assign _T_60990 = _T_60989[10:0]; // @[Modules.scala 71:109:@9178.4]
  assign buffer_3_699 = $signed(_T_60990); // @[Modules.scala 71:109:@9179.4]
  assign _T_60992 = $signed(buffer_3_616) + $signed(buffer_3_617); // @[Modules.scala 71:109:@9181.4]
  assign _T_60993 = _T_60992[10:0]; // @[Modules.scala 71:109:@9182.4]
  assign buffer_3_700 = $signed(_T_60993); // @[Modules.scala 71:109:@9183.4]
  assign _T_60995 = $signed(buffer_3_618) + $signed(buffer_3_619); // @[Modules.scala 71:109:@9185.4]
  assign _T_60996 = _T_60995[10:0]; // @[Modules.scala 71:109:@9186.4]
  assign buffer_3_701 = $signed(_T_60996); // @[Modules.scala 71:109:@9187.4]
  assign _T_60998 = $signed(buffer_3_620) + $signed(buffer_3_621); // @[Modules.scala 71:109:@9189.4]
  assign _T_60999 = _T_60998[10:0]; // @[Modules.scala 71:109:@9190.4]
  assign buffer_3_702 = $signed(_T_60999); // @[Modules.scala 71:109:@9191.4]
  assign _T_61001 = $signed(buffer_3_622) + $signed(buffer_3_623); // @[Modules.scala 71:109:@9193.4]
  assign _T_61002 = _T_61001[10:0]; // @[Modules.scala 71:109:@9194.4]
  assign buffer_3_703 = $signed(_T_61002); // @[Modules.scala 71:109:@9195.4]
  assign _T_61004 = $signed(buffer_3_624) + $signed(buffer_3_625); // @[Modules.scala 71:109:@9197.4]
  assign _T_61005 = _T_61004[10:0]; // @[Modules.scala 71:109:@9198.4]
  assign buffer_3_704 = $signed(_T_61005); // @[Modules.scala 71:109:@9199.4]
  assign _T_61007 = $signed(buffer_3_626) + $signed(buffer_0_593); // @[Modules.scala 71:109:@9201.4]
  assign _T_61008 = _T_61007[10:0]; // @[Modules.scala 71:109:@9202.4]
  assign buffer_3_705 = $signed(_T_61008); // @[Modules.scala 71:109:@9203.4]
  assign _T_61010 = $signed(buffer_0_593) + $signed(buffer_3_629); // @[Modules.scala 71:109:@9205.4]
  assign _T_61011 = _T_61010[10:0]; // @[Modules.scala 71:109:@9206.4]
  assign buffer_3_706 = $signed(_T_61011); // @[Modules.scala 71:109:@9207.4]
  assign _T_61013 = $signed(buffer_3_630) + $signed(buffer_0_593); // @[Modules.scala 71:109:@9209.4]
  assign _T_61014 = _T_61013[10:0]; // @[Modules.scala 71:109:@9210.4]
  assign buffer_3_707 = $signed(_T_61014); // @[Modules.scala 71:109:@9211.4]
  assign _T_61016 = $signed(buffer_2_632) + $signed(buffer_3_633); // @[Modules.scala 71:109:@9213.4]
  assign _T_61017 = _T_61016[10:0]; // @[Modules.scala 71:109:@9214.4]
  assign buffer_3_708 = $signed(_T_61017); // @[Modules.scala 71:109:@9215.4]
  assign _T_61019 = $signed(buffer_3_634) + $signed(buffer_3_635); // @[Modules.scala 71:109:@9217.4]
  assign _T_61020 = _T_61019[10:0]; // @[Modules.scala 71:109:@9218.4]
  assign buffer_3_709 = $signed(_T_61020); // @[Modules.scala 71:109:@9219.4]
  assign _T_61022 = $signed(buffer_3_636) + $signed(buffer_3_637); // @[Modules.scala 71:109:@9221.4]
  assign _T_61023 = _T_61022[10:0]; // @[Modules.scala 71:109:@9222.4]
  assign buffer_3_710 = $signed(_T_61023); // @[Modules.scala 71:109:@9223.4]
  assign _T_61025 = $signed(buffer_3_638) + $signed(buffer_3_639); // @[Modules.scala 71:109:@9225.4]
  assign _T_61026 = _T_61025[10:0]; // @[Modules.scala 71:109:@9226.4]
  assign buffer_3_711 = $signed(_T_61026); // @[Modules.scala 71:109:@9227.4]
  assign _T_61028 = $signed(buffer_3_640) + $signed(buffer_3_641); // @[Modules.scala 71:109:@9229.4]
  assign _T_61029 = _T_61028[10:0]; // @[Modules.scala 71:109:@9230.4]
  assign buffer_3_712 = $signed(_T_61029); // @[Modules.scala 71:109:@9231.4]
  assign _T_61031 = $signed(buffer_0_593) + $signed(buffer_3_643); // @[Modules.scala 71:109:@9233.4]
  assign _T_61032 = _T_61031[10:0]; // @[Modules.scala 71:109:@9234.4]
  assign buffer_3_713 = $signed(_T_61032); // @[Modules.scala 71:109:@9235.4]
  assign _T_61034 = $signed(buffer_3_644) + $signed(buffer_0_593); // @[Modules.scala 71:109:@9237.4]
  assign _T_61035 = _T_61034[10:0]; // @[Modules.scala 71:109:@9238.4]
  assign buffer_3_714 = $signed(_T_61035); // @[Modules.scala 71:109:@9239.4]
  assign _T_61037 = $signed(buffer_3_646) + $signed(buffer_3_647); // @[Modules.scala 71:109:@9241.4]
  assign _T_61038 = _T_61037[10:0]; // @[Modules.scala 71:109:@9242.4]
  assign buffer_3_715 = $signed(_T_61038); // @[Modules.scala 71:109:@9243.4]
  assign _T_61040 = $signed(buffer_3_648) + $signed(buffer_3_649); // @[Modules.scala 71:109:@9245.4]
  assign _T_61041 = _T_61040[10:0]; // @[Modules.scala 71:109:@9246.4]
  assign buffer_3_716 = $signed(_T_61041); // @[Modules.scala 71:109:@9247.4]
  assign _T_61043 = $signed(buffer_3_650) + $signed(buffer_3_651); // @[Modules.scala 71:109:@9249.4]
  assign _T_61044 = _T_61043[10:0]; // @[Modules.scala 71:109:@9250.4]
  assign buffer_3_717 = $signed(_T_61044); // @[Modules.scala 71:109:@9251.4]
  assign _T_61046 = $signed(buffer_0_593) + $signed(buffer_3_653); // @[Modules.scala 71:109:@9253.4]
  assign _T_61047 = _T_61046[10:0]; // @[Modules.scala 71:109:@9254.4]
  assign buffer_3_718 = $signed(_T_61047); // @[Modules.scala 71:109:@9255.4]
  assign _T_61049 = $signed(buffer_3_654) + $signed(buffer_3_655); // @[Modules.scala 71:109:@9257.4]
  assign _T_61050 = _T_61049[10:0]; // @[Modules.scala 71:109:@9258.4]
  assign buffer_3_719 = $signed(_T_61050); // @[Modules.scala 71:109:@9259.4]
  assign _T_61052 = $signed(buffer_3_656) + $signed(buffer_3_657); // @[Modules.scala 71:109:@9261.4]
  assign _T_61053 = _T_61052[10:0]; // @[Modules.scala 71:109:@9262.4]
  assign buffer_3_720 = $signed(_T_61053); // @[Modules.scala 71:109:@9263.4]
  assign _T_61055 = $signed(buffer_3_658) + $signed(buffer_3_659); // @[Modules.scala 71:109:@9265.4]
  assign _T_61056 = _T_61055[10:0]; // @[Modules.scala 71:109:@9266.4]
  assign buffer_3_721 = $signed(_T_61056); // @[Modules.scala 71:109:@9267.4]
  assign _T_61058 = $signed(buffer_3_660) + $signed(buffer_3_661); // @[Modules.scala 71:109:@9269.4]
  assign _T_61059 = _T_61058[10:0]; // @[Modules.scala 71:109:@9270.4]
  assign buffer_3_722 = $signed(_T_61059); // @[Modules.scala 71:109:@9271.4]
  assign _T_61061 = $signed(buffer_3_662) + $signed(buffer_3_663); // @[Modules.scala 71:109:@9273.4]
  assign _T_61062 = _T_61061[10:0]; // @[Modules.scala 71:109:@9274.4]
  assign buffer_3_723 = $signed(_T_61062); // @[Modules.scala 71:109:@9275.4]
  assign _T_61064 = $signed(buffer_3_664) + $signed(buffer_3_665); // @[Modules.scala 71:109:@9277.4]
  assign _T_61065 = _T_61064[10:0]; // @[Modules.scala 71:109:@9278.4]
  assign buffer_3_724 = $signed(_T_61065); // @[Modules.scala 71:109:@9279.4]
  assign _T_61067 = $signed(buffer_3_666) + $signed(buffer_3_667); // @[Modules.scala 71:109:@9281.4]
  assign _T_61068 = _T_61067[10:0]; // @[Modules.scala 71:109:@9282.4]
  assign buffer_3_725 = $signed(_T_61068); // @[Modules.scala 71:109:@9283.4]
  assign _T_61070 = $signed(buffer_3_668) + $signed(buffer_3_669); // @[Modules.scala 71:109:@9285.4]
  assign _T_61071 = _T_61070[10:0]; // @[Modules.scala 71:109:@9286.4]
  assign buffer_3_726 = $signed(_T_61071); // @[Modules.scala 71:109:@9287.4]
  assign _T_61073 = $signed(buffer_3_670) + $signed(buffer_3_671); // @[Modules.scala 71:109:@9289.4]
  assign _T_61074 = _T_61073[10:0]; // @[Modules.scala 71:109:@9290.4]
  assign buffer_3_727 = $signed(_T_61074); // @[Modules.scala 71:109:@9291.4]
  assign _T_61076 = $signed(buffer_3_672) + $signed(buffer_3_673); // @[Modules.scala 71:109:@9293.4]
  assign _T_61077 = _T_61076[10:0]; // @[Modules.scala 71:109:@9294.4]
  assign buffer_3_728 = $signed(_T_61077); // @[Modules.scala 71:109:@9295.4]
  assign _T_61079 = $signed(buffer_0_593) + $signed(buffer_3_675); // @[Modules.scala 71:109:@9297.4]
  assign _T_61080 = _T_61079[10:0]; // @[Modules.scala 71:109:@9298.4]
  assign buffer_3_729 = $signed(_T_61080); // @[Modules.scala 71:109:@9299.4]
  assign _T_61082 = $signed(buffer_3_676) + $signed(buffer_3_677); // @[Modules.scala 71:109:@9301.4]
  assign _T_61083 = _T_61082[10:0]; // @[Modules.scala 71:109:@9302.4]
  assign buffer_3_730 = $signed(_T_61083); // @[Modules.scala 71:109:@9303.4]
  assign _T_61085 = $signed(buffer_3_678) + $signed(buffer_3_679); // @[Modules.scala 71:109:@9305.4]
  assign _T_61086 = _T_61085[10:0]; // @[Modules.scala 71:109:@9306.4]
  assign buffer_3_731 = $signed(_T_61086); // @[Modules.scala 71:109:@9307.4]
  assign _T_61088 = $signed(buffer_3_680) + $signed(buffer_3_681); // @[Modules.scala 71:109:@9309.4]
  assign _T_61089 = _T_61088[10:0]; // @[Modules.scala 71:109:@9310.4]
  assign buffer_3_732 = $signed(_T_61089); // @[Modules.scala 71:109:@9311.4]
  assign _T_61091 = $signed(buffer_3_682) + $signed(buffer_3_683); // @[Modules.scala 71:109:@9313.4]
  assign _T_61092 = _T_61091[10:0]; // @[Modules.scala 71:109:@9314.4]
  assign buffer_3_733 = $signed(_T_61092); // @[Modules.scala 71:109:@9315.4]
  assign _T_61094 = $signed(buffer_3_684) + $signed(buffer_3_685); // @[Modules.scala 71:109:@9317.4]
  assign _T_61095 = _T_61094[10:0]; // @[Modules.scala 71:109:@9318.4]
  assign buffer_3_734 = $signed(_T_61095); // @[Modules.scala 71:109:@9319.4]
  assign _T_61097 = $signed(buffer_3_686) + $signed(buffer_3_687); // @[Modules.scala 78:156:@9322.4]
  assign _T_61098 = _T_61097[10:0]; // @[Modules.scala 78:156:@9323.4]
  assign buffer_3_736 = $signed(_T_61098); // @[Modules.scala 78:156:@9324.4]
  assign _T_61100 = $signed(buffer_3_736) + $signed(buffer_3_688); // @[Modules.scala 78:156:@9326.4]
  assign _T_61101 = _T_61100[10:0]; // @[Modules.scala 78:156:@9327.4]
  assign buffer_3_737 = $signed(_T_61101); // @[Modules.scala 78:156:@9328.4]
  assign _T_61103 = $signed(buffer_3_737) + $signed(buffer_3_689); // @[Modules.scala 78:156:@9330.4]
  assign _T_61104 = _T_61103[10:0]; // @[Modules.scala 78:156:@9331.4]
  assign buffer_3_738 = $signed(_T_61104); // @[Modules.scala 78:156:@9332.4]
  assign _T_61106 = $signed(buffer_3_738) + $signed(buffer_0_701); // @[Modules.scala 78:156:@9334.4]
  assign _T_61107 = _T_61106[10:0]; // @[Modules.scala 78:156:@9335.4]
  assign buffer_3_739 = $signed(_T_61107); // @[Modules.scala 78:156:@9336.4]
  assign _T_61109 = $signed(buffer_3_739) + $signed(buffer_3_691); // @[Modules.scala 78:156:@9338.4]
  assign _T_61110 = _T_61109[10:0]; // @[Modules.scala 78:156:@9339.4]
  assign buffer_3_740 = $signed(_T_61110); // @[Modules.scala 78:156:@9340.4]
  assign _T_61112 = $signed(buffer_3_740) + $signed(buffer_3_692); // @[Modules.scala 78:156:@9342.4]
  assign _T_61113 = _T_61112[10:0]; // @[Modules.scala 78:156:@9343.4]
  assign buffer_3_741 = $signed(_T_61113); // @[Modules.scala 78:156:@9344.4]
  assign _T_61115 = $signed(buffer_3_741) + $signed(buffer_3_693); // @[Modules.scala 78:156:@9346.4]
  assign _T_61116 = _T_61115[10:0]; // @[Modules.scala 78:156:@9347.4]
  assign buffer_3_742 = $signed(_T_61116); // @[Modules.scala 78:156:@9348.4]
  assign _T_61118 = $signed(buffer_3_742) + $signed(buffer_3_694); // @[Modules.scala 78:156:@9350.4]
  assign _T_61119 = _T_61118[10:0]; // @[Modules.scala 78:156:@9351.4]
  assign buffer_3_743 = $signed(_T_61119); // @[Modules.scala 78:156:@9352.4]
  assign _T_61121 = $signed(buffer_3_743) + $signed(buffer_3_695); // @[Modules.scala 78:156:@9354.4]
  assign _T_61122 = _T_61121[10:0]; // @[Modules.scala 78:156:@9355.4]
  assign buffer_3_744 = $signed(_T_61122); // @[Modules.scala 78:156:@9356.4]
  assign _T_61124 = $signed(buffer_3_744) + $signed(buffer_3_696); // @[Modules.scala 78:156:@9358.4]
  assign _T_61125 = _T_61124[10:0]; // @[Modules.scala 78:156:@9359.4]
  assign buffer_3_745 = $signed(_T_61125); // @[Modules.scala 78:156:@9360.4]
  assign _T_61127 = $signed(buffer_3_745) + $signed(buffer_3_697); // @[Modules.scala 78:156:@9362.4]
  assign _T_61128 = _T_61127[10:0]; // @[Modules.scala 78:156:@9363.4]
  assign buffer_3_746 = $signed(_T_61128); // @[Modules.scala 78:156:@9364.4]
  assign _T_61130 = $signed(buffer_3_746) + $signed(buffer_3_698); // @[Modules.scala 78:156:@9366.4]
  assign _T_61131 = _T_61130[10:0]; // @[Modules.scala 78:156:@9367.4]
  assign buffer_3_747 = $signed(_T_61131); // @[Modules.scala 78:156:@9368.4]
  assign _T_61133 = $signed(buffer_3_747) + $signed(buffer_3_699); // @[Modules.scala 78:156:@9370.4]
  assign _T_61134 = _T_61133[10:0]; // @[Modules.scala 78:156:@9371.4]
  assign buffer_3_748 = $signed(_T_61134); // @[Modules.scala 78:156:@9372.4]
  assign _T_61136 = $signed(buffer_3_748) + $signed(buffer_3_700); // @[Modules.scala 78:156:@9374.4]
  assign _T_61137 = _T_61136[10:0]; // @[Modules.scala 78:156:@9375.4]
  assign buffer_3_749 = $signed(_T_61137); // @[Modules.scala 78:156:@9376.4]
  assign _T_61139 = $signed(buffer_3_749) + $signed(buffer_3_701); // @[Modules.scala 78:156:@9378.4]
  assign _T_61140 = _T_61139[10:0]; // @[Modules.scala 78:156:@9379.4]
  assign buffer_3_750 = $signed(_T_61140); // @[Modules.scala 78:156:@9380.4]
  assign _T_61142 = $signed(buffer_3_750) + $signed(buffer_3_702); // @[Modules.scala 78:156:@9382.4]
  assign _T_61143 = _T_61142[10:0]; // @[Modules.scala 78:156:@9383.4]
  assign buffer_3_751 = $signed(_T_61143); // @[Modules.scala 78:156:@9384.4]
  assign _T_61145 = $signed(buffer_3_751) + $signed(buffer_3_703); // @[Modules.scala 78:156:@9386.4]
  assign _T_61146 = _T_61145[10:0]; // @[Modules.scala 78:156:@9387.4]
  assign buffer_3_752 = $signed(_T_61146); // @[Modules.scala 78:156:@9388.4]
  assign _T_61148 = $signed(buffer_3_752) + $signed(buffer_3_704); // @[Modules.scala 78:156:@9390.4]
  assign _T_61149 = _T_61148[10:0]; // @[Modules.scala 78:156:@9391.4]
  assign buffer_3_753 = $signed(_T_61149); // @[Modules.scala 78:156:@9392.4]
  assign _T_61151 = $signed(buffer_3_753) + $signed(buffer_3_705); // @[Modules.scala 78:156:@9394.4]
  assign _T_61152 = _T_61151[10:0]; // @[Modules.scala 78:156:@9395.4]
  assign buffer_3_754 = $signed(_T_61152); // @[Modules.scala 78:156:@9396.4]
  assign _T_61154 = $signed(buffer_3_754) + $signed(buffer_3_706); // @[Modules.scala 78:156:@9398.4]
  assign _T_61155 = _T_61154[10:0]; // @[Modules.scala 78:156:@9399.4]
  assign buffer_3_755 = $signed(_T_61155); // @[Modules.scala 78:156:@9400.4]
  assign _T_61157 = $signed(buffer_3_755) + $signed(buffer_3_707); // @[Modules.scala 78:156:@9402.4]
  assign _T_61158 = _T_61157[10:0]; // @[Modules.scala 78:156:@9403.4]
  assign buffer_3_756 = $signed(_T_61158); // @[Modules.scala 78:156:@9404.4]
  assign _T_61160 = $signed(buffer_3_756) + $signed(buffer_3_708); // @[Modules.scala 78:156:@9406.4]
  assign _T_61161 = _T_61160[10:0]; // @[Modules.scala 78:156:@9407.4]
  assign buffer_3_757 = $signed(_T_61161); // @[Modules.scala 78:156:@9408.4]
  assign _T_61163 = $signed(buffer_3_757) + $signed(buffer_3_709); // @[Modules.scala 78:156:@9410.4]
  assign _T_61164 = _T_61163[10:0]; // @[Modules.scala 78:156:@9411.4]
  assign buffer_3_758 = $signed(_T_61164); // @[Modules.scala 78:156:@9412.4]
  assign _T_61166 = $signed(buffer_3_758) + $signed(buffer_3_710); // @[Modules.scala 78:156:@9414.4]
  assign _T_61167 = _T_61166[10:0]; // @[Modules.scala 78:156:@9415.4]
  assign buffer_3_759 = $signed(_T_61167); // @[Modules.scala 78:156:@9416.4]
  assign _T_61169 = $signed(buffer_3_759) + $signed(buffer_3_711); // @[Modules.scala 78:156:@9418.4]
  assign _T_61170 = _T_61169[10:0]; // @[Modules.scala 78:156:@9419.4]
  assign buffer_3_760 = $signed(_T_61170); // @[Modules.scala 78:156:@9420.4]
  assign _T_61172 = $signed(buffer_3_760) + $signed(buffer_3_712); // @[Modules.scala 78:156:@9422.4]
  assign _T_61173 = _T_61172[10:0]; // @[Modules.scala 78:156:@9423.4]
  assign buffer_3_761 = $signed(_T_61173); // @[Modules.scala 78:156:@9424.4]
  assign _T_61175 = $signed(buffer_3_761) + $signed(buffer_3_713); // @[Modules.scala 78:156:@9426.4]
  assign _T_61176 = _T_61175[10:0]; // @[Modules.scala 78:156:@9427.4]
  assign buffer_3_762 = $signed(_T_61176); // @[Modules.scala 78:156:@9428.4]
  assign _T_61178 = $signed(buffer_3_762) + $signed(buffer_3_714); // @[Modules.scala 78:156:@9430.4]
  assign _T_61179 = _T_61178[10:0]; // @[Modules.scala 78:156:@9431.4]
  assign buffer_3_763 = $signed(_T_61179); // @[Modules.scala 78:156:@9432.4]
  assign _T_61181 = $signed(buffer_3_763) + $signed(buffer_3_715); // @[Modules.scala 78:156:@9434.4]
  assign _T_61182 = _T_61181[10:0]; // @[Modules.scala 78:156:@9435.4]
  assign buffer_3_764 = $signed(_T_61182); // @[Modules.scala 78:156:@9436.4]
  assign _T_61184 = $signed(buffer_3_764) + $signed(buffer_3_716); // @[Modules.scala 78:156:@9438.4]
  assign _T_61185 = _T_61184[10:0]; // @[Modules.scala 78:156:@9439.4]
  assign buffer_3_765 = $signed(_T_61185); // @[Modules.scala 78:156:@9440.4]
  assign _T_61187 = $signed(buffer_3_765) + $signed(buffer_3_717); // @[Modules.scala 78:156:@9442.4]
  assign _T_61188 = _T_61187[10:0]; // @[Modules.scala 78:156:@9443.4]
  assign buffer_3_766 = $signed(_T_61188); // @[Modules.scala 78:156:@9444.4]
  assign _T_61190 = $signed(buffer_3_766) + $signed(buffer_3_718); // @[Modules.scala 78:156:@9446.4]
  assign _T_61191 = _T_61190[10:0]; // @[Modules.scala 78:156:@9447.4]
  assign buffer_3_767 = $signed(_T_61191); // @[Modules.scala 78:156:@9448.4]
  assign _T_61193 = $signed(buffer_3_767) + $signed(buffer_3_719); // @[Modules.scala 78:156:@9450.4]
  assign _T_61194 = _T_61193[10:0]; // @[Modules.scala 78:156:@9451.4]
  assign buffer_3_768 = $signed(_T_61194); // @[Modules.scala 78:156:@9452.4]
  assign _T_61196 = $signed(buffer_3_768) + $signed(buffer_3_720); // @[Modules.scala 78:156:@9454.4]
  assign _T_61197 = _T_61196[10:0]; // @[Modules.scala 78:156:@9455.4]
  assign buffer_3_769 = $signed(_T_61197); // @[Modules.scala 78:156:@9456.4]
  assign _T_61199 = $signed(buffer_3_769) + $signed(buffer_3_721); // @[Modules.scala 78:156:@9458.4]
  assign _T_61200 = _T_61199[10:0]; // @[Modules.scala 78:156:@9459.4]
  assign buffer_3_770 = $signed(_T_61200); // @[Modules.scala 78:156:@9460.4]
  assign _T_61202 = $signed(buffer_3_770) + $signed(buffer_3_722); // @[Modules.scala 78:156:@9462.4]
  assign _T_61203 = _T_61202[10:0]; // @[Modules.scala 78:156:@9463.4]
  assign buffer_3_771 = $signed(_T_61203); // @[Modules.scala 78:156:@9464.4]
  assign _T_61205 = $signed(buffer_3_771) + $signed(buffer_3_723); // @[Modules.scala 78:156:@9466.4]
  assign _T_61206 = _T_61205[10:0]; // @[Modules.scala 78:156:@9467.4]
  assign buffer_3_772 = $signed(_T_61206); // @[Modules.scala 78:156:@9468.4]
  assign _T_61208 = $signed(buffer_3_772) + $signed(buffer_3_724); // @[Modules.scala 78:156:@9470.4]
  assign _T_61209 = _T_61208[10:0]; // @[Modules.scala 78:156:@9471.4]
  assign buffer_3_773 = $signed(_T_61209); // @[Modules.scala 78:156:@9472.4]
  assign _T_61211 = $signed(buffer_3_773) + $signed(buffer_3_725); // @[Modules.scala 78:156:@9474.4]
  assign _T_61212 = _T_61211[10:0]; // @[Modules.scala 78:156:@9475.4]
  assign buffer_3_774 = $signed(_T_61212); // @[Modules.scala 78:156:@9476.4]
  assign _T_61214 = $signed(buffer_3_774) + $signed(buffer_3_726); // @[Modules.scala 78:156:@9478.4]
  assign _T_61215 = _T_61214[10:0]; // @[Modules.scala 78:156:@9479.4]
  assign buffer_3_775 = $signed(_T_61215); // @[Modules.scala 78:156:@9480.4]
  assign _T_61217 = $signed(buffer_3_775) + $signed(buffer_3_727); // @[Modules.scala 78:156:@9482.4]
  assign _T_61218 = _T_61217[10:0]; // @[Modules.scala 78:156:@9483.4]
  assign buffer_3_776 = $signed(_T_61218); // @[Modules.scala 78:156:@9484.4]
  assign _T_61220 = $signed(buffer_3_776) + $signed(buffer_3_728); // @[Modules.scala 78:156:@9486.4]
  assign _T_61221 = _T_61220[10:0]; // @[Modules.scala 78:156:@9487.4]
  assign buffer_3_777 = $signed(_T_61221); // @[Modules.scala 78:156:@9488.4]
  assign _T_61223 = $signed(buffer_3_777) + $signed(buffer_3_729); // @[Modules.scala 78:156:@9490.4]
  assign _T_61224 = _T_61223[10:0]; // @[Modules.scala 78:156:@9491.4]
  assign buffer_3_778 = $signed(_T_61224); // @[Modules.scala 78:156:@9492.4]
  assign _T_61226 = $signed(buffer_3_778) + $signed(buffer_3_730); // @[Modules.scala 78:156:@9494.4]
  assign _T_61227 = _T_61226[10:0]; // @[Modules.scala 78:156:@9495.4]
  assign buffer_3_779 = $signed(_T_61227); // @[Modules.scala 78:156:@9496.4]
  assign _T_61229 = $signed(buffer_3_779) + $signed(buffer_3_731); // @[Modules.scala 78:156:@9498.4]
  assign _T_61230 = _T_61229[10:0]; // @[Modules.scala 78:156:@9499.4]
  assign buffer_3_780 = $signed(_T_61230); // @[Modules.scala 78:156:@9500.4]
  assign _T_61232 = $signed(buffer_3_780) + $signed(buffer_3_732); // @[Modules.scala 78:156:@9502.4]
  assign _T_61233 = _T_61232[10:0]; // @[Modules.scala 78:156:@9503.4]
  assign buffer_3_781 = $signed(_T_61233); // @[Modules.scala 78:156:@9504.4]
  assign _T_61235 = $signed(buffer_3_781) + $signed(buffer_3_733); // @[Modules.scala 78:156:@9506.4]
  assign _T_61236 = _T_61235[10:0]; // @[Modules.scala 78:156:@9507.4]
  assign buffer_3_782 = $signed(_T_61236); // @[Modules.scala 78:156:@9508.4]
  assign _T_61238 = $signed(buffer_3_782) + $signed(buffer_3_734); // @[Modules.scala 78:156:@9510.4]
  assign _T_61239 = _T_61238[10:0]; // @[Modules.scala 78:156:@9511.4]
  assign buffer_3_783 = $signed(_T_61239); // @[Modules.scala 78:156:@9512.4]
  assign _T_61268 = $signed(io_in_44) + $signed(io_in_45); // @[Modules.scala 37:46:@9558.4]
  assign _T_61269 = _T_61268[4:0]; // @[Modules.scala 37:46:@9559.4]
  assign _T_61270 = $signed(_T_61269); // @[Modules.scala 37:46:@9560.4]
  assign _T_61361 = $signed(io_in_138) + $signed(io_in_139); // @[Modules.scala 37:46:@9686.4]
  assign _T_61362 = _T_61361[4:0]; // @[Modules.scala 37:46:@9687.4]
  assign _T_61363 = $signed(_T_61362); // @[Modules.scala 37:46:@9688.4]
  assign _T_61365 = $signed(io_in_144) + $signed(io_in_145); // @[Modules.scala 37:46:@9692.4]
  assign _T_61366 = _T_61365[4:0]; // @[Modules.scala 37:46:@9693.4]
  assign _T_61367 = $signed(_T_61366); // @[Modules.scala 37:46:@9694.4]
  assign _T_61377 = $signed(io_in_152) + $signed(io_in_153); // @[Modules.scala 37:46:@9708.4]
  assign _T_61378 = _T_61377[4:0]; // @[Modules.scala 37:46:@9709.4]
  assign _T_61379 = $signed(_T_61378); // @[Modules.scala 37:46:@9710.4]
  assign _T_61383 = $signed(io_in_156) + $signed(io_in_157); // @[Modules.scala 37:46:@9716.4]
  assign _T_61384 = _T_61383[4:0]; // @[Modules.scala 37:46:@9717.4]
  assign _T_61385 = $signed(_T_61384); // @[Modules.scala 37:46:@9718.4]
  assign _T_61395 = $signed(io_in_168) + $signed(io_in_169); // @[Modules.scala 37:46:@9734.4]
  assign _T_61396 = _T_61395[4:0]; // @[Modules.scala 37:46:@9735.4]
  assign _T_61397 = $signed(_T_61396); // @[Modules.scala 37:46:@9736.4]
  assign _T_61413 = $signed(io_in_188) + $signed(io_in_189); // @[Modules.scala 37:46:@9759.4]
  assign _T_61414 = _T_61413[4:0]; // @[Modules.scala 37:46:@9760.4]
  assign _T_61415 = $signed(_T_61414); // @[Modules.scala 37:46:@9761.4]
  assign _T_61447 = $signed(io_in_232) + $signed(io_in_233); // @[Modules.scala 37:46:@9808.4]
  assign _T_61448 = _T_61447[4:0]; // @[Modules.scala 37:46:@9809.4]
  assign _T_61449 = $signed(_T_61448); // @[Modules.scala 37:46:@9810.4]
  assign _T_61456 = $signed(io_in_244) + $signed(io_in_245); // @[Modules.scala 37:46:@9820.4]
  assign _T_61457 = _T_61456[4:0]; // @[Modules.scala 37:46:@9821.4]
  assign _T_61458 = $signed(_T_61457); // @[Modules.scala 37:46:@9822.4]
  assign _T_61470 = $signed(io_in_258) + $signed(io_in_259); // @[Modules.scala 37:46:@9839.4]
  assign _T_61471 = _T_61470[4:0]; // @[Modules.scala 37:46:@9840.4]
  assign _T_61472 = $signed(_T_61471); // @[Modules.scala 37:46:@9841.4]
  assign _T_61473 = $signed(io_in_260) + $signed(io_in_261); // @[Modules.scala 37:46:@9843.4]
  assign _T_61474 = _T_61473[4:0]; // @[Modules.scala 37:46:@9844.4]
  assign _T_61475 = $signed(_T_61474); // @[Modules.scala 37:46:@9845.4]
  assign _T_61496 = $signed(io_in_298) + $signed(io_in_299); // @[Modules.scala 37:46:@9877.4]
  assign _T_61497 = _T_61496[4:0]; // @[Modules.scala 37:46:@9878.4]
  assign _T_61498 = $signed(_T_61497); // @[Modules.scala 37:46:@9879.4]
  assign _T_61500 = $signed(io_in_302) + $signed(io_in_303); // @[Modules.scala 37:46:@9882.4]
  assign _T_61501 = _T_61500[4:0]; // @[Modules.scala 37:46:@9883.4]
  assign _T_61502 = $signed(_T_61501); // @[Modules.scala 37:46:@9884.4]
  assign _T_61554 = $signed(io_in_388) + $signed(io_in_389); // @[Modules.scala 37:46:@9961.4]
  assign _T_61555 = _T_61554[4:0]; // @[Modules.scala 37:46:@9962.4]
  assign _T_61556 = $signed(_T_61555); // @[Modules.scala 37:46:@9963.4]
  assign _T_61570 = $signed(io_in_416) + $signed(io_in_417); // @[Modules.scala 37:46:@9990.4]
  assign _T_61571 = _T_61570[4:0]; // @[Modules.scala 37:46:@9991.4]
  assign _T_61572 = $signed(_T_61571); // @[Modules.scala 37:46:@9992.4]
  assign _T_61573 = $signed(io_in_420) + $signed(io_in_421); // @[Modules.scala 37:46:@9995.4]
  assign _T_61574 = _T_61573[4:0]; // @[Modules.scala 37:46:@9996.4]
  assign _T_61575 = $signed(_T_61574); // @[Modules.scala 37:46:@9997.4]
  assign _T_61635 = $signed(io_in_492) + $signed(io_in_493); // @[Modules.scala 37:46:@10091.4]
  assign _T_61636 = _T_61635[4:0]; // @[Modules.scala 37:46:@10092.4]
  assign _T_61637 = $signed(_T_61636); // @[Modules.scala 37:46:@10093.4]
  assign _T_61686 = $signed(io_in_546) + $signed(io_in_547); // @[Modules.scala 37:46:@10166.4]
  assign _T_61687 = _T_61686[4:0]; // @[Modules.scala 37:46:@10167.4]
  assign _T_61688 = $signed(_T_61687); // @[Modules.scala 37:46:@10168.4]
  assign _T_61729 = $signed(io_in_580) + $signed(io_in_581); // @[Modules.scala 37:46:@10225.4]
  assign _T_61730 = _T_61729[4:0]; // @[Modules.scala 37:46:@10226.4]
  assign _T_61731 = $signed(_T_61730); // @[Modules.scala 37:46:@10227.4]
  assign _T_61766 = $signed(io_in_614) + $signed(io_in_615); // @[Modules.scala 37:46:@10278.4]
  assign _T_61767 = _T_61766[4:0]; // @[Modules.scala 37:46:@10279.4]
  assign _T_61768 = $signed(_T_61767); // @[Modules.scala 37:46:@10280.4]
  assign _T_61775 = $signed(io_in_622) + $signed(io_in_623); // @[Modules.scala 37:46:@10291.4]
  assign _T_61776 = _T_61775[4:0]; // @[Modules.scala 37:46:@10292.4]
  assign _T_61777 = $signed(_T_61776); // @[Modules.scala 37:46:@10293.4]
  assign _T_61821 = $signed(io_in_672) + $signed(io_in_673); // @[Modules.scala 37:46:@10358.4]
  assign _T_61822 = _T_61821[4:0]; // @[Modules.scala 37:46:@10359.4]
  assign _T_61823 = $signed(_T_61822); // @[Modules.scala 37:46:@10360.4]
  assign _T_61861 = $signed(io_in_726) + $signed(io_in_727); // @[Modules.scala 37:46:@10412.4]
  assign _T_61862 = _T_61861[4:0]; // @[Modules.scala 37:46:@10413.4]
  assign _T_61863 = $signed(_T_61862); // @[Modules.scala 37:46:@10414.4]
  assign buffer_4_1 = {{6{io_in_3[4]}},io_in_3}; // @[Modules.scala 32:22:@8.4]
  assign _T_61887 = $signed(buffer_3_0) + $signed(buffer_4_1); // @[Modules.scala 65:57:@10450.4]
  assign _T_61888 = _T_61887[10:0]; // @[Modules.scala 65:57:@10451.4]
  assign buffer_4_392 = $signed(_T_61888); // @[Modules.scala 65:57:@10452.4]
  assign _T_61890 = $signed(buffer_0_2) + $signed(buffer_1_3); // @[Modules.scala 65:57:@10454.4]
  assign _T_61891 = _T_61890[10:0]; // @[Modules.scala 65:57:@10455.4]
  assign buffer_4_393 = $signed(_T_61891); // @[Modules.scala 65:57:@10456.4]
  assign buffer_4_5 = {{6{io_in_11[4]}},io_in_11}; // @[Modules.scala 32:22:@8.4]
  assign _T_61893 = $signed(11'sh0) + $signed(buffer_4_5); // @[Modules.scala 65:57:@10458.4]
  assign _T_61894 = _T_61893[10:0]; // @[Modules.scala 65:57:@10459.4]
  assign buffer_4_394 = $signed(_T_61894); // @[Modules.scala 65:57:@10460.4]
  assign _T_61896 = $signed(11'sh0) + $signed(buffer_1_7); // @[Modules.scala 65:57:@10462.4]
  assign _T_61897 = _T_61896[10:0]; // @[Modules.scala 65:57:@10463.4]
  assign buffer_4_395 = $signed(_T_61897); // @[Modules.scala 65:57:@10464.4]
  assign _T_61899 = $signed(11'sh0) + $signed(buffer_1_9); // @[Modules.scala 65:57:@10466.4]
  assign _T_61900 = _T_61899[10:0]; // @[Modules.scala 65:57:@10467.4]
  assign buffer_4_396 = $signed(_T_61900); // @[Modules.scala 65:57:@10468.4]
  assign _T_61902 = $signed(buffer_0_10) + $signed(11'sh0); // @[Modules.scala 65:57:@10470.4]
  assign _T_61903 = _T_61902[10:0]; // @[Modules.scala 65:57:@10471.4]
  assign buffer_4_397 = $signed(_T_61903); // @[Modules.scala 65:57:@10472.4]
  assign buffer_4_13 = {{6{io_in_27[4]}},io_in_27}; // @[Modules.scala 32:22:@8.4]
  assign _T_61905 = $signed(buffer_3_12) + $signed(buffer_4_13); // @[Modules.scala 65:57:@10474.4]
  assign _T_61906 = _T_61905[10:0]; // @[Modules.scala 65:57:@10475.4]
  assign buffer_4_398 = $signed(_T_61906); // @[Modules.scala 65:57:@10476.4]
  assign buffer_4_14 = {{6{io_in_29[4]}},io_in_29}; // @[Modules.scala 32:22:@8.4]
  assign _T_61908 = $signed(buffer_4_14) + $signed(buffer_2_15); // @[Modules.scala 65:57:@10478.4]
  assign _T_61909 = _T_61908[10:0]; // @[Modules.scala 65:57:@10479.4]
  assign buffer_4_399 = $signed(_T_61909); // @[Modules.scala 65:57:@10480.4]
  assign _T_61917 = $signed(buffer_1_20) + $signed(11'sh0); // @[Modules.scala 65:57:@10490.4]
  assign _T_61918 = _T_61917[10:0]; // @[Modules.scala 65:57:@10491.4]
  assign buffer_4_402 = $signed(_T_61918); // @[Modules.scala 65:57:@10492.4]
  assign buffer_4_22 = {{6{_T_61270[4]}},_T_61270}; // @[Modules.scala 32:22:@8.4]
  assign _T_61920 = $signed(buffer_4_22) + $signed(11'sh0); // @[Modules.scala 65:57:@10494.4]
  assign _T_61921 = _T_61920[10:0]; // @[Modules.scala 65:57:@10495.4]
  assign buffer_4_403 = $signed(_T_61921); // @[Modules.scala 65:57:@10496.4]
  assign _T_61926 = $signed(11'sh0) + $signed(buffer_0_27); // @[Modules.scala 65:57:@10502.4]
  assign _T_61927 = _T_61926[10:0]; // @[Modules.scala 65:57:@10503.4]
  assign buffer_4_405 = $signed(_T_61927); // @[Modules.scala 65:57:@10504.4]
  assign _T_61950 = $signed(buffer_1_42) + $signed(11'sh0); // @[Modules.scala 65:57:@10534.4]
  assign _T_61951 = _T_61950[10:0]; // @[Modules.scala 65:57:@10535.4]
  assign buffer_4_413 = $signed(_T_61951); // @[Modules.scala 65:57:@10536.4]
  assign buffer_4_44 = {{6{io_in_89[4]}},io_in_89}; // @[Modules.scala 32:22:@8.4]
  assign _T_61953 = $signed(buffer_4_44) + $signed(buffer_0_45); // @[Modules.scala 65:57:@10538.4]
  assign _T_61954 = _T_61953[10:0]; // @[Modules.scala 65:57:@10539.4]
  assign buffer_4_414 = $signed(_T_61954); // @[Modules.scala 65:57:@10540.4]
  assign buffer_4_58 = {{6{io_in_117[4]}},io_in_117}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_59 = {{6{io_in_119[4]}},io_in_119}; // @[Modules.scala 32:22:@8.4]
  assign _T_61974 = $signed(buffer_4_58) + $signed(buffer_4_59); // @[Modules.scala 65:57:@10566.4]
  assign _T_61975 = _T_61974[10:0]; // @[Modules.scala 65:57:@10567.4]
  assign buffer_4_421 = $signed(_T_61975); // @[Modules.scala 65:57:@10568.4]
  assign buffer_4_61 = {{6{io_in_122[4]}},io_in_122}; // @[Modules.scala 32:22:@8.4]
  assign _T_61977 = $signed(buffer_3_60) + $signed(buffer_4_61); // @[Modules.scala 65:57:@10570.4]
  assign _T_61978 = _T_61977[10:0]; // @[Modules.scala 65:57:@10571.4]
  assign buffer_4_422 = $signed(_T_61978); // @[Modules.scala 65:57:@10572.4]
  assign _T_61980 = $signed(11'sh0) + $signed(buffer_3_63); // @[Modules.scala 65:57:@10574.4]
  assign _T_61981 = _T_61980[10:0]; // @[Modules.scala 65:57:@10575.4]
  assign buffer_4_423 = $signed(_T_61981); // @[Modules.scala 65:57:@10576.4]
  assign buffer_4_64 = {{6{io_in_128[4]}},io_in_128}; // @[Modules.scala 32:22:@8.4]
  assign _T_61983 = $signed(buffer_4_64) + $signed(11'sh0); // @[Modules.scala 65:57:@10578.4]
  assign _T_61984 = _T_61983[10:0]; // @[Modules.scala 65:57:@10579.4]
  assign buffer_4_424 = $signed(_T_61984); // @[Modules.scala 65:57:@10580.4]
  assign buffer_4_69 = {{6{_T_61363[4]}},_T_61363}; // @[Modules.scala 32:22:@8.4]
  assign _T_61989 = $signed(buffer_1_68) + $signed(buffer_4_69); // @[Modules.scala 65:57:@10586.4]
  assign _T_61990 = _T_61989[10:0]; // @[Modules.scala 65:57:@10587.4]
  assign buffer_4_426 = $signed(_T_61990); // @[Modules.scala 65:57:@10588.4]
  assign _T_61992 = $signed(buffer_2_70) + $signed(11'sh0); // @[Modules.scala 65:57:@10590.4]
  assign _T_61993 = _T_61992[10:0]; // @[Modules.scala 65:57:@10591.4]
  assign buffer_4_427 = $signed(_T_61993); // @[Modules.scala 65:57:@10592.4]
  assign buffer_4_72 = {{6{_T_61367[4]}},_T_61367}; // @[Modules.scala 32:22:@8.4]
  assign _T_61995 = $signed(buffer_4_72) + $signed(buffer_0_73); // @[Modules.scala 65:57:@10594.4]
  assign _T_61996 = _T_61995[10:0]; // @[Modules.scala 65:57:@10595.4]
  assign buffer_4_428 = $signed(_T_61996); // @[Modules.scala 65:57:@10596.4]
  assign buffer_4_76 = {{6{_T_61379[4]}},_T_61379}; // @[Modules.scala 32:22:@8.4]
  assign _T_62001 = $signed(buffer_4_76) + $signed(buffer_3_77); // @[Modules.scala 65:57:@10602.4]
  assign _T_62002 = _T_62001[10:0]; // @[Modules.scala 65:57:@10603.4]
  assign buffer_4_430 = $signed(_T_62002); // @[Modules.scala 65:57:@10604.4]
  assign buffer_4_78 = {{6{_T_61385[4]}},_T_61385}; // @[Modules.scala 32:22:@8.4]
  assign _T_62004 = $signed(buffer_4_78) + $signed(buffer_3_79); // @[Modules.scala 65:57:@10606.4]
  assign _T_62005 = _T_62004[10:0]; // @[Modules.scala 65:57:@10607.4]
  assign buffer_4_431 = $signed(_T_62005); // @[Modules.scala 65:57:@10608.4]
  assign buffer_4_80 = {{6{io_in_160[4]}},io_in_160}; // @[Modules.scala 32:22:@8.4]
  assign _T_62007 = $signed(buffer_4_80) + $signed(buffer_1_81); // @[Modules.scala 65:57:@10610.4]
  assign _T_62008 = _T_62007[10:0]; // @[Modules.scala 65:57:@10611.4]
  assign buffer_4_432 = $signed(_T_62008); // @[Modules.scala 65:57:@10612.4]
  assign buffer_4_84 = {{6{_T_61397[4]}},_T_61397}; // @[Modules.scala 32:22:@8.4]
  assign _T_62013 = $signed(buffer_4_84) + $signed(11'sh0); // @[Modules.scala 65:57:@10618.4]
  assign _T_62014 = _T_62013[10:0]; // @[Modules.scala 65:57:@10619.4]
  assign buffer_4_434 = $signed(_T_62014); // @[Modules.scala 65:57:@10620.4]
  assign buffer_4_92 = {{6{io_in_185[4]}},io_in_185}; // @[Modules.scala 32:22:@8.4]
  assign _T_62025 = $signed(buffer_4_92) + $signed(buffer_0_93); // @[Modules.scala 65:57:@10634.4]
  assign _T_62026 = _T_62025[10:0]; // @[Modules.scala 65:57:@10635.4]
  assign buffer_4_438 = $signed(_T_62026); // @[Modules.scala 65:57:@10636.4]
  assign buffer_4_94 = {{6{_T_61415[4]}},_T_61415}; // @[Modules.scala 32:22:@8.4]
  assign _T_62028 = $signed(buffer_4_94) + $signed(buffer_2_95); // @[Modules.scala 65:57:@10638.4]
  assign _T_62029 = _T_62028[10:0]; // @[Modules.scala 65:57:@10639.4]
  assign buffer_4_439 = $signed(_T_62029); // @[Modules.scala 65:57:@10640.4]
  assign _T_62034 = $signed(buffer_1_98) + $signed(11'sh0); // @[Modules.scala 65:57:@10646.4]
  assign _T_62035 = _T_62034[10:0]; // @[Modules.scala 65:57:@10647.4]
  assign buffer_4_441 = $signed(_T_62035); // @[Modules.scala 65:57:@10648.4]
  assign buffer_4_101 = {{6{io_in_203[4]}},io_in_203}; // @[Modules.scala 32:22:@8.4]
  assign _T_62037 = $signed(buffer_1_100) + $signed(buffer_4_101); // @[Modules.scala 65:57:@10650.4]
  assign _T_62038 = _T_62037[10:0]; // @[Modules.scala 65:57:@10651.4]
  assign buffer_4_442 = $signed(_T_62038); // @[Modules.scala 65:57:@10652.4]
  assign buffer_4_102 = {{6{io_in_204[4]}},io_in_204}; // @[Modules.scala 32:22:@8.4]
  assign _T_62040 = $signed(buffer_4_102) + $signed(buffer_1_103); // @[Modules.scala 65:57:@10654.4]
  assign _T_62041 = _T_62040[10:0]; // @[Modules.scala 65:57:@10655.4]
  assign buffer_4_443 = $signed(_T_62041); // @[Modules.scala 65:57:@10656.4]
  assign buffer_4_114 = {{6{io_in_229[4]}},io_in_229}; // @[Modules.scala 32:22:@8.4]
  assign _T_62058 = $signed(buffer_4_114) + $signed(11'sh0); // @[Modules.scala 65:57:@10678.4]
  assign _T_62059 = _T_62058[10:0]; // @[Modules.scala 65:57:@10679.4]
  assign buffer_4_449 = $signed(_T_62059); // @[Modules.scala 65:57:@10680.4]
  assign buffer_4_116 = {{6{_T_61449[4]}},_T_61449}; // @[Modules.scala 32:22:@8.4]
  assign _T_62061 = $signed(buffer_4_116) + $signed(buffer_3_117); // @[Modules.scala 65:57:@10682.4]
  assign _T_62062 = _T_62061[10:0]; // @[Modules.scala 65:57:@10683.4]
  assign buffer_4_450 = $signed(_T_62062); // @[Modules.scala 65:57:@10684.4]
  assign buffer_4_121 = {{6{io_in_243[4]}},io_in_243}; // @[Modules.scala 32:22:@8.4]
  assign _T_62067 = $signed(11'sh0) + $signed(buffer_4_121); // @[Modules.scala 65:57:@10690.4]
  assign _T_62068 = _T_62067[10:0]; // @[Modules.scala 65:57:@10691.4]
  assign buffer_4_452 = $signed(_T_62068); // @[Modules.scala 65:57:@10692.4]
  assign buffer_4_122 = {{6{_T_61458[4]}},_T_61458}; // @[Modules.scala 32:22:@8.4]
  assign _T_62070 = $signed(buffer_4_122) + $signed(buffer_3_123); // @[Modules.scala 65:57:@10694.4]
  assign _T_62071 = _T_62070[10:0]; // @[Modules.scala 65:57:@10695.4]
  assign buffer_4_453 = $signed(_T_62071); // @[Modules.scala 65:57:@10696.4]
  assign buffer_4_128 = {{6{io_in_257[4]}},io_in_257}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_129 = {{6{_T_61472[4]}},_T_61472}; // @[Modules.scala 32:22:@8.4]
  assign _T_62079 = $signed(buffer_4_128) + $signed(buffer_4_129); // @[Modules.scala 65:57:@10706.4]
  assign _T_62080 = _T_62079[10:0]; // @[Modules.scala 65:57:@10707.4]
  assign buffer_4_456 = $signed(_T_62080); // @[Modules.scala 65:57:@10708.4]
  assign buffer_4_130 = {{6{_T_61475[4]}},_T_61475}; // @[Modules.scala 32:22:@8.4]
  assign _T_62082 = $signed(buffer_4_130) + $signed(buffer_0_131); // @[Modules.scala 65:57:@10710.4]
  assign _T_62083 = _T_62082[10:0]; // @[Modules.scala 65:57:@10711.4]
  assign buffer_4_457 = $signed(_T_62083); // @[Modules.scala 65:57:@10712.4]
  assign _T_62097 = $signed(buffer_1_140) + $signed(11'sh0); // @[Modules.scala 65:57:@10730.4]
  assign _T_62098 = _T_62097[10:0]; // @[Modules.scala 65:57:@10731.4]
  assign buffer_4_462 = $signed(_T_62098); // @[Modules.scala 65:57:@10732.4]
  assign _T_62100 = $signed(buffer_3_142) + $signed(buffer_2_143); // @[Modules.scala 65:57:@10734.4]
  assign _T_62101 = _T_62100[10:0]; // @[Modules.scala 65:57:@10735.4]
  assign buffer_4_463 = $signed(_T_62101); // @[Modules.scala 65:57:@10736.4]
  assign buffer_4_148 = {{6{io_in_297[4]}},io_in_297}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_149 = {{6{_T_61498[4]}},_T_61498}; // @[Modules.scala 32:22:@8.4]
  assign _T_62109 = $signed(buffer_4_148) + $signed(buffer_4_149); // @[Modules.scala 65:57:@10746.4]
  assign _T_62110 = _T_62109[10:0]; // @[Modules.scala 65:57:@10747.4]
  assign buffer_4_466 = $signed(_T_62110); // @[Modules.scala 65:57:@10748.4]
  assign buffer_4_151 = {{6{_T_61502[4]}},_T_61502}; // @[Modules.scala 32:22:@8.4]
  assign _T_62112 = $signed(11'sh0) + $signed(buffer_4_151); // @[Modules.scala 65:57:@10750.4]
  assign _T_62113 = _T_62112[10:0]; // @[Modules.scala 65:57:@10751.4]
  assign buffer_4_467 = $signed(_T_62113); // @[Modules.scala 65:57:@10752.4]
  assign buffer_4_154 = {{6{io_in_308[4]}},io_in_308}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_155 = {{6{io_in_311[4]}},io_in_311}; // @[Modules.scala 32:22:@8.4]
  assign _T_62118 = $signed(buffer_4_154) + $signed(buffer_4_155); // @[Modules.scala 65:57:@10758.4]
  assign _T_62119 = _T_62118[10:0]; // @[Modules.scala 65:57:@10759.4]
  assign buffer_4_469 = $signed(_T_62119); // @[Modules.scala 65:57:@10760.4]
  assign _T_62127 = $signed(buffer_2_160) + $signed(11'sh0); // @[Modules.scala 65:57:@10770.4]
  assign _T_62128 = _T_62127[10:0]; // @[Modules.scala 65:57:@10771.4]
  assign buffer_4_472 = $signed(_T_62128); // @[Modules.scala 65:57:@10772.4]
  assign _T_62136 = $signed(buffer_1_166) + $signed(buffer_3_167); // @[Modules.scala 65:57:@10782.4]
  assign _T_62137 = _T_62136[10:0]; // @[Modules.scala 65:57:@10783.4]
  assign buffer_4_475 = $signed(_T_62137); // @[Modules.scala 65:57:@10784.4]
  assign buffer_4_172 = {{6{io_in_344[4]}},io_in_344}; // @[Modules.scala 32:22:@8.4]
  assign _T_62145 = $signed(buffer_4_172) + $signed(buffer_0_173); // @[Modules.scala 65:57:@10794.4]
  assign _T_62146 = _T_62145[10:0]; // @[Modules.scala 65:57:@10795.4]
  assign buffer_4_478 = $signed(_T_62146); // @[Modules.scala 65:57:@10796.4]
  assign buffer_4_176 = {{6{io_in_352[4]}},io_in_352}; // @[Modules.scala 32:22:@8.4]
  assign _T_62151 = $signed(buffer_4_176) + $signed(11'sh0); // @[Modules.scala 65:57:@10802.4]
  assign _T_62152 = _T_62151[10:0]; // @[Modules.scala 65:57:@10803.4]
  assign buffer_4_480 = $signed(_T_62152); // @[Modules.scala 65:57:@10804.4]
  assign _T_62157 = $signed(buffer_1_180) + $signed(buffer_2_181); // @[Modules.scala 65:57:@10810.4]
  assign _T_62158 = _T_62157[10:0]; // @[Modules.scala 65:57:@10811.4]
  assign buffer_4_482 = $signed(_T_62158); // @[Modules.scala 65:57:@10812.4]
  assign buffer_4_182 = {{6{io_in_364[4]}},io_in_364}; // @[Modules.scala 32:22:@8.4]
  assign _T_62160 = $signed(buffer_4_182) + $signed(11'sh0); // @[Modules.scala 65:57:@10814.4]
  assign _T_62161 = _T_62160[10:0]; // @[Modules.scala 65:57:@10815.4]
  assign buffer_4_483 = $signed(_T_62161); // @[Modules.scala 65:57:@10816.4]
  assign buffer_4_185 = {{6{io_in_370[4]}},io_in_370}; // @[Modules.scala 32:22:@8.4]
  assign _T_62163 = $signed(11'sh0) + $signed(buffer_4_185); // @[Modules.scala 65:57:@10818.4]
  assign _T_62164 = _T_62163[10:0]; // @[Modules.scala 65:57:@10819.4]
  assign buffer_4_484 = $signed(_T_62164); // @[Modules.scala 65:57:@10820.4]
  assign buffer_4_190 = {{6{io_in_380[4]}},io_in_380}; // @[Modules.scala 32:22:@8.4]
  assign _T_62172 = $signed(buffer_4_190) + $signed(11'sh0); // @[Modules.scala 65:57:@10830.4]
  assign _T_62173 = _T_62172[10:0]; // @[Modules.scala 65:57:@10831.4]
  assign buffer_4_487 = $signed(_T_62173); // @[Modules.scala 65:57:@10832.4]
  assign _T_62175 = $signed(11'sh0) + $signed(buffer_0_193); // @[Modules.scala 65:57:@10834.4]
  assign _T_62176 = _T_62175[10:0]; // @[Modules.scala 65:57:@10835.4]
  assign buffer_4_488 = $signed(_T_62176); // @[Modules.scala 65:57:@10836.4]
  assign buffer_4_194 = {{6{_T_61556[4]}},_T_61556}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_195 = {{6{io_in_390[4]}},io_in_390}; // @[Modules.scala 32:22:@8.4]
  assign _T_62178 = $signed(buffer_4_194) + $signed(buffer_4_195); // @[Modules.scala 65:57:@10838.4]
  assign _T_62179 = _T_62178[10:0]; // @[Modules.scala 65:57:@10839.4]
  assign buffer_4_489 = $signed(_T_62179); // @[Modules.scala 65:57:@10840.4]
  assign buffer_4_196 = {{6{io_in_392[4]}},io_in_392}; // @[Modules.scala 32:22:@8.4]
  assign _T_62181 = $signed(buffer_4_196) + $signed(11'sh0); // @[Modules.scala 65:57:@10842.4]
  assign _T_62182 = _T_62181[10:0]; // @[Modules.scala 65:57:@10843.4]
  assign buffer_4_490 = $signed(_T_62182); // @[Modules.scala 65:57:@10844.4]
  assign buffer_4_199 = {{6{io_in_399[4]}},io_in_399}; // @[Modules.scala 32:22:@8.4]
  assign _T_62184 = $signed(buffer_1_198) + $signed(buffer_4_199); // @[Modules.scala 65:57:@10846.4]
  assign _T_62185 = _T_62184[10:0]; // @[Modules.scala 65:57:@10847.4]
  assign buffer_4_491 = $signed(_T_62185); // @[Modules.scala 65:57:@10848.4]
  assign _T_62187 = $signed(buffer_3_200) + $signed(buffer_0_201); // @[Modules.scala 65:57:@10850.4]
  assign _T_62188 = _T_62187[10:0]; // @[Modules.scala 65:57:@10851.4]
  assign buffer_4_492 = $signed(_T_62188); // @[Modules.scala 65:57:@10852.4]
  assign buffer_4_203 = {{6{io_in_407[4]}},io_in_407}; // @[Modules.scala 32:22:@8.4]
  assign _T_62190 = $signed(buffer_0_202) + $signed(buffer_4_203); // @[Modules.scala 65:57:@10854.4]
  assign _T_62191 = _T_62190[10:0]; // @[Modules.scala 65:57:@10855.4]
  assign buffer_4_493 = $signed(_T_62191); // @[Modules.scala 65:57:@10856.4]
  assign _T_62193 = $signed(buffer_0_204) + $signed(buffer_3_205); // @[Modules.scala 65:57:@10858.4]
  assign _T_62194 = _T_62193[10:0]; // @[Modules.scala 65:57:@10859.4]
  assign buffer_4_494 = $signed(_T_62194); // @[Modules.scala 65:57:@10860.4]
  assign buffer_4_206 = {{6{io_in_412[4]}},io_in_412}; // @[Modules.scala 32:22:@8.4]
  assign _T_62196 = $signed(buffer_4_206) + $signed(buffer_0_207); // @[Modules.scala 65:57:@10862.4]
  assign _T_62197 = _T_62196[10:0]; // @[Modules.scala 65:57:@10863.4]
  assign buffer_4_495 = $signed(_T_62197); // @[Modules.scala 65:57:@10864.4]
  assign buffer_4_208 = {{6{_T_61572[4]}},_T_61572}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_209 = {{6{io_in_418[4]}},io_in_418}; // @[Modules.scala 32:22:@8.4]
  assign _T_62199 = $signed(buffer_4_208) + $signed(buffer_4_209); // @[Modules.scala 65:57:@10866.4]
  assign _T_62200 = _T_62199[10:0]; // @[Modules.scala 65:57:@10867.4]
  assign buffer_4_496 = $signed(_T_62200); // @[Modules.scala 65:57:@10868.4]
  assign buffer_4_210 = {{6{_T_61575[4]}},_T_61575}; // @[Modules.scala 32:22:@8.4]
  assign _T_62202 = $signed(buffer_4_210) + $signed(buffer_2_211); // @[Modules.scala 65:57:@10870.4]
  assign _T_62203 = _T_62202[10:0]; // @[Modules.scala 65:57:@10871.4]
  assign buffer_4_497 = $signed(_T_62203); // @[Modules.scala 65:57:@10872.4]
  assign buffer_4_216 = {{6{io_in_432[4]}},io_in_432}; // @[Modules.scala 32:22:@8.4]
  assign _T_62211 = $signed(buffer_4_216) + $signed(buffer_0_217); // @[Modules.scala 65:57:@10882.4]
  assign _T_62212 = _T_62211[10:0]; // @[Modules.scala 65:57:@10883.4]
  assign buffer_4_500 = $signed(_T_62212); // @[Modules.scala 65:57:@10884.4]
  assign buffer_4_218 = {{6{io_in_436[4]}},io_in_436}; // @[Modules.scala 32:22:@8.4]
  assign _T_62214 = $signed(buffer_4_218) + $signed(buffer_1_219); // @[Modules.scala 65:57:@10886.4]
  assign _T_62215 = _T_62214[10:0]; // @[Modules.scala 65:57:@10887.4]
  assign buffer_4_501 = $signed(_T_62215); // @[Modules.scala 65:57:@10888.4]
  assign _T_62217 = $signed(buffer_3_220) + $signed(buffer_1_221); // @[Modules.scala 65:57:@10890.4]
  assign _T_62218 = _T_62217[10:0]; // @[Modules.scala 65:57:@10891.4]
  assign buffer_4_502 = $signed(_T_62218); // @[Modules.scala 65:57:@10892.4]
  assign buffer_4_227 = {{6{io_in_454[4]}},io_in_454}; // @[Modules.scala 32:22:@8.4]
  assign _T_62226 = $signed(buffer_0_226) + $signed(buffer_4_227); // @[Modules.scala 65:57:@10902.4]
  assign _T_62227 = _T_62226[10:0]; // @[Modules.scala 65:57:@10903.4]
  assign buffer_4_505 = $signed(_T_62227); // @[Modules.scala 65:57:@10904.4]
  assign buffer_4_231 = {{6{io_in_463[4]}},io_in_463}; // @[Modules.scala 32:22:@8.4]
  assign _T_62232 = $signed(buffer_2_230) + $signed(buffer_4_231); // @[Modules.scala 65:57:@10910.4]
  assign _T_62233 = _T_62232[10:0]; // @[Modules.scala 65:57:@10911.4]
  assign buffer_4_507 = $signed(_T_62233); // @[Modules.scala 65:57:@10912.4]
  assign _T_62235 = $signed(buffer_2_232) + $signed(buffer_1_233); // @[Modules.scala 65:57:@10914.4]
  assign _T_62236 = _T_62235[10:0]; // @[Modules.scala 65:57:@10915.4]
  assign buffer_4_508 = $signed(_T_62236); // @[Modules.scala 65:57:@10916.4]
  assign _T_62244 = $signed(buffer_2_238) + $signed(buffer_1_239); // @[Modules.scala 65:57:@10926.4]
  assign _T_62245 = _T_62244[10:0]; // @[Modules.scala 65:57:@10927.4]
  assign buffer_4_511 = $signed(_T_62245); // @[Modules.scala 65:57:@10928.4]
  assign _T_62247 = $signed(buffer_3_240) + $signed(buffer_0_241); // @[Modules.scala 65:57:@10930.4]
  assign _T_62248 = _T_62247[10:0]; // @[Modules.scala 65:57:@10931.4]
  assign buffer_4_512 = $signed(_T_62248); // @[Modules.scala 65:57:@10932.4]
  assign buffer_4_243 = {{6{io_in_487[4]}},io_in_487}; // @[Modules.scala 32:22:@8.4]
  assign _T_62250 = $signed(buffer_0_242) + $signed(buffer_4_243); // @[Modules.scala 65:57:@10934.4]
  assign _T_62251 = _T_62250[10:0]; // @[Modules.scala 65:57:@10935.4]
  assign buffer_4_513 = $signed(_T_62251); // @[Modules.scala 65:57:@10936.4]
  assign buffer_4_246 = {{6{_T_61637[4]}},_T_61637}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_247 = {{6{io_in_495[4]}},io_in_495}; // @[Modules.scala 32:22:@8.4]
  assign _T_62256 = $signed(buffer_4_246) + $signed(buffer_4_247); // @[Modules.scala 65:57:@10942.4]
  assign _T_62257 = _T_62256[10:0]; // @[Modules.scala 65:57:@10943.4]
  assign buffer_4_515 = $signed(_T_62257); // @[Modules.scala 65:57:@10944.4]
  assign _T_62265 = $signed(11'sh0) + $signed(buffer_1_253); // @[Modules.scala 65:57:@10954.4]
  assign _T_62266 = _T_62265[10:0]; // @[Modules.scala 65:57:@10955.4]
  assign buffer_4_518 = $signed(_T_62266); // @[Modules.scala 65:57:@10956.4]
  assign buffer_4_256 = {{6{io_in_512[4]}},io_in_512}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_257 = {{6{io_in_514[4]}},io_in_514}; // @[Modules.scala 32:22:@8.4]
  assign _T_62271 = $signed(buffer_4_256) + $signed(buffer_4_257); // @[Modules.scala 65:57:@10962.4]
  assign _T_62272 = _T_62271[10:0]; // @[Modules.scala 65:57:@10963.4]
  assign buffer_4_520 = $signed(_T_62272); // @[Modules.scala 65:57:@10964.4]
  assign buffer_4_259 = {{6{io_in_519[4]}},io_in_519}; // @[Modules.scala 32:22:@8.4]
  assign _T_62274 = $signed(buffer_0_258) + $signed(buffer_4_259); // @[Modules.scala 65:57:@10966.4]
  assign _T_62275 = _T_62274[10:0]; // @[Modules.scala 65:57:@10967.4]
  assign buffer_4_521 = $signed(_T_62275); // @[Modules.scala 65:57:@10968.4]
  assign buffer_4_260 = {{6{io_in_520[4]}},io_in_520}; // @[Modules.scala 32:22:@8.4]
  assign _T_62277 = $signed(buffer_4_260) + $signed(buffer_1_261); // @[Modules.scala 65:57:@10970.4]
  assign _T_62278 = _T_62277[10:0]; // @[Modules.scala 65:57:@10971.4]
  assign buffer_4_522 = $signed(_T_62278); // @[Modules.scala 65:57:@10972.4]
  assign _T_62280 = $signed(buffer_1_262) + $signed(buffer_0_263); // @[Modules.scala 65:57:@10974.4]
  assign _T_62281 = _T_62280[10:0]; // @[Modules.scala 65:57:@10975.4]
  assign buffer_4_523 = $signed(_T_62281); // @[Modules.scala 65:57:@10976.4]
  assign _T_62286 = $signed(11'sh0) + $signed(buffer_0_267); // @[Modules.scala 65:57:@10982.4]
  assign _T_62287 = _T_62286[10:0]; // @[Modules.scala 65:57:@10983.4]
  assign buffer_4_525 = $signed(_T_62287); // @[Modules.scala 65:57:@10984.4]
  assign buffer_4_272 = {{6{io_in_544[4]}},io_in_544}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_273 = {{6{_T_61688[4]}},_T_61688}; // @[Modules.scala 32:22:@8.4]
  assign _T_62295 = $signed(buffer_4_272) + $signed(buffer_4_273); // @[Modules.scala 65:57:@10994.4]
  assign _T_62296 = _T_62295[10:0]; // @[Modules.scala 65:57:@10995.4]
  assign buffer_4_528 = $signed(_T_62296); // @[Modules.scala 65:57:@10996.4]
  assign _T_62304 = $signed(buffer_3_278) + $signed(11'sh0); // @[Modules.scala 65:57:@11006.4]
  assign _T_62305 = _T_62304[10:0]; // @[Modules.scala 65:57:@11007.4]
  assign buffer_4_531 = $signed(_T_62305); // @[Modules.scala 65:57:@11008.4]
  assign _T_62316 = $signed(buffer_1_286) + $signed(buffer_0_287); // @[Modules.scala 65:57:@11022.4]
  assign _T_62317 = _T_62316[10:0]; // @[Modules.scala 65:57:@11023.4]
  assign buffer_4_535 = $signed(_T_62317); // @[Modules.scala 65:57:@11024.4]
  assign buffer_4_290 = {{6{_T_61731[4]}},_T_61731}; // @[Modules.scala 32:22:@8.4]
  assign _T_62322 = $signed(buffer_4_290) + $signed(buffer_3_291); // @[Modules.scala 65:57:@11030.4]
  assign _T_62323 = _T_62322[10:0]; // @[Modules.scala 65:57:@11031.4]
  assign buffer_4_537 = $signed(_T_62323); // @[Modules.scala 65:57:@11032.4]
  assign buffer_4_292 = {{6{io_in_584[4]}},io_in_584}; // @[Modules.scala 32:22:@8.4]
  assign _T_62325 = $signed(buffer_4_292) + $signed(11'sh0); // @[Modules.scala 65:57:@11034.4]
  assign _T_62326 = _T_62325[10:0]; // @[Modules.scala 65:57:@11035.4]
  assign buffer_4_538 = $signed(_T_62326); // @[Modules.scala 65:57:@11036.4]
  assign _T_62328 = $signed(buffer_0_294) + $signed(buffer_1_295); // @[Modules.scala 65:57:@11038.4]
  assign _T_62329 = _T_62328[10:0]; // @[Modules.scala 65:57:@11039.4]
  assign buffer_4_539 = $signed(_T_62329); // @[Modules.scala 65:57:@11040.4]
  assign _T_62334 = $signed(buffer_2_298) + $signed(buffer_1_299); // @[Modules.scala 65:57:@11046.4]
  assign _T_62335 = _T_62334[10:0]; // @[Modules.scala 65:57:@11047.4]
  assign buffer_4_541 = $signed(_T_62335); // @[Modules.scala 65:57:@11048.4]
  assign _T_62343 = $signed(buffer_2_304) + $signed(buffer_3_305); // @[Modules.scala 65:57:@11058.4]
  assign _T_62344 = _T_62343[10:0]; // @[Modules.scala 65:57:@11059.4]
  assign buffer_4_544 = $signed(_T_62344); // @[Modules.scala 65:57:@11060.4]
  assign buffer_4_306 = {{6{io_in_612[4]}},io_in_612}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_307 = {{6{_T_61768[4]}},_T_61768}; // @[Modules.scala 32:22:@8.4]
  assign _T_62346 = $signed(buffer_4_306) + $signed(buffer_4_307); // @[Modules.scala 65:57:@11062.4]
  assign _T_62347 = _T_62346[10:0]; // @[Modules.scala 65:57:@11063.4]
  assign buffer_4_545 = $signed(_T_62347); // @[Modules.scala 65:57:@11064.4]
  assign buffer_4_311 = {{6{_T_61777[4]}},_T_61777}; // @[Modules.scala 32:22:@8.4]
  assign _T_62352 = $signed(buffer_3_310) + $signed(buffer_4_311); // @[Modules.scala 65:57:@11070.4]
  assign _T_62353 = _T_62352[10:0]; // @[Modules.scala 65:57:@11071.4]
  assign buffer_4_547 = $signed(_T_62353); // @[Modules.scala 65:57:@11072.4]
  assign _T_62355 = $signed(11'sh0) + $signed(buffer_1_313); // @[Modules.scala 65:57:@11074.4]
  assign _T_62356 = _T_62355[10:0]; // @[Modules.scala 65:57:@11075.4]
  assign buffer_4_548 = $signed(_T_62356); // @[Modules.scala 65:57:@11076.4]
  assign buffer_4_316 = {{6{io_in_633[4]}},io_in_633}; // @[Modules.scala 32:22:@8.4]
  assign _T_62361 = $signed(buffer_4_316) + $signed(buffer_2_317); // @[Modules.scala 65:57:@11082.4]
  assign _T_62362 = _T_62361[10:0]; // @[Modules.scala 65:57:@11083.4]
  assign buffer_4_550 = $signed(_T_62362); // @[Modules.scala 65:57:@11084.4]
  assign _T_62367 = $signed(11'sh0) + $signed(buffer_0_321); // @[Modules.scala 65:57:@11090.4]
  assign _T_62368 = _T_62367[10:0]; // @[Modules.scala 65:57:@11091.4]
  assign buffer_4_552 = $signed(_T_62368); // @[Modules.scala 65:57:@11092.4]
  assign buffer_4_324 = {{6{io_in_648[4]}},io_in_648}; // @[Modules.scala 32:22:@8.4]
  assign _T_62373 = $signed(buffer_4_324) + $signed(11'sh0); // @[Modules.scala 65:57:@11098.4]
  assign _T_62374 = _T_62373[10:0]; // @[Modules.scala 65:57:@11099.4]
  assign buffer_4_554 = $signed(_T_62374); // @[Modules.scala 65:57:@11100.4]
  assign buffer_4_330 = {{6{io_in_660[4]}},io_in_660}; // @[Modules.scala 32:22:@8.4]
  assign _T_62382 = $signed(buffer_4_330) + $signed(buffer_1_331); // @[Modules.scala 65:57:@11110.4]
  assign _T_62383 = _T_62382[10:0]; // @[Modules.scala 65:57:@11111.4]
  assign buffer_4_557 = $signed(_T_62383); // @[Modules.scala 65:57:@11112.4]
  assign _T_62385 = $signed(buffer_0_332) + $signed(11'sh0); // @[Modules.scala 65:57:@11114.4]
  assign _T_62386 = _T_62385[10:0]; // @[Modules.scala 65:57:@11115.4]
  assign buffer_4_558 = $signed(_T_62386); // @[Modules.scala 65:57:@11116.4]
  assign buffer_4_334 = {{6{io_in_669[4]}},io_in_669}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_335 = {{6{io_in_671[4]}},io_in_671}; // @[Modules.scala 32:22:@8.4]
  assign _T_62388 = $signed(buffer_4_334) + $signed(buffer_4_335); // @[Modules.scala 65:57:@11118.4]
  assign _T_62389 = _T_62388[10:0]; // @[Modules.scala 65:57:@11119.4]
  assign buffer_4_559 = $signed(_T_62389); // @[Modules.scala 65:57:@11120.4]
  assign buffer_4_336 = {{6{_T_61823[4]}},_T_61823}; // @[Modules.scala 32:22:@8.4]
  assign _T_62391 = $signed(buffer_4_336) + $signed(buffer_1_337); // @[Modules.scala 65:57:@11122.4]
  assign _T_62392 = _T_62391[10:0]; // @[Modules.scala 65:57:@11123.4]
  assign buffer_4_560 = $signed(_T_62392); // @[Modules.scala 65:57:@11124.4]
  assign buffer_4_338 = {{6{io_in_676[4]}},io_in_676}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_339 = {{6{io_in_679[4]}},io_in_679}; // @[Modules.scala 32:22:@8.4]
  assign _T_62394 = $signed(buffer_4_338) + $signed(buffer_4_339); // @[Modules.scala 65:57:@11126.4]
  assign _T_62395 = _T_62394[10:0]; // @[Modules.scala 65:57:@11127.4]
  assign buffer_4_561 = $signed(_T_62395); // @[Modules.scala 65:57:@11128.4]
  assign _T_62400 = $signed(buffer_1_342) + $signed(buffer_3_343); // @[Modules.scala 65:57:@11134.4]
  assign _T_62401 = _T_62400[10:0]; // @[Modules.scala 65:57:@11135.4]
  assign buffer_4_563 = $signed(_T_62401); // @[Modules.scala 65:57:@11136.4]
  assign _T_62403 = $signed(buffer_0_344) + $signed(11'sh0); // @[Modules.scala 65:57:@11138.4]
  assign _T_62404 = _T_62403[10:0]; // @[Modules.scala 65:57:@11139.4]
  assign buffer_4_564 = $signed(_T_62404); // @[Modules.scala 65:57:@11140.4]
  assign buffer_4_348 = {{6{io_in_697[4]}},io_in_697}; // @[Modules.scala 32:22:@8.4]
  assign buffer_4_349 = {{6{io_in_698[4]}},io_in_698}; // @[Modules.scala 32:22:@8.4]
  assign _T_62409 = $signed(buffer_4_348) + $signed(buffer_4_349); // @[Modules.scala 65:57:@11146.4]
  assign _T_62410 = _T_62409[10:0]; // @[Modules.scala 65:57:@11147.4]
  assign buffer_4_566 = $signed(_T_62410); // @[Modules.scala 65:57:@11148.4]
  assign buffer_4_352 = {{6{io_in_704[4]}},io_in_704}; // @[Modules.scala 32:22:@8.4]
  assign _T_62415 = $signed(buffer_4_352) + $signed(11'sh0); // @[Modules.scala 65:57:@11154.4]
  assign _T_62416 = _T_62415[10:0]; // @[Modules.scala 65:57:@11155.4]
  assign buffer_4_568 = $signed(_T_62416); // @[Modules.scala 65:57:@11156.4]
  assign buffer_4_363 = {{6{_T_61863[4]}},_T_61863}; // @[Modules.scala 32:22:@8.4]
  assign _T_62430 = $signed(11'sh0) + $signed(buffer_4_363); // @[Modules.scala 65:57:@11174.4]
  assign _T_62431 = _T_62430[10:0]; // @[Modules.scala 65:57:@11175.4]
  assign buffer_4_573 = $signed(_T_62431); // @[Modules.scala 65:57:@11176.4]
  assign buffer_4_376 = {{6{io_in_753[4]}},io_in_753}; // @[Modules.scala 32:22:@8.4]
  assign _T_62451 = $signed(buffer_4_376) + $signed(buffer_3_377); // @[Modules.scala 65:57:@11202.4]
  assign _T_62452 = _T_62451[10:0]; // @[Modules.scala 65:57:@11203.4]
  assign buffer_4_580 = $signed(_T_62452); // @[Modules.scala 65:57:@11204.4]
  assign _T_62454 = $signed(buffer_1_378) + $signed(11'sh0); // @[Modules.scala 65:57:@11206.4]
  assign _T_62455 = _T_62454[10:0]; // @[Modules.scala 65:57:@11207.4]
  assign buffer_4_581 = $signed(_T_62455); // @[Modules.scala 65:57:@11208.4]
  assign _T_62457 = $signed(buffer_1_380) + $signed(11'sh0); // @[Modules.scala 65:57:@11210.4]
  assign _T_62458 = _T_62457[10:0]; // @[Modules.scala 65:57:@11211.4]
  assign buffer_4_582 = $signed(_T_62458); // @[Modules.scala 65:57:@11212.4]
  assign buffer_4_383 = {{6{io_in_767[4]}},io_in_767}; // @[Modules.scala 32:22:@8.4]
  assign _T_62460 = $signed(11'sh0) + $signed(buffer_4_383); // @[Modules.scala 65:57:@11214.4]
  assign _T_62461 = _T_62460[10:0]; // @[Modules.scala 65:57:@11215.4]
  assign buffer_4_583 = $signed(_T_62461); // @[Modules.scala 65:57:@11216.4]
  assign _T_62463 = $signed(buffer_0_384) + $signed(11'sh0); // @[Modules.scala 65:57:@11218.4]
  assign _T_62464 = _T_62463[10:0]; // @[Modules.scala 65:57:@11219.4]
  assign buffer_4_584 = $signed(_T_62464); // @[Modules.scala 65:57:@11220.4]
  assign buffer_4_386 = {{6{io_in_772[4]}},io_in_772}; // @[Modules.scala 32:22:@8.4]
  assign _T_62466 = $signed(buffer_4_386) + $signed(11'sh0); // @[Modules.scala 65:57:@11222.4]
  assign _T_62467 = _T_62466[10:0]; // @[Modules.scala 65:57:@11223.4]
  assign buffer_4_585 = $signed(_T_62467); // @[Modules.scala 65:57:@11224.4]
  assign _T_62472 = $signed(11'sh0) + $signed(buffer_2_391); // @[Modules.scala 65:57:@11230.4]
  assign _T_62473 = _T_62472[10:0]; // @[Modules.scala 65:57:@11231.4]
  assign buffer_4_587 = $signed(_T_62473); // @[Modules.scala 65:57:@11232.4]
  assign _T_62475 = $signed(buffer_4_392) + $signed(buffer_4_393); // @[Modules.scala 68:83:@11234.4]
  assign _T_62476 = _T_62475[10:0]; // @[Modules.scala 68:83:@11235.4]
  assign buffer_4_588 = $signed(_T_62476); // @[Modules.scala 68:83:@11236.4]
  assign _T_62478 = $signed(buffer_4_394) + $signed(buffer_4_395); // @[Modules.scala 68:83:@11238.4]
  assign _T_62479 = _T_62478[10:0]; // @[Modules.scala 68:83:@11239.4]
  assign buffer_4_589 = $signed(_T_62479); // @[Modules.scala 68:83:@11240.4]
  assign _T_62481 = $signed(buffer_4_396) + $signed(buffer_4_397); // @[Modules.scala 68:83:@11242.4]
  assign _T_62482 = _T_62481[10:0]; // @[Modules.scala 68:83:@11243.4]
  assign buffer_4_590 = $signed(_T_62482); // @[Modules.scala 68:83:@11244.4]
  assign _T_62484 = $signed(buffer_4_398) + $signed(buffer_4_399); // @[Modules.scala 68:83:@11246.4]
  assign _T_62485 = _T_62484[10:0]; // @[Modules.scala 68:83:@11247.4]
  assign buffer_4_591 = $signed(_T_62485); // @[Modules.scala 68:83:@11248.4]
  assign _T_62487 = $signed(buffer_0_400) + $signed(buffer_1_401); // @[Modules.scala 68:83:@11250.4]
  assign _T_62488 = _T_62487[10:0]; // @[Modules.scala 68:83:@11251.4]
  assign buffer_4_592 = $signed(_T_62488); // @[Modules.scala 68:83:@11252.4]
  assign _T_62490 = $signed(buffer_4_402) + $signed(buffer_4_403); // @[Modules.scala 68:83:@11254.4]
  assign _T_62491 = _T_62490[10:0]; // @[Modules.scala 68:83:@11255.4]
  assign buffer_4_593 = $signed(_T_62491); // @[Modules.scala 68:83:@11256.4]
  assign _T_62493 = $signed(buffer_1_404) + $signed(buffer_4_405); // @[Modules.scala 68:83:@11258.4]
  assign _T_62494 = _T_62493[10:0]; // @[Modules.scala 68:83:@11259.4]
  assign buffer_4_594 = $signed(_T_62494); // @[Modules.scala 68:83:@11260.4]
  assign _T_62496 = $signed(buffer_2_406) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11262.4]
  assign _T_62497 = _T_62496[10:0]; // @[Modules.scala 68:83:@11263.4]
  assign buffer_4_595 = $signed(_T_62497); // @[Modules.scala 68:83:@11264.4]
  assign _T_62505 = $signed(buffer_2_412) + $signed(buffer_4_413); // @[Modules.scala 68:83:@11274.4]
  assign _T_62506 = _T_62505[10:0]; // @[Modules.scala 68:83:@11275.4]
  assign buffer_4_598 = $signed(_T_62506); // @[Modules.scala 68:83:@11276.4]
  assign _T_62508 = $signed(buffer_4_414) + $signed(buffer_1_415); // @[Modules.scala 68:83:@11278.4]
  assign _T_62509 = _T_62508[10:0]; // @[Modules.scala 68:83:@11279.4]
  assign buffer_4_599 = $signed(_T_62509); // @[Modules.scala 68:83:@11280.4]
  assign _T_62517 = $signed(buffer_0_395) + $signed(buffer_4_421); // @[Modules.scala 68:83:@11290.4]
  assign _T_62518 = _T_62517[10:0]; // @[Modules.scala 68:83:@11291.4]
  assign buffer_4_602 = $signed(_T_62518); // @[Modules.scala 68:83:@11292.4]
  assign _T_62520 = $signed(buffer_4_422) + $signed(buffer_4_423); // @[Modules.scala 68:83:@11294.4]
  assign _T_62521 = _T_62520[10:0]; // @[Modules.scala 68:83:@11295.4]
  assign buffer_4_603 = $signed(_T_62521); // @[Modules.scala 68:83:@11296.4]
  assign _T_62523 = $signed(buffer_4_424) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11298.4]
  assign _T_62524 = _T_62523[10:0]; // @[Modules.scala 68:83:@11299.4]
  assign buffer_4_604 = $signed(_T_62524); // @[Modules.scala 68:83:@11300.4]
  assign _T_62526 = $signed(buffer_4_426) + $signed(buffer_4_427); // @[Modules.scala 68:83:@11302.4]
  assign _T_62527 = _T_62526[10:0]; // @[Modules.scala 68:83:@11303.4]
  assign buffer_4_605 = $signed(_T_62527); // @[Modules.scala 68:83:@11304.4]
  assign _T_62529 = $signed(buffer_4_428) + $signed(buffer_3_429); // @[Modules.scala 68:83:@11306.4]
  assign _T_62530 = _T_62529[10:0]; // @[Modules.scala 68:83:@11307.4]
  assign buffer_4_606 = $signed(_T_62530); // @[Modules.scala 68:83:@11308.4]
  assign _T_62532 = $signed(buffer_4_430) + $signed(buffer_4_431); // @[Modules.scala 68:83:@11310.4]
  assign _T_62533 = _T_62532[10:0]; // @[Modules.scala 68:83:@11311.4]
  assign buffer_4_607 = $signed(_T_62533); // @[Modules.scala 68:83:@11312.4]
  assign _T_62535 = $signed(buffer_4_432) + $signed(buffer_2_433); // @[Modules.scala 68:83:@11314.4]
  assign _T_62536 = _T_62535[10:0]; // @[Modules.scala 68:83:@11315.4]
  assign buffer_4_608 = $signed(_T_62536); // @[Modules.scala 68:83:@11316.4]
  assign _T_62538 = $signed(buffer_4_434) + $signed(buffer_3_435); // @[Modules.scala 68:83:@11318.4]
  assign _T_62539 = _T_62538[10:0]; // @[Modules.scala 68:83:@11319.4]
  assign buffer_4_609 = $signed(_T_62539); // @[Modules.scala 68:83:@11320.4]
  assign _T_62541 = $signed(buffer_1_436) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11322.4]
  assign _T_62542 = _T_62541[10:0]; // @[Modules.scala 68:83:@11323.4]
  assign buffer_4_610 = $signed(_T_62542); // @[Modules.scala 68:83:@11324.4]
  assign _T_62544 = $signed(buffer_4_438) + $signed(buffer_4_439); // @[Modules.scala 68:83:@11326.4]
  assign _T_62545 = _T_62544[10:0]; // @[Modules.scala 68:83:@11327.4]
  assign buffer_4_611 = $signed(_T_62545); // @[Modules.scala 68:83:@11328.4]
  assign _T_62547 = $signed(buffer_2_440) + $signed(buffer_4_441); // @[Modules.scala 68:83:@11330.4]
  assign _T_62548 = _T_62547[10:0]; // @[Modules.scala 68:83:@11331.4]
  assign buffer_4_612 = $signed(_T_62548); // @[Modules.scala 68:83:@11332.4]
  assign _T_62550 = $signed(buffer_4_442) + $signed(buffer_4_443); // @[Modules.scala 68:83:@11334.4]
  assign _T_62551 = _T_62550[10:0]; // @[Modules.scala 68:83:@11335.4]
  assign buffer_4_613 = $signed(_T_62551); // @[Modules.scala 68:83:@11336.4]
  assign _T_62559 = $signed(buffer_1_448) + $signed(buffer_4_449); // @[Modules.scala 68:83:@11346.4]
  assign _T_62560 = _T_62559[10:0]; // @[Modules.scala 68:83:@11347.4]
  assign buffer_4_616 = $signed(_T_62560); // @[Modules.scala 68:83:@11348.4]
  assign _T_62562 = $signed(buffer_4_450) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11350.4]
  assign _T_62563 = _T_62562[10:0]; // @[Modules.scala 68:83:@11351.4]
  assign buffer_4_617 = $signed(_T_62563); // @[Modules.scala 68:83:@11352.4]
  assign _T_62565 = $signed(buffer_4_452) + $signed(buffer_4_453); // @[Modules.scala 68:83:@11354.4]
  assign _T_62566 = _T_62565[10:0]; // @[Modules.scala 68:83:@11355.4]
  assign buffer_4_618 = $signed(_T_62566); // @[Modules.scala 68:83:@11356.4]
  assign _T_62571 = $signed(buffer_4_456) + $signed(buffer_4_457); // @[Modules.scala 68:83:@11362.4]
  assign _T_62572 = _T_62571[10:0]; // @[Modules.scala 68:83:@11363.4]
  assign buffer_4_620 = $signed(_T_62572); // @[Modules.scala 68:83:@11364.4]
  assign _T_62580 = $signed(buffer_4_462) + $signed(buffer_4_463); // @[Modules.scala 68:83:@11374.4]
  assign _T_62581 = _T_62580[10:0]; // @[Modules.scala 68:83:@11375.4]
  assign buffer_4_623 = $signed(_T_62581); // @[Modules.scala 68:83:@11376.4]
  assign _T_62586 = $signed(buffer_4_466) + $signed(buffer_4_467); // @[Modules.scala 68:83:@11382.4]
  assign _T_62587 = _T_62586[10:0]; // @[Modules.scala 68:83:@11383.4]
  assign buffer_4_625 = $signed(_T_62587); // @[Modules.scala 68:83:@11384.4]
  assign _T_62589 = $signed(buffer_1_468) + $signed(buffer_4_469); // @[Modules.scala 68:83:@11386.4]
  assign _T_62590 = _T_62589[10:0]; // @[Modules.scala 68:83:@11387.4]
  assign buffer_4_626 = $signed(_T_62590); // @[Modules.scala 68:83:@11388.4]
  assign _T_62592 = $signed(buffer_0_395) + $signed(buffer_1_471); // @[Modules.scala 68:83:@11390.4]
  assign _T_62593 = _T_62592[10:0]; // @[Modules.scala 68:83:@11391.4]
  assign buffer_4_627 = $signed(_T_62593); // @[Modules.scala 68:83:@11392.4]
  assign _T_62595 = $signed(buffer_4_472) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11394.4]
  assign _T_62596 = _T_62595[10:0]; // @[Modules.scala 68:83:@11395.4]
  assign buffer_4_628 = $signed(_T_62596); // @[Modules.scala 68:83:@11396.4]
  assign _T_62598 = $signed(buffer_1_474) + $signed(buffer_4_475); // @[Modules.scala 68:83:@11398.4]
  assign _T_62599 = _T_62598[10:0]; // @[Modules.scala 68:83:@11399.4]
  assign buffer_4_629 = $signed(_T_62599); // @[Modules.scala 68:83:@11400.4]
  assign _T_62601 = $signed(buffer_0_476) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11402.4]
  assign _T_62602 = _T_62601[10:0]; // @[Modules.scala 68:83:@11403.4]
  assign buffer_4_630 = $signed(_T_62602); // @[Modules.scala 68:83:@11404.4]
  assign _T_62604 = $signed(buffer_4_478) + $signed(buffer_1_479); // @[Modules.scala 68:83:@11406.4]
  assign _T_62605 = _T_62604[10:0]; // @[Modules.scala 68:83:@11407.4]
  assign buffer_4_631 = $signed(_T_62605); // @[Modules.scala 68:83:@11408.4]
  assign _T_62607 = $signed(buffer_4_480) + $signed(buffer_1_481); // @[Modules.scala 68:83:@11410.4]
  assign _T_62608 = _T_62607[10:0]; // @[Modules.scala 68:83:@11411.4]
  assign buffer_4_632 = $signed(_T_62608); // @[Modules.scala 68:83:@11412.4]
  assign _T_62610 = $signed(buffer_4_482) + $signed(buffer_4_483); // @[Modules.scala 68:83:@11414.4]
  assign _T_62611 = _T_62610[10:0]; // @[Modules.scala 68:83:@11415.4]
  assign buffer_4_633 = $signed(_T_62611); // @[Modules.scala 68:83:@11416.4]
  assign _T_62613 = $signed(buffer_4_484) + $signed(buffer_0_485); // @[Modules.scala 68:83:@11418.4]
  assign _T_62614 = _T_62613[10:0]; // @[Modules.scala 68:83:@11419.4]
  assign buffer_4_634 = $signed(_T_62614); // @[Modules.scala 68:83:@11420.4]
  assign _T_62616 = $signed(buffer_1_486) + $signed(buffer_4_487); // @[Modules.scala 68:83:@11422.4]
  assign _T_62617 = _T_62616[10:0]; // @[Modules.scala 68:83:@11423.4]
  assign buffer_4_635 = $signed(_T_62617); // @[Modules.scala 68:83:@11424.4]
  assign _T_62619 = $signed(buffer_4_488) + $signed(buffer_4_489); // @[Modules.scala 68:83:@11426.4]
  assign _T_62620 = _T_62619[10:0]; // @[Modules.scala 68:83:@11427.4]
  assign buffer_4_636 = $signed(_T_62620); // @[Modules.scala 68:83:@11428.4]
  assign _T_62622 = $signed(buffer_4_490) + $signed(buffer_4_491); // @[Modules.scala 68:83:@11430.4]
  assign _T_62623 = _T_62622[10:0]; // @[Modules.scala 68:83:@11431.4]
  assign buffer_4_637 = $signed(_T_62623); // @[Modules.scala 68:83:@11432.4]
  assign _T_62625 = $signed(buffer_4_492) + $signed(buffer_4_493); // @[Modules.scala 68:83:@11434.4]
  assign _T_62626 = _T_62625[10:0]; // @[Modules.scala 68:83:@11435.4]
  assign buffer_4_638 = $signed(_T_62626); // @[Modules.scala 68:83:@11436.4]
  assign _T_62628 = $signed(buffer_4_494) + $signed(buffer_4_495); // @[Modules.scala 68:83:@11438.4]
  assign _T_62629 = _T_62628[10:0]; // @[Modules.scala 68:83:@11439.4]
  assign buffer_4_639 = $signed(_T_62629); // @[Modules.scala 68:83:@11440.4]
  assign _T_62631 = $signed(buffer_4_496) + $signed(buffer_4_497); // @[Modules.scala 68:83:@11442.4]
  assign _T_62632 = _T_62631[10:0]; // @[Modules.scala 68:83:@11443.4]
  assign buffer_4_640 = $signed(_T_62632); // @[Modules.scala 68:83:@11444.4]
  assign _T_62634 = $signed(buffer_3_498) + $signed(buffer_0_499); // @[Modules.scala 68:83:@11446.4]
  assign _T_62635 = _T_62634[10:0]; // @[Modules.scala 68:83:@11447.4]
  assign buffer_4_641 = $signed(_T_62635); // @[Modules.scala 68:83:@11448.4]
  assign _T_62637 = $signed(buffer_4_500) + $signed(buffer_4_501); // @[Modules.scala 68:83:@11450.4]
  assign _T_62638 = _T_62637[10:0]; // @[Modules.scala 68:83:@11451.4]
  assign buffer_4_642 = $signed(_T_62638); // @[Modules.scala 68:83:@11452.4]
  assign _T_62640 = $signed(buffer_4_502) + $signed(buffer_3_503); // @[Modules.scala 68:83:@11454.4]
  assign _T_62641 = _T_62640[10:0]; // @[Modules.scala 68:83:@11455.4]
  assign buffer_4_643 = $signed(_T_62641); // @[Modules.scala 68:83:@11456.4]
  assign _T_62643 = $signed(buffer_1_504) + $signed(buffer_4_505); // @[Modules.scala 68:83:@11458.4]
  assign _T_62644 = _T_62643[10:0]; // @[Modules.scala 68:83:@11459.4]
  assign buffer_4_644 = $signed(_T_62644); // @[Modules.scala 68:83:@11460.4]
  assign _T_62646 = $signed(buffer_1_506) + $signed(buffer_4_507); // @[Modules.scala 68:83:@11462.4]
  assign _T_62647 = _T_62646[10:0]; // @[Modules.scala 68:83:@11463.4]
  assign buffer_4_645 = $signed(_T_62647); // @[Modules.scala 68:83:@11464.4]
  assign _T_62649 = $signed(buffer_4_508) + $signed(buffer_1_509); // @[Modules.scala 68:83:@11466.4]
  assign _T_62650 = _T_62649[10:0]; // @[Modules.scala 68:83:@11467.4]
  assign buffer_4_646 = $signed(_T_62650); // @[Modules.scala 68:83:@11468.4]
  assign _T_62652 = $signed(buffer_3_510) + $signed(buffer_4_511); // @[Modules.scala 68:83:@11470.4]
  assign _T_62653 = _T_62652[10:0]; // @[Modules.scala 68:83:@11471.4]
  assign buffer_4_647 = $signed(_T_62653); // @[Modules.scala 68:83:@11472.4]
  assign _T_62655 = $signed(buffer_4_512) + $signed(buffer_4_513); // @[Modules.scala 68:83:@11474.4]
  assign _T_62656 = _T_62655[10:0]; // @[Modules.scala 68:83:@11475.4]
  assign buffer_4_648 = $signed(_T_62656); // @[Modules.scala 68:83:@11476.4]
  assign _T_62658 = $signed(buffer_0_395) + $signed(buffer_4_515); // @[Modules.scala 68:83:@11478.4]
  assign _T_62659 = _T_62658[10:0]; // @[Modules.scala 68:83:@11479.4]
  assign buffer_4_649 = $signed(_T_62659); // @[Modules.scala 68:83:@11480.4]
  assign _T_62664 = $signed(buffer_4_518) + $signed(buffer_3_519); // @[Modules.scala 68:83:@11486.4]
  assign _T_62665 = _T_62664[10:0]; // @[Modules.scala 68:83:@11487.4]
  assign buffer_4_651 = $signed(_T_62665); // @[Modules.scala 68:83:@11488.4]
  assign _T_62667 = $signed(buffer_4_520) + $signed(buffer_4_521); // @[Modules.scala 68:83:@11490.4]
  assign _T_62668 = _T_62667[10:0]; // @[Modules.scala 68:83:@11491.4]
  assign buffer_4_652 = $signed(_T_62668); // @[Modules.scala 68:83:@11492.4]
  assign _T_62670 = $signed(buffer_4_522) + $signed(buffer_4_523); // @[Modules.scala 68:83:@11494.4]
  assign _T_62671 = _T_62670[10:0]; // @[Modules.scala 68:83:@11495.4]
  assign buffer_4_653 = $signed(_T_62671); // @[Modules.scala 68:83:@11496.4]
  assign _T_62673 = $signed(buffer_0_524) + $signed(buffer_4_525); // @[Modules.scala 68:83:@11498.4]
  assign _T_62674 = _T_62673[10:0]; // @[Modules.scala 68:83:@11499.4]
  assign buffer_4_654 = $signed(_T_62674); // @[Modules.scala 68:83:@11500.4]
  assign _T_62679 = $signed(buffer_4_528) + $signed(buffer_1_529); // @[Modules.scala 68:83:@11506.4]
  assign _T_62680 = _T_62679[10:0]; // @[Modules.scala 68:83:@11507.4]
  assign buffer_4_656 = $signed(_T_62680); // @[Modules.scala 68:83:@11508.4]
  assign _T_62682 = $signed(buffer_3_530) + $signed(buffer_4_531); // @[Modules.scala 68:83:@11510.4]
  assign _T_62683 = _T_62682[10:0]; // @[Modules.scala 68:83:@11511.4]
  assign buffer_4_657 = $signed(_T_62683); // @[Modules.scala 68:83:@11512.4]
  assign _T_62685 = $signed(buffer_1_532) + $signed(buffer_3_533); // @[Modules.scala 68:83:@11514.4]
  assign _T_62686 = _T_62685[10:0]; // @[Modules.scala 68:83:@11515.4]
  assign buffer_4_658 = $signed(_T_62686); // @[Modules.scala 68:83:@11516.4]
  assign _T_62688 = $signed(buffer_1_534) + $signed(buffer_4_535); // @[Modules.scala 68:83:@11518.4]
  assign _T_62689 = _T_62688[10:0]; // @[Modules.scala 68:83:@11519.4]
  assign buffer_4_659 = $signed(_T_62689); // @[Modules.scala 68:83:@11520.4]
  assign _T_62691 = $signed(buffer_2_536) + $signed(buffer_4_537); // @[Modules.scala 68:83:@11522.4]
  assign _T_62692 = _T_62691[10:0]; // @[Modules.scala 68:83:@11523.4]
  assign buffer_4_660 = $signed(_T_62692); // @[Modules.scala 68:83:@11524.4]
  assign _T_62694 = $signed(buffer_4_538) + $signed(buffer_4_539); // @[Modules.scala 68:83:@11526.4]
  assign _T_62695 = _T_62694[10:0]; // @[Modules.scala 68:83:@11527.4]
  assign buffer_4_661 = $signed(_T_62695); // @[Modules.scala 68:83:@11528.4]
  assign _T_62697 = $signed(buffer_3_540) + $signed(buffer_4_541); // @[Modules.scala 68:83:@11530.4]
  assign _T_62698 = _T_62697[10:0]; // @[Modules.scala 68:83:@11531.4]
  assign buffer_4_662 = $signed(_T_62698); // @[Modules.scala 68:83:@11532.4]
  assign _T_62703 = $signed(buffer_4_544) + $signed(buffer_4_545); // @[Modules.scala 68:83:@11538.4]
  assign _T_62704 = _T_62703[10:0]; // @[Modules.scala 68:83:@11539.4]
  assign buffer_4_664 = $signed(_T_62704); // @[Modules.scala 68:83:@11540.4]
  assign _T_62706 = $signed(buffer_0_546) + $signed(buffer_4_547); // @[Modules.scala 68:83:@11542.4]
  assign _T_62707 = _T_62706[10:0]; // @[Modules.scala 68:83:@11543.4]
  assign buffer_4_665 = $signed(_T_62707); // @[Modules.scala 68:83:@11544.4]
  assign _T_62709 = $signed(buffer_4_548) + $signed(buffer_1_549); // @[Modules.scala 68:83:@11546.4]
  assign _T_62710 = _T_62709[10:0]; // @[Modules.scala 68:83:@11547.4]
  assign buffer_4_666 = $signed(_T_62710); // @[Modules.scala 68:83:@11548.4]
  assign _T_62712 = $signed(buffer_4_550) + $signed(buffer_3_551); // @[Modules.scala 68:83:@11550.4]
  assign _T_62713 = _T_62712[10:0]; // @[Modules.scala 68:83:@11551.4]
  assign buffer_4_667 = $signed(_T_62713); // @[Modules.scala 68:83:@11552.4]
  assign _T_62715 = $signed(buffer_4_552) + $signed(buffer_0_553); // @[Modules.scala 68:83:@11554.4]
  assign _T_62716 = _T_62715[10:0]; // @[Modules.scala 68:83:@11555.4]
  assign buffer_4_668 = $signed(_T_62716); // @[Modules.scala 68:83:@11556.4]
  assign _T_62718 = $signed(buffer_4_554) + $signed(buffer_1_555); // @[Modules.scala 68:83:@11558.4]
  assign _T_62719 = _T_62718[10:0]; // @[Modules.scala 68:83:@11559.4]
  assign buffer_4_669 = $signed(_T_62719); // @[Modules.scala 68:83:@11560.4]
  assign _T_62721 = $signed(buffer_1_556) + $signed(buffer_4_557); // @[Modules.scala 68:83:@11562.4]
  assign _T_62722 = _T_62721[10:0]; // @[Modules.scala 68:83:@11563.4]
  assign buffer_4_670 = $signed(_T_62722); // @[Modules.scala 68:83:@11564.4]
  assign _T_62724 = $signed(buffer_4_558) + $signed(buffer_4_559); // @[Modules.scala 68:83:@11566.4]
  assign _T_62725 = _T_62724[10:0]; // @[Modules.scala 68:83:@11567.4]
  assign buffer_4_671 = $signed(_T_62725); // @[Modules.scala 68:83:@11568.4]
  assign _T_62727 = $signed(buffer_4_560) + $signed(buffer_4_561); // @[Modules.scala 68:83:@11570.4]
  assign _T_62728 = _T_62727[10:0]; // @[Modules.scala 68:83:@11571.4]
  assign buffer_4_672 = $signed(_T_62728); // @[Modules.scala 68:83:@11572.4]
  assign _T_62730 = $signed(buffer_3_562) + $signed(buffer_4_563); // @[Modules.scala 68:83:@11574.4]
  assign _T_62731 = _T_62730[10:0]; // @[Modules.scala 68:83:@11575.4]
  assign buffer_4_673 = $signed(_T_62731); // @[Modules.scala 68:83:@11576.4]
  assign _T_62733 = $signed(buffer_4_564) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11578.4]
  assign _T_62734 = _T_62733[10:0]; // @[Modules.scala 68:83:@11579.4]
  assign buffer_4_674 = $signed(_T_62734); // @[Modules.scala 68:83:@11580.4]
  assign _T_62736 = $signed(buffer_4_566) + $signed(buffer_1_567); // @[Modules.scala 68:83:@11582.4]
  assign _T_62737 = _T_62736[10:0]; // @[Modules.scala 68:83:@11583.4]
  assign buffer_4_675 = $signed(_T_62737); // @[Modules.scala 68:83:@11584.4]
  assign _T_62739 = $signed(buffer_4_568) + $signed(buffer_0_395); // @[Modules.scala 68:83:@11586.4]
  assign _T_62740 = _T_62739[10:0]; // @[Modules.scala 68:83:@11587.4]
  assign buffer_4_676 = $signed(_T_62740); // @[Modules.scala 68:83:@11588.4]
  assign _T_62745 = $signed(buffer_0_395) + $signed(buffer_4_573); // @[Modules.scala 68:83:@11594.4]
  assign _T_62746 = _T_62745[10:0]; // @[Modules.scala 68:83:@11595.4]
  assign buffer_4_678 = $signed(_T_62746); // @[Modules.scala 68:83:@11596.4]
  assign _T_62748 = $signed(buffer_3_574) + $signed(buffer_2_575); // @[Modules.scala 68:83:@11598.4]
  assign _T_62749 = _T_62748[10:0]; // @[Modules.scala 68:83:@11599.4]
  assign buffer_4_679 = $signed(_T_62749); // @[Modules.scala 68:83:@11600.4]
  assign _T_62757 = $signed(buffer_4_580) + $signed(buffer_4_581); // @[Modules.scala 68:83:@11610.4]
  assign _T_62758 = _T_62757[10:0]; // @[Modules.scala 68:83:@11611.4]
  assign buffer_4_682 = $signed(_T_62758); // @[Modules.scala 68:83:@11612.4]
  assign _T_62760 = $signed(buffer_4_582) + $signed(buffer_4_583); // @[Modules.scala 68:83:@11614.4]
  assign _T_62761 = _T_62760[10:0]; // @[Modules.scala 68:83:@11615.4]
  assign buffer_4_683 = $signed(_T_62761); // @[Modules.scala 68:83:@11616.4]
  assign _T_62763 = $signed(buffer_4_584) + $signed(buffer_4_585); // @[Modules.scala 68:83:@11618.4]
  assign _T_62764 = _T_62763[10:0]; // @[Modules.scala 68:83:@11619.4]
  assign buffer_4_684 = $signed(_T_62764); // @[Modules.scala 68:83:@11620.4]
  assign _T_62766 = $signed(buffer_0_395) + $signed(buffer_4_587); // @[Modules.scala 68:83:@11622.4]
  assign _T_62767 = _T_62766[10:0]; // @[Modules.scala 68:83:@11623.4]
  assign buffer_4_685 = $signed(_T_62767); // @[Modules.scala 68:83:@11624.4]
  assign _T_62769 = $signed(buffer_4_588) + $signed(buffer_4_589); // @[Modules.scala 71:109:@11626.4]
  assign _T_62770 = _T_62769[10:0]; // @[Modules.scala 71:109:@11627.4]
  assign buffer_4_686 = $signed(_T_62770); // @[Modules.scala 71:109:@11628.4]
  assign _T_62772 = $signed(buffer_4_590) + $signed(buffer_4_591); // @[Modules.scala 71:109:@11630.4]
  assign _T_62773 = _T_62772[10:0]; // @[Modules.scala 71:109:@11631.4]
  assign buffer_4_687 = $signed(_T_62773); // @[Modules.scala 71:109:@11632.4]
  assign _T_62775 = $signed(buffer_4_592) + $signed(buffer_4_593); // @[Modules.scala 71:109:@11634.4]
  assign _T_62776 = _T_62775[10:0]; // @[Modules.scala 71:109:@11635.4]
  assign buffer_4_688 = $signed(_T_62776); // @[Modules.scala 71:109:@11636.4]
  assign _T_62778 = $signed(buffer_4_594) + $signed(buffer_4_595); // @[Modules.scala 71:109:@11638.4]
  assign _T_62779 = _T_62778[10:0]; // @[Modules.scala 71:109:@11639.4]
  assign buffer_4_689 = $signed(_T_62779); // @[Modules.scala 71:109:@11640.4]
  assign _T_62784 = $signed(buffer_4_598) + $signed(buffer_4_599); // @[Modules.scala 71:109:@11646.4]
  assign _T_62785 = _T_62784[10:0]; // @[Modules.scala 71:109:@11647.4]
  assign buffer_4_691 = $signed(_T_62785); // @[Modules.scala 71:109:@11648.4]
  assign _T_62790 = $signed(buffer_4_602) + $signed(buffer_4_603); // @[Modules.scala 71:109:@11654.4]
  assign _T_62791 = _T_62790[10:0]; // @[Modules.scala 71:109:@11655.4]
  assign buffer_4_693 = $signed(_T_62791); // @[Modules.scala 71:109:@11656.4]
  assign _T_62793 = $signed(buffer_4_604) + $signed(buffer_4_605); // @[Modules.scala 71:109:@11658.4]
  assign _T_62794 = _T_62793[10:0]; // @[Modules.scala 71:109:@11659.4]
  assign buffer_4_694 = $signed(_T_62794); // @[Modules.scala 71:109:@11660.4]
  assign _T_62796 = $signed(buffer_4_606) + $signed(buffer_4_607); // @[Modules.scala 71:109:@11662.4]
  assign _T_62797 = _T_62796[10:0]; // @[Modules.scala 71:109:@11663.4]
  assign buffer_4_695 = $signed(_T_62797); // @[Modules.scala 71:109:@11664.4]
  assign _T_62799 = $signed(buffer_4_608) + $signed(buffer_4_609); // @[Modules.scala 71:109:@11666.4]
  assign _T_62800 = _T_62799[10:0]; // @[Modules.scala 71:109:@11667.4]
  assign buffer_4_696 = $signed(_T_62800); // @[Modules.scala 71:109:@11668.4]
  assign _T_62802 = $signed(buffer_4_610) + $signed(buffer_4_611); // @[Modules.scala 71:109:@11670.4]
  assign _T_62803 = _T_62802[10:0]; // @[Modules.scala 71:109:@11671.4]
  assign buffer_4_697 = $signed(_T_62803); // @[Modules.scala 71:109:@11672.4]
  assign _T_62805 = $signed(buffer_4_612) + $signed(buffer_4_613); // @[Modules.scala 71:109:@11674.4]
  assign _T_62806 = _T_62805[10:0]; // @[Modules.scala 71:109:@11675.4]
  assign buffer_4_698 = $signed(_T_62806); // @[Modules.scala 71:109:@11676.4]
  assign _T_62808 = $signed(buffer_0_593) + $signed(buffer_2_615); // @[Modules.scala 71:109:@11678.4]
  assign _T_62809 = _T_62808[10:0]; // @[Modules.scala 71:109:@11679.4]
  assign buffer_4_699 = $signed(_T_62809); // @[Modules.scala 71:109:@11680.4]
  assign _T_62811 = $signed(buffer_4_616) + $signed(buffer_4_617); // @[Modules.scala 71:109:@11682.4]
  assign _T_62812 = _T_62811[10:0]; // @[Modules.scala 71:109:@11683.4]
  assign buffer_4_700 = $signed(_T_62812); // @[Modules.scala 71:109:@11684.4]
  assign _T_62814 = $signed(buffer_4_618) + $signed(buffer_2_619); // @[Modules.scala 71:109:@11686.4]
  assign _T_62815 = _T_62814[10:0]; // @[Modules.scala 71:109:@11687.4]
  assign buffer_4_701 = $signed(_T_62815); // @[Modules.scala 71:109:@11688.4]
  assign _T_62817 = $signed(buffer_4_620) + $signed(buffer_0_593); // @[Modules.scala 71:109:@11690.4]
  assign _T_62818 = _T_62817[10:0]; // @[Modules.scala 71:109:@11691.4]
  assign buffer_4_702 = $signed(_T_62818); // @[Modules.scala 71:109:@11692.4]
  assign _T_62820 = $signed(buffer_3_622) + $signed(buffer_4_623); // @[Modules.scala 71:109:@11694.4]
  assign _T_62821 = _T_62820[10:0]; // @[Modules.scala 71:109:@11695.4]
  assign buffer_4_703 = $signed(_T_62821); // @[Modules.scala 71:109:@11696.4]
  assign _T_62823 = $signed(buffer_0_624) + $signed(buffer_4_625); // @[Modules.scala 71:109:@11698.4]
  assign _T_62824 = _T_62823[10:0]; // @[Modules.scala 71:109:@11699.4]
  assign buffer_4_704 = $signed(_T_62824); // @[Modules.scala 71:109:@11700.4]
  assign _T_62826 = $signed(buffer_4_626) + $signed(buffer_4_627); // @[Modules.scala 71:109:@11702.4]
  assign _T_62827 = _T_62826[10:0]; // @[Modules.scala 71:109:@11703.4]
  assign buffer_4_705 = $signed(_T_62827); // @[Modules.scala 71:109:@11704.4]
  assign _T_62829 = $signed(buffer_4_628) + $signed(buffer_4_629); // @[Modules.scala 71:109:@11706.4]
  assign _T_62830 = _T_62829[10:0]; // @[Modules.scala 71:109:@11707.4]
  assign buffer_4_706 = $signed(_T_62830); // @[Modules.scala 71:109:@11708.4]
  assign _T_62832 = $signed(buffer_4_630) + $signed(buffer_4_631); // @[Modules.scala 71:109:@11710.4]
  assign _T_62833 = _T_62832[10:0]; // @[Modules.scala 71:109:@11711.4]
  assign buffer_4_707 = $signed(_T_62833); // @[Modules.scala 71:109:@11712.4]
  assign _T_62835 = $signed(buffer_4_632) + $signed(buffer_4_633); // @[Modules.scala 71:109:@11714.4]
  assign _T_62836 = _T_62835[10:0]; // @[Modules.scala 71:109:@11715.4]
  assign buffer_4_708 = $signed(_T_62836); // @[Modules.scala 71:109:@11716.4]
  assign _T_62838 = $signed(buffer_4_634) + $signed(buffer_4_635); // @[Modules.scala 71:109:@11718.4]
  assign _T_62839 = _T_62838[10:0]; // @[Modules.scala 71:109:@11719.4]
  assign buffer_4_709 = $signed(_T_62839); // @[Modules.scala 71:109:@11720.4]
  assign _T_62841 = $signed(buffer_4_636) + $signed(buffer_4_637); // @[Modules.scala 71:109:@11722.4]
  assign _T_62842 = _T_62841[10:0]; // @[Modules.scala 71:109:@11723.4]
  assign buffer_4_710 = $signed(_T_62842); // @[Modules.scala 71:109:@11724.4]
  assign _T_62844 = $signed(buffer_4_638) + $signed(buffer_4_639); // @[Modules.scala 71:109:@11726.4]
  assign _T_62845 = _T_62844[10:0]; // @[Modules.scala 71:109:@11727.4]
  assign buffer_4_711 = $signed(_T_62845); // @[Modules.scala 71:109:@11728.4]
  assign _T_62847 = $signed(buffer_4_640) + $signed(buffer_4_641); // @[Modules.scala 71:109:@11730.4]
  assign _T_62848 = _T_62847[10:0]; // @[Modules.scala 71:109:@11731.4]
  assign buffer_4_712 = $signed(_T_62848); // @[Modules.scala 71:109:@11732.4]
  assign _T_62850 = $signed(buffer_4_642) + $signed(buffer_4_643); // @[Modules.scala 71:109:@11734.4]
  assign _T_62851 = _T_62850[10:0]; // @[Modules.scala 71:109:@11735.4]
  assign buffer_4_713 = $signed(_T_62851); // @[Modules.scala 71:109:@11736.4]
  assign _T_62853 = $signed(buffer_4_644) + $signed(buffer_4_645); // @[Modules.scala 71:109:@11738.4]
  assign _T_62854 = _T_62853[10:0]; // @[Modules.scala 71:109:@11739.4]
  assign buffer_4_714 = $signed(_T_62854); // @[Modules.scala 71:109:@11740.4]
  assign _T_62856 = $signed(buffer_4_646) + $signed(buffer_4_647); // @[Modules.scala 71:109:@11742.4]
  assign _T_62857 = _T_62856[10:0]; // @[Modules.scala 71:109:@11743.4]
  assign buffer_4_715 = $signed(_T_62857); // @[Modules.scala 71:109:@11744.4]
  assign _T_62859 = $signed(buffer_4_648) + $signed(buffer_4_649); // @[Modules.scala 71:109:@11746.4]
  assign _T_62860 = _T_62859[10:0]; // @[Modules.scala 71:109:@11747.4]
  assign buffer_4_716 = $signed(_T_62860); // @[Modules.scala 71:109:@11748.4]
  assign _T_62862 = $signed(buffer_3_650) + $signed(buffer_4_651); // @[Modules.scala 71:109:@11750.4]
  assign _T_62863 = _T_62862[10:0]; // @[Modules.scala 71:109:@11751.4]
  assign buffer_4_717 = $signed(_T_62863); // @[Modules.scala 71:109:@11752.4]
  assign _T_62865 = $signed(buffer_4_652) + $signed(buffer_4_653); // @[Modules.scala 71:109:@11754.4]
  assign _T_62866 = _T_62865[10:0]; // @[Modules.scala 71:109:@11755.4]
  assign buffer_4_718 = $signed(_T_62866); // @[Modules.scala 71:109:@11756.4]
  assign _T_62868 = $signed(buffer_4_654) + $signed(buffer_1_655); // @[Modules.scala 71:109:@11758.4]
  assign _T_62869 = _T_62868[10:0]; // @[Modules.scala 71:109:@11759.4]
  assign buffer_4_719 = $signed(_T_62869); // @[Modules.scala 71:109:@11760.4]
  assign _T_62871 = $signed(buffer_4_656) + $signed(buffer_4_657); // @[Modules.scala 71:109:@11762.4]
  assign _T_62872 = _T_62871[10:0]; // @[Modules.scala 71:109:@11763.4]
  assign buffer_4_720 = $signed(_T_62872); // @[Modules.scala 71:109:@11764.4]
  assign _T_62874 = $signed(buffer_4_658) + $signed(buffer_4_659); // @[Modules.scala 71:109:@11766.4]
  assign _T_62875 = _T_62874[10:0]; // @[Modules.scala 71:109:@11767.4]
  assign buffer_4_721 = $signed(_T_62875); // @[Modules.scala 71:109:@11768.4]
  assign _T_62877 = $signed(buffer_4_660) + $signed(buffer_4_661); // @[Modules.scala 71:109:@11770.4]
  assign _T_62878 = _T_62877[10:0]; // @[Modules.scala 71:109:@11771.4]
  assign buffer_4_722 = $signed(_T_62878); // @[Modules.scala 71:109:@11772.4]
  assign _T_62880 = $signed(buffer_4_662) + $signed(buffer_0_663); // @[Modules.scala 71:109:@11774.4]
  assign _T_62881 = _T_62880[10:0]; // @[Modules.scala 71:109:@11775.4]
  assign buffer_4_723 = $signed(_T_62881); // @[Modules.scala 71:109:@11776.4]
  assign _T_62883 = $signed(buffer_4_664) + $signed(buffer_4_665); // @[Modules.scala 71:109:@11778.4]
  assign _T_62884 = _T_62883[10:0]; // @[Modules.scala 71:109:@11779.4]
  assign buffer_4_724 = $signed(_T_62884); // @[Modules.scala 71:109:@11780.4]
  assign _T_62886 = $signed(buffer_4_666) + $signed(buffer_4_667); // @[Modules.scala 71:109:@11782.4]
  assign _T_62887 = _T_62886[10:0]; // @[Modules.scala 71:109:@11783.4]
  assign buffer_4_725 = $signed(_T_62887); // @[Modules.scala 71:109:@11784.4]
  assign _T_62889 = $signed(buffer_4_668) + $signed(buffer_4_669); // @[Modules.scala 71:109:@11786.4]
  assign _T_62890 = _T_62889[10:0]; // @[Modules.scala 71:109:@11787.4]
  assign buffer_4_726 = $signed(_T_62890); // @[Modules.scala 71:109:@11788.4]
  assign _T_62892 = $signed(buffer_4_670) + $signed(buffer_4_671); // @[Modules.scala 71:109:@11790.4]
  assign _T_62893 = _T_62892[10:0]; // @[Modules.scala 71:109:@11791.4]
  assign buffer_4_727 = $signed(_T_62893); // @[Modules.scala 71:109:@11792.4]
  assign _T_62895 = $signed(buffer_4_672) + $signed(buffer_4_673); // @[Modules.scala 71:109:@11794.4]
  assign _T_62896 = _T_62895[10:0]; // @[Modules.scala 71:109:@11795.4]
  assign buffer_4_728 = $signed(_T_62896); // @[Modules.scala 71:109:@11796.4]
  assign _T_62898 = $signed(buffer_4_674) + $signed(buffer_4_675); // @[Modules.scala 71:109:@11798.4]
  assign _T_62899 = _T_62898[10:0]; // @[Modules.scala 71:109:@11799.4]
  assign buffer_4_729 = $signed(_T_62899); // @[Modules.scala 71:109:@11800.4]
  assign _T_62901 = $signed(buffer_4_676) + $signed(buffer_0_593); // @[Modules.scala 71:109:@11802.4]
  assign _T_62902 = _T_62901[10:0]; // @[Modules.scala 71:109:@11803.4]
  assign buffer_4_730 = $signed(_T_62902); // @[Modules.scala 71:109:@11804.4]
  assign _T_62904 = $signed(buffer_4_678) + $signed(buffer_4_679); // @[Modules.scala 71:109:@11806.4]
  assign _T_62905 = _T_62904[10:0]; // @[Modules.scala 71:109:@11807.4]
  assign buffer_4_731 = $signed(_T_62905); // @[Modules.scala 71:109:@11808.4]
  assign _T_62910 = $signed(buffer_4_682) + $signed(buffer_4_683); // @[Modules.scala 71:109:@11814.4]
  assign _T_62911 = _T_62910[10:0]; // @[Modules.scala 71:109:@11815.4]
  assign buffer_4_733 = $signed(_T_62911); // @[Modules.scala 71:109:@11816.4]
  assign _T_62913 = $signed(buffer_4_684) + $signed(buffer_4_685); // @[Modules.scala 71:109:@11818.4]
  assign _T_62914 = _T_62913[10:0]; // @[Modules.scala 71:109:@11819.4]
  assign buffer_4_734 = $signed(_T_62914); // @[Modules.scala 71:109:@11820.4]
  assign _T_62916 = $signed(buffer_4_686) + $signed(buffer_4_687); // @[Modules.scala 78:156:@11823.4]
  assign _T_62917 = _T_62916[10:0]; // @[Modules.scala 78:156:@11824.4]
  assign buffer_4_736 = $signed(_T_62917); // @[Modules.scala 78:156:@11825.4]
  assign _T_62919 = $signed(buffer_4_736) + $signed(buffer_4_688); // @[Modules.scala 78:156:@11827.4]
  assign _T_62920 = _T_62919[10:0]; // @[Modules.scala 78:156:@11828.4]
  assign buffer_4_737 = $signed(_T_62920); // @[Modules.scala 78:156:@11829.4]
  assign _T_62922 = $signed(buffer_4_737) + $signed(buffer_4_689); // @[Modules.scala 78:156:@11831.4]
  assign _T_62923 = _T_62922[10:0]; // @[Modules.scala 78:156:@11832.4]
  assign buffer_4_738 = $signed(_T_62923); // @[Modules.scala 78:156:@11833.4]
  assign _T_62925 = $signed(buffer_4_738) + $signed(buffer_1_690); // @[Modules.scala 78:156:@11835.4]
  assign _T_62926 = _T_62925[10:0]; // @[Modules.scala 78:156:@11836.4]
  assign buffer_4_739 = $signed(_T_62926); // @[Modules.scala 78:156:@11837.4]
  assign _T_62928 = $signed(buffer_4_739) + $signed(buffer_4_691); // @[Modules.scala 78:156:@11839.4]
  assign _T_62929 = _T_62928[10:0]; // @[Modules.scala 78:156:@11840.4]
  assign buffer_4_740 = $signed(_T_62929); // @[Modules.scala 78:156:@11841.4]
  assign _T_62931 = $signed(buffer_4_740) + $signed(buffer_1_692); // @[Modules.scala 78:156:@11843.4]
  assign _T_62932 = _T_62931[10:0]; // @[Modules.scala 78:156:@11844.4]
  assign buffer_4_741 = $signed(_T_62932); // @[Modules.scala 78:156:@11845.4]
  assign _T_62934 = $signed(buffer_4_741) + $signed(buffer_4_693); // @[Modules.scala 78:156:@11847.4]
  assign _T_62935 = _T_62934[10:0]; // @[Modules.scala 78:156:@11848.4]
  assign buffer_4_742 = $signed(_T_62935); // @[Modules.scala 78:156:@11849.4]
  assign _T_62937 = $signed(buffer_4_742) + $signed(buffer_4_694); // @[Modules.scala 78:156:@11851.4]
  assign _T_62938 = _T_62937[10:0]; // @[Modules.scala 78:156:@11852.4]
  assign buffer_4_743 = $signed(_T_62938); // @[Modules.scala 78:156:@11853.4]
  assign _T_62940 = $signed(buffer_4_743) + $signed(buffer_4_695); // @[Modules.scala 78:156:@11855.4]
  assign _T_62941 = _T_62940[10:0]; // @[Modules.scala 78:156:@11856.4]
  assign buffer_4_744 = $signed(_T_62941); // @[Modules.scala 78:156:@11857.4]
  assign _T_62943 = $signed(buffer_4_744) + $signed(buffer_4_696); // @[Modules.scala 78:156:@11859.4]
  assign _T_62944 = _T_62943[10:0]; // @[Modules.scala 78:156:@11860.4]
  assign buffer_4_745 = $signed(_T_62944); // @[Modules.scala 78:156:@11861.4]
  assign _T_62946 = $signed(buffer_4_745) + $signed(buffer_4_697); // @[Modules.scala 78:156:@11863.4]
  assign _T_62947 = _T_62946[10:0]; // @[Modules.scala 78:156:@11864.4]
  assign buffer_4_746 = $signed(_T_62947); // @[Modules.scala 78:156:@11865.4]
  assign _T_62949 = $signed(buffer_4_746) + $signed(buffer_4_698); // @[Modules.scala 78:156:@11867.4]
  assign _T_62950 = _T_62949[10:0]; // @[Modules.scala 78:156:@11868.4]
  assign buffer_4_747 = $signed(_T_62950); // @[Modules.scala 78:156:@11869.4]
  assign _T_62952 = $signed(buffer_4_747) + $signed(buffer_4_699); // @[Modules.scala 78:156:@11871.4]
  assign _T_62953 = _T_62952[10:0]; // @[Modules.scala 78:156:@11872.4]
  assign buffer_4_748 = $signed(_T_62953); // @[Modules.scala 78:156:@11873.4]
  assign _T_62955 = $signed(buffer_4_748) + $signed(buffer_4_700); // @[Modules.scala 78:156:@11875.4]
  assign _T_62956 = _T_62955[10:0]; // @[Modules.scala 78:156:@11876.4]
  assign buffer_4_749 = $signed(_T_62956); // @[Modules.scala 78:156:@11877.4]
  assign _T_62958 = $signed(buffer_4_749) + $signed(buffer_4_701); // @[Modules.scala 78:156:@11879.4]
  assign _T_62959 = _T_62958[10:0]; // @[Modules.scala 78:156:@11880.4]
  assign buffer_4_750 = $signed(_T_62959); // @[Modules.scala 78:156:@11881.4]
  assign _T_62961 = $signed(buffer_4_750) + $signed(buffer_4_702); // @[Modules.scala 78:156:@11883.4]
  assign _T_62962 = _T_62961[10:0]; // @[Modules.scala 78:156:@11884.4]
  assign buffer_4_751 = $signed(_T_62962); // @[Modules.scala 78:156:@11885.4]
  assign _T_62964 = $signed(buffer_4_751) + $signed(buffer_4_703); // @[Modules.scala 78:156:@11887.4]
  assign _T_62965 = _T_62964[10:0]; // @[Modules.scala 78:156:@11888.4]
  assign buffer_4_752 = $signed(_T_62965); // @[Modules.scala 78:156:@11889.4]
  assign _T_62967 = $signed(buffer_4_752) + $signed(buffer_4_704); // @[Modules.scala 78:156:@11891.4]
  assign _T_62968 = _T_62967[10:0]; // @[Modules.scala 78:156:@11892.4]
  assign buffer_4_753 = $signed(_T_62968); // @[Modules.scala 78:156:@11893.4]
  assign _T_62970 = $signed(buffer_4_753) + $signed(buffer_4_705); // @[Modules.scala 78:156:@11895.4]
  assign _T_62971 = _T_62970[10:0]; // @[Modules.scala 78:156:@11896.4]
  assign buffer_4_754 = $signed(_T_62971); // @[Modules.scala 78:156:@11897.4]
  assign _T_62973 = $signed(buffer_4_754) + $signed(buffer_4_706); // @[Modules.scala 78:156:@11899.4]
  assign _T_62974 = _T_62973[10:0]; // @[Modules.scala 78:156:@11900.4]
  assign buffer_4_755 = $signed(_T_62974); // @[Modules.scala 78:156:@11901.4]
  assign _T_62976 = $signed(buffer_4_755) + $signed(buffer_4_707); // @[Modules.scala 78:156:@11903.4]
  assign _T_62977 = _T_62976[10:0]; // @[Modules.scala 78:156:@11904.4]
  assign buffer_4_756 = $signed(_T_62977); // @[Modules.scala 78:156:@11905.4]
  assign _T_62979 = $signed(buffer_4_756) + $signed(buffer_4_708); // @[Modules.scala 78:156:@11907.4]
  assign _T_62980 = _T_62979[10:0]; // @[Modules.scala 78:156:@11908.4]
  assign buffer_4_757 = $signed(_T_62980); // @[Modules.scala 78:156:@11909.4]
  assign _T_62982 = $signed(buffer_4_757) + $signed(buffer_4_709); // @[Modules.scala 78:156:@11911.4]
  assign _T_62983 = _T_62982[10:0]; // @[Modules.scala 78:156:@11912.4]
  assign buffer_4_758 = $signed(_T_62983); // @[Modules.scala 78:156:@11913.4]
  assign _T_62985 = $signed(buffer_4_758) + $signed(buffer_4_710); // @[Modules.scala 78:156:@11915.4]
  assign _T_62986 = _T_62985[10:0]; // @[Modules.scala 78:156:@11916.4]
  assign buffer_4_759 = $signed(_T_62986); // @[Modules.scala 78:156:@11917.4]
  assign _T_62988 = $signed(buffer_4_759) + $signed(buffer_4_711); // @[Modules.scala 78:156:@11919.4]
  assign _T_62989 = _T_62988[10:0]; // @[Modules.scala 78:156:@11920.4]
  assign buffer_4_760 = $signed(_T_62989); // @[Modules.scala 78:156:@11921.4]
  assign _T_62991 = $signed(buffer_4_760) + $signed(buffer_4_712); // @[Modules.scala 78:156:@11923.4]
  assign _T_62992 = _T_62991[10:0]; // @[Modules.scala 78:156:@11924.4]
  assign buffer_4_761 = $signed(_T_62992); // @[Modules.scala 78:156:@11925.4]
  assign _T_62994 = $signed(buffer_4_761) + $signed(buffer_4_713); // @[Modules.scala 78:156:@11927.4]
  assign _T_62995 = _T_62994[10:0]; // @[Modules.scala 78:156:@11928.4]
  assign buffer_4_762 = $signed(_T_62995); // @[Modules.scala 78:156:@11929.4]
  assign _T_62997 = $signed(buffer_4_762) + $signed(buffer_4_714); // @[Modules.scala 78:156:@11931.4]
  assign _T_62998 = _T_62997[10:0]; // @[Modules.scala 78:156:@11932.4]
  assign buffer_4_763 = $signed(_T_62998); // @[Modules.scala 78:156:@11933.4]
  assign _T_63000 = $signed(buffer_4_763) + $signed(buffer_4_715); // @[Modules.scala 78:156:@11935.4]
  assign _T_63001 = _T_63000[10:0]; // @[Modules.scala 78:156:@11936.4]
  assign buffer_4_764 = $signed(_T_63001); // @[Modules.scala 78:156:@11937.4]
  assign _T_63003 = $signed(buffer_4_764) + $signed(buffer_4_716); // @[Modules.scala 78:156:@11939.4]
  assign _T_63004 = _T_63003[10:0]; // @[Modules.scala 78:156:@11940.4]
  assign buffer_4_765 = $signed(_T_63004); // @[Modules.scala 78:156:@11941.4]
  assign _T_63006 = $signed(buffer_4_765) + $signed(buffer_4_717); // @[Modules.scala 78:156:@11943.4]
  assign _T_63007 = _T_63006[10:0]; // @[Modules.scala 78:156:@11944.4]
  assign buffer_4_766 = $signed(_T_63007); // @[Modules.scala 78:156:@11945.4]
  assign _T_63009 = $signed(buffer_4_766) + $signed(buffer_4_718); // @[Modules.scala 78:156:@11947.4]
  assign _T_63010 = _T_63009[10:0]; // @[Modules.scala 78:156:@11948.4]
  assign buffer_4_767 = $signed(_T_63010); // @[Modules.scala 78:156:@11949.4]
  assign _T_63012 = $signed(buffer_4_767) + $signed(buffer_4_719); // @[Modules.scala 78:156:@11951.4]
  assign _T_63013 = _T_63012[10:0]; // @[Modules.scala 78:156:@11952.4]
  assign buffer_4_768 = $signed(_T_63013); // @[Modules.scala 78:156:@11953.4]
  assign _T_63015 = $signed(buffer_4_768) + $signed(buffer_4_720); // @[Modules.scala 78:156:@11955.4]
  assign _T_63016 = _T_63015[10:0]; // @[Modules.scala 78:156:@11956.4]
  assign buffer_4_769 = $signed(_T_63016); // @[Modules.scala 78:156:@11957.4]
  assign _T_63018 = $signed(buffer_4_769) + $signed(buffer_4_721); // @[Modules.scala 78:156:@11959.4]
  assign _T_63019 = _T_63018[10:0]; // @[Modules.scala 78:156:@11960.4]
  assign buffer_4_770 = $signed(_T_63019); // @[Modules.scala 78:156:@11961.4]
  assign _T_63021 = $signed(buffer_4_770) + $signed(buffer_4_722); // @[Modules.scala 78:156:@11963.4]
  assign _T_63022 = _T_63021[10:0]; // @[Modules.scala 78:156:@11964.4]
  assign buffer_4_771 = $signed(_T_63022); // @[Modules.scala 78:156:@11965.4]
  assign _T_63024 = $signed(buffer_4_771) + $signed(buffer_4_723); // @[Modules.scala 78:156:@11967.4]
  assign _T_63025 = _T_63024[10:0]; // @[Modules.scala 78:156:@11968.4]
  assign buffer_4_772 = $signed(_T_63025); // @[Modules.scala 78:156:@11969.4]
  assign _T_63027 = $signed(buffer_4_772) + $signed(buffer_4_724); // @[Modules.scala 78:156:@11971.4]
  assign _T_63028 = _T_63027[10:0]; // @[Modules.scala 78:156:@11972.4]
  assign buffer_4_773 = $signed(_T_63028); // @[Modules.scala 78:156:@11973.4]
  assign _T_63030 = $signed(buffer_4_773) + $signed(buffer_4_725); // @[Modules.scala 78:156:@11975.4]
  assign _T_63031 = _T_63030[10:0]; // @[Modules.scala 78:156:@11976.4]
  assign buffer_4_774 = $signed(_T_63031); // @[Modules.scala 78:156:@11977.4]
  assign _T_63033 = $signed(buffer_4_774) + $signed(buffer_4_726); // @[Modules.scala 78:156:@11979.4]
  assign _T_63034 = _T_63033[10:0]; // @[Modules.scala 78:156:@11980.4]
  assign buffer_4_775 = $signed(_T_63034); // @[Modules.scala 78:156:@11981.4]
  assign _T_63036 = $signed(buffer_4_775) + $signed(buffer_4_727); // @[Modules.scala 78:156:@11983.4]
  assign _T_63037 = _T_63036[10:0]; // @[Modules.scala 78:156:@11984.4]
  assign buffer_4_776 = $signed(_T_63037); // @[Modules.scala 78:156:@11985.4]
  assign _T_63039 = $signed(buffer_4_776) + $signed(buffer_4_728); // @[Modules.scala 78:156:@11987.4]
  assign _T_63040 = _T_63039[10:0]; // @[Modules.scala 78:156:@11988.4]
  assign buffer_4_777 = $signed(_T_63040); // @[Modules.scala 78:156:@11989.4]
  assign _T_63042 = $signed(buffer_4_777) + $signed(buffer_4_729); // @[Modules.scala 78:156:@11991.4]
  assign _T_63043 = _T_63042[10:0]; // @[Modules.scala 78:156:@11992.4]
  assign buffer_4_778 = $signed(_T_63043); // @[Modules.scala 78:156:@11993.4]
  assign _T_63045 = $signed(buffer_4_778) + $signed(buffer_4_730); // @[Modules.scala 78:156:@11995.4]
  assign _T_63046 = _T_63045[10:0]; // @[Modules.scala 78:156:@11996.4]
  assign buffer_4_779 = $signed(_T_63046); // @[Modules.scala 78:156:@11997.4]
  assign _T_63048 = $signed(buffer_4_779) + $signed(buffer_4_731); // @[Modules.scala 78:156:@11999.4]
  assign _T_63049 = _T_63048[10:0]; // @[Modules.scala 78:156:@12000.4]
  assign buffer_4_780 = $signed(_T_63049); // @[Modules.scala 78:156:@12001.4]
  assign _T_63051 = $signed(buffer_4_780) + $signed(buffer_0_701); // @[Modules.scala 78:156:@12003.4]
  assign _T_63052 = _T_63051[10:0]; // @[Modules.scala 78:156:@12004.4]
  assign buffer_4_781 = $signed(_T_63052); // @[Modules.scala 78:156:@12005.4]
  assign _T_63054 = $signed(buffer_4_781) + $signed(buffer_4_733); // @[Modules.scala 78:156:@12007.4]
  assign _T_63055 = _T_63054[10:0]; // @[Modules.scala 78:156:@12008.4]
  assign buffer_4_782 = $signed(_T_63055); // @[Modules.scala 78:156:@12009.4]
  assign _T_63057 = $signed(buffer_4_782) + $signed(buffer_4_734); // @[Modules.scala 78:156:@12011.4]
  assign _T_63058 = _T_63057[10:0]; // @[Modules.scala 78:156:@12012.4]
  assign buffer_4_783 = $signed(_T_63058); // @[Modules.scala 78:156:@12013.4]
  assign _T_63098 = $signed(io_in_84) + $signed(io_in_85); // @[Modules.scala 37:46:@12076.4]
  assign _T_63099 = _T_63098[4:0]; // @[Modules.scala 37:46:@12077.4]
  assign _T_63100 = $signed(_T_63099); // @[Modules.scala 37:46:@12078.4]
  assign _T_63118 = $signed(io_in_116) + $signed(io_in_117); // @[Modules.scala 37:46:@12107.4]
  assign _T_63119 = _T_63118[4:0]; // @[Modules.scala 37:46:@12108.4]
  assign _T_63120 = $signed(_T_63119); // @[Modules.scala 37:46:@12109.4]
  assign _T_63141 = $signed(io_in_142) + $signed(io_in_143); // @[Modules.scala 37:46:@12141.4]
  assign _T_63142 = _T_63141[4:0]; // @[Modules.scala 37:46:@12142.4]
  assign _T_63143 = $signed(_T_63142); // @[Modules.scala 37:46:@12143.4]
  assign _T_63177 = $signed(io_in_182) + $signed(io_in_183); // @[Modules.scala 37:46:@12194.4]
  assign _T_63178 = _T_63177[4:0]; // @[Modules.scala 37:46:@12195.4]
  assign _T_63179 = $signed(_T_63178); // @[Modules.scala 37:46:@12196.4]
  assign _T_63180 = $signed(io_in_184) + $signed(io_in_185); // @[Modules.scala 37:46:@12198.4]
  assign _T_63181 = _T_63180[4:0]; // @[Modules.scala 37:46:@12199.4]
  assign _T_63182 = $signed(_T_63181); // @[Modules.scala 37:46:@12200.4]
  assign _T_63206 = $signed(io_in_230) + $signed(io_in_231); // @[Modules.scala 37:46:@12242.4]
  assign _T_63207 = _T_63206[4:0]; // @[Modules.scala 37:46:@12243.4]
  assign _T_63208 = $signed(_T_63207); // @[Modules.scala 37:46:@12244.4]
  assign _T_63253 = $signed(io_in_294) + $signed(io_in_295); // @[Modules.scala 37:46:@12310.4]
  assign _T_63254 = _T_63253[4:0]; // @[Modules.scala 37:46:@12311.4]
  assign _T_63255 = $signed(_T_63254); // @[Modules.scala 37:46:@12312.4]
  assign _T_63259 = $signed(io_in_300) + $signed(io_in_301); // @[Modules.scala 37:46:@12319.4]
  assign _T_63260 = _T_63259[4:0]; // @[Modules.scala 37:46:@12320.4]
  assign _T_63261 = $signed(_T_63260); // @[Modules.scala 37:46:@12321.4]
  assign _T_63269 = $signed(io_in_322) + $signed(io_in_323); // @[Modules.scala 37:46:@12333.4]
  assign _T_63270 = _T_63269[4:0]; // @[Modules.scala 37:46:@12334.4]
  assign _T_63271 = $signed(_T_63270); // @[Modules.scala 37:46:@12335.4]
  assign _T_63272 = $signed(io_in_326) + $signed(io_in_327); // @[Modules.scala 37:46:@12338.4]
  assign _T_63273 = _T_63272[4:0]; // @[Modules.scala 37:46:@12339.4]
  assign _T_63274 = $signed(_T_63273); // @[Modules.scala 37:46:@12340.4]
  assign _T_63278 = $signed(io_in_330) + $signed(io_in_331); // @[Modules.scala 37:46:@12346.4]
  assign _T_63279 = _T_63278[4:0]; // @[Modules.scala 37:46:@12347.4]
  assign _T_63280 = $signed(_T_63279); // @[Modules.scala 37:46:@12348.4]
  assign _T_63282 = $signed(io_in_336) + $signed(io_in_337); // @[Modules.scala 37:46:@12352.4]
  assign _T_63283 = _T_63282[4:0]; // @[Modules.scala 37:46:@12353.4]
  assign _T_63284 = $signed(_T_63283); // @[Modules.scala 37:46:@12354.4]
  assign _T_63425 = $signed(io_in_558) + $signed(io_in_559); // @[Modules.scala 37:46:@12568.4]
  assign _T_63426 = _T_63425[4:0]; // @[Modules.scala 37:46:@12569.4]
  assign _T_63427 = $signed(_T_63426); // @[Modules.scala 37:46:@12570.4]
  assign _T_63560 = $signed(io_in_742) + $signed(io_in_743); // @[Modules.scala 37:46:@12777.4]
  assign _T_63561 = _T_63560[4:0]; // @[Modules.scala 37:46:@12778.4]
  assign _T_63562 = $signed(_T_63561); // @[Modules.scala 37:46:@12779.4]
  assign _T_63572 = $signed(io_in_750) + $signed(io_in_751); // @[Modules.scala 37:46:@12793.4]
  assign _T_63573 = _T_63572[4:0]; // @[Modules.scala 37:46:@12794.4]
  assign _T_63574 = $signed(_T_63573); // @[Modules.scala 37:46:@12795.4]
  assign _T_63596 = $signed(io_in_778) + $signed(io_in_779); // @[Modules.scala 37:46:@12828.4]
  assign _T_63597 = _T_63596[4:0]; // @[Modules.scala 37:46:@12829.4]
  assign _T_63598 = $signed(_T_63597); // @[Modules.scala 37:46:@12830.4]
  assign _T_63602 = $signed(11'sh0) + $signed(buffer_3_1); // @[Modules.scala 65:57:@12837.4]
  assign _T_63603 = _T_63602[10:0]; // @[Modules.scala 65:57:@12838.4]
  assign buffer_5_392 = $signed(_T_63603); // @[Modules.scala 65:57:@12839.4]
  assign _T_63605 = $signed(buffer_2_2) + $signed(buffer_1_3); // @[Modules.scala 65:57:@12841.4]
  assign _T_63606 = _T_63605[10:0]; // @[Modules.scala 65:57:@12842.4]
  assign buffer_5_393 = $signed(_T_63606); // @[Modules.scala 65:57:@12843.4]
  assign _T_63608 = $signed(buffer_0_4) + $signed(buffer_3_5); // @[Modules.scala 65:57:@12845.4]
  assign _T_63609 = _T_63608[10:0]; // @[Modules.scala 65:57:@12846.4]
  assign buffer_5_394 = $signed(_T_63609); // @[Modules.scala 65:57:@12847.4]
  assign buffer_5_10 = {{6{io_in_21[4]}},io_in_21}; // @[Modules.scala 32:22:@8.4]
  assign _T_63617 = $signed(buffer_5_10) + $signed(11'sh0); // @[Modules.scala 65:57:@12857.4]
  assign _T_63618 = _T_63617[10:0]; // @[Modules.scala 65:57:@12858.4]
  assign buffer_5_397 = $signed(_T_63618); // @[Modules.scala 65:57:@12859.4]
  assign _T_63623 = $signed(11'sh0) + $signed(buffer_1_15); // @[Modules.scala 65:57:@12865.4]
  assign _T_63624 = _T_63623[10:0]; // @[Modules.scala 65:57:@12866.4]
  assign buffer_5_399 = $signed(_T_63624); // @[Modules.scala 65:57:@12867.4]
  assign buffer_5_16 = {{6{io_in_33[4]}},io_in_33}; // @[Modules.scala 32:22:@8.4]
  assign _T_63626 = $signed(buffer_5_16) + $signed(11'sh0); // @[Modules.scala 65:57:@12869.4]
  assign _T_63627 = _T_63626[10:0]; // @[Modules.scala 65:57:@12870.4]
  assign buffer_5_400 = $signed(_T_63627); // @[Modules.scala 65:57:@12871.4]
  assign buffer_5_21 = {{6{io_in_43[4]}},io_in_43}; // @[Modules.scala 32:22:@8.4]
  assign _T_63632 = $signed(11'sh0) + $signed(buffer_5_21); // @[Modules.scala 65:57:@12877.4]
  assign _T_63633 = _T_63632[10:0]; // @[Modules.scala 65:57:@12878.4]
  assign buffer_5_402 = $signed(_T_63633); // @[Modules.scala 65:57:@12879.4]
  assign _T_63644 = $signed(buffer_0_28) + $signed(buffer_2_29); // @[Modules.scala 65:57:@12893.4]
  assign _T_63645 = _T_63644[10:0]; // @[Modules.scala 65:57:@12894.4]
  assign buffer_5_406 = $signed(_T_63645); // @[Modules.scala 65:57:@12895.4]
  assign _T_63653 = $signed(11'sh0) + $signed(buffer_2_35); // @[Modules.scala 65:57:@12905.4]
  assign _T_63654 = _T_63653[10:0]; // @[Modules.scala 65:57:@12906.4]
  assign buffer_5_409 = $signed(_T_63654); // @[Modules.scala 65:57:@12907.4]
  assign buffer_5_36 = {{6{io_in_73[4]}},io_in_73}; // @[Modules.scala 32:22:@8.4]
  assign _T_63656 = $signed(buffer_5_36) + $signed(11'sh0); // @[Modules.scala 65:57:@12909.4]
  assign _T_63657 = _T_63656[10:0]; // @[Modules.scala 65:57:@12910.4]
  assign buffer_5_410 = $signed(_T_63657); // @[Modules.scala 65:57:@12911.4]
  assign _T_63662 = $signed(buffer_1_40) + $signed(buffer_0_41); // @[Modules.scala 65:57:@12917.4]
  assign _T_63663 = _T_63662[10:0]; // @[Modules.scala 65:57:@12918.4]
  assign buffer_5_412 = $signed(_T_63663); // @[Modules.scala 65:57:@12919.4]
  assign buffer_5_42 = {{6{_T_63100[4]}},_T_63100}; // @[Modules.scala 32:22:@8.4]
  assign _T_63665 = $signed(buffer_5_42) + $signed(11'sh0); // @[Modules.scala 65:57:@12921.4]
  assign _T_63666 = _T_63665[10:0]; // @[Modules.scala 65:57:@12922.4]
  assign buffer_5_413 = $signed(_T_63666); // @[Modules.scala 65:57:@12923.4]
  assign _T_63677 = $signed(buffer_2_50) + $signed(11'sh0); // @[Modules.scala 65:57:@12937.4]
  assign _T_63678 = _T_63677[10:0]; // @[Modules.scala 65:57:@12938.4]
  assign buffer_5_417 = $signed(_T_63678); // @[Modules.scala 65:57:@12939.4]
  assign _T_63683 = $signed(buffer_3_54) + $signed(11'sh0); // @[Modules.scala 65:57:@12945.4]
  assign _T_63684 = _T_63683[10:0]; // @[Modules.scala 65:57:@12946.4]
  assign buffer_5_419 = $signed(_T_63684); // @[Modules.scala 65:57:@12947.4]
  assign buffer_5_57 = {{6{io_in_114[4]}},io_in_114}; // @[Modules.scala 32:22:@8.4]
  assign _T_63686 = $signed(buffer_0_56) + $signed(buffer_5_57); // @[Modules.scala 65:57:@12949.4]
  assign _T_63687 = _T_63686[10:0]; // @[Modules.scala 65:57:@12950.4]
  assign buffer_5_420 = $signed(_T_63687); // @[Modules.scala 65:57:@12951.4]
  assign buffer_5_58 = {{6{_T_63120[4]}},_T_63120}; // @[Modules.scala 32:22:@8.4]
  assign _T_63689 = $signed(buffer_5_58) + $signed(buffer_0_59); // @[Modules.scala 65:57:@12953.4]
  assign _T_63690 = _T_63689[10:0]; // @[Modules.scala 65:57:@12954.4]
  assign buffer_5_421 = $signed(_T_63690); // @[Modules.scala 65:57:@12955.4]
  assign _T_63698 = $signed(buffer_1_64) + $signed(11'sh0); // @[Modules.scala 65:57:@12965.4]
  assign _T_63699 = _T_63698[10:0]; // @[Modules.scala 65:57:@12966.4]
  assign buffer_5_424 = $signed(_T_63699); // @[Modules.scala 65:57:@12967.4]
  assign buffer_5_66 = {{6{io_in_132[4]}},io_in_132}; // @[Modules.scala 32:22:@8.4]
  assign _T_63701 = $signed(buffer_5_66) + $signed(11'sh0); // @[Modules.scala 65:57:@12969.4]
  assign _T_63702 = _T_63701[10:0]; // @[Modules.scala 65:57:@12970.4]
  assign buffer_5_425 = $signed(_T_63702); // @[Modules.scala 65:57:@12971.4]
  assign buffer_5_68 = {{6{io_in_137[4]}},io_in_137}; // @[Modules.scala 32:22:@8.4]
  assign _T_63704 = $signed(buffer_5_68) + $signed(buffer_3_69); // @[Modules.scala 65:57:@12973.4]
  assign _T_63705 = _T_63704[10:0]; // @[Modules.scala 65:57:@12974.4]
  assign buffer_5_426 = $signed(_T_63705); // @[Modules.scala 65:57:@12975.4]
  assign buffer_5_71 = {{6{_T_63143[4]}},_T_63143}; // @[Modules.scala 32:22:@8.4]
  assign _T_63707 = $signed(buffer_2_70) + $signed(buffer_5_71); // @[Modules.scala 65:57:@12977.4]
  assign _T_63708 = _T_63707[10:0]; // @[Modules.scala 65:57:@12978.4]
  assign buffer_5_427 = $signed(_T_63708); // @[Modules.scala 65:57:@12979.4]
  assign buffer_5_73 = {{6{io_in_147[4]}},io_in_147}; // @[Modules.scala 32:22:@8.4]
  assign _T_63710 = $signed(buffer_4_72) + $signed(buffer_5_73); // @[Modules.scala 65:57:@12981.4]
  assign _T_63711 = _T_63710[10:0]; // @[Modules.scala 65:57:@12982.4]
  assign buffer_5_428 = $signed(_T_63711); // @[Modules.scala 65:57:@12983.4]
  assign buffer_5_80 = {{6{io_in_161[4]}},io_in_161}; // @[Modules.scala 32:22:@8.4]
  assign _T_63722 = $signed(buffer_5_80) + $signed(11'sh0); // @[Modules.scala 65:57:@12997.4]
  assign _T_63723 = _T_63722[10:0]; // @[Modules.scala 65:57:@12998.4]
  assign buffer_5_432 = $signed(_T_63723); // @[Modules.scala 65:57:@12999.4]
  assign buffer_5_82 = {{6{io_in_165[4]}},io_in_165}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_83 = {{6{io_in_166[4]}},io_in_166}; // @[Modules.scala 32:22:@8.4]
  assign _T_63725 = $signed(buffer_5_82) + $signed(buffer_5_83); // @[Modules.scala 65:57:@13001.4]
  assign _T_63726 = _T_63725[10:0]; // @[Modules.scala 65:57:@13002.4]
  assign buffer_5_433 = $signed(_T_63726); // @[Modules.scala 65:57:@13003.4]
  assign _T_63728 = $signed(11'sh0) + $signed(buffer_1_85); // @[Modules.scala 65:57:@13005.4]
  assign _T_63729 = _T_63728[10:0]; // @[Modules.scala 65:57:@13006.4]
  assign buffer_5_434 = $signed(_T_63729); // @[Modules.scala 65:57:@13007.4]
  assign buffer_5_87 = {{6{io_in_174[4]}},io_in_174}; // @[Modules.scala 32:22:@8.4]
  assign _T_63731 = $signed(buffer_3_86) + $signed(buffer_5_87); // @[Modules.scala 65:57:@13009.4]
  assign _T_63732 = _T_63731[10:0]; // @[Modules.scala 65:57:@13010.4]
  assign buffer_5_435 = $signed(_T_63732); // @[Modules.scala 65:57:@13011.4]
  assign buffer_5_91 = {{6{_T_63179[4]}},_T_63179}; // @[Modules.scala 32:22:@8.4]
  assign _T_63737 = $signed(buffer_3_90) + $signed(buffer_5_91); // @[Modules.scala 65:57:@13017.4]
  assign _T_63738 = _T_63737[10:0]; // @[Modules.scala 65:57:@13018.4]
  assign buffer_5_437 = $signed(_T_63738); // @[Modules.scala 65:57:@13019.4]
  assign buffer_5_92 = {{6{_T_63182[4]}},_T_63182}; // @[Modules.scala 32:22:@8.4]
  assign _T_63740 = $signed(buffer_5_92) + $signed(buffer_3_93); // @[Modules.scala 65:57:@13021.4]
  assign _T_63741 = _T_63740[10:0]; // @[Modules.scala 65:57:@13022.4]
  assign buffer_5_438 = $signed(_T_63741); // @[Modules.scala 65:57:@13023.4]
  assign _T_63743 = $signed(buffer_1_94) + $signed(11'sh0); // @[Modules.scala 65:57:@13025.4]
  assign _T_63744 = _T_63743[10:0]; // @[Modules.scala 65:57:@13026.4]
  assign buffer_5_439 = $signed(_T_63744); // @[Modules.scala 65:57:@13027.4]
  assign _T_63746 = $signed(buffer_1_96) + $signed(11'sh0); // @[Modules.scala 65:57:@13029.4]
  assign _T_63747 = _T_63746[10:0]; // @[Modules.scala 65:57:@13030.4]
  assign buffer_5_440 = $signed(_T_63747); // @[Modules.scala 65:57:@13031.4]
  assign buffer_5_101 = {{6{io_in_202[4]}},io_in_202}; // @[Modules.scala 32:22:@8.4]
  assign _T_63752 = $signed(buffer_3_100) + $signed(buffer_5_101); // @[Modules.scala 65:57:@13037.4]
  assign _T_63753 = _T_63752[10:0]; // @[Modules.scala 65:57:@13038.4]
  assign buffer_5_442 = $signed(_T_63753); // @[Modules.scala 65:57:@13039.4]
  assign _T_63755 = $signed(buffer_4_102) + $signed(buffer_0_103); // @[Modules.scala 65:57:@13041.4]
  assign _T_63756 = _T_63755[10:0]; // @[Modules.scala 65:57:@13042.4]
  assign buffer_5_443 = $signed(_T_63756); // @[Modules.scala 65:57:@13043.4]
  assign _T_63758 = $signed(buffer_3_104) + $signed(buffer_0_105); // @[Modules.scala 65:57:@13045.4]
  assign _T_63759 = _T_63758[10:0]; // @[Modules.scala 65:57:@13046.4]
  assign buffer_5_444 = $signed(_T_63759); // @[Modules.scala 65:57:@13047.4]
  assign _T_63761 = $signed(buffer_3_106) + $signed(buffer_1_107); // @[Modules.scala 65:57:@13049.4]
  assign _T_63762 = _T_63761[10:0]; // @[Modules.scala 65:57:@13050.4]
  assign buffer_5_445 = $signed(_T_63762); // @[Modules.scala 65:57:@13051.4]
  assign buffer_5_108 = {{6{io_in_216[4]}},io_in_216}; // @[Modules.scala 32:22:@8.4]
  assign _T_63764 = $signed(buffer_5_108) + $signed(11'sh0); // @[Modules.scala 65:57:@13053.4]
  assign _T_63765 = _T_63764[10:0]; // @[Modules.scala 65:57:@13054.4]
  assign buffer_5_446 = $signed(_T_63765); // @[Modules.scala 65:57:@13055.4]
  assign buffer_5_111 = {{6{io_in_222[4]}},io_in_222}; // @[Modules.scala 32:22:@8.4]
  assign _T_63767 = $signed(11'sh0) + $signed(buffer_5_111); // @[Modules.scala 65:57:@13057.4]
  assign _T_63768 = _T_63767[10:0]; // @[Modules.scala 65:57:@13058.4]
  assign buffer_5_447 = $signed(_T_63768); // @[Modules.scala 65:57:@13059.4]
  assign buffer_5_113 = {{6{io_in_227[4]}},io_in_227}; // @[Modules.scala 32:22:@8.4]
  assign _T_63770 = $signed(11'sh0) + $signed(buffer_5_113); // @[Modules.scala 65:57:@13061.4]
  assign _T_63771 = _T_63770[10:0]; // @[Modules.scala 65:57:@13062.4]
  assign buffer_5_448 = $signed(_T_63771); // @[Modules.scala 65:57:@13063.4]
  assign buffer_5_115 = {{6{_T_63208[4]}},_T_63208}; // @[Modules.scala 32:22:@8.4]
  assign _T_63773 = $signed(buffer_3_114) + $signed(buffer_5_115); // @[Modules.scala 65:57:@13065.4]
  assign _T_63774 = _T_63773[10:0]; // @[Modules.scala 65:57:@13066.4]
  assign buffer_5_449 = $signed(_T_63774); // @[Modules.scala 65:57:@13067.4]
  assign _T_63785 = $signed(buffer_4_122) + $signed(11'sh0); // @[Modules.scala 65:57:@13081.4]
  assign _T_63786 = _T_63785[10:0]; // @[Modules.scala 65:57:@13082.4]
  assign buffer_5_453 = $signed(_T_63786); // @[Modules.scala 65:57:@13083.4]
  assign _T_63788 = $signed(11'sh0) + $signed(buffer_1_125); // @[Modules.scala 65:57:@13085.4]
  assign _T_63789 = _T_63788[10:0]; // @[Modules.scala 65:57:@13086.4]
  assign buffer_5_454 = $signed(_T_63789); // @[Modules.scala 65:57:@13087.4]
  assign buffer_5_126 = {{6{io_in_252[4]}},io_in_252}; // @[Modules.scala 32:22:@8.4]
  assign _T_63791 = $signed(buffer_5_126) + $signed(11'sh0); // @[Modules.scala 65:57:@13089.4]
  assign _T_63792 = _T_63791[10:0]; // @[Modules.scala 65:57:@13090.4]
  assign buffer_5_455 = $signed(_T_63792); // @[Modules.scala 65:57:@13091.4]
  assign _T_63797 = $signed(buffer_2_130) + $signed(11'sh0); // @[Modules.scala 65:57:@13097.4]
  assign _T_63798 = _T_63797[10:0]; // @[Modules.scala 65:57:@13098.4]
  assign buffer_5_457 = $signed(_T_63798); // @[Modules.scala 65:57:@13099.4]
  assign buffer_5_132 = {{6{io_in_265[4]}},io_in_265}; // @[Modules.scala 32:22:@8.4]
  assign _T_63800 = $signed(buffer_5_132) + $signed(buffer_1_133); // @[Modules.scala 65:57:@13101.4]
  assign _T_63801 = _T_63800[10:0]; // @[Modules.scala 65:57:@13102.4]
  assign buffer_5_458 = $signed(_T_63801); // @[Modules.scala 65:57:@13103.4]
  assign buffer_5_135 = {{6{io_in_270[4]}},io_in_270}; // @[Modules.scala 32:22:@8.4]
  assign _T_63803 = $signed(buffer_3_134) + $signed(buffer_5_135); // @[Modules.scala 65:57:@13105.4]
  assign _T_63804 = _T_63803[10:0]; // @[Modules.scala 65:57:@13106.4]
  assign buffer_5_459 = $signed(_T_63804); // @[Modules.scala 65:57:@13107.4]
  assign buffer_5_136 = {{6{io_in_272[4]}},io_in_272}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_137 = {{6{io_in_274[4]}},io_in_274}; // @[Modules.scala 32:22:@8.4]
  assign _T_63806 = $signed(buffer_5_136) + $signed(buffer_5_137); // @[Modules.scala 65:57:@13109.4]
  assign _T_63807 = _T_63806[10:0]; // @[Modules.scala 65:57:@13110.4]
  assign buffer_5_460 = $signed(_T_63807); // @[Modules.scala 65:57:@13111.4]
  assign buffer_5_139 = {{6{io_in_278[4]}},io_in_278}; // @[Modules.scala 32:22:@8.4]
  assign _T_63809 = $signed(11'sh0) + $signed(buffer_5_139); // @[Modules.scala 65:57:@13113.4]
  assign _T_63810 = _T_63809[10:0]; // @[Modules.scala 65:57:@13114.4]
  assign buffer_5_461 = $signed(_T_63810); // @[Modules.scala 65:57:@13115.4]
  assign buffer_5_140 = {{6{io_in_280[4]}},io_in_280}; // @[Modules.scala 32:22:@8.4]
  assign _T_63812 = $signed(buffer_5_140) + $signed(11'sh0); // @[Modules.scala 65:57:@13117.4]
  assign _T_63813 = _T_63812[10:0]; // @[Modules.scala 65:57:@13118.4]
  assign buffer_5_462 = $signed(_T_63813); // @[Modules.scala 65:57:@13119.4]
  assign buffer_5_143 = {{6{io_in_286[4]}},io_in_286}; // @[Modules.scala 32:22:@8.4]
  assign _T_63815 = $signed(11'sh0) + $signed(buffer_5_143); // @[Modules.scala 65:57:@13121.4]
  assign _T_63816 = _T_63815[10:0]; // @[Modules.scala 65:57:@13122.4]
  assign buffer_5_463 = $signed(_T_63816); // @[Modules.scala 65:57:@13123.4]
  assign buffer_5_147 = {{6{_T_63255[4]}},_T_63255}; // @[Modules.scala 32:22:@8.4]
  assign _T_63821 = $signed(11'sh0) + $signed(buffer_5_147); // @[Modules.scala 65:57:@13129.4]
  assign _T_63822 = _T_63821[10:0]; // @[Modules.scala 65:57:@13130.4]
  assign buffer_5_465 = $signed(_T_63822); // @[Modules.scala 65:57:@13131.4]
  assign buffer_5_148 = {{6{io_in_296[4]}},io_in_296}; // @[Modules.scala 32:22:@8.4]
  assign _T_63824 = $signed(buffer_5_148) + $signed(buffer_4_149); // @[Modules.scala 65:57:@13133.4]
  assign _T_63825 = _T_63824[10:0]; // @[Modules.scala 65:57:@13134.4]
  assign buffer_5_466 = $signed(_T_63825); // @[Modules.scala 65:57:@13135.4]
  assign buffer_5_150 = {{6{_T_63261[4]}},_T_63261}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_151 = {{6{io_in_302[4]}},io_in_302}; // @[Modules.scala 32:22:@8.4]
  assign _T_63827 = $signed(buffer_5_150) + $signed(buffer_5_151); // @[Modules.scala 65:57:@13137.4]
  assign _T_63828 = _T_63827[10:0]; // @[Modules.scala 65:57:@13138.4]
  assign buffer_5_467 = $signed(_T_63828); // @[Modules.scala 65:57:@13139.4]
  assign buffer_5_153 = {{6{io_in_307[4]}},io_in_307}; // @[Modules.scala 32:22:@8.4]
  assign _T_63830 = $signed(11'sh0) + $signed(buffer_5_153); // @[Modules.scala 65:57:@13141.4]
  assign _T_63831 = _T_63830[10:0]; // @[Modules.scala 65:57:@13142.4]
  assign buffer_5_468 = $signed(_T_63831); // @[Modules.scala 65:57:@13143.4]
  assign _T_63833 = $signed(buffer_4_154) + $signed(11'sh0); // @[Modules.scala 65:57:@13145.4]
  assign _T_63834 = _T_63833[10:0]; // @[Modules.scala 65:57:@13146.4]
  assign buffer_5_469 = $signed(_T_63834); // @[Modules.scala 65:57:@13147.4]
  assign buffer_5_161 = {{6{_T_63271[4]}},_T_63271}; // @[Modules.scala 32:22:@8.4]
  assign _T_63842 = $signed(11'sh0) + $signed(buffer_5_161); // @[Modules.scala 65:57:@13157.4]
  assign _T_63843 = _T_63842[10:0]; // @[Modules.scala 65:57:@13158.4]
  assign buffer_5_472 = $signed(_T_63843); // @[Modules.scala 65:57:@13159.4]
  assign buffer_5_162 = {{6{io_in_324[4]}},io_in_324}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_163 = {{6{_T_63274[4]}},_T_63274}; // @[Modules.scala 32:22:@8.4]
  assign _T_63845 = $signed(buffer_5_162) + $signed(buffer_5_163); // @[Modules.scala 65:57:@13161.4]
  assign _T_63846 = _T_63845[10:0]; // @[Modules.scala 65:57:@13162.4]
  assign buffer_5_473 = $signed(_T_63846); // @[Modules.scala 65:57:@13163.4]
  assign buffer_5_165 = {{6{_T_63280[4]}},_T_63280}; // @[Modules.scala 32:22:@8.4]
  assign _T_63848 = $signed(buffer_0_164) + $signed(buffer_5_165); // @[Modules.scala 65:57:@13165.4]
  assign _T_63849 = _T_63848[10:0]; // @[Modules.scala 65:57:@13166.4]
  assign buffer_5_474 = $signed(_T_63849); // @[Modules.scala 65:57:@13167.4]
  assign buffer_5_168 = {{6{_T_63284[4]}},_T_63284}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_169 = {{6{io_in_339[4]}},io_in_339}; // @[Modules.scala 32:22:@8.4]
  assign _T_63854 = $signed(buffer_5_168) + $signed(buffer_5_169); // @[Modules.scala 65:57:@13173.4]
  assign _T_63855 = _T_63854[10:0]; // @[Modules.scala 65:57:@13174.4]
  assign buffer_5_476 = $signed(_T_63855); // @[Modules.scala 65:57:@13175.4]
  assign buffer_5_170 = {{6{io_in_340[4]}},io_in_340}; // @[Modules.scala 32:22:@8.4]
  assign _T_63857 = $signed(buffer_5_170) + $signed(11'sh0); // @[Modules.scala 65:57:@13177.4]
  assign _T_63858 = _T_63857[10:0]; // @[Modules.scala 65:57:@13178.4]
  assign buffer_5_477 = $signed(_T_63858); // @[Modules.scala 65:57:@13179.4]
  assign _T_63863 = $signed(11'sh0) + $signed(buffer_0_175); // @[Modules.scala 65:57:@13185.4]
  assign _T_63864 = _T_63863[10:0]; // @[Modules.scala 65:57:@13186.4]
  assign buffer_5_479 = $signed(_T_63864); // @[Modules.scala 65:57:@13187.4]
  assign buffer_5_177 = {{6{io_in_355[4]}},io_in_355}; // @[Modules.scala 32:22:@8.4]
  assign _T_63866 = $signed(buffer_0_176) + $signed(buffer_5_177); // @[Modules.scala 65:57:@13189.4]
  assign _T_63867 = _T_63866[10:0]; // @[Modules.scala 65:57:@13190.4]
  assign buffer_5_480 = $signed(_T_63867); // @[Modules.scala 65:57:@13191.4]
  assign buffer_5_178 = {{6{io_in_356[4]}},io_in_356}; // @[Modules.scala 32:22:@8.4]
  assign _T_63869 = $signed(buffer_5_178) + $signed(11'sh0); // @[Modules.scala 65:57:@13193.4]
  assign _T_63870 = _T_63869[10:0]; // @[Modules.scala 65:57:@13194.4]
  assign buffer_5_481 = $signed(_T_63870); // @[Modules.scala 65:57:@13195.4]
  assign buffer_5_183 = {{6{io_in_367[4]}},io_in_367}; // @[Modules.scala 32:22:@8.4]
  assign _T_63875 = $signed(11'sh0) + $signed(buffer_5_183); // @[Modules.scala 65:57:@13201.4]
  assign _T_63876 = _T_63875[10:0]; // @[Modules.scala 65:57:@13202.4]
  assign buffer_5_483 = $signed(_T_63876); // @[Modules.scala 65:57:@13203.4]
  assign buffer_5_186 = {{6{io_in_372[4]}},io_in_372}; // @[Modules.scala 32:22:@8.4]
  assign _T_63881 = $signed(buffer_5_186) + $signed(11'sh0); // @[Modules.scala 65:57:@13209.4]
  assign _T_63882 = _T_63881[10:0]; // @[Modules.scala 65:57:@13210.4]
  assign buffer_5_485 = $signed(_T_63882); // @[Modules.scala 65:57:@13211.4]
  assign buffer_5_188 = {{6{io_in_377[4]}},io_in_377}; // @[Modules.scala 32:22:@8.4]
  assign _T_63884 = $signed(buffer_5_188) + $signed(buffer_0_189); // @[Modules.scala 65:57:@13213.4]
  assign _T_63885 = _T_63884[10:0]; // @[Modules.scala 65:57:@13214.4]
  assign buffer_5_486 = $signed(_T_63885); // @[Modules.scala 65:57:@13215.4]
  assign buffer_5_194 = {{6{io_in_389[4]}},io_in_389}; // @[Modules.scala 32:22:@8.4]
  assign _T_63893 = $signed(buffer_5_194) + $signed(buffer_3_195); // @[Modules.scala 65:57:@13225.4]
  assign _T_63894 = _T_63893[10:0]; // @[Modules.scala 65:57:@13226.4]
  assign buffer_5_489 = $signed(_T_63894); // @[Modules.scala 65:57:@13227.4]
  assign buffer_5_197 = {{6{io_in_395[4]}},io_in_395}; // @[Modules.scala 32:22:@8.4]
  assign _T_63896 = $signed(11'sh0) + $signed(buffer_5_197); // @[Modules.scala 65:57:@13229.4]
  assign _T_63897 = _T_63896[10:0]; // @[Modules.scala 65:57:@13230.4]
  assign buffer_5_490 = $signed(_T_63897); // @[Modules.scala 65:57:@13231.4]
  assign _T_63914 = $signed(11'sh0) + $signed(buffer_3_209); // @[Modules.scala 65:57:@13253.4]
  assign _T_63915 = _T_63914[10:0]; // @[Modules.scala 65:57:@13254.4]
  assign buffer_5_496 = $signed(_T_63915); // @[Modules.scala 65:57:@13255.4]
  assign buffer_5_211 = {{6{io_in_423[4]}},io_in_423}; // @[Modules.scala 32:22:@8.4]
  assign _T_63917 = $signed(11'sh0) + $signed(buffer_5_211); // @[Modules.scala 65:57:@13257.4]
  assign _T_63918 = _T_63917[10:0]; // @[Modules.scala 65:57:@13258.4]
  assign buffer_5_497 = $signed(_T_63918); // @[Modules.scala 65:57:@13259.4]
  assign buffer_5_212 = {{6{io_in_424[4]}},io_in_424}; // @[Modules.scala 32:22:@8.4]
  assign _T_63920 = $signed(buffer_5_212) + $signed(buffer_3_213); // @[Modules.scala 65:57:@13261.4]
  assign _T_63921 = _T_63920[10:0]; // @[Modules.scala 65:57:@13262.4]
  assign buffer_5_498 = $signed(_T_63921); // @[Modules.scala 65:57:@13263.4]
  assign buffer_5_218 = {{6{io_in_437[4]}},io_in_437}; // @[Modules.scala 32:22:@8.4]
  assign _T_63929 = $signed(buffer_5_218) + $signed(11'sh0); // @[Modules.scala 65:57:@13273.4]
  assign _T_63930 = _T_63929[10:0]; // @[Modules.scala 65:57:@13274.4]
  assign buffer_5_501 = $signed(_T_63930); // @[Modules.scala 65:57:@13275.4]
  assign buffer_5_222 = {{6{io_in_445[4]}},io_in_445}; // @[Modules.scala 32:22:@8.4]
  assign _T_63935 = $signed(buffer_5_222) + $signed(buffer_3_223); // @[Modules.scala 65:57:@13281.4]
  assign _T_63936 = _T_63935[10:0]; // @[Modules.scala 65:57:@13282.4]
  assign buffer_5_503 = $signed(_T_63936); // @[Modules.scala 65:57:@13283.4]
  assign _T_63941 = $signed(buffer_3_226) + $signed(11'sh0); // @[Modules.scala 65:57:@13289.4]
  assign _T_63942 = _T_63941[10:0]; // @[Modules.scala 65:57:@13290.4]
  assign buffer_5_505 = $signed(_T_63942); // @[Modules.scala 65:57:@13291.4]
  assign buffer_5_231 = {{6{io_in_462[4]}},io_in_462}; // @[Modules.scala 32:22:@8.4]
  assign _T_63947 = $signed(buffer_2_230) + $signed(buffer_5_231); // @[Modules.scala 65:57:@13297.4]
  assign _T_63948 = _T_63947[10:0]; // @[Modules.scala 65:57:@13298.4]
  assign buffer_5_507 = $signed(_T_63948); // @[Modules.scala 65:57:@13299.4]
  assign buffer_5_232 = {{6{io_in_464[4]}},io_in_464}; // @[Modules.scala 32:22:@8.4]
  assign _T_63950 = $signed(buffer_5_232) + $signed(11'sh0); // @[Modules.scala 65:57:@13301.4]
  assign _T_63951 = _T_63950[10:0]; // @[Modules.scala 65:57:@13302.4]
  assign buffer_5_508 = $signed(_T_63951); // @[Modules.scala 65:57:@13303.4]
  assign buffer_5_236 = {{6{io_in_473[4]}},io_in_473}; // @[Modules.scala 32:22:@8.4]
  assign _T_63956 = $signed(buffer_5_236) + $signed(buffer_3_237); // @[Modules.scala 65:57:@13309.4]
  assign _T_63957 = _T_63956[10:0]; // @[Modules.scala 65:57:@13310.4]
  assign buffer_5_510 = $signed(_T_63957); // @[Modules.scala 65:57:@13311.4]
  assign _T_63962 = $signed(buffer_3_240) + $signed(11'sh0); // @[Modules.scala 65:57:@13317.4]
  assign _T_63963 = _T_63962[10:0]; // @[Modules.scala 65:57:@13318.4]
  assign buffer_5_512 = $signed(_T_63963); // @[Modules.scala 65:57:@13319.4]
  assign buffer_5_242 = {{6{io_in_484[4]}},io_in_484}; // @[Modules.scala 32:22:@8.4]
  assign _T_63965 = $signed(buffer_5_242) + $signed(11'sh0); // @[Modules.scala 65:57:@13321.4]
  assign _T_63966 = _T_63965[10:0]; // @[Modules.scala 65:57:@13322.4]
  assign buffer_5_513 = $signed(_T_63966); // @[Modules.scala 65:57:@13323.4]
  assign _T_63971 = $signed(11'sh0) + $signed(buffer_4_247); // @[Modules.scala 65:57:@13329.4]
  assign _T_63972 = _T_63971[10:0]; // @[Modules.scala 65:57:@13330.4]
  assign buffer_5_515 = $signed(_T_63972); // @[Modules.scala 65:57:@13331.4]
  assign buffer_5_255 = {{6{io_in_510[4]}},io_in_510}; // @[Modules.scala 32:22:@8.4]
  assign _T_63983 = $signed(buffer_3_254) + $signed(buffer_5_255); // @[Modules.scala 65:57:@13345.4]
  assign _T_63984 = _T_63983[10:0]; // @[Modules.scala 65:57:@13346.4]
  assign buffer_5_519 = $signed(_T_63984); // @[Modules.scala 65:57:@13347.4]
  assign buffer_5_256 = {{6{io_in_513[4]}},io_in_513}; // @[Modules.scala 32:22:@8.4]
  assign _T_63986 = $signed(buffer_5_256) + $signed(buffer_0_257); // @[Modules.scala 65:57:@13349.4]
  assign _T_63987 = _T_63986[10:0]; // @[Modules.scala 65:57:@13350.4]
  assign buffer_5_520 = $signed(_T_63987); // @[Modules.scala 65:57:@13351.4]
  assign _T_63989 = $signed(buffer_2_258) + $signed(buffer_0_259); // @[Modules.scala 65:57:@13353.4]
  assign _T_63990 = _T_63989[10:0]; // @[Modules.scala 65:57:@13354.4]
  assign buffer_5_521 = $signed(_T_63990); // @[Modules.scala 65:57:@13355.4]
  assign _T_63992 = $signed(buffer_1_260) + $signed(buffer_0_261); // @[Modules.scala 65:57:@13357.4]
  assign _T_63993 = _T_63992[10:0]; // @[Modules.scala 65:57:@13358.4]
  assign buffer_5_522 = $signed(_T_63993); // @[Modules.scala 65:57:@13359.4]
  assign buffer_5_268 = {{6{io_in_536[4]}},io_in_536}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_269 = {{6{io_in_539[4]}},io_in_539}; // @[Modules.scala 32:22:@8.4]
  assign _T_64004 = $signed(buffer_5_268) + $signed(buffer_5_269); // @[Modules.scala 65:57:@13373.4]
  assign _T_64005 = _T_64004[10:0]; // @[Modules.scala 65:57:@13374.4]
  assign buffer_5_526 = $signed(_T_64005); // @[Modules.scala 65:57:@13375.4]
  assign buffer_5_270 = {{6{io_in_541[4]}},io_in_541}; // @[Modules.scala 32:22:@8.4]
  assign _T_64007 = $signed(buffer_5_270) + $signed(11'sh0); // @[Modules.scala 65:57:@13377.4]
  assign _T_64008 = _T_64007[10:0]; // @[Modules.scala 65:57:@13378.4]
  assign buffer_5_527 = $signed(_T_64008); // @[Modules.scala 65:57:@13379.4]
  assign _T_64010 = $signed(11'sh0) + $signed(buffer_1_273); // @[Modules.scala 65:57:@13381.4]
  assign _T_64011 = _T_64010[10:0]; // @[Modules.scala 65:57:@13382.4]
  assign buffer_5_528 = $signed(_T_64011); // @[Modules.scala 65:57:@13383.4]
  assign _T_64013 = $signed(buffer_2_274) + $signed(buffer_1_275); // @[Modules.scala 65:57:@13385.4]
  assign _T_64014 = _T_64013[10:0]; // @[Modules.scala 65:57:@13386.4]
  assign buffer_5_529 = $signed(_T_64014); // @[Modules.scala 65:57:@13387.4]
  assign buffer_5_277 = {{6{io_in_555[4]}},io_in_555}; // @[Modules.scala 32:22:@8.4]
  assign _T_64016 = $signed(buffer_0_276) + $signed(buffer_5_277); // @[Modules.scala 65:57:@13389.4]
  assign _T_64017 = _T_64016[10:0]; // @[Modules.scala 65:57:@13390.4]
  assign buffer_5_530 = $signed(_T_64017); // @[Modules.scala 65:57:@13391.4]
  assign buffer_5_279 = {{6{_T_63427[4]}},_T_63427}; // @[Modules.scala 32:22:@8.4]
  assign _T_64019 = $signed(buffer_3_278) + $signed(buffer_5_279); // @[Modules.scala 65:57:@13393.4]
  assign _T_64020 = _T_64019[10:0]; // @[Modules.scala 65:57:@13394.4]
  assign buffer_5_531 = $signed(_T_64020); // @[Modules.scala 65:57:@13395.4]
  assign buffer_5_281 = {{6{io_in_563[4]}},io_in_563}; // @[Modules.scala 32:22:@8.4]
  assign _T_64022 = $signed(11'sh0) + $signed(buffer_5_281); // @[Modules.scala 65:57:@13397.4]
  assign _T_64023 = _T_64022[10:0]; // @[Modules.scala 65:57:@13398.4]
  assign buffer_5_532 = $signed(_T_64023); // @[Modules.scala 65:57:@13399.4]
  assign buffer_5_282 = {{6{io_in_564[4]}},io_in_564}; // @[Modules.scala 32:22:@8.4]
  assign _T_64025 = $signed(buffer_5_282) + $signed(buffer_3_283); // @[Modules.scala 65:57:@13401.4]
  assign _T_64026 = _T_64025[10:0]; // @[Modules.scala 65:57:@13402.4]
  assign buffer_5_533 = $signed(_T_64026); // @[Modules.scala 65:57:@13403.4]
  assign buffer_5_289 = {{6{io_in_579[4]}},io_in_579}; // @[Modules.scala 32:22:@8.4]
  assign _T_64034 = $signed(11'sh0) + $signed(buffer_5_289); // @[Modules.scala 65:57:@13413.4]
  assign _T_64035 = _T_64034[10:0]; // @[Modules.scala 65:57:@13414.4]
  assign buffer_5_536 = $signed(_T_64035); // @[Modules.scala 65:57:@13415.4]
  assign buffer_5_290 = {{6{io_in_581[4]}},io_in_581}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_291 = {{6{io_in_583[4]}},io_in_583}; // @[Modules.scala 32:22:@8.4]
  assign _T_64037 = $signed(buffer_5_290) + $signed(buffer_5_291); // @[Modules.scala 65:57:@13417.4]
  assign _T_64038 = _T_64037[10:0]; // @[Modules.scala 65:57:@13418.4]
  assign buffer_5_537 = $signed(_T_64038); // @[Modules.scala 65:57:@13419.4]
  assign _T_64049 = $signed(buffer_2_298) + $signed(11'sh0); // @[Modules.scala 65:57:@13433.4]
  assign _T_64050 = _T_64049[10:0]; // @[Modules.scala 65:57:@13434.4]
  assign buffer_5_541 = $signed(_T_64050); // @[Modules.scala 65:57:@13435.4]
  assign buffer_5_302 = {{6{io_in_604[4]}},io_in_604}; // @[Modules.scala 32:22:@8.4]
  assign _T_64055 = $signed(buffer_5_302) + $signed(buffer_0_303); // @[Modules.scala 65:57:@13441.4]
  assign _T_64056 = _T_64055[10:0]; // @[Modules.scala 65:57:@13442.4]
  assign buffer_5_543 = $signed(_T_64056); // @[Modules.scala 65:57:@13443.4]
  assign buffer_5_313 = {{6{io_in_626[4]}},io_in_626}; // @[Modules.scala 32:22:@8.4]
  assign _T_64070 = $signed(11'sh0) + $signed(buffer_5_313); // @[Modules.scala 65:57:@13461.4]
  assign _T_64071 = _T_64070[10:0]; // @[Modules.scala 65:57:@13462.4]
  assign buffer_5_548 = $signed(_T_64071); // @[Modules.scala 65:57:@13463.4]
  assign buffer_5_314 = {{6{io_in_628[4]}},io_in_628}; // @[Modules.scala 32:22:@8.4]
  assign _T_64073 = $signed(buffer_5_314) + $signed(buffer_3_315); // @[Modules.scala 65:57:@13465.4]
  assign _T_64074 = _T_64073[10:0]; // @[Modules.scala 65:57:@13466.4]
  assign buffer_5_549 = $signed(_T_64074); // @[Modules.scala 65:57:@13467.4]
  assign _T_64076 = $signed(buffer_3_316) + $signed(11'sh0); // @[Modules.scala 65:57:@13469.4]
  assign _T_64077 = _T_64076[10:0]; // @[Modules.scala 65:57:@13470.4]
  assign buffer_5_550 = $signed(_T_64077); // @[Modules.scala 65:57:@13471.4]
  assign buffer_5_320 = {{6{io_in_640[4]}},io_in_640}; // @[Modules.scala 32:22:@8.4]
  assign _T_64082 = $signed(buffer_5_320) + $signed(buffer_0_321); // @[Modules.scala 65:57:@13477.4]
  assign _T_64083 = _T_64082[10:0]; // @[Modules.scala 65:57:@13478.4]
  assign buffer_5_552 = $signed(_T_64083); // @[Modules.scala 65:57:@13479.4]
  assign _T_64088 = $signed(buffer_4_324) + $signed(buffer_1_325); // @[Modules.scala 65:57:@13485.4]
  assign _T_64089 = _T_64088[10:0]; // @[Modules.scala 65:57:@13486.4]
  assign buffer_5_554 = $signed(_T_64089); // @[Modules.scala 65:57:@13487.4]
  assign buffer_5_326 = {{6{io_in_652[4]}},io_in_652}; // @[Modules.scala 32:22:@8.4]
  assign _T_64091 = $signed(buffer_5_326) + $signed(11'sh0); // @[Modules.scala 65:57:@13489.4]
  assign _T_64092 = _T_64091[10:0]; // @[Modules.scala 65:57:@13490.4]
  assign buffer_5_555 = $signed(_T_64092); // @[Modules.scala 65:57:@13491.4]
  assign buffer_5_328 = {{6{io_in_657[4]}},io_in_657}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_329 = {{6{io_in_658[4]}},io_in_658}; // @[Modules.scala 32:22:@8.4]
  assign _T_64094 = $signed(buffer_5_328) + $signed(buffer_5_329); // @[Modules.scala 65:57:@13493.4]
  assign _T_64095 = _T_64094[10:0]; // @[Modules.scala 65:57:@13494.4]
  assign buffer_5_556 = $signed(_T_64095); // @[Modules.scala 65:57:@13495.4]
  assign _T_64097 = $signed(buffer_2_330) + $signed(buffer_0_331); // @[Modules.scala 65:57:@13497.4]
  assign _T_64098 = _T_64097[10:0]; // @[Modules.scala 65:57:@13498.4]
  assign buffer_5_557 = $signed(_T_64098); // @[Modules.scala 65:57:@13499.4]
  assign buffer_5_332 = {{6{io_in_665[4]}},io_in_665}; // @[Modules.scala 32:22:@8.4]
  assign _T_64100 = $signed(buffer_5_332) + $signed(buffer_0_333); // @[Modules.scala 65:57:@13501.4]
  assign _T_64101 = _T_64100[10:0]; // @[Modules.scala 65:57:@13502.4]
  assign buffer_5_558 = $signed(_T_64101); // @[Modules.scala 65:57:@13503.4]
  assign _T_64106 = $signed(buffer_0_336) + $signed(buffer_1_337); // @[Modules.scala 65:57:@13509.4]
  assign _T_64107 = _T_64106[10:0]; // @[Modules.scala 65:57:@13510.4]
  assign buffer_5_560 = $signed(_T_64107); // @[Modules.scala 65:57:@13511.4]
  assign buffer_5_339 = {{6{io_in_678[4]}},io_in_678}; // @[Modules.scala 32:22:@8.4]
  assign _T_64109 = $signed(buffer_0_338) + $signed(buffer_5_339); // @[Modules.scala 65:57:@13513.4]
  assign _T_64110 = _T_64109[10:0]; // @[Modules.scala 65:57:@13514.4]
  assign buffer_5_561 = $signed(_T_64110); // @[Modules.scala 65:57:@13515.4]
  assign buffer_5_340 = {{6{io_in_680[4]}},io_in_680}; // @[Modules.scala 32:22:@8.4]
  assign buffer_5_341 = {{6{io_in_683[4]}},io_in_683}; // @[Modules.scala 32:22:@8.4]
  assign _T_64112 = $signed(buffer_5_340) + $signed(buffer_5_341); // @[Modules.scala 65:57:@13517.4]
  assign _T_64113 = _T_64112[10:0]; // @[Modules.scala 65:57:@13518.4]
  assign buffer_5_562 = $signed(_T_64113); // @[Modules.scala 65:57:@13519.4]
  assign buffer_5_343 = {{6{io_in_687[4]}},io_in_687}; // @[Modules.scala 32:22:@8.4]
  assign _T_64115 = $signed(buffer_3_342) + $signed(buffer_5_343); // @[Modules.scala 65:57:@13521.4]
  assign _T_64116 = _T_64115[10:0]; // @[Modules.scala 65:57:@13522.4]
  assign buffer_5_563 = $signed(_T_64116); // @[Modules.scala 65:57:@13523.4]
  assign _T_64124 = $signed(buffer_1_348) + $signed(buffer_3_349); // @[Modules.scala 65:57:@13533.4]
  assign _T_64125 = _T_64124[10:0]; // @[Modules.scala 65:57:@13534.4]
  assign buffer_5_566 = $signed(_T_64125); // @[Modules.scala 65:57:@13535.4]
  assign buffer_5_350 = {{6{io_in_700[4]}},io_in_700}; // @[Modules.scala 32:22:@8.4]
  assign _T_64127 = $signed(buffer_5_350) + $signed(11'sh0); // @[Modules.scala 65:57:@13537.4]
  assign _T_64128 = _T_64127[10:0]; // @[Modules.scala 65:57:@13538.4]
  assign buffer_5_567 = $signed(_T_64128); // @[Modules.scala 65:57:@13539.4]
  assign buffer_5_352 = {{6{io_in_705[4]}},io_in_705}; // @[Modules.scala 32:22:@8.4]
  assign _T_64130 = $signed(buffer_5_352) + $signed(buffer_0_353); // @[Modules.scala 65:57:@13541.4]
  assign _T_64131 = _T_64130[10:0]; // @[Modules.scala 65:57:@13542.4]
  assign buffer_5_568 = $signed(_T_64131); // @[Modules.scala 65:57:@13543.4]
  assign buffer_5_361 = {{6{io_in_722[4]}},io_in_722}; // @[Modules.scala 32:22:@8.4]
  assign _T_64142 = $signed(buffer_0_360) + $signed(buffer_5_361); // @[Modules.scala 65:57:@13557.4]
  assign _T_64143 = _T_64142[10:0]; // @[Modules.scala 65:57:@13558.4]
  assign buffer_5_572 = $signed(_T_64143); // @[Modules.scala 65:57:@13559.4]
  assign buffer_5_367 = {{6{io_in_734[4]}},io_in_734}; // @[Modules.scala 32:22:@8.4]
  assign _T_64151 = $signed(buffer_0_366) + $signed(buffer_5_367); // @[Modules.scala 65:57:@13569.4]
  assign _T_64152 = _T_64151[10:0]; // @[Modules.scala 65:57:@13570.4]
  assign buffer_5_575 = $signed(_T_64152); // @[Modules.scala 65:57:@13571.4]
  assign buffer_5_371 = {{6{_T_63562[4]}},_T_63562}; // @[Modules.scala 32:22:@8.4]
  assign _T_64157 = $signed(buffer_3_370) + $signed(buffer_5_371); // @[Modules.scala 65:57:@13577.4]
  assign _T_64158 = _T_64157[10:0]; // @[Modules.scala 65:57:@13578.4]
  assign buffer_5_577 = $signed(_T_64158); // @[Modules.scala 65:57:@13579.4]
  assign buffer_5_375 = {{6{_T_63574[4]}},_T_63574}; // @[Modules.scala 32:22:@8.4]
  assign _T_64163 = $signed(buffer_0_374) + $signed(buffer_5_375); // @[Modules.scala 65:57:@13585.4]
  assign _T_64164 = _T_64163[10:0]; // @[Modules.scala 65:57:@13586.4]
  assign buffer_5_579 = $signed(_T_64164); // @[Modules.scala 65:57:@13587.4]
  assign buffer_5_383 = {{6{io_in_766[4]}},io_in_766}; // @[Modules.scala 32:22:@8.4]
  assign _T_64175 = $signed(11'sh0) + $signed(buffer_5_383); // @[Modules.scala 65:57:@13601.4]
  assign _T_64176 = _T_64175[10:0]; // @[Modules.scala 65:57:@13602.4]
  assign buffer_5_583 = $signed(_T_64176); // @[Modules.scala 65:57:@13603.4]
  assign buffer_5_389 = {{6{_T_63598[4]}},_T_63598}; // @[Modules.scala 32:22:@8.4]
  assign _T_64184 = $signed(buffer_0_388) + $signed(buffer_5_389); // @[Modules.scala 65:57:@13613.4]
  assign _T_64185 = _T_64184[10:0]; // @[Modules.scala 65:57:@13614.4]
  assign buffer_5_586 = $signed(_T_64185); // @[Modules.scala 65:57:@13615.4]
  assign _T_64190 = $signed(buffer_5_392) + $signed(buffer_5_393); // @[Modules.scala 68:83:@13621.4]
  assign _T_64191 = _T_64190[10:0]; // @[Modules.scala 68:83:@13622.4]
  assign buffer_5_588 = $signed(_T_64191); // @[Modules.scala 68:83:@13623.4]
  assign _T_64193 = $signed(buffer_5_394) + $signed(buffer_4_395); // @[Modules.scala 68:83:@13625.4]
  assign _T_64194 = _T_64193[10:0]; // @[Modules.scala 68:83:@13626.4]
  assign buffer_5_589 = $signed(_T_64194); // @[Modules.scala 68:83:@13627.4]
  assign _T_64196 = $signed(buffer_0_396) + $signed(buffer_5_397); // @[Modules.scala 68:83:@13629.4]
  assign _T_64197 = _T_64196[10:0]; // @[Modules.scala 68:83:@13630.4]
  assign buffer_5_590 = $signed(_T_64197); // @[Modules.scala 68:83:@13631.4]
  assign _T_64199 = $signed(buffer_4_398) + $signed(buffer_5_399); // @[Modules.scala 68:83:@13633.4]
  assign _T_64200 = _T_64199[10:0]; // @[Modules.scala 68:83:@13634.4]
  assign buffer_5_591 = $signed(_T_64200); // @[Modules.scala 68:83:@13635.4]
  assign _T_64202 = $signed(buffer_5_400) + $signed(buffer_0_395); // @[Modules.scala 68:83:@13637.4]
  assign _T_64203 = _T_64202[10:0]; // @[Modules.scala 68:83:@13638.4]
  assign buffer_5_592 = $signed(_T_64203); // @[Modules.scala 68:83:@13639.4]
  assign _T_64205 = $signed(buffer_5_402) + $signed(buffer_4_403); // @[Modules.scala 68:83:@13641.4]
  assign _T_64206 = _T_64205[10:0]; // @[Modules.scala 68:83:@13642.4]
  assign buffer_5_593 = $signed(_T_64206); // @[Modules.scala 68:83:@13643.4]
  assign _T_64208 = $signed(buffer_0_395) + $signed(buffer_4_405); // @[Modules.scala 68:83:@13645.4]
  assign _T_64209 = _T_64208[10:0]; // @[Modules.scala 68:83:@13646.4]
  assign buffer_5_594 = $signed(_T_64209); // @[Modules.scala 68:83:@13647.4]
  assign _T_64211 = $signed(buffer_5_406) + $signed(buffer_3_407); // @[Modules.scala 68:83:@13649.4]
  assign _T_64212 = _T_64211[10:0]; // @[Modules.scala 68:83:@13650.4]
  assign buffer_5_595 = $signed(_T_64212); // @[Modules.scala 68:83:@13651.4]
  assign _T_64214 = $signed(buffer_0_395) + $signed(buffer_5_409); // @[Modules.scala 68:83:@13653.4]
  assign _T_64215 = _T_64214[10:0]; // @[Modules.scala 68:83:@13654.4]
  assign buffer_5_596 = $signed(_T_64215); // @[Modules.scala 68:83:@13655.4]
  assign _T_64217 = $signed(buffer_5_410) + $signed(buffer_0_395); // @[Modules.scala 68:83:@13657.4]
  assign _T_64218 = _T_64217[10:0]; // @[Modules.scala 68:83:@13658.4]
  assign buffer_5_597 = $signed(_T_64218); // @[Modules.scala 68:83:@13659.4]
  assign _T_64220 = $signed(buffer_5_412) + $signed(buffer_5_413); // @[Modules.scala 68:83:@13661.4]
  assign _T_64221 = _T_64220[10:0]; // @[Modules.scala 68:83:@13662.4]
  assign buffer_5_598 = $signed(_T_64221); // @[Modules.scala 68:83:@13663.4]
  assign _T_64226 = $signed(buffer_3_416) + $signed(buffer_5_417); // @[Modules.scala 68:83:@13669.4]
  assign _T_64227 = _T_64226[10:0]; // @[Modules.scala 68:83:@13670.4]
  assign buffer_5_600 = $signed(_T_64227); // @[Modules.scala 68:83:@13671.4]
  assign _T_64229 = $signed(buffer_0_395) + $signed(buffer_5_419); // @[Modules.scala 68:83:@13673.4]
  assign _T_64230 = _T_64229[10:0]; // @[Modules.scala 68:83:@13674.4]
  assign buffer_5_601 = $signed(_T_64230); // @[Modules.scala 68:83:@13675.4]
  assign _T_64232 = $signed(buffer_5_420) + $signed(buffer_5_421); // @[Modules.scala 68:83:@13677.4]
  assign _T_64233 = _T_64232[10:0]; // @[Modules.scala 68:83:@13678.4]
  assign buffer_5_602 = $signed(_T_64233); // @[Modules.scala 68:83:@13679.4]
  assign _T_64238 = $signed(buffer_5_424) + $signed(buffer_5_425); // @[Modules.scala 68:83:@13685.4]
  assign _T_64239 = _T_64238[10:0]; // @[Modules.scala 68:83:@13686.4]
  assign buffer_5_604 = $signed(_T_64239); // @[Modules.scala 68:83:@13687.4]
  assign _T_64241 = $signed(buffer_5_426) + $signed(buffer_5_427); // @[Modules.scala 68:83:@13689.4]
  assign _T_64242 = _T_64241[10:0]; // @[Modules.scala 68:83:@13690.4]
  assign buffer_5_605 = $signed(_T_64242); // @[Modules.scala 68:83:@13691.4]
  assign _T_64244 = $signed(buffer_5_428) + $signed(buffer_3_429); // @[Modules.scala 68:83:@13693.4]
  assign _T_64245 = _T_64244[10:0]; // @[Modules.scala 68:83:@13694.4]
  assign buffer_5_606 = $signed(_T_64245); // @[Modules.scala 68:83:@13695.4]
  assign _T_64247 = $signed(buffer_4_430) + $signed(buffer_1_431); // @[Modules.scala 68:83:@13697.4]
  assign _T_64248 = _T_64247[10:0]; // @[Modules.scala 68:83:@13698.4]
  assign buffer_5_607 = $signed(_T_64248); // @[Modules.scala 68:83:@13699.4]
  assign _T_64250 = $signed(buffer_5_432) + $signed(buffer_5_433); // @[Modules.scala 68:83:@13701.4]
  assign _T_64251 = _T_64250[10:0]; // @[Modules.scala 68:83:@13702.4]
  assign buffer_5_608 = $signed(_T_64251); // @[Modules.scala 68:83:@13703.4]
  assign _T_64253 = $signed(buffer_5_434) + $signed(buffer_5_435); // @[Modules.scala 68:83:@13705.4]
  assign _T_64254 = _T_64253[10:0]; // @[Modules.scala 68:83:@13706.4]
  assign buffer_5_609 = $signed(_T_64254); // @[Modules.scala 68:83:@13707.4]
  assign _T_64256 = $signed(buffer_3_436) + $signed(buffer_5_437); // @[Modules.scala 68:83:@13709.4]
  assign _T_64257 = _T_64256[10:0]; // @[Modules.scala 68:83:@13710.4]
  assign buffer_5_610 = $signed(_T_64257); // @[Modules.scala 68:83:@13711.4]
  assign _T_64259 = $signed(buffer_5_438) + $signed(buffer_5_439); // @[Modules.scala 68:83:@13713.4]
  assign _T_64260 = _T_64259[10:0]; // @[Modules.scala 68:83:@13714.4]
  assign buffer_5_611 = $signed(_T_64260); // @[Modules.scala 68:83:@13715.4]
  assign _T_64262 = $signed(buffer_5_440) + $signed(buffer_3_441); // @[Modules.scala 68:83:@13717.4]
  assign _T_64263 = _T_64262[10:0]; // @[Modules.scala 68:83:@13718.4]
  assign buffer_5_612 = $signed(_T_64263); // @[Modules.scala 68:83:@13719.4]
  assign _T_64265 = $signed(buffer_5_442) + $signed(buffer_5_443); // @[Modules.scala 68:83:@13721.4]
  assign _T_64266 = _T_64265[10:0]; // @[Modules.scala 68:83:@13722.4]
  assign buffer_5_613 = $signed(_T_64266); // @[Modules.scala 68:83:@13723.4]
  assign _T_64268 = $signed(buffer_5_444) + $signed(buffer_5_445); // @[Modules.scala 68:83:@13725.4]
  assign _T_64269 = _T_64268[10:0]; // @[Modules.scala 68:83:@13726.4]
  assign buffer_5_614 = $signed(_T_64269); // @[Modules.scala 68:83:@13727.4]
  assign _T_64271 = $signed(buffer_5_446) + $signed(buffer_5_447); // @[Modules.scala 68:83:@13729.4]
  assign _T_64272 = _T_64271[10:0]; // @[Modules.scala 68:83:@13730.4]
  assign buffer_5_615 = $signed(_T_64272); // @[Modules.scala 68:83:@13731.4]
  assign _T_64274 = $signed(buffer_5_448) + $signed(buffer_5_449); // @[Modules.scala 68:83:@13733.4]
  assign _T_64275 = _T_64274[10:0]; // @[Modules.scala 68:83:@13734.4]
  assign buffer_5_616 = $signed(_T_64275); // @[Modules.scala 68:83:@13735.4]
  assign _T_64277 = $signed(buffer_4_450) + $signed(buffer_3_451); // @[Modules.scala 68:83:@13737.4]
  assign _T_64278 = _T_64277[10:0]; // @[Modules.scala 68:83:@13738.4]
  assign buffer_5_617 = $signed(_T_64278); // @[Modules.scala 68:83:@13739.4]
  assign _T_64280 = $signed(buffer_3_452) + $signed(buffer_5_453); // @[Modules.scala 68:83:@13741.4]
  assign _T_64281 = _T_64280[10:0]; // @[Modules.scala 68:83:@13742.4]
  assign buffer_5_618 = $signed(_T_64281); // @[Modules.scala 68:83:@13743.4]
  assign _T_64283 = $signed(buffer_5_454) + $signed(buffer_5_455); // @[Modules.scala 68:83:@13745.4]
  assign _T_64284 = _T_64283[10:0]; // @[Modules.scala 68:83:@13746.4]
  assign buffer_5_619 = $signed(_T_64284); // @[Modules.scala 68:83:@13747.4]
  assign _T_64286 = $signed(buffer_3_456) + $signed(buffer_5_457); // @[Modules.scala 68:83:@13749.4]
  assign _T_64287 = _T_64286[10:0]; // @[Modules.scala 68:83:@13750.4]
  assign buffer_5_620 = $signed(_T_64287); // @[Modules.scala 68:83:@13751.4]
  assign _T_64289 = $signed(buffer_5_458) + $signed(buffer_5_459); // @[Modules.scala 68:83:@13753.4]
  assign _T_64290 = _T_64289[10:0]; // @[Modules.scala 68:83:@13754.4]
  assign buffer_5_621 = $signed(_T_64290); // @[Modules.scala 68:83:@13755.4]
  assign _T_64292 = $signed(buffer_5_460) + $signed(buffer_5_461); // @[Modules.scala 68:83:@13757.4]
  assign _T_64293 = _T_64292[10:0]; // @[Modules.scala 68:83:@13758.4]
  assign buffer_5_622 = $signed(_T_64293); // @[Modules.scala 68:83:@13759.4]
  assign _T_64295 = $signed(buffer_5_462) + $signed(buffer_5_463); // @[Modules.scala 68:83:@13761.4]
  assign _T_64296 = _T_64295[10:0]; // @[Modules.scala 68:83:@13762.4]
  assign buffer_5_623 = $signed(_T_64296); // @[Modules.scala 68:83:@13763.4]
  assign _T_64298 = $signed(buffer_0_395) + $signed(buffer_5_465); // @[Modules.scala 68:83:@13765.4]
  assign _T_64299 = _T_64298[10:0]; // @[Modules.scala 68:83:@13766.4]
  assign buffer_5_624 = $signed(_T_64299); // @[Modules.scala 68:83:@13767.4]
  assign _T_64301 = $signed(buffer_5_466) + $signed(buffer_5_467); // @[Modules.scala 68:83:@13769.4]
  assign _T_64302 = _T_64301[10:0]; // @[Modules.scala 68:83:@13770.4]
  assign buffer_5_625 = $signed(_T_64302); // @[Modules.scala 68:83:@13771.4]
  assign _T_64304 = $signed(buffer_5_468) + $signed(buffer_5_469); // @[Modules.scala 68:83:@13773.4]
  assign _T_64305 = _T_64304[10:0]; // @[Modules.scala 68:83:@13774.4]
  assign buffer_5_626 = $signed(_T_64305); // @[Modules.scala 68:83:@13775.4]
  assign _T_64310 = $signed(buffer_5_472) + $signed(buffer_5_473); // @[Modules.scala 68:83:@13781.4]
  assign _T_64311 = _T_64310[10:0]; // @[Modules.scala 68:83:@13782.4]
  assign buffer_5_628 = $signed(_T_64311); // @[Modules.scala 68:83:@13783.4]
  assign _T_64313 = $signed(buffer_5_474) + $signed(buffer_3_475); // @[Modules.scala 68:83:@13785.4]
  assign _T_64314 = _T_64313[10:0]; // @[Modules.scala 68:83:@13786.4]
  assign buffer_5_629 = $signed(_T_64314); // @[Modules.scala 68:83:@13787.4]
  assign _T_64316 = $signed(buffer_5_476) + $signed(buffer_5_477); // @[Modules.scala 68:83:@13789.4]
  assign _T_64317 = _T_64316[10:0]; // @[Modules.scala 68:83:@13790.4]
  assign buffer_5_630 = $signed(_T_64317); // @[Modules.scala 68:83:@13791.4]
  assign _T_64319 = $signed(buffer_0_395) + $signed(buffer_5_479); // @[Modules.scala 68:83:@13793.4]
  assign _T_64320 = _T_64319[10:0]; // @[Modules.scala 68:83:@13794.4]
  assign buffer_5_631 = $signed(_T_64320); // @[Modules.scala 68:83:@13795.4]
  assign _T_64322 = $signed(buffer_5_480) + $signed(buffer_5_481); // @[Modules.scala 68:83:@13797.4]
  assign _T_64323 = _T_64322[10:0]; // @[Modules.scala 68:83:@13798.4]
  assign buffer_5_632 = $signed(_T_64323); // @[Modules.scala 68:83:@13799.4]
  assign _T_64325 = $signed(buffer_2_482) + $signed(buffer_5_483); // @[Modules.scala 68:83:@13801.4]
  assign _T_64326 = _T_64325[10:0]; // @[Modules.scala 68:83:@13802.4]
  assign buffer_5_633 = $signed(_T_64326); // @[Modules.scala 68:83:@13803.4]
  assign _T_64328 = $signed(buffer_0_395) + $signed(buffer_5_485); // @[Modules.scala 68:83:@13805.4]
  assign _T_64329 = _T_64328[10:0]; // @[Modules.scala 68:83:@13806.4]
  assign buffer_5_634 = $signed(_T_64329); // @[Modules.scala 68:83:@13807.4]
  assign _T_64331 = $signed(buffer_5_486) + $signed(buffer_0_487); // @[Modules.scala 68:83:@13809.4]
  assign _T_64332 = _T_64331[10:0]; // @[Modules.scala 68:83:@13810.4]
  assign buffer_5_635 = $signed(_T_64332); // @[Modules.scala 68:83:@13811.4]
  assign _T_64334 = $signed(buffer_0_395) + $signed(buffer_5_489); // @[Modules.scala 68:83:@13813.4]
  assign _T_64335 = _T_64334[10:0]; // @[Modules.scala 68:83:@13814.4]
  assign buffer_5_636 = $signed(_T_64335); // @[Modules.scala 68:83:@13815.4]
  assign _T_64337 = $signed(buffer_5_490) + $signed(buffer_0_395); // @[Modules.scala 68:83:@13817.4]
  assign _T_64338 = _T_64337[10:0]; // @[Modules.scala 68:83:@13818.4]
  assign buffer_5_637 = $signed(_T_64338); // @[Modules.scala 68:83:@13819.4]
  assign _T_64340 = $signed(buffer_0_395) + $signed(buffer_0_493); // @[Modules.scala 68:83:@13821.4]
  assign _T_64341 = _T_64340[10:0]; // @[Modules.scala 68:83:@13822.4]
  assign buffer_5_638 = $signed(_T_64341); // @[Modules.scala 68:83:@13823.4]
  assign _T_64343 = $signed(buffer_4_494) + $signed(buffer_0_395); // @[Modules.scala 68:83:@13825.4]
  assign _T_64344 = _T_64343[10:0]; // @[Modules.scala 68:83:@13826.4]
  assign buffer_5_639 = $signed(_T_64344); // @[Modules.scala 68:83:@13827.4]
  assign _T_64346 = $signed(buffer_5_496) + $signed(buffer_5_497); // @[Modules.scala 68:83:@13829.4]
  assign _T_64347 = _T_64346[10:0]; // @[Modules.scala 68:83:@13830.4]
  assign buffer_5_640 = $signed(_T_64347); // @[Modules.scala 68:83:@13831.4]
  assign _T_64349 = $signed(buffer_5_498) + $signed(buffer_0_395); // @[Modules.scala 68:83:@13833.4]
  assign _T_64350 = _T_64349[10:0]; // @[Modules.scala 68:83:@13834.4]
  assign buffer_5_641 = $signed(_T_64350); // @[Modules.scala 68:83:@13835.4]
  assign _T_64352 = $signed(buffer_0_500) + $signed(buffer_5_501); // @[Modules.scala 68:83:@13837.4]
  assign _T_64353 = _T_64352[10:0]; // @[Modules.scala 68:83:@13838.4]
  assign buffer_5_642 = $signed(_T_64353); // @[Modules.scala 68:83:@13839.4]
  assign _T_64355 = $signed(buffer_0_395) + $signed(buffer_5_503); // @[Modules.scala 68:83:@13841.4]
  assign _T_64356 = _T_64355[10:0]; // @[Modules.scala 68:83:@13842.4]
  assign buffer_5_643 = $signed(_T_64356); // @[Modules.scala 68:83:@13843.4]
  assign _T_64358 = $signed(buffer_3_504) + $signed(buffer_5_505); // @[Modules.scala 68:83:@13845.4]
  assign _T_64359 = _T_64358[10:0]; // @[Modules.scala 68:83:@13846.4]
  assign buffer_5_644 = $signed(_T_64359); // @[Modules.scala 68:83:@13847.4]
  assign _T_64361 = $signed(buffer_1_506) + $signed(buffer_5_507); // @[Modules.scala 68:83:@13849.4]
  assign _T_64362 = _T_64361[10:0]; // @[Modules.scala 68:83:@13850.4]
  assign buffer_5_645 = $signed(_T_64362); // @[Modules.scala 68:83:@13851.4]
  assign _T_64364 = $signed(buffer_5_508) + $signed(buffer_0_395); // @[Modules.scala 68:83:@13853.4]
  assign _T_64365 = _T_64364[10:0]; // @[Modules.scala 68:83:@13854.4]
  assign buffer_5_646 = $signed(_T_64365); // @[Modules.scala 68:83:@13855.4]
  assign _T_64367 = $signed(buffer_5_510) + $signed(buffer_3_511); // @[Modules.scala 68:83:@13857.4]
  assign _T_64368 = _T_64367[10:0]; // @[Modules.scala 68:83:@13858.4]
  assign buffer_5_647 = $signed(_T_64368); // @[Modules.scala 68:83:@13859.4]
  assign _T_64370 = $signed(buffer_5_512) + $signed(buffer_5_513); // @[Modules.scala 68:83:@13861.4]
  assign _T_64371 = _T_64370[10:0]; // @[Modules.scala 68:83:@13862.4]
  assign buffer_5_648 = $signed(_T_64371); // @[Modules.scala 68:83:@13863.4]
  assign _T_64373 = $signed(buffer_2_514) + $signed(buffer_5_515); // @[Modules.scala 68:83:@13865.4]
  assign _T_64374 = _T_64373[10:0]; // @[Modules.scala 68:83:@13866.4]
  assign buffer_5_649 = $signed(_T_64374); // @[Modules.scala 68:83:@13867.4]
  assign _T_64376 = $signed(buffer_0_395) + $signed(buffer_3_517); // @[Modules.scala 68:83:@13869.4]
  assign _T_64377 = _T_64376[10:0]; // @[Modules.scala 68:83:@13870.4]
  assign buffer_5_650 = $signed(_T_64377); // @[Modules.scala 68:83:@13871.4]
  assign _T_64379 = $signed(buffer_3_518) + $signed(buffer_5_519); // @[Modules.scala 68:83:@13873.4]
  assign _T_64380 = _T_64379[10:0]; // @[Modules.scala 68:83:@13874.4]
  assign buffer_5_651 = $signed(_T_64380); // @[Modules.scala 68:83:@13875.4]
  assign _T_64382 = $signed(buffer_5_520) + $signed(buffer_5_521); // @[Modules.scala 68:83:@13877.4]
  assign _T_64383 = _T_64382[10:0]; // @[Modules.scala 68:83:@13878.4]
  assign buffer_5_652 = $signed(_T_64383); // @[Modules.scala 68:83:@13879.4]
  assign _T_64385 = $signed(buffer_5_522) + $signed(buffer_1_523); // @[Modules.scala 68:83:@13881.4]
  assign _T_64386 = _T_64385[10:0]; // @[Modules.scala 68:83:@13882.4]
  assign buffer_5_653 = $signed(_T_64386); // @[Modules.scala 68:83:@13883.4]
  assign _T_64388 = $signed(buffer_3_524) + $signed(buffer_4_525); // @[Modules.scala 68:83:@13885.4]
  assign _T_64389 = _T_64388[10:0]; // @[Modules.scala 68:83:@13886.4]
  assign buffer_5_654 = $signed(_T_64389); // @[Modules.scala 68:83:@13887.4]
  assign _T_64391 = $signed(buffer_5_526) + $signed(buffer_5_527); // @[Modules.scala 68:83:@13889.4]
  assign _T_64392 = _T_64391[10:0]; // @[Modules.scala 68:83:@13890.4]
  assign buffer_5_655 = $signed(_T_64392); // @[Modules.scala 68:83:@13891.4]
  assign _T_64394 = $signed(buffer_5_528) + $signed(buffer_5_529); // @[Modules.scala 68:83:@13893.4]
  assign _T_64395 = _T_64394[10:0]; // @[Modules.scala 68:83:@13894.4]
  assign buffer_5_656 = $signed(_T_64395); // @[Modules.scala 68:83:@13895.4]
  assign _T_64397 = $signed(buffer_5_530) + $signed(buffer_5_531); // @[Modules.scala 68:83:@13897.4]
  assign _T_64398 = _T_64397[10:0]; // @[Modules.scala 68:83:@13898.4]
  assign buffer_5_657 = $signed(_T_64398); // @[Modules.scala 68:83:@13899.4]
  assign _T_64400 = $signed(buffer_5_532) + $signed(buffer_5_533); // @[Modules.scala 68:83:@13901.4]
  assign _T_64401 = _T_64400[10:0]; // @[Modules.scala 68:83:@13902.4]
  assign buffer_5_658 = $signed(_T_64401); // @[Modules.scala 68:83:@13903.4]
  assign _T_64406 = $signed(buffer_5_536) + $signed(buffer_5_537); // @[Modules.scala 68:83:@13909.4]
  assign _T_64407 = _T_64406[10:0]; // @[Modules.scala 68:83:@13910.4]
  assign buffer_5_660 = $signed(_T_64407); // @[Modules.scala 68:83:@13911.4]
  assign _T_64409 = $signed(buffer_3_538) + $signed(buffer_4_539); // @[Modules.scala 68:83:@13913.4]
  assign _T_64410 = _T_64409[10:0]; // @[Modules.scala 68:83:@13914.4]
  assign buffer_5_661 = $signed(_T_64410); // @[Modules.scala 68:83:@13915.4]
  assign _T_64412 = $signed(buffer_1_540) + $signed(buffer_5_541); // @[Modules.scala 68:83:@13917.4]
  assign _T_64413 = _T_64412[10:0]; // @[Modules.scala 68:83:@13918.4]
  assign buffer_5_662 = $signed(_T_64413); // @[Modules.scala 68:83:@13919.4]
  assign _T_64415 = $signed(buffer_0_395) + $signed(buffer_5_543); // @[Modules.scala 68:83:@13921.4]
  assign _T_64416 = _T_64415[10:0]; // @[Modules.scala 68:83:@13922.4]
  assign buffer_5_663 = $signed(_T_64416); // @[Modules.scala 68:83:@13923.4]
  assign _T_64418 = $signed(buffer_2_544) + $signed(buffer_0_545); // @[Modules.scala 68:83:@13925.4]
  assign _T_64419 = _T_64418[10:0]; // @[Modules.scala 68:83:@13926.4]
  assign buffer_5_664 = $signed(_T_64419); // @[Modules.scala 68:83:@13927.4]
  assign _T_64421 = $signed(buffer_1_546) + $signed(buffer_4_547); // @[Modules.scala 68:83:@13929.4]
  assign _T_64422 = _T_64421[10:0]; // @[Modules.scala 68:83:@13930.4]
  assign buffer_5_665 = $signed(_T_64422); // @[Modules.scala 68:83:@13931.4]
  assign _T_64424 = $signed(buffer_5_548) + $signed(buffer_5_549); // @[Modules.scala 68:83:@13933.4]
  assign _T_64425 = _T_64424[10:0]; // @[Modules.scala 68:83:@13934.4]
  assign buffer_5_666 = $signed(_T_64425); // @[Modules.scala 68:83:@13935.4]
  assign _T_64427 = $signed(buffer_5_550) + $signed(buffer_0_551); // @[Modules.scala 68:83:@13937.4]
  assign _T_64428 = _T_64427[10:0]; // @[Modules.scala 68:83:@13938.4]
  assign buffer_5_667 = $signed(_T_64428); // @[Modules.scala 68:83:@13939.4]
  assign _T_64430 = $signed(buffer_5_552) + $signed(buffer_1_553); // @[Modules.scala 68:83:@13941.4]
  assign _T_64431 = _T_64430[10:0]; // @[Modules.scala 68:83:@13942.4]
  assign buffer_5_668 = $signed(_T_64431); // @[Modules.scala 68:83:@13943.4]
  assign _T_64433 = $signed(buffer_5_554) + $signed(buffer_5_555); // @[Modules.scala 68:83:@13945.4]
  assign _T_64434 = _T_64433[10:0]; // @[Modules.scala 68:83:@13946.4]
  assign buffer_5_669 = $signed(_T_64434); // @[Modules.scala 68:83:@13947.4]
  assign _T_64436 = $signed(buffer_5_556) + $signed(buffer_5_557); // @[Modules.scala 68:83:@13949.4]
  assign _T_64437 = _T_64436[10:0]; // @[Modules.scala 68:83:@13950.4]
  assign buffer_5_670 = $signed(_T_64437); // @[Modules.scala 68:83:@13951.4]
  assign _T_64439 = $signed(buffer_5_558) + $signed(buffer_0_559); // @[Modules.scala 68:83:@13953.4]
  assign _T_64440 = _T_64439[10:0]; // @[Modules.scala 68:83:@13954.4]
  assign buffer_5_671 = $signed(_T_64440); // @[Modules.scala 68:83:@13955.4]
  assign _T_64442 = $signed(buffer_5_560) + $signed(buffer_5_561); // @[Modules.scala 68:83:@13957.4]
  assign _T_64443 = _T_64442[10:0]; // @[Modules.scala 68:83:@13958.4]
  assign buffer_5_672 = $signed(_T_64443); // @[Modules.scala 68:83:@13959.4]
  assign _T_64445 = $signed(buffer_5_562) + $signed(buffer_5_563); // @[Modules.scala 68:83:@13961.4]
  assign _T_64446 = _T_64445[10:0]; // @[Modules.scala 68:83:@13962.4]
  assign buffer_5_673 = $signed(_T_64446); // @[Modules.scala 68:83:@13963.4]
  assign _T_64451 = $signed(buffer_5_566) + $signed(buffer_5_567); // @[Modules.scala 68:83:@13969.4]
  assign _T_64452 = _T_64451[10:0]; // @[Modules.scala 68:83:@13970.4]
  assign buffer_5_675 = $signed(_T_64452); // @[Modules.scala 68:83:@13971.4]
  assign _T_64454 = $signed(buffer_5_568) + $signed(buffer_3_569); // @[Modules.scala 68:83:@13973.4]
  assign _T_64455 = _T_64454[10:0]; // @[Modules.scala 68:83:@13974.4]
  assign buffer_5_676 = $signed(_T_64455); // @[Modules.scala 68:83:@13975.4]
  assign _T_64460 = $signed(buffer_5_572) + $signed(buffer_0_573); // @[Modules.scala 68:83:@13981.4]
  assign _T_64461 = _T_64460[10:0]; // @[Modules.scala 68:83:@13982.4]
  assign buffer_5_678 = $signed(_T_64461); // @[Modules.scala 68:83:@13983.4]
  assign _T_64463 = $signed(buffer_2_574) + $signed(buffer_5_575); // @[Modules.scala 68:83:@13985.4]
  assign _T_64464 = _T_64463[10:0]; // @[Modules.scala 68:83:@13986.4]
  assign buffer_5_679 = $signed(_T_64464); // @[Modules.scala 68:83:@13987.4]
  assign _T_64466 = $signed(buffer_3_576) + $signed(buffer_5_577); // @[Modules.scala 68:83:@13989.4]
  assign _T_64467 = _T_64466[10:0]; // @[Modules.scala 68:83:@13990.4]
  assign buffer_5_680 = $signed(_T_64467); // @[Modules.scala 68:83:@13991.4]
  assign _T_64469 = $signed(buffer_3_578) + $signed(buffer_5_579); // @[Modules.scala 68:83:@13993.4]
  assign _T_64470 = _T_64469[10:0]; // @[Modules.scala 68:83:@13994.4]
  assign buffer_5_681 = $signed(_T_64470); // @[Modules.scala 68:83:@13995.4]
  assign _T_64472 = $signed(buffer_3_580) + $signed(buffer_1_581); // @[Modules.scala 68:83:@13997.4]
  assign _T_64473 = _T_64472[10:0]; // @[Modules.scala 68:83:@13998.4]
  assign buffer_5_682 = $signed(_T_64473); // @[Modules.scala 68:83:@13999.4]
  assign _T_64475 = $signed(buffer_0_395) + $signed(buffer_5_583); // @[Modules.scala 68:83:@14001.4]
  assign _T_64476 = _T_64475[10:0]; // @[Modules.scala 68:83:@14002.4]
  assign buffer_5_683 = $signed(_T_64476); // @[Modules.scala 68:83:@14003.4]
  assign _T_64481 = $signed(buffer_5_586) + $signed(buffer_3_587); // @[Modules.scala 68:83:@14009.4]
  assign _T_64482 = _T_64481[10:0]; // @[Modules.scala 68:83:@14010.4]
  assign buffer_5_685 = $signed(_T_64482); // @[Modules.scala 68:83:@14011.4]
  assign _T_64484 = $signed(buffer_5_588) + $signed(buffer_5_589); // @[Modules.scala 71:109:@14013.4]
  assign _T_64485 = _T_64484[10:0]; // @[Modules.scala 71:109:@14014.4]
  assign buffer_5_686 = $signed(_T_64485); // @[Modules.scala 71:109:@14015.4]
  assign _T_64487 = $signed(buffer_5_590) + $signed(buffer_5_591); // @[Modules.scala 71:109:@14017.4]
  assign _T_64488 = _T_64487[10:0]; // @[Modules.scala 71:109:@14018.4]
  assign buffer_5_687 = $signed(_T_64488); // @[Modules.scala 71:109:@14019.4]
  assign _T_64490 = $signed(buffer_5_592) + $signed(buffer_5_593); // @[Modules.scala 71:109:@14021.4]
  assign _T_64491 = _T_64490[10:0]; // @[Modules.scala 71:109:@14022.4]
  assign buffer_5_688 = $signed(_T_64491); // @[Modules.scala 71:109:@14023.4]
  assign _T_64493 = $signed(buffer_5_594) + $signed(buffer_5_595); // @[Modules.scala 71:109:@14025.4]
  assign _T_64494 = _T_64493[10:0]; // @[Modules.scala 71:109:@14026.4]
  assign buffer_5_689 = $signed(_T_64494); // @[Modules.scala 71:109:@14027.4]
  assign _T_64496 = $signed(buffer_5_596) + $signed(buffer_5_597); // @[Modules.scala 71:109:@14029.4]
  assign _T_64497 = _T_64496[10:0]; // @[Modules.scala 71:109:@14030.4]
  assign buffer_5_690 = $signed(_T_64497); // @[Modules.scala 71:109:@14031.4]
  assign _T_64499 = $signed(buffer_5_598) + $signed(buffer_0_599); // @[Modules.scala 71:109:@14033.4]
  assign _T_64500 = _T_64499[10:0]; // @[Modules.scala 71:109:@14034.4]
  assign buffer_5_691 = $signed(_T_64500); // @[Modules.scala 71:109:@14035.4]
  assign _T_64502 = $signed(buffer_5_600) + $signed(buffer_5_601); // @[Modules.scala 71:109:@14037.4]
  assign _T_64503 = _T_64502[10:0]; // @[Modules.scala 71:109:@14038.4]
  assign buffer_5_692 = $signed(_T_64503); // @[Modules.scala 71:109:@14039.4]
  assign _T_64505 = $signed(buffer_5_602) + $signed(buffer_3_603); // @[Modules.scala 71:109:@14041.4]
  assign _T_64506 = _T_64505[10:0]; // @[Modules.scala 71:109:@14042.4]
  assign buffer_5_693 = $signed(_T_64506); // @[Modules.scala 71:109:@14043.4]
  assign _T_64508 = $signed(buffer_5_604) + $signed(buffer_5_605); // @[Modules.scala 71:109:@14045.4]
  assign _T_64509 = _T_64508[10:0]; // @[Modules.scala 71:109:@14046.4]
  assign buffer_5_694 = $signed(_T_64509); // @[Modules.scala 71:109:@14047.4]
  assign _T_64511 = $signed(buffer_5_606) + $signed(buffer_5_607); // @[Modules.scala 71:109:@14049.4]
  assign _T_64512 = _T_64511[10:0]; // @[Modules.scala 71:109:@14050.4]
  assign buffer_5_695 = $signed(_T_64512); // @[Modules.scala 71:109:@14051.4]
  assign _T_64514 = $signed(buffer_5_608) + $signed(buffer_5_609); // @[Modules.scala 71:109:@14053.4]
  assign _T_64515 = _T_64514[10:0]; // @[Modules.scala 71:109:@14054.4]
  assign buffer_5_696 = $signed(_T_64515); // @[Modules.scala 71:109:@14055.4]
  assign _T_64517 = $signed(buffer_5_610) + $signed(buffer_5_611); // @[Modules.scala 71:109:@14057.4]
  assign _T_64518 = _T_64517[10:0]; // @[Modules.scala 71:109:@14058.4]
  assign buffer_5_697 = $signed(_T_64518); // @[Modules.scala 71:109:@14059.4]
  assign _T_64520 = $signed(buffer_5_612) + $signed(buffer_5_613); // @[Modules.scala 71:109:@14061.4]
  assign _T_64521 = _T_64520[10:0]; // @[Modules.scala 71:109:@14062.4]
  assign buffer_5_698 = $signed(_T_64521); // @[Modules.scala 71:109:@14063.4]
  assign _T_64523 = $signed(buffer_5_614) + $signed(buffer_5_615); // @[Modules.scala 71:109:@14065.4]
  assign _T_64524 = _T_64523[10:0]; // @[Modules.scala 71:109:@14066.4]
  assign buffer_5_699 = $signed(_T_64524); // @[Modules.scala 71:109:@14067.4]
  assign _T_64526 = $signed(buffer_5_616) + $signed(buffer_5_617); // @[Modules.scala 71:109:@14069.4]
  assign _T_64527 = _T_64526[10:0]; // @[Modules.scala 71:109:@14070.4]
  assign buffer_5_700 = $signed(_T_64527); // @[Modules.scala 71:109:@14071.4]
  assign _T_64529 = $signed(buffer_5_618) + $signed(buffer_5_619); // @[Modules.scala 71:109:@14073.4]
  assign _T_64530 = _T_64529[10:0]; // @[Modules.scala 71:109:@14074.4]
  assign buffer_5_701 = $signed(_T_64530); // @[Modules.scala 71:109:@14075.4]
  assign _T_64532 = $signed(buffer_5_620) + $signed(buffer_5_621); // @[Modules.scala 71:109:@14077.4]
  assign _T_64533 = _T_64532[10:0]; // @[Modules.scala 71:109:@14078.4]
  assign buffer_5_702 = $signed(_T_64533); // @[Modules.scala 71:109:@14079.4]
  assign _T_64535 = $signed(buffer_5_622) + $signed(buffer_5_623); // @[Modules.scala 71:109:@14081.4]
  assign _T_64536 = _T_64535[10:0]; // @[Modules.scala 71:109:@14082.4]
  assign buffer_5_703 = $signed(_T_64536); // @[Modules.scala 71:109:@14083.4]
  assign _T_64538 = $signed(buffer_5_624) + $signed(buffer_5_625); // @[Modules.scala 71:109:@14085.4]
  assign _T_64539 = _T_64538[10:0]; // @[Modules.scala 71:109:@14086.4]
  assign buffer_5_704 = $signed(_T_64539); // @[Modules.scala 71:109:@14087.4]
  assign _T_64541 = $signed(buffer_5_626) + $signed(buffer_0_593); // @[Modules.scala 71:109:@14089.4]
  assign _T_64542 = _T_64541[10:0]; // @[Modules.scala 71:109:@14090.4]
  assign buffer_5_705 = $signed(_T_64542); // @[Modules.scala 71:109:@14091.4]
  assign _T_64544 = $signed(buffer_5_628) + $signed(buffer_5_629); // @[Modules.scala 71:109:@14093.4]
  assign _T_64545 = _T_64544[10:0]; // @[Modules.scala 71:109:@14094.4]
  assign buffer_5_706 = $signed(_T_64545); // @[Modules.scala 71:109:@14095.4]
  assign _T_64547 = $signed(buffer_5_630) + $signed(buffer_5_631); // @[Modules.scala 71:109:@14097.4]
  assign _T_64548 = _T_64547[10:0]; // @[Modules.scala 71:109:@14098.4]
  assign buffer_5_707 = $signed(_T_64548); // @[Modules.scala 71:109:@14099.4]
  assign _T_64550 = $signed(buffer_5_632) + $signed(buffer_5_633); // @[Modules.scala 71:109:@14101.4]
  assign _T_64551 = _T_64550[10:0]; // @[Modules.scala 71:109:@14102.4]
  assign buffer_5_708 = $signed(_T_64551); // @[Modules.scala 71:109:@14103.4]
  assign _T_64553 = $signed(buffer_5_634) + $signed(buffer_5_635); // @[Modules.scala 71:109:@14105.4]
  assign _T_64554 = _T_64553[10:0]; // @[Modules.scala 71:109:@14106.4]
  assign buffer_5_709 = $signed(_T_64554); // @[Modules.scala 71:109:@14107.4]
  assign _T_64556 = $signed(buffer_5_636) + $signed(buffer_5_637); // @[Modules.scala 71:109:@14109.4]
  assign _T_64557 = _T_64556[10:0]; // @[Modules.scala 71:109:@14110.4]
  assign buffer_5_710 = $signed(_T_64557); // @[Modules.scala 71:109:@14111.4]
  assign _T_64559 = $signed(buffer_5_638) + $signed(buffer_5_639); // @[Modules.scala 71:109:@14113.4]
  assign _T_64560 = _T_64559[10:0]; // @[Modules.scala 71:109:@14114.4]
  assign buffer_5_711 = $signed(_T_64560); // @[Modules.scala 71:109:@14115.4]
  assign _T_64562 = $signed(buffer_5_640) + $signed(buffer_5_641); // @[Modules.scala 71:109:@14117.4]
  assign _T_64563 = _T_64562[10:0]; // @[Modules.scala 71:109:@14118.4]
  assign buffer_5_712 = $signed(_T_64563); // @[Modules.scala 71:109:@14119.4]
  assign _T_64565 = $signed(buffer_5_642) + $signed(buffer_5_643); // @[Modules.scala 71:109:@14121.4]
  assign _T_64566 = _T_64565[10:0]; // @[Modules.scala 71:109:@14122.4]
  assign buffer_5_713 = $signed(_T_64566); // @[Modules.scala 71:109:@14123.4]
  assign _T_64568 = $signed(buffer_5_644) + $signed(buffer_5_645); // @[Modules.scala 71:109:@14125.4]
  assign _T_64569 = _T_64568[10:0]; // @[Modules.scala 71:109:@14126.4]
  assign buffer_5_714 = $signed(_T_64569); // @[Modules.scala 71:109:@14127.4]
  assign _T_64571 = $signed(buffer_5_646) + $signed(buffer_5_647); // @[Modules.scala 71:109:@14129.4]
  assign _T_64572 = _T_64571[10:0]; // @[Modules.scala 71:109:@14130.4]
  assign buffer_5_715 = $signed(_T_64572); // @[Modules.scala 71:109:@14131.4]
  assign _T_64574 = $signed(buffer_5_648) + $signed(buffer_5_649); // @[Modules.scala 71:109:@14133.4]
  assign _T_64575 = _T_64574[10:0]; // @[Modules.scala 71:109:@14134.4]
  assign buffer_5_716 = $signed(_T_64575); // @[Modules.scala 71:109:@14135.4]
  assign _T_64577 = $signed(buffer_5_650) + $signed(buffer_5_651); // @[Modules.scala 71:109:@14137.4]
  assign _T_64578 = _T_64577[10:0]; // @[Modules.scala 71:109:@14138.4]
  assign buffer_5_717 = $signed(_T_64578); // @[Modules.scala 71:109:@14139.4]
  assign _T_64580 = $signed(buffer_5_652) + $signed(buffer_5_653); // @[Modules.scala 71:109:@14141.4]
  assign _T_64581 = _T_64580[10:0]; // @[Modules.scala 71:109:@14142.4]
  assign buffer_5_718 = $signed(_T_64581); // @[Modules.scala 71:109:@14143.4]
  assign _T_64583 = $signed(buffer_5_654) + $signed(buffer_5_655); // @[Modules.scala 71:109:@14145.4]
  assign _T_64584 = _T_64583[10:0]; // @[Modules.scala 71:109:@14146.4]
  assign buffer_5_719 = $signed(_T_64584); // @[Modules.scala 71:109:@14147.4]
  assign _T_64586 = $signed(buffer_5_656) + $signed(buffer_5_657); // @[Modules.scala 71:109:@14149.4]
  assign _T_64587 = _T_64586[10:0]; // @[Modules.scala 71:109:@14150.4]
  assign buffer_5_720 = $signed(_T_64587); // @[Modules.scala 71:109:@14151.4]
  assign _T_64589 = $signed(buffer_5_658) + $signed(buffer_0_593); // @[Modules.scala 71:109:@14153.4]
  assign _T_64590 = _T_64589[10:0]; // @[Modules.scala 71:109:@14154.4]
  assign buffer_5_721 = $signed(_T_64590); // @[Modules.scala 71:109:@14155.4]
  assign _T_64592 = $signed(buffer_5_660) + $signed(buffer_5_661); // @[Modules.scala 71:109:@14157.4]
  assign _T_64593 = _T_64592[10:0]; // @[Modules.scala 71:109:@14158.4]
  assign buffer_5_722 = $signed(_T_64593); // @[Modules.scala 71:109:@14159.4]
  assign _T_64595 = $signed(buffer_5_662) + $signed(buffer_5_663); // @[Modules.scala 71:109:@14161.4]
  assign _T_64596 = _T_64595[10:0]; // @[Modules.scala 71:109:@14162.4]
  assign buffer_5_723 = $signed(_T_64596); // @[Modules.scala 71:109:@14163.4]
  assign _T_64598 = $signed(buffer_5_664) + $signed(buffer_5_665); // @[Modules.scala 71:109:@14165.4]
  assign _T_64599 = _T_64598[10:0]; // @[Modules.scala 71:109:@14166.4]
  assign buffer_5_724 = $signed(_T_64599); // @[Modules.scala 71:109:@14167.4]
  assign _T_64601 = $signed(buffer_5_666) + $signed(buffer_5_667); // @[Modules.scala 71:109:@14169.4]
  assign _T_64602 = _T_64601[10:0]; // @[Modules.scala 71:109:@14170.4]
  assign buffer_5_725 = $signed(_T_64602); // @[Modules.scala 71:109:@14171.4]
  assign _T_64604 = $signed(buffer_5_668) + $signed(buffer_5_669); // @[Modules.scala 71:109:@14173.4]
  assign _T_64605 = _T_64604[10:0]; // @[Modules.scala 71:109:@14174.4]
  assign buffer_5_726 = $signed(_T_64605); // @[Modules.scala 71:109:@14175.4]
  assign _T_64607 = $signed(buffer_5_670) + $signed(buffer_5_671); // @[Modules.scala 71:109:@14177.4]
  assign _T_64608 = _T_64607[10:0]; // @[Modules.scala 71:109:@14178.4]
  assign buffer_5_727 = $signed(_T_64608); // @[Modules.scala 71:109:@14179.4]
  assign _T_64610 = $signed(buffer_5_672) + $signed(buffer_5_673); // @[Modules.scala 71:109:@14181.4]
  assign _T_64611 = _T_64610[10:0]; // @[Modules.scala 71:109:@14182.4]
  assign buffer_5_728 = $signed(_T_64611); // @[Modules.scala 71:109:@14183.4]
  assign _T_64613 = $signed(buffer_0_674) + $signed(buffer_5_675); // @[Modules.scala 71:109:@14185.4]
  assign _T_64614 = _T_64613[10:0]; // @[Modules.scala 71:109:@14186.4]
  assign buffer_5_729 = $signed(_T_64614); // @[Modules.scala 71:109:@14187.4]
  assign _T_64616 = $signed(buffer_5_676) + $signed(buffer_0_677); // @[Modules.scala 71:109:@14189.4]
  assign _T_64617 = _T_64616[10:0]; // @[Modules.scala 71:109:@14190.4]
  assign buffer_5_730 = $signed(_T_64617); // @[Modules.scala 71:109:@14191.4]
  assign _T_64619 = $signed(buffer_5_678) + $signed(buffer_5_679); // @[Modules.scala 71:109:@14193.4]
  assign _T_64620 = _T_64619[10:0]; // @[Modules.scala 71:109:@14194.4]
  assign buffer_5_731 = $signed(_T_64620); // @[Modules.scala 71:109:@14195.4]
  assign _T_64622 = $signed(buffer_5_680) + $signed(buffer_5_681); // @[Modules.scala 71:109:@14197.4]
  assign _T_64623 = _T_64622[10:0]; // @[Modules.scala 71:109:@14198.4]
  assign buffer_5_732 = $signed(_T_64623); // @[Modules.scala 71:109:@14199.4]
  assign _T_64625 = $signed(buffer_5_682) + $signed(buffer_5_683); // @[Modules.scala 71:109:@14201.4]
  assign _T_64626 = _T_64625[10:0]; // @[Modules.scala 71:109:@14202.4]
  assign buffer_5_733 = $signed(_T_64626); // @[Modules.scala 71:109:@14203.4]
  assign _T_64628 = $signed(buffer_3_684) + $signed(buffer_5_685); // @[Modules.scala 71:109:@14205.4]
  assign _T_64629 = _T_64628[10:0]; // @[Modules.scala 71:109:@14206.4]
  assign buffer_5_734 = $signed(_T_64629); // @[Modules.scala 71:109:@14207.4]
  assign _T_64631 = $signed(buffer_5_686) + $signed(buffer_5_687); // @[Modules.scala 78:156:@14210.4]
  assign _T_64632 = _T_64631[10:0]; // @[Modules.scala 78:156:@14211.4]
  assign buffer_5_736 = $signed(_T_64632); // @[Modules.scala 78:156:@14212.4]
  assign _T_64634 = $signed(buffer_5_736) + $signed(buffer_5_688); // @[Modules.scala 78:156:@14214.4]
  assign _T_64635 = _T_64634[10:0]; // @[Modules.scala 78:156:@14215.4]
  assign buffer_5_737 = $signed(_T_64635); // @[Modules.scala 78:156:@14216.4]
  assign _T_64637 = $signed(buffer_5_737) + $signed(buffer_5_689); // @[Modules.scala 78:156:@14218.4]
  assign _T_64638 = _T_64637[10:0]; // @[Modules.scala 78:156:@14219.4]
  assign buffer_5_738 = $signed(_T_64638); // @[Modules.scala 78:156:@14220.4]
  assign _T_64640 = $signed(buffer_5_738) + $signed(buffer_5_690); // @[Modules.scala 78:156:@14222.4]
  assign _T_64641 = _T_64640[10:0]; // @[Modules.scala 78:156:@14223.4]
  assign buffer_5_739 = $signed(_T_64641); // @[Modules.scala 78:156:@14224.4]
  assign _T_64643 = $signed(buffer_5_739) + $signed(buffer_5_691); // @[Modules.scala 78:156:@14226.4]
  assign _T_64644 = _T_64643[10:0]; // @[Modules.scala 78:156:@14227.4]
  assign buffer_5_740 = $signed(_T_64644); // @[Modules.scala 78:156:@14228.4]
  assign _T_64646 = $signed(buffer_5_740) + $signed(buffer_5_692); // @[Modules.scala 78:156:@14230.4]
  assign _T_64647 = _T_64646[10:0]; // @[Modules.scala 78:156:@14231.4]
  assign buffer_5_741 = $signed(_T_64647); // @[Modules.scala 78:156:@14232.4]
  assign _T_64649 = $signed(buffer_5_741) + $signed(buffer_5_693); // @[Modules.scala 78:156:@14234.4]
  assign _T_64650 = _T_64649[10:0]; // @[Modules.scala 78:156:@14235.4]
  assign buffer_5_742 = $signed(_T_64650); // @[Modules.scala 78:156:@14236.4]
  assign _T_64652 = $signed(buffer_5_742) + $signed(buffer_5_694); // @[Modules.scala 78:156:@14238.4]
  assign _T_64653 = _T_64652[10:0]; // @[Modules.scala 78:156:@14239.4]
  assign buffer_5_743 = $signed(_T_64653); // @[Modules.scala 78:156:@14240.4]
  assign _T_64655 = $signed(buffer_5_743) + $signed(buffer_5_695); // @[Modules.scala 78:156:@14242.4]
  assign _T_64656 = _T_64655[10:0]; // @[Modules.scala 78:156:@14243.4]
  assign buffer_5_744 = $signed(_T_64656); // @[Modules.scala 78:156:@14244.4]
  assign _T_64658 = $signed(buffer_5_744) + $signed(buffer_5_696); // @[Modules.scala 78:156:@14246.4]
  assign _T_64659 = _T_64658[10:0]; // @[Modules.scala 78:156:@14247.4]
  assign buffer_5_745 = $signed(_T_64659); // @[Modules.scala 78:156:@14248.4]
  assign _T_64661 = $signed(buffer_5_745) + $signed(buffer_5_697); // @[Modules.scala 78:156:@14250.4]
  assign _T_64662 = _T_64661[10:0]; // @[Modules.scala 78:156:@14251.4]
  assign buffer_5_746 = $signed(_T_64662); // @[Modules.scala 78:156:@14252.4]
  assign _T_64664 = $signed(buffer_5_746) + $signed(buffer_5_698); // @[Modules.scala 78:156:@14254.4]
  assign _T_64665 = _T_64664[10:0]; // @[Modules.scala 78:156:@14255.4]
  assign buffer_5_747 = $signed(_T_64665); // @[Modules.scala 78:156:@14256.4]
  assign _T_64667 = $signed(buffer_5_747) + $signed(buffer_5_699); // @[Modules.scala 78:156:@14258.4]
  assign _T_64668 = _T_64667[10:0]; // @[Modules.scala 78:156:@14259.4]
  assign buffer_5_748 = $signed(_T_64668); // @[Modules.scala 78:156:@14260.4]
  assign _T_64670 = $signed(buffer_5_748) + $signed(buffer_5_700); // @[Modules.scala 78:156:@14262.4]
  assign _T_64671 = _T_64670[10:0]; // @[Modules.scala 78:156:@14263.4]
  assign buffer_5_749 = $signed(_T_64671); // @[Modules.scala 78:156:@14264.4]
  assign _T_64673 = $signed(buffer_5_749) + $signed(buffer_5_701); // @[Modules.scala 78:156:@14266.4]
  assign _T_64674 = _T_64673[10:0]; // @[Modules.scala 78:156:@14267.4]
  assign buffer_5_750 = $signed(_T_64674); // @[Modules.scala 78:156:@14268.4]
  assign _T_64676 = $signed(buffer_5_750) + $signed(buffer_5_702); // @[Modules.scala 78:156:@14270.4]
  assign _T_64677 = _T_64676[10:0]; // @[Modules.scala 78:156:@14271.4]
  assign buffer_5_751 = $signed(_T_64677); // @[Modules.scala 78:156:@14272.4]
  assign _T_64679 = $signed(buffer_5_751) + $signed(buffer_5_703); // @[Modules.scala 78:156:@14274.4]
  assign _T_64680 = _T_64679[10:0]; // @[Modules.scala 78:156:@14275.4]
  assign buffer_5_752 = $signed(_T_64680); // @[Modules.scala 78:156:@14276.4]
  assign _T_64682 = $signed(buffer_5_752) + $signed(buffer_5_704); // @[Modules.scala 78:156:@14278.4]
  assign _T_64683 = _T_64682[10:0]; // @[Modules.scala 78:156:@14279.4]
  assign buffer_5_753 = $signed(_T_64683); // @[Modules.scala 78:156:@14280.4]
  assign _T_64685 = $signed(buffer_5_753) + $signed(buffer_5_705); // @[Modules.scala 78:156:@14282.4]
  assign _T_64686 = _T_64685[10:0]; // @[Modules.scala 78:156:@14283.4]
  assign buffer_5_754 = $signed(_T_64686); // @[Modules.scala 78:156:@14284.4]
  assign _T_64688 = $signed(buffer_5_754) + $signed(buffer_5_706); // @[Modules.scala 78:156:@14286.4]
  assign _T_64689 = _T_64688[10:0]; // @[Modules.scala 78:156:@14287.4]
  assign buffer_5_755 = $signed(_T_64689); // @[Modules.scala 78:156:@14288.4]
  assign _T_64691 = $signed(buffer_5_755) + $signed(buffer_5_707); // @[Modules.scala 78:156:@14290.4]
  assign _T_64692 = _T_64691[10:0]; // @[Modules.scala 78:156:@14291.4]
  assign buffer_5_756 = $signed(_T_64692); // @[Modules.scala 78:156:@14292.4]
  assign _T_64694 = $signed(buffer_5_756) + $signed(buffer_5_708); // @[Modules.scala 78:156:@14294.4]
  assign _T_64695 = _T_64694[10:0]; // @[Modules.scala 78:156:@14295.4]
  assign buffer_5_757 = $signed(_T_64695); // @[Modules.scala 78:156:@14296.4]
  assign _T_64697 = $signed(buffer_5_757) + $signed(buffer_5_709); // @[Modules.scala 78:156:@14298.4]
  assign _T_64698 = _T_64697[10:0]; // @[Modules.scala 78:156:@14299.4]
  assign buffer_5_758 = $signed(_T_64698); // @[Modules.scala 78:156:@14300.4]
  assign _T_64700 = $signed(buffer_5_758) + $signed(buffer_5_710); // @[Modules.scala 78:156:@14302.4]
  assign _T_64701 = _T_64700[10:0]; // @[Modules.scala 78:156:@14303.4]
  assign buffer_5_759 = $signed(_T_64701); // @[Modules.scala 78:156:@14304.4]
  assign _T_64703 = $signed(buffer_5_759) + $signed(buffer_5_711); // @[Modules.scala 78:156:@14306.4]
  assign _T_64704 = _T_64703[10:0]; // @[Modules.scala 78:156:@14307.4]
  assign buffer_5_760 = $signed(_T_64704); // @[Modules.scala 78:156:@14308.4]
  assign _T_64706 = $signed(buffer_5_760) + $signed(buffer_5_712); // @[Modules.scala 78:156:@14310.4]
  assign _T_64707 = _T_64706[10:0]; // @[Modules.scala 78:156:@14311.4]
  assign buffer_5_761 = $signed(_T_64707); // @[Modules.scala 78:156:@14312.4]
  assign _T_64709 = $signed(buffer_5_761) + $signed(buffer_5_713); // @[Modules.scala 78:156:@14314.4]
  assign _T_64710 = _T_64709[10:0]; // @[Modules.scala 78:156:@14315.4]
  assign buffer_5_762 = $signed(_T_64710); // @[Modules.scala 78:156:@14316.4]
  assign _T_64712 = $signed(buffer_5_762) + $signed(buffer_5_714); // @[Modules.scala 78:156:@14318.4]
  assign _T_64713 = _T_64712[10:0]; // @[Modules.scala 78:156:@14319.4]
  assign buffer_5_763 = $signed(_T_64713); // @[Modules.scala 78:156:@14320.4]
  assign _T_64715 = $signed(buffer_5_763) + $signed(buffer_5_715); // @[Modules.scala 78:156:@14322.4]
  assign _T_64716 = _T_64715[10:0]; // @[Modules.scala 78:156:@14323.4]
  assign buffer_5_764 = $signed(_T_64716); // @[Modules.scala 78:156:@14324.4]
  assign _T_64718 = $signed(buffer_5_764) + $signed(buffer_5_716); // @[Modules.scala 78:156:@14326.4]
  assign _T_64719 = _T_64718[10:0]; // @[Modules.scala 78:156:@14327.4]
  assign buffer_5_765 = $signed(_T_64719); // @[Modules.scala 78:156:@14328.4]
  assign _T_64721 = $signed(buffer_5_765) + $signed(buffer_5_717); // @[Modules.scala 78:156:@14330.4]
  assign _T_64722 = _T_64721[10:0]; // @[Modules.scala 78:156:@14331.4]
  assign buffer_5_766 = $signed(_T_64722); // @[Modules.scala 78:156:@14332.4]
  assign _T_64724 = $signed(buffer_5_766) + $signed(buffer_5_718); // @[Modules.scala 78:156:@14334.4]
  assign _T_64725 = _T_64724[10:0]; // @[Modules.scala 78:156:@14335.4]
  assign buffer_5_767 = $signed(_T_64725); // @[Modules.scala 78:156:@14336.4]
  assign _T_64727 = $signed(buffer_5_767) + $signed(buffer_5_719); // @[Modules.scala 78:156:@14338.4]
  assign _T_64728 = _T_64727[10:0]; // @[Modules.scala 78:156:@14339.4]
  assign buffer_5_768 = $signed(_T_64728); // @[Modules.scala 78:156:@14340.4]
  assign _T_64730 = $signed(buffer_5_768) + $signed(buffer_5_720); // @[Modules.scala 78:156:@14342.4]
  assign _T_64731 = _T_64730[10:0]; // @[Modules.scala 78:156:@14343.4]
  assign buffer_5_769 = $signed(_T_64731); // @[Modules.scala 78:156:@14344.4]
  assign _T_64733 = $signed(buffer_5_769) + $signed(buffer_5_721); // @[Modules.scala 78:156:@14346.4]
  assign _T_64734 = _T_64733[10:0]; // @[Modules.scala 78:156:@14347.4]
  assign buffer_5_770 = $signed(_T_64734); // @[Modules.scala 78:156:@14348.4]
  assign _T_64736 = $signed(buffer_5_770) + $signed(buffer_5_722); // @[Modules.scala 78:156:@14350.4]
  assign _T_64737 = _T_64736[10:0]; // @[Modules.scala 78:156:@14351.4]
  assign buffer_5_771 = $signed(_T_64737); // @[Modules.scala 78:156:@14352.4]
  assign _T_64739 = $signed(buffer_5_771) + $signed(buffer_5_723); // @[Modules.scala 78:156:@14354.4]
  assign _T_64740 = _T_64739[10:0]; // @[Modules.scala 78:156:@14355.4]
  assign buffer_5_772 = $signed(_T_64740); // @[Modules.scala 78:156:@14356.4]
  assign _T_64742 = $signed(buffer_5_772) + $signed(buffer_5_724); // @[Modules.scala 78:156:@14358.4]
  assign _T_64743 = _T_64742[10:0]; // @[Modules.scala 78:156:@14359.4]
  assign buffer_5_773 = $signed(_T_64743); // @[Modules.scala 78:156:@14360.4]
  assign _T_64745 = $signed(buffer_5_773) + $signed(buffer_5_725); // @[Modules.scala 78:156:@14362.4]
  assign _T_64746 = _T_64745[10:0]; // @[Modules.scala 78:156:@14363.4]
  assign buffer_5_774 = $signed(_T_64746); // @[Modules.scala 78:156:@14364.4]
  assign _T_64748 = $signed(buffer_5_774) + $signed(buffer_5_726); // @[Modules.scala 78:156:@14366.4]
  assign _T_64749 = _T_64748[10:0]; // @[Modules.scala 78:156:@14367.4]
  assign buffer_5_775 = $signed(_T_64749); // @[Modules.scala 78:156:@14368.4]
  assign _T_64751 = $signed(buffer_5_775) + $signed(buffer_5_727); // @[Modules.scala 78:156:@14370.4]
  assign _T_64752 = _T_64751[10:0]; // @[Modules.scala 78:156:@14371.4]
  assign buffer_5_776 = $signed(_T_64752); // @[Modules.scala 78:156:@14372.4]
  assign _T_64754 = $signed(buffer_5_776) + $signed(buffer_5_728); // @[Modules.scala 78:156:@14374.4]
  assign _T_64755 = _T_64754[10:0]; // @[Modules.scala 78:156:@14375.4]
  assign buffer_5_777 = $signed(_T_64755); // @[Modules.scala 78:156:@14376.4]
  assign _T_64757 = $signed(buffer_5_777) + $signed(buffer_5_729); // @[Modules.scala 78:156:@14378.4]
  assign _T_64758 = _T_64757[10:0]; // @[Modules.scala 78:156:@14379.4]
  assign buffer_5_778 = $signed(_T_64758); // @[Modules.scala 78:156:@14380.4]
  assign _T_64760 = $signed(buffer_5_778) + $signed(buffer_5_730); // @[Modules.scala 78:156:@14382.4]
  assign _T_64761 = _T_64760[10:0]; // @[Modules.scala 78:156:@14383.4]
  assign buffer_5_779 = $signed(_T_64761); // @[Modules.scala 78:156:@14384.4]
  assign _T_64763 = $signed(buffer_5_779) + $signed(buffer_5_731); // @[Modules.scala 78:156:@14386.4]
  assign _T_64764 = _T_64763[10:0]; // @[Modules.scala 78:156:@14387.4]
  assign buffer_5_780 = $signed(_T_64764); // @[Modules.scala 78:156:@14388.4]
  assign _T_64766 = $signed(buffer_5_780) + $signed(buffer_5_732); // @[Modules.scala 78:156:@14390.4]
  assign _T_64767 = _T_64766[10:0]; // @[Modules.scala 78:156:@14391.4]
  assign buffer_5_781 = $signed(_T_64767); // @[Modules.scala 78:156:@14392.4]
  assign _T_64769 = $signed(buffer_5_781) + $signed(buffer_5_733); // @[Modules.scala 78:156:@14394.4]
  assign _T_64770 = _T_64769[10:0]; // @[Modules.scala 78:156:@14395.4]
  assign buffer_5_782 = $signed(_T_64770); // @[Modules.scala 78:156:@14396.4]
  assign _T_64772 = $signed(buffer_5_782) + $signed(buffer_5_734); // @[Modules.scala 78:156:@14398.4]
  assign _T_64773 = _T_64772[10:0]; // @[Modules.scala 78:156:@14399.4]
  assign buffer_5_783 = $signed(_T_64773); // @[Modules.scala 78:156:@14400.4]
  assign _T_64873 = $signed(io_in_204) + $signed(io_in_205); // @[Modules.scala 37:46:@14544.4]
  assign _T_64874 = _T_64873[4:0]; // @[Modules.scala 37:46:@14545.4]
  assign _T_64875 = $signed(_T_64874); // @[Modules.scala 37:46:@14546.4]
  assign _T_64909 = $signed(io_in_262) + $signed(io_in_263); // @[Modules.scala 37:46:@14603.4]
  assign _T_64910 = _T_64909[4:0]; // @[Modules.scala 37:46:@14604.4]
  assign _T_64911 = $signed(_T_64910); // @[Modules.scala 37:46:@14605.4]
  assign _T_64948 = $signed(io_in_324) + $signed(io_in_325); // @[Modules.scala 37:46:@14664.4]
  assign _T_64949 = _T_64948[4:0]; // @[Modules.scala 37:46:@14665.4]
  assign _T_64950 = $signed(_T_64949); // @[Modules.scala 37:46:@14666.4]
  assign _T_64960 = $signed(io_in_338) + $signed(io_in_339); // @[Modules.scala 37:46:@14680.4]
  assign _T_64961 = _T_64960[4:0]; // @[Modules.scala 37:46:@14681.4]
  assign _T_64962 = $signed(_T_64961); // @[Modules.scala 37:46:@14682.4]
  assign _T_64963 = $signed(io_in_340) + $signed(io_in_341); // @[Modules.scala 37:46:@14684.4]
  assign _T_64964 = _T_64963[4:0]; // @[Modules.scala 37:46:@14685.4]
  assign _T_64965 = $signed(_T_64964); // @[Modules.scala 37:46:@14686.4]
  assign _T_65020 = $signed(io_in_438) + $signed(io_in_439); // @[Modules.scala 37:46:@14784.4]
  assign _T_65021 = _T_65020[4:0]; // @[Modules.scala 37:46:@14785.4]
  assign _T_65022 = $signed(_T_65021); // @[Modules.scala 37:46:@14786.4]
  assign _T_65058 = $signed(io_in_504) + $signed(io_in_505); // @[Modules.scala 37:46:@14844.4]
  assign _T_65059 = _T_65058[4:0]; // @[Modules.scala 37:46:@14845.4]
  assign _T_65060 = $signed(_T_65059); // @[Modules.scala 37:46:@14846.4]
  assign _T_65102 = $signed(io_in_588) + $signed(io_in_589); // @[Modules.scala 37:46:@14892.4]
  assign _T_65103 = _T_65102[4:0]; // @[Modules.scala 37:46:@14893.4]
  assign _T_65104 = $signed(_T_65103); // @[Modules.scala 37:46:@14894.4]
  assign _T_65226 = $signed(buffer_0_2) + $signed(11'sh0); // @[Modules.scala 65:57:@15066.4]
  assign _T_65227 = _T_65226[10:0]; // @[Modules.scala 65:57:@15067.4]
  assign buffer_6_393 = $signed(_T_65227); // @[Modules.scala 65:57:@15068.4]
  assign _T_65229 = $signed(buffer_2_4) + $signed(buffer_3_5); // @[Modules.scala 65:57:@15070.4]
  assign _T_65230 = _T_65229[10:0]; // @[Modules.scala 65:57:@15071.4]
  assign buffer_6_394 = $signed(_T_65230); // @[Modules.scala 65:57:@15072.4]
  assign _T_65262 = $signed(buffer_3_26) + $signed(buffer_0_27); // @[Modules.scala 65:57:@15114.4]
  assign _T_65263 = _T_65262[10:0]; // @[Modules.scala 65:57:@15115.4]
  assign buffer_6_405 = $signed(_T_65263); // @[Modules.scala 65:57:@15116.4]
  assign _T_65265 = $signed(buffer_2_28) + $signed(buffer_3_29); // @[Modules.scala 65:57:@15118.4]
  assign _T_65266 = _T_65265[10:0]; // @[Modules.scala 65:57:@15119.4]
  assign buffer_6_406 = $signed(_T_65266); // @[Modules.scala 65:57:@15120.4]
  assign _T_65286 = $signed(buffer_5_42) + $signed(buffer_3_43); // @[Modules.scala 65:57:@15146.4]
  assign _T_65287 = _T_65286[10:0]; // @[Modules.scala 65:57:@15147.4]
  assign buffer_6_413 = $signed(_T_65287); // @[Modules.scala 65:57:@15148.4]
  assign buffer_6_53 = {{6{io_in_106[4]}},io_in_106}; // @[Modules.scala 32:22:@8.4]
  assign _T_65301 = $signed(11'sh0) + $signed(buffer_6_53); // @[Modules.scala 65:57:@15166.4]
  assign _T_65302 = _T_65301[10:0]; // @[Modules.scala 65:57:@15167.4]
  assign buffer_6_418 = $signed(_T_65302); // @[Modules.scala 65:57:@15168.4]
  assign _T_65304 = $signed(11'sh0) + $signed(buffer_0_55); // @[Modules.scala 65:57:@15170.4]
  assign _T_65305 = _T_65304[10:0]; // @[Modules.scala 65:57:@15171.4]
  assign buffer_6_419 = $signed(_T_65305); // @[Modules.scala 65:57:@15172.4]
  assign buffer_6_73 = {{6{io_in_146[4]}},io_in_146}; // @[Modules.scala 32:22:@8.4]
  assign _T_65331 = $signed(buffer_3_72) + $signed(buffer_6_73); // @[Modules.scala 65:57:@15206.4]
  assign _T_65332 = _T_65331[10:0]; // @[Modules.scala 65:57:@15207.4]
  assign buffer_6_428 = $signed(_T_65332); // @[Modules.scala 65:57:@15208.4]
  assign buffer_6_74 = {{6{io_in_149[4]}},io_in_149}; // @[Modules.scala 32:22:@8.4]
  assign _T_65334 = $signed(buffer_6_74) + $signed(11'sh0); // @[Modules.scala 65:57:@15210.4]
  assign _T_65335 = _T_65334[10:0]; // @[Modules.scala 65:57:@15211.4]
  assign buffer_6_429 = $signed(_T_65335); // @[Modules.scala 65:57:@15212.4]
  assign _T_65346 = $signed(buffer_2_82) + $signed(11'sh0); // @[Modules.scala 65:57:@15226.4]
  assign _T_65347 = _T_65346[10:0]; // @[Modules.scala 65:57:@15227.4]
  assign buffer_6_433 = $signed(_T_65347); // @[Modules.scala 65:57:@15228.4]
  assign buffer_6_86 = {{6{io_in_173[4]}},io_in_173}; // @[Modules.scala 32:22:@8.4]
  assign _T_65352 = $signed(buffer_6_86) + $signed(buffer_1_87); // @[Modules.scala 65:57:@15234.4]
  assign _T_65353 = _T_65352[10:0]; // @[Modules.scala 65:57:@15235.4]
  assign buffer_6_435 = $signed(_T_65353); // @[Modules.scala 65:57:@15236.4]
  assign _T_65355 = $signed(11'sh0) + $signed(buffer_1_89); // @[Modules.scala 65:57:@15238.4]
  assign _T_65356 = _T_65355[10:0]; // @[Modules.scala 65:57:@15239.4]
  assign buffer_6_436 = $signed(_T_65356); // @[Modules.scala 65:57:@15240.4]
  assign buffer_6_94 = {{6{io_in_189[4]}},io_in_189}; // @[Modules.scala 32:22:@8.4]
  assign _T_65364 = $signed(buffer_6_94) + $signed(11'sh0); // @[Modules.scala 65:57:@15250.4]
  assign _T_65365 = _T_65364[10:0]; // @[Modules.scala 65:57:@15251.4]
  assign buffer_6_439 = $signed(_T_65365); // @[Modules.scala 65:57:@15252.4]
  assign buffer_6_97 = {{6{io_in_194[4]}},io_in_194}; // @[Modules.scala 32:22:@8.4]
  assign _T_65367 = $signed(buffer_1_96) + $signed(buffer_6_97); // @[Modules.scala 65:57:@15254.4]
  assign _T_65368 = _T_65367[10:0]; // @[Modules.scala 65:57:@15255.4]
  assign buffer_6_440 = $signed(_T_65368); // @[Modules.scala 65:57:@15256.4]
  assign _T_65370 = $signed(11'sh0) + $signed(buffer_3_99); // @[Modules.scala 65:57:@15258.4]
  assign _T_65371 = _T_65370[10:0]; // @[Modules.scala 65:57:@15259.4]
  assign buffer_6_441 = $signed(_T_65371); // @[Modules.scala 65:57:@15260.4]
  assign _T_65373 = $signed(buffer_3_100) + $signed(buffer_4_101); // @[Modules.scala 65:57:@15262.4]
  assign _T_65374 = _T_65373[10:0]; // @[Modules.scala 65:57:@15263.4]
  assign buffer_6_442 = $signed(_T_65374); // @[Modules.scala 65:57:@15264.4]
  assign buffer_6_102 = {{6{_T_64875[4]}},_T_64875}; // @[Modules.scala 32:22:@8.4]
  assign _T_65376 = $signed(buffer_6_102) + $signed(buffer_3_103); // @[Modules.scala 65:57:@15266.4]
  assign _T_65377 = _T_65376[10:0]; // @[Modules.scala 65:57:@15267.4]
  assign buffer_6_443 = $signed(_T_65377); // @[Modules.scala 65:57:@15268.4]
  assign _T_65379 = $signed(buffer_3_104) + $signed(11'sh0); // @[Modules.scala 65:57:@15270.4]
  assign _T_65380 = _T_65379[10:0]; // @[Modules.scala 65:57:@15271.4]
  assign buffer_6_444 = $signed(_T_65380); // @[Modules.scala 65:57:@15272.4]
  assign buffer_6_107 = {{6{io_in_214[4]}},io_in_214}; // @[Modules.scala 32:22:@8.4]
  assign _T_65382 = $signed(buffer_3_106) + $signed(buffer_6_107); // @[Modules.scala 65:57:@15274.4]
  assign _T_65383 = _T_65382[10:0]; // @[Modules.scala 65:57:@15275.4]
  assign buffer_6_445 = $signed(_T_65383); // @[Modules.scala 65:57:@15276.4]
  assign _T_65385 = $signed(buffer_5_108) + $signed(buffer_3_109); // @[Modules.scala 65:57:@15278.4]
  assign _T_65386 = _T_65385[10:0]; // @[Modules.scala 65:57:@15279.4]
  assign buffer_6_446 = $signed(_T_65386); // @[Modules.scala 65:57:@15280.4]
  assign _T_65391 = $signed(11'sh0) + $signed(buffer_3_113); // @[Modules.scala 65:57:@15286.4]
  assign _T_65392 = _T_65391[10:0]; // @[Modules.scala 65:57:@15287.4]
  assign buffer_6_448 = $signed(_T_65392); // @[Modules.scala 65:57:@15288.4]
  assign _T_65397 = $signed(buffer_3_116) + $signed(buffer_2_117); // @[Modules.scala 65:57:@15294.4]
  assign _T_65398 = _T_65397[10:0]; // @[Modules.scala 65:57:@15295.4]
  assign buffer_6_450 = $signed(_T_65398); // @[Modules.scala 65:57:@15296.4]
  assign buffer_6_120 = {{6{io_in_241[4]}},io_in_241}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_121 = {{6{io_in_242[4]}},io_in_242}; // @[Modules.scala 32:22:@8.4]
  assign _T_65403 = $signed(buffer_6_120) + $signed(buffer_6_121); // @[Modules.scala 65:57:@15302.4]
  assign _T_65404 = _T_65403[10:0]; // @[Modules.scala 65:57:@15303.4]
  assign buffer_6_452 = $signed(_T_65404); // @[Modules.scala 65:57:@15304.4]
  assign buffer_6_123 = {{6{io_in_246[4]}},io_in_246}; // @[Modules.scala 32:22:@8.4]
  assign _T_65406 = $signed(buffer_3_122) + $signed(buffer_6_123); // @[Modules.scala 65:57:@15306.4]
  assign _T_65407 = _T_65406[10:0]; // @[Modules.scala 65:57:@15307.4]
  assign buffer_6_453 = $signed(_T_65407); // @[Modules.scala 65:57:@15308.4]
  assign _T_65412 = $signed(11'sh0) + $signed(buffer_3_127); // @[Modules.scala 65:57:@15314.4]
  assign _T_65413 = _T_65412[10:0]; // @[Modules.scala 65:57:@15315.4]
  assign buffer_6_455 = $signed(_T_65413); // @[Modules.scala 65:57:@15316.4]
  assign buffer_6_129 = {{6{io_in_258[4]}},io_in_258}; // @[Modules.scala 32:22:@8.4]
  assign _T_65415 = $signed(buffer_4_128) + $signed(buffer_6_129); // @[Modules.scala 65:57:@15318.4]
  assign _T_65416 = _T_65415[10:0]; // @[Modules.scala 65:57:@15319.4]
  assign buffer_6_456 = $signed(_T_65416); // @[Modules.scala 65:57:@15320.4]
  assign buffer_6_131 = {{6{_T_64911[4]}},_T_64911}; // @[Modules.scala 32:22:@8.4]
  assign _T_65418 = $signed(buffer_4_130) + $signed(buffer_6_131); // @[Modules.scala 65:57:@15322.4]
  assign _T_65419 = _T_65418[10:0]; // @[Modules.scala 65:57:@15323.4]
  assign buffer_6_457 = $signed(_T_65419); // @[Modules.scala 65:57:@15324.4]
  assign _T_65427 = $signed(buffer_5_136) + $signed(11'sh0); // @[Modules.scala 65:57:@15334.4]
  assign _T_65428 = _T_65427[10:0]; // @[Modules.scala 65:57:@15335.4]
  assign buffer_6_460 = $signed(_T_65428); // @[Modules.scala 65:57:@15336.4]
  assign _T_65433 = $signed(11'sh0) + $signed(buffer_3_141); // @[Modules.scala 65:57:@15342.4]
  assign _T_65434 = _T_65433[10:0]; // @[Modules.scala 65:57:@15343.4]
  assign buffer_6_462 = $signed(_T_65434); // @[Modules.scala 65:57:@15344.4]
  assign buffer_6_145 = {{6{io_in_290[4]}},io_in_290}; // @[Modules.scala 32:22:@8.4]
  assign _T_65439 = $signed(buffer_0_144) + $signed(buffer_6_145); // @[Modules.scala 65:57:@15350.4]
  assign _T_65440 = _T_65439[10:0]; // @[Modules.scala 65:57:@15351.4]
  assign buffer_6_464 = $signed(_T_65440); // @[Modules.scala 65:57:@15352.4]
  assign _T_65442 = $signed(buffer_1_146) + $signed(buffer_3_147); // @[Modules.scala 65:57:@15354.4]
  assign _T_65443 = _T_65442[10:0]; // @[Modules.scala 65:57:@15355.4]
  assign buffer_6_465 = $signed(_T_65443); // @[Modules.scala 65:57:@15356.4]
  assign _T_65445 = $signed(buffer_3_148) + $signed(buffer_4_149); // @[Modules.scala 65:57:@15358.4]
  assign _T_65446 = _T_65445[10:0]; // @[Modules.scala 65:57:@15359.4]
  assign buffer_6_466 = $signed(_T_65446); // @[Modules.scala 65:57:@15360.4]
  assign buffer_6_150 = {{6{io_in_301[4]}},io_in_301}; // @[Modules.scala 32:22:@8.4]
  assign _T_65448 = $signed(buffer_6_150) + $signed(11'sh0); // @[Modules.scala 65:57:@15362.4]
  assign _T_65449 = _T_65448[10:0]; // @[Modules.scala 65:57:@15363.4]
  assign buffer_6_467 = $signed(_T_65449); // @[Modules.scala 65:57:@15364.4]
  assign _T_65454 = $signed(buffer_3_154) + $signed(buffer_4_155); // @[Modules.scala 65:57:@15370.4]
  assign _T_65455 = _T_65454[10:0]; // @[Modules.scala 65:57:@15371.4]
  assign buffer_6_469 = $signed(_T_65455); // @[Modules.scala 65:57:@15372.4]
  assign buffer_6_156 = {{6{io_in_313[4]}},io_in_313}; // @[Modules.scala 32:22:@8.4]
  assign _T_65457 = $signed(buffer_6_156) + $signed(buffer_0_157); // @[Modules.scala 65:57:@15374.4]
  assign _T_65458 = _T_65457[10:0]; // @[Modules.scala 65:57:@15375.4]
  assign buffer_6_470 = $signed(_T_65458); // @[Modules.scala 65:57:@15376.4]
  assign buffer_6_158 = {{6{io_in_317[4]}},io_in_317}; // @[Modules.scala 32:22:@8.4]
  assign _T_65460 = $signed(buffer_6_158) + $signed(buffer_0_159); // @[Modules.scala 65:57:@15378.4]
  assign _T_65461 = _T_65460[10:0]; // @[Modules.scala 65:57:@15379.4]
  assign buffer_6_471 = $signed(_T_65461); // @[Modules.scala 65:57:@15380.4]
  assign buffer_6_161 = {{6{io_in_323[4]}},io_in_323}; // @[Modules.scala 32:22:@8.4]
  assign _T_65463 = $signed(buffer_2_160) + $signed(buffer_6_161); // @[Modules.scala 65:57:@15382.4]
  assign _T_65464 = _T_65463[10:0]; // @[Modules.scala 65:57:@15383.4]
  assign buffer_6_472 = $signed(_T_65464); // @[Modules.scala 65:57:@15384.4]
  assign buffer_6_162 = {{6{_T_64950[4]}},_T_64950}; // @[Modules.scala 32:22:@8.4]
  assign _T_65466 = $signed(buffer_6_162) + $signed(buffer_5_163); // @[Modules.scala 65:57:@15386.4]
  assign _T_65467 = _T_65466[10:0]; // @[Modules.scala 65:57:@15387.4]
  assign buffer_6_473 = $signed(_T_65467); // @[Modules.scala 65:57:@15388.4]
  assign buffer_6_169 = {{6{_T_64962[4]}},_T_64962}; // @[Modules.scala 32:22:@8.4]
  assign _T_65475 = $signed(buffer_3_168) + $signed(buffer_6_169); // @[Modules.scala 65:57:@15398.4]
  assign _T_65476 = _T_65475[10:0]; // @[Modules.scala 65:57:@15399.4]
  assign buffer_6_476 = $signed(_T_65476); // @[Modules.scala 65:57:@15400.4]
  assign buffer_6_170 = {{6{_T_64965[4]}},_T_64965}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_171 = {{6{io_in_343[4]}},io_in_343}; // @[Modules.scala 32:22:@8.4]
  assign _T_65478 = $signed(buffer_6_170) + $signed(buffer_6_171); // @[Modules.scala 65:57:@15402.4]
  assign _T_65479 = _T_65478[10:0]; // @[Modules.scala 65:57:@15403.4]
  assign buffer_6_477 = $signed(_T_65479); // @[Modules.scala 65:57:@15404.4]
  assign buffer_6_173 = {{6{io_in_347[4]}},io_in_347}; // @[Modules.scala 32:22:@8.4]
  assign _T_65481 = $signed(buffer_0_172) + $signed(buffer_6_173); // @[Modules.scala 65:57:@15406.4]
  assign _T_65482 = _T_65481[10:0]; // @[Modules.scala 65:57:@15407.4]
  assign buffer_6_478 = $signed(_T_65482); // @[Modules.scala 65:57:@15408.4]
  assign buffer_6_175 = {{6{io_in_351[4]}},io_in_351}; // @[Modules.scala 32:22:@8.4]
  assign _T_65484 = $signed(11'sh0) + $signed(buffer_6_175); // @[Modules.scala 65:57:@15410.4]
  assign _T_65485 = _T_65484[10:0]; // @[Modules.scala 65:57:@15411.4]
  assign buffer_6_479 = $signed(_T_65485); // @[Modules.scala 65:57:@15412.4]
  assign buffer_6_178 = {{6{io_in_357[4]}},io_in_357}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_179 = {{6{io_in_358[4]}},io_in_358}; // @[Modules.scala 32:22:@8.4]
  assign _T_65490 = $signed(buffer_6_178) + $signed(buffer_6_179); // @[Modules.scala 65:57:@15418.4]
  assign _T_65491 = _T_65490[10:0]; // @[Modules.scala 65:57:@15419.4]
  assign buffer_6_481 = $signed(_T_65491); // @[Modules.scala 65:57:@15420.4]
  assign _T_65496 = $signed(buffer_4_182) + $signed(buffer_5_183); // @[Modules.scala 65:57:@15426.4]
  assign _T_65497 = _T_65496[10:0]; // @[Modules.scala 65:57:@15427.4]
  assign buffer_6_483 = $signed(_T_65497); // @[Modules.scala 65:57:@15428.4]
  assign _T_65502 = $signed(buffer_5_186) + $signed(buffer_0_187); // @[Modules.scala 65:57:@15434.4]
  assign _T_65503 = _T_65502[10:0]; // @[Modules.scala 65:57:@15435.4]
  assign buffer_6_485 = $signed(_T_65503); // @[Modules.scala 65:57:@15436.4]
  assign buffer_6_189 = {{6{io_in_379[4]}},io_in_379}; // @[Modules.scala 32:22:@8.4]
  assign _T_65505 = $signed(11'sh0) + $signed(buffer_6_189); // @[Modules.scala 65:57:@15438.4]
  assign _T_65506 = _T_65505[10:0]; // @[Modules.scala 65:57:@15439.4]
  assign buffer_6_486 = $signed(_T_65506); // @[Modules.scala 65:57:@15440.4]
  assign buffer_6_196 = {{6{io_in_393[4]}},io_in_393}; // @[Modules.scala 32:22:@8.4]
  assign _T_65517 = $signed(buffer_6_196) + $signed(buffer_5_197); // @[Modules.scala 65:57:@15454.4]
  assign _T_65518 = _T_65517[10:0]; // @[Modules.scala 65:57:@15455.4]
  assign buffer_6_490 = $signed(_T_65518); // @[Modules.scala 65:57:@15456.4]
  assign _T_65523 = $signed(buffer_3_200) + $signed(11'sh0); // @[Modules.scala 65:57:@15462.4]
  assign _T_65524 = _T_65523[10:0]; // @[Modules.scala 65:57:@15463.4]
  assign buffer_6_492 = $signed(_T_65524); // @[Modules.scala 65:57:@15464.4]
  assign _T_65526 = $signed(11'sh0) + $signed(buffer_4_203); // @[Modules.scala 65:57:@15466.4]
  assign _T_65527 = _T_65526[10:0]; // @[Modules.scala 65:57:@15467.4]
  assign buffer_6_493 = $signed(_T_65527); // @[Modules.scala 65:57:@15468.4]
  assign buffer_6_207 = {{6{io_in_414[4]}},io_in_414}; // @[Modules.scala 32:22:@8.4]
  assign _T_65532 = $signed(buffer_4_206) + $signed(buffer_6_207); // @[Modules.scala 65:57:@15474.4]
  assign _T_65533 = _T_65532[10:0]; // @[Modules.scala 65:57:@15475.4]
  assign buffer_6_495 = $signed(_T_65533); // @[Modules.scala 65:57:@15476.4]
  assign _T_65535 = $signed(buffer_3_208) + $signed(buffer_0_209); // @[Modules.scala 65:57:@15478.4]
  assign _T_65536 = _T_65535[10:0]; // @[Modules.scala 65:57:@15479.4]
  assign buffer_6_496 = $signed(_T_65536); // @[Modules.scala 65:57:@15480.4]
  assign _T_65538 = $signed(buffer_0_210) + $signed(buffer_5_211); // @[Modules.scala 65:57:@15482.4]
  assign _T_65539 = _T_65538[10:0]; // @[Modules.scala 65:57:@15483.4]
  assign buffer_6_497 = $signed(_T_65539); // @[Modules.scala 65:57:@15484.4]
  assign buffer_6_213 = {{6{io_in_426[4]}},io_in_426}; // @[Modules.scala 32:22:@8.4]
  assign _T_65541 = $signed(buffer_3_212) + $signed(buffer_6_213); // @[Modules.scala 65:57:@15486.4]
  assign _T_65542 = _T_65541[10:0]; // @[Modules.scala 65:57:@15487.4]
  assign buffer_6_498 = $signed(_T_65542); // @[Modules.scala 65:57:@15488.4]
  assign buffer_6_214 = {{6{io_in_428[4]}},io_in_428}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_215 = {{6{io_in_431[4]}},io_in_431}; // @[Modules.scala 32:22:@8.4]
  assign _T_65544 = $signed(buffer_6_214) + $signed(buffer_6_215); // @[Modules.scala 65:57:@15490.4]
  assign _T_65545 = _T_65544[10:0]; // @[Modules.scala 65:57:@15491.4]
  assign buffer_6_499 = $signed(_T_65545); // @[Modules.scala 65:57:@15492.4]
  assign buffer_6_217 = {{6{io_in_435[4]}},io_in_435}; // @[Modules.scala 32:22:@8.4]
  assign _T_65547 = $signed(buffer_4_216) + $signed(buffer_6_217); // @[Modules.scala 65:57:@15494.4]
  assign _T_65548 = _T_65547[10:0]; // @[Modules.scala 65:57:@15495.4]
  assign buffer_6_500 = $signed(_T_65548); // @[Modules.scala 65:57:@15496.4]
  assign buffer_6_219 = {{6{_T_65022[4]}},_T_65022}; // @[Modules.scala 32:22:@8.4]
  assign _T_65550 = $signed(buffer_0_218) + $signed(buffer_6_219); // @[Modules.scala 65:57:@15498.4]
  assign _T_65551 = _T_65550[10:0]; // @[Modules.scala 65:57:@15499.4]
  assign buffer_6_501 = $signed(_T_65551); // @[Modules.scala 65:57:@15500.4]
  assign buffer_6_221 = {{6{io_in_442[4]}},io_in_442}; // @[Modules.scala 32:22:@8.4]
  assign _T_65553 = $signed(buffer_0_220) + $signed(buffer_6_221); // @[Modules.scala 65:57:@15502.4]
  assign _T_65554 = _T_65553[10:0]; // @[Modules.scala 65:57:@15503.4]
  assign buffer_6_502 = $signed(_T_65554); // @[Modules.scala 65:57:@15504.4]
  assign _T_65559 = $signed(buffer_3_224) + $signed(11'sh0); // @[Modules.scala 65:57:@15510.4]
  assign _T_65560 = _T_65559[10:0]; // @[Modules.scala 65:57:@15511.4]
  assign buffer_6_504 = $signed(_T_65560); // @[Modules.scala 65:57:@15512.4]
  assign buffer_6_229 = {{6{io_in_459[4]}},io_in_459}; // @[Modules.scala 32:22:@8.4]
  assign _T_65565 = $signed(buffer_2_228) + $signed(buffer_6_229); // @[Modules.scala 65:57:@15518.4]
  assign _T_65566 = _T_65565[10:0]; // @[Modules.scala 65:57:@15519.4]
  assign buffer_6_506 = $signed(_T_65566); // @[Modules.scala 65:57:@15520.4]
  assign _T_65568 = $signed(11'sh0) + $signed(buffer_0_231); // @[Modules.scala 65:57:@15522.4]
  assign _T_65569 = _T_65568[10:0]; // @[Modules.scala 65:57:@15523.4]
  assign buffer_6_507 = $signed(_T_65569); // @[Modules.scala 65:57:@15524.4]
  assign buffer_6_233 = {{6{io_in_466[4]}},io_in_466}; // @[Modules.scala 32:22:@8.4]
  assign _T_65571 = $signed(buffer_0_232) + $signed(buffer_6_233); // @[Modules.scala 65:57:@15526.4]
  assign _T_65572 = _T_65571[10:0]; // @[Modules.scala 65:57:@15527.4]
  assign buffer_6_508 = $signed(_T_65572); // @[Modules.scala 65:57:@15528.4]
  assign buffer_6_235 = {{6{io_in_470[4]}},io_in_470}; // @[Modules.scala 32:22:@8.4]
  assign _T_65574 = $signed(buffer_0_234) + $signed(buffer_6_235); // @[Modules.scala 65:57:@15530.4]
  assign _T_65575 = _T_65574[10:0]; // @[Modules.scala 65:57:@15531.4]
  assign buffer_6_509 = $signed(_T_65575); // @[Modules.scala 65:57:@15532.4]
  assign _T_65580 = $signed(buffer_1_238) + $signed(buffer_0_239); // @[Modules.scala 65:57:@15538.4]
  assign _T_65581 = _T_65580[10:0]; // @[Modules.scala 65:57:@15539.4]
  assign buffer_6_511 = $signed(_T_65581); // @[Modules.scala 65:57:@15540.4]
  assign buffer_6_241 = {{6{io_in_483[4]}},io_in_483}; // @[Modules.scala 32:22:@8.4]
  assign _T_65583 = $signed(11'sh0) + $signed(buffer_6_241); // @[Modules.scala 65:57:@15542.4]
  assign _T_65584 = _T_65583[10:0]; // @[Modules.scala 65:57:@15543.4]
  assign buffer_6_512 = $signed(_T_65584); // @[Modules.scala 65:57:@15544.4]
  assign _T_65586 = $signed(buffer_5_242) + $signed(buffer_0_243); // @[Modules.scala 65:57:@15546.4]
  assign _T_65587 = _T_65586[10:0]; // @[Modules.scala 65:57:@15547.4]
  assign buffer_6_513 = $signed(_T_65587); // @[Modules.scala 65:57:@15548.4]
  assign _T_65592 = $signed(buffer_4_246) + $signed(buffer_0_247); // @[Modules.scala 65:57:@15554.4]
  assign _T_65593 = _T_65592[10:0]; // @[Modules.scala 65:57:@15555.4]
  assign buffer_6_515 = $signed(_T_65593); // @[Modules.scala 65:57:@15556.4]
  assign buffer_6_252 = {{6{_T_65060[4]}},_T_65060}; // @[Modules.scala 32:22:@8.4]
  assign buffer_6_253 = {{6{io_in_506[4]}},io_in_506}; // @[Modules.scala 32:22:@8.4]
  assign _T_65601 = $signed(buffer_6_252) + $signed(buffer_6_253); // @[Modules.scala 65:57:@15566.4]
  assign _T_65602 = _T_65601[10:0]; // @[Modules.scala 65:57:@15567.4]
  assign buffer_6_518 = $signed(_T_65602); // @[Modules.scala 65:57:@15568.4]
  assign _T_65610 = $signed(11'sh0) + $signed(buffer_0_259); // @[Modules.scala 65:57:@15578.4]
  assign _T_65611 = _T_65610[10:0]; // @[Modules.scala 65:57:@15579.4]
  assign buffer_6_521 = $signed(_T_65611); // @[Modules.scala 65:57:@15580.4]
  assign buffer_6_294 = {{6{_T_65104[4]}},_T_65104}; // @[Modules.scala 32:22:@8.4]
  assign _T_65664 = $signed(buffer_6_294) + $signed(11'sh0); // @[Modules.scala 65:57:@15650.4]
  assign _T_65665 = _T_65664[10:0]; // @[Modules.scala 65:57:@15651.4]
  assign buffer_6_539 = $signed(_T_65665); // @[Modules.scala 65:57:@15652.4]
  assign buffer_6_306 = {{6{io_in_613[4]}},io_in_613}; // @[Modules.scala 32:22:@8.4]
  assign _T_65682 = $signed(buffer_6_306) + $signed(buffer_0_307); // @[Modules.scala 65:57:@15674.4]
  assign _T_65683 = _T_65682[10:0]; // @[Modules.scala 65:57:@15675.4]
  assign buffer_6_545 = $signed(_T_65683); // @[Modules.scala 65:57:@15676.4]
  assign buffer_6_312 = {{6{io_in_625[4]}},io_in_625}; // @[Modules.scala 32:22:@8.4]
  assign _T_65691 = $signed(buffer_6_312) + $signed(11'sh0); // @[Modules.scala 65:57:@15686.4]
  assign _T_65692 = _T_65691[10:0]; // @[Modules.scala 65:57:@15687.4]
  assign buffer_6_548 = $signed(_T_65692); // @[Modules.scala 65:57:@15688.4]
  assign buffer_6_315 = {{6{io_in_631[4]}},io_in_631}; // @[Modules.scala 32:22:@8.4]
  assign _T_65694 = $signed(buffer_5_314) + $signed(buffer_6_315); // @[Modules.scala 65:57:@15690.4]
  assign _T_65695 = _T_65694[10:0]; // @[Modules.scala 65:57:@15691.4]
  assign buffer_6_549 = $signed(_T_65695); // @[Modules.scala 65:57:@15692.4]
  assign _T_65709 = $signed(11'sh0) + $signed(buffer_1_325); // @[Modules.scala 65:57:@15710.4]
  assign _T_65710 = _T_65709[10:0]; // @[Modules.scala 65:57:@15711.4]
  assign buffer_6_554 = $signed(_T_65710); // @[Modules.scala 65:57:@15712.4]
  assign buffer_6_327 = {{6{io_in_654[4]}},io_in_654}; // @[Modules.scala 32:22:@8.4]
  assign _T_65712 = $signed(buffer_5_326) + $signed(buffer_6_327); // @[Modules.scala 65:57:@15714.4]
  assign _T_65713 = _T_65712[10:0]; // @[Modules.scala 65:57:@15715.4]
  assign buffer_6_555 = $signed(_T_65713); // @[Modules.scala 65:57:@15716.4]
  assign _T_65724 = $signed(11'sh0) + $signed(buffer_4_335); // @[Modules.scala 65:57:@15730.4]
  assign _T_65725 = _T_65724[10:0]; // @[Modules.scala 65:57:@15731.4]
  assign buffer_6_559 = $signed(_T_65725); // @[Modules.scala 65:57:@15732.4]
  assign _T_65727 = $signed(buffer_4_336) + $signed(11'sh0); // @[Modules.scala 65:57:@15734.4]
  assign _T_65728 = _T_65727[10:0]; // @[Modules.scala 65:57:@15735.4]
  assign buffer_6_560 = $signed(_T_65728); // @[Modules.scala 65:57:@15736.4]
  assign _T_65739 = $signed(buffer_2_344) + $signed(11'sh0); // @[Modules.scala 65:57:@15750.4]
  assign _T_65740 = _T_65739[10:0]; // @[Modules.scala 65:57:@15751.4]
  assign buffer_6_564 = $signed(_T_65740); // @[Modules.scala 65:57:@15752.4]
  assign _T_65742 = $signed(buffer_0_346) + $signed(buffer_1_347); // @[Modules.scala 65:57:@15754.4]
  assign _T_65743 = _T_65742[10:0]; // @[Modules.scala 65:57:@15755.4]
  assign buffer_6_565 = $signed(_T_65743); // @[Modules.scala 65:57:@15756.4]
  assign _T_65754 = $signed(buffer_0_354) + $signed(buffer_1_355); // @[Modules.scala 65:57:@15770.4]
  assign _T_65755 = _T_65754[10:0]; // @[Modules.scala 65:57:@15771.4]
  assign buffer_6_569 = $signed(_T_65755); // @[Modules.scala 65:57:@15772.4]
  assign buffer_6_357 = {{6{io_in_714[4]}},io_in_714}; // @[Modules.scala 32:22:@8.4]
  assign _T_65757 = $signed(11'sh0) + $signed(buffer_6_357); // @[Modules.scala 65:57:@15774.4]
  assign _T_65758 = _T_65757[10:0]; // @[Modules.scala 65:57:@15775.4]
  assign buffer_6_570 = $signed(_T_65758); // @[Modules.scala 65:57:@15776.4]
  assign buffer_6_359 = {{6{io_in_719[4]}},io_in_719}; // @[Modules.scala 32:22:@8.4]
  assign _T_65760 = $signed(11'sh0) + $signed(buffer_6_359); // @[Modules.scala 65:57:@15778.4]
  assign _T_65761 = _T_65760[10:0]; // @[Modules.scala 65:57:@15779.4]
  assign buffer_6_571 = $signed(_T_65761); // @[Modules.scala 65:57:@15780.4]
  assign _T_65769 = $signed(buffer_0_364) + $signed(buffer_2_365); // @[Modules.scala 65:57:@15790.4]
  assign _T_65770 = _T_65769[10:0]; // @[Modules.scala 65:57:@15791.4]
  assign buffer_6_574 = $signed(_T_65770); // @[Modules.scala 65:57:@15792.4]
  assign _T_65784 = $signed(buffer_0_374) + $signed(11'sh0); // @[Modules.scala 65:57:@15810.4]
  assign _T_65785 = _T_65784[10:0]; // @[Modules.scala 65:57:@15811.4]
  assign buffer_6_579 = $signed(_T_65785); // @[Modules.scala 65:57:@15812.4]
  assign buffer_6_384 = {{6{io_in_769[4]}},io_in_769}; // @[Modules.scala 32:22:@8.4]
  assign _T_65799 = $signed(buffer_6_384) + $signed(buffer_3_385); // @[Modules.scala 65:57:@15830.4]
  assign _T_65800 = _T_65799[10:0]; // @[Modules.scala 65:57:@15831.4]
  assign buffer_6_584 = $signed(_T_65800); // @[Modules.scala 65:57:@15832.4]
  assign buffer_6_388 = {{6{io_in_777[4]}},io_in_777}; // @[Modules.scala 32:22:@8.4]
  assign _T_65805 = $signed(buffer_6_388) + $signed(buffer_5_389); // @[Modules.scala 65:57:@15838.4]
  assign _T_65806 = _T_65805[10:0]; // @[Modules.scala 65:57:@15839.4]
  assign buffer_6_586 = $signed(_T_65806); // @[Modules.scala 65:57:@15840.4]
  assign _T_65811 = $signed(buffer_0_392) + $signed(buffer_6_393); // @[Modules.scala 68:83:@15846.4]
  assign _T_65812 = _T_65811[10:0]; // @[Modules.scala 68:83:@15847.4]
  assign buffer_6_588 = $signed(_T_65812); // @[Modules.scala 68:83:@15848.4]
  assign _T_65814 = $signed(buffer_6_394) + $signed(buffer_0_395); // @[Modules.scala 68:83:@15850.4]
  assign _T_65815 = _T_65814[10:0]; // @[Modules.scala 68:83:@15851.4]
  assign buffer_6_589 = $signed(_T_65815); // @[Modules.scala 68:83:@15852.4]
  assign _T_65817 = $signed(buffer_1_396) + $signed(buffer_4_397); // @[Modules.scala 68:83:@15854.4]
  assign _T_65818 = _T_65817[10:0]; // @[Modules.scala 68:83:@15855.4]
  assign buffer_6_590 = $signed(_T_65818); // @[Modules.scala 68:83:@15856.4]
  assign _T_65820 = $signed(buffer_1_398) + $signed(buffer_0_399); // @[Modules.scala 68:83:@15858.4]
  assign _T_65821 = _T_65820[10:0]; // @[Modules.scala 68:83:@15859.4]
  assign buffer_6_591 = $signed(_T_65821); // @[Modules.scala 68:83:@15860.4]
  assign _T_65823 = $signed(buffer_3_400) + $signed(buffer_0_395); // @[Modules.scala 68:83:@15862.4]
  assign _T_65824 = _T_65823[10:0]; // @[Modules.scala 68:83:@15863.4]
  assign buffer_6_592 = $signed(_T_65824); // @[Modules.scala 68:83:@15864.4]
  assign _T_65829 = $signed(buffer_0_395) + $signed(buffer_6_405); // @[Modules.scala 68:83:@15870.4]
  assign _T_65830 = _T_65829[10:0]; // @[Modules.scala 68:83:@15871.4]
  assign buffer_6_594 = $signed(_T_65830); // @[Modules.scala 68:83:@15872.4]
  assign _T_65832 = $signed(buffer_6_406) + $signed(buffer_0_395); // @[Modules.scala 68:83:@15874.4]
  assign _T_65833 = _T_65832[10:0]; // @[Modules.scala 68:83:@15875.4]
  assign buffer_6_595 = $signed(_T_65833); // @[Modules.scala 68:83:@15876.4]
  assign _T_65841 = $signed(buffer_2_412) + $signed(buffer_6_413); // @[Modules.scala 68:83:@15886.4]
  assign _T_65842 = _T_65841[10:0]; // @[Modules.scala 68:83:@15887.4]
  assign buffer_6_598 = $signed(_T_65842); // @[Modules.scala 68:83:@15888.4]
  assign _T_65850 = $signed(buffer_6_418) + $signed(buffer_6_419); // @[Modules.scala 68:83:@15898.4]
  assign _T_65851 = _T_65850[10:0]; // @[Modules.scala 68:83:@15899.4]
  assign buffer_6_601 = $signed(_T_65851); // @[Modules.scala 68:83:@15900.4]
  assign _T_65853 = $signed(buffer_5_420) + $signed(buffer_0_395); // @[Modules.scala 68:83:@15902.4]
  assign _T_65854 = _T_65853[10:0]; // @[Modules.scala 68:83:@15903.4]
  assign buffer_6_602 = $signed(_T_65854); // @[Modules.scala 68:83:@15904.4]
  assign _T_65859 = $signed(buffer_0_395) + $signed(buffer_0_425); // @[Modules.scala 68:83:@15910.4]
  assign _T_65860 = _T_65859[10:0]; // @[Modules.scala 68:83:@15911.4]
  assign buffer_6_604 = $signed(_T_65860); // @[Modules.scala 68:83:@15912.4]
  assign _T_65862 = $signed(buffer_0_426) + $signed(buffer_4_427); // @[Modules.scala 68:83:@15914.4]
  assign _T_65863 = _T_65862[10:0]; // @[Modules.scala 68:83:@15915.4]
  assign buffer_6_605 = $signed(_T_65863); // @[Modules.scala 68:83:@15916.4]
  assign _T_65865 = $signed(buffer_6_428) + $signed(buffer_6_429); // @[Modules.scala 68:83:@15918.4]
  assign _T_65866 = _T_65865[10:0]; // @[Modules.scala 68:83:@15919.4]
  assign buffer_6_606 = $signed(_T_65866); // @[Modules.scala 68:83:@15920.4]
  assign _T_65871 = $signed(buffer_0_432) + $signed(buffer_6_433); // @[Modules.scala 68:83:@15926.4]
  assign _T_65872 = _T_65871[10:0]; // @[Modules.scala 68:83:@15927.4]
  assign buffer_6_608 = $signed(_T_65872); // @[Modules.scala 68:83:@15928.4]
  assign _T_65874 = $signed(buffer_2_434) + $signed(buffer_6_435); // @[Modules.scala 68:83:@15930.4]
  assign _T_65875 = _T_65874[10:0]; // @[Modules.scala 68:83:@15931.4]
  assign buffer_6_609 = $signed(_T_65875); // @[Modules.scala 68:83:@15932.4]
  assign _T_65877 = $signed(buffer_6_436) + $signed(buffer_1_437); // @[Modules.scala 68:83:@15934.4]
  assign _T_65878 = _T_65877[10:0]; // @[Modules.scala 68:83:@15935.4]
  assign buffer_6_610 = $signed(_T_65878); // @[Modules.scala 68:83:@15936.4]
  assign _T_65880 = $signed(buffer_3_438) + $signed(buffer_6_439); // @[Modules.scala 68:83:@15938.4]
  assign _T_65881 = _T_65880[10:0]; // @[Modules.scala 68:83:@15939.4]
  assign buffer_6_611 = $signed(_T_65881); // @[Modules.scala 68:83:@15940.4]
  assign _T_65883 = $signed(buffer_6_440) + $signed(buffer_6_441); // @[Modules.scala 68:83:@15942.4]
  assign _T_65884 = _T_65883[10:0]; // @[Modules.scala 68:83:@15943.4]
  assign buffer_6_612 = $signed(_T_65884); // @[Modules.scala 68:83:@15944.4]
  assign _T_65886 = $signed(buffer_6_442) + $signed(buffer_6_443); // @[Modules.scala 68:83:@15946.4]
  assign _T_65887 = _T_65886[10:0]; // @[Modules.scala 68:83:@15947.4]
  assign buffer_6_613 = $signed(_T_65887); // @[Modules.scala 68:83:@15948.4]
  assign _T_65889 = $signed(buffer_6_444) + $signed(buffer_6_445); // @[Modules.scala 68:83:@15950.4]
  assign _T_65890 = _T_65889[10:0]; // @[Modules.scala 68:83:@15951.4]
  assign buffer_6_614 = $signed(_T_65890); // @[Modules.scala 68:83:@15952.4]
  assign _T_65892 = $signed(buffer_6_446) + $signed(buffer_5_447); // @[Modules.scala 68:83:@15954.4]
  assign _T_65893 = _T_65892[10:0]; // @[Modules.scala 68:83:@15955.4]
  assign buffer_6_615 = $signed(_T_65893); // @[Modules.scala 68:83:@15956.4]
  assign _T_65895 = $signed(buffer_6_448) + $signed(buffer_3_449); // @[Modules.scala 68:83:@15958.4]
  assign _T_65896 = _T_65895[10:0]; // @[Modules.scala 68:83:@15959.4]
  assign buffer_6_616 = $signed(_T_65896); // @[Modules.scala 68:83:@15960.4]
  assign _T_65898 = $signed(buffer_6_450) + $signed(buffer_3_451); // @[Modules.scala 68:83:@15962.4]
  assign _T_65899 = _T_65898[10:0]; // @[Modules.scala 68:83:@15963.4]
  assign buffer_6_617 = $signed(_T_65899); // @[Modules.scala 68:83:@15964.4]
  assign _T_65901 = $signed(buffer_6_452) + $signed(buffer_6_453); // @[Modules.scala 68:83:@15966.4]
  assign _T_65902 = _T_65901[10:0]; // @[Modules.scala 68:83:@15967.4]
  assign buffer_6_618 = $signed(_T_65902); // @[Modules.scala 68:83:@15968.4]
  assign _T_65904 = $signed(buffer_0_395) + $signed(buffer_6_455); // @[Modules.scala 68:83:@15970.4]
  assign _T_65905 = _T_65904[10:0]; // @[Modules.scala 68:83:@15971.4]
  assign buffer_6_619 = $signed(_T_65905); // @[Modules.scala 68:83:@15972.4]
  assign _T_65907 = $signed(buffer_6_456) + $signed(buffer_6_457); // @[Modules.scala 68:83:@15974.4]
  assign _T_65908 = _T_65907[10:0]; // @[Modules.scala 68:83:@15975.4]
  assign buffer_6_620 = $signed(_T_65908); // @[Modules.scala 68:83:@15976.4]
  assign _T_65913 = $signed(buffer_6_460) + $signed(buffer_0_395); // @[Modules.scala 68:83:@15982.4]
  assign _T_65914 = _T_65913[10:0]; // @[Modules.scala 68:83:@15983.4]
  assign buffer_6_622 = $signed(_T_65914); // @[Modules.scala 68:83:@15984.4]
  assign _T_65916 = $signed(buffer_6_462) + $signed(buffer_0_395); // @[Modules.scala 68:83:@15986.4]
  assign _T_65917 = _T_65916[10:0]; // @[Modules.scala 68:83:@15987.4]
  assign buffer_6_623 = $signed(_T_65917); // @[Modules.scala 68:83:@15988.4]
  assign _T_65919 = $signed(buffer_6_464) + $signed(buffer_6_465); // @[Modules.scala 68:83:@15990.4]
  assign _T_65920 = _T_65919[10:0]; // @[Modules.scala 68:83:@15991.4]
  assign buffer_6_624 = $signed(_T_65920); // @[Modules.scala 68:83:@15992.4]
  assign _T_65922 = $signed(buffer_6_466) + $signed(buffer_6_467); // @[Modules.scala 68:83:@15994.4]
  assign _T_65923 = _T_65922[10:0]; // @[Modules.scala 68:83:@15995.4]
  assign buffer_6_625 = $signed(_T_65923); // @[Modules.scala 68:83:@15996.4]
  assign _T_65925 = $signed(buffer_0_395) + $signed(buffer_6_469); // @[Modules.scala 68:83:@15998.4]
  assign _T_65926 = _T_65925[10:0]; // @[Modules.scala 68:83:@15999.4]
  assign buffer_6_626 = $signed(_T_65926); // @[Modules.scala 68:83:@16000.4]
  assign _T_65928 = $signed(buffer_6_470) + $signed(buffer_6_471); // @[Modules.scala 68:83:@16002.4]
  assign _T_65929 = _T_65928[10:0]; // @[Modules.scala 68:83:@16003.4]
  assign buffer_6_627 = $signed(_T_65929); // @[Modules.scala 68:83:@16004.4]
  assign _T_65931 = $signed(buffer_6_472) + $signed(buffer_6_473); // @[Modules.scala 68:83:@16006.4]
  assign _T_65932 = _T_65931[10:0]; // @[Modules.scala 68:83:@16007.4]
  assign buffer_6_628 = $signed(_T_65932); // @[Modules.scala 68:83:@16008.4]
  assign _T_65934 = $signed(buffer_0_474) + $signed(buffer_0_395); // @[Modules.scala 68:83:@16010.4]
  assign _T_65935 = _T_65934[10:0]; // @[Modules.scala 68:83:@16011.4]
  assign buffer_6_629 = $signed(_T_65935); // @[Modules.scala 68:83:@16012.4]
  assign _T_65937 = $signed(buffer_6_476) + $signed(buffer_6_477); // @[Modules.scala 68:83:@16014.4]
  assign _T_65938 = _T_65937[10:0]; // @[Modules.scala 68:83:@16015.4]
  assign buffer_6_630 = $signed(_T_65938); // @[Modules.scala 68:83:@16016.4]
  assign _T_65940 = $signed(buffer_6_478) + $signed(buffer_6_479); // @[Modules.scala 68:83:@16018.4]
  assign _T_65941 = _T_65940[10:0]; // @[Modules.scala 68:83:@16019.4]
  assign buffer_6_631 = $signed(_T_65941); // @[Modules.scala 68:83:@16020.4]
  assign _T_65943 = $signed(buffer_0_480) + $signed(buffer_6_481); // @[Modules.scala 68:83:@16022.4]
  assign _T_65944 = _T_65943[10:0]; // @[Modules.scala 68:83:@16023.4]
  assign buffer_6_632 = $signed(_T_65944); // @[Modules.scala 68:83:@16024.4]
  assign _T_65946 = $signed(buffer_0_482) + $signed(buffer_6_483); // @[Modules.scala 68:83:@16026.4]
  assign _T_65947 = _T_65946[10:0]; // @[Modules.scala 68:83:@16027.4]
  assign buffer_6_633 = $signed(_T_65947); // @[Modules.scala 68:83:@16028.4]
  assign _T_65949 = $signed(buffer_0_484) + $signed(buffer_6_485); // @[Modules.scala 68:83:@16030.4]
  assign _T_65950 = _T_65949[10:0]; // @[Modules.scala 68:83:@16031.4]
  assign buffer_6_634 = $signed(_T_65950); // @[Modules.scala 68:83:@16032.4]
  assign _T_65952 = $signed(buffer_6_486) + $signed(buffer_0_487); // @[Modules.scala 68:83:@16034.4]
  assign _T_65953 = _T_65952[10:0]; // @[Modules.scala 68:83:@16035.4]
  assign buffer_6_635 = $signed(_T_65953); // @[Modules.scala 68:83:@16036.4]
  assign _T_65955 = $signed(buffer_2_488) + $signed(buffer_5_489); // @[Modules.scala 68:83:@16038.4]
  assign _T_65956 = _T_65955[10:0]; // @[Modules.scala 68:83:@16039.4]
  assign buffer_6_636 = $signed(_T_65956); // @[Modules.scala 68:83:@16040.4]
  assign _T_65958 = $signed(buffer_6_490) + $signed(buffer_0_491); // @[Modules.scala 68:83:@16042.4]
  assign _T_65959 = _T_65958[10:0]; // @[Modules.scala 68:83:@16043.4]
  assign buffer_6_637 = $signed(_T_65959); // @[Modules.scala 68:83:@16044.4]
  assign _T_65961 = $signed(buffer_6_492) + $signed(buffer_6_493); // @[Modules.scala 68:83:@16046.4]
  assign _T_65962 = _T_65961[10:0]; // @[Modules.scala 68:83:@16047.4]
  assign buffer_6_638 = $signed(_T_65962); // @[Modules.scala 68:83:@16048.4]
  assign _T_65964 = $signed(buffer_0_494) + $signed(buffer_6_495); // @[Modules.scala 68:83:@16050.4]
  assign _T_65965 = _T_65964[10:0]; // @[Modules.scala 68:83:@16051.4]
  assign buffer_6_639 = $signed(_T_65965); // @[Modules.scala 68:83:@16052.4]
  assign _T_65967 = $signed(buffer_6_496) + $signed(buffer_6_497); // @[Modules.scala 68:83:@16054.4]
  assign _T_65968 = _T_65967[10:0]; // @[Modules.scala 68:83:@16055.4]
  assign buffer_6_640 = $signed(_T_65968); // @[Modules.scala 68:83:@16056.4]
  assign _T_65970 = $signed(buffer_6_498) + $signed(buffer_6_499); // @[Modules.scala 68:83:@16058.4]
  assign _T_65971 = _T_65970[10:0]; // @[Modules.scala 68:83:@16059.4]
  assign buffer_6_641 = $signed(_T_65971); // @[Modules.scala 68:83:@16060.4]
  assign _T_65973 = $signed(buffer_6_500) + $signed(buffer_6_501); // @[Modules.scala 68:83:@16062.4]
  assign _T_65974 = _T_65973[10:0]; // @[Modules.scala 68:83:@16063.4]
  assign buffer_6_642 = $signed(_T_65974); // @[Modules.scala 68:83:@16064.4]
  assign _T_65976 = $signed(buffer_6_502) + $signed(buffer_0_395); // @[Modules.scala 68:83:@16066.4]
  assign _T_65977 = _T_65976[10:0]; // @[Modules.scala 68:83:@16067.4]
  assign buffer_6_643 = $signed(_T_65977); // @[Modules.scala 68:83:@16068.4]
  assign _T_65979 = $signed(buffer_6_504) + $signed(buffer_3_505); // @[Modules.scala 68:83:@16070.4]
  assign _T_65980 = _T_65979[10:0]; // @[Modules.scala 68:83:@16071.4]
  assign buffer_6_644 = $signed(_T_65980); // @[Modules.scala 68:83:@16072.4]
  assign _T_65982 = $signed(buffer_6_506) + $signed(buffer_6_507); // @[Modules.scala 68:83:@16074.4]
  assign _T_65983 = _T_65982[10:0]; // @[Modules.scala 68:83:@16075.4]
  assign buffer_6_645 = $signed(_T_65983); // @[Modules.scala 68:83:@16076.4]
  assign _T_65985 = $signed(buffer_6_508) + $signed(buffer_6_509); // @[Modules.scala 68:83:@16078.4]
  assign _T_65986 = _T_65985[10:0]; // @[Modules.scala 68:83:@16079.4]
  assign buffer_6_646 = $signed(_T_65986); // @[Modules.scala 68:83:@16080.4]
  assign _T_65988 = $signed(buffer_0_395) + $signed(buffer_6_511); // @[Modules.scala 68:83:@16082.4]
  assign _T_65989 = _T_65988[10:0]; // @[Modules.scala 68:83:@16083.4]
  assign buffer_6_647 = $signed(_T_65989); // @[Modules.scala 68:83:@16084.4]
  assign _T_65991 = $signed(buffer_6_512) + $signed(buffer_6_513); // @[Modules.scala 68:83:@16086.4]
  assign _T_65992 = _T_65991[10:0]; // @[Modules.scala 68:83:@16087.4]
  assign buffer_6_648 = $signed(_T_65992); // @[Modules.scala 68:83:@16088.4]
  assign _T_65994 = $signed(buffer_2_514) + $signed(buffer_6_515); // @[Modules.scala 68:83:@16090.4]
  assign _T_65995 = _T_65994[10:0]; // @[Modules.scala 68:83:@16091.4]
  assign buffer_6_649 = $signed(_T_65995); // @[Modules.scala 68:83:@16092.4]
  assign _T_66000 = $signed(buffer_6_518) + $signed(buffer_0_395); // @[Modules.scala 68:83:@16098.4]
  assign _T_66001 = _T_66000[10:0]; // @[Modules.scala 68:83:@16099.4]
  assign buffer_6_651 = $signed(_T_66001); // @[Modules.scala 68:83:@16100.4]
  assign _T_66003 = $signed(buffer_0_395) + $signed(buffer_6_521); // @[Modules.scala 68:83:@16102.4]
  assign _T_66004 = _T_66003[10:0]; // @[Modules.scala 68:83:@16103.4]
  assign buffer_6_652 = $signed(_T_66004); // @[Modules.scala 68:83:@16104.4]
  assign _T_66018 = $signed(buffer_0_395) + $signed(buffer_2_531); // @[Modules.scala 68:83:@16122.4]
  assign _T_66019 = _T_66018[10:0]; // @[Modules.scala 68:83:@16123.4]
  assign buffer_6_657 = $signed(_T_66019); // @[Modules.scala 68:83:@16124.4]
  assign _T_66030 = $signed(buffer_0_395) + $signed(buffer_6_539); // @[Modules.scala 68:83:@16138.4]
  assign _T_66031 = _T_66030[10:0]; // @[Modules.scala 68:83:@16139.4]
  assign buffer_6_661 = $signed(_T_66031); // @[Modules.scala 68:83:@16140.4]
  assign _T_66039 = $signed(buffer_0_395) + $signed(buffer_6_545); // @[Modules.scala 68:83:@16150.4]
  assign _T_66040 = _T_66039[10:0]; // @[Modules.scala 68:83:@16151.4]
  assign buffer_6_664 = $signed(_T_66040); // @[Modules.scala 68:83:@16152.4]
  assign _T_66045 = $signed(buffer_6_548) + $signed(buffer_6_549); // @[Modules.scala 68:83:@16158.4]
  assign _T_66046 = _T_66045[10:0]; // @[Modules.scala 68:83:@16159.4]
  assign buffer_6_666 = $signed(_T_66046); // @[Modules.scala 68:83:@16160.4]
  assign _T_66051 = $signed(buffer_0_552) + $signed(buffer_0_395); // @[Modules.scala 68:83:@16166.4]
  assign _T_66052 = _T_66051[10:0]; // @[Modules.scala 68:83:@16167.4]
  assign buffer_6_668 = $signed(_T_66052); // @[Modules.scala 68:83:@16168.4]
  assign _T_66054 = $signed(buffer_6_554) + $signed(buffer_6_555); // @[Modules.scala 68:83:@16170.4]
  assign _T_66055 = _T_66054[10:0]; // @[Modules.scala 68:83:@16171.4]
  assign buffer_6_669 = $signed(_T_66055); // @[Modules.scala 68:83:@16172.4]
  assign _T_66060 = $signed(buffer_0_395) + $signed(buffer_6_559); // @[Modules.scala 68:83:@16178.4]
  assign _T_66061 = _T_66060[10:0]; // @[Modules.scala 68:83:@16179.4]
  assign buffer_6_671 = $signed(_T_66061); // @[Modules.scala 68:83:@16180.4]
  assign _T_66063 = $signed(buffer_6_560) + $signed(buffer_5_561); // @[Modules.scala 68:83:@16182.4]
  assign _T_66064 = _T_66063[10:0]; // @[Modules.scala 68:83:@16183.4]
  assign buffer_6_672 = $signed(_T_66064); // @[Modules.scala 68:83:@16184.4]
  assign _T_66069 = $signed(buffer_6_564) + $signed(buffer_6_565); // @[Modules.scala 68:83:@16190.4]
  assign _T_66070 = _T_66069[10:0]; // @[Modules.scala 68:83:@16191.4]
  assign buffer_6_674 = $signed(_T_66070); // @[Modules.scala 68:83:@16192.4]
  assign _T_66072 = $signed(buffer_2_566) + $signed(buffer_3_567); // @[Modules.scala 68:83:@16194.4]
  assign _T_66073 = _T_66072[10:0]; // @[Modules.scala 68:83:@16195.4]
  assign buffer_6_675 = $signed(_T_66073); // @[Modules.scala 68:83:@16196.4]
  assign _T_66075 = $signed(buffer_0_568) + $signed(buffer_6_569); // @[Modules.scala 68:83:@16198.4]
  assign _T_66076 = _T_66075[10:0]; // @[Modules.scala 68:83:@16199.4]
  assign buffer_6_676 = $signed(_T_66076); // @[Modules.scala 68:83:@16200.4]
  assign _T_66078 = $signed(buffer_6_570) + $signed(buffer_6_571); // @[Modules.scala 68:83:@16202.4]
  assign _T_66079 = _T_66078[10:0]; // @[Modules.scala 68:83:@16203.4]
  assign buffer_6_677 = $signed(_T_66079); // @[Modules.scala 68:83:@16204.4]
  assign _T_66081 = $signed(buffer_0_572) + $signed(buffer_0_395); // @[Modules.scala 68:83:@16206.4]
  assign _T_66082 = _T_66081[10:0]; // @[Modules.scala 68:83:@16207.4]
  assign buffer_6_678 = $signed(_T_66082); // @[Modules.scala 68:83:@16208.4]
  assign _T_66084 = $signed(buffer_6_574) + $signed(buffer_0_575); // @[Modules.scala 68:83:@16210.4]
  assign _T_66085 = _T_66084[10:0]; // @[Modules.scala 68:83:@16211.4]
  assign buffer_6_679 = $signed(_T_66085); // @[Modules.scala 68:83:@16212.4]
  assign _T_66090 = $signed(buffer_3_578) + $signed(buffer_6_579); // @[Modules.scala 68:83:@16218.4]
  assign _T_66091 = _T_66090[10:0]; // @[Modules.scala 68:83:@16219.4]
  assign buffer_6_681 = $signed(_T_66091); // @[Modules.scala 68:83:@16220.4]
  assign _T_66093 = $signed(buffer_3_580) + $signed(buffer_4_581); // @[Modules.scala 68:83:@16222.4]
  assign _T_66094 = _T_66093[10:0]; // @[Modules.scala 68:83:@16223.4]
  assign buffer_6_682 = $signed(_T_66094); // @[Modules.scala 68:83:@16224.4]
  assign _T_66099 = $signed(buffer_6_584) + $signed(buffer_0_395); // @[Modules.scala 68:83:@16230.4]
  assign _T_66100 = _T_66099[10:0]; // @[Modules.scala 68:83:@16231.4]
  assign buffer_6_684 = $signed(_T_66100); // @[Modules.scala 68:83:@16232.4]
  assign _T_66102 = $signed(buffer_6_586) + $signed(buffer_4_587); // @[Modules.scala 68:83:@16234.4]
  assign _T_66103 = _T_66102[10:0]; // @[Modules.scala 68:83:@16235.4]
  assign buffer_6_685 = $signed(_T_66103); // @[Modules.scala 68:83:@16236.4]
  assign _T_66105 = $signed(buffer_6_588) + $signed(buffer_6_589); // @[Modules.scala 71:109:@16238.4]
  assign _T_66106 = _T_66105[10:0]; // @[Modules.scala 71:109:@16239.4]
  assign buffer_6_686 = $signed(_T_66106); // @[Modules.scala 71:109:@16240.4]
  assign _T_66108 = $signed(buffer_6_590) + $signed(buffer_6_591); // @[Modules.scala 71:109:@16242.4]
  assign _T_66109 = _T_66108[10:0]; // @[Modules.scala 71:109:@16243.4]
  assign buffer_6_687 = $signed(_T_66109); // @[Modules.scala 71:109:@16244.4]
  assign _T_66111 = $signed(buffer_6_592) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16246.4]
  assign _T_66112 = _T_66111[10:0]; // @[Modules.scala 71:109:@16247.4]
  assign buffer_6_688 = $signed(_T_66112); // @[Modules.scala 71:109:@16248.4]
  assign _T_66114 = $signed(buffer_6_594) + $signed(buffer_6_595); // @[Modules.scala 71:109:@16250.4]
  assign _T_66115 = _T_66114[10:0]; // @[Modules.scala 71:109:@16251.4]
  assign buffer_6_689 = $signed(_T_66115); // @[Modules.scala 71:109:@16252.4]
  assign _T_66120 = $signed(buffer_6_598) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16258.4]
  assign _T_66121 = _T_66120[10:0]; // @[Modules.scala 71:109:@16259.4]
  assign buffer_6_691 = $signed(_T_66121); // @[Modules.scala 71:109:@16260.4]
  assign _T_66123 = $signed(buffer_0_593) + $signed(buffer_6_601); // @[Modules.scala 71:109:@16262.4]
  assign _T_66124 = _T_66123[10:0]; // @[Modules.scala 71:109:@16263.4]
  assign buffer_6_692 = $signed(_T_66124); // @[Modules.scala 71:109:@16264.4]
  assign _T_66126 = $signed(buffer_6_602) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16266.4]
  assign _T_66127 = _T_66126[10:0]; // @[Modules.scala 71:109:@16267.4]
  assign buffer_6_693 = $signed(_T_66127); // @[Modules.scala 71:109:@16268.4]
  assign _T_66129 = $signed(buffer_6_604) + $signed(buffer_6_605); // @[Modules.scala 71:109:@16270.4]
  assign _T_66130 = _T_66129[10:0]; // @[Modules.scala 71:109:@16271.4]
  assign buffer_6_694 = $signed(_T_66130); // @[Modules.scala 71:109:@16272.4]
  assign _T_66132 = $signed(buffer_6_606) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16274.4]
  assign _T_66133 = _T_66132[10:0]; // @[Modules.scala 71:109:@16275.4]
  assign buffer_6_695 = $signed(_T_66133); // @[Modules.scala 71:109:@16276.4]
  assign _T_66135 = $signed(buffer_6_608) + $signed(buffer_6_609); // @[Modules.scala 71:109:@16278.4]
  assign _T_66136 = _T_66135[10:0]; // @[Modules.scala 71:109:@16279.4]
  assign buffer_6_696 = $signed(_T_66136); // @[Modules.scala 71:109:@16280.4]
  assign _T_66138 = $signed(buffer_6_610) + $signed(buffer_6_611); // @[Modules.scala 71:109:@16282.4]
  assign _T_66139 = _T_66138[10:0]; // @[Modules.scala 71:109:@16283.4]
  assign buffer_6_697 = $signed(_T_66139); // @[Modules.scala 71:109:@16284.4]
  assign _T_66141 = $signed(buffer_6_612) + $signed(buffer_6_613); // @[Modules.scala 71:109:@16286.4]
  assign _T_66142 = _T_66141[10:0]; // @[Modules.scala 71:109:@16287.4]
  assign buffer_6_698 = $signed(_T_66142); // @[Modules.scala 71:109:@16288.4]
  assign _T_66144 = $signed(buffer_6_614) + $signed(buffer_6_615); // @[Modules.scala 71:109:@16290.4]
  assign _T_66145 = _T_66144[10:0]; // @[Modules.scala 71:109:@16291.4]
  assign buffer_6_699 = $signed(_T_66145); // @[Modules.scala 71:109:@16292.4]
  assign _T_66147 = $signed(buffer_6_616) + $signed(buffer_6_617); // @[Modules.scala 71:109:@16294.4]
  assign _T_66148 = _T_66147[10:0]; // @[Modules.scala 71:109:@16295.4]
  assign buffer_6_700 = $signed(_T_66148); // @[Modules.scala 71:109:@16296.4]
  assign _T_66150 = $signed(buffer_6_618) + $signed(buffer_6_619); // @[Modules.scala 71:109:@16298.4]
  assign _T_66151 = _T_66150[10:0]; // @[Modules.scala 71:109:@16299.4]
  assign buffer_6_701 = $signed(_T_66151); // @[Modules.scala 71:109:@16300.4]
  assign _T_66153 = $signed(buffer_6_620) + $signed(buffer_3_621); // @[Modules.scala 71:109:@16302.4]
  assign _T_66154 = _T_66153[10:0]; // @[Modules.scala 71:109:@16303.4]
  assign buffer_6_702 = $signed(_T_66154); // @[Modules.scala 71:109:@16304.4]
  assign _T_66156 = $signed(buffer_6_622) + $signed(buffer_6_623); // @[Modules.scala 71:109:@16306.4]
  assign _T_66157 = _T_66156[10:0]; // @[Modules.scala 71:109:@16307.4]
  assign buffer_6_703 = $signed(_T_66157); // @[Modules.scala 71:109:@16308.4]
  assign _T_66159 = $signed(buffer_6_624) + $signed(buffer_6_625); // @[Modules.scala 71:109:@16310.4]
  assign _T_66160 = _T_66159[10:0]; // @[Modules.scala 71:109:@16311.4]
  assign buffer_6_704 = $signed(_T_66160); // @[Modules.scala 71:109:@16312.4]
  assign _T_66162 = $signed(buffer_6_626) + $signed(buffer_6_627); // @[Modules.scala 71:109:@16314.4]
  assign _T_66163 = _T_66162[10:0]; // @[Modules.scala 71:109:@16315.4]
  assign buffer_6_705 = $signed(_T_66163); // @[Modules.scala 71:109:@16316.4]
  assign _T_66165 = $signed(buffer_6_628) + $signed(buffer_6_629); // @[Modules.scala 71:109:@16318.4]
  assign _T_66166 = _T_66165[10:0]; // @[Modules.scala 71:109:@16319.4]
  assign buffer_6_706 = $signed(_T_66166); // @[Modules.scala 71:109:@16320.4]
  assign _T_66168 = $signed(buffer_6_630) + $signed(buffer_6_631); // @[Modules.scala 71:109:@16322.4]
  assign _T_66169 = _T_66168[10:0]; // @[Modules.scala 71:109:@16323.4]
  assign buffer_6_707 = $signed(_T_66169); // @[Modules.scala 71:109:@16324.4]
  assign _T_66171 = $signed(buffer_6_632) + $signed(buffer_6_633); // @[Modules.scala 71:109:@16326.4]
  assign _T_66172 = _T_66171[10:0]; // @[Modules.scala 71:109:@16327.4]
  assign buffer_6_708 = $signed(_T_66172); // @[Modules.scala 71:109:@16328.4]
  assign _T_66174 = $signed(buffer_6_634) + $signed(buffer_6_635); // @[Modules.scala 71:109:@16330.4]
  assign _T_66175 = _T_66174[10:0]; // @[Modules.scala 71:109:@16331.4]
  assign buffer_6_709 = $signed(_T_66175); // @[Modules.scala 71:109:@16332.4]
  assign _T_66177 = $signed(buffer_6_636) + $signed(buffer_6_637); // @[Modules.scala 71:109:@16334.4]
  assign _T_66178 = _T_66177[10:0]; // @[Modules.scala 71:109:@16335.4]
  assign buffer_6_710 = $signed(_T_66178); // @[Modules.scala 71:109:@16336.4]
  assign _T_66180 = $signed(buffer_6_638) + $signed(buffer_6_639); // @[Modules.scala 71:109:@16338.4]
  assign _T_66181 = _T_66180[10:0]; // @[Modules.scala 71:109:@16339.4]
  assign buffer_6_711 = $signed(_T_66181); // @[Modules.scala 71:109:@16340.4]
  assign _T_66183 = $signed(buffer_6_640) + $signed(buffer_6_641); // @[Modules.scala 71:109:@16342.4]
  assign _T_66184 = _T_66183[10:0]; // @[Modules.scala 71:109:@16343.4]
  assign buffer_6_712 = $signed(_T_66184); // @[Modules.scala 71:109:@16344.4]
  assign _T_66186 = $signed(buffer_6_642) + $signed(buffer_6_643); // @[Modules.scala 71:109:@16346.4]
  assign _T_66187 = _T_66186[10:0]; // @[Modules.scala 71:109:@16347.4]
  assign buffer_6_713 = $signed(_T_66187); // @[Modules.scala 71:109:@16348.4]
  assign _T_66189 = $signed(buffer_6_644) + $signed(buffer_6_645); // @[Modules.scala 71:109:@16350.4]
  assign _T_66190 = _T_66189[10:0]; // @[Modules.scala 71:109:@16351.4]
  assign buffer_6_714 = $signed(_T_66190); // @[Modules.scala 71:109:@16352.4]
  assign _T_66192 = $signed(buffer_6_646) + $signed(buffer_6_647); // @[Modules.scala 71:109:@16354.4]
  assign _T_66193 = _T_66192[10:0]; // @[Modules.scala 71:109:@16355.4]
  assign buffer_6_715 = $signed(_T_66193); // @[Modules.scala 71:109:@16356.4]
  assign _T_66195 = $signed(buffer_6_648) + $signed(buffer_6_649); // @[Modules.scala 71:109:@16358.4]
  assign _T_66196 = _T_66195[10:0]; // @[Modules.scala 71:109:@16359.4]
  assign buffer_6_716 = $signed(_T_66196); // @[Modules.scala 71:109:@16360.4]
  assign _T_66198 = $signed(buffer_0_593) + $signed(buffer_6_651); // @[Modules.scala 71:109:@16362.4]
  assign _T_66199 = _T_66198[10:0]; // @[Modules.scala 71:109:@16363.4]
  assign buffer_6_717 = $signed(_T_66199); // @[Modules.scala 71:109:@16364.4]
  assign _T_66201 = $signed(buffer_6_652) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16366.4]
  assign _T_66202 = _T_66201[10:0]; // @[Modules.scala 71:109:@16367.4]
  assign buffer_6_718 = $signed(_T_66202); // @[Modules.scala 71:109:@16368.4]
  assign _T_66207 = $signed(buffer_0_593) + $signed(buffer_6_657); // @[Modules.scala 71:109:@16374.4]
  assign _T_66208 = _T_66207[10:0]; // @[Modules.scala 71:109:@16375.4]
  assign buffer_6_720 = $signed(_T_66208); // @[Modules.scala 71:109:@16376.4]
  assign _T_66213 = $signed(buffer_0_593) + $signed(buffer_6_661); // @[Modules.scala 71:109:@16382.4]
  assign _T_66214 = _T_66213[10:0]; // @[Modules.scala 71:109:@16383.4]
  assign buffer_6_722 = $signed(_T_66214); // @[Modules.scala 71:109:@16384.4]
  assign _T_66219 = $signed(buffer_6_664) + $signed(buffer_2_665); // @[Modules.scala 71:109:@16390.4]
  assign _T_66220 = _T_66219[10:0]; // @[Modules.scala 71:109:@16391.4]
  assign buffer_6_724 = $signed(_T_66220); // @[Modules.scala 71:109:@16392.4]
  assign _T_66222 = $signed(buffer_6_666) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16394.4]
  assign _T_66223 = _T_66222[10:0]; // @[Modules.scala 71:109:@16395.4]
  assign buffer_6_725 = $signed(_T_66223); // @[Modules.scala 71:109:@16396.4]
  assign _T_66225 = $signed(buffer_6_668) + $signed(buffer_6_669); // @[Modules.scala 71:109:@16398.4]
  assign _T_66226 = _T_66225[10:0]; // @[Modules.scala 71:109:@16399.4]
  assign buffer_6_726 = $signed(_T_66226); // @[Modules.scala 71:109:@16400.4]
  assign _T_66228 = $signed(buffer_0_593) + $signed(buffer_6_671); // @[Modules.scala 71:109:@16402.4]
  assign _T_66229 = _T_66228[10:0]; // @[Modules.scala 71:109:@16403.4]
  assign buffer_6_727 = $signed(_T_66229); // @[Modules.scala 71:109:@16404.4]
  assign _T_66231 = $signed(buffer_6_672) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16406.4]
  assign _T_66232 = _T_66231[10:0]; // @[Modules.scala 71:109:@16407.4]
  assign buffer_6_728 = $signed(_T_66232); // @[Modules.scala 71:109:@16408.4]
  assign _T_66234 = $signed(buffer_6_674) + $signed(buffer_6_675); // @[Modules.scala 71:109:@16410.4]
  assign _T_66235 = _T_66234[10:0]; // @[Modules.scala 71:109:@16411.4]
  assign buffer_6_729 = $signed(_T_66235); // @[Modules.scala 71:109:@16412.4]
  assign _T_66237 = $signed(buffer_6_676) + $signed(buffer_6_677); // @[Modules.scala 71:109:@16414.4]
  assign _T_66238 = _T_66237[10:0]; // @[Modules.scala 71:109:@16415.4]
  assign buffer_6_730 = $signed(_T_66238); // @[Modules.scala 71:109:@16416.4]
  assign _T_66240 = $signed(buffer_6_678) + $signed(buffer_6_679); // @[Modules.scala 71:109:@16418.4]
  assign _T_66241 = _T_66240[10:0]; // @[Modules.scala 71:109:@16419.4]
  assign buffer_6_731 = $signed(_T_66241); // @[Modules.scala 71:109:@16420.4]
  assign _T_66243 = $signed(buffer_5_680) + $signed(buffer_6_681); // @[Modules.scala 71:109:@16422.4]
  assign _T_66244 = _T_66243[10:0]; // @[Modules.scala 71:109:@16423.4]
  assign buffer_6_732 = $signed(_T_66244); // @[Modules.scala 71:109:@16424.4]
  assign _T_66246 = $signed(buffer_6_682) + $signed(buffer_0_593); // @[Modules.scala 71:109:@16426.4]
  assign _T_66247 = _T_66246[10:0]; // @[Modules.scala 71:109:@16427.4]
  assign buffer_6_733 = $signed(_T_66247); // @[Modules.scala 71:109:@16428.4]
  assign _T_66249 = $signed(buffer_6_684) + $signed(buffer_6_685); // @[Modules.scala 71:109:@16430.4]
  assign _T_66250 = _T_66249[10:0]; // @[Modules.scala 71:109:@16431.4]
  assign buffer_6_734 = $signed(_T_66250); // @[Modules.scala 71:109:@16432.4]
  assign _T_66252 = $signed(buffer_6_686) + $signed(buffer_6_687); // @[Modules.scala 78:156:@16435.4]
  assign _T_66253 = _T_66252[10:0]; // @[Modules.scala 78:156:@16436.4]
  assign buffer_6_736 = $signed(_T_66253); // @[Modules.scala 78:156:@16437.4]
  assign _T_66255 = $signed(buffer_6_736) + $signed(buffer_6_688); // @[Modules.scala 78:156:@16439.4]
  assign _T_66256 = _T_66255[10:0]; // @[Modules.scala 78:156:@16440.4]
  assign buffer_6_737 = $signed(_T_66256); // @[Modules.scala 78:156:@16441.4]
  assign _T_66258 = $signed(buffer_6_737) + $signed(buffer_6_689); // @[Modules.scala 78:156:@16443.4]
  assign _T_66259 = _T_66258[10:0]; // @[Modules.scala 78:156:@16444.4]
  assign buffer_6_738 = $signed(_T_66259); // @[Modules.scala 78:156:@16445.4]
  assign _T_66261 = $signed(buffer_6_738) + $signed(buffer_0_701); // @[Modules.scala 78:156:@16447.4]
  assign _T_66262 = _T_66261[10:0]; // @[Modules.scala 78:156:@16448.4]
  assign buffer_6_739 = $signed(_T_66262); // @[Modules.scala 78:156:@16449.4]
  assign _T_66264 = $signed(buffer_6_739) + $signed(buffer_6_691); // @[Modules.scala 78:156:@16451.4]
  assign _T_66265 = _T_66264[10:0]; // @[Modules.scala 78:156:@16452.4]
  assign buffer_6_740 = $signed(_T_66265); // @[Modules.scala 78:156:@16453.4]
  assign _T_66267 = $signed(buffer_6_740) + $signed(buffer_6_692); // @[Modules.scala 78:156:@16455.4]
  assign _T_66268 = _T_66267[10:0]; // @[Modules.scala 78:156:@16456.4]
  assign buffer_6_741 = $signed(_T_66268); // @[Modules.scala 78:156:@16457.4]
  assign _T_66270 = $signed(buffer_6_741) + $signed(buffer_6_693); // @[Modules.scala 78:156:@16459.4]
  assign _T_66271 = _T_66270[10:0]; // @[Modules.scala 78:156:@16460.4]
  assign buffer_6_742 = $signed(_T_66271); // @[Modules.scala 78:156:@16461.4]
  assign _T_66273 = $signed(buffer_6_742) + $signed(buffer_6_694); // @[Modules.scala 78:156:@16463.4]
  assign _T_66274 = _T_66273[10:0]; // @[Modules.scala 78:156:@16464.4]
  assign buffer_6_743 = $signed(_T_66274); // @[Modules.scala 78:156:@16465.4]
  assign _T_66276 = $signed(buffer_6_743) + $signed(buffer_6_695); // @[Modules.scala 78:156:@16467.4]
  assign _T_66277 = _T_66276[10:0]; // @[Modules.scala 78:156:@16468.4]
  assign buffer_6_744 = $signed(_T_66277); // @[Modules.scala 78:156:@16469.4]
  assign _T_66279 = $signed(buffer_6_744) + $signed(buffer_6_696); // @[Modules.scala 78:156:@16471.4]
  assign _T_66280 = _T_66279[10:0]; // @[Modules.scala 78:156:@16472.4]
  assign buffer_6_745 = $signed(_T_66280); // @[Modules.scala 78:156:@16473.4]
  assign _T_66282 = $signed(buffer_6_745) + $signed(buffer_6_697); // @[Modules.scala 78:156:@16475.4]
  assign _T_66283 = _T_66282[10:0]; // @[Modules.scala 78:156:@16476.4]
  assign buffer_6_746 = $signed(_T_66283); // @[Modules.scala 78:156:@16477.4]
  assign _T_66285 = $signed(buffer_6_746) + $signed(buffer_6_698); // @[Modules.scala 78:156:@16479.4]
  assign _T_66286 = _T_66285[10:0]; // @[Modules.scala 78:156:@16480.4]
  assign buffer_6_747 = $signed(_T_66286); // @[Modules.scala 78:156:@16481.4]
  assign _T_66288 = $signed(buffer_6_747) + $signed(buffer_6_699); // @[Modules.scala 78:156:@16483.4]
  assign _T_66289 = _T_66288[10:0]; // @[Modules.scala 78:156:@16484.4]
  assign buffer_6_748 = $signed(_T_66289); // @[Modules.scala 78:156:@16485.4]
  assign _T_66291 = $signed(buffer_6_748) + $signed(buffer_6_700); // @[Modules.scala 78:156:@16487.4]
  assign _T_66292 = _T_66291[10:0]; // @[Modules.scala 78:156:@16488.4]
  assign buffer_6_749 = $signed(_T_66292); // @[Modules.scala 78:156:@16489.4]
  assign _T_66294 = $signed(buffer_6_749) + $signed(buffer_6_701); // @[Modules.scala 78:156:@16491.4]
  assign _T_66295 = _T_66294[10:0]; // @[Modules.scala 78:156:@16492.4]
  assign buffer_6_750 = $signed(_T_66295); // @[Modules.scala 78:156:@16493.4]
  assign _T_66297 = $signed(buffer_6_750) + $signed(buffer_6_702); // @[Modules.scala 78:156:@16495.4]
  assign _T_66298 = _T_66297[10:0]; // @[Modules.scala 78:156:@16496.4]
  assign buffer_6_751 = $signed(_T_66298); // @[Modules.scala 78:156:@16497.4]
  assign _T_66300 = $signed(buffer_6_751) + $signed(buffer_6_703); // @[Modules.scala 78:156:@16499.4]
  assign _T_66301 = _T_66300[10:0]; // @[Modules.scala 78:156:@16500.4]
  assign buffer_6_752 = $signed(_T_66301); // @[Modules.scala 78:156:@16501.4]
  assign _T_66303 = $signed(buffer_6_752) + $signed(buffer_6_704); // @[Modules.scala 78:156:@16503.4]
  assign _T_66304 = _T_66303[10:0]; // @[Modules.scala 78:156:@16504.4]
  assign buffer_6_753 = $signed(_T_66304); // @[Modules.scala 78:156:@16505.4]
  assign _T_66306 = $signed(buffer_6_753) + $signed(buffer_6_705); // @[Modules.scala 78:156:@16507.4]
  assign _T_66307 = _T_66306[10:0]; // @[Modules.scala 78:156:@16508.4]
  assign buffer_6_754 = $signed(_T_66307); // @[Modules.scala 78:156:@16509.4]
  assign _T_66309 = $signed(buffer_6_754) + $signed(buffer_6_706); // @[Modules.scala 78:156:@16511.4]
  assign _T_66310 = _T_66309[10:0]; // @[Modules.scala 78:156:@16512.4]
  assign buffer_6_755 = $signed(_T_66310); // @[Modules.scala 78:156:@16513.4]
  assign _T_66312 = $signed(buffer_6_755) + $signed(buffer_6_707); // @[Modules.scala 78:156:@16515.4]
  assign _T_66313 = _T_66312[10:0]; // @[Modules.scala 78:156:@16516.4]
  assign buffer_6_756 = $signed(_T_66313); // @[Modules.scala 78:156:@16517.4]
  assign _T_66315 = $signed(buffer_6_756) + $signed(buffer_6_708); // @[Modules.scala 78:156:@16519.4]
  assign _T_66316 = _T_66315[10:0]; // @[Modules.scala 78:156:@16520.4]
  assign buffer_6_757 = $signed(_T_66316); // @[Modules.scala 78:156:@16521.4]
  assign _T_66318 = $signed(buffer_6_757) + $signed(buffer_6_709); // @[Modules.scala 78:156:@16523.4]
  assign _T_66319 = _T_66318[10:0]; // @[Modules.scala 78:156:@16524.4]
  assign buffer_6_758 = $signed(_T_66319); // @[Modules.scala 78:156:@16525.4]
  assign _T_66321 = $signed(buffer_6_758) + $signed(buffer_6_710); // @[Modules.scala 78:156:@16527.4]
  assign _T_66322 = _T_66321[10:0]; // @[Modules.scala 78:156:@16528.4]
  assign buffer_6_759 = $signed(_T_66322); // @[Modules.scala 78:156:@16529.4]
  assign _T_66324 = $signed(buffer_6_759) + $signed(buffer_6_711); // @[Modules.scala 78:156:@16531.4]
  assign _T_66325 = _T_66324[10:0]; // @[Modules.scala 78:156:@16532.4]
  assign buffer_6_760 = $signed(_T_66325); // @[Modules.scala 78:156:@16533.4]
  assign _T_66327 = $signed(buffer_6_760) + $signed(buffer_6_712); // @[Modules.scala 78:156:@16535.4]
  assign _T_66328 = _T_66327[10:0]; // @[Modules.scala 78:156:@16536.4]
  assign buffer_6_761 = $signed(_T_66328); // @[Modules.scala 78:156:@16537.4]
  assign _T_66330 = $signed(buffer_6_761) + $signed(buffer_6_713); // @[Modules.scala 78:156:@16539.4]
  assign _T_66331 = _T_66330[10:0]; // @[Modules.scala 78:156:@16540.4]
  assign buffer_6_762 = $signed(_T_66331); // @[Modules.scala 78:156:@16541.4]
  assign _T_66333 = $signed(buffer_6_762) + $signed(buffer_6_714); // @[Modules.scala 78:156:@16543.4]
  assign _T_66334 = _T_66333[10:0]; // @[Modules.scala 78:156:@16544.4]
  assign buffer_6_763 = $signed(_T_66334); // @[Modules.scala 78:156:@16545.4]
  assign _T_66336 = $signed(buffer_6_763) + $signed(buffer_6_715); // @[Modules.scala 78:156:@16547.4]
  assign _T_66337 = _T_66336[10:0]; // @[Modules.scala 78:156:@16548.4]
  assign buffer_6_764 = $signed(_T_66337); // @[Modules.scala 78:156:@16549.4]
  assign _T_66339 = $signed(buffer_6_764) + $signed(buffer_6_716); // @[Modules.scala 78:156:@16551.4]
  assign _T_66340 = _T_66339[10:0]; // @[Modules.scala 78:156:@16552.4]
  assign buffer_6_765 = $signed(_T_66340); // @[Modules.scala 78:156:@16553.4]
  assign _T_66342 = $signed(buffer_6_765) + $signed(buffer_6_717); // @[Modules.scala 78:156:@16555.4]
  assign _T_66343 = _T_66342[10:0]; // @[Modules.scala 78:156:@16556.4]
  assign buffer_6_766 = $signed(_T_66343); // @[Modules.scala 78:156:@16557.4]
  assign _T_66345 = $signed(buffer_6_766) + $signed(buffer_6_718); // @[Modules.scala 78:156:@16559.4]
  assign _T_66346 = _T_66345[10:0]; // @[Modules.scala 78:156:@16560.4]
  assign buffer_6_767 = $signed(_T_66346); // @[Modules.scala 78:156:@16561.4]
  assign _T_66348 = $signed(buffer_6_767) + $signed(buffer_0_701); // @[Modules.scala 78:156:@16563.4]
  assign _T_66349 = _T_66348[10:0]; // @[Modules.scala 78:156:@16564.4]
  assign buffer_6_768 = $signed(_T_66349); // @[Modules.scala 78:156:@16565.4]
  assign _T_66351 = $signed(buffer_6_768) + $signed(buffer_6_720); // @[Modules.scala 78:156:@16567.4]
  assign _T_66352 = _T_66351[10:0]; // @[Modules.scala 78:156:@16568.4]
  assign buffer_6_769 = $signed(_T_66352); // @[Modules.scala 78:156:@16569.4]
  assign _T_66354 = $signed(buffer_6_769) + $signed(buffer_0_701); // @[Modules.scala 78:156:@16571.4]
  assign _T_66355 = _T_66354[10:0]; // @[Modules.scala 78:156:@16572.4]
  assign buffer_6_770 = $signed(_T_66355); // @[Modules.scala 78:156:@16573.4]
  assign _T_66357 = $signed(buffer_6_770) + $signed(buffer_6_722); // @[Modules.scala 78:156:@16575.4]
  assign _T_66358 = _T_66357[10:0]; // @[Modules.scala 78:156:@16576.4]
  assign buffer_6_771 = $signed(_T_66358); // @[Modules.scala 78:156:@16577.4]
  assign _T_66360 = $signed(buffer_6_771) + $signed(buffer_0_701); // @[Modules.scala 78:156:@16579.4]
  assign _T_66361 = _T_66360[10:0]; // @[Modules.scala 78:156:@16580.4]
  assign buffer_6_772 = $signed(_T_66361); // @[Modules.scala 78:156:@16581.4]
  assign _T_66363 = $signed(buffer_6_772) + $signed(buffer_6_724); // @[Modules.scala 78:156:@16583.4]
  assign _T_66364 = _T_66363[10:0]; // @[Modules.scala 78:156:@16584.4]
  assign buffer_6_773 = $signed(_T_66364); // @[Modules.scala 78:156:@16585.4]
  assign _T_66366 = $signed(buffer_6_773) + $signed(buffer_6_725); // @[Modules.scala 78:156:@16587.4]
  assign _T_66367 = _T_66366[10:0]; // @[Modules.scala 78:156:@16588.4]
  assign buffer_6_774 = $signed(_T_66367); // @[Modules.scala 78:156:@16589.4]
  assign _T_66369 = $signed(buffer_6_774) + $signed(buffer_6_726); // @[Modules.scala 78:156:@16591.4]
  assign _T_66370 = _T_66369[10:0]; // @[Modules.scala 78:156:@16592.4]
  assign buffer_6_775 = $signed(_T_66370); // @[Modules.scala 78:156:@16593.4]
  assign _T_66372 = $signed(buffer_6_775) + $signed(buffer_6_727); // @[Modules.scala 78:156:@16595.4]
  assign _T_66373 = _T_66372[10:0]; // @[Modules.scala 78:156:@16596.4]
  assign buffer_6_776 = $signed(_T_66373); // @[Modules.scala 78:156:@16597.4]
  assign _T_66375 = $signed(buffer_6_776) + $signed(buffer_6_728); // @[Modules.scala 78:156:@16599.4]
  assign _T_66376 = _T_66375[10:0]; // @[Modules.scala 78:156:@16600.4]
  assign buffer_6_777 = $signed(_T_66376); // @[Modules.scala 78:156:@16601.4]
  assign _T_66378 = $signed(buffer_6_777) + $signed(buffer_6_729); // @[Modules.scala 78:156:@16603.4]
  assign _T_66379 = _T_66378[10:0]; // @[Modules.scala 78:156:@16604.4]
  assign buffer_6_778 = $signed(_T_66379); // @[Modules.scala 78:156:@16605.4]
  assign _T_66381 = $signed(buffer_6_778) + $signed(buffer_6_730); // @[Modules.scala 78:156:@16607.4]
  assign _T_66382 = _T_66381[10:0]; // @[Modules.scala 78:156:@16608.4]
  assign buffer_6_779 = $signed(_T_66382); // @[Modules.scala 78:156:@16609.4]
  assign _T_66384 = $signed(buffer_6_779) + $signed(buffer_6_731); // @[Modules.scala 78:156:@16611.4]
  assign _T_66385 = _T_66384[10:0]; // @[Modules.scala 78:156:@16612.4]
  assign buffer_6_780 = $signed(_T_66385); // @[Modules.scala 78:156:@16613.4]
  assign _T_66387 = $signed(buffer_6_780) + $signed(buffer_6_732); // @[Modules.scala 78:156:@16615.4]
  assign _T_66388 = _T_66387[10:0]; // @[Modules.scala 78:156:@16616.4]
  assign buffer_6_781 = $signed(_T_66388); // @[Modules.scala 78:156:@16617.4]
  assign _T_66390 = $signed(buffer_6_781) + $signed(buffer_6_733); // @[Modules.scala 78:156:@16619.4]
  assign _T_66391 = _T_66390[10:0]; // @[Modules.scala 78:156:@16620.4]
  assign buffer_6_782 = $signed(_T_66391); // @[Modules.scala 78:156:@16621.4]
  assign _T_66393 = $signed(buffer_6_782) + $signed(buffer_6_734); // @[Modules.scala 78:156:@16623.4]
  assign _T_66394 = _T_66393[10:0]; // @[Modules.scala 78:156:@16624.4]
  assign buffer_6_783 = $signed(_T_66394); // @[Modules.scala 78:156:@16625.4]
  assign _T_66396 = $signed(io_in_0) + $signed(io_in_1); // @[Modules.scala 37:46:@16628.4]
  assign _T_66397 = _T_66396[4:0]; // @[Modules.scala 37:46:@16629.4]
  assign _T_66398 = $signed(_T_66397); // @[Modules.scala 37:46:@16630.4]
  assign _T_66427 = $signed(io_in_54) + $signed(io_in_55); // @[Modules.scala 37:46:@16679.4]
  assign _T_66428 = _T_66427[4:0]; // @[Modules.scala 37:46:@16680.4]
  assign _T_66429 = $signed(_T_66428); // @[Modules.scala 37:46:@16681.4]
  assign _T_66557 = $signed(io_in_216) + $signed(io_in_217); // @[Modules.scala 37:46:@16871.4]
  assign _T_66558 = _T_66557[4:0]; // @[Modules.scala 37:46:@16872.4]
  assign _T_66559 = $signed(_T_66558); // @[Modules.scala 37:46:@16873.4]
  assign _T_66599 = $signed(io_in_284) + $signed(io_in_285); // @[Modules.scala 37:46:@16932.4]
  assign _T_66600 = _T_66599[4:0]; // @[Modules.scala 37:46:@16933.4]
  assign _T_66601 = $signed(_T_66600); // @[Modules.scala 37:46:@16934.4]
  assign _T_66602 = $signed(io_in_286) + $signed(io_in_287); // @[Modules.scala 37:46:@16936.4]
  assign _T_66603 = _T_66602[4:0]; // @[Modules.scala 37:46:@16937.4]
  assign _T_66604 = $signed(_T_66603); // @[Modules.scala 37:46:@16938.4]
  assign _T_66618 = $signed(io_in_312) + $signed(io_in_313); // @[Modules.scala 37:46:@16958.4]
  assign _T_66619 = _T_66618[4:0]; // @[Modules.scala 37:46:@16959.4]
  assign _T_66620 = $signed(_T_66619); // @[Modules.scala 37:46:@16960.4]
  assign _T_66648 = $signed(io_in_364) + $signed(io_in_365); // @[Modules.scala 37:46:@17002.4]
  assign _T_66649 = _T_66648[4:0]; // @[Modules.scala 37:46:@17003.4]
  assign _T_66650 = $signed(_T_66649); // @[Modules.scala 37:46:@17004.4]
  assign _T_66927 = $signed(io_in_780) + $signed(io_in_781); // @[Modules.scala 37:46:@17405.4]
  assign _T_66928 = _T_66927[4:0]; // @[Modules.scala 37:46:@17406.4]
  assign _T_66929 = $signed(_T_66928); // @[Modules.scala 37:46:@17407.4]
  assign buffer_7_0 = {{6{_T_66398[4]}},_T_66398}; // @[Modules.scala 32:22:@8.4]
  assign _T_66930 = $signed(buffer_7_0) + $signed(11'sh0); // @[Modules.scala 65:57:@17410.4]
  assign _T_66931 = _T_66930[10:0]; // @[Modules.scala 65:57:@17411.4]
  assign buffer_7_392 = $signed(_T_66931); // @[Modules.scala 65:57:@17412.4]
  assign _T_66933 = $signed(buffer_2_2) + $signed(buffer_0_3); // @[Modules.scala 65:57:@17414.4]
  assign _T_66934 = _T_66933[10:0]; // @[Modules.scala 65:57:@17415.4]
  assign buffer_7_393 = $signed(_T_66934); // @[Modules.scala 65:57:@17416.4]
  assign buffer_7_8 = {{6{io_in_17[4]}},io_in_17}; // @[Modules.scala 32:22:@8.4]
  assign _T_66942 = $signed(buffer_7_8) + $signed(buffer_2_9); // @[Modules.scala 65:57:@17426.4]
  assign _T_66943 = _T_66942[10:0]; // @[Modules.scala 65:57:@17427.4]
  assign buffer_7_396 = $signed(_T_66943); // @[Modules.scala 65:57:@17428.4]
  assign _T_66945 = $signed(11'sh0) + $signed(buffer_0_11); // @[Modules.scala 65:57:@17430.4]
  assign _T_66946 = _T_66945[10:0]; // @[Modules.scala 65:57:@17431.4]
  assign buffer_7_397 = $signed(_T_66946); // @[Modules.scala 65:57:@17432.4]
  assign _T_66951 = $signed(buffer_1_14) + $signed(11'sh0); // @[Modules.scala 65:57:@17438.4]
  assign _T_66952 = _T_66951[10:0]; // @[Modules.scala 65:57:@17439.4]
  assign buffer_7_399 = $signed(_T_66952); // @[Modules.scala 65:57:@17440.4]
  assign buffer_7_17 = {{6{io_in_35[4]}},io_in_35}; // @[Modules.scala 32:22:@8.4]
  assign _T_66954 = $signed(buffer_5_16) + $signed(buffer_7_17); // @[Modules.scala 65:57:@17442.4]
  assign _T_66955 = _T_66954[10:0]; // @[Modules.scala 65:57:@17443.4]
  assign buffer_7_400 = $signed(_T_66955); // @[Modules.scala 65:57:@17444.4]
  assign buffer_7_27 = {{6{_T_66429[4]}},_T_66429}; // @[Modules.scala 32:22:@8.4]
  assign _T_66969 = $signed(buffer_3_26) + $signed(buffer_7_27); // @[Modules.scala 65:57:@17462.4]
  assign _T_66970 = _T_66969[10:0]; // @[Modules.scala 65:57:@17463.4]
  assign buffer_7_405 = $signed(_T_66970); // @[Modules.scala 65:57:@17464.4]
  assign _T_66975 = $signed(buffer_3_30) + $signed(buffer_1_31); // @[Modules.scala 65:57:@17470.4]
  assign _T_66976 = _T_66975[10:0]; // @[Modules.scala 65:57:@17471.4]
  assign buffer_7_407 = $signed(_T_66976); // @[Modules.scala 65:57:@17472.4]
  assign _T_67002 = $signed(11'sh0) + $signed(buffer_0_49); // @[Modules.scala 65:57:@17506.4]
  assign _T_67003 = _T_67002[10:0]; // @[Modules.scala 65:57:@17507.4]
  assign buffer_7_416 = $signed(_T_67003); // @[Modules.scala 65:57:@17508.4]
  assign _T_67017 = $signed(buffer_4_58) + $signed(buffer_0_59); // @[Modules.scala 65:57:@17526.4]
  assign _T_67018 = _T_67017[10:0]; // @[Modules.scala 65:57:@17527.4]
  assign buffer_7_421 = $signed(_T_67018); // @[Modules.scala 65:57:@17528.4]
  assign _T_67020 = $signed(buffer_3_60) + $signed(11'sh0); // @[Modules.scala 65:57:@17530.4]
  assign _T_67021 = _T_67020[10:0]; // @[Modules.scala 65:57:@17531.4]
  assign buffer_7_422 = $signed(_T_67021); // @[Modules.scala 65:57:@17532.4]
  assign buffer_7_63 = {{6{io_in_126[4]}},io_in_126}; // @[Modules.scala 32:22:@8.4]
  assign _T_67023 = $signed(11'sh0) + $signed(buffer_7_63); // @[Modules.scala 65:57:@17534.4]
  assign _T_67024 = _T_67023[10:0]; // @[Modules.scala 65:57:@17535.4]
  assign buffer_7_423 = $signed(_T_67024); // @[Modules.scala 65:57:@17536.4]
  assign _T_67029 = $signed(11'sh0) + $signed(buffer_0_67); // @[Modules.scala 65:57:@17542.4]
  assign _T_67030 = _T_67029[10:0]; // @[Modules.scala 65:57:@17543.4]
  assign buffer_7_425 = $signed(_T_67030); // @[Modules.scala 65:57:@17544.4]
  assign _T_67038 = $signed(11'sh0) + $signed(buffer_5_73); // @[Modules.scala 65:57:@17554.4]
  assign _T_67039 = _T_67038[10:0]; // @[Modules.scala 65:57:@17555.4]
  assign buffer_7_428 = $signed(_T_67039); // @[Modules.scala 65:57:@17556.4]
  assign _T_67041 = $signed(buffer_6_74) + $signed(buffer_1_75); // @[Modules.scala 65:57:@17558.4]
  assign _T_67042 = _T_67041[10:0]; // @[Modules.scala 65:57:@17559.4]
  assign buffer_7_429 = $signed(_T_67042); // @[Modules.scala 65:57:@17560.4]
  assign buffer_7_76 = {{6{io_in_152[4]}},io_in_152}; // @[Modules.scala 32:22:@8.4]
  assign _T_67044 = $signed(buffer_7_76) + $signed(buffer_3_77); // @[Modules.scala 65:57:@17562.4]
  assign _T_67045 = _T_67044[10:0]; // @[Modules.scala 65:57:@17563.4]
  assign buffer_7_430 = $signed(_T_67045); // @[Modules.scala 65:57:@17564.4]
  assign buffer_7_87 = {{6{io_in_175[4]}},io_in_175}; // @[Modules.scala 32:22:@8.4]
  assign _T_67059 = $signed(buffer_3_86) + $signed(buffer_7_87); // @[Modules.scala 65:57:@17582.4]
  assign _T_67060 = _T_67059[10:0]; // @[Modules.scala 65:57:@17583.4]
  assign buffer_7_435 = $signed(_T_67060); // @[Modules.scala 65:57:@17584.4]
  assign buffer_7_89 = {{6{io_in_179[4]}},io_in_179}; // @[Modules.scala 32:22:@8.4]
  assign _T_67062 = $signed(11'sh0) + $signed(buffer_7_89); // @[Modules.scala 65:57:@17586.4]
  assign _T_67063 = _T_67062[10:0]; // @[Modules.scala 65:57:@17587.4]
  assign buffer_7_436 = $signed(_T_67063); // @[Modules.scala 65:57:@17588.4]
  assign _T_67071 = $signed(buffer_6_94) + $signed(buffer_2_95); // @[Modules.scala 65:57:@17598.4]
  assign _T_67072 = _T_67071[10:0]; // @[Modules.scala 65:57:@17599.4]
  assign buffer_7_439 = $signed(_T_67072); // @[Modules.scala 65:57:@17600.4]
  assign buffer_7_108 = {{6{_T_66559[4]}},_T_66559}; // @[Modules.scala 32:22:@8.4]
  assign _T_67092 = $signed(buffer_7_108) + $signed(buffer_2_109); // @[Modules.scala 65:57:@17626.4]
  assign _T_67093 = _T_67092[10:0]; // @[Modules.scala 65:57:@17627.4]
  assign buffer_7_446 = $signed(_T_67093); // @[Modules.scala 65:57:@17628.4]
  assign _T_67101 = $signed(11'sh0) + $signed(buffer_3_115); // @[Modules.scala 65:57:@17638.4]
  assign _T_67102 = _T_67101[10:0]; // @[Modules.scala 65:57:@17639.4]
  assign buffer_7_449 = $signed(_T_67102); // @[Modules.scala 65:57:@17640.4]
  assign buffer_7_116 = {{6{io_in_233[4]}},io_in_233}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_117 = {{6{io_in_234[4]}},io_in_234}; // @[Modules.scala 32:22:@8.4]
  assign _T_67104 = $signed(buffer_7_116) + $signed(buffer_7_117); // @[Modules.scala 65:57:@17642.4]
  assign _T_67105 = _T_67104[10:0]; // @[Modules.scala 65:57:@17643.4]
  assign buffer_7_450 = $signed(_T_67105); // @[Modules.scala 65:57:@17644.4]
  assign _T_67113 = $signed(buffer_3_122) + $signed(buffer_1_123); // @[Modules.scala 65:57:@17654.4]
  assign _T_67114 = _T_67113[10:0]; // @[Modules.scala 65:57:@17655.4]
  assign buffer_7_453 = $signed(_T_67114); // @[Modules.scala 65:57:@17656.4]
  assign _T_67131 = $signed(11'sh0) + $signed(buffer_5_135); // @[Modules.scala 65:57:@17678.4]
  assign _T_67132 = _T_67131[10:0]; // @[Modules.scala 65:57:@17679.4]
  assign buffer_7_459 = $signed(_T_67132); // @[Modules.scala 65:57:@17680.4]
  assign buffer_7_136 = {{6{io_in_273[4]}},io_in_273}; // @[Modules.scala 32:22:@8.4]
  assign _T_67134 = $signed(buffer_7_136) + $signed(buffer_3_137); // @[Modules.scala 65:57:@17682.4]
  assign _T_67135 = _T_67134[10:0]; // @[Modules.scala 65:57:@17683.4]
  assign buffer_7_460 = $signed(_T_67135); // @[Modules.scala 65:57:@17684.4]
  assign buffer_7_142 = {{6{_T_66601[4]}},_T_66601}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_143 = {{6{_T_66604[4]}},_T_66604}; // @[Modules.scala 32:22:@8.4]
  assign _T_67143 = $signed(buffer_7_142) + $signed(buffer_7_143); // @[Modules.scala 65:57:@17694.4]
  assign _T_67144 = _T_67143[10:0]; // @[Modules.scala 65:57:@17695.4]
  assign buffer_7_463 = $signed(_T_67144); // @[Modules.scala 65:57:@17696.4]
  assign buffer_7_144 = {{6{io_in_288[4]}},io_in_288}; // @[Modules.scala 32:22:@8.4]
  assign _T_67146 = $signed(buffer_7_144) + $signed(buffer_6_145); // @[Modules.scala 65:57:@17698.4]
  assign _T_67147 = _T_67146[10:0]; // @[Modules.scala 65:57:@17699.4]
  assign buffer_7_464 = $signed(_T_67147); // @[Modules.scala 65:57:@17700.4]
  assign buffer_7_146 = {{6{io_in_292[4]}},io_in_292}; // @[Modules.scala 32:22:@8.4]
  assign _T_67149 = $signed(buffer_7_146) + $signed(11'sh0); // @[Modules.scala 65:57:@17702.4]
  assign _T_67150 = _T_67149[10:0]; // @[Modules.scala 65:57:@17703.4]
  assign buffer_7_465 = $signed(_T_67150); // @[Modules.scala 65:57:@17704.4]
  assign buffer_7_156 = {{6{_T_66620[4]}},_T_66620}; // @[Modules.scala 32:22:@8.4]
  assign _T_67164 = $signed(buffer_7_156) + $signed(buffer_0_157); // @[Modules.scala 65:57:@17722.4]
  assign _T_67165 = _T_67164[10:0]; // @[Modules.scala 65:57:@17723.4]
  assign buffer_7_470 = $signed(_T_67165); // @[Modules.scala 65:57:@17724.4]
  assign _T_67167 = $signed(buffer_6_158) + $signed(11'sh0); // @[Modules.scala 65:57:@17726.4]
  assign _T_67168 = _T_67167[10:0]; // @[Modules.scala 65:57:@17727.4]
  assign buffer_7_471 = $signed(_T_67168); // @[Modules.scala 65:57:@17728.4]
  assign _T_67197 = $signed(buffer_6_178) + $signed(11'sh0); // @[Modules.scala 65:57:@17766.4]
  assign _T_67198 = _T_67197[10:0]; // @[Modules.scala 65:57:@17767.4]
  assign buffer_7_481 = $signed(_T_67198); // @[Modules.scala 65:57:@17768.4]
  assign buffer_7_182 = {{6{_T_66650[4]}},_T_66650}; // @[Modules.scala 32:22:@8.4]
  assign _T_67203 = $signed(buffer_7_182) + $signed(buffer_5_183); // @[Modules.scala 65:57:@17774.4]
  assign _T_67204 = _T_67203[10:0]; // @[Modules.scala 65:57:@17775.4]
  assign buffer_7_483 = $signed(_T_67204); // @[Modules.scala 65:57:@17776.4]
  assign buffer_7_191 = {{6{io_in_383[4]}},io_in_383}; // @[Modules.scala 32:22:@8.4]
  assign _T_67215 = $signed(11'sh0) + $signed(buffer_7_191); // @[Modules.scala 65:57:@17790.4]
  assign _T_67216 = _T_67215[10:0]; // @[Modules.scala 65:57:@17791.4]
  assign buffer_7_487 = $signed(_T_67216); // @[Modules.scala 65:57:@17792.4]
  assign _T_67224 = $signed(buffer_4_196) + $signed(buffer_5_197); // @[Modules.scala 65:57:@17802.4]
  assign _T_67225 = _T_67224[10:0]; // @[Modules.scala 65:57:@17803.4]
  assign buffer_7_490 = $signed(_T_67225); // @[Modules.scala 65:57:@17804.4]
  assign buffer_7_198 = {{6{io_in_396[4]}},io_in_396}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_199 = {{6{io_in_398[4]}},io_in_398}; // @[Modules.scala 32:22:@8.4]
  assign _T_67227 = $signed(buffer_7_198) + $signed(buffer_7_199); // @[Modules.scala 65:57:@17806.4]
  assign _T_67228 = _T_67227[10:0]; // @[Modules.scala 65:57:@17807.4]
  assign buffer_7_491 = $signed(_T_67228); // @[Modules.scala 65:57:@17808.4]
  assign _T_67230 = $signed(11'sh0) + $signed(buffer_0_201); // @[Modules.scala 65:57:@17810.4]
  assign _T_67231 = _T_67230[10:0]; // @[Modules.scala 65:57:@17811.4]
  assign buffer_7_492 = $signed(_T_67231); // @[Modules.scala 65:57:@17812.4]
  assign _T_67236 = $signed(buffer_1_204) + $signed(buffer_3_205); // @[Modules.scala 65:57:@17818.4]
  assign _T_67237 = _T_67236[10:0]; // @[Modules.scala 65:57:@17819.4]
  assign buffer_7_494 = $signed(_T_67237); // @[Modules.scala 65:57:@17820.4]
  assign _T_67245 = $signed(buffer_3_210) + $signed(buffer_5_211); // @[Modules.scala 65:57:@17830.4]
  assign _T_67246 = _T_67245[10:0]; // @[Modules.scala 65:57:@17831.4]
  assign buffer_7_497 = $signed(_T_67246); // @[Modules.scala 65:57:@17832.4]
  assign _T_67248 = $signed(buffer_3_212) + $signed(buffer_0_213); // @[Modules.scala 65:57:@17834.4]
  assign _T_67249 = _T_67248[10:0]; // @[Modules.scala 65:57:@17835.4]
  assign buffer_7_498 = $signed(_T_67249); // @[Modules.scala 65:57:@17836.4]
  assign _T_67251 = $signed(buffer_0_214) + $signed(buffer_6_215); // @[Modules.scala 65:57:@17838.4]
  assign _T_67252 = _T_67251[10:0]; // @[Modules.scala 65:57:@17839.4]
  assign buffer_7_499 = $signed(_T_67252); // @[Modules.scala 65:57:@17840.4]
  assign _T_67257 = $signed(buffer_4_218) + $signed(buffer_0_219); // @[Modules.scala 65:57:@17846.4]
  assign _T_67258 = _T_67257[10:0]; // @[Modules.scala 65:57:@17847.4]
  assign buffer_7_501 = $signed(_T_67258); // @[Modules.scala 65:57:@17848.4]
  assign buffer_7_225 = {{6{io_in_451[4]}},io_in_451}; // @[Modules.scala 32:22:@8.4]
  assign _T_67266 = $signed(11'sh0) + $signed(buffer_7_225); // @[Modules.scala 65:57:@17858.4]
  assign _T_67267 = _T_67266[10:0]; // @[Modules.scala 65:57:@17859.4]
  assign buffer_7_504 = $signed(_T_67267); // @[Modules.scala 65:57:@17860.4]
  assign _T_67272 = $signed(11'sh0) + $signed(buffer_0_229); // @[Modules.scala 65:57:@17866.4]
  assign _T_67273 = _T_67272[10:0]; // @[Modules.scala 65:57:@17867.4]
  assign buffer_7_506 = $signed(_T_67273); // @[Modules.scala 65:57:@17868.4]
  assign buffer_7_234 = {{6{io_in_469[4]}},io_in_469}; // @[Modules.scala 32:22:@8.4]
  assign _T_67281 = $signed(buffer_7_234) + $signed(11'sh0); // @[Modules.scala 65:57:@17878.4]
  assign _T_67282 = _T_67281[10:0]; // @[Modules.scala 65:57:@17879.4]
  assign buffer_7_509 = $signed(_T_67282); // @[Modules.scala 65:57:@17880.4]
  assign buffer_7_240 = {{6{io_in_480[4]}},io_in_480}; // @[Modules.scala 32:22:@8.4]
  assign _T_67290 = $signed(buffer_7_240) + $signed(buffer_0_241); // @[Modules.scala 65:57:@17890.4]
  assign _T_67291 = _T_67290[10:0]; // @[Modules.scala 65:57:@17891.4]
  assign buffer_7_512 = $signed(_T_67291); // @[Modules.scala 65:57:@17892.4]
  assign _T_67299 = $signed(buffer_0_246) + $signed(11'sh0); // @[Modules.scala 65:57:@17902.4]
  assign _T_67300 = _T_67299[10:0]; // @[Modules.scala 65:57:@17903.4]
  assign buffer_7_515 = $signed(_T_67300); // @[Modules.scala 65:57:@17904.4]
  assign buffer_7_251 = {{6{io_in_502[4]}},io_in_502}; // @[Modules.scala 32:22:@8.4]
  assign _T_67305 = $signed(buffer_3_250) + $signed(buffer_7_251); // @[Modules.scala 65:57:@17910.4]
  assign _T_67306 = _T_67305[10:0]; // @[Modules.scala 65:57:@17911.4]
  assign buffer_7_517 = $signed(_T_67306); // @[Modules.scala 65:57:@17912.4]
  assign _T_67320 = $signed(11'sh0) + $signed(buffer_1_261); // @[Modules.scala 65:57:@17930.4]
  assign _T_67321 = _T_67320[10:0]; // @[Modules.scala 65:57:@17931.4]
  assign buffer_7_522 = $signed(_T_67321); // @[Modules.scala 65:57:@17932.4]
  assign buffer_7_262 = {{6{io_in_524[4]}},io_in_524}; // @[Modules.scala 32:22:@8.4]
  assign buffer_7_263 = {{6{io_in_527[4]}},io_in_527}; // @[Modules.scala 32:22:@8.4]
  assign _T_67323 = $signed(buffer_7_262) + $signed(buffer_7_263); // @[Modules.scala 65:57:@17934.4]
  assign _T_67324 = _T_67323[10:0]; // @[Modules.scala 65:57:@17935.4]
  assign buffer_7_523 = $signed(_T_67324); // @[Modules.scala 65:57:@17936.4]
  assign buffer_7_269 = {{6{io_in_538[4]}},io_in_538}; // @[Modules.scala 32:22:@8.4]
  assign _T_67332 = $signed(11'sh0) + $signed(buffer_7_269); // @[Modules.scala 65:57:@17946.4]
  assign _T_67333 = _T_67332[10:0]; // @[Modules.scala 65:57:@17947.4]
  assign buffer_7_526 = $signed(_T_67333); // @[Modules.scala 65:57:@17948.4]
  assign _T_67338 = $signed(buffer_1_272) + $signed(buffer_4_273); // @[Modules.scala 65:57:@17954.4]
  assign _T_67339 = _T_67338[10:0]; // @[Modules.scala 65:57:@17955.4]
  assign buffer_7_528 = $signed(_T_67339); // @[Modules.scala 65:57:@17956.4]
  assign _T_67341 = $signed(buffer_1_274) + $signed(buffer_0_275); // @[Modules.scala 65:57:@17958.4]
  assign _T_67342 = _T_67341[10:0]; // @[Modules.scala 65:57:@17959.4]
  assign buffer_7_529 = $signed(_T_67342); // @[Modules.scala 65:57:@17960.4]
  assign buffer_7_276 = {{6{io_in_553[4]}},io_in_553}; // @[Modules.scala 32:22:@8.4]
  assign _T_67344 = $signed(buffer_7_276) + $signed(buffer_3_277); // @[Modules.scala 65:57:@17962.4]
  assign _T_67345 = _T_67344[10:0]; // @[Modules.scala 65:57:@17963.4]
  assign buffer_7_530 = $signed(_T_67345); // @[Modules.scala 65:57:@17964.4]
  assign _T_67353 = $signed(11'sh0) + $signed(buffer_3_283); // @[Modules.scala 65:57:@17974.4]
  assign _T_67354 = _T_67353[10:0]; // @[Modules.scala 65:57:@17975.4]
  assign buffer_7_533 = $signed(_T_67354); // @[Modules.scala 65:57:@17976.4]
  assign buffer_7_293 = {{6{io_in_586[4]}},io_in_586}; // @[Modules.scala 32:22:@8.4]
  assign _T_67368 = $signed(buffer_4_292) + $signed(buffer_7_293); // @[Modules.scala 65:57:@17994.4]
  assign _T_67369 = _T_67368[10:0]; // @[Modules.scala 65:57:@17995.4]
  assign buffer_7_538 = $signed(_T_67369); // @[Modules.scala 65:57:@17996.4]
  assign buffer_7_299 = {{6{io_in_599[4]}},io_in_599}; // @[Modules.scala 32:22:@8.4]
  assign _T_67377 = $signed(buffer_2_298) + $signed(buffer_7_299); // @[Modules.scala 65:57:@18006.4]
  assign _T_67378 = _T_67377[10:0]; // @[Modules.scala 65:57:@18007.4]
  assign buffer_7_541 = $signed(_T_67378); // @[Modules.scala 65:57:@18008.4]
  assign buffer_7_301 = {{6{io_in_603[4]}},io_in_603}; // @[Modules.scala 32:22:@8.4]
  assign _T_67380 = $signed(buffer_2_300) + $signed(buffer_7_301); // @[Modules.scala 65:57:@18010.4]
  assign _T_67381 = _T_67380[10:0]; // @[Modules.scala 65:57:@18011.4]
  assign buffer_7_542 = $signed(_T_67381); // @[Modules.scala 65:57:@18012.4]
  assign _T_67389 = $signed(buffer_4_306) + $signed(11'sh0); // @[Modules.scala 65:57:@18022.4]
  assign _T_67390 = _T_67389[10:0]; // @[Modules.scala 65:57:@18023.4]
  assign buffer_7_545 = $signed(_T_67390); // @[Modules.scala 65:57:@18024.4]
  assign buffer_7_311 = {{6{io_in_622[4]}},io_in_622}; // @[Modules.scala 32:22:@8.4]
  assign _T_67395 = $signed(buffer_3_310) + $signed(buffer_7_311); // @[Modules.scala 65:57:@18030.4]
  assign _T_67396 = _T_67395[10:0]; // @[Modules.scala 65:57:@18031.4]
  assign buffer_7_547 = $signed(_T_67396); // @[Modules.scala 65:57:@18032.4]
  assign _T_67398 = $signed(buffer_6_312) + $signed(buffer_3_313); // @[Modules.scala 65:57:@18034.4]
  assign _T_67399 = _T_67398[10:0]; // @[Modules.scala 65:57:@18035.4]
  assign buffer_7_548 = $signed(_T_67399); // @[Modules.scala 65:57:@18036.4]
  assign _T_67404 = $signed(11'sh0) + $signed(buffer_2_317); // @[Modules.scala 65:57:@18042.4]
  assign _T_67405 = _T_67404[10:0]; // @[Modules.scala 65:57:@18043.4]
  assign buffer_7_550 = $signed(_T_67405); // @[Modules.scala 65:57:@18044.4]
  assign _T_67413 = $signed(buffer_2_322) + $signed(11'sh0); // @[Modules.scala 65:57:@18054.4]
  assign _T_67414 = _T_67413[10:0]; // @[Modules.scala 65:57:@18055.4]
  assign buffer_7_553 = $signed(_T_67414); // @[Modules.scala 65:57:@18056.4]
  assign _T_67422 = $signed(11'sh0) + $signed(buffer_5_329); // @[Modules.scala 65:57:@18066.4]
  assign _T_67423 = _T_67422[10:0]; // @[Modules.scala 65:57:@18067.4]
  assign buffer_7_556 = $signed(_T_67423); // @[Modules.scala 65:57:@18068.4]
  assign _T_67428 = $signed(buffer_0_332) + $signed(buffer_3_333); // @[Modules.scala 65:57:@18074.4]
  assign _T_67429 = _T_67428[10:0]; // @[Modules.scala 65:57:@18075.4]
  assign buffer_7_558 = $signed(_T_67429); // @[Modules.scala 65:57:@18076.4]
  assign _T_67431 = $signed(buffer_0_334) + $signed(buffer_2_335); // @[Modules.scala 65:57:@18078.4]
  assign _T_67432 = _T_67431[10:0]; // @[Modules.scala 65:57:@18079.4]
  assign buffer_7_559 = $signed(_T_67432); // @[Modules.scala 65:57:@18080.4]
  assign _T_67434 = $signed(buffer_4_336) + $signed(buffer_0_337); // @[Modules.scala 65:57:@18082.4]
  assign _T_67435 = _T_67434[10:0]; // @[Modules.scala 65:57:@18083.4]
  assign buffer_7_560 = $signed(_T_67435); // @[Modules.scala 65:57:@18084.4]
  assign _T_67443 = $signed(buffer_2_342) + $signed(buffer_3_343); // @[Modules.scala 65:57:@18094.4]
  assign _T_67444 = _T_67443[10:0]; // @[Modules.scala 65:57:@18095.4]
  assign buffer_7_563 = $signed(_T_67444); // @[Modules.scala 65:57:@18096.4]
  assign buffer_7_345 = {{6{io_in_691[4]}},io_in_691}; // @[Modules.scala 32:22:@8.4]
  assign _T_67446 = $signed(11'sh0) + $signed(buffer_7_345); // @[Modules.scala 65:57:@18098.4]
  assign _T_67447 = _T_67446[10:0]; // @[Modules.scala 65:57:@18099.4]
  assign buffer_7_564 = $signed(_T_67447); // @[Modules.scala 65:57:@18100.4]
  assign _T_67452 = $signed(buffer_4_348) + $signed(11'sh0); // @[Modules.scala 65:57:@18106.4]
  assign _T_67453 = _T_67452[10:0]; // @[Modules.scala 65:57:@18107.4]
  assign buffer_7_566 = $signed(_T_67453); // @[Modules.scala 65:57:@18108.4]
  assign _T_67473 = $signed(11'sh0) + $signed(buffer_1_363); // @[Modules.scala 65:57:@18134.4]
  assign _T_67474 = _T_67473[10:0]; // @[Modules.scala 65:57:@18135.4]
  assign buffer_7_573 = $signed(_T_67474); // @[Modules.scala 65:57:@18136.4]
  assign _T_67494 = $signed(buffer_4_376) + $signed(buffer_0_377); // @[Modules.scala 65:57:@18162.4]
  assign _T_67495 = _T_67494[10:0]; // @[Modules.scala 65:57:@18163.4]
  assign buffer_7_580 = $signed(_T_67495); // @[Modules.scala 65:57:@18164.4]
  assign buffer_7_380 = {{6{io_in_761[4]}},io_in_761}; // @[Modules.scala 32:22:@8.4]
  assign _T_67500 = $signed(buffer_7_380) + $signed(11'sh0); // @[Modules.scala 65:57:@18170.4]
  assign _T_67501 = _T_67500[10:0]; // @[Modules.scala 65:57:@18171.4]
  assign buffer_7_582 = $signed(_T_67501); // @[Modules.scala 65:57:@18172.4]
  assign buffer_7_390 = {{6{_T_66929[4]}},_T_66929}; // @[Modules.scala 32:22:@8.4]
  assign _T_67515 = $signed(buffer_7_390) + $signed(buffer_2_391); // @[Modules.scala 65:57:@18190.4]
  assign _T_67516 = _T_67515[10:0]; // @[Modules.scala 65:57:@18191.4]
  assign buffer_7_587 = $signed(_T_67516); // @[Modules.scala 65:57:@18192.4]
  assign _T_67518 = $signed(buffer_7_392) + $signed(buffer_7_393); // @[Modules.scala 68:83:@18194.4]
  assign _T_67519 = _T_67518[10:0]; // @[Modules.scala 68:83:@18195.4]
  assign buffer_7_588 = $signed(_T_67519); // @[Modules.scala 68:83:@18196.4]
  assign _T_67524 = $signed(buffer_7_396) + $signed(buffer_7_397); // @[Modules.scala 68:83:@18202.4]
  assign _T_67525 = _T_67524[10:0]; // @[Modules.scala 68:83:@18203.4]
  assign buffer_7_590 = $signed(_T_67525); // @[Modules.scala 68:83:@18204.4]
  assign _T_67527 = $signed(buffer_2_398) + $signed(buffer_7_399); // @[Modules.scala 68:83:@18206.4]
  assign _T_67528 = _T_67527[10:0]; // @[Modules.scala 68:83:@18207.4]
  assign buffer_7_591 = $signed(_T_67528); // @[Modules.scala 68:83:@18208.4]
  assign _T_67530 = $signed(buffer_7_400) + $signed(buffer_1_401); // @[Modules.scala 68:83:@18210.4]
  assign _T_67531 = _T_67530[10:0]; // @[Modules.scala 68:83:@18211.4]
  assign buffer_7_592 = $signed(_T_67531); // @[Modules.scala 68:83:@18212.4]
  assign _T_67533 = $signed(buffer_2_402) + $signed(buffer_4_403); // @[Modules.scala 68:83:@18214.4]
  assign _T_67534 = _T_67533[10:0]; // @[Modules.scala 68:83:@18215.4]
  assign buffer_7_593 = $signed(_T_67534); // @[Modules.scala 68:83:@18216.4]
  assign _T_67536 = $signed(buffer_1_404) + $signed(buffer_7_405); // @[Modules.scala 68:83:@18218.4]
  assign _T_67537 = _T_67536[10:0]; // @[Modules.scala 68:83:@18219.4]
  assign buffer_7_594 = $signed(_T_67537); // @[Modules.scala 68:83:@18220.4]
  assign _T_67539 = $signed(buffer_0_406) + $signed(buffer_7_407); // @[Modules.scala 68:83:@18222.4]
  assign _T_67540 = _T_67539[10:0]; // @[Modules.scala 68:83:@18223.4]
  assign buffer_7_595 = $signed(_T_67540); // @[Modules.scala 68:83:@18224.4]
  assign _T_67548 = $signed(buffer_3_412) + $signed(buffer_1_413); // @[Modules.scala 68:83:@18234.4]
  assign _T_67549 = _T_67548[10:0]; // @[Modules.scala 68:83:@18235.4]
  assign buffer_7_598 = $signed(_T_67549); // @[Modules.scala 68:83:@18236.4]
  assign _T_67551 = $signed(buffer_2_414) + $signed(buffer_1_415); // @[Modules.scala 68:83:@18238.4]
  assign _T_67552 = _T_67551[10:0]; // @[Modules.scala 68:83:@18239.4]
  assign buffer_7_599 = $signed(_T_67552); // @[Modules.scala 68:83:@18240.4]
  assign _T_67554 = $signed(buffer_7_416) + $signed(buffer_2_417); // @[Modules.scala 68:83:@18242.4]
  assign _T_67555 = _T_67554[10:0]; // @[Modules.scala 68:83:@18243.4]
  assign buffer_7_600 = $signed(_T_67555); // @[Modules.scala 68:83:@18244.4]
  assign _T_67557 = $signed(buffer_0_418) + $signed(buffer_6_419); // @[Modules.scala 68:83:@18246.4]
  assign _T_67558 = _T_67557[10:0]; // @[Modules.scala 68:83:@18247.4]
  assign buffer_7_601 = $signed(_T_67558); // @[Modules.scala 68:83:@18248.4]
  assign _T_67560 = $signed(buffer_0_420) + $signed(buffer_7_421); // @[Modules.scala 68:83:@18250.4]
  assign _T_67561 = _T_67560[10:0]; // @[Modules.scala 68:83:@18251.4]
  assign buffer_7_602 = $signed(_T_67561); // @[Modules.scala 68:83:@18252.4]
  assign _T_67563 = $signed(buffer_7_422) + $signed(buffer_7_423); // @[Modules.scala 68:83:@18254.4]
  assign _T_67564 = _T_67563[10:0]; // @[Modules.scala 68:83:@18255.4]
  assign buffer_7_603 = $signed(_T_67564); // @[Modules.scala 68:83:@18256.4]
  assign _T_67566 = $signed(buffer_4_424) + $signed(buffer_7_425); // @[Modules.scala 68:83:@18258.4]
  assign _T_67567 = _T_67566[10:0]; // @[Modules.scala 68:83:@18259.4]
  assign buffer_7_604 = $signed(_T_67567); // @[Modules.scala 68:83:@18260.4]
  assign _T_67569 = $signed(buffer_4_426) + $signed(buffer_2_427); // @[Modules.scala 68:83:@18262.4]
  assign _T_67570 = _T_67569[10:0]; // @[Modules.scala 68:83:@18263.4]
  assign buffer_7_605 = $signed(_T_67570); // @[Modules.scala 68:83:@18264.4]
  assign _T_67572 = $signed(buffer_7_428) + $signed(buffer_7_429); // @[Modules.scala 68:83:@18266.4]
  assign _T_67573 = _T_67572[10:0]; // @[Modules.scala 68:83:@18267.4]
  assign buffer_7_606 = $signed(_T_67573); // @[Modules.scala 68:83:@18268.4]
  assign _T_67575 = $signed(buffer_7_430) + $signed(buffer_4_431); // @[Modules.scala 68:83:@18270.4]
  assign _T_67576 = _T_67575[10:0]; // @[Modules.scala 68:83:@18271.4]
  assign buffer_7_607 = $signed(_T_67576); // @[Modules.scala 68:83:@18272.4]
  assign _T_67581 = $signed(buffer_2_434) + $signed(buffer_7_435); // @[Modules.scala 68:83:@18278.4]
  assign _T_67582 = _T_67581[10:0]; // @[Modules.scala 68:83:@18279.4]
  assign buffer_7_609 = $signed(_T_67582); // @[Modules.scala 68:83:@18280.4]
  assign _T_67584 = $signed(buffer_7_436) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18282.4]
  assign _T_67585 = _T_67584[10:0]; // @[Modules.scala 68:83:@18283.4]
  assign buffer_7_610 = $signed(_T_67585); // @[Modules.scala 68:83:@18284.4]
  assign _T_67587 = $signed(buffer_0_395) + $signed(buffer_7_439); // @[Modules.scala 68:83:@18286.4]
  assign _T_67588 = _T_67587[10:0]; // @[Modules.scala 68:83:@18287.4]
  assign buffer_7_611 = $signed(_T_67588); // @[Modules.scala 68:83:@18288.4]
  assign _T_67590 = $signed(buffer_2_440) + $signed(buffer_0_441); // @[Modules.scala 68:83:@18290.4]
  assign _T_67591 = _T_67590[10:0]; // @[Modules.scala 68:83:@18291.4]
  assign buffer_7_612 = $signed(_T_67591); // @[Modules.scala 68:83:@18292.4]
  assign _T_67593 = $signed(buffer_1_442) + $signed(buffer_5_443); // @[Modules.scala 68:83:@18294.4]
  assign _T_67594 = _T_67593[10:0]; // @[Modules.scala 68:83:@18295.4]
  assign buffer_7_613 = $signed(_T_67594); // @[Modules.scala 68:83:@18296.4]
  assign _T_67599 = $signed(buffer_7_446) + $signed(buffer_2_447); // @[Modules.scala 68:83:@18302.4]
  assign _T_67600 = _T_67599[10:0]; // @[Modules.scala 68:83:@18303.4]
  assign buffer_7_615 = $signed(_T_67600); // @[Modules.scala 68:83:@18304.4]
  assign _T_67602 = $signed(buffer_0_395) + $signed(buffer_7_449); // @[Modules.scala 68:83:@18306.4]
  assign _T_67603 = _T_67602[10:0]; // @[Modules.scala 68:83:@18307.4]
  assign buffer_7_616 = $signed(_T_67603); // @[Modules.scala 68:83:@18308.4]
  assign _T_67605 = $signed(buffer_7_450) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18310.4]
  assign _T_67606 = _T_67605[10:0]; // @[Modules.scala 68:83:@18311.4]
  assign buffer_7_617 = $signed(_T_67606); // @[Modules.scala 68:83:@18312.4]
  assign _T_67608 = $signed(buffer_4_452) + $signed(buffer_7_453); // @[Modules.scala 68:83:@18314.4]
  assign _T_67609 = _T_67608[10:0]; // @[Modules.scala 68:83:@18315.4]
  assign buffer_7_618 = $signed(_T_67609); // @[Modules.scala 68:83:@18316.4]
  assign _T_67617 = $signed(buffer_0_395) + $signed(buffer_7_459); // @[Modules.scala 68:83:@18326.4]
  assign _T_67618 = _T_67617[10:0]; // @[Modules.scala 68:83:@18327.4]
  assign buffer_7_621 = $signed(_T_67618); // @[Modules.scala 68:83:@18328.4]
  assign _T_67620 = $signed(buffer_7_460) + $signed(buffer_1_461); // @[Modules.scala 68:83:@18330.4]
  assign _T_67621 = _T_67620[10:0]; // @[Modules.scala 68:83:@18331.4]
  assign buffer_7_622 = $signed(_T_67621); // @[Modules.scala 68:83:@18332.4]
  assign _T_67623 = $signed(buffer_0_395) + $signed(buffer_7_463); // @[Modules.scala 68:83:@18334.4]
  assign _T_67624 = _T_67623[10:0]; // @[Modules.scala 68:83:@18335.4]
  assign buffer_7_623 = $signed(_T_67624); // @[Modules.scala 68:83:@18336.4]
  assign _T_67626 = $signed(buffer_7_464) + $signed(buffer_7_465); // @[Modules.scala 68:83:@18338.4]
  assign _T_67627 = _T_67626[10:0]; // @[Modules.scala 68:83:@18339.4]
  assign buffer_7_624 = $signed(_T_67627); // @[Modules.scala 68:83:@18340.4]
  assign _T_67635 = $signed(buffer_7_470) + $signed(buffer_7_471); // @[Modules.scala 68:83:@18350.4]
  assign _T_67636 = _T_67635[10:0]; // @[Modules.scala 68:83:@18351.4]
  assign buffer_7_627 = $signed(_T_67636); // @[Modules.scala 68:83:@18352.4]
  assign _T_67644 = $signed(buffer_0_395) + $signed(buffer_6_477); // @[Modules.scala 68:83:@18362.4]
  assign _T_67645 = _T_67644[10:0]; // @[Modules.scala 68:83:@18363.4]
  assign buffer_7_630 = $signed(_T_67645); // @[Modules.scala 68:83:@18364.4]
  assign _T_67650 = $signed(buffer_0_395) + $signed(buffer_7_481); // @[Modules.scala 68:83:@18370.4]
  assign _T_67651 = _T_67650[10:0]; // @[Modules.scala 68:83:@18371.4]
  assign buffer_7_632 = $signed(_T_67651); // @[Modules.scala 68:83:@18372.4]
  assign _T_67653 = $signed(buffer_2_482) + $signed(buffer_7_483); // @[Modules.scala 68:83:@18374.4]
  assign _T_67654 = _T_67653[10:0]; // @[Modules.scala 68:83:@18375.4]
  assign buffer_7_633 = $signed(_T_67654); // @[Modules.scala 68:83:@18376.4]
  assign _T_67659 = $signed(buffer_0_486) + $signed(buffer_7_487); // @[Modules.scala 68:83:@18382.4]
  assign _T_67660 = _T_67659[10:0]; // @[Modules.scala 68:83:@18383.4]
  assign buffer_7_635 = $signed(_T_67660); // @[Modules.scala 68:83:@18384.4]
  assign _T_67665 = $signed(buffer_7_490) + $signed(buffer_7_491); // @[Modules.scala 68:83:@18390.4]
  assign _T_67666 = _T_67665[10:0]; // @[Modules.scala 68:83:@18391.4]
  assign buffer_7_637 = $signed(_T_67666); // @[Modules.scala 68:83:@18392.4]
  assign _T_67668 = $signed(buffer_7_492) + $signed(buffer_0_493); // @[Modules.scala 68:83:@18394.4]
  assign _T_67669 = _T_67668[10:0]; // @[Modules.scala 68:83:@18395.4]
  assign buffer_7_638 = $signed(_T_67669); // @[Modules.scala 68:83:@18396.4]
  assign _T_67671 = $signed(buffer_7_494) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18398.4]
  assign _T_67672 = _T_67671[10:0]; // @[Modules.scala 68:83:@18399.4]
  assign buffer_7_639 = $signed(_T_67672); // @[Modules.scala 68:83:@18400.4]
  assign _T_67674 = $signed(buffer_5_496) + $signed(buffer_7_497); // @[Modules.scala 68:83:@18402.4]
  assign _T_67675 = _T_67674[10:0]; // @[Modules.scala 68:83:@18403.4]
  assign buffer_7_640 = $signed(_T_67675); // @[Modules.scala 68:83:@18404.4]
  assign _T_67677 = $signed(buffer_7_498) + $signed(buffer_7_499); // @[Modules.scala 68:83:@18406.4]
  assign _T_67678 = _T_67677[10:0]; // @[Modules.scala 68:83:@18407.4]
  assign buffer_7_641 = $signed(_T_67678); // @[Modules.scala 68:83:@18408.4]
  assign _T_67680 = $signed(buffer_0_500) + $signed(buffer_7_501); // @[Modules.scala 68:83:@18410.4]
  assign _T_67681 = _T_67680[10:0]; // @[Modules.scala 68:83:@18411.4]
  assign buffer_7_642 = $signed(_T_67681); // @[Modules.scala 68:83:@18412.4]
  assign _T_67683 = $signed(buffer_3_502) + $signed(buffer_5_503); // @[Modules.scala 68:83:@18414.4]
  assign _T_67684 = _T_67683[10:0]; // @[Modules.scala 68:83:@18415.4]
  assign buffer_7_643 = $signed(_T_67684); // @[Modules.scala 68:83:@18416.4]
  assign _T_67686 = $signed(buffer_7_504) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18418.4]
  assign _T_67687 = _T_67686[10:0]; // @[Modules.scala 68:83:@18419.4]
  assign buffer_7_644 = $signed(_T_67687); // @[Modules.scala 68:83:@18420.4]
  assign _T_67689 = $signed(buffer_7_506) + $signed(buffer_2_507); // @[Modules.scala 68:83:@18422.4]
  assign _T_67690 = _T_67689[10:0]; // @[Modules.scala 68:83:@18423.4]
  assign buffer_7_645 = $signed(_T_67690); // @[Modules.scala 68:83:@18424.4]
  assign _T_67692 = $signed(buffer_5_508) + $signed(buffer_7_509); // @[Modules.scala 68:83:@18426.4]
  assign _T_67693 = _T_67692[10:0]; // @[Modules.scala 68:83:@18427.4]
  assign buffer_7_646 = $signed(_T_67693); // @[Modules.scala 68:83:@18428.4]
  assign _T_67695 = $signed(buffer_3_510) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18430.4]
  assign _T_67696 = _T_67695[10:0]; // @[Modules.scala 68:83:@18431.4]
  assign buffer_7_647 = $signed(_T_67696); // @[Modules.scala 68:83:@18432.4]
  assign _T_67698 = $signed(buffer_7_512) + $signed(buffer_2_513); // @[Modules.scala 68:83:@18434.4]
  assign _T_67699 = _T_67698[10:0]; // @[Modules.scala 68:83:@18435.4]
  assign buffer_7_648 = $signed(_T_67699); // @[Modules.scala 68:83:@18436.4]
  assign _T_67701 = $signed(buffer_2_514) + $signed(buffer_7_515); // @[Modules.scala 68:83:@18438.4]
  assign _T_67702 = _T_67701[10:0]; // @[Modules.scala 68:83:@18439.4]
  assign buffer_7_649 = $signed(_T_67702); // @[Modules.scala 68:83:@18440.4]
  assign _T_67704 = $signed(buffer_0_395) + $signed(buffer_7_517); // @[Modules.scala 68:83:@18442.4]
  assign _T_67705 = _T_67704[10:0]; // @[Modules.scala 68:83:@18443.4]
  assign buffer_7_650 = $signed(_T_67705); // @[Modules.scala 68:83:@18444.4]
  assign _T_67707 = $signed(buffer_0_395) + $signed(buffer_3_519); // @[Modules.scala 68:83:@18446.4]
  assign _T_67708 = _T_67707[10:0]; // @[Modules.scala 68:83:@18447.4]
  assign buffer_7_651 = $signed(_T_67708); // @[Modules.scala 68:83:@18448.4]
  assign _T_67710 = $signed(buffer_0_520) + $signed(buffer_5_521); // @[Modules.scala 68:83:@18450.4]
  assign _T_67711 = _T_67710[10:0]; // @[Modules.scala 68:83:@18451.4]
  assign buffer_7_652 = $signed(_T_67711); // @[Modules.scala 68:83:@18452.4]
  assign _T_67713 = $signed(buffer_7_522) + $signed(buffer_7_523); // @[Modules.scala 68:83:@18454.4]
  assign _T_67714 = _T_67713[10:0]; // @[Modules.scala 68:83:@18455.4]
  assign buffer_7_653 = $signed(_T_67714); // @[Modules.scala 68:83:@18456.4]
  assign _T_67716 = $signed(buffer_3_524) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18458.4]
  assign _T_67717 = _T_67716[10:0]; // @[Modules.scala 68:83:@18459.4]
  assign buffer_7_654 = $signed(_T_67717); // @[Modules.scala 68:83:@18460.4]
  assign _T_67719 = $signed(buffer_7_526) + $signed(buffer_1_527); // @[Modules.scala 68:83:@18462.4]
  assign _T_67720 = _T_67719[10:0]; // @[Modules.scala 68:83:@18463.4]
  assign buffer_7_655 = $signed(_T_67720); // @[Modules.scala 68:83:@18464.4]
  assign _T_67722 = $signed(buffer_7_528) + $signed(buffer_7_529); // @[Modules.scala 68:83:@18466.4]
  assign _T_67723 = _T_67722[10:0]; // @[Modules.scala 68:83:@18467.4]
  assign buffer_7_656 = $signed(_T_67723); // @[Modules.scala 68:83:@18468.4]
  assign _T_67725 = $signed(buffer_7_530) + $signed(buffer_5_531); // @[Modules.scala 68:83:@18470.4]
  assign _T_67726 = _T_67725[10:0]; // @[Modules.scala 68:83:@18471.4]
  assign buffer_7_657 = $signed(_T_67726); // @[Modules.scala 68:83:@18472.4]
  assign _T_67728 = $signed(buffer_2_532) + $signed(buffer_7_533); // @[Modules.scala 68:83:@18474.4]
  assign _T_67729 = _T_67728[10:0]; // @[Modules.scala 68:83:@18475.4]
  assign buffer_7_658 = $signed(_T_67729); // @[Modules.scala 68:83:@18476.4]
  assign _T_67734 = $signed(buffer_2_536) + $signed(buffer_3_537); // @[Modules.scala 68:83:@18482.4]
  assign _T_67735 = _T_67734[10:0]; // @[Modules.scala 68:83:@18483.4]
  assign buffer_7_660 = $signed(_T_67735); // @[Modules.scala 68:83:@18484.4]
  assign _T_67737 = $signed(buffer_7_538) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18486.4]
  assign _T_67738 = _T_67737[10:0]; // @[Modules.scala 68:83:@18487.4]
  assign buffer_7_661 = $signed(_T_67738); // @[Modules.scala 68:83:@18488.4]
  assign _T_67740 = $signed(buffer_2_540) + $signed(buffer_7_541); // @[Modules.scala 68:83:@18490.4]
  assign _T_67741 = _T_67740[10:0]; // @[Modules.scala 68:83:@18491.4]
  assign buffer_7_662 = $signed(_T_67741); // @[Modules.scala 68:83:@18492.4]
  assign _T_67743 = $signed(buffer_7_542) + $signed(buffer_3_543); // @[Modules.scala 68:83:@18494.4]
  assign _T_67744 = _T_67743[10:0]; // @[Modules.scala 68:83:@18495.4]
  assign buffer_7_663 = $signed(_T_67744); // @[Modules.scala 68:83:@18496.4]
  assign _T_67746 = $signed(buffer_3_544) + $signed(buffer_7_545); // @[Modules.scala 68:83:@18498.4]
  assign _T_67747 = _T_67746[10:0]; // @[Modules.scala 68:83:@18499.4]
  assign buffer_7_664 = $signed(_T_67747); // @[Modules.scala 68:83:@18500.4]
  assign _T_67749 = $signed(buffer_0_395) + $signed(buffer_7_547); // @[Modules.scala 68:83:@18502.4]
  assign _T_67750 = _T_67749[10:0]; // @[Modules.scala 68:83:@18503.4]
  assign buffer_7_665 = $signed(_T_67750); // @[Modules.scala 68:83:@18504.4]
  assign _T_67752 = $signed(buffer_7_548) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18506.4]
  assign _T_67753 = _T_67752[10:0]; // @[Modules.scala 68:83:@18507.4]
  assign buffer_7_666 = $signed(_T_67753); // @[Modules.scala 68:83:@18508.4]
  assign _T_67755 = $signed(buffer_7_550) + $signed(buffer_3_551); // @[Modules.scala 68:83:@18510.4]
  assign _T_67756 = _T_67755[10:0]; // @[Modules.scala 68:83:@18511.4]
  assign buffer_7_667 = $signed(_T_67756); // @[Modules.scala 68:83:@18512.4]
  assign _T_67758 = $signed(buffer_3_552) + $signed(buffer_7_553); // @[Modules.scala 68:83:@18514.4]
  assign _T_67759 = _T_67758[10:0]; // @[Modules.scala 68:83:@18515.4]
  assign buffer_7_668 = $signed(_T_67759); // @[Modules.scala 68:83:@18516.4]
  assign _T_67761 = $signed(buffer_0_395) + $signed(buffer_5_555); // @[Modules.scala 68:83:@18518.4]
  assign _T_67762 = _T_67761[10:0]; // @[Modules.scala 68:83:@18519.4]
  assign buffer_7_669 = $signed(_T_67762); // @[Modules.scala 68:83:@18520.4]
  assign _T_67764 = $signed(buffer_7_556) + $signed(buffer_4_557); // @[Modules.scala 68:83:@18522.4]
  assign _T_67765 = _T_67764[10:0]; // @[Modules.scala 68:83:@18523.4]
  assign buffer_7_670 = $signed(_T_67765); // @[Modules.scala 68:83:@18524.4]
  assign _T_67767 = $signed(buffer_7_558) + $signed(buffer_7_559); // @[Modules.scala 68:83:@18526.4]
  assign _T_67768 = _T_67767[10:0]; // @[Modules.scala 68:83:@18527.4]
  assign buffer_7_671 = $signed(_T_67768); // @[Modules.scala 68:83:@18528.4]
  assign _T_67770 = $signed(buffer_7_560) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18530.4]
  assign _T_67771 = _T_67770[10:0]; // @[Modules.scala 68:83:@18531.4]
  assign buffer_7_672 = $signed(_T_67771); // @[Modules.scala 68:83:@18532.4]
  assign _T_67773 = $signed(buffer_0_395) + $signed(buffer_7_563); // @[Modules.scala 68:83:@18534.4]
  assign _T_67774 = _T_67773[10:0]; // @[Modules.scala 68:83:@18535.4]
  assign buffer_7_673 = $signed(_T_67774); // @[Modules.scala 68:83:@18536.4]
  assign _T_67776 = $signed(buffer_7_564) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18538.4]
  assign _T_67777 = _T_67776[10:0]; // @[Modules.scala 68:83:@18539.4]
  assign buffer_7_674 = $signed(_T_67777); // @[Modules.scala 68:83:@18540.4]
  assign _T_67779 = $signed(buffer_7_566) + $signed(buffer_0_395); // @[Modules.scala 68:83:@18542.4]
  assign _T_67780 = _T_67779[10:0]; // @[Modules.scala 68:83:@18543.4]
  assign buffer_7_675 = $signed(_T_67780); // @[Modules.scala 68:83:@18544.4]
  assign _T_67788 = $signed(buffer_0_395) + $signed(buffer_7_573); // @[Modules.scala 68:83:@18554.4]
  assign _T_67789 = _T_67788[10:0]; // @[Modules.scala 68:83:@18555.4]
  assign buffer_7_678 = $signed(_T_67789); // @[Modules.scala 68:83:@18556.4]
  assign _T_67800 = $signed(buffer_7_580) + $signed(buffer_1_581); // @[Modules.scala 68:83:@18570.4]
  assign _T_67801 = _T_67800[10:0]; // @[Modules.scala 68:83:@18571.4]
  assign buffer_7_682 = $signed(_T_67801); // @[Modules.scala 68:83:@18572.4]
  assign _T_67803 = $signed(buffer_7_582) + $signed(buffer_4_583); // @[Modules.scala 68:83:@18574.4]
  assign _T_67804 = _T_67803[10:0]; // @[Modules.scala 68:83:@18575.4]
  assign buffer_7_683 = $signed(_T_67804); // @[Modules.scala 68:83:@18576.4]
  assign _T_67809 = $signed(buffer_0_395) + $signed(buffer_7_587); // @[Modules.scala 68:83:@18582.4]
  assign _T_67810 = _T_67809[10:0]; // @[Modules.scala 68:83:@18583.4]
  assign buffer_7_685 = $signed(_T_67810); // @[Modules.scala 68:83:@18584.4]
  assign _T_67812 = $signed(buffer_7_588) + $signed(buffer_2_589); // @[Modules.scala 71:109:@18586.4]
  assign _T_67813 = _T_67812[10:0]; // @[Modules.scala 71:109:@18587.4]
  assign buffer_7_686 = $signed(_T_67813); // @[Modules.scala 71:109:@18588.4]
  assign _T_67815 = $signed(buffer_7_590) + $signed(buffer_7_591); // @[Modules.scala 71:109:@18590.4]
  assign _T_67816 = _T_67815[10:0]; // @[Modules.scala 71:109:@18591.4]
  assign buffer_7_687 = $signed(_T_67816); // @[Modules.scala 71:109:@18592.4]
  assign _T_67818 = $signed(buffer_7_592) + $signed(buffer_7_593); // @[Modules.scala 71:109:@18594.4]
  assign _T_67819 = _T_67818[10:0]; // @[Modules.scala 71:109:@18595.4]
  assign buffer_7_688 = $signed(_T_67819); // @[Modules.scala 71:109:@18596.4]
  assign _T_67821 = $signed(buffer_7_594) + $signed(buffer_7_595); // @[Modules.scala 71:109:@18598.4]
  assign _T_67822 = _T_67821[10:0]; // @[Modules.scala 71:109:@18599.4]
  assign buffer_7_689 = $signed(_T_67822); // @[Modules.scala 71:109:@18600.4]
  assign _T_67827 = $signed(buffer_7_598) + $signed(buffer_7_599); // @[Modules.scala 71:109:@18606.4]
  assign _T_67828 = _T_67827[10:0]; // @[Modules.scala 71:109:@18607.4]
  assign buffer_7_691 = $signed(_T_67828); // @[Modules.scala 71:109:@18608.4]
  assign _T_67830 = $signed(buffer_7_600) + $signed(buffer_7_601); // @[Modules.scala 71:109:@18610.4]
  assign _T_67831 = _T_67830[10:0]; // @[Modules.scala 71:109:@18611.4]
  assign buffer_7_692 = $signed(_T_67831); // @[Modules.scala 71:109:@18612.4]
  assign _T_67833 = $signed(buffer_7_602) + $signed(buffer_7_603); // @[Modules.scala 71:109:@18614.4]
  assign _T_67834 = _T_67833[10:0]; // @[Modules.scala 71:109:@18615.4]
  assign buffer_7_693 = $signed(_T_67834); // @[Modules.scala 71:109:@18616.4]
  assign _T_67836 = $signed(buffer_7_604) + $signed(buffer_7_605); // @[Modules.scala 71:109:@18618.4]
  assign _T_67837 = _T_67836[10:0]; // @[Modules.scala 71:109:@18619.4]
  assign buffer_7_694 = $signed(_T_67837); // @[Modules.scala 71:109:@18620.4]
  assign _T_67839 = $signed(buffer_7_606) + $signed(buffer_7_607); // @[Modules.scala 71:109:@18622.4]
  assign _T_67840 = _T_67839[10:0]; // @[Modules.scala 71:109:@18623.4]
  assign buffer_7_695 = $signed(_T_67840); // @[Modules.scala 71:109:@18624.4]
  assign _T_67842 = $signed(buffer_2_608) + $signed(buffer_7_609); // @[Modules.scala 71:109:@18626.4]
  assign _T_67843 = _T_67842[10:0]; // @[Modules.scala 71:109:@18627.4]
  assign buffer_7_696 = $signed(_T_67843); // @[Modules.scala 71:109:@18628.4]
  assign _T_67845 = $signed(buffer_7_610) + $signed(buffer_7_611); // @[Modules.scala 71:109:@18630.4]
  assign _T_67846 = _T_67845[10:0]; // @[Modules.scala 71:109:@18631.4]
  assign buffer_7_697 = $signed(_T_67846); // @[Modules.scala 71:109:@18632.4]
  assign _T_67848 = $signed(buffer_7_612) + $signed(buffer_7_613); // @[Modules.scala 71:109:@18634.4]
  assign _T_67849 = _T_67848[10:0]; // @[Modules.scala 71:109:@18635.4]
  assign buffer_7_698 = $signed(_T_67849); // @[Modules.scala 71:109:@18636.4]
  assign _T_67851 = $signed(buffer_0_593) + $signed(buffer_7_615); // @[Modules.scala 71:109:@18638.4]
  assign _T_67852 = _T_67851[10:0]; // @[Modules.scala 71:109:@18639.4]
  assign buffer_7_699 = $signed(_T_67852); // @[Modules.scala 71:109:@18640.4]
  assign _T_67854 = $signed(buffer_7_616) + $signed(buffer_7_617); // @[Modules.scala 71:109:@18642.4]
  assign _T_67855 = _T_67854[10:0]; // @[Modules.scala 71:109:@18643.4]
  assign buffer_7_700 = $signed(_T_67855); // @[Modules.scala 71:109:@18644.4]
  assign _T_67857 = $signed(buffer_7_618) + $signed(buffer_2_619); // @[Modules.scala 71:109:@18646.4]
  assign _T_67858 = _T_67857[10:0]; // @[Modules.scala 71:109:@18647.4]
  assign buffer_7_701 = $signed(_T_67858); // @[Modules.scala 71:109:@18648.4]
  assign _T_67860 = $signed(buffer_2_620) + $signed(buffer_7_621); // @[Modules.scala 71:109:@18650.4]
  assign _T_67861 = _T_67860[10:0]; // @[Modules.scala 71:109:@18651.4]
  assign buffer_7_702 = $signed(_T_67861); // @[Modules.scala 71:109:@18652.4]
  assign _T_67863 = $signed(buffer_7_622) + $signed(buffer_7_623); // @[Modules.scala 71:109:@18654.4]
  assign _T_67864 = _T_67863[10:0]; // @[Modules.scala 71:109:@18655.4]
  assign buffer_7_703 = $signed(_T_67864); // @[Modules.scala 71:109:@18656.4]
  assign _T_67866 = $signed(buffer_7_624) + $signed(buffer_0_593); // @[Modules.scala 71:109:@18658.4]
  assign _T_67867 = _T_67866[10:0]; // @[Modules.scala 71:109:@18659.4]
  assign buffer_7_704 = $signed(_T_67867); // @[Modules.scala 71:109:@18660.4]
  assign _T_67869 = $signed(buffer_1_626) + $signed(buffer_7_627); // @[Modules.scala 71:109:@18662.4]
  assign _T_67870 = _T_67869[10:0]; // @[Modules.scala 71:109:@18663.4]
  assign buffer_7_705 = $signed(_T_67870); // @[Modules.scala 71:109:@18664.4]
  assign _T_67872 = $signed(buffer_4_628) + $signed(buffer_2_629); // @[Modules.scala 71:109:@18666.4]
  assign _T_67873 = _T_67872[10:0]; // @[Modules.scala 71:109:@18667.4]
  assign buffer_7_706 = $signed(_T_67873); // @[Modules.scala 71:109:@18668.4]
  assign _T_67875 = $signed(buffer_7_630) + $signed(buffer_1_631); // @[Modules.scala 71:109:@18670.4]
  assign _T_67876 = _T_67875[10:0]; // @[Modules.scala 71:109:@18671.4]
  assign buffer_7_707 = $signed(_T_67876); // @[Modules.scala 71:109:@18672.4]
  assign _T_67878 = $signed(buffer_7_632) + $signed(buffer_7_633); // @[Modules.scala 71:109:@18674.4]
  assign _T_67879 = _T_67878[10:0]; // @[Modules.scala 71:109:@18675.4]
  assign buffer_7_708 = $signed(_T_67879); // @[Modules.scala 71:109:@18676.4]
  assign _T_67881 = $signed(buffer_4_634) + $signed(buffer_7_635); // @[Modules.scala 71:109:@18678.4]
  assign _T_67882 = _T_67881[10:0]; // @[Modules.scala 71:109:@18679.4]
  assign buffer_7_709 = $signed(_T_67882); // @[Modules.scala 71:109:@18680.4]
  assign _T_67884 = $signed(buffer_3_636) + $signed(buffer_7_637); // @[Modules.scala 71:109:@18682.4]
  assign _T_67885 = _T_67884[10:0]; // @[Modules.scala 71:109:@18683.4]
  assign buffer_7_710 = $signed(_T_67885); // @[Modules.scala 71:109:@18684.4]
  assign _T_67887 = $signed(buffer_7_638) + $signed(buffer_7_639); // @[Modules.scala 71:109:@18686.4]
  assign _T_67888 = _T_67887[10:0]; // @[Modules.scala 71:109:@18687.4]
  assign buffer_7_711 = $signed(_T_67888); // @[Modules.scala 71:109:@18688.4]
  assign _T_67890 = $signed(buffer_7_640) + $signed(buffer_7_641); // @[Modules.scala 71:109:@18690.4]
  assign _T_67891 = _T_67890[10:0]; // @[Modules.scala 71:109:@18691.4]
  assign buffer_7_712 = $signed(_T_67891); // @[Modules.scala 71:109:@18692.4]
  assign _T_67893 = $signed(buffer_7_642) + $signed(buffer_7_643); // @[Modules.scala 71:109:@18694.4]
  assign _T_67894 = _T_67893[10:0]; // @[Modules.scala 71:109:@18695.4]
  assign buffer_7_713 = $signed(_T_67894); // @[Modules.scala 71:109:@18696.4]
  assign _T_67896 = $signed(buffer_7_644) + $signed(buffer_7_645); // @[Modules.scala 71:109:@18698.4]
  assign _T_67897 = _T_67896[10:0]; // @[Modules.scala 71:109:@18699.4]
  assign buffer_7_714 = $signed(_T_67897); // @[Modules.scala 71:109:@18700.4]
  assign _T_67899 = $signed(buffer_7_646) + $signed(buffer_7_647); // @[Modules.scala 71:109:@18702.4]
  assign _T_67900 = _T_67899[10:0]; // @[Modules.scala 71:109:@18703.4]
  assign buffer_7_715 = $signed(_T_67900); // @[Modules.scala 71:109:@18704.4]
  assign _T_67902 = $signed(buffer_7_648) + $signed(buffer_7_649); // @[Modules.scala 71:109:@18706.4]
  assign _T_67903 = _T_67902[10:0]; // @[Modules.scala 71:109:@18707.4]
  assign buffer_7_716 = $signed(_T_67903); // @[Modules.scala 71:109:@18708.4]
  assign _T_67905 = $signed(buffer_7_650) + $signed(buffer_7_651); // @[Modules.scala 71:109:@18710.4]
  assign _T_67906 = _T_67905[10:0]; // @[Modules.scala 71:109:@18711.4]
  assign buffer_7_717 = $signed(_T_67906); // @[Modules.scala 71:109:@18712.4]
  assign _T_67908 = $signed(buffer_7_652) + $signed(buffer_7_653); // @[Modules.scala 71:109:@18714.4]
  assign _T_67909 = _T_67908[10:0]; // @[Modules.scala 71:109:@18715.4]
  assign buffer_7_718 = $signed(_T_67909); // @[Modules.scala 71:109:@18716.4]
  assign _T_67911 = $signed(buffer_7_654) + $signed(buffer_7_655); // @[Modules.scala 71:109:@18718.4]
  assign _T_67912 = _T_67911[10:0]; // @[Modules.scala 71:109:@18719.4]
  assign buffer_7_719 = $signed(_T_67912); // @[Modules.scala 71:109:@18720.4]
  assign _T_67914 = $signed(buffer_7_656) + $signed(buffer_7_657); // @[Modules.scala 71:109:@18722.4]
  assign _T_67915 = _T_67914[10:0]; // @[Modules.scala 71:109:@18723.4]
  assign buffer_7_720 = $signed(_T_67915); // @[Modules.scala 71:109:@18724.4]
  assign _T_67917 = $signed(buffer_7_658) + $signed(buffer_3_659); // @[Modules.scala 71:109:@18726.4]
  assign _T_67918 = _T_67917[10:0]; // @[Modules.scala 71:109:@18727.4]
  assign buffer_7_721 = $signed(_T_67918); // @[Modules.scala 71:109:@18728.4]
  assign _T_67920 = $signed(buffer_7_660) + $signed(buffer_7_661); // @[Modules.scala 71:109:@18730.4]
  assign _T_67921 = _T_67920[10:0]; // @[Modules.scala 71:109:@18731.4]
  assign buffer_7_722 = $signed(_T_67921); // @[Modules.scala 71:109:@18732.4]
  assign _T_67923 = $signed(buffer_7_662) + $signed(buffer_7_663); // @[Modules.scala 71:109:@18734.4]
  assign _T_67924 = _T_67923[10:0]; // @[Modules.scala 71:109:@18735.4]
  assign buffer_7_723 = $signed(_T_67924); // @[Modules.scala 71:109:@18736.4]
  assign _T_67926 = $signed(buffer_7_664) + $signed(buffer_7_665); // @[Modules.scala 71:109:@18738.4]
  assign _T_67927 = _T_67926[10:0]; // @[Modules.scala 71:109:@18739.4]
  assign buffer_7_724 = $signed(_T_67927); // @[Modules.scala 71:109:@18740.4]
  assign _T_67929 = $signed(buffer_7_666) + $signed(buffer_7_667); // @[Modules.scala 71:109:@18742.4]
  assign _T_67930 = _T_67929[10:0]; // @[Modules.scala 71:109:@18743.4]
  assign buffer_7_725 = $signed(_T_67930); // @[Modules.scala 71:109:@18744.4]
  assign _T_67932 = $signed(buffer_7_668) + $signed(buffer_7_669); // @[Modules.scala 71:109:@18746.4]
  assign _T_67933 = _T_67932[10:0]; // @[Modules.scala 71:109:@18747.4]
  assign buffer_7_726 = $signed(_T_67933); // @[Modules.scala 71:109:@18748.4]
  assign _T_67935 = $signed(buffer_7_670) + $signed(buffer_7_671); // @[Modules.scala 71:109:@18750.4]
  assign _T_67936 = _T_67935[10:0]; // @[Modules.scala 71:109:@18751.4]
  assign buffer_7_727 = $signed(_T_67936); // @[Modules.scala 71:109:@18752.4]
  assign _T_67938 = $signed(buffer_7_672) + $signed(buffer_7_673); // @[Modules.scala 71:109:@18754.4]
  assign _T_67939 = _T_67938[10:0]; // @[Modules.scala 71:109:@18755.4]
  assign buffer_7_728 = $signed(_T_67939); // @[Modules.scala 71:109:@18756.4]
  assign _T_67941 = $signed(buffer_7_674) + $signed(buffer_7_675); // @[Modules.scala 71:109:@18758.4]
  assign _T_67942 = _T_67941[10:0]; // @[Modules.scala 71:109:@18759.4]
  assign buffer_7_729 = $signed(_T_67942); // @[Modules.scala 71:109:@18760.4]
  assign _T_67947 = $signed(buffer_7_678) + $signed(buffer_0_593); // @[Modules.scala 71:109:@18766.4]
  assign _T_67948 = _T_67947[10:0]; // @[Modules.scala 71:109:@18767.4]
  assign buffer_7_731 = $signed(_T_67948); // @[Modules.scala 71:109:@18768.4]
  assign _T_67953 = $signed(buffer_7_682) + $signed(buffer_7_683); // @[Modules.scala 71:109:@18774.4]
  assign _T_67954 = _T_67953[10:0]; // @[Modules.scala 71:109:@18775.4]
  assign buffer_7_733 = $signed(_T_67954); // @[Modules.scala 71:109:@18776.4]
  assign _T_67956 = $signed(buffer_0_593) + $signed(buffer_7_685); // @[Modules.scala 71:109:@18778.4]
  assign _T_67957 = _T_67956[10:0]; // @[Modules.scala 71:109:@18779.4]
  assign buffer_7_734 = $signed(_T_67957); // @[Modules.scala 71:109:@18780.4]
  assign _T_67959 = $signed(buffer_7_686) + $signed(buffer_7_687); // @[Modules.scala 78:156:@18783.4]
  assign _T_67960 = _T_67959[10:0]; // @[Modules.scala 78:156:@18784.4]
  assign buffer_7_736 = $signed(_T_67960); // @[Modules.scala 78:156:@18785.4]
  assign _T_67962 = $signed(buffer_7_736) + $signed(buffer_7_688); // @[Modules.scala 78:156:@18787.4]
  assign _T_67963 = _T_67962[10:0]; // @[Modules.scala 78:156:@18788.4]
  assign buffer_7_737 = $signed(_T_67963); // @[Modules.scala 78:156:@18789.4]
  assign _T_67965 = $signed(buffer_7_737) + $signed(buffer_7_689); // @[Modules.scala 78:156:@18791.4]
  assign _T_67966 = _T_67965[10:0]; // @[Modules.scala 78:156:@18792.4]
  assign buffer_7_738 = $signed(_T_67966); // @[Modules.scala 78:156:@18793.4]
  assign _T_67968 = $signed(buffer_7_738) + $signed(buffer_1_690); // @[Modules.scala 78:156:@18795.4]
  assign _T_67969 = _T_67968[10:0]; // @[Modules.scala 78:156:@18796.4]
  assign buffer_7_739 = $signed(_T_67969); // @[Modules.scala 78:156:@18797.4]
  assign _T_67971 = $signed(buffer_7_739) + $signed(buffer_7_691); // @[Modules.scala 78:156:@18799.4]
  assign _T_67972 = _T_67971[10:0]; // @[Modules.scala 78:156:@18800.4]
  assign buffer_7_740 = $signed(_T_67972); // @[Modules.scala 78:156:@18801.4]
  assign _T_67974 = $signed(buffer_7_740) + $signed(buffer_7_692); // @[Modules.scala 78:156:@18803.4]
  assign _T_67975 = _T_67974[10:0]; // @[Modules.scala 78:156:@18804.4]
  assign buffer_7_741 = $signed(_T_67975); // @[Modules.scala 78:156:@18805.4]
  assign _T_67977 = $signed(buffer_7_741) + $signed(buffer_7_693); // @[Modules.scala 78:156:@18807.4]
  assign _T_67978 = _T_67977[10:0]; // @[Modules.scala 78:156:@18808.4]
  assign buffer_7_742 = $signed(_T_67978); // @[Modules.scala 78:156:@18809.4]
  assign _T_67980 = $signed(buffer_7_742) + $signed(buffer_7_694); // @[Modules.scala 78:156:@18811.4]
  assign _T_67981 = _T_67980[10:0]; // @[Modules.scala 78:156:@18812.4]
  assign buffer_7_743 = $signed(_T_67981); // @[Modules.scala 78:156:@18813.4]
  assign _T_67983 = $signed(buffer_7_743) + $signed(buffer_7_695); // @[Modules.scala 78:156:@18815.4]
  assign _T_67984 = _T_67983[10:0]; // @[Modules.scala 78:156:@18816.4]
  assign buffer_7_744 = $signed(_T_67984); // @[Modules.scala 78:156:@18817.4]
  assign _T_67986 = $signed(buffer_7_744) + $signed(buffer_7_696); // @[Modules.scala 78:156:@18819.4]
  assign _T_67987 = _T_67986[10:0]; // @[Modules.scala 78:156:@18820.4]
  assign buffer_7_745 = $signed(_T_67987); // @[Modules.scala 78:156:@18821.4]
  assign _T_67989 = $signed(buffer_7_745) + $signed(buffer_7_697); // @[Modules.scala 78:156:@18823.4]
  assign _T_67990 = _T_67989[10:0]; // @[Modules.scala 78:156:@18824.4]
  assign buffer_7_746 = $signed(_T_67990); // @[Modules.scala 78:156:@18825.4]
  assign _T_67992 = $signed(buffer_7_746) + $signed(buffer_7_698); // @[Modules.scala 78:156:@18827.4]
  assign _T_67993 = _T_67992[10:0]; // @[Modules.scala 78:156:@18828.4]
  assign buffer_7_747 = $signed(_T_67993); // @[Modules.scala 78:156:@18829.4]
  assign _T_67995 = $signed(buffer_7_747) + $signed(buffer_7_699); // @[Modules.scala 78:156:@18831.4]
  assign _T_67996 = _T_67995[10:0]; // @[Modules.scala 78:156:@18832.4]
  assign buffer_7_748 = $signed(_T_67996); // @[Modules.scala 78:156:@18833.4]
  assign _T_67998 = $signed(buffer_7_748) + $signed(buffer_7_700); // @[Modules.scala 78:156:@18835.4]
  assign _T_67999 = _T_67998[10:0]; // @[Modules.scala 78:156:@18836.4]
  assign buffer_7_749 = $signed(_T_67999); // @[Modules.scala 78:156:@18837.4]
  assign _T_68001 = $signed(buffer_7_749) + $signed(buffer_7_701); // @[Modules.scala 78:156:@18839.4]
  assign _T_68002 = _T_68001[10:0]; // @[Modules.scala 78:156:@18840.4]
  assign buffer_7_750 = $signed(_T_68002); // @[Modules.scala 78:156:@18841.4]
  assign _T_68004 = $signed(buffer_7_750) + $signed(buffer_7_702); // @[Modules.scala 78:156:@18843.4]
  assign _T_68005 = _T_68004[10:0]; // @[Modules.scala 78:156:@18844.4]
  assign buffer_7_751 = $signed(_T_68005); // @[Modules.scala 78:156:@18845.4]
  assign _T_68007 = $signed(buffer_7_751) + $signed(buffer_7_703); // @[Modules.scala 78:156:@18847.4]
  assign _T_68008 = _T_68007[10:0]; // @[Modules.scala 78:156:@18848.4]
  assign buffer_7_752 = $signed(_T_68008); // @[Modules.scala 78:156:@18849.4]
  assign _T_68010 = $signed(buffer_7_752) + $signed(buffer_7_704); // @[Modules.scala 78:156:@18851.4]
  assign _T_68011 = _T_68010[10:0]; // @[Modules.scala 78:156:@18852.4]
  assign buffer_7_753 = $signed(_T_68011); // @[Modules.scala 78:156:@18853.4]
  assign _T_68013 = $signed(buffer_7_753) + $signed(buffer_7_705); // @[Modules.scala 78:156:@18855.4]
  assign _T_68014 = _T_68013[10:0]; // @[Modules.scala 78:156:@18856.4]
  assign buffer_7_754 = $signed(_T_68014); // @[Modules.scala 78:156:@18857.4]
  assign _T_68016 = $signed(buffer_7_754) + $signed(buffer_7_706); // @[Modules.scala 78:156:@18859.4]
  assign _T_68017 = _T_68016[10:0]; // @[Modules.scala 78:156:@18860.4]
  assign buffer_7_755 = $signed(_T_68017); // @[Modules.scala 78:156:@18861.4]
  assign _T_68019 = $signed(buffer_7_755) + $signed(buffer_7_707); // @[Modules.scala 78:156:@18863.4]
  assign _T_68020 = _T_68019[10:0]; // @[Modules.scala 78:156:@18864.4]
  assign buffer_7_756 = $signed(_T_68020); // @[Modules.scala 78:156:@18865.4]
  assign _T_68022 = $signed(buffer_7_756) + $signed(buffer_7_708); // @[Modules.scala 78:156:@18867.4]
  assign _T_68023 = _T_68022[10:0]; // @[Modules.scala 78:156:@18868.4]
  assign buffer_7_757 = $signed(_T_68023); // @[Modules.scala 78:156:@18869.4]
  assign _T_68025 = $signed(buffer_7_757) + $signed(buffer_7_709); // @[Modules.scala 78:156:@18871.4]
  assign _T_68026 = _T_68025[10:0]; // @[Modules.scala 78:156:@18872.4]
  assign buffer_7_758 = $signed(_T_68026); // @[Modules.scala 78:156:@18873.4]
  assign _T_68028 = $signed(buffer_7_758) + $signed(buffer_7_710); // @[Modules.scala 78:156:@18875.4]
  assign _T_68029 = _T_68028[10:0]; // @[Modules.scala 78:156:@18876.4]
  assign buffer_7_759 = $signed(_T_68029); // @[Modules.scala 78:156:@18877.4]
  assign _T_68031 = $signed(buffer_7_759) + $signed(buffer_7_711); // @[Modules.scala 78:156:@18879.4]
  assign _T_68032 = _T_68031[10:0]; // @[Modules.scala 78:156:@18880.4]
  assign buffer_7_760 = $signed(_T_68032); // @[Modules.scala 78:156:@18881.4]
  assign _T_68034 = $signed(buffer_7_760) + $signed(buffer_7_712); // @[Modules.scala 78:156:@18883.4]
  assign _T_68035 = _T_68034[10:0]; // @[Modules.scala 78:156:@18884.4]
  assign buffer_7_761 = $signed(_T_68035); // @[Modules.scala 78:156:@18885.4]
  assign _T_68037 = $signed(buffer_7_761) + $signed(buffer_7_713); // @[Modules.scala 78:156:@18887.4]
  assign _T_68038 = _T_68037[10:0]; // @[Modules.scala 78:156:@18888.4]
  assign buffer_7_762 = $signed(_T_68038); // @[Modules.scala 78:156:@18889.4]
  assign _T_68040 = $signed(buffer_7_762) + $signed(buffer_7_714); // @[Modules.scala 78:156:@18891.4]
  assign _T_68041 = _T_68040[10:0]; // @[Modules.scala 78:156:@18892.4]
  assign buffer_7_763 = $signed(_T_68041); // @[Modules.scala 78:156:@18893.4]
  assign _T_68043 = $signed(buffer_7_763) + $signed(buffer_7_715); // @[Modules.scala 78:156:@18895.4]
  assign _T_68044 = _T_68043[10:0]; // @[Modules.scala 78:156:@18896.4]
  assign buffer_7_764 = $signed(_T_68044); // @[Modules.scala 78:156:@18897.4]
  assign _T_68046 = $signed(buffer_7_764) + $signed(buffer_7_716); // @[Modules.scala 78:156:@18899.4]
  assign _T_68047 = _T_68046[10:0]; // @[Modules.scala 78:156:@18900.4]
  assign buffer_7_765 = $signed(_T_68047); // @[Modules.scala 78:156:@18901.4]
  assign _T_68049 = $signed(buffer_7_765) + $signed(buffer_7_717); // @[Modules.scala 78:156:@18903.4]
  assign _T_68050 = _T_68049[10:0]; // @[Modules.scala 78:156:@18904.4]
  assign buffer_7_766 = $signed(_T_68050); // @[Modules.scala 78:156:@18905.4]
  assign _T_68052 = $signed(buffer_7_766) + $signed(buffer_7_718); // @[Modules.scala 78:156:@18907.4]
  assign _T_68053 = _T_68052[10:0]; // @[Modules.scala 78:156:@18908.4]
  assign buffer_7_767 = $signed(_T_68053); // @[Modules.scala 78:156:@18909.4]
  assign _T_68055 = $signed(buffer_7_767) + $signed(buffer_7_719); // @[Modules.scala 78:156:@18911.4]
  assign _T_68056 = _T_68055[10:0]; // @[Modules.scala 78:156:@18912.4]
  assign buffer_7_768 = $signed(_T_68056); // @[Modules.scala 78:156:@18913.4]
  assign _T_68058 = $signed(buffer_7_768) + $signed(buffer_7_720); // @[Modules.scala 78:156:@18915.4]
  assign _T_68059 = _T_68058[10:0]; // @[Modules.scala 78:156:@18916.4]
  assign buffer_7_769 = $signed(_T_68059); // @[Modules.scala 78:156:@18917.4]
  assign _T_68061 = $signed(buffer_7_769) + $signed(buffer_7_721); // @[Modules.scala 78:156:@18919.4]
  assign _T_68062 = _T_68061[10:0]; // @[Modules.scala 78:156:@18920.4]
  assign buffer_7_770 = $signed(_T_68062); // @[Modules.scala 78:156:@18921.4]
  assign _T_68064 = $signed(buffer_7_770) + $signed(buffer_7_722); // @[Modules.scala 78:156:@18923.4]
  assign _T_68065 = _T_68064[10:0]; // @[Modules.scala 78:156:@18924.4]
  assign buffer_7_771 = $signed(_T_68065); // @[Modules.scala 78:156:@18925.4]
  assign _T_68067 = $signed(buffer_7_771) + $signed(buffer_7_723); // @[Modules.scala 78:156:@18927.4]
  assign _T_68068 = _T_68067[10:0]; // @[Modules.scala 78:156:@18928.4]
  assign buffer_7_772 = $signed(_T_68068); // @[Modules.scala 78:156:@18929.4]
  assign _T_68070 = $signed(buffer_7_772) + $signed(buffer_7_724); // @[Modules.scala 78:156:@18931.4]
  assign _T_68071 = _T_68070[10:0]; // @[Modules.scala 78:156:@18932.4]
  assign buffer_7_773 = $signed(_T_68071); // @[Modules.scala 78:156:@18933.4]
  assign _T_68073 = $signed(buffer_7_773) + $signed(buffer_7_725); // @[Modules.scala 78:156:@18935.4]
  assign _T_68074 = _T_68073[10:0]; // @[Modules.scala 78:156:@18936.4]
  assign buffer_7_774 = $signed(_T_68074); // @[Modules.scala 78:156:@18937.4]
  assign _T_68076 = $signed(buffer_7_774) + $signed(buffer_7_726); // @[Modules.scala 78:156:@18939.4]
  assign _T_68077 = _T_68076[10:0]; // @[Modules.scala 78:156:@18940.4]
  assign buffer_7_775 = $signed(_T_68077); // @[Modules.scala 78:156:@18941.4]
  assign _T_68079 = $signed(buffer_7_775) + $signed(buffer_7_727); // @[Modules.scala 78:156:@18943.4]
  assign _T_68080 = _T_68079[10:0]; // @[Modules.scala 78:156:@18944.4]
  assign buffer_7_776 = $signed(_T_68080); // @[Modules.scala 78:156:@18945.4]
  assign _T_68082 = $signed(buffer_7_776) + $signed(buffer_7_728); // @[Modules.scala 78:156:@18947.4]
  assign _T_68083 = _T_68082[10:0]; // @[Modules.scala 78:156:@18948.4]
  assign buffer_7_777 = $signed(_T_68083); // @[Modules.scala 78:156:@18949.4]
  assign _T_68085 = $signed(buffer_7_777) + $signed(buffer_7_729); // @[Modules.scala 78:156:@18951.4]
  assign _T_68086 = _T_68085[10:0]; // @[Modules.scala 78:156:@18952.4]
  assign buffer_7_778 = $signed(_T_68086); // @[Modules.scala 78:156:@18953.4]
  assign _T_68088 = $signed(buffer_7_778) + $signed(buffer_0_701); // @[Modules.scala 78:156:@18955.4]
  assign _T_68089 = _T_68088[10:0]; // @[Modules.scala 78:156:@18956.4]
  assign buffer_7_779 = $signed(_T_68089); // @[Modules.scala 78:156:@18957.4]
  assign _T_68091 = $signed(buffer_7_779) + $signed(buffer_7_731); // @[Modules.scala 78:156:@18959.4]
  assign _T_68092 = _T_68091[10:0]; // @[Modules.scala 78:156:@18960.4]
  assign buffer_7_780 = $signed(_T_68092); // @[Modules.scala 78:156:@18961.4]
  assign _T_68094 = $signed(buffer_7_780) + $signed(buffer_0_701); // @[Modules.scala 78:156:@18963.4]
  assign _T_68095 = _T_68094[10:0]; // @[Modules.scala 78:156:@18964.4]
  assign buffer_7_781 = $signed(_T_68095); // @[Modules.scala 78:156:@18965.4]
  assign _T_68097 = $signed(buffer_7_781) + $signed(buffer_7_733); // @[Modules.scala 78:156:@18967.4]
  assign _T_68098 = _T_68097[10:0]; // @[Modules.scala 78:156:@18968.4]
  assign buffer_7_782 = $signed(_T_68098); // @[Modules.scala 78:156:@18969.4]
  assign _T_68100 = $signed(buffer_7_782) + $signed(buffer_7_734); // @[Modules.scala 78:156:@18971.4]
  assign _T_68101 = _T_68100[10:0]; // @[Modules.scala 78:156:@18972.4]
  assign buffer_7_783 = $signed(_T_68101); // @[Modules.scala 78:156:@18973.4]
  assign _T_68334 = $signed(io_in_362) + $signed(io_in_363); // @[Modules.scala 37:46:@19298.4]
  assign _T_68335 = _T_68334[4:0]; // @[Modules.scala 37:46:@19299.4]
  assign _T_68336 = $signed(_T_68335); // @[Modules.scala 37:46:@19300.4]
  assign _T_68355 = $signed(io_in_394) + $signed(io_in_395); // @[Modules.scala 37:46:@19329.4]
  assign _T_68356 = _T_68355[4:0]; // @[Modules.scala 37:46:@19330.4]
  assign _T_68357 = $signed(_T_68356); // @[Modules.scala 37:46:@19331.4]
  assign _T_68626 = $signed(buffer_1_4) + $signed(buffer_2_5); // @[Modules.scala 65:57:@19724.4]
  assign _T_68627 = _T_68626[10:0]; // @[Modules.scala 65:57:@19725.4]
  assign buffer_8_394 = $signed(_T_68627); // @[Modules.scala 65:57:@19726.4]
  assign _T_68635 = $signed(buffer_0_10) + $signed(buffer_2_11); // @[Modules.scala 65:57:@19736.4]
  assign _T_68636 = _T_68635[10:0]; // @[Modules.scala 65:57:@19737.4]
  assign buffer_8_397 = $signed(_T_68636); // @[Modules.scala 65:57:@19738.4]
  assign _T_68641 = $signed(buffer_3_14) + $signed(buffer_0_15); // @[Modules.scala 65:57:@19744.4]
  assign _T_68642 = _T_68641[10:0]; // @[Modules.scala 65:57:@19745.4]
  assign buffer_8_399 = $signed(_T_68642); // @[Modules.scala 65:57:@19746.4]
  assign _T_68686 = $signed(buffer_4_44) + $signed(11'sh0); // @[Modules.scala 65:57:@19804.4]
  assign _T_68687 = _T_68686[10:0]; // @[Modules.scala 65:57:@19805.4]
  assign buffer_8_414 = $signed(_T_68687); // @[Modules.scala 65:57:@19806.4]
  assign buffer_8_55 = {{6{io_in_111[4]}},io_in_111}; // @[Modules.scala 32:22:@8.4]
  assign _T_68701 = $signed(11'sh0) + $signed(buffer_8_55); // @[Modules.scala 65:57:@19824.4]
  assign _T_68702 = _T_68701[10:0]; // @[Modules.scala 65:57:@19825.4]
  assign buffer_8_419 = $signed(_T_68702); // @[Modules.scala 65:57:@19826.4]
  assign _T_68704 = $signed(11'sh0) + $signed(buffer_3_57); // @[Modules.scala 65:57:@19828.4]
  assign _T_68705 = _T_68704[10:0]; // @[Modules.scala 65:57:@19829.4]
  assign buffer_8_420 = $signed(_T_68705); // @[Modules.scala 65:57:@19830.4]
  assign buffer_8_60 = {{6{io_in_121[4]}},io_in_121}; // @[Modules.scala 32:22:@8.4]
  assign buffer_8_61 = {{6{io_in_123[4]}},io_in_123}; // @[Modules.scala 32:22:@8.4]
  assign _T_68710 = $signed(buffer_8_60) + $signed(buffer_8_61); // @[Modules.scala 65:57:@19836.4]
  assign _T_68711 = _T_68710[10:0]; // @[Modules.scala 65:57:@19837.4]
  assign buffer_8_422 = $signed(_T_68711); // @[Modules.scala 65:57:@19838.4]
  assign buffer_8_62 = {{6{io_in_125[4]}},io_in_125}; // @[Modules.scala 32:22:@8.4]
  assign _T_68713 = $signed(buffer_8_62) + $signed(buffer_7_63); // @[Modules.scala 65:57:@19840.4]
  assign _T_68714 = _T_68713[10:0]; // @[Modules.scala 65:57:@19841.4]
  assign buffer_8_423 = $signed(_T_68714); // @[Modules.scala 65:57:@19842.4]
  assign _T_68725 = $signed(buffer_0_70) + $signed(buffer_5_71); // @[Modules.scala 65:57:@19856.4]
  assign _T_68726 = _T_68725[10:0]; // @[Modules.scala 65:57:@19857.4]
  assign buffer_8_427 = $signed(_T_68726); // @[Modules.scala 65:57:@19858.4]
  assign _T_68743 = $signed(buffer_0_82) + $signed(11'sh0); // @[Modules.scala 65:57:@19880.4]
  assign _T_68744 = _T_68743[10:0]; // @[Modules.scala 65:57:@19881.4]
  assign buffer_8_433 = $signed(_T_68744); // @[Modules.scala 65:57:@19882.4]
  assign buffer_8_96 = {{6{io_in_192[4]}},io_in_192}; // @[Modules.scala 32:22:@8.4]
  assign _T_68764 = $signed(buffer_8_96) + $signed(buffer_6_97); // @[Modules.scala 65:57:@19908.4]
  assign _T_68765 = _T_68764[10:0]; // @[Modules.scala 65:57:@19909.4]
  assign buffer_8_440 = $signed(_T_68765); // @[Modules.scala 65:57:@19910.4]
  assign _T_68773 = $signed(buffer_6_102) + $signed(buffer_1_103); // @[Modules.scala 65:57:@19920.4]
  assign _T_68774 = _T_68773[10:0]; // @[Modules.scala 65:57:@19921.4]
  assign buffer_8_443 = $signed(_T_68774); // @[Modules.scala 65:57:@19922.4]
  assign _T_68779 = $signed(11'sh0) + $signed(buffer_1_107); // @[Modules.scala 65:57:@19928.4]
  assign _T_68780 = _T_68779[10:0]; // @[Modules.scala 65:57:@19929.4]
  assign buffer_8_445 = $signed(_T_68780); // @[Modules.scala 65:57:@19930.4]
  assign buffer_8_112 = {{6{io_in_225[4]}},io_in_225}; // @[Modules.scala 32:22:@8.4]
  assign _T_68788 = $signed(buffer_8_112) + $signed(buffer_3_113); // @[Modules.scala 65:57:@19940.4]
  assign _T_68789 = _T_68788[10:0]; // @[Modules.scala 65:57:@19941.4]
  assign buffer_8_448 = $signed(_T_68789); // @[Modules.scala 65:57:@19942.4]
  assign buffer_8_115 = {{6{io_in_230[4]}},io_in_230}; // @[Modules.scala 32:22:@8.4]
  assign _T_68791 = $signed(buffer_3_114) + $signed(buffer_8_115); // @[Modules.scala 65:57:@19944.4]
  assign _T_68792 = _T_68791[10:0]; // @[Modules.scala 65:57:@19945.4]
  assign buffer_8_449 = $signed(_T_68792); // @[Modules.scala 65:57:@19946.4]
  assign buffer_8_118 = {{6{io_in_236[4]}},io_in_236}; // @[Modules.scala 32:22:@8.4]
  assign _T_68797 = $signed(buffer_8_118) + $signed(11'sh0); // @[Modules.scala 65:57:@19952.4]
  assign _T_68798 = _T_68797[10:0]; // @[Modules.scala 65:57:@19953.4]
  assign buffer_8_451 = $signed(_T_68798); // @[Modules.scala 65:57:@19954.4]
  assign _T_68800 = $signed(11'sh0) + $signed(buffer_3_121); // @[Modules.scala 65:57:@19956.4]
  assign _T_68801 = _T_68800[10:0]; // @[Modules.scala 65:57:@19957.4]
  assign buffer_8_452 = $signed(_T_68801); // @[Modules.scala 65:57:@19958.4]
  assign _T_68803 = $signed(buffer_4_122) + $signed(buffer_6_123); // @[Modules.scala 65:57:@19960.4]
  assign _T_68804 = _T_68803[10:0]; // @[Modules.scala 65:57:@19961.4]
  assign buffer_8_453 = $signed(_T_68804); // @[Modules.scala 65:57:@19962.4]
  assign buffer_8_127 = {{6{io_in_254[4]}},io_in_254}; // @[Modules.scala 32:22:@8.4]
  assign _T_68809 = $signed(buffer_5_126) + $signed(buffer_8_127); // @[Modules.scala 65:57:@19968.4]
  assign _T_68810 = _T_68809[10:0]; // @[Modules.scala 65:57:@19969.4]
  assign buffer_8_455 = $signed(_T_68810); // @[Modules.scala 65:57:@19970.4]
  assign buffer_8_128 = {{6{io_in_256[4]}},io_in_256}; // @[Modules.scala 32:22:@8.4]
  assign _T_68812 = $signed(buffer_8_128) + $signed(11'sh0); // @[Modules.scala 65:57:@19972.4]
  assign _T_68813 = _T_68812[10:0]; // @[Modules.scala 65:57:@19973.4]
  assign buffer_8_456 = $signed(_T_68813); // @[Modules.scala 65:57:@19974.4]
  assign _T_68824 = $signed(buffer_3_136) + $signed(buffer_5_137); // @[Modules.scala 65:57:@19988.4]
  assign _T_68825 = _T_68824[10:0]; // @[Modules.scala 65:57:@19989.4]
  assign buffer_8_460 = $signed(_T_68825); // @[Modules.scala 65:57:@19990.4]
  assign buffer_8_141 = {{6{io_in_282[4]}},io_in_282}; // @[Modules.scala 32:22:@8.4]
  assign _T_68830 = $signed(buffer_5_140) + $signed(buffer_8_141); // @[Modules.scala 65:57:@19996.4]
  assign _T_68831 = _T_68830[10:0]; // @[Modules.scala 65:57:@19997.4]
  assign buffer_8_462 = $signed(_T_68831); // @[Modules.scala 65:57:@19998.4]
  assign _T_68851 = $signed(buffer_4_154) + $signed(buffer_3_155); // @[Modules.scala 65:57:@20024.4]
  assign _T_68852 = _T_68851[10:0]; // @[Modules.scala 65:57:@20025.4]
  assign buffer_8_469 = $signed(_T_68852); // @[Modules.scala 65:57:@20026.4]
  assign _T_68863 = $signed(buffer_6_162) + $signed(11'sh0); // @[Modules.scala 65:57:@20040.4]
  assign _T_68864 = _T_68863[10:0]; // @[Modules.scala 65:57:@20041.4]
  assign buffer_8_473 = $signed(_T_68864); // @[Modules.scala 65:57:@20042.4]
  assign _T_68872 = $signed(buffer_0_168) + $signed(buffer_5_169); // @[Modules.scala 65:57:@20052.4]
  assign _T_68873 = _T_68872[10:0]; // @[Modules.scala 65:57:@20053.4]
  assign buffer_8_476 = $signed(_T_68873); // @[Modules.scala 65:57:@20054.4]
  assign _T_68884 = $signed(11'sh0) + $signed(buffer_5_177); // @[Modules.scala 65:57:@20068.4]
  assign _T_68885 = _T_68884[10:0]; // @[Modules.scala 65:57:@20069.4]
  assign buffer_8_480 = $signed(_T_68885); // @[Modules.scala 65:57:@20070.4]
  assign buffer_8_181 = {{6{_T_68336[4]}},_T_68336}; // @[Modules.scala 32:22:@8.4]
  assign _T_68890 = $signed(11'sh0) + $signed(buffer_8_181); // @[Modules.scala 65:57:@20076.4]
  assign _T_68891 = _T_68890[10:0]; // @[Modules.scala 65:57:@20077.4]
  assign buffer_8_482 = $signed(_T_68891); // @[Modules.scala 65:57:@20078.4]
  assign buffer_8_189 = {{6{io_in_378[4]}},io_in_378}; // @[Modules.scala 32:22:@8.4]
  assign _T_68902 = $signed(buffer_0_188) + $signed(buffer_8_189); // @[Modules.scala 65:57:@20092.4]
  assign _T_68903 = _T_68902[10:0]; // @[Modules.scala 65:57:@20093.4]
  assign buffer_8_486 = $signed(_T_68903); // @[Modules.scala 65:57:@20094.4]
  assign buffer_8_192 = {{6{io_in_384[4]}},io_in_384}; // @[Modules.scala 32:22:@8.4]
  assign _T_68908 = $signed(buffer_8_192) + $signed(11'sh0); // @[Modules.scala 65:57:@20100.4]
  assign _T_68909 = _T_68908[10:0]; // @[Modules.scala 65:57:@20101.4]
  assign buffer_8_488 = $signed(_T_68909); // @[Modules.scala 65:57:@20102.4]
  assign buffer_8_197 = {{6{_T_68357[4]}},_T_68357}; // @[Modules.scala 32:22:@8.4]
  assign _T_68914 = $signed(buffer_6_196) + $signed(buffer_8_197); // @[Modules.scala 65:57:@20108.4]
  assign _T_68915 = _T_68914[10:0]; // @[Modules.scala 65:57:@20109.4]
  assign buffer_8_490 = $signed(_T_68915); // @[Modules.scala 65:57:@20110.4]
  assign _T_68920 = $signed(buffer_0_200) + $signed(buffer_3_201); // @[Modules.scala 65:57:@20116.4]
  assign _T_68921 = _T_68920[10:0]; // @[Modules.scala 65:57:@20117.4]
  assign buffer_8_492 = $signed(_T_68921); // @[Modules.scala 65:57:@20118.4]
  assign buffer_8_204 = {{6{io_in_409[4]}},io_in_409}; // @[Modules.scala 32:22:@8.4]
  assign _T_68926 = $signed(buffer_8_204) + $signed(buffer_0_205); // @[Modules.scala 65:57:@20124.4]
  assign _T_68927 = _T_68926[10:0]; // @[Modules.scala 65:57:@20125.4]
  assign buffer_8_494 = $signed(_T_68927); // @[Modules.scala 65:57:@20126.4]
  assign _T_68929 = $signed(buffer_4_206) + $signed(11'sh0); // @[Modules.scala 65:57:@20128.4]
  assign _T_68930 = _T_68929[10:0]; // @[Modules.scala 65:57:@20129.4]
  assign buffer_8_495 = $signed(_T_68930); // @[Modules.scala 65:57:@20130.4]
  assign _T_68950 = $signed(11'sh0) + $signed(buffer_6_221); // @[Modules.scala 65:57:@20156.4]
  assign _T_68951 = _T_68950[10:0]; // @[Modules.scala 65:57:@20157.4]
  assign buffer_8_502 = $signed(_T_68951); // @[Modules.scala 65:57:@20158.4]
  assign _T_68953 = $signed(11'sh0) + $signed(buffer_3_223); // @[Modules.scala 65:57:@20160.4]
  assign _T_68954 = _T_68953[10:0]; // @[Modules.scala 65:57:@20161.4]
  assign buffer_8_503 = $signed(_T_68954); // @[Modules.scala 65:57:@20162.4]
  assign _T_68956 = $signed(buffer_3_224) + $signed(buffer_7_225); // @[Modules.scala 65:57:@20164.4]
  assign _T_68957 = _T_68956[10:0]; // @[Modules.scala 65:57:@20165.4]
  assign buffer_8_504 = $signed(_T_68957); // @[Modules.scala 65:57:@20166.4]
  assign buffer_8_239 = {{6{io_in_479[4]}},io_in_479}; // @[Modules.scala 32:22:@8.4]
  assign _T_68977 = $signed(buffer_2_238) + $signed(buffer_8_239); // @[Modules.scala 65:57:@20192.4]
  assign _T_68978 = _T_68977[10:0]; // @[Modules.scala 65:57:@20193.4]
  assign buffer_8_511 = $signed(_T_68978); // @[Modules.scala 65:57:@20194.4]
  assign _T_68989 = $signed(buffer_4_246) + $signed(11'sh0); // @[Modules.scala 65:57:@20208.4]
  assign _T_68990 = _T_68989[10:0]; // @[Modules.scala 65:57:@20209.4]
  assign buffer_8_515 = $signed(_T_68990); // @[Modules.scala 65:57:@20210.4]
  assign buffer_8_248 = {{6{io_in_497[4]}},io_in_497}; // @[Modules.scala 32:22:@8.4]
  assign _T_68992 = $signed(buffer_8_248) + $signed(buffer_0_249); // @[Modules.scala 65:57:@20212.4]
  assign _T_68993 = _T_68992[10:0]; // @[Modules.scala 65:57:@20213.4]
  assign buffer_8_516 = $signed(_T_68993); // @[Modules.scala 65:57:@20214.4]
  assign _T_68998 = $signed(buffer_1_252) + $signed(buffer_0_253); // @[Modules.scala 65:57:@20220.4]
  assign _T_68999 = _T_68998[10:0]; // @[Modules.scala 65:57:@20221.4]
  assign buffer_8_518 = $signed(_T_68999); // @[Modules.scala 65:57:@20222.4]
  assign buffer_8_254 = {{6{io_in_509[4]}},io_in_509}; // @[Modules.scala 32:22:@8.4]
  assign _T_69001 = $signed(buffer_8_254) + $signed(buffer_1_255); // @[Modules.scala 65:57:@20224.4]
  assign _T_69002 = _T_69001[10:0]; // @[Modules.scala 65:57:@20225.4]
  assign buffer_8_519 = $signed(_T_69002); // @[Modules.scala 65:57:@20226.4]
  assign _T_69019 = $signed(11'sh0) + $signed(buffer_1_267); // @[Modules.scala 65:57:@20248.4]
  assign _T_69020 = _T_69019[10:0]; // @[Modules.scala 65:57:@20249.4]
  assign buffer_8_525 = $signed(_T_69020); // @[Modules.scala 65:57:@20250.4]
  assign _T_69022 = $signed(buffer_1_268) + $signed(buffer_7_269); // @[Modules.scala 65:57:@20252.4]
  assign _T_69023 = _T_69022[10:0]; // @[Modules.scala 65:57:@20253.4]
  assign buffer_8_526 = $signed(_T_69023); // @[Modules.scala 65:57:@20254.4]
  assign _T_69028 = $signed(buffer_2_272) + $signed(buffer_3_273); // @[Modules.scala 65:57:@20260.4]
  assign _T_69029 = _T_69028[10:0]; // @[Modules.scala 65:57:@20261.4]
  assign buffer_8_528 = $signed(_T_69029); // @[Modules.scala 65:57:@20262.4]
  assign _T_69034 = $signed(buffer_7_276) + $signed(buffer_5_277); // @[Modules.scala 65:57:@20268.4]
  assign _T_69035 = _T_69034[10:0]; // @[Modules.scala 65:57:@20269.4]
  assign buffer_8_530 = $signed(_T_69035); // @[Modules.scala 65:57:@20270.4]
  assign _T_69040 = $signed(11'sh0) + $signed(buffer_1_281); // @[Modules.scala 65:57:@20276.4]
  assign _T_69041 = _T_69040[10:0]; // @[Modules.scala 65:57:@20277.4]
  assign buffer_8_532 = $signed(_T_69041); // @[Modules.scala 65:57:@20278.4]
  assign _T_69043 = $signed(buffer_5_282) + $signed(buffer_1_283); // @[Modules.scala 65:57:@20280.4]
  assign _T_69044 = _T_69043[10:0]; // @[Modules.scala 65:57:@20281.4]
  assign buffer_8_533 = $signed(_T_69044); // @[Modules.scala 65:57:@20282.4]
  assign buffer_8_284 = {{6{io_in_569[4]}},io_in_569}; // @[Modules.scala 32:22:@8.4]
  assign _T_69046 = $signed(buffer_8_284) + $signed(11'sh0); // @[Modules.scala 65:57:@20284.4]
  assign _T_69047 = _T_69046[10:0]; // @[Modules.scala 65:57:@20285.4]
  assign buffer_8_534 = $signed(_T_69047); // @[Modules.scala 65:57:@20286.4]
  assign _T_69058 = $signed(buffer_0_292) + $signed(buffer_7_293); // @[Modules.scala 65:57:@20300.4]
  assign _T_69059 = _T_69058[10:0]; // @[Modules.scala 65:57:@20301.4]
  assign buffer_8_538 = $signed(_T_69059); // @[Modules.scala 65:57:@20302.4]
  assign buffer_8_298 = {{6{io_in_597[4]}},io_in_597}; // @[Modules.scala 32:22:@8.4]
  assign _T_69067 = $signed(buffer_8_298) + $signed(11'sh0); // @[Modules.scala 65:57:@20312.4]
  assign _T_69068 = _T_69067[10:0]; // @[Modules.scala 65:57:@20313.4]
  assign buffer_8_541 = $signed(_T_69068); // @[Modules.scala 65:57:@20314.4]
  assign _T_69070 = $signed(11'sh0) + $signed(buffer_7_301); // @[Modules.scala 65:57:@20316.4]
  assign _T_69071 = _T_69070[10:0]; // @[Modules.scala 65:57:@20317.4]
  assign buffer_8_542 = $signed(_T_69071); // @[Modules.scala 65:57:@20318.4]
  assign buffer_8_303 = {{6{io_in_607[4]}},io_in_607}; // @[Modules.scala 32:22:@8.4]
  assign _T_69073 = $signed(11'sh0) + $signed(buffer_8_303); // @[Modules.scala 65:57:@20320.4]
  assign _T_69074 = _T_69073[10:0]; // @[Modules.scala 65:57:@20321.4]
  assign buffer_8_543 = $signed(_T_69074); // @[Modules.scala 65:57:@20322.4]
  assign buffer_8_311 = {{6{io_in_623[4]}},io_in_623}; // @[Modules.scala 32:22:@8.4]
  assign _T_69085 = $signed(buffer_3_310) + $signed(buffer_8_311); // @[Modules.scala 65:57:@20336.4]
  assign _T_69086 = _T_69085[10:0]; // @[Modules.scala 65:57:@20337.4]
  assign buffer_8_547 = $signed(_T_69086); // @[Modules.scala 65:57:@20338.4]
  assign _T_69088 = $signed(buffer_1_312) + $signed(11'sh0); // @[Modules.scala 65:57:@20340.4]
  assign _T_69089 = _T_69088[10:0]; // @[Modules.scala 65:57:@20341.4]
  assign buffer_8_548 = $signed(_T_69089); // @[Modules.scala 65:57:@20342.4]
  assign _T_69091 = $signed(11'sh0) + $signed(buffer_6_315); // @[Modules.scala 65:57:@20344.4]
  assign _T_69092 = _T_69091[10:0]; // @[Modules.scala 65:57:@20345.4]
  assign buffer_8_549 = $signed(_T_69092); // @[Modules.scala 65:57:@20346.4]
  assign _T_69106 = $signed(buffer_1_324) + $signed(buffer_2_325); // @[Modules.scala 65:57:@20364.4]
  assign _T_69107 = _T_69106[10:0]; // @[Modules.scala 65:57:@20365.4]
  assign buffer_8_554 = $signed(_T_69107); // @[Modules.scala 65:57:@20366.4]
  assign buffer_8_327 = {{6{io_in_655[4]}},io_in_655}; // @[Modules.scala 32:22:@8.4]
  assign _T_69109 = $signed(buffer_3_326) + $signed(buffer_8_327); // @[Modules.scala 65:57:@20368.4]
  assign _T_69110 = _T_69109[10:0]; // @[Modules.scala 65:57:@20369.4]
  assign buffer_8_555 = $signed(_T_69110); // @[Modules.scala 65:57:@20370.4]
  assign _T_69115 = $signed(buffer_4_330) + $signed(buffer_0_331); // @[Modules.scala 65:57:@20376.4]
  assign _T_69116 = _T_69115[10:0]; // @[Modules.scala 65:57:@20377.4]
  assign buffer_8_557 = $signed(_T_69116); // @[Modules.scala 65:57:@20378.4]
  assign _T_69121 = $signed(buffer_4_334) + $signed(buffer_3_335); // @[Modules.scala 65:57:@20384.4]
  assign _T_69122 = _T_69121[10:0]; // @[Modules.scala 65:57:@20385.4]
  assign buffer_8_559 = $signed(_T_69122); // @[Modules.scala 65:57:@20386.4]
  assign _T_69127 = $signed(buffer_4_338) + $signed(11'sh0); // @[Modules.scala 65:57:@20392.4]
  assign _T_69128 = _T_69127[10:0]; // @[Modules.scala 65:57:@20393.4]
  assign buffer_8_561 = $signed(_T_69128); // @[Modules.scala 65:57:@20394.4]
  assign _T_69145 = $signed(buffer_5_350) + $signed(buffer_3_351); // @[Modules.scala 65:57:@20416.4]
  assign _T_69146 = _T_69145[10:0]; // @[Modules.scala 65:57:@20417.4]
  assign buffer_8_567 = $signed(_T_69146); // @[Modules.scala 65:57:@20418.4]
  assign _T_69184 = $signed(11'sh0) + $signed(buffer_3_377); // @[Modules.scala 65:57:@20468.4]
  assign _T_69185 = _T_69184[10:0]; // @[Modules.scala 65:57:@20469.4]
  assign buffer_8_580 = $signed(_T_69185); // @[Modules.scala 65:57:@20470.4]
  assign buffer_8_379 = {{6{io_in_759[4]}},io_in_759}; // @[Modules.scala 32:22:@8.4]
  assign _T_69187 = $signed(buffer_1_378) + $signed(buffer_8_379); // @[Modules.scala 65:57:@20472.4]
  assign _T_69188 = _T_69187[10:0]; // @[Modules.scala 65:57:@20473.4]
  assign buffer_8_581 = $signed(_T_69188); // @[Modules.scala 65:57:@20474.4]
  assign buffer_8_382 = {{6{io_in_764[4]}},io_in_764}; // @[Modules.scala 32:22:@8.4]
  assign _T_69193 = $signed(buffer_8_382) + $signed(11'sh0); // @[Modules.scala 65:57:@20480.4]
  assign _T_69194 = _T_69193[10:0]; // @[Modules.scala 65:57:@20481.4]
  assign buffer_8_583 = $signed(_T_69194); // @[Modules.scala 65:57:@20482.4]
  assign _T_69202 = $signed(11'sh0) + $signed(buffer_5_389); // @[Modules.scala 65:57:@20492.4]
  assign _T_69203 = _T_69202[10:0]; // @[Modules.scala 65:57:@20493.4]
  assign buffer_8_586 = $signed(_T_69203); // @[Modules.scala 65:57:@20494.4]
  assign _T_69211 = $signed(buffer_8_394) + $signed(buffer_4_395); // @[Modules.scala 68:83:@20504.4]
  assign _T_69212 = _T_69211[10:0]; // @[Modules.scala 68:83:@20505.4]
  assign buffer_8_589 = $signed(_T_69212); // @[Modules.scala 68:83:@20506.4]
  assign _T_69214 = $signed(buffer_3_396) + $signed(buffer_8_397); // @[Modules.scala 68:83:@20508.4]
  assign _T_69215 = _T_69214[10:0]; // @[Modules.scala 68:83:@20509.4]
  assign buffer_8_590 = $signed(_T_69215); // @[Modules.scala 68:83:@20510.4]
  assign _T_69217 = $signed(buffer_3_398) + $signed(buffer_8_399); // @[Modules.scala 68:83:@20512.4]
  assign _T_69218 = _T_69217[10:0]; // @[Modules.scala 68:83:@20513.4]
  assign buffer_8_591 = $signed(_T_69218); // @[Modules.scala 68:83:@20514.4]
  assign _T_69226 = $signed(buffer_0_395) + $signed(buffer_7_405); // @[Modules.scala 68:83:@20524.4]
  assign _T_69227 = _T_69226[10:0]; // @[Modules.scala 68:83:@20525.4]
  assign buffer_8_594 = $signed(_T_69227); // @[Modules.scala 68:83:@20526.4]
  assign _T_69238 = $signed(buffer_0_412) + $signed(buffer_6_413); // @[Modules.scala 68:83:@20540.4]
  assign _T_69239 = _T_69238[10:0]; // @[Modules.scala 68:83:@20541.4]
  assign buffer_8_598 = $signed(_T_69239); // @[Modules.scala 68:83:@20542.4]
  assign _T_69241 = $signed(buffer_8_414) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20544.4]
  assign _T_69242 = _T_69241[10:0]; // @[Modules.scala 68:83:@20545.4]
  assign buffer_8_599 = $signed(_T_69242); // @[Modules.scala 68:83:@20546.4]
  assign _T_69247 = $signed(buffer_0_395) + $signed(buffer_8_419); // @[Modules.scala 68:83:@20552.4]
  assign _T_69248 = _T_69247[10:0]; // @[Modules.scala 68:83:@20553.4]
  assign buffer_8_601 = $signed(_T_69248); // @[Modules.scala 68:83:@20554.4]
  assign _T_69250 = $signed(buffer_8_420) + $signed(buffer_5_421); // @[Modules.scala 68:83:@20556.4]
  assign _T_69251 = _T_69250[10:0]; // @[Modules.scala 68:83:@20557.4]
  assign buffer_8_602 = $signed(_T_69251); // @[Modules.scala 68:83:@20558.4]
  assign _T_69253 = $signed(buffer_8_422) + $signed(buffer_8_423); // @[Modules.scala 68:83:@20560.4]
  assign _T_69254 = _T_69253[10:0]; // @[Modules.scala 68:83:@20561.4]
  assign buffer_8_603 = $signed(_T_69254); // @[Modules.scala 68:83:@20562.4]
  assign _T_69259 = $signed(buffer_0_395) + $signed(buffer_8_427); // @[Modules.scala 68:83:@20568.4]
  assign _T_69260 = _T_69259[10:0]; // @[Modules.scala 68:83:@20569.4]
  assign buffer_8_605 = $signed(_T_69260); // @[Modules.scala 68:83:@20570.4]
  assign _T_69268 = $signed(buffer_1_432) + $signed(buffer_8_433); // @[Modules.scala 68:83:@20580.4]
  assign _T_69269 = _T_69268[10:0]; // @[Modules.scala 68:83:@20581.4]
  assign buffer_8_608 = $signed(_T_69269); // @[Modules.scala 68:83:@20582.4]
  assign _T_69274 = $signed(buffer_3_436) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20588.4]
  assign _T_69275 = _T_69274[10:0]; // @[Modules.scala 68:83:@20589.4]
  assign buffer_8_610 = $signed(_T_69275); // @[Modules.scala 68:83:@20590.4]
  assign _T_69277 = $signed(buffer_0_395) + $signed(buffer_4_439); // @[Modules.scala 68:83:@20592.4]
  assign _T_69278 = _T_69277[10:0]; // @[Modules.scala 68:83:@20593.4]
  assign buffer_8_611 = $signed(_T_69278); // @[Modules.scala 68:83:@20594.4]
  assign _T_69280 = $signed(buffer_8_440) + $signed(buffer_3_441); // @[Modules.scala 68:83:@20596.4]
  assign _T_69281 = _T_69280[10:0]; // @[Modules.scala 68:83:@20597.4]
  assign buffer_8_612 = $signed(_T_69281); // @[Modules.scala 68:83:@20598.4]
  assign _T_69283 = $signed(buffer_3_442) + $signed(buffer_8_443); // @[Modules.scala 68:83:@20600.4]
  assign _T_69284 = _T_69283[10:0]; // @[Modules.scala 68:83:@20601.4]
  assign buffer_8_613 = $signed(_T_69284); // @[Modules.scala 68:83:@20602.4]
  assign _T_69286 = $signed(buffer_0_395) + $signed(buffer_8_445); // @[Modules.scala 68:83:@20604.4]
  assign _T_69287 = _T_69286[10:0]; // @[Modules.scala 68:83:@20605.4]
  assign buffer_8_614 = $signed(_T_69287); // @[Modules.scala 68:83:@20606.4]
  assign _T_69289 = $signed(buffer_2_446) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20608.4]
  assign _T_69290 = _T_69289[10:0]; // @[Modules.scala 68:83:@20609.4]
  assign buffer_8_615 = $signed(_T_69290); // @[Modules.scala 68:83:@20610.4]
  assign _T_69292 = $signed(buffer_8_448) + $signed(buffer_8_449); // @[Modules.scala 68:83:@20612.4]
  assign _T_69293 = _T_69292[10:0]; // @[Modules.scala 68:83:@20613.4]
  assign buffer_8_616 = $signed(_T_69293); // @[Modules.scala 68:83:@20614.4]
  assign _T_69295 = $signed(buffer_0_395) + $signed(buffer_8_451); // @[Modules.scala 68:83:@20616.4]
  assign _T_69296 = _T_69295[10:0]; // @[Modules.scala 68:83:@20617.4]
  assign buffer_8_617 = $signed(_T_69296); // @[Modules.scala 68:83:@20618.4]
  assign _T_69298 = $signed(buffer_8_452) + $signed(buffer_8_453); // @[Modules.scala 68:83:@20620.4]
  assign _T_69299 = _T_69298[10:0]; // @[Modules.scala 68:83:@20621.4]
  assign buffer_8_618 = $signed(_T_69299); // @[Modules.scala 68:83:@20622.4]
  assign _T_69301 = $signed(buffer_0_395) + $signed(buffer_8_455); // @[Modules.scala 68:83:@20624.4]
  assign _T_69302 = _T_69301[10:0]; // @[Modules.scala 68:83:@20625.4]
  assign buffer_8_619 = $signed(_T_69302); // @[Modules.scala 68:83:@20626.4]
  assign _T_69304 = $signed(buffer_8_456) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20628.4]
  assign _T_69305 = _T_69304[10:0]; // @[Modules.scala 68:83:@20629.4]
  assign buffer_8_620 = $signed(_T_69305); // @[Modules.scala 68:83:@20630.4]
  assign _T_69307 = $signed(buffer_0_395) + $signed(buffer_5_459); // @[Modules.scala 68:83:@20632.4]
  assign _T_69308 = _T_69307[10:0]; // @[Modules.scala 68:83:@20633.4]
  assign buffer_8_621 = $signed(_T_69308); // @[Modules.scala 68:83:@20634.4]
  assign _T_69310 = $signed(buffer_8_460) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20636.4]
  assign _T_69311 = _T_69310[10:0]; // @[Modules.scala 68:83:@20637.4]
  assign buffer_8_622 = $signed(_T_69311); // @[Modules.scala 68:83:@20638.4]
  assign _T_69313 = $signed(buffer_8_462) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20640.4]
  assign _T_69314 = _T_69313[10:0]; // @[Modules.scala 68:83:@20641.4]
  assign buffer_8_623 = $signed(_T_69314); // @[Modules.scala 68:83:@20642.4]
  assign _T_69319 = $signed(buffer_3_466) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20648.4]
  assign _T_69320 = _T_69319[10:0]; // @[Modules.scala 68:83:@20649.4]
  assign buffer_8_625 = $signed(_T_69320); // @[Modules.scala 68:83:@20650.4]
  assign _T_69322 = $signed(buffer_5_468) + $signed(buffer_8_469); // @[Modules.scala 68:83:@20652.4]
  assign _T_69323 = _T_69322[10:0]; // @[Modules.scala 68:83:@20653.4]
  assign buffer_8_626 = $signed(_T_69323); // @[Modules.scala 68:83:@20654.4]
  assign _T_69328 = $signed(buffer_5_472) + $signed(buffer_8_473); // @[Modules.scala 68:83:@20660.4]
  assign _T_69329 = _T_69328[10:0]; // @[Modules.scala 68:83:@20661.4]
  assign buffer_8_628 = $signed(_T_69329); // @[Modules.scala 68:83:@20662.4]
  assign _T_69331 = $signed(buffer_0_395) + $signed(buffer_0_475); // @[Modules.scala 68:83:@20664.4]
  assign _T_69332 = _T_69331[10:0]; // @[Modules.scala 68:83:@20665.4]
  assign buffer_8_629 = $signed(_T_69332); // @[Modules.scala 68:83:@20666.4]
  assign _T_69334 = $signed(buffer_8_476) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20668.4]
  assign _T_69335 = _T_69334[10:0]; // @[Modules.scala 68:83:@20669.4]
  assign buffer_8_630 = $signed(_T_69335); // @[Modules.scala 68:83:@20670.4]
  assign _T_69340 = $signed(buffer_8_480) + $signed(buffer_5_481); // @[Modules.scala 68:83:@20676.4]
  assign _T_69341 = _T_69340[10:0]; // @[Modules.scala 68:83:@20677.4]
  assign buffer_8_632 = $signed(_T_69341); // @[Modules.scala 68:83:@20678.4]
  assign _T_69343 = $signed(buffer_8_482) + $signed(buffer_4_483); // @[Modules.scala 68:83:@20680.4]
  assign _T_69344 = _T_69343[10:0]; // @[Modules.scala 68:83:@20681.4]
  assign buffer_8_633 = $signed(_T_69344); // @[Modules.scala 68:83:@20682.4]
  assign _T_69346 = $signed(buffer_0_395) + $signed(buffer_0_485); // @[Modules.scala 68:83:@20684.4]
  assign _T_69347 = _T_69346[10:0]; // @[Modules.scala 68:83:@20685.4]
  assign buffer_8_634 = $signed(_T_69347); // @[Modules.scala 68:83:@20686.4]
  assign _T_69349 = $signed(buffer_8_486) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20688.4]
  assign _T_69350 = _T_69349[10:0]; // @[Modules.scala 68:83:@20689.4]
  assign buffer_8_635 = $signed(_T_69350); // @[Modules.scala 68:83:@20690.4]
  assign _T_69352 = $signed(buffer_8_488) + $signed(buffer_5_489); // @[Modules.scala 68:83:@20692.4]
  assign _T_69353 = _T_69352[10:0]; // @[Modules.scala 68:83:@20693.4]
  assign buffer_8_636 = $signed(_T_69353); // @[Modules.scala 68:83:@20694.4]
  assign _T_69355 = $signed(buffer_8_490) + $signed(buffer_0_491); // @[Modules.scala 68:83:@20696.4]
  assign _T_69356 = _T_69355[10:0]; // @[Modules.scala 68:83:@20697.4]
  assign buffer_8_637 = $signed(_T_69356); // @[Modules.scala 68:83:@20698.4]
  assign _T_69358 = $signed(buffer_8_492) + $signed(buffer_0_493); // @[Modules.scala 68:83:@20700.4]
  assign _T_69359 = _T_69358[10:0]; // @[Modules.scala 68:83:@20701.4]
  assign buffer_8_638 = $signed(_T_69359); // @[Modules.scala 68:83:@20702.4]
  assign _T_69361 = $signed(buffer_8_494) + $signed(buffer_8_495); // @[Modules.scala 68:83:@20704.4]
  assign _T_69362 = _T_69361[10:0]; // @[Modules.scala 68:83:@20705.4]
  assign buffer_8_639 = $signed(_T_69362); // @[Modules.scala 68:83:@20706.4]
  assign _T_69367 = $signed(buffer_7_498) + $signed(buffer_2_499); // @[Modules.scala 68:83:@20712.4]
  assign _T_69368 = _T_69367[10:0]; // @[Modules.scala 68:83:@20713.4]
  assign buffer_8_641 = $signed(_T_69368); // @[Modules.scala 68:83:@20714.4]
  assign _T_69370 = $signed(buffer_0_500) + $signed(buffer_6_501); // @[Modules.scala 68:83:@20716.4]
  assign _T_69371 = _T_69370[10:0]; // @[Modules.scala 68:83:@20717.4]
  assign buffer_8_642 = $signed(_T_69371); // @[Modules.scala 68:83:@20718.4]
  assign _T_69373 = $signed(buffer_8_502) + $signed(buffer_8_503); // @[Modules.scala 68:83:@20720.4]
  assign _T_69374 = _T_69373[10:0]; // @[Modules.scala 68:83:@20721.4]
  assign buffer_8_643 = $signed(_T_69374); // @[Modules.scala 68:83:@20722.4]
  assign _T_69376 = $signed(buffer_8_504) + $signed(buffer_3_505); // @[Modules.scala 68:83:@20724.4]
  assign _T_69377 = _T_69376[10:0]; // @[Modules.scala 68:83:@20725.4]
  assign buffer_8_644 = $signed(_T_69377); // @[Modules.scala 68:83:@20726.4]
  assign _T_69382 = $signed(buffer_0_508) + $signed(buffer_7_509); // @[Modules.scala 68:83:@20732.4]
  assign _T_69383 = _T_69382[10:0]; // @[Modules.scala 68:83:@20733.4]
  assign buffer_8_646 = $signed(_T_69383); // @[Modules.scala 68:83:@20734.4]
  assign _T_69385 = $signed(buffer_5_510) + $signed(buffer_8_511); // @[Modules.scala 68:83:@20736.4]
  assign _T_69386 = _T_69385[10:0]; // @[Modules.scala 68:83:@20737.4]
  assign buffer_8_647 = $signed(_T_69386); // @[Modules.scala 68:83:@20738.4]
  assign _T_69388 = $signed(buffer_4_512) + $signed(buffer_5_513); // @[Modules.scala 68:83:@20740.4]
  assign _T_69389 = _T_69388[10:0]; // @[Modules.scala 68:83:@20741.4]
  assign buffer_8_648 = $signed(_T_69389); // @[Modules.scala 68:83:@20742.4]
  assign _T_69391 = $signed(buffer_2_514) + $signed(buffer_8_515); // @[Modules.scala 68:83:@20744.4]
  assign _T_69392 = _T_69391[10:0]; // @[Modules.scala 68:83:@20745.4]
  assign buffer_8_649 = $signed(_T_69392); // @[Modules.scala 68:83:@20746.4]
  assign _T_69394 = $signed(buffer_8_516) + $signed(buffer_3_517); // @[Modules.scala 68:83:@20748.4]
  assign _T_69395 = _T_69394[10:0]; // @[Modules.scala 68:83:@20749.4]
  assign buffer_8_650 = $signed(_T_69395); // @[Modules.scala 68:83:@20750.4]
  assign _T_69397 = $signed(buffer_8_518) + $signed(buffer_8_519); // @[Modules.scala 68:83:@20752.4]
  assign _T_69398 = _T_69397[10:0]; // @[Modules.scala 68:83:@20753.4]
  assign buffer_8_651 = $signed(_T_69398); // @[Modules.scala 68:83:@20754.4]
  assign _T_69400 = $signed(buffer_0_395) + $signed(buffer_5_521); // @[Modules.scala 68:83:@20756.4]
  assign _T_69401 = _T_69400[10:0]; // @[Modules.scala 68:83:@20757.4]
  assign buffer_8_652 = $signed(_T_69401); // @[Modules.scala 68:83:@20758.4]
  assign _T_69403 = $signed(buffer_0_395) + $signed(buffer_7_523); // @[Modules.scala 68:83:@20760.4]
  assign _T_69404 = _T_69403[10:0]; // @[Modules.scala 68:83:@20761.4]
  assign buffer_8_653 = $signed(_T_69404); // @[Modules.scala 68:83:@20762.4]
  assign _T_69406 = $signed(buffer_3_524) + $signed(buffer_8_525); // @[Modules.scala 68:83:@20764.4]
  assign _T_69407 = _T_69406[10:0]; // @[Modules.scala 68:83:@20765.4]
  assign buffer_8_654 = $signed(_T_69407); // @[Modules.scala 68:83:@20766.4]
  assign _T_69409 = $signed(buffer_8_526) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20768.4]
  assign _T_69410 = _T_69409[10:0]; // @[Modules.scala 68:83:@20769.4]
  assign buffer_8_655 = $signed(_T_69410); // @[Modules.scala 68:83:@20770.4]
  assign _T_69412 = $signed(buffer_8_528) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20772.4]
  assign _T_69413 = _T_69412[10:0]; // @[Modules.scala 68:83:@20773.4]
  assign buffer_8_656 = $signed(_T_69413); // @[Modules.scala 68:83:@20774.4]
  assign _T_69415 = $signed(buffer_8_530) + $signed(buffer_5_531); // @[Modules.scala 68:83:@20776.4]
  assign _T_69416 = _T_69415[10:0]; // @[Modules.scala 68:83:@20777.4]
  assign buffer_8_657 = $signed(_T_69416); // @[Modules.scala 68:83:@20778.4]
  assign _T_69418 = $signed(buffer_8_532) + $signed(buffer_8_533); // @[Modules.scala 68:83:@20780.4]
  assign _T_69419 = _T_69418[10:0]; // @[Modules.scala 68:83:@20781.4]
  assign buffer_8_658 = $signed(_T_69419); // @[Modules.scala 68:83:@20782.4]
  assign _T_69421 = $signed(buffer_8_534) + $signed(buffer_0_395); // @[Modules.scala 68:83:@20784.4]
  assign _T_69422 = _T_69421[10:0]; // @[Modules.scala 68:83:@20785.4]
  assign buffer_8_659 = $signed(_T_69422); // @[Modules.scala 68:83:@20786.4]
  assign _T_69424 = $signed(buffer_0_536) + $signed(buffer_4_537); // @[Modules.scala 68:83:@20788.4]
  assign _T_69425 = _T_69424[10:0]; // @[Modules.scala 68:83:@20789.4]
  assign buffer_8_660 = $signed(_T_69425); // @[Modules.scala 68:83:@20790.4]
  assign _T_69427 = $signed(buffer_8_538) + $signed(buffer_1_539); // @[Modules.scala 68:83:@20792.4]
  assign _T_69428 = _T_69427[10:0]; // @[Modules.scala 68:83:@20793.4]
  assign buffer_8_661 = $signed(_T_69428); // @[Modules.scala 68:83:@20794.4]
  assign _T_69430 = $signed(buffer_1_540) + $signed(buffer_8_541); // @[Modules.scala 68:83:@20796.4]
  assign _T_69431 = _T_69430[10:0]; // @[Modules.scala 68:83:@20797.4]
  assign buffer_8_662 = $signed(_T_69431); // @[Modules.scala 68:83:@20798.4]
  assign _T_69433 = $signed(buffer_8_542) + $signed(buffer_8_543); // @[Modules.scala 68:83:@20800.4]
  assign _T_69434 = _T_69433[10:0]; // @[Modules.scala 68:83:@20801.4]
  assign buffer_8_663 = $signed(_T_69434); // @[Modules.scala 68:83:@20802.4]
  assign _T_69439 = $signed(buffer_1_546) + $signed(buffer_8_547); // @[Modules.scala 68:83:@20808.4]
  assign _T_69440 = _T_69439[10:0]; // @[Modules.scala 68:83:@20809.4]
  assign buffer_8_665 = $signed(_T_69440); // @[Modules.scala 68:83:@20810.4]
  assign _T_69442 = $signed(buffer_8_548) + $signed(buffer_8_549); // @[Modules.scala 68:83:@20812.4]
  assign _T_69443 = _T_69442[10:0]; // @[Modules.scala 68:83:@20813.4]
  assign buffer_8_666 = $signed(_T_69443); // @[Modules.scala 68:83:@20814.4]
  assign _T_69451 = $signed(buffer_8_554) + $signed(buffer_8_555); // @[Modules.scala 68:83:@20824.4]
  assign _T_69452 = _T_69451[10:0]; // @[Modules.scala 68:83:@20825.4]
  assign buffer_8_669 = $signed(_T_69452); // @[Modules.scala 68:83:@20826.4]
  assign _T_69454 = $signed(buffer_0_395) + $signed(buffer_8_557); // @[Modules.scala 68:83:@20828.4]
  assign _T_69455 = _T_69454[10:0]; // @[Modules.scala 68:83:@20829.4]
  assign buffer_8_670 = $signed(_T_69455); // @[Modules.scala 68:83:@20830.4]
  assign _T_69457 = $signed(buffer_0_395) + $signed(buffer_8_559); // @[Modules.scala 68:83:@20832.4]
  assign _T_69458 = _T_69457[10:0]; // @[Modules.scala 68:83:@20833.4]
  assign buffer_8_671 = $signed(_T_69458); // @[Modules.scala 68:83:@20834.4]
  assign _T_69460 = $signed(buffer_5_560) + $signed(buffer_8_561); // @[Modules.scala 68:83:@20836.4]
  assign _T_69461 = _T_69460[10:0]; // @[Modules.scala 68:83:@20837.4]
  assign buffer_8_672 = $signed(_T_69461); // @[Modules.scala 68:83:@20838.4]
  assign _T_69469 = $signed(buffer_4_566) + $signed(buffer_8_567); // @[Modules.scala 68:83:@20848.4]
  assign _T_69470 = _T_69469[10:0]; // @[Modules.scala 68:83:@20849.4]
  assign buffer_8_675 = $signed(_T_69470); // @[Modules.scala 68:83:@20850.4]
  assign _T_69490 = $signed(buffer_8_580) + $signed(buffer_8_581); // @[Modules.scala 68:83:@20876.4]
  assign _T_69491 = _T_69490[10:0]; // @[Modules.scala 68:83:@20877.4]
  assign buffer_8_682 = $signed(_T_69491); // @[Modules.scala 68:83:@20878.4]
  assign _T_69493 = $signed(buffer_4_582) + $signed(buffer_8_583); // @[Modules.scala 68:83:@20880.4]
  assign _T_69494 = _T_69493[10:0]; // @[Modules.scala 68:83:@20881.4]
  assign buffer_8_683 = $signed(_T_69494); // @[Modules.scala 68:83:@20882.4]
  assign _T_69499 = $signed(buffer_8_586) + $signed(buffer_1_587); // @[Modules.scala 68:83:@20888.4]
  assign _T_69500 = _T_69499[10:0]; // @[Modules.scala 68:83:@20889.4]
  assign buffer_8_685 = $signed(_T_69500); // @[Modules.scala 68:83:@20890.4]
  assign _T_69502 = $signed(buffer_4_588) + $signed(buffer_8_589); // @[Modules.scala 71:109:@20892.4]
  assign _T_69503 = _T_69502[10:0]; // @[Modules.scala 71:109:@20893.4]
  assign buffer_8_686 = $signed(_T_69503); // @[Modules.scala 71:109:@20894.4]
  assign _T_69505 = $signed(buffer_8_590) + $signed(buffer_8_591); // @[Modules.scala 71:109:@20896.4]
  assign _T_69506 = _T_69505[10:0]; // @[Modules.scala 71:109:@20897.4]
  assign buffer_8_687 = $signed(_T_69506); // @[Modules.scala 71:109:@20898.4]
  assign _T_69511 = $signed(buffer_8_594) + $signed(buffer_0_595); // @[Modules.scala 71:109:@20904.4]
  assign _T_69512 = _T_69511[10:0]; // @[Modules.scala 71:109:@20905.4]
  assign buffer_8_689 = $signed(_T_69512); // @[Modules.scala 71:109:@20906.4]
  assign _T_69517 = $signed(buffer_8_598) + $signed(buffer_8_599); // @[Modules.scala 71:109:@20912.4]
  assign _T_69518 = _T_69517[10:0]; // @[Modules.scala 71:109:@20913.4]
  assign buffer_8_691 = $signed(_T_69518); // @[Modules.scala 71:109:@20914.4]
  assign _T_69520 = $signed(buffer_0_593) + $signed(buffer_8_601); // @[Modules.scala 71:109:@20916.4]
  assign _T_69521 = _T_69520[10:0]; // @[Modules.scala 71:109:@20917.4]
  assign buffer_8_692 = $signed(_T_69521); // @[Modules.scala 71:109:@20918.4]
  assign _T_69523 = $signed(buffer_8_602) + $signed(buffer_8_603); // @[Modules.scala 71:109:@20920.4]
  assign _T_69524 = _T_69523[10:0]; // @[Modules.scala 71:109:@20921.4]
  assign buffer_8_693 = $signed(_T_69524); // @[Modules.scala 71:109:@20922.4]
  assign _T_69526 = $signed(buffer_0_593) + $signed(buffer_8_605); // @[Modules.scala 71:109:@20924.4]
  assign _T_69527 = _T_69526[10:0]; // @[Modules.scala 71:109:@20925.4]
  assign buffer_8_694 = $signed(_T_69527); // @[Modules.scala 71:109:@20926.4]
  assign _T_69532 = $signed(buffer_8_608) + $signed(buffer_3_609); // @[Modules.scala 71:109:@20932.4]
  assign _T_69533 = _T_69532[10:0]; // @[Modules.scala 71:109:@20933.4]
  assign buffer_8_696 = $signed(_T_69533); // @[Modules.scala 71:109:@20934.4]
  assign _T_69535 = $signed(buffer_8_610) + $signed(buffer_8_611); // @[Modules.scala 71:109:@20936.4]
  assign _T_69536 = _T_69535[10:0]; // @[Modules.scala 71:109:@20937.4]
  assign buffer_8_697 = $signed(_T_69536); // @[Modules.scala 71:109:@20938.4]
  assign _T_69538 = $signed(buffer_8_612) + $signed(buffer_8_613); // @[Modules.scala 71:109:@20940.4]
  assign _T_69539 = _T_69538[10:0]; // @[Modules.scala 71:109:@20941.4]
  assign buffer_8_698 = $signed(_T_69539); // @[Modules.scala 71:109:@20942.4]
  assign _T_69541 = $signed(buffer_8_614) + $signed(buffer_8_615); // @[Modules.scala 71:109:@20944.4]
  assign _T_69542 = _T_69541[10:0]; // @[Modules.scala 71:109:@20945.4]
  assign buffer_8_699 = $signed(_T_69542); // @[Modules.scala 71:109:@20946.4]
  assign _T_69544 = $signed(buffer_8_616) + $signed(buffer_8_617); // @[Modules.scala 71:109:@20948.4]
  assign _T_69545 = _T_69544[10:0]; // @[Modules.scala 71:109:@20949.4]
  assign buffer_8_700 = $signed(_T_69545); // @[Modules.scala 71:109:@20950.4]
  assign _T_69547 = $signed(buffer_8_618) + $signed(buffer_8_619); // @[Modules.scala 71:109:@20952.4]
  assign _T_69548 = _T_69547[10:0]; // @[Modules.scala 71:109:@20953.4]
  assign buffer_8_701 = $signed(_T_69548); // @[Modules.scala 71:109:@20954.4]
  assign _T_69550 = $signed(buffer_8_620) + $signed(buffer_8_621); // @[Modules.scala 71:109:@20956.4]
  assign _T_69551 = _T_69550[10:0]; // @[Modules.scala 71:109:@20957.4]
  assign buffer_8_702 = $signed(_T_69551); // @[Modules.scala 71:109:@20958.4]
  assign _T_69553 = $signed(buffer_8_622) + $signed(buffer_8_623); // @[Modules.scala 71:109:@20960.4]
  assign _T_69554 = _T_69553[10:0]; // @[Modules.scala 71:109:@20961.4]
  assign buffer_8_703 = $signed(_T_69554); // @[Modules.scala 71:109:@20962.4]
  assign _T_69556 = $signed(buffer_5_624) + $signed(buffer_8_625); // @[Modules.scala 71:109:@20964.4]
  assign _T_69557 = _T_69556[10:0]; // @[Modules.scala 71:109:@20965.4]
  assign buffer_8_704 = $signed(_T_69557); // @[Modules.scala 71:109:@20966.4]
  assign _T_69559 = $signed(buffer_8_626) + $signed(buffer_0_593); // @[Modules.scala 71:109:@20968.4]
  assign _T_69560 = _T_69559[10:0]; // @[Modules.scala 71:109:@20969.4]
  assign buffer_8_705 = $signed(_T_69560); // @[Modules.scala 71:109:@20970.4]
  assign _T_69562 = $signed(buffer_8_628) + $signed(buffer_8_629); // @[Modules.scala 71:109:@20972.4]
  assign _T_69563 = _T_69562[10:0]; // @[Modules.scala 71:109:@20973.4]
  assign buffer_8_706 = $signed(_T_69563); // @[Modules.scala 71:109:@20974.4]
  assign _T_69565 = $signed(buffer_8_630) + $signed(buffer_5_631); // @[Modules.scala 71:109:@20976.4]
  assign _T_69566 = _T_69565[10:0]; // @[Modules.scala 71:109:@20977.4]
  assign buffer_8_707 = $signed(_T_69566); // @[Modules.scala 71:109:@20978.4]
  assign _T_69568 = $signed(buffer_8_632) + $signed(buffer_8_633); // @[Modules.scala 71:109:@20980.4]
  assign _T_69569 = _T_69568[10:0]; // @[Modules.scala 71:109:@20981.4]
  assign buffer_8_708 = $signed(_T_69569); // @[Modules.scala 71:109:@20982.4]
  assign _T_69571 = $signed(buffer_8_634) + $signed(buffer_8_635); // @[Modules.scala 71:109:@20984.4]
  assign _T_69572 = _T_69571[10:0]; // @[Modules.scala 71:109:@20985.4]
  assign buffer_8_709 = $signed(_T_69572); // @[Modules.scala 71:109:@20986.4]
  assign _T_69574 = $signed(buffer_8_636) + $signed(buffer_8_637); // @[Modules.scala 71:109:@20988.4]
  assign _T_69575 = _T_69574[10:0]; // @[Modules.scala 71:109:@20989.4]
  assign buffer_8_710 = $signed(_T_69575); // @[Modules.scala 71:109:@20990.4]
  assign _T_69577 = $signed(buffer_8_638) + $signed(buffer_8_639); // @[Modules.scala 71:109:@20992.4]
  assign _T_69578 = _T_69577[10:0]; // @[Modules.scala 71:109:@20993.4]
  assign buffer_8_711 = $signed(_T_69578); // @[Modules.scala 71:109:@20994.4]
  assign _T_69580 = $signed(buffer_3_640) + $signed(buffer_8_641); // @[Modules.scala 71:109:@20996.4]
  assign _T_69581 = _T_69580[10:0]; // @[Modules.scala 71:109:@20997.4]
  assign buffer_8_712 = $signed(_T_69581); // @[Modules.scala 71:109:@20998.4]
  assign _T_69583 = $signed(buffer_8_642) + $signed(buffer_8_643); // @[Modules.scala 71:109:@21000.4]
  assign _T_69584 = _T_69583[10:0]; // @[Modules.scala 71:109:@21001.4]
  assign buffer_8_713 = $signed(_T_69584); // @[Modules.scala 71:109:@21002.4]
  assign _T_69586 = $signed(buffer_8_644) + $signed(buffer_2_645); // @[Modules.scala 71:109:@21004.4]
  assign _T_69587 = _T_69586[10:0]; // @[Modules.scala 71:109:@21005.4]
  assign buffer_8_714 = $signed(_T_69587); // @[Modules.scala 71:109:@21006.4]
  assign _T_69589 = $signed(buffer_8_646) + $signed(buffer_8_647); // @[Modules.scala 71:109:@21008.4]
  assign _T_69590 = _T_69589[10:0]; // @[Modules.scala 71:109:@21009.4]
  assign buffer_8_715 = $signed(_T_69590); // @[Modules.scala 71:109:@21010.4]
  assign _T_69592 = $signed(buffer_8_648) + $signed(buffer_8_649); // @[Modules.scala 71:109:@21012.4]
  assign _T_69593 = _T_69592[10:0]; // @[Modules.scala 71:109:@21013.4]
  assign buffer_8_716 = $signed(_T_69593); // @[Modules.scala 71:109:@21014.4]
  assign _T_69595 = $signed(buffer_8_650) + $signed(buffer_8_651); // @[Modules.scala 71:109:@21016.4]
  assign _T_69596 = _T_69595[10:0]; // @[Modules.scala 71:109:@21017.4]
  assign buffer_8_717 = $signed(_T_69596); // @[Modules.scala 71:109:@21018.4]
  assign _T_69598 = $signed(buffer_8_652) + $signed(buffer_8_653); // @[Modules.scala 71:109:@21020.4]
  assign _T_69599 = _T_69598[10:0]; // @[Modules.scala 71:109:@21021.4]
  assign buffer_8_718 = $signed(_T_69599); // @[Modules.scala 71:109:@21022.4]
  assign _T_69601 = $signed(buffer_8_654) + $signed(buffer_8_655); // @[Modules.scala 71:109:@21024.4]
  assign _T_69602 = _T_69601[10:0]; // @[Modules.scala 71:109:@21025.4]
  assign buffer_8_719 = $signed(_T_69602); // @[Modules.scala 71:109:@21026.4]
  assign _T_69604 = $signed(buffer_8_656) + $signed(buffer_8_657); // @[Modules.scala 71:109:@21028.4]
  assign _T_69605 = _T_69604[10:0]; // @[Modules.scala 71:109:@21029.4]
  assign buffer_8_720 = $signed(_T_69605); // @[Modules.scala 71:109:@21030.4]
  assign _T_69607 = $signed(buffer_8_658) + $signed(buffer_8_659); // @[Modules.scala 71:109:@21032.4]
  assign _T_69608 = _T_69607[10:0]; // @[Modules.scala 71:109:@21033.4]
  assign buffer_8_721 = $signed(_T_69608); // @[Modules.scala 71:109:@21034.4]
  assign _T_69610 = $signed(buffer_8_660) + $signed(buffer_8_661); // @[Modules.scala 71:109:@21036.4]
  assign _T_69611 = _T_69610[10:0]; // @[Modules.scala 71:109:@21037.4]
  assign buffer_8_722 = $signed(_T_69611); // @[Modules.scala 71:109:@21038.4]
  assign _T_69613 = $signed(buffer_8_662) + $signed(buffer_8_663); // @[Modules.scala 71:109:@21040.4]
  assign _T_69614 = _T_69613[10:0]; // @[Modules.scala 71:109:@21041.4]
  assign buffer_8_723 = $signed(_T_69614); // @[Modules.scala 71:109:@21042.4]
  assign _T_69616 = $signed(buffer_3_664) + $signed(buffer_8_665); // @[Modules.scala 71:109:@21044.4]
  assign _T_69617 = _T_69616[10:0]; // @[Modules.scala 71:109:@21045.4]
  assign buffer_8_724 = $signed(_T_69617); // @[Modules.scala 71:109:@21046.4]
  assign _T_69619 = $signed(buffer_8_666) + $signed(buffer_4_667); // @[Modules.scala 71:109:@21048.4]
  assign _T_69620 = _T_69619[10:0]; // @[Modules.scala 71:109:@21049.4]
  assign buffer_8_725 = $signed(_T_69620); // @[Modules.scala 71:109:@21050.4]
  assign _T_69622 = $signed(buffer_3_668) + $signed(buffer_8_669); // @[Modules.scala 71:109:@21052.4]
  assign _T_69623 = _T_69622[10:0]; // @[Modules.scala 71:109:@21053.4]
  assign buffer_8_726 = $signed(_T_69623); // @[Modules.scala 71:109:@21054.4]
  assign _T_69625 = $signed(buffer_8_670) + $signed(buffer_8_671); // @[Modules.scala 71:109:@21056.4]
  assign _T_69626 = _T_69625[10:0]; // @[Modules.scala 71:109:@21057.4]
  assign buffer_8_727 = $signed(_T_69626); // @[Modules.scala 71:109:@21058.4]
  assign _T_69628 = $signed(buffer_8_672) + $signed(buffer_0_593); // @[Modules.scala 71:109:@21060.4]
  assign _T_69629 = _T_69628[10:0]; // @[Modules.scala 71:109:@21061.4]
  assign buffer_8_728 = $signed(_T_69629); // @[Modules.scala 71:109:@21062.4]
  assign _T_69631 = $signed(buffer_0_593) + $signed(buffer_8_675); // @[Modules.scala 71:109:@21064.4]
  assign _T_69632 = _T_69631[10:0]; // @[Modules.scala 71:109:@21065.4]
  assign buffer_8_729 = $signed(_T_69632); // @[Modules.scala 71:109:@21066.4]
  assign _T_69637 = $signed(buffer_4_678) + $signed(buffer_0_593); // @[Modules.scala 71:109:@21072.4]
  assign _T_69638 = _T_69637[10:0]; // @[Modules.scala 71:109:@21073.4]
  assign buffer_8_731 = $signed(_T_69638); // @[Modules.scala 71:109:@21074.4]
  assign _T_69643 = $signed(buffer_8_682) + $signed(buffer_8_683); // @[Modules.scala 71:109:@21080.4]
  assign _T_69644 = _T_69643[10:0]; // @[Modules.scala 71:109:@21081.4]
  assign buffer_8_733 = $signed(_T_69644); // @[Modules.scala 71:109:@21082.4]
  assign _T_69646 = $signed(buffer_0_593) + $signed(buffer_8_685); // @[Modules.scala 71:109:@21084.4]
  assign _T_69647 = _T_69646[10:0]; // @[Modules.scala 71:109:@21085.4]
  assign buffer_8_734 = $signed(_T_69647); // @[Modules.scala 71:109:@21086.4]
  assign _T_69649 = $signed(buffer_8_686) + $signed(buffer_8_687); // @[Modules.scala 78:156:@21089.4]
  assign _T_69650 = _T_69649[10:0]; // @[Modules.scala 78:156:@21090.4]
  assign buffer_8_736 = $signed(_T_69650); // @[Modules.scala 78:156:@21091.4]
  assign _T_69652 = $signed(buffer_8_736) + $signed(buffer_0_701); // @[Modules.scala 78:156:@21093.4]
  assign _T_69653 = _T_69652[10:0]; // @[Modules.scala 78:156:@21094.4]
  assign buffer_8_737 = $signed(_T_69653); // @[Modules.scala 78:156:@21095.4]
  assign _T_69655 = $signed(buffer_8_737) + $signed(buffer_8_689); // @[Modules.scala 78:156:@21097.4]
  assign _T_69656 = _T_69655[10:0]; // @[Modules.scala 78:156:@21098.4]
  assign buffer_8_738 = $signed(_T_69656); // @[Modules.scala 78:156:@21099.4]
  assign _T_69658 = $signed(buffer_8_738) + $signed(buffer_0_701); // @[Modules.scala 78:156:@21101.4]
  assign _T_69659 = _T_69658[10:0]; // @[Modules.scala 78:156:@21102.4]
  assign buffer_8_739 = $signed(_T_69659); // @[Modules.scala 78:156:@21103.4]
  assign _T_69661 = $signed(buffer_8_739) + $signed(buffer_8_691); // @[Modules.scala 78:156:@21105.4]
  assign _T_69662 = _T_69661[10:0]; // @[Modules.scala 78:156:@21106.4]
  assign buffer_8_740 = $signed(_T_69662); // @[Modules.scala 78:156:@21107.4]
  assign _T_69664 = $signed(buffer_8_740) + $signed(buffer_8_692); // @[Modules.scala 78:156:@21109.4]
  assign _T_69665 = _T_69664[10:0]; // @[Modules.scala 78:156:@21110.4]
  assign buffer_8_741 = $signed(_T_69665); // @[Modules.scala 78:156:@21111.4]
  assign _T_69667 = $signed(buffer_8_741) + $signed(buffer_8_693); // @[Modules.scala 78:156:@21113.4]
  assign _T_69668 = _T_69667[10:0]; // @[Modules.scala 78:156:@21114.4]
  assign buffer_8_742 = $signed(_T_69668); // @[Modules.scala 78:156:@21115.4]
  assign _T_69670 = $signed(buffer_8_742) + $signed(buffer_8_694); // @[Modules.scala 78:156:@21117.4]
  assign _T_69671 = _T_69670[10:0]; // @[Modules.scala 78:156:@21118.4]
  assign buffer_8_743 = $signed(_T_69671); // @[Modules.scala 78:156:@21119.4]
  assign _T_69673 = $signed(buffer_8_743) + $signed(buffer_4_695); // @[Modules.scala 78:156:@21121.4]
  assign _T_69674 = _T_69673[10:0]; // @[Modules.scala 78:156:@21122.4]
  assign buffer_8_744 = $signed(_T_69674); // @[Modules.scala 78:156:@21123.4]
  assign _T_69676 = $signed(buffer_8_744) + $signed(buffer_8_696); // @[Modules.scala 78:156:@21125.4]
  assign _T_69677 = _T_69676[10:0]; // @[Modules.scala 78:156:@21126.4]
  assign buffer_8_745 = $signed(_T_69677); // @[Modules.scala 78:156:@21127.4]
  assign _T_69679 = $signed(buffer_8_745) + $signed(buffer_8_697); // @[Modules.scala 78:156:@21129.4]
  assign _T_69680 = _T_69679[10:0]; // @[Modules.scala 78:156:@21130.4]
  assign buffer_8_746 = $signed(_T_69680); // @[Modules.scala 78:156:@21131.4]
  assign _T_69682 = $signed(buffer_8_746) + $signed(buffer_8_698); // @[Modules.scala 78:156:@21133.4]
  assign _T_69683 = _T_69682[10:0]; // @[Modules.scala 78:156:@21134.4]
  assign buffer_8_747 = $signed(_T_69683); // @[Modules.scala 78:156:@21135.4]
  assign _T_69685 = $signed(buffer_8_747) + $signed(buffer_8_699); // @[Modules.scala 78:156:@21137.4]
  assign _T_69686 = _T_69685[10:0]; // @[Modules.scala 78:156:@21138.4]
  assign buffer_8_748 = $signed(_T_69686); // @[Modules.scala 78:156:@21139.4]
  assign _T_69688 = $signed(buffer_8_748) + $signed(buffer_8_700); // @[Modules.scala 78:156:@21141.4]
  assign _T_69689 = _T_69688[10:0]; // @[Modules.scala 78:156:@21142.4]
  assign buffer_8_749 = $signed(_T_69689); // @[Modules.scala 78:156:@21143.4]
  assign _T_69691 = $signed(buffer_8_749) + $signed(buffer_8_701); // @[Modules.scala 78:156:@21145.4]
  assign _T_69692 = _T_69691[10:0]; // @[Modules.scala 78:156:@21146.4]
  assign buffer_8_750 = $signed(_T_69692); // @[Modules.scala 78:156:@21147.4]
  assign _T_69694 = $signed(buffer_8_750) + $signed(buffer_8_702); // @[Modules.scala 78:156:@21149.4]
  assign _T_69695 = _T_69694[10:0]; // @[Modules.scala 78:156:@21150.4]
  assign buffer_8_751 = $signed(_T_69695); // @[Modules.scala 78:156:@21151.4]
  assign _T_69697 = $signed(buffer_8_751) + $signed(buffer_8_703); // @[Modules.scala 78:156:@21153.4]
  assign _T_69698 = _T_69697[10:0]; // @[Modules.scala 78:156:@21154.4]
  assign buffer_8_752 = $signed(_T_69698); // @[Modules.scala 78:156:@21155.4]
  assign _T_69700 = $signed(buffer_8_752) + $signed(buffer_8_704); // @[Modules.scala 78:156:@21157.4]
  assign _T_69701 = _T_69700[10:0]; // @[Modules.scala 78:156:@21158.4]
  assign buffer_8_753 = $signed(_T_69701); // @[Modules.scala 78:156:@21159.4]
  assign _T_69703 = $signed(buffer_8_753) + $signed(buffer_8_705); // @[Modules.scala 78:156:@21161.4]
  assign _T_69704 = _T_69703[10:0]; // @[Modules.scala 78:156:@21162.4]
  assign buffer_8_754 = $signed(_T_69704); // @[Modules.scala 78:156:@21163.4]
  assign _T_69706 = $signed(buffer_8_754) + $signed(buffer_8_706); // @[Modules.scala 78:156:@21165.4]
  assign _T_69707 = _T_69706[10:0]; // @[Modules.scala 78:156:@21166.4]
  assign buffer_8_755 = $signed(_T_69707); // @[Modules.scala 78:156:@21167.4]
  assign _T_69709 = $signed(buffer_8_755) + $signed(buffer_8_707); // @[Modules.scala 78:156:@21169.4]
  assign _T_69710 = _T_69709[10:0]; // @[Modules.scala 78:156:@21170.4]
  assign buffer_8_756 = $signed(_T_69710); // @[Modules.scala 78:156:@21171.4]
  assign _T_69712 = $signed(buffer_8_756) + $signed(buffer_8_708); // @[Modules.scala 78:156:@21173.4]
  assign _T_69713 = _T_69712[10:0]; // @[Modules.scala 78:156:@21174.4]
  assign buffer_8_757 = $signed(_T_69713); // @[Modules.scala 78:156:@21175.4]
  assign _T_69715 = $signed(buffer_8_757) + $signed(buffer_8_709); // @[Modules.scala 78:156:@21177.4]
  assign _T_69716 = _T_69715[10:0]; // @[Modules.scala 78:156:@21178.4]
  assign buffer_8_758 = $signed(_T_69716); // @[Modules.scala 78:156:@21179.4]
  assign _T_69718 = $signed(buffer_8_758) + $signed(buffer_8_710); // @[Modules.scala 78:156:@21181.4]
  assign _T_69719 = _T_69718[10:0]; // @[Modules.scala 78:156:@21182.4]
  assign buffer_8_759 = $signed(_T_69719); // @[Modules.scala 78:156:@21183.4]
  assign _T_69721 = $signed(buffer_8_759) + $signed(buffer_8_711); // @[Modules.scala 78:156:@21185.4]
  assign _T_69722 = _T_69721[10:0]; // @[Modules.scala 78:156:@21186.4]
  assign buffer_8_760 = $signed(_T_69722); // @[Modules.scala 78:156:@21187.4]
  assign _T_69724 = $signed(buffer_8_760) + $signed(buffer_8_712); // @[Modules.scala 78:156:@21189.4]
  assign _T_69725 = _T_69724[10:0]; // @[Modules.scala 78:156:@21190.4]
  assign buffer_8_761 = $signed(_T_69725); // @[Modules.scala 78:156:@21191.4]
  assign _T_69727 = $signed(buffer_8_761) + $signed(buffer_8_713); // @[Modules.scala 78:156:@21193.4]
  assign _T_69728 = _T_69727[10:0]; // @[Modules.scala 78:156:@21194.4]
  assign buffer_8_762 = $signed(_T_69728); // @[Modules.scala 78:156:@21195.4]
  assign _T_69730 = $signed(buffer_8_762) + $signed(buffer_8_714); // @[Modules.scala 78:156:@21197.4]
  assign _T_69731 = _T_69730[10:0]; // @[Modules.scala 78:156:@21198.4]
  assign buffer_8_763 = $signed(_T_69731); // @[Modules.scala 78:156:@21199.4]
  assign _T_69733 = $signed(buffer_8_763) + $signed(buffer_8_715); // @[Modules.scala 78:156:@21201.4]
  assign _T_69734 = _T_69733[10:0]; // @[Modules.scala 78:156:@21202.4]
  assign buffer_8_764 = $signed(_T_69734); // @[Modules.scala 78:156:@21203.4]
  assign _T_69736 = $signed(buffer_8_764) + $signed(buffer_8_716); // @[Modules.scala 78:156:@21205.4]
  assign _T_69737 = _T_69736[10:0]; // @[Modules.scala 78:156:@21206.4]
  assign buffer_8_765 = $signed(_T_69737); // @[Modules.scala 78:156:@21207.4]
  assign _T_69739 = $signed(buffer_8_765) + $signed(buffer_8_717); // @[Modules.scala 78:156:@21209.4]
  assign _T_69740 = _T_69739[10:0]; // @[Modules.scala 78:156:@21210.4]
  assign buffer_8_766 = $signed(_T_69740); // @[Modules.scala 78:156:@21211.4]
  assign _T_69742 = $signed(buffer_8_766) + $signed(buffer_8_718); // @[Modules.scala 78:156:@21213.4]
  assign _T_69743 = _T_69742[10:0]; // @[Modules.scala 78:156:@21214.4]
  assign buffer_8_767 = $signed(_T_69743); // @[Modules.scala 78:156:@21215.4]
  assign _T_69745 = $signed(buffer_8_767) + $signed(buffer_8_719); // @[Modules.scala 78:156:@21217.4]
  assign _T_69746 = _T_69745[10:0]; // @[Modules.scala 78:156:@21218.4]
  assign buffer_8_768 = $signed(_T_69746); // @[Modules.scala 78:156:@21219.4]
  assign _T_69748 = $signed(buffer_8_768) + $signed(buffer_8_720); // @[Modules.scala 78:156:@21221.4]
  assign _T_69749 = _T_69748[10:0]; // @[Modules.scala 78:156:@21222.4]
  assign buffer_8_769 = $signed(_T_69749); // @[Modules.scala 78:156:@21223.4]
  assign _T_69751 = $signed(buffer_8_769) + $signed(buffer_8_721); // @[Modules.scala 78:156:@21225.4]
  assign _T_69752 = _T_69751[10:0]; // @[Modules.scala 78:156:@21226.4]
  assign buffer_8_770 = $signed(_T_69752); // @[Modules.scala 78:156:@21227.4]
  assign _T_69754 = $signed(buffer_8_770) + $signed(buffer_8_722); // @[Modules.scala 78:156:@21229.4]
  assign _T_69755 = _T_69754[10:0]; // @[Modules.scala 78:156:@21230.4]
  assign buffer_8_771 = $signed(_T_69755); // @[Modules.scala 78:156:@21231.4]
  assign _T_69757 = $signed(buffer_8_771) + $signed(buffer_8_723); // @[Modules.scala 78:156:@21233.4]
  assign _T_69758 = _T_69757[10:0]; // @[Modules.scala 78:156:@21234.4]
  assign buffer_8_772 = $signed(_T_69758); // @[Modules.scala 78:156:@21235.4]
  assign _T_69760 = $signed(buffer_8_772) + $signed(buffer_8_724); // @[Modules.scala 78:156:@21237.4]
  assign _T_69761 = _T_69760[10:0]; // @[Modules.scala 78:156:@21238.4]
  assign buffer_8_773 = $signed(_T_69761); // @[Modules.scala 78:156:@21239.4]
  assign _T_69763 = $signed(buffer_8_773) + $signed(buffer_8_725); // @[Modules.scala 78:156:@21241.4]
  assign _T_69764 = _T_69763[10:0]; // @[Modules.scala 78:156:@21242.4]
  assign buffer_8_774 = $signed(_T_69764); // @[Modules.scala 78:156:@21243.4]
  assign _T_69766 = $signed(buffer_8_774) + $signed(buffer_8_726); // @[Modules.scala 78:156:@21245.4]
  assign _T_69767 = _T_69766[10:0]; // @[Modules.scala 78:156:@21246.4]
  assign buffer_8_775 = $signed(_T_69767); // @[Modules.scala 78:156:@21247.4]
  assign _T_69769 = $signed(buffer_8_775) + $signed(buffer_8_727); // @[Modules.scala 78:156:@21249.4]
  assign _T_69770 = _T_69769[10:0]; // @[Modules.scala 78:156:@21250.4]
  assign buffer_8_776 = $signed(_T_69770); // @[Modules.scala 78:156:@21251.4]
  assign _T_69772 = $signed(buffer_8_776) + $signed(buffer_8_728); // @[Modules.scala 78:156:@21253.4]
  assign _T_69773 = _T_69772[10:0]; // @[Modules.scala 78:156:@21254.4]
  assign buffer_8_777 = $signed(_T_69773); // @[Modules.scala 78:156:@21255.4]
  assign _T_69775 = $signed(buffer_8_777) + $signed(buffer_8_729); // @[Modules.scala 78:156:@21257.4]
  assign _T_69776 = _T_69775[10:0]; // @[Modules.scala 78:156:@21258.4]
  assign buffer_8_778 = $signed(_T_69776); // @[Modules.scala 78:156:@21259.4]
  assign _T_69778 = $signed(buffer_8_778) + $signed(buffer_0_701); // @[Modules.scala 78:156:@21261.4]
  assign _T_69779 = _T_69778[10:0]; // @[Modules.scala 78:156:@21262.4]
  assign buffer_8_779 = $signed(_T_69779); // @[Modules.scala 78:156:@21263.4]
  assign _T_69781 = $signed(buffer_8_779) + $signed(buffer_8_731); // @[Modules.scala 78:156:@21265.4]
  assign _T_69782 = _T_69781[10:0]; // @[Modules.scala 78:156:@21266.4]
  assign buffer_8_780 = $signed(_T_69782); // @[Modules.scala 78:156:@21267.4]
  assign _T_69784 = $signed(buffer_8_780) + $signed(buffer_0_701); // @[Modules.scala 78:156:@21269.4]
  assign _T_69785 = _T_69784[10:0]; // @[Modules.scala 78:156:@21270.4]
  assign buffer_8_781 = $signed(_T_69785); // @[Modules.scala 78:156:@21271.4]
  assign _T_69787 = $signed(buffer_8_781) + $signed(buffer_8_733); // @[Modules.scala 78:156:@21273.4]
  assign _T_69788 = _T_69787[10:0]; // @[Modules.scala 78:156:@21274.4]
  assign buffer_8_782 = $signed(_T_69788); // @[Modules.scala 78:156:@21275.4]
  assign _T_69790 = $signed(buffer_8_782) + $signed(buffer_8_734); // @[Modules.scala 78:156:@21277.4]
  assign _T_69791 = _T_69790[10:0]; // @[Modules.scala 78:156:@21278.4]
  assign buffer_8_783 = $signed(_T_69791); // @[Modules.scala 78:156:@21279.4]
  assign _T_69794 = $signed(io_in_2) + $signed(io_in_3); // @[Modules.scala 37:46:@21283.4]
  assign _T_69795 = _T_69794[4:0]; // @[Modules.scala 37:46:@21284.4]
  assign _T_69796 = $signed(_T_69795); // @[Modules.scala 37:46:@21285.4]
  assign _T_69803 = $signed(io_in_18) + $signed(io_in_19); // @[Modules.scala 37:46:@21294.4]
  assign _T_69804 = _T_69803[4:0]; // @[Modules.scala 37:46:@21295.4]
  assign _T_69805 = $signed(_T_69804); // @[Modules.scala 37:46:@21296.4]
  assign buffer_9_1 = {{6{_T_69796[4]}},_T_69796}; // @[Modules.scala 32:22:@8.4]
  assign _T_70417 = $signed(11'sh0) + $signed(buffer_9_1); // @[Modules.scala 65:57:@22199.4]
  assign _T_70418 = _T_70417[10:0]; // @[Modules.scala 65:57:@22200.4]
  assign buffer_9_392 = $signed(_T_70418); // @[Modules.scala 65:57:@22201.4]
  assign _T_70420 = $signed(11'sh0) + $signed(buffer_0_3); // @[Modules.scala 65:57:@22203.4]
  assign _T_70421 = _T_70420[10:0]; // @[Modules.scala 65:57:@22204.4]
  assign buffer_9_393 = $signed(_T_70421); // @[Modules.scala 65:57:@22205.4]
  assign buffer_9_9 = {{6{_T_69805[4]}},_T_69805}; // @[Modules.scala 32:22:@8.4]
  assign _T_70429 = $signed(11'sh0) + $signed(buffer_9_9); // @[Modules.scala 65:57:@22215.4]
  assign _T_70430 = _T_70429[10:0]; // @[Modules.scala 65:57:@22216.4]
  assign buffer_9_396 = $signed(_T_70430); // @[Modules.scala 65:57:@22217.4]
  assign _T_70435 = $signed(buffer_3_12) + $signed(11'sh0); // @[Modules.scala 65:57:@22223.4]
  assign _T_70436 = _T_70435[10:0]; // @[Modules.scala 65:57:@22224.4]
  assign buffer_9_398 = $signed(_T_70436); // @[Modules.scala 65:57:@22225.4]
  assign _T_70450 = $signed(buffer_4_22) + $signed(buffer_1_23); // @[Modules.scala 65:57:@22243.4]
  assign _T_70451 = _T_70450[10:0]; // @[Modules.scala 65:57:@22244.4]
  assign buffer_9_403 = $signed(_T_70451); // @[Modules.scala 65:57:@22245.4]
  assign buffer_9_41 = {{6{io_in_83[4]}},io_in_83}; // @[Modules.scala 32:22:@8.4]
  assign _T_70477 = $signed(buffer_1_40) + $signed(buffer_9_41); // @[Modules.scala 65:57:@22279.4]
  assign _T_70478 = _T_70477[10:0]; // @[Modules.scala 65:57:@22280.4]
  assign buffer_9_412 = $signed(_T_70478); // @[Modules.scala 65:57:@22281.4]
  assign _T_70501 = $signed(buffer_0_56) + $signed(buffer_3_57); // @[Modules.scala 65:57:@22311.4]
  assign _T_70502 = _T_70501[10:0]; // @[Modules.scala 65:57:@22312.4]
  assign buffer_9_420 = $signed(_T_70502); // @[Modules.scala 65:57:@22313.4]
  assign _T_70519 = $signed(11'sh0) + $signed(buffer_4_69); // @[Modules.scala 65:57:@22335.4]
  assign _T_70520 = _T_70519[10:0]; // @[Modules.scala 65:57:@22336.4]
  assign buffer_9_426 = $signed(_T_70520); // @[Modules.scala 65:57:@22337.4]
  assign buffer_9_75 = {{6{io_in_151[4]}},io_in_151}; // @[Modules.scala 32:22:@8.4]
  assign _T_70528 = $signed(buffer_0_74) + $signed(buffer_9_75); // @[Modules.scala 65:57:@22347.4]
  assign _T_70529 = _T_70528[10:0]; // @[Modules.scala 65:57:@22348.4]
  assign buffer_9_429 = $signed(_T_70529); // @[Modules.scala 65:57:@22349.4]
  assign _T_70531 = $signed(buffer_7_76) + $signed(11'sh0); // @[Modules.scala 65:57:@22351.4]
  assign _T_70532 = _T_70531[10:0]; // @[Modules.scala 65:57:@22352.4]
  assign buffer_9_430 = $signed(_T_70532); // @[Modules.scala 65:57:@22353.4]
  assign buffer_9_78 = {{6{io_in_157[4]}},io_in_157}; // @[Modules.scala 32:22:@8.4]
  assign _T_70534 = $signed(buffer_9_78) + $signed(buffer_2_79); // @[Modules.scala 65:57:@22355.4]
  assign _T_70535 = _T_70534[10:0]; // @[Modules.scala 65:57:@22356.4]
  assign buffer_9_431 = $signed(_T_70535); // @[Modules.scala 65:57:@22357.4]
  assign buffer_9_85 = {{6{io_in_171[4]}},io_in_171}; // @[Modules.scala 32:22:@8.4]
  assign _T_70543 = $signed(buffer_4_84) + $signed(buffer_9_85); // @[Modules.scala 65:57:@22367.4]
  assign _T_70544 = _T_70543[10:0]; // @[Modules.scala 65:57:@22368.4]
  assign buffer_9_434 = $signed(_T_70544); // @[Modules.scala 65:57:@22369.4]
  assign buffer_9_91 = {{6{io_in_183[4]}},io_in_183}; // @[Modules.scala 32:22:@8.4]
  assign _T_70552 = $signed(buffer_3_90) + $signed(buffer_9_91); // @[Modules.scala 65:57:@22379.4]
  assign _T_70553 = _T_70552[10:0]; // @[Modules.scala 65:57:@22380.4]
  assign buffer_9_437 = $signed(_T_70553); // @[Modules.scala 65:57:@22381.4]
  assign _T_70561 = $signed(buffer_1_96) + $signed(buffer_2_97); // @[Modules.scala 65:57:@22391.4]
  assign _T_70562 = _T_70561[10:0]; // @[Modules.scala 65:57:@22392.4]
  assign buffer_9_440 = $signed(_T_70562); // @[Modules.scala 65:57:@22393.4]
  assign _T_70570 = $signed(buffer_4_102) + $signed(11'sh0); // @[Modules.scala 65:57:@22403.4]
  assign _T_70571 = _T_70570[10:0]; // @[Modules.scala 65:57:@22404.4]
  assign buffer_9_443 = $signed(_T_70571); // @[Modules.scala 65:57:@22405.4]
  assign _T_70576 = $signed(buffer_1_106) + $signed(11'sh0); // @[Modules.scala 65:57:@22411.4]
  assign _T_70577 = _T_70576[10:0]; // @[Modules.scala 65:57:@22412.4]
  assign buffer_9_445 = $signed(_T_70577); // @[Modules.scala 65:57:@22413.4]
  assign _T_70579 = $signed(buffer_7_108) + $signed(11'sh0); // @[Modules.scala 65:57:@22415.4]
  assign _T_70580 = _T_70579[10:0]; // @[Modules.scala 65:57:@22416.4]
  assign buffer_9_446 = $signed(_T_70580); // @[Modules.scala 65:57:@22417.4]
  assign _T_70582 = $signed(11'sh0) + $signed(buffer_2_111); // @[Modules.scala 65:57:@22419.4]
  assign _T_70583 = _T_70582[10:0]; // @[Modules.scala 65:57:@22420.4]
  assign buffer_9_447 = $signed(_T_70583); // @[Modules.scala 65:57:@22421.4]
  assign _T_70585 = $signed(buffer_1_112) + $signed(buffer_5_113); // @[Modules.scala 65:57:@22423.4]
  assign _T_70586 = _T_70585[10:0]; // @[Modules.scala 65:57:@22424.4]
  assign buffer_9_448 = $signed(_T_70586); // @[Modules.scala 65:57:@22425.4]
  assign buffer_9_114 = {{6{io_in_228[4]}},io_in_228}; // @[Modules.scala 32:22:@8.4]
  assign _T_70588 = $signed(buffer_9_114) + $signed(buffer_8_115); // @[Modules.scala 65:57:@22427.4]
  assign _T_70589 = _T_70588[10:0]; // @[Modules.scala 65:57:@22428.4]
  assign buffer_9_449 = $signed(_T_70589); // @[Modules.scala 65:57:@22429.4]
  assign _T_70594 = $signed(buffer_0_118) + $signed(buffer_3_119); // @[Modules.scala 65:57:@22435.4]
  assign _T_70595 = _T_70594[10:0]; // @[Modules.scala 65:57:@22436.4]
  assign buffer_9_451 = $signed(_T_70595); // @[Modules.scala 65:57:@22437.4]
  assign buffer_9_122 = {{6{io_in_245[4]}},io_in_245}; // @[Modules.scala 32:22:@8.4]
  assign _T_70600 = $signed(buffer_9_122) + $signed(11'sh0); // @[Modules.scala 65:57:@22443.4]
  assign _T_70601 = _T_70600[10:0]; // @[Modules.scala 65:57:@22444.4]
  assign buffer_9_453 = $signed(_T_70601); // @[Modules.scala 65:57:@22445.4]
  assign _T_70609 = $signed(buffer_8_128) + $signed(buffer_4_129); // @[Modules.scala 65:57:@22455.4]
  assign _T_70610 = _T_70609[10:0]; // @[Modules.scala 65:57:@22456.4]
  assign buffer_9_456 = $signed(_T_70610); // @[Modules.scala 65:57:@22457.4]
  assign buffer_9_133 = {{6{io_in_266[4]}},io_in_266}; // @[Modules.scala 32:22:@8.4]
  assign _T_70615 = $signed(11'sh0) + $signed(buffer_9_133); // @[Modules.scala 65:57:@22463.4]
  assign _T_70616 = _T_70615[10:0]; // @[Modules.scala 65:57:@22464.4]
  assign buffer_9_458 = $signed(_T_70616); // @[Modules.scala 65:57:@22465.4]
  assign _T_70624 = $signed(11'sh0) + $signed(buffer_1_139); // @[Modules.scala 65:57:@22475.4]
  assign _T_70625 = _T_70624[10:0]; // @[Modules.scala 65:57:@22476.4]
  assign buffer_9_461 = $signed(_T_70625); // @[Modules.scala 65:57:@22477.4]
  assign _T_70627 = $signed(buffer_3_140) + $signed(buffer_1_141); // @[Modules.scala 65:57:@22479.4]
  assign _T_70628 = _T_70627[10:0]; // @[Modules.scala 65:57:@22480.4]
  assign buffer_9_462 = $signed(_T_70628); // @[Modules.scala 65:57:@22481.4]
  assign _T_70630 = $signed(buffer_3_142) + $signed(buffer_5_143); // @[Modules.scala 65:57:@22483.4]
  assign _T_70631 = _T_70630[10:0]; // @[Modules.scala 65:57:@22484.4]
  assign buffer_9_463 = $signed(_T_70631); // @[Modules.scala 65:57:@22485.4]
  assign _T_70642 = $signed(buffer_6_150) + $signed(buffer_4_151); // @[Modules.scala 65:57:@22499.4]
  assign _T_70643 = _T_70642[10:0]; // @[Modules.scala 65:57:@22500.4]
  assign buffer_9_467 = $signed(_T_70643); // @[Modules.scala 65:57:@22501.4]
  assign buffer_9_152 = {{6{io_in_304[4]}},io_in_304}; // @[Modules.scala 32:22:@8.4]
  assign _T_70645 = $signed(buffer_9_152) + $signed(buffer_5_153); // @[Modules.scala 65:57:@22503.4]
  assign _T_70646 = _T_70645[10:0]; // @[Modules.scala 65:57:@22504.4]
  assign buffer_9_468 = $signed(_T_70646); // @[Modules.scala 65:57:@22505.4]
  assign buffer_9_156 = {{6{io_in_312[4]}},io_in_312}; // @[Modules.scala 32:22:@8.4]
  assign _T_70651 = $signed(buffer_9_156) + $signed(11'sh0); // @[Modules.scala 65:57:@22511.4]
  assign _T_70652 = _T_70651[10:0]; // @[Modules.scala 65:57:@22512.4]
  assign buffer_9_470 = $signed(_T_70652); // @[Modules.scala 65:57:@22513.4]
  assign buffer_9_160 = {{6{io_in_321[4]}},io_in_321}; // @[Modules.scala 32:22:@8.4]
  assign _T_70657 = $signed(buffer_9_160) + $signed(buffer_5_161); // @[Modules.scala 65:57:@22519.4]
  assign _T_70658 = _T_70657[10:0]; // @[Modules.scala 65:57:@22520.4]
  assign buffer_9_472 = $signed(_T_70658); // @[Modules.scala 65:57:@22521.4]
  assign buffer_9_174 = {{6{io_in_349[4]}},io_in_349}; // @[Modules.scala 32:22:@8.4]
  assign _T_70678 = $signed(buffer_9_174) + $signed(buffer_0_175); // @[Modules.scala 65:57:@22547.4]
  assign _T_70679 = _T_70678[10:0]; // @[Modules.scala 65:57:@22548.4]
  assign buffer_9_479 = $signed(_T_70679); // @[Modules.scala 65:57:@22549.4]
  assign _T_70681 = $signed(11'sh0) + $signed(buffer_0_177); // @[Modules.scala 65:57:@22551.4]
  assign _T_70682 = _T_70681[10:0]; // @[Modules.scala 65:57:@22552.4]
  assign buffer_9_480 = $signed(_T_70682); // @[Modules.scala 65:57:@22553.4]
  assign _T_70684 = $signed(buffer_0_178) + $signed(11'sh0); // @[Modules.scala 65:57:@22555.4]
  assign _T_70685 = _T_70684[10:0]; // @[Modules.scala 65:57:@22556.4]
  assign buffer_9_481 = $signed(_T_70685); // @[Modules.scala 65:57:@22557.4]
  assign buffer_9_191 = {{6{io_in_382[4]}},io_in_382}; // @[Modules.scala 32:22:@8.4]
  assign _T_70702 = $signed(buffer_4_190) + $signed(buffer_9_191); // @[Modules.scala 65:57:@22579.4]
  assign _T_70703 = _T_70702[10:0]; // @[Modules.scala 65:57:@22580.4]
  assign buffer_9_487 = $signed(_T_70703); // @[Modules.scala 65:57:@22581.4]
  assign _T_70708 = $signed(buffer_4_194) + $signed(buffer_3_195); // @[Modules.scala 65:57:@22587.4]
  assign _T_70709 = _T_70708[10:0]; // @[Modules.scala 65:57:@22588.4]
  assign buffer_9_489 = $signed(_T_70709); // @[Modules.scala 65:57:@22589.4]
  assign _T_70711 = $signed(buffer_6_196) + $signed(buffer_3_197); // @[Modules.scala 65:57:@22591.4]
  assign _T_70712 = _T_70711[10:0]; // @[Modules.scala 65:57:@22592.4]
  assign buffer_9_490 = $signed(_T_70712); // @[Modules.scala 65:57:@22593.4]
  assign buffer_9_200 = {{6{io_in_400[4]}},io_in_400}; // @[Modules.scala 32:22:@8.4]
  assign _T_70717 = $signed(buffer_9_200) + $signed(11'sh0); // @[Modules.scala 65:57:@22599.4]
  assign _T_70718 = _T_70717[10:0]; // @[Modules.scala 65:57:@22600.4]
  assign buffer_9_492 = $signed(_T_70718); // @[Modules.scala 65:57:@22601.4]
  assign _T_70738 = $signed(11'sh0) + $signed(buffer_6_215); // @[Modules.scala 65:57:@22627.4]
  assign _T_70739 = _T_70738[10:0]; // @[Modules.scala 65:57:@22628.4]
  assign buffer_9_499 = $signed(_T_70739); // @[Modules.scala 65:57:@22629.4]
  assign _T_70753 = $signed(buffer_0_224) + $signed(buffer_1_225); // @[Modules.scala 65:57:@22647.4]
  assign _T_70754 = _T_70753[10:0]; // @[Modules.scala 65:57:@22648.4]
  assign buffer_9_504 = $signed(_T_70754); // @[Modules.scala 65:57:@22649.4]
  assign buffer_9_226 = {{6{io_in_452[4]}},io_in_452}; // @[Modules.scala 32:22:@8.4]
  assign _T_70756 = $signed(buffer_9_226) + $signed(11'sh0); // @[Modules.scala 65:57:@22651.4]
  assign _T_70757 = _T_70756[10:0]; // @[Modules.scala 65:57:@22652.4]
  assign buffer_9_505 = $signed(_T_70757); // @[Modules.scala 65:57:@22653.4]
  assign _T_70759 = $signed(11'sh0) + $signed(buffer_6_229); // @[Modules.scala 65:57:@22655.4]
  assign _T_70760 = _T_70759[10:0]; // @[Modules.scala 65:57:@22656.4]
  assign buffer_9_506 = $signed(_T_70760); // @[Modules.scala 65:57:@22657.4]
  assign _T_70777 = $signed(buffer_7_240) + $signed(11'sh0); // @[Modules.scala 65:57:@22679.4]
  assign _T_70778 = _T_70777[10:0]; // @[Modules.scala 65:57:@22680.4]
  assign buffer_9_512 = $signed(_T_70778); // @[Modules.scala 65:57:@22681.4]
  assign buffer_9_245 = {{6{io_in_490[4]}},io_in_490}; // @[Modules.scala 32:22:@8.4]
  assign _T_70783 = $signed(buffer_2_244) + $signed(buffer_9_245); // @[Modules.scala 65:57:@22687.4]
  assign _T_70784 = _T_70783[10:0]; // @[Modules.scala 65:57:@22688.4]
  assign buffer_9_514 = $signed(_T_70784); // @[Modules.scala 65:57:@22689.4]
  assign _T_70798 = $signed(buffer_3_254) + $signed(11'sh0); // @[Modules.scala 65:57:@22707.4]
  assign _T_70799 = _T_70798[10:0]; // @[Modules.scala 65:57:@22708.4]
  assign buffer_9_519 = $signed(_T_70799); // @[Modules.scala 65:57:@22709.4]
  assign _T_70819 = $signed(buffer_1_268) + $signed(buffer_5_269); // @[Modules.scala 65:57:@22735.4]
  assign _T_70820 = _T_70819[10:0]; // @[Modules.scala 65:57:@22736.4]
  assign buffer_9_526 = $signed(_T_70820); // @[Modules.scala 65:57:@22737.4]
  assign buffer_9_283 = {{6{io_in_567[4]}},io_in_567}; // @[Modules.scala 32:22:@8.4]
  assign _T_70840 = $signed(buffer_1_282) + $signed(buffer_9_283); // @[Modules.scala 65:57:@22763.4]
  assign _T_70841 = _T_70840[10:0]; // @[Modules.scala 65:57:@22764.4]
  assign buffer_9_533 = $signed(_T_70841); // @[Modules.scala 65:57:@22765.4]
  assign _T_70843 = $signed(buffer_8_284) + $signed(buffer_1_285); // @[Modules.scala 65:57:@22767.4]
  assign _T_70844 = _T_70843[10:0]; // @[Modules.scala 65:57:@22768.4]
  assign buffer_9_534 = $signed(_T_70844); // @[Modules.scala 65:57:@22769.4]
  assign _T_70846 = $signed(buffer_3_286) + $signed(buffer_1_287); // @[Modules.scala 65:57:@22771.4]
  assign _T_70847 = _T_70846[10:0]; // @[Modules.scala 65:57:@22772.4]
  assign buffer_9_535 = $signed(_T_70847); // @[Modules.scala 65:57:@22773.4]
  assign _T_70864 = $signed(buffer_1_298) + $signed(buffer_2_299); // @[Modules.scala 65:57:@22795.4]
  assign _T_70865 = _T_70864[10:0]; // @[Modules.scala 65:57:@22796.4]
  assign buffer_9_541 = $signed(_T_70865); // @[Modules.scala 65:57:@22797.4]
  assign buffer_9_300 = {{6{io_in_600[4]}},io_in_600}; // @[Modules.scala 32:22:@8.4]
  assign _T_70867 = $signed(buffer_9_300) + $signed(buffer_0_301); // @[Modules.scala 65:57:@22799.4]
  assign _T_70868 = _T_70867[10:0]; // @[Modules.scala 65:57:@22800.4]
  assign buffer_9_542 = $signed(_T_70868); // @[Modules.scala 65:57:@22801.4]
  assign buffer_9_304 = {{6{io_in_608[4]}},io_in_608}; // @[Modules.scala 32:22:@8.4]
  assign buffer_9_305 = {{6{io_in_611[4]}},io_in_611}; // @[Modules.scala 32:22:@8.4]
  assign _T_70873 = $signed(buffer_9_304) + $signed(buffer_9_305); // @[Modules.scala 65:57:@22807.4]
  assign _T_70874 = _T_70873[10:0]; // @[Modules.scala 65:57:@22808.4]
  assign buffer_9_544 = $signed(_T_70874); // @[Modules.scala 65:57:@22809.4]
  assign _T_70885 = $signed(buffer_1_312) + $signed(buffer_5_313); // @[Modules.scala 65:57:@22823.4]
  assign _T_70886 = _T_70885[10:0]; // @[Modules.scala 65:57:@22824.4]
  assign buffer_9_548 = $signed(_T_70886); // @[Modules.scala 65:57:@22825.4]
  assign _T_70891 = $signed(buffer_4_316) + $signed(11'sh0); // @[Modules.scala 65:57:@22831.4]
  assign _T_70892 = _T_70891[10:0]; // @[Modules.scala 65:57:@22832.4]
  assign buffer_9_550 = $signed(_T_70892); // @[Modules.scala 65:57:@22833.4]
  assign _T_70894 = $signed(buffer_1_318) + $signed(buffer_0_319); // @[Modules.scala 65:57:@22835.4]
  assign _T_70895 = _T_70894[10:0]; // @[Modules.scala 65:57:@22836.4]
  assign buffer_9_551 = $signed(_T_70895); // @[Modules.scala 65:57:@22837.4]
  assign buffer_9_320 = {{6{io_in_641[4]}},io_in_641}; // @[Modules.scala 32:22:@8.4]
  assign _T_70897 = $signed(buffer_9_320) + $signed(buffer_3_321); // @[Modules.scala 65:57:@22839.4]
  assign _T_70898 = _T_70897[10:0]; // @[Modules.scala 65:57:@22840.4]
  assign buffer_9_552 = $signed(_T_70898); // @[Modules.scala 65:57:@22841.4]
  assign _T_70906 = $signed(buffer_1_326) + $signed(buffer_8_327); // @[Modules.scala 65:57:@22851.4]
  assign _T_70907 = _T_70906[10:0]; // @[Modules.scala 65:57:@22852.4]
  assign buffer_9_555 = $signed(_T_70907); // @[Modules.scala 65:57:@22853.4]
  assign _T_70915 = $signed(buffer_5_332) + $signed(11'sh0); // @[Modules.scala 65:57:@22863.4]
  assign _T_70916 = _T_70915[10:0]; // @[Modules.scala 65:57:@22864.4]
  assign buffer_9_558 = $signed(_T_70916); // @[Modules.scala 65:57:@22865.4]
  assign buffer_9_346 = {{6{io_in_693[4]}},io_in_693}; // @[Modules.scala 32:22:@8.4]
  assign buffer_9_347 = {{6{io_in_694[4]}},io_in_694}; // @[Modules.scala 32:22:@8.4]
  assign _T_70936 = $signed(buffer_9_346) + $signed(buffer_9_347); // @[Modules.scala 65:57:@22891.4]
  assign _T_70937 = _T_70936[10:0]; // @[Modules.scala 65:57:@22892.4]
  assign buffer_9_565 = $signed(_T_70937); // @[Modules.scala 65:57:@22893.4]
  assign _T_70939 = $signed(buffer_0_348) + $signed(buffer_3_349); // @[Modules.scala 65:57:@22895.4]
  assign _T_70940 = _T_70939[10:0]; // @[Modules.scala 65:57:@22896.4]
  assign buffer_9_566 = $signed(_T_70940); // @[Modules.scala 65:57:@22897.4]
  assign _T_70942 = $signed(buffer_5_350) + $signed(buffer_0_351); // @[Modules.scala 65:57:@22899.4]
  assign _T_70943 = _T_70942[10:0]; // @[Modules.scala 65:57:@22900.4]
  assign buffer_9_567 = $signed(_T_70943); // @[Modules.scala 65:57:@22901.4]
  assign buffer_9_354 = {{6{io_in_708[4]}},io_in_708}; // @[Modules.scala 32:22:@8.4]
  assign _T_70948 = $signed(buffer_9_354) + $signed(11'sh0); // @[Modules.scala 65:57:@22907.4]
  assign _T_70949 = _T_70948[10:0]; // @[Modules.scala 65:57:@22908.4]
  assign buffer_9_569 = $signed(_T_70949); // @[Modules.scala 65:57:@22909.4]
  assign buffer_9_356 = {{6{io_in_712[4]}},io_in_712}; // @[Modules.scala 32:22:@8.4]
  assign _T_70951 = $signed(buffer_9_356) + $signed(11'sh0); // @[Modules.scala 65:57:@22911.4]
  assign _T_70952 = _T_70951[10:0]; // @[Modules.scala 65:57:@22912.4]
  assign buffer_9_570 = $signed(_T_70952); // @[Modules.scala 65:57:@22913.4]
  assign buffer_9_358 = {{6{io_in_717[4]}},io_in_717}; // @[Modules.scala 32:22:@8.4]
  assign _T_70954 = $signed(buffer_9_358) + $signed(buffer_6_359); // @[Modules.scala 65:57:@22915.4]
  assign _T_70955 = _T_70954[10:0]; // @[Modules.scala 65:57:@22916.4]
  assign buffer_9_571 = $signed(_T_70955); // @[Modules.scala 65:57:@22917.4]
  assign buffer_9_362 = {{6{io_in_725[4]}},io_in_725}; // @[Modules.scala 32:22:@8.4]
  assign _T_70960 = $signed(buffer_9_362) + $signed(buffer_1_363); // @[Modules.scala 65:57:@22923.4]
  assign _T_70961 = _T_70960[10:0]; // @[Modules.scala 65:57:@22924.4]
  assign buffer_9_573 = $signed(_T_70961); // @[Modules.scala 65:57:@22925.4]
  assign buffer_9_364 = {{6{io_in_729[4]}},io_in_729}; // @[Modules.scala 32:22:@8.4]
  assign _T_70963 = $signed(buffer_9_364) + $signed(buffer_3_365); // @[Modules.scala 65:57:@22927.4]
  assign _T_70964 = _T_70963[10:0]; // @[Modules.scala 65:57:@22928.4]
  assign buffer_9_574 = $signed(_T_70964); // @[Modules.scala 65:57:@22929.4]
  assign _T_70975 = $signed(11'sh0) + $signed(buffer_3_373); // @[Modules.scala 65:57:@22943.4]
  assign _T_70976 = _T_70975[10:0]; // @[Modules.scala 65:57:@22944.4]
  assign buffer_9_578 = $signed(_T_70976); // @[Modules.scala 65:57:@22945.4]
  assign _T_70978 = $signed(buffer_0_374) + $signed(buffer_2_375); // @[Modules.scala 65:57:@22947.4]
  assign _T_70979 = _T_70978[10:0]; // @[Modules.scala 65:57:@22948.4]
  assign buffer_9_579 = $signed(_T_70979); // @[Modules.scala 65:57:@22949.4]
  assign _T_70981 = $signed(buffer_0_376) + $signed(11'sh0); // @[Modules.scala 65:57:@22951.4]
  assign _T_70982 = _T_70981[10:0]; // @[Modules.scala 65:57:@22952.4]
  assign buffer_9_580 = $signed(_T_70982); // @[Modules.scala 65:57:@22953.4]
  assign buffer_9_379 = {{6{io_in_758[4]}},io_in_758}; // @[Modules.scala 32:22:@8.4]
  assign _T_70984 = $signed(buffer_3_378) + $signed(buffer_9_379); // @[Modules.scala 65:57:@22955.4]
  assign _T_70985 = _T_70984[10:0]; // @[Modules.scala 65:57:@22956.4]
  assign buffer_9_581 = $signed(_T_70985); // @[Modules.scala 65:57:@22957.4]
  assign buffer_9_381 = {{6{io_in_763[4]}},io_in_763}; // @[Modules.scala 32:22:@8.4]
  assign _T_70987 = $signed(11'sh0) + $signed(buffer_9_381); // @[Modules.scala 65:57:@22959.4]
  assign _T_70988 = _T_70987[10:0]; // @[Modules.scala 65:57:@22960.4]
  assign buffer_9_582 = $signed(_T_70988); // @[Modules.scala 65:57:@22961.4]
  assign _T_70990 = $signed(buffer_3_382) + $signed(buffer_4_383); // @[Modules.scala 65:57:@22963.4]
  assign _T_70991 = _T_70990[10:0]; // @[Modules.scala 65:57:@22964.4]
  assign buffer_9_583 = $signed(_T_70991); // @[Modules.scala 65:57:@22965.4]
  assign buffer_9_387 = {{6{io_in_774[4]}},io_in_774}; // @[Modules.scala 32:22:@8.4]
  assign _T_70996 = $signed(buffer_3_386) + $signed(buffer_9_387); // @[Modules.scala 65:57:@22971.4]
  assign _T_70997 = _T_70996[10:0]; // @[Modules.scala 65:57:@22972.4]
  assign buffer_9_585 = $signed(_T_70997); // @[Modules.scala 65:57:@22973.4]
  assign _T_71005 = $signed(buffer_9_392) + $signed(buffer_9_393); // @[Modules.scala 68:83:@22983.4]
  assign _T_71006 = _T_71005[10:0]; // @[Modules.scala 68:83:@22984.4]
  assign buffer_9_588 = $signed(_T_71006); // @[Modules.scala 68:83:@22985.4]
  assign _T_71011 = $signed(buffer_9_396) + $signed(buffer_5_397); // @[Modules.scala 68:83:@22991.4]
  assign _T_71012 = _T_71011[10:0]; // @[Modules.scala 68:83:@22992.4]
  assign buffer_9_590 = $signed(_T_71012); // @[Modules.scala 68:83:@22993.4]
  assign _T_71014 = $signed(buffer_9_398) + $signed(buffer_3_399); // @[Modules.scala 68:83:@22995.4]
  assign _T_71015 = _T_71014[10:0]; // @[Modules.scala 68:83:@22996.4]
  assign buffer_9_591 = $signed(_T_71015); // @[Modules.scala 68:83:@22997.4]
  assign _T_71020 = $signed(buffer_1_402) + $signed(buffer_9_403); // @[Modules.scala 68:83:@23003.4]
  assign _T_71021 = _T_71020[10:0]; // @[Modules.scala 68:83:@23004.4]
  assign buffer_9_593 = $signed(_T_71021); // @[Modules.scala 68:83:@23005.4]
  assign _T_71023 = $signed(buffer_1_404) + $signed(buffer_6_405); // @[Modules.scala 68:83:@23007.4]
  assign _T_71024 = _T_71023[10:0]; // @[Modules.scala 68:83:@23008.4]
  assign buffer_9_594 = $signed(_T_71024); // @[Modules.scala 68:83:@23009.4]
  assign _T_71026 = $signed(buffer_2_406) + $signed(buffer_1_407); // @[Modules.scala 68:83:@23011.4]
  assign _T_71027 = _T_71026[10:0]; // @[Modules.scala 68:83:@23012.4]
  assign buffer_9_595 = $signed(_T_71027); // @[Modules.scala 68:83:@23013.4]
  assign _T_71035 = $signed(buffer_9_412) + $signed(buffer_1_413); // @[Modules.scala 68:83:@23023.4]
  assign _T_71036 = _T_71035[10:0]; // @[Modules.scala 68:83:@23024.4]
  assign buffer_9_598 = $signed(_T_71036); // @[Modules.scala 68:83:@23025.4]
  assign _T_71047 = $signed(buffer_9_420) + $signed(buffer_7_421); // @[Modules.scala 68:83:@23039.4]
  assign _T_71048 = _T_71047[10:0]; // @[Modules.scala 68:83:@23040.4]
  assign buffer_9_602 = $signed(_T_71048); // @[Modules.scala 68:83:@23041.4]
  assign _T_71053 = $signed(buffer_1_424) + $signed(buffer_0_395); // @[Modules.scala 68:83:@23047.4]
  assign _T_71054 = _T_71053[10:0]; // @[Modules.scala 68:83:@23048.4]
  assign buffer_9_604 = $signed(_T_71054); // @[Modules.scala 68:83:@23049.4]
  assign _T_71056 = $signed(buffer_9_426) + $signed(buffer_5_427); // @[Modules.scala 68:83:@23051.4]
  assign _T_71057 = _T_71056[10:0]; // @[Modules.scala 68:83:@23052.4]
  assign buffer_9_605 = $signed(_T_71057); // @[Modules.scala 68:83:@23053.4]
  assign _T_71059 = $signed(buffer_4_428) + $signed(buffer_9_429); // @[Modules.scala 68:83:@23055.4]
  assign _T_71060 = _T_71059[10:0]; // @[Modules.scala 68:83:@23056.4]
  assign buffer_9_606 = $signed(_T_71060); // @[Modules.scala 68:83:@23057.4]
  assign _T_71062 = $signed(buffer_9_430) + $signed(buffer_9_431); // @[Modules.scala 68:83:@23059.4]
  assign _T_71063 = _T_71062[10:0]; // @[Modules.scala 68:83:@23060.4]
  assign buffer_9_607 = $signed(_T_71063); // @[Modules.scala 68:83:@23061.4]
  assign _T_71065 = $signed(buffer_0_395) + $signed(buffer_1_433); // @[Modules.scala 68:83:@23063.4]
  assign _T_71066 = _T_71065[10:0]; // @[Modules.scala 68:83:@23064.4]
  assign buffer_9_608 = $signed(_T_71066); // @[Modules.scala 68:83:@23065.4]
  assign _T_71068 = $signed(buffer_9_434) + $signed(buffer_1_435); // @[Modules.scala 68:83:@23067.4]
  assign _T_71069 = _T_71068[10:0]; // @[Modules.scala 68:83:@23068.4]
  assign buffer_9_609 = $signed(_T_71069); // @[Modules.scala 68:83:@23069.4]
  assign _T_71071 = $signed(buffer_7_436) + $signed(buffer_9_437); // @[Modules.scala 68:83:@23071.4]
  assign _T_71072 = _T_71071[10:0]; // @[Modules.scala 68:83:@23072.4]
  assign buffer_9_610 = $signed(_T_71072); // @[Modules.scala 68:83:@23073.4]
  assign _T_71074 = $signed(buffer_3_438) + $signed(buffer_0_395); // @[Modules.scala 68:83:@23075.4]
  assign _T_71075 = _T_71074[10:0]; // @[Modules.scala 68:83:@23076.4]
  assign buffer_9_611 = $signed(_T_71075); // @[Modules.scala 68:83:@23077.4]
  assign _T_71077 = $signed(buffer_9_440) + $signed(buffer_1_441); // @[Modules.scala 68:83:@23079.4]
  assign _T_71078 = _T_71077[10:0]; // @[Modules.scala 68:83:@23080.4]
  assign buffer_9_612 = $signed(_T_71078); // @[Modules.scala 68:83:@23081.4]
  assign _T_71080 = $signed(buffer_5_442) + $signed(buffer_9_443); // @[Modules.scala 68:83:@23083.4]
  assign _T_71081 = _T_71080[10:0]; // @[Modules.scala 68:83:@23084.4]
  assign buffer_9_613 = $signed(_T_71081); // @[Modules.scala 68:83:@23085.4]
  assign _T_71083 = $signed(buffer_2_444) + $signed(buffer_9_445); // @[Modules.scala 68:83:@23087.4]
  assign _T_71084 = _T_71083[10:0]; // @[Modules.scala 68:83:@23088.4]
  assign buffer_9_614 = $signed(_T_71084); // @[Modules.scala 68:83:@23089.4]
  assign _T_71086 = $signed(buffer_9_446) + $signed(buffer_9_447); // @[Modules.scala 68:83:@23091.4]
  assign _T_71087 = _T_71086[10:0]; // @[Modules.scala 68:83:@23092.4]
  assign buffer_9_615 = $signed(_T_71087); // @[Modules.scala 68:83:@23093.4]
  assign _T_71089 = $signed(buffer_9_448) + $signed(buffer_9_449); // @[Modules.scala 68:83:@23095.4]
  assign _T_71090 = _T_71089[10:0]; // @[Modules.scala 68:83:@23096.4]
  assign buffer_9_616 = $signed(_T_71090); // @[Modules.scala 68:83:@23097.4]
  assign _T_71092 = $signed(buffer_7_450) + $signed(buffer_9_451); // @[Modules.scala 68:83:@23099.4]
  assign _T_71093 = _T_71092[10:0]; // @[Modules.scala 68:83:@23100.4]
  assign buffer_9_617 = $signed(_T_71093); // @[Modules.scala 68:83:@23101.4]
  assign _T_71095 = $signed(buffer_4_452) + $signed(buffer_9_453); // @[Modules.scala 68:83:@23103.4]
  assign _T_71096 = _T_71095[10:0]; // @[Modules.scala 68:83:@23104.4]
  assign buffer_9_618 = $signed(_T_71096); // @[Modules.scala 68:83:@23105.4]
  assign _T_71101 = $signed(buffer_9_456) + $signed(buffer_1_457); // @[Modules.scala 68:83:@23111.4]
  assign _T_71102 = _T_71101[10:0]; // @[Modules.scala 68:83:@23112.4]
  assign buffer_9_620 = $signed(_T_71102); // @[Modules.scala 68:83:@23113.4]
  assign _T_71104 = $signed(buffer_9_458) + $signed(buffer_0_395); // @[Modules.scala 68:83:@23115.4]
  assign _T_71105 = _T_71104[10:0]; // @[Modules.scala 68:83:@23116.4]
  assign buffer_9_621 = $signed(_T_71105); // @[Modules.scala 68:83:@23117.4]
  assign _T_71107 = $signed(buffer_0_395) + $signed(buffer_9_461); // @[Modules.scala 68:83:@23119.4]
  assign _T_71108 = _T_71107[10:0]; // @[Modules.scala 68:83:@23120.4]
  assign buffer_9_622 = $signed(_T_71108); // @[Modules.scala 68:83:@23121.4]
  assign _T_71110 = $signed(buffer_9_462) + $signed(buffer_9_463); // @[Modules.scala 68:83:@23123.4]
  assign _T_71111 = _T_71110[10:0]; // @[Modules.scala 68:83:@23124.4]
  assign buffer_9_623 = $signed(_T_71111); // @[Modules.scala 68:83:@23125.4]
  assign _T_71116 = $signed(buffer_0_395) + $signed(buffer_9_467); // @[Modules.scala 68:83:@23131.4]
  assign _T_71117 = _T_71116[10:0]; // @[Modules.scala 68:83:@23132.4]
  assign buffer_9_625 = $signed(_T_71117); // @[Modules.scala 68:83:@23133.4]
  assign _T_71119 = $signed(buffer_9_468) + $signed(buffer_8_469); // @[Modules.scala 68:83:@23135.4]
  assign _T_71120 = _T_71119[10:0]; // @[Modules.scala 68:83:@23136.4]
  assign buffer_9_626 = $signed(_T_71120); // @[Modules.scala 68:83:@23137.4]
  assign _T_71122 = $signed(buffer_9_470) + $signed(buffer_0_395); // @[Modules.scala 68:83:@23139.4]
  assign _T_71123 = _T_71122[10:0]; // @[Modules.scala 68:83:@23140.4]
  assign buffer_9_627 = $signed(_T_71123); // @[Modules.scala 68:83:@23141.4]
  assign _T_71125 = $signed(buffer_9_472) + $signed(buffer_6_473); // @[Modules.scala 68:83:@23143.4]
  assign _T_71126 = _T_71125[10:0]; // @[Modules.scala 68:83:@23144.4]
  assign buffer_9_628 = $signed(_T_71126); // @[Modules.scala 68:83:@23145.4]
  assign _T_71128 = $signed(buffer_5_474) + $signed(buffer_1_475); // @[Modules.scala 68:83:@23147.4]
  assign _T_71129 = _T_71128[10:0]; // @[Modules.scala 68:83:@23148.4]
  assign buffer_9_629 = $signed(_T_71129); // @[Modules.scala 68:83:@23149.4]
  assign _T_71134 = $signed(buffer_0_395) + $signed(buffer_9_479); // @[Modules.scala 68:83:@23155.4]
  assign _T_71135 = _T_71134[10:0]; // @[Modules.scala 68:83:@23156.4]
  assign buffer_9_631 = $signed(_T_71135); // @[Modules.scala 68:83:@23157.4]
  assign _T_71137 = $signed(buffer_9_480) + $signed(buffer_9_481); // @[Modules.scala 68:83:@23159.4]
  assign _T_71138 = _T_71137[10:0]; // @[Modules.scala 68:83:@23160.4]
  assign buffer_9_632 = $signed(_T_71138); // @[Modules.scala 68:83:@23161.4]
  assign _T_71146 = $signed(buffer_0_486) + $signed(buffer_9_487); // @[Modules.scala 68:83:@23171.4]
  assign _T_71147 = _T_71146[10:0]; // @[Modules.scala 68:83:@23172.4]
  assign buffer_9_635 = $signed(_T_71147); // @[Modules.scala 68:83:@23173.4]
  assign _T_71149 = $signed(buffer_0_395) + $signed(buffer_9_489); // @[Modules.scala 68:83:@23175.4]
  assign _T_71150 = _T_71149[10:0]; // @[Modules.scala 68:83:@23176.4]
  assign buffer_9_636 = $signed(_T_71150); // @[Modules.scala 68:83:@23177.4]
  assign _T_71152 = $signed(buffer_9_490) + $signed(buffer_0_395); // @[Modules.scala 68:83:@23179.4]
  assign _T_71153 = _T_71152[10:0]; // @[Modules.scala 68:83:@23180.4]
  assign buffer_9_637 = $signed(_T_71153); // @[Modules.scala 68:83:@23181.4]
  assign _T_71155 = $signed(buffer_9_492) + $signed(buffer_0_493); // @[Modules.scala 68:83:@23183.4]
  assign _T_71156 = _T_71155[10:0]; // @[Modules.scala 68:83:@23184.4]
  assign buffer_9_638 = $signed(_T_71156); // @[Modules.scala 68:83:@23185.4]
  assign _T_71161 = $signed(buffer_3_496) + $signed(buffer_2_497); // @[Modules.scala 68:83:@23191.4]
  assign _T_71162 = _T_71161[10:0]; // @[Modules.scala 68:83:@23192.4]
  assign buffer_9_640 = $signed(_T_71162); // @[Modules.scala 68:83:@23193.4]
  assign _T_71164 = $signed(buffer_0_395) + $signed(buffer_9_499); // @[Modules.scala 68:83:@23195.4]
  assign _T_71165 = _T_71164[10:0]; // @[Modules.scala 68:83:@23196.4]
  assign buffer_9_641 = $signed(_T_71165); // @[Modules.scala 68:83:@23197.4]
  assign _T_71173 = $signed(buffer_9_504) + $signed(buffer_9_505); // @[Modules.scala 68:83:@23207.4]
  assign _T_71174 = _T_71173[10:0]; // @[Modules.scala 68:83:@23208.4]
  assign buffer_9_644 = $signed(_T_71174); // @[Modules.scala 68:83:@23209.4]
  assign _T_71176 = $signed(buffer_9_506) + $signed(buffer_2_507); // @[Modules.scala 68:83:@23211.4]
  assign _T_71177 = _T_71176[10:0]; // @[Modules.scala 68:83:@23212.4]
  assign buffer_9_645 = $signed(_T_71177); // @[Modules.scala 68:83:@23213.4]
  assign _T_71185 = $signed(buffer_9_512) + $signed(buffer_2_513); // @[Modules.scala 68:83:@23223.4]
  assign _T_71186 = _T_71185[10:0]; // @[Modules.scala 68:83:@23224.4]
  assign buffer_9_648 = $signed(_T_71186); // @[Modules.scala 68:83:@23225.4]
  assign _T_71188 = $signed(buffer_9_514) + $signed(buffer_1_515); // @[Modules.scala 68:83:@23227.4]
  assign _T_71189 = _T_71188[10:0]; // @[Modules.scala 68:83:@23228.4]
  assign buffer_9_649 = $signed(_T_71189); // @[Modules.scala 68:83:@23229.4]
  assign _T_71194 = $signed(buffer_1_518) + $signed(buffer_9_519); // @[Modules.scala 68:83:@23235.4]
  assign _T_71195 = _T_71194[10:0]; // @[Modules.scala 68:83:@23236.4]
  assign buffer_9_651 = $signed(_T_71195); // @[Modules.scala 68:83:@23237.4]
  assign _T_71206 = $signed(buffer_9_526) + $signed(buffer_1_527); // @[Modules.scala 68:83:@23251.4]
  assign _T_71207 = _T_71206[10:0]; // @[Modules.scala 68:83:@23252.4]
  assign buffer_9_655 = $signed(_T_71207); // @[Modules.scala 68:83:@23253.4]
  assign _T_71215 = $signed(buffer_8_532) + $signed(buffer_9_533); // @[Modules.scala 68:83:@23263.4]
  assign _T_71216 = _T_71215[10:0]; // @[Modules.scala 68:83:@23264.4]
  assign buffer_9_658 = $signed(_T_71216); // @[Modules.scala 68:83:@23265.4]
  assign _T_71218 = $signed(buffer_9_534) + $signed(buffer_9_535); // @[Modules.scala 68:83:@23267.4]
  assign _T_71219 = _T_71218[10:0]; // @[Modules.scala 68:83:@23268.4]
  assign buffer_9_659 = $signed(_T_71219); // @[Modules.scala 68:83:@23269.4]
  assign _T_71224 = $signed(buffer_8_538) + $signed(buffer_4_539); // @[Modules.scala 68:83:@23275.4]
  assign _T_71225 = _T_71224[10:0]; // @[Modules.scala 68:83:@23276.4]
  assign buffer_9_661 = $signed(_T_71225); // @[Modules.scala 68:83:@23277.4]
  assign _T_71227 = $signed(buffer_3_540) + $signed(buffer_9_541); // @[Modules.scala 68:83:@23279.4]
  assign _T_71228 = _T_71227[10:0]; // @[Modules.scala 68:83:@23280.4]
  assign buffer_9_662 = $signed(_T_71228); // @[Modules.scala 68:83:@23281.4]
  assign _T_71230 = $signed(buffer_9_542) + $signed(buffer_0_543); // @[Modules.scala 68:83:@23283.4]
  assign _T_71231 = _T_71230[10:0]; // @[Modules.scala 68:83:@23284.4]
  assign buffer_9_663 = $signed(_T_71231); // @[Modules.scala 68:83:@23285.4]
  assign _T_71233 = $signed(buffer_9_544) + $signed(buffer_3_545); // @[Modules.scala 68:83:@23287.4]
  assign _T_71234 = _T_71233[10:0]; // @[Modules.scala 68:83:@23288.4]
  assign buffer_9_664 = $signed(_T_71234); // @[Modules.scala 68:83:@23289.4]
  assign _T_71239 = $signed(buffer_9_548) + $signed(buffer_5_549); // @[Modules.scala 68:83:@23295.4]
  assign _T_71240 = _T_71239[10:0]; // @[Modules.scala 68:83:@23296.4]
  assign buffer_9_666 = $signed(_T_71240); // @[Modules.scala 68:83:@23297.4]
  assign _T_71242 = $signed(buffer_9_550) + $signed(buffer_9_551); // @[Modules.scala 68:83:@23299.4]
  assign _T_71243 = _T_71242[10:0]; // @[Modules.scala 68:83:@23300.4]
  assign buffer_9_667 = $signed(_T_71243); // @[Modules.scala 68:83:@23301.4]
  assign _T_71245 = $signed(buffer_9_552) + $signed(buffer_1_553); // @[Modules.scala 68:83:@23303.4]
  assign _T_71246 = _T_71245[10:0]; // @[Modules.scala 68:83:@23304.4]
  assign buffer_9_668 = $signed(_T_71246); // @[Modules.scala 68:83:@23305.4]
  assign _T_71248 = $signed(buffer_1_554) + $signed(buffer_9_555); // @[Modules.scala 68:83:@23307.4]
  assign _T_71249 = _T_71248[10:0]; // @[Modules.scala 68:83:@23308.4]
  assign buffer_9_669 = $signed(_T_71249); // @[Modules.scala 68:83:@23309.4]
  assign _T_71254 = $signed(buffer_9_558) + $signed(buffer_8_559); // @[Modules.scala 68:83:@23315.4]
  assign _T_71255 = _T_71254[10:0]; // @[Modules.scala 68:83:@23316.4]
  assign buffer_9_671 = $signed(_T_71255); // @[Modules.scala 68:83:@23317.4]
  assign _T_71257 = $signed(buffer_5_560) + $signed(buffer_0_561); // @[Modules.scala 68:83:@23319.4]
  assign _T_71258 = _T_71257[10:0]; // @[Modules.scala 68:83:@23320.4]
  assign buffer_9_672 = $signed(_T_71258); // @[Modules.scala 68:83:@23321.4]
  assign _T_71263 = $signed(buffer_4_564) + $signed(buffer_9_565); // @[Modules.scala 68:83:@23327.4]
  assign _T_71264 = _T_71263[10:0]; // @[Modules.scala 68:83:@23328.4]
  assign buffer_9_674 = $signed(_T_71264); // @[Modules.scala 68:83:@23329.4]
  assign _T_71266 = $signed(buffer_9_566) + $signed(buffer_9_567); // @[Modules.scala 68:83:@23331.4]
  assign _T_71267 = _T_71266[10:0]; // @[Modules.scala 68:83:@23332.4]
  assign buffer_9_675 = $signed(_T_71267); // @[Modules.scala 68:83:@23333.4]
  assign _T_71269 = $signed(buffer_0_395) + $signed(buffer_9_569); // @[Modules.scala 68:83:@23335.4]
  assign _T_71270 = _T_71269[10:0]; // @[Modules.scala 68:83:@23336.4]
  assign buffer_9_676 = $signed(_T_71270); // @[Modules.scala 68:83:@23337.4]
  assign _T_71272 = $signed(buffer_9_570) + $signed(buffer_9_571); // @[Modules.scala 68:83:@23339.4]
  assign _T_71273 = _T_71272[10:0]; // @[Modules.scala 68:83:@23340.4]
  assign buffer_9_677 = $signed(_T_71273); // @[Modules.scala 68:83:@23341.4]
  assign _T_71275 = $signed(buffer_0_395) + $signed(buffer_9_573); // @[Modules.scala 68:83:@23343.4]
  assign _T_71276 = _T_71275[10:0]; // @[Modules.scala 68:83:@23344.4]
  assign buffer_9_678 = $signed(_T_71276); // @[Modules.scala 68:83:@23345.4]
  assign _T_71278 = $signed(buffer_9_574) + $signed(buffer_0_395); // @[Modules.scala 68:83:@23347.4]
  assign _T_71279 = _T_71278[10:0]; // @[Modules.scala 68:83:@23348.4]
  assign buffer_9_679 = $signed(_T_71279); // @[Modules.scala 68:83:@23349.4]
  assign _T_71284 = $signed(buffer_9_578) + $signed(buffer_9_579); // @[Modules.scala 68:83:@23355.4]
  assign _T_71285 = _T_71284[10:0]; // @[Modules.scala 68:83:@23356.4]
  assign buffer_9_681 = $signed(_T_71285); // @[Modules.scala 68:83:@23357.4]
  assign _T_71287 = $signed(buffer_9_580) + $signed(buffer_9_581); // @[Modules.scala 68:83:@23359.4]
  assign _T_71288 = _T_71287[10:0]; // @[Modules.scala 68:83:@23360.4]
  assign buffer_9_682 = $signed(_T_71288); // @[Modules.scala 68:83:@23361.4]
  assign _T_71290 = $signed(buffer_9_582) + $signed(buffer_9_583); // @[Modules.scala 68:83:@23363.4]
  assign _T_71291 = _T_71290[10:0]; // @[Modules.scala 68:83:@23364.4]
  assign buffer_9_683 = $signed(_T_71291); // @[Modules.scala 68:83:@23365.4]
  assign _T_71293 = $signed(buffer_3_584) + $signed(buffer_9_585); // @[Modules.scala 68:83:@23367.4]
  assign _T_71294 = _T_71293[10:0]; // @[Modules.scala 68:83:@23368.4]
  assign buffer_9_684 = $signed(_T_71294); // @[Modules.scala 68:83:@23369.4]
  assign _T_71299 = $signed(buffer_9_588) + $signed(buffer_0_593); // @[Modules.scala 71:109:@23375.4]
  assign _T_71300 = _T_71299[10:0]; // @[Modules.scala 71:109:@23376.4]
  assign buffer_9_686 = $signed(_T_71300); // @[Modules.scala 71:109:@23377.4]
  assign _T_71302 = $signed(buffer_9_590) + $signed(buffer_9_591); // @[Modules.scala 71:109:@23379.4]
  assign _T_71303 = _T_71302[10:0]; // @[Modules.scala 71:109:@23380.4]
  assign buffer_9_687 = $signed(_T_71303); // @[Modules.scala 71:109:@23381.4]
  assign _T_71305 = $signed(buffer_2_592) + $signed(buffer_9_593); // @[Modules.scala 71:109:@23383.4]
  assign _T_71306 = _T_71305[10:0]; // @[Modules.scala 71:109:@23384.4]
  assign buffer_9_688 = $signed(_T_71306); // @[Modules.scala 71:109:@23385.4]
  assign _T_71308 = $signed(buffer_9_594) + $signed(buffer_9_595); // @[Modules.scala 71:109:@23387.4]
  assign _T_71309 = _T_71308[10:0]; // @[Modules.scala 71:109:@23388.4]
  assign buffer_9_689 = $signed(_T_71309); // @[Modules.scala 71:109:@23389.4]
  assign _T_71314 = $signed(buffer_9_598) + $signed(buffer_1_599); // @[Modules.scala 71:109:@23395.4]
  assign _T_71315 = _T_71314[10:0]; // @[Modules.scala 71:109:@23396.4]
  assign buffer_9_691 = $signed(_T_71315); // @[Modules.scala 71:109:@23397.4]
  assign _T_71320 = $signed(buffer_9_602) + $signed(buffer_3_603); // @[Modules.scala 71:109:@23403.4]
  assign _T_71321 = _T_71320[10:0]; // @[Modules.scala 71:109:@23404.4]
  assign buffer_9_693 = $signed(_T_71321); // @[Modules.scala 71:109:@23405.4]
  assign _T_71323 = $signed(buffer_9_604) + $signed(buffer_9_605); // @[Modules.scala 71:109:@23407.4]
  assign _T_71324 = _T_71323[10:0]; // @[Modules.scala 71:109:@23408.4]
  assign buffer_9_694 = $signed(_T_71324); // @[Modules.scala 71:109:@23409.4]
  assign _T_71326 = $signed(buffer_9_606) + $signed(buffer_9_607); // @[Modules.scala 71:109:@23411.4]
  assign _T_71327 = _T_71326[10:0]; // @[Modules.scala 71:109:@23412.4]
  assign buffer_9_695 = $signed(_T_71327); // @[Modules.scala 71:109:@23413.4]
  assign _T_71329 = $signed(buffer_9_608) + $signed(buffer_9_609); // @[Modules.scala 71:109:@23415.4]
  assign _T_71330 = _T_71329[10:0]; // @[Modules.scala 71:109:@23416.4]
  assign buffer_9_696 = $signed(_T_71330); // @[Modules.scala 71:109:@23417.4]
  assign _T_71332 = $signed(buffer_9_610) + $signed(buffer_9_611); // @[Modules.scala 71:109:@23419.4]
  assign _T_71333 = _T_71332[10:0]; // @[Modules.scala 71:109:@23420.4]
  assign buffer_9_697 = $signed(_T_71333); // @[Modules.scala 71:109:@23421.4]
  assign _T_71335 = $signed(buffer_9_612) + $signed(buffer_9_613); // @[Modules.scala 71:109:@23423.4]
  assign _T_71336 = _T_71335[10:0]; // @[Modules.scala 71:109:@23424.4]
  assign buffer_9_698 = $signed(_T_71336); // @[Modules.scala 71:109:@23425.4]
  assign _T_71338 = $signed(buffer_9_614) + $signed(buffer_9_615); // @[Modules.scala 71:109:@23427.4]
  assign _T_71339 = _T_71338[10:0]; // @[Modules.scala 71:109:@23428.4]
  assign buffer_9_699 = $signed(_T_71339); // @[Modules.scala 71:109:@23429.4]
  assign _T_71341 = $signed(buffer_9_616) + $signed(buffer_9_617); // @[Modules.scala 71:109:@23431.4]
  assign _T_71342 = _T_71341[10:0]; // @[Modules.scala 71:109:@23432.4]
  assign buffer_9_700 = $signed(_T_71342); // @[Modules.scala 71:109:@23433.4]
  assign _T_71344 = $signed(buffer_9_618) + $signed(buffer_5_619); // @[Modules.scala 71:109:@23435.4]
  assign _T_71345 = _T_71344[10:0]; // @[Modules.scala 71:109:@23436.4]
  assign buffer_9_701 = $signed(_T_71345); // @[Modules.scala 71:109:@23437.4]
  assign _T_71347 = $signed(buffer_9_620) + $signed(buffer_9_621); // @[Modules.scala 71:109:@23439.4]
  assign _T_71348 = _T_71347[10:0]; // @[Modules.scala 71:109:@23440.4]
  assign buffer_9_702 = $signed(_T_71348); // @[Modules.scala 71:109:@23441.4]
  assign _T_71350 = $signed(buffer_9_622) + $signed(buffer_9_623); // @[Modules.scala 71:109:@23443.4]
  assign _T_71351 = _T_71350[10:0]; // @[Modules.scala 71:109:@23444.4]
  assign buffer_9_703 = $signed(_T_71351); // @[Modules.scala 71:109:@23445.4]
  assign _T_71353 = $signed(buffer_5_624) + $signed(buffer_9_625); // @[Modules.scala 71:109:@23447.4]
  assign _T_71354 = _T_71353[10:0]; // @[Modules.scala 71:109:@23448.4]
  assign buffer_9_704 = $signed(_T_71354); // @[Modules.scala 71:109:@23449.4]
  assign _T_71356 = $signed(buffer_9_626) + $signed(buffer_9_627); // @[Modules.scala 71:109:@23451.4]
  assign _T_71357 = _T_71356[10:0]; // @[Modules.scala 71:109:@23452.4]
  assign buffer_9_705 = $signed(_T_71357); // @[Modules.scala 71:109:@23453.4]
  assign _T_71359 = $signed(buffer_9_628) + $signed(buffer_9_629); // @[Modules.scala 71:109:@23455.4]
  assign _T_71360 = _T_71359[10:0]; // @[Modules.scala 71:109:@23456.4]
  assign buffer_9_706 = $signed(_T_71360); // @[Modules.scala 71:109:@23457.4]
  assign _T_71362 = $signed(buffer_8_630) + $signed(buffer_9_631); // @[Modules.scala 71:109:@23459.4]
  assign _T_71363 = _T_71362[10:0]; // @[Modules.scala 71:109:@23460.4]
  assign buffer_9_707 = $signed(_T_71363); // @[Modules.scala 71:109:@23461.4]
  assign _T_71365 = $signed(buffer_9_632) + $signed(buffer_4_633); // @[Modules.scala 71:109:@23463.4]
  assign _T_71366 = _T_71365[10:0]; // @[Modules.scala 71:109:@23464.4]
  assign buffer_9_708 = $signed(_T_71366); // @[Modules.scala 71:109:@23465.4]
  assign _T_71368 = $signed(buffer_0_593) + $signed(buffer_9_635); // @[Modules.scala 71:109:@23467.4]
  assign _T_71369 = _T_71368[10:0]; // @[Modules.scala 71:109:@23468.4]
  assign buffer_9_709 = $signed(_T_71369); // @[Modules.scala 71:109:@23469.4]
  assign _T_71371 = $signed(buffer_9_636) + $signed(buffer_9_637); // @[Modules.scala 71:109:@23471.4]
  assign _T_71372 = _T_71371[10:0]; // @[Modules.scala 71:109:@23472.4]
  assign buffer_9_710 = $signed(_T_71372); // @[Modules.scala 71:109:@23473.4]
  assign _T_71374 = $signed(buffer_9_638) + $signed(buffer_5_639); // @[Modules.scala 71:109:@23475.4]
  assign _T_71375 = _T_71374[10:0]; // @[Modules.scala 71:109:@23476.4]
  assign buffer_9_711 = $signed(_T_71375); // @[Modules.scala 71:109:@23477.4]
  assign _T_71377 = $signed(buffer_9_640) + $signed(buffer_9_641); // @[Modules.scala 71:109:@23479.4]
  assign _T_71378 = _T_71377[10:0]; // @[Modules.scala 71:109:@23480.4]
  assign buffer_9_712 = $signed(_T_71378); // @[Modules.scala 71:109:@23481.4]
  assign _T_71380 = $signed(buffer_2_642) + $signed(buffer_3_643); // @[Modules.scala 71:109:@23483.4]
  assign _T_71381 = _T_71380[10:0]; // @[Modules.scala 71:109:@23484.4]
  assign buffer_9_713 = $signed(_T_71381); // @[Modules.scala 71:109:@23485.4]
  assign _T_71383 = $signed(buffer_9_644) + $signed(buffer_9_645); // @[Modules.scala 71:109:@23487.4]
  assign _T_71384 = _T_71383[10:0]; // @[Modules.scala 71:109:@23488.4]
  assign buffer_9_714 = $signed(_T_71384); // @[Modules.scala 71:109:@23489.4]
  assign _T_71386 = $signed(buffer_0_593) + $signed(buffer_4_647); // @[Modules.scala 71:109:@23491.4]
  assign _T_71387 = _T_71386[10:0]; // @[Modules.scala 71:109:@23492.4]
  assign buffer_9_715 = $signed(_T_71387); // @[Modules.scala 71:109:@23493.4]
  assign _T_71389 = $signed(buffer_9_648) + $signed(buffer_9_649); // @[Modules.scala 71:109:@23495.4]
  assign _T_71390 = _T_71389[10:0]; // @[Modules.scala 71:109:@23496.4]
  assign buffer_9_716 = $signed(_T_71390); // @[Modules.scala 71:109:@23497.4]
  assign _T_71392 = $signed(buffer_3_650) + $signed(buffer_9_651); // @[Modules.scala 71:109:@23499.4]
  assign _T_71393 = _T_71392[10:0]; // @[Modules.scala 71:109:@23500.4]
  assign buffer_9_717 = $signed(_T_71393); // @[Modules.scala 71:109:@23501.4]
  assign _T_71395 = $signed(buffer_7_652) + $signed(buffer_3_653); // @[Modules.scala 71:109:@23503.4]
  assign _T_71396 = _T_71395[10:0]; // @[Modules.scala 71:109:@23504.4]
  assign buffer_9_718 = $signed(_T_71396); // @[Modules.scala 71:109:@23505.4]
  assign _T_71398 = $signed(buffer_8_654) + $signed(buffer_9_655); // @[Modules.scala 71:109:@23507.4]
  assign _T_71399 = _T_71398[10:0]; // @[Modules.scala 71:109:@23508.4]
  assign buffer_9_719 = $signed(_T_71399); // @[Modules.scala 71:109:@23509.4]
  assign _T_71401 = $signed(buffer_1_656) + $signed(buffer_3_657); // @[Modules.scala 71:109:@23511.4]
  assign _T_71402 = _T_71401[10:0]; // @[Modules.scala 71:109:@23512.4]
  assign buffer_9_720 = $signed(_T_71402); // @[Modules.scala 71:109:@23513.4]
  assign _T_71404 = $signed(buffer_9_658) + $signed(buffer_9_659); // @[Modules.scala 71:109:@23515.4]
  assign _T_71405 = _T_71404[10:0]; // @[Modules.scala 71:109:@23516.4]
  assign buffer_9_721 = $signed(_T_71405); // @[Modules.scala 71:109:@23517.4]
  assign _T_71407 = $signed(buffer_7_660) + $signed(buffer_9_661); // @[Modules.scala 71:109:@23519.4]
  assign _T_71408 = _T_71407[10:0]; // @[Modules.scala 71:109:@23520.4]
  assign buffer_9_722 = $signed(_T_71408); // @[Modules.scala 71:109:@23521.4]
  assign _T_71410 = $signed(buffer_9_662) + $signed(buffer_9_663); // @[Modules.scala 71:109:@23523.4]
  assign _T_71411 = _T_71410[10:0]; // @[Modules.scala 71:109:@23524.4]
  assign buffer_9_723 = $signed(_T_71411); // @[Modules.scala 71:109:@23525.4]
  assign _T_71413 = $signed(buffer_9_664) + $signed(buffer_4_665); // @[Modules.scala 71:109:@23527.4]
  assign _T_71414 = _T_71413[10:0]; // @[Modules.scala 71:109:@23528.4]
  assign buffer_9_724 = $signed(_T_71414); // @[Modules.scala 71:109:@23529.4]
  assign _T_71416 = $signed(buffer_9_666) + $signed(buffer_9_667); // @[Modules.scala 71:109:@23531.4]
  assign _T_71417 = _T_71416[10:0]; // @[Modules.scala 71:109:@23532.4]
  assign buffer_9_725 = $signed(_T_71417); // @[Modules.scala 71:109:@23533.4]
  assign _T_71419 = $signed(buffer_9_668) + $signed(buffer_9_669); // @[Modules.scala 71:109:@23535.4]
  assign _T_71420 = _T_71419[10:0]; // @[Modules.scala 71:109:@23536.4]
  assign buffer_9_726 = $signed(_T_71420); // @[Modules.scala 71:109:@23537.4]
  assign _T_71422 = $signed(buffer_4_670) + $signed(buffer_9_671); // @[Modules.scala 71:109:@23539.4]
  assign _T_71423 = _T_71422[10:0]; // @[Modules.scala 71:109:@23540.4]
  assign buffer_9_727 = $signed(_T_71423); // @[Modules.scala 71:109:@23541.4]
  assign _T_71425 = $signed(buffer_9_672) + $signed(buffer_4_673); // @[Modules.scala 71:109:@23543.4]
  assign _T_71426 = _T_71425[10:0]; // @[Modules.scala 71:109:@23544.4]
  assign buffer_9_728 = $signed(_T_71426); // @[Modules.scala 71:109:@23545.4]
  assign _T_71428 = $signed(buffer_9_674) + $signed(buffer_9_675); // @[Modules.scala 71:109:@23547.4]
  assign _T_71429 = _T_71428[10:0]; // @[Modules.scala 71:109:@23548.4]
  assign buffer_9_729 = $signed(_T_71429); // @[Modules.scala 71:109:@23549.4]
  assign _T_71431 = $signed(buffer_9_676) + $signed(buffer_9_677); // @[Modules.scala 71:109:@23551.4]
  assign _T_71432 = _T_71431[10:0]; // @[Modules.scala 71:109:@23552.4]
  assign buffer_9_730 = $signed(_T_71432); // @[Modules.scala 71:109:@23553.4]
  assign _T_71434 = $signed(buffer_9_678) + $signed(buffer_9_679); // @[Modules.scala 71:109:@23555.4]
  assign _T_71435 = _T_71434[10:0]; // @[Modules.scala 71:109:@23556.4]
  assign buffer_9_731 = $signed(_T_71435); // @[Modules.scala 71:109:@23557.4]
  assign _T_71437 = $signed(buffer_0_593) + $signed(buffer_9_681); // @[Modules.scala 71:109:@23559.4]
  assign _T_71438 = _T_71437[10:0]; // @[Modules.scala 71:109:@23560.4]
  assign buffer_9_732 = $signed(_T_71438); // @[Modules.scala 71:109:@23561.4]
  assign _T_71440 = $signed(buffer_9_682) + $signed(buffer_9_683); // @[Modules.scala 71:109:@23563.4]
  assign _T_71441 = _T_71440[10:0]; // @[Modules.scala 71:109:@23564.4]
  assign buffer_9_733 = $signed(_T_71441); // @[Modules.scala 71:109:@23565.4]
  assign _T_71443 = $signed(buffer_9_684) + $signed(buffer_5_685); // @[Modules.scala 71:109:@23567.4]
  assign _T_71444 = _T_71443[10:0]; // @[Modules.scala 71:109:@23568.4]
  assign buffer_9_734 = $signed(_T_71444); // @[Modules.scala 71:109:@23569.4]
  assign _T_71446 = $signed(buffer_9_686) + $signed(buffer_9_687); // @[Modules.scala 78:156:@23572.4]
  assign _T_71447 = _T_71446[10:0]; // @[Modules.scala 78:156:@23573.4]
  assign buffer_9_736 = $signed(_T_71447); // @[Modules.scala 78:156:@23574.4]
  assign _T_71449 = $signed(buffer_9_736) + $signed(buffer_9_688); // @[Modules.scala 78:156:@23576.4]
  assign _T_71450 = _T_71449[10:0]; // @[Modules.scala 78:156:@23577.4]
  assign buffer_9_737 = $signed(_T_71450); // @[Modules.scala 78:156:@23578.4]
  assign _T_71452 = $signed(buffer_9_737) + $signed(buffer_9_689); // @[Modules.scala 78:156:@23580.4]
  assign _T_71453 = _T_71452[10:0]; // @[Modules.scala 78:156:@23581.4]
  assign buffer_9_738 = $signed(_T_71453); // @[Modules.scala 78:156:@23582.4]
  assign _T_71455 = $signed(buffer_9_738) + $signed(buffer_1_690); // @[Modules.scala 78:156:@23584.4]
  assign _T_71456 = _T_71455[10:0]; // @[Modules.scala 78:156:@23585.4]
  assign buffer_9_739 = $signed(_T_71456); // @[Modules.scala 78:156:@23586.4]
  assign _T_71458 = $signed(buffer_9_739) + $signed(buffer_9_691); // @[Modules.scala 78:156:@23588.4]
  assign _T_71459 = _T_71458[10:0]; // @[Modules.scala 78:156:@23589.4]
  assign buffer_9_740 = $signed(_T_71459); // @[Modules.scala 78:156:@23590.4]
  assign _T_71461 = $signed(buffer_9_740) + $signed(buffer_1_692); // @[Modules.scala 78:156:@23592.4]
  assign _T_71462 = _T_71461[10:0]; // @[Modules.scala 78:156:@23593.4]
  assign buffer_9_741 = $signed(_T_71462); // @[Modules.scala 78:156:@23594.4]
  assign _T_71464 = $signed(buffer_9_741) + $signed(buffer_9_693); // @[Modules.scala 78:156:@23596.4]
  assign _T_71465 = _T_71464[10:0]; // @[Modules.scala 78:156:@23597.4]
  assign buffer_9_742 = $signed(_T_71465); // @[Modules.scala 78:156:@23598.4]
  assign _T_71467 = $signed(buffer_9_742) + $signed(buffer_9_694); // @[Modules.scala 78:156:@23600.4]
  assign _T_71468 = _T_71467[10:0]; // @[Modules.scala 78:156:@23601.4]
  assign buffer_9_743 = $signed(_T_71468); // @[Modules.scala 78:156:@23602.4]
  assign _T_71470 = $signed(buffer_9_743) + $signed(buffer_9_695); // @[Modules.scala 78:156:@23604.4]
  assign _T_71471 = _T_71470[10:0]; // @[Modules.scala 78:156:@23605.4]
  assign buffer_9_744 = $signed(_T_71471); // @[Modules.scala 78:156:@23606.4]
  assign _T_71473 = $signed(buffer_9_744) + $signed(buffer_9_696); // @[Modules.scala 78:156:@23608.4]
  assign _T_71474 = _T_71473[10:0]; // @[Modules.scala 78:156:@23609.4]
  assign buffer_9_745 = $signed(_T_71474); // @[Modules.scala 78:156:@23610.4]
  assign _T_71476 = $signed(buffer_9_745) + $signed(buffer_9_697); // @[Modules.scala 78:156:@23612.4]
  assign _T_71477 = _T_71476[10:0]; // @[Modules.scala 78:156:@23613.4]
  assign buffer_9_746 = $signed(_T_71477); // @[Modules.scala 78:156:@23614.4]
  assign _T_71479 = $signed(buffer_9_746) + $signed(buffer_9_698); // @[Modules.scala 78:156:@23616.4]
  assign _T_71480 = _T_71479[10:0]; // @[Modules.scala 78:156:@23617.4]
  assign buffer_9_747 = $signed(_T_71480); // @[Modules.scala 78:156:@23618.4]
  assign _T_71482 = $signed(buffer_9_747) + $signed(buffer_9_699); // @[Modules.scala 78:156:@23620.4]
  assign _T_71483 = _T_71482[10:0]; // @[Modules.scala 78:156:@23621.4]
  assign buffer_9_748 = $signed(_T_71483); // @[Modules.scala 78:156:@23622.4]
  assign _T_71485 = $signed(buffer_9_748) + $signed(buffer_9_700); // @[Modules.scala 78:156:@23624.4]
  assign _T_71486 = _T_71485[10:0]; // @[Modules.scala 78:156:@23625.4]
  assign buffer_9_749 = $signed(_T_71486); // @[Modules.scala 78:156:@23626.4]
  assign _T_71488 = $signed(buffer_9_749) + $signed(buffer_9_701); // @[Modules.scala 78:156:@23628.4]
  assign _T_71489 = _T_71488[10:0]; // @[Modules.scala 78:156:@23629.4]
  assign buffer_9_750 = $signed(_T_71489); // @[Modules.scala 78:156:@23630.4]
  assign _T_71491 = $signed(buffer_9_750) + $signed(buffer_9_702); // @[Modules.scala 78:156:@23632.4]
  assign _T_71492 = _T_71491[10:0]; // @[Modules.scala 78:156:@23633.4]
  assign buffer_9_751 = $signed(_T_71492); // @[Modules.scala 78:156:@23634.4]
  assign _T_71494 = $signed(buffer_9_751) + $signed(buffer_9_703); // @[Modules.scala 78:156:@23636.4]
  assign _T_71495 = _T_71494[10:0]; // @[Modules.scala 78:156:@23637.4]
  assign buffer_9_752 = $signed(_T_71495); // @[Modules.scala 78:156:@23638.4]
  assign _T_71497 = $signed(buffer_9_752) + $signed(buffer_9_704); // @[Modules.scala 78:156:@23640.4]
  assign _T_71498 = _T_71497[10:0]; // @[Modules.scala 78:156:@23641.4]
  assign buffer_9_753 = $signed(_T_71498); // @[Modules.scala 78:156:@23642.4]
  assign _T_71500 = $signed(buffer_9_753) + $signed(buffer_9_705); // @[Modules.scala 78:156:@23644.4]
  assign _T_71501 = _T_71500[10:0]; // @[Modules.scala 78:156:@23645.4]
  assign buffer_9_754 = $signed(_T_71501); // @[Modules.scala 78:156:@23646.4]
  assign _T_71503 = $signed(buffer_9_754) + $signed(buffer_9_706); // @[Modules.scala 78:156:@23648.4]
  assign _T_71504 = _T_71503[10:0]; // @[Modules.scala 78:156:@23649.4]
  assign buffer_9_755 = $signed(_T_71504); // @[Modules.scala 78:156:@23650.4]
  assign _T_71506 = $signed(buffer_9_755) + $signed(buffer_9_707); // @[Modules.scala 78:156:@23652.4]
  assign _T_71507 = _T_71506[10:0]; // @[Modules.scala 78:156:@23653.4]
  assign buffer_9_756 = $signed(_T_71507); // @[Modules.scala 78:156:@23654.4]
  assign _T_71509 = $signed(buffer_9_756) + $signed(buffer_9_708); // @[Modules.scala 78:156:@23656.4]
  assign _T_71510 = _T_71509[10:0]; // @[Modules.scala 78:156:@23657.4]
  assign buffer_9_757 = $signed(_T_71510); // @[Modules.scala 78:156:@23658.4]
  assign _T_71512 = $signed(buffer_9_757) + $signed(buffer_9_709); // @[Modules.scala 78:156:@23660.4]
  assign _T_71513 = _T_71512[10:0]; // @[Modules.scala 78:156:@23661.4]
  assign buffer_9_758 = $signed(_T_71513); // @[Modules.scala 78:156:@23662.4]
  assign _T_71515 = $signed(buffer_9_758) + $signed(buffer_9_710); // @[Modules.scala 78:156:@23664.4]
  assign _T_71516 = _T_71515[10:0]; // @[Modules.scala 78:156:@23665.4]
  assign buffer_9_759 = $signed(_T_71516); // @[Modules.scala 78:156:@23666.4]
  assign _T_71518 = $signed(buffer_9_759) + $signed(buffer_9_711); // @[Modules.scala 78:156:@23668.4]
  assign _T_71519 = _T_71518[10:0]; // @[Modules.scala 78:156:@23669.4]
  assign buffer_9_760 = $signed(_T_71519); // @[Modules.scala 78:156:@23670.4]
  assign _T_71521 = $signed(buffer_9_760) + $signed(buffer_9_712); // @[Modules.scala 78:156:@23672.4]
  assign _T_71522 = _T_71521[10:0]; // @[Modules.scala 78:156:@23673.4]
  assign buffer_9_761 = $signed(_T_71522); // @[Modules.scala 78:156:@23674.4]
  assign _T_71524 = $signed(buffer_9_761) + $signed(buffer_9_713); // @[Modules.scala 78:156:@23676.4]
  assign _T_71525 = _T_71524[10:0]; // @[Modules.scala 78:156:@23677.4]
  assign buffer_9_762 = $signed(_T_71525); // @[Modules.scala 78:156:@23678.4]
  assign _T_71527 = $signed(buffer_9_762) + $signed(buffer_9_714); // @[Modules.scala 78:156:@23680.4]
  assign _T_71528 = _T_71527[10:0]; // @[Modules.scala 78:156:@23681.4]
  assign buffer_9_763 = $signed(_T_71528); // @[Modules.scala 78:156:@23682.4]
  assign _T_71530 = $signed(buffer_9_763) + $signed(buffer_9_715); // @[Modules.scala 78:156:@23684.4]
  assign _T_71531 = _T_71530[10:0]; // @[Modules.scala 78:156:@23685.4]
  assign buffer_9_764 = $signed(_T_71531); // @[Modules.scala 78:156:@23686.4]
  assign _T_71533 = $signed(buffer_9_764) + $signed(buffer_9_716); // @[Modules.scala 78:156:@23688.4]
  assign _T_71534 = _T_71533[10:0]; // @[Modules.scala 78:156:@23689.4]
  assign buffer_9_765 = $signed(_T_71534); // @[Modules.scala 78:156:@23690.4]
  assign _T_71536 = $signed(buffer_9_765) + $signed(buffer_9_717); // @[Modules.scala 78:156:@23692.4]
  assign _T_71537 = _T_71536[10:0]; // @[Modules.scala 78:156:@23693.4]
  assign buffer_9_766 = $signed(_T_71537); // @[Modules.scala 78:156:@23694.4]
  assign _T_71539 = $signed(buffer_9_766) + $signed(buffer_9_718); // @[Modules.scala 78:156:@23696.4]
  assign _T_71540 = _T_71539[10:0]; // @[Modules.scala 78:156:@23697.4]
  assign buffer_9_767 = $signed(_T_71540); // @[Modules.scala 78:156:@23698.4]
  assign _T_71542 = $signed(buffer_9_767) + $signed(buffer_9_719); // @[Modules.scala 78:156:@23700.4]
  assign _T_71543 = _T_71542[10:0]; // @[Modules.scala 78:156:@23701.4]
  assign buffer_9_768 = $signed(_T_71543); // @[Modules.scala 78:156:@23702.4]
  assign _T_71545 = $signed(buffer_9_768) + $signed(buffer_9_720); // @[Modules.scala 78:156:@23704.4]
  assign _T_71546 = _T_71545[10:0]; // @[Modules.scala 78:156:@23705.4]
  assign buffer_9_769 = $signed(_T_71546); // @[Modules.scala 78:156:@23706.4]
  assign _T_71548 = $signed(buffer_9_769) + $signed(buffer_9_721); // @[Modules.scala 78:156:@23708.4]
  assign _T_71549 = _T_71548[10:0]; // @[Modules.scala 78:156:@23709.4]
  assign buffer_9_770 = $signed(_T_71549); // @[Modules.scala 78:156:@23710.4]
  assign _T_71551 = $signed(buffer_9_770) + $signed(buffer_9_722); // @[Modules.scala 78:156:@23712.4]
  assign _T_71552 = _T_71551[10:0]; // @[Modules.scala 78:156:@23713.4]
  assign buffer_9_771 = $signed(_T_71552); // @[Modules.scala 78:156:@23714.4]
  assign _T_71554 = $signed(buffer_9_771) + $signed(buffer_9_723); // @[Modules.scala 78:156:@23716.4]
  assign _T_71555 = _T_71554[10:0]; // @[Modules.scala 78:156:@23717.4]
  assign buffer_9_772 = $signed(_T_71555); // @[Modules.scala 78:156:@23718.4]
  assign _T_71557 = $signed(buffer_9_772) + $signed(buffer_9_724); // @[Modules.scala 78:156:@23720.4]
  assign _T_71558 = _T_71557[10:0]; // @[Modules.scala 78:156:@23721.4]
  assign buffer_9_773 = $signed(_T_71558); // @[Modules.scala 78:156:@23722.4]
  assign _T_71560 = $signed(buffer_9_773) + $signed(buffer_9_725); // @[Modules.scala 78:156:@23724.4]
  assign _T_71561 = _T_71560[10:0]; // @[Modules.scala 78:156:@23725.4]
  assign buffer_9_774 = $signed(_T_71561); // @[Modules.scala 78:156:@23726.4]
  assign _T_71563 = $signed(buffer_9_774) + $signed(buffer_9_726); // @[Modules.scala 78:156:@23728.4]
  assign _T_71564 = _T_71563[10:0]; // @[Modules.scala 78:156:@23729.4]
  assign buffer_9_775 = $signed(_T_71564); // @[Modules.scala 78:156:@23730.4]
  assign _T_71566 = $signed(buffer_9_775) + $signed(buffer_9_727); // @[Modules.scala 78:156:@23732.4]
  assign _T_71567 = _T_71566[10:0]; // @[Modules.scala 78:156:@23733.4]
  assign buffer_9_776 = $signed(_T_71567); // @[Modules.scala 78:156:@23734.4]
  assign _T_71569 = $signed(buffer_9_776) + $signed(buffer_9_728); // @[Modules.scala 78:156:@23736.4]
  assign _T_71570 = _T_71569[10:0]; // @[Modules.scala 78:156:@23737.4]
  assign buffer_9_777 = $signed(_T_71570); // @[Modules.scala 78:156:@23738.4]
  assign _T_71572 = $signed(buffer_9_777) + $signed(buffer_9_729); // @[Modules.scala 78:156:@23740.4]
  assign _T_71573 = _T_71572[10:0]; // @[Modules.scala 78:156:@23741.4]
  assign buffer_9_778 = $signed(_T_71573); // @[Modules.scala 78:156:@23742.4]
  assign _T_71575 = $signed(buffer_9_778) + $signed(buffer_9_730); // @[Modules.scala 78:156:@23744.4]
  assign _T_71576 = _T_71575[10:0]; // @[Modules.scala 78:156:@23745.4]
  assign buffer_9_779 = $signed(_T_71576); // @[Modules.scala 78:156:@23746.4]
  assign _T_71578 = $signed(buffer_9_779) + $signed(buffer_9_731); // @[Modules.scala 78:156:@23748.4]
  assign _T_71579 = _T_71578[10:0]; // @[Modules.scala 78:156:@23749.4]
  assign buffer_9_780 = $signed(_T_71579); // @[Modules.scala 78:156:@23750.4]
  assign _T_71581 = $signed(buffer_9_780) + $signed(buffer_9_732); // @[Modules.scala 78:156:@23752.4]
  assign _T_71582 = _T_71581[10:0]; // @[Modules.scala 78:156:@23753.4]
  assign buffer_9_781 = $signed(_T_71582); // @[Modules.scala 78:156:@23754.4]
  assign _T_71584 = $signed(buffer_9_781) + $signed(buffer_9_733); // @[Modules.scala 78:156:@23756.4]
  assign _T_71585 = _T_71584[10:0]; // @[Modules.scala 78:156:@23757.4]
  assign buffer_9_782 = $signed(_T_71585); // @[Modules.scala 78:156:@23758.4]
  assign _T_71587 = $signed(buffer_9_782) + $signed(buffer_9_734); // @[Modules.scala 78:156:@23760.4]
  assign _T_71588 = _T_71587[10:0]; // @[Modules.scala 78:156:@23761.4]
  assign buffer_9_783 = $signed(_T_71588); // @[Modules.scala 78:156:@23762.4]
  assign _T_71705 = $signed(io_in_112) + $signed(io_in_113); // @[Modules.scala 37:46:@23929.4]
  assign _T_71706 = _T_71705[4:0]; // @[Modules.scala 37:46:@23930.4]
  assign _T_71707 = $signed(_T_71706); // @[Modules.scala 37:46:@23931.4]
  assign _T_71839 = $signed(io_in_308) + $signed(io_in_309); // @[Modules.scala 37:46:@24117.4]
  assign _T_71840 = _T_71839[4:0]; // @[Modules.scala 37:46:@24118.4]
  assign _T_71841 = $signed(_T_71840); // @[Modules.scala 37:46:@24119.4]
  assign _T_72129 = $signed(io_in_644) + $signed(io_in_645); // @[Modules.scala 37:46:@24534.4]
  assign _T_72130 = _T_72129[4:0]; // @[Modules.scala 37:46:@24535.4]
  assign _T_72131 = $signed(_T_72130); // @[Modules.scala 37:46:@24536.4]
  assign _T_72240 = $signed(11'sh0) + $signed(buffer_1_3); // @[Modules.scala 65:57:@24686.4]
  assign _T_72241 = _T_72240[10:0]; // @[Modules.scala 65:57:@24687.4]
  assign buffer_10_393 = $signed(_T_72241); // @[Modules.scala 65:57:@24688.4]
  assign _T_72243 = $signed(buffer_1_4) + $signed(buffer_3_5); // @[Modules.scala 65:57:@24690.4]
  assign _T_72244 = _T_72243[10:0]; // @[Modules.scala 65:57:@24691.4]
  assign buffer_10_394 = $signed(_T_72244); // @[Modules.scala 65:57:@24692.4]
  assign _T_72255 = $signed(buffer_0_12) + $signed(buffer_3_13); // @[Modules.scala 65:57:@24706.4]
  assign _T_72256 = _T_72255[10:0]; // @[Modules.scala 65:57:@24707.4]
  assign buffer_10_398 = $signed(_T_72256); // @[Modules.scala 65:57:@24708.4]
  assign _T_72276 = $signed(buffer_1_26) + $signed(buffer_0_27); // @[Modules.scala 65:57:@24734.4]
  assign _T_72277 = _T_72276[10:0]; // @[Modules.scala 65:57:@24735.4]
  assign buffer_10_405 = $signed(_T_72277); // @[Modules.scala 65:57:@24736.4]
  assign _T_72282 = $signed(11'sh0) + $signed(buffer_1_31); // @[Modules.scala 65:57:@24742.4]
  assign _T_72283 = _T_72282[10:0]; // @[Modules.scala 65:57:@24743.4]
  assign buffer_10_407 = $signed(_T_72283); // @[Modules.scala 65:57:@24744.4]
  assign _T_72300 = $signed(buffer_0_42) + $signed(buffer_1_43); // @[Modules.scala 65:57:@24766.4]
  assign _T_72301 = _T_72300[10:0]; // @[Modules.scala 65:57:@24767.4]
  assign buffer_10_413 = $signed(_T_72301); // @[Modules.scala 65:57:@24768.4]
  assign _T_72318 = $signed(buffer_0_54) + $signed(buffer_3_55); // @[Modules.scala 65:57:@24790.4]
  assign _T_72319 = _T_72318[10:0]; // @[Modules.scala 65:57:@24791.4]
  assign buffer_10_419 = $signed(_T_72319); // @[Modules.scala 65:57:@24792.4]
  assign buffer_10_56 = {{6{_T_71707[4]}},_T_71707}; // @[Modules.scala 32:22:@8.4]
  assign _T_72321 = $signed(buffer_10_56) + $signed(buffer_1_57); // @[Modules.scala 65:57:@24794.4]
  assign _T_72322 = _T_72321[10:0]; // @[Modules.scala 65:57:@24795.4]
  assign buffer_10_420 = $signed(_T_72322); // @[Modules.scala 65:57:@24796.4]
  assign _T_72333 = $signed(buffer_4_64) + $signed(buffer_1_65); // @[Modules.scala 65:57:@24810.4]
  assign _T_72334 = _T_72333[10:0]; // @[Modules.scala 65:57:@24811.4]
  assign buffer_10_424 = $signed(_T_72334); // @[Modules.scala 65:57:@24812.4]
  assign _T_72339 = $signed(buffer_5_68) + $signed(buffer_4_69); // @[Modules.scala 65:57:@24818.4]
  assign _T_72340 = _T_72339[10:0]; // @[Modules.scala 65:57:@24819.4]
  assign buffer_10_426 = $signed(_T_72340); // @[Modules.scala 65:57:@24820.4]
  assign _T_72342 = $signed(buffer_1_70) + $signed(buffer_5_71); // @[Modules.scala 65:57:@24822.4]
  assign _T_72343 = _T_72342[10:0]; // @[Modules.scala 65:57:@24823.4]
  assign buffer_10_427 = $signed(_T_72343); // @[Modules.scala 65:57:@24824.4]
  assign _T_72348 = $signed(buffer_1_74) + $signed(buffer_3_75); // @[Modules.scala 65:57:@24830.4]
  assign _T_72349 = _T_72348[10:0]; // @[Modules.scala 65:57:@24831.4]
  assign buffer_10_429 = $signed(_T_72349); // @[Modules.scala 65:57:@24832.4]
  assign buffer_10_77 = {{6{io_in_155[4]}},io_in_155}; // @[Modules.scala 32:22:@8.4]
  assign _T_72351 = $signed(buffer_4_76) + $signed(buffer_10_77); // @[Modules.scala 65:57:@24834.4]
  assign _T_72352 = _T_72351[10:0]; // @[Modules.scala 65:57:@24835.4]
  assign buffer_10_430 = $signed(_T_72352); // @[Modules.scala 65:57:@24836.4]
  assign _T_72354 = $signed(buffer_4_78) + $signed(11'sh0); // @[Modules.scala 65:57:@24838.4]
  assign _T_72355 = _T_72354[10:0]; // @[Modules.scala 65:57:@24839.4]
  assign buffer_10_431 = $signed(_T_72355); // @[Modules.scala 65:57:@24840.4]
  assign _T_72357 = $signed(buffer_4_80) + $signed(buffer_0_81); // @[Modules.scala 65:57:@24842.4]
  assign _T_72358 = _T_72357[10:0]; // @[Modules.scala 65:57:@24843.4]
  assign buffer_10_432 = $signed(_T_72358); // @[Modules.scala 65:57:@24844.4]
  assign _T_72360 = $signed(buffer_0_82) + $signed(buffer_1_83); // @[Modules.scala 65:57:@24846.4]
  assign _T_72361 = _T_72360[10:0]; // @[Modules.scala 65:57:@24847.4]
  assign buffer_10_433 = $signed(_T_72361); // @[Modules.scala 65:57:@24848.4]
  assign _T_72363 = $signed(buffer_4_84) + $signed(buffer_1_85); // @[Modules.scala 65:57:@24850.4]
  assign _T_72364 = _T_72363[10:0]; // @[Modules.scala 65:57:@24851.4]
  assign buffer_10_434 = $signed(_T_72364); // @[Modules.scala 65:57:@24852.4]
  assign _T_72366 = $signed(buffer_0_86) + $signed(buffer_7_87); // @[Modules.scala 65:57:@24854.4]
  assign _T_72367 = _T_72366[10:0]; // @[Modules.scala 65:57:@24855.4]
  assign buffer_10_435 = $signed(_T_72367); // @[Modules.scala 65:57:@24856.4]
  assign buffer_10_88 = {{6{io_in_176[4]}},io_in_176}; // @[Modules.scala 32:22:@8.4]
  assign _T_72369 = $signed(buffer_10_88) + $signed(buffer_7_89); // @[Modules.scala 65:57:@24858.4]
  assign _T_72370 = _T_72369[10:0]; // @[Modules.scala 65:57:@24859.4]
  assign buffer_10_436 = $signed(_T_72370); // @[Modules.scala 65:57:@24860.4]
  assign _T_72381 = $signed(11'sh0) + $signed(buffer_2_97); // @[Modules.scala 65:57:@24874.4]
  assign _T_72382 = _T_72381[10:0]; // @[Modules.scala 65:57:@24875.4]
  assign buffer_10_440 = $signed(_T_72382); // @[Modules.scala 65:57:@24876.4]
  assign buffer_10_100 = {{6{io_in_200[4]}},io_in_200}; // @[Modules.scala 32:22:@8.4]
  assign _T_72387 = $signed(buffer_10_100) + $signed(buffer_1_101); // @[Modules.scala 65:57:@24882.4]
  assign _T_72388 = _T_72387[10:0]; // @[Modules.scala 65:57:@24883.4]
  assign buffer_10_442 = $signed(_T_72388); // @[Modules.scala 65:57:@24884.4]
  assign _T_72390 = $signed(11'sh0) + $signed(buffer_1_103); // @[Modules.scala 65:57:@24886.4]
  assign _T_72391 = _T_72390[10:0]; // @[Modules.scala 65:57:@24887.4]
  assign buffer_10_443 = $signed(_T_72391); // @[Modules.scala 65:57:@24888.4]
  assign _T_72393 = $signed(11'sh0) + $signed(buffer_3_105); // @[Modules.scala 65:57:@24890.4]
  assign _T_72394 = _T_72393[10:0]; // @[Modules.scala 65:57:@24891.4]
  assign buffer_10_444 = $signed(_T_72394); // @[Modules.scala 65:57:@24892.4]
  assign _T_72408 = $signed(buffer_3_114) + $signed(11'sh0); // @[Modules.scala 65:57:@24910.4]
  assign _T_72409 = _T_72408[10:0]; // @[Modules.scala 65:57:@24911.4]
  assign buffer_10_449 = $signed(_T_72409); // @[Modules.scala 65:57:@24912.4]
  assign buffer_10_119 = {{6{io_in_238[4]}},io_in_238}; // @[Modules.scala 32:22:@8.4]
  assign _T_72414 = $signed(11'sh0) + $signed(buffer_10_119); // @[Modules.scala 65:57:@24918.4]
  assign _T_72415 = _T_72414[10:0]; // @[Modules.scala 65:57:@24919.4]
  assign buffer_10_451 = $signed(_T_72415); // @[Modules.scala 65:57:@24920.4]
  assign buffer_10_154 = {{6{_T_71841[4]}},_T_71841}; // @[Modules.scala 32:22:@8.4]
  assign _T_72468 = $signed(buffer_10_154) + $signed(buffer_3_155); // @[Modules.scala 65:57:@24990.4]
  assign _T_72469 = _T_72468[10:0]; // @[Modules.scala 65:57:@24991.4]
  assign buffer_10_469 = $signed(_T_72469); // @[Modules.scala 65:57:@24992.4]
  assign _T_72480 = $signed(buffer_5_162) + $signed(11'sh0); // @[Modules.scala 65:57:@25006.4]
  assign _T_72481 = _T_72480[10:0]; // @[Modules.scala 65:57:@25007.4]
  assign buffer_10_473 = $signed(_T_72481); // @[Modules.scala 65:57:@25008.4]
  assign _T_72486 = $signed(buffer_2_166) + $signed(buffer_0_167); // @[Modules.scala 65:57:@25014.4]
  assign _T_72487 = _T_72486[10:0]; // @[Modules.scala 65:57:@25015.4]
  assign buffer_10_475 = $signed(_T_72487); // @[Modules.scala 65:57:@25016.4]
  assign _T_72501 = $signed(buffer_0_176) + $signed(buffer_2_177); // @[Modules.scala 65:57:@25034.4]
  assign _T_72502 = _T_72501[10:0]; // @[Modules.scala 65:57:@25035.4]
  assign buffer_10_480 = $signed(_T_72502); // @[Modules.scala 65:57:@25036.4]
  assign _T_72522 = $signed(11'sh0) + $signed(buffer_0_191); // @[Modules.scala 65:57:@25062.4]
  assign _T_72523 = _T_72522[10:0]; // @[Modules.scala 65:57:@25063.4]
  assign buffer_10_487 = $signed(_T_72523); // @[Modules.scala 65:57:@25064.4]
  assign buffer_10_193 = {{6{io_in_387[4]}},io_in_387}; // @[Modules.scala 32:22:@8.4]
  assign _T_72525 = $signed(buffer_0_192) + $signed(buffer_10_193); // @[Modules.scala 65:57:@25066.4]
  assign _T_72526 = _T_72525[10:0]; // @[Modules.scala 65:57:@25067.4]
  assign buffer_10_488 = $signed(_T_72526); // @[Modules.scala 65:57:@25068.4]
  assign buffer_10_203 = {{6{io_in_406[4]}},io_in_406}; // @[Modules.scala 32:22:@8.4]
  assign _T_72540 = $signed(buffer_0_202) + $signed(buffer_10_203); // @[Modules.scala 65:57:@25086.4]
  assign _T_72541 = _T_72540[10:0]; // @[Modules.scala 65:57:@25087.4]
  assign buffer_10_493 = $signed(_T_72541); // @[Modules.scala 65:57:@25088.4]
  assign _T_72546 = $signed(11'sh0) + $signed(buffer_0_207); // @[Modules.scala 65:57:@25094.4]
  assign _T_72547 = _T_72546[10:0]; // @[Modules.scala 65:57:@25095.4]
  assign buffer_10_495 = $signed(_T_72547); // @[Modules.scala 65:57:@25096.4]
  assign _T_72549 = $signed(buffer_4_208) + $signed(buffer_3_209); // @[Modules.scala 65:57:@25098.4]
  assign _T_72550 = _T_72549[10:0]; // @[Modules.scala 65:57:@25099.4]
  assign buffer_10_496 = $signed(_T_72550); // @[Modules.scala 65:57:@25100.4]
  assign _T_72567 = $signed(buffer_1_220) + $signed(buffer_6_221); // @[Modules.scala 65:57:@25122.4]
  assign _T_72568 = _T_72567[10:0]; // @[Modules.scala 65:57:@25123.4]
  assign buffer_10_502 = $signed(_T_72568); // @[Modules.scala 65:57:@25124.4]
  assign _T_72576 = $signed(buffer_9_226) + $signed(buffer_4_227); // @[Modules.scala 65:57:@25134.4]
  assign _T_72577 = _T_72576[10:0]; // @[Modules.scala 65:57:@25135.4]
  assign buffer_10_505 = $signed(_T_72577); // @[Modules.scala 65:57:@25136.4]
  assign buffer_10_230 = {{6{io_in_461[4]}},io_in_461}; // @[Modules.scala 32:22:@8.4]
  assign _T_72582 = $signed(buffer_10_230) + $signed(buffer_5_231); // @[Modules.scala 65:57:@25142.4]
  assign _T_72583 = _T_72582[10:0]; // @[Modules.scala 65:57:@25143.4]
  assign buffer_10_507 = $signed(_T_72583); // @[Modules.scala 65:57:@25144.4]
  assign _T_72588 = $signed(buffer_1_234) + $signed(buffer_6_235); // @[Modules.scala 65:57:@25150.4]
  assign _T_72589 = _T_72588[10:0]; // @[Modules.scala 65:57:@25151.4]
  assign buffer_10_509 = $signed(_T_72589); // @[Modules.scala 65:57:@25152.4]
  assign _T_72603 = $signed(11'sh0) + $signed(buffer_9_245); // @[Modules.scala 65:57:@25170.4]
  assign _T_72604 = _T_72603[10:0]; // @[Modules.scala 65:57:@25171.4]
  assign buffer_10_514 = $signed(_T_72604); // @[Modules.scala 65:57:@25172.4]
  assign _T_72606 = $signed(buffer_4_246) + $signed(buffer_1_247); // @[Modules.scala 65:57:@25174.4]
  assign _T_72607 = _T_72606[10:0]; // @[Modules.scala 65:57:@25175.4]
  assign buffer_10_515 = $signed(_T_72607); // @[Modules.scala 65:57:@25176.4]
  assign buffer_10_255 = {{6{io_in_511[4]}},io_in_511}; // @[Modules.scala 32:22:@8.4]
  assign _T_72618 = $signed(buffer_1_254) + $signed(buffer_10_255); // @[Modules.scala 65:57:@25190.4]
  assign _T_72619 = _T_72618[10:0]; // @[Modules.scala 65:57:@25191.4]
  assign buffer_10_519 = $signed(_T_72619); // @[Modules.scala 65:57:@25192.4]
  assign _T_72621 = $signed(buffer_4_256) + $signed(buffer_0_257); // @[Modules.scala 65:57:@25194.4]
  assign _T_72622 = _T_72621[10:0]; // @[Modules.scala 65:57:@25195.4]
  assign buffer_10_520 = $signed(_T_72622); // @[Modules.scala 65:57:@25196.4]
  assign _T_72624 = $signed(buffer_2_258) + $signed(11'sh0); // @[Modules.scala 65:57:@25198.4]
  assign _T_72625 = _T_72624[10:0]; // @[Modules.scala 65:57:@25199.4]
  assign buffer_10_521 = $signed(_T_72625); // @[Modules.scala 65:57:@25200.4]
  assign _T_72642 = $signed(buffer_5_270) + $signed(buffer_1_271); // @[Modules.scala 65:57:@25222.4]
  assign _T_72643 = _T_72642[10:0]; // @[Modules.scala 65:57:@25223.4]
  assign buffer_10_527 = $signed(_T_72643); // @[Modules.scala 65:57:@25224.4]
  assign _T_72663 = $signed(buffer_1_284) + $signed(buffer_0_285); // @[Modules.scala 65:57:@25250.4]
  assign _T_72664 = _T_72663[10:0]; // @[Modules.scala 65:57:@25251.4]
  assign buffer_10_534 = $signed(_T_72664); // @[Modules.scala 65:57:@25252.4]
  assign _T_72672 = $signed(buffer_4_290) + $signed(buffer_5_291); // @[Modules.scala 65:57:@25262.4]
  assign _T_72673 = _T_72672[10:0]; // @[Modules.scala 65:57:@25263.4]
  assign buffer_10_537 = $signed(_T_72673); // @[Modules.scala 65:57:@25264.4]
  assign _T_72693 = $signed(buffer_2_304) + $signed(buffer_9_305); // @[Modules.scala 65:57:@25290.4]
  assign _T_72694 = _T_72693[10:0]; // @[Modules.scala 65:57:@25291.4]
  assign buffer_10_544 = $signed(_T_72694); // @[Modules.scala 65:57:@25292.4]
  assign _T_72696 = $signed(buffer_0_306) + $signed(buffer_4_307); // @[Modules.scala 65:57:@25294.4]
  assign _T_72697 = _T_72696[10:0]; // @[Modules.scala 65:57:@25295.4]
  assign buffer_10_545 = $signed(_T_72697); // @[Modules.scala 65:57:@25296.4]
  assign buffer_10_318 = {{6{io_in_636[4]}},io_in_636}; // @[Modules.scala 32:22:@8.4]
  assign _T_72714 = $signed(buffer_10_318) + $signed(buffer_0_319); // @[Modules.scala 65:57:@25318.4]
  assign _T_72715 = _T_72714[10:0]; // @[Modules.scala 65:57:@25319.4]
  assign buffer_10_551 = $signed(_T_72715); // @[Modules.scala 65:57:@25320.4]
  assign _T_72717 = $signed(buffer_9_320) + $signed(buffer_1_321); // @[Modules.scala 65:57:@25322.4]
  assign _T_72718 = _T_72717[10:0]; // @[Modules.scala 65:57:@25323.4]
  assign buffer_10_552 = $signed(_T_72718); // @[Modules.scala 65:57:@25324.4]
  assign buffer_10_322 = {{6{_T_72131[4]}},_T_72131}; // @[Modules.scala 32:22:@8.4]
  assign _T_72720 = $signed(buffer_10_322) + $signed(buffer_0_323); // @[Modules.scala 65:57:@25326.4]
  assign _T_72721 = _T_72720[10:0]; // @[Modules.scala 65:57:@25327.4]
  assign buffer_10_553 = $signed(_T_72721); // @[Modules.scala 65:57:@25328.4]
  assign _T_72726 = $signed(buffer_1_326) + $signed(buffer_6_327); // @[Modules.scala 65:57:@25334.4]
  assign _T_72727 = _T_72726[10:0]; // @[Modules.scala 65:57:@25335.4]
  assign buffer_10_555 = $signed(_T_72727); // @[Modules.scala 65:57:@25336.4]
  assign _T_72750 = $signed(buffer_2_342) + $signed(buffer_1_343); // @[Modules.scala 65:57:@25366.4]
  assign _T_72751 = _T_72750[10:0]; // @[Modules.scala 65:57:@25367.4]
  assign buffer_10_563 = $signed(_T_72751); // @[Modules.scala 65:57:@25368.4]
  assign buffer_10_353 = {{6{io_in_706[4]}},io_in_706}; // @[Modules.scala 32:22:@8.4]
  assign _T_72765 = $signed(11'sh0) + $signed(buffer_10_353); // @[Modules.scala 65:57:@25386.4]
  assign _T_72766 = _T_72765[10:0]; // @[Modules.scala 65:57:@25387.4]
  assign buffer_10_568 = $signed(_T_72766); // @[Modules.scala 65:57:@25388.4]
  assign buffer_10_368 = {{6{io_in_737[4]}},io_in_737}; // @[Modules.scala 32:22:@8.4]
  assign _T_72789 = $signed(buffer_10_368) + $signed(11'sh0); // @[Modules.scala 65:57:@25418.4]
  assign _T_72790 = _T_72789[10:0]; // @[Modules.scala 65:57:@25419.4]
  assign buffer_10_576 = $signed(_T_72790); // @[Modules.scala 65:57:@25420.4]
  assign _T_72801 = $signed(buffer_4_376) + $signed(11'sh0); // @[Modules.scala 65:57:@25434.4]
  assign _T_72802 = _T_72801[10:0]; // @[Modules.scala 65:57:@25435.4]
  assign buffer_10_580 = $signed(_T_72802); // @[Modules.scala 65:57:@25436.4]
  assign _T_72804 = $signed(buffer_3_378) + $signed(buffer_1_379); // @[Modules.scala 65:57:@25438.4]
  assign _T_72805 = _T_72804[10:0]; // @[Modules.scala 65:57:@25439.4]
  assign buffer_10_581 = $signed(_T_72805); // @[Modules.scala 65:57:@25440.4]
  assign _T_72807 = $signed(buffer_7_380) + $signed(buffer_1_381); // @[Modules.scala 65:57:@25442.4]
  assign _T_72808 = _T_72807[10:0]; // @[Modules.scala 65:57:@25443.4]
  assign buffer_10_582 = $signed(_T_72808); // @[Modules.scala 65:57:@25444.4]
  assign _T_72822 = $signed(buffer_7_390) + $signed(buffer_0_391); // @[Modules.scala 65:57:@25462.4]
  assign _T_72823 = _T_72822[10:0]; // @[Modules.scala 65:57:@25463.4]
  assign buffer_10_587 = $signed(_T_72823); // @[Modules.scala 65:57:@25464.4]
  assign _T_72825 = $signed(buffer_0_392) + $signed(buffer_10_393); // @[Modules.scala 68:83:@25466.4]
  assign _T_72826 = _T_72825[10:0]; // @[Modules.scala 68:83:@25467.4]
  assign buffer_10_588 = $signed(_T_72826); // @[Modules.scala 68:83:@25468.4]
  assign _T_72828 = $signed(buffer_10_394) + $signed(buffer_4_395); // @[Modules.scala 68:83:@25470.4]
  assign _T_72829 = _T_72828[10:0]; // @[Modules.scala 68:83:@25471.4]
  assign buffer_10_589 = $signed(_T_72829); // @[Modules.scala 68:83:@25472.4]
  assign _T_72834 = $signed(buffer_10_398) + $signed(buffer_1_399); // @[Modules.scala 68:83:@25478.4]
  assign _T_72835 = _T_72834[10:0]; // @[Modules.scala 68:83:@25479.4]
  assign buffer_10_591 = $signed(_T_72835); // @[Modules.scala 68:83:@25480.4]
  assign _T_72843 = $signed(buffer_1_404) + $signed(buffer_10_405); // @[Modules.scala 68:83:@25490.4]
  assign _T_72844 = _T_72843[10:0]; // @[Modules.scala 68:83:@25491.4]
  assign buffer_10_594 = $signed(_T_72844); // @[Modules.scala 68:83:@25492.4]
  assign _T_72846 = $signed(buffer_2_406) + $signed(buffer_10_407); // @[Modules.scala 68:83:@25494.4]
  assign _T_72847 = _T_72846[10:0]; // @[Modules.scala 68:83:@25495.4]
  assign buffer_10_595 = $signed(_T_72847); // @[Modules.scala 68:83:@25496.4]
  assign _T_72855 = $signed(buffer_9_412) + $signed(buffer_10_413); // @[Modules.scala 68:83:@25506.4]
  assign _T_72856 = _T_72855[10:0]; // @[Modules.scala 68:83:@25507.4]
  assign buffer_10_598 = $signed(_T_72856); // @[Modules.scala 68:83:@25508.4]
  assign _T_72864 = $signed(buffer_0_418) + $signed(buffer_10_419); // @[Modules.scala 68:83:@25518.4]
  assign _T_72865 = _T_72864[10:0]; // @[Modules.scala 68:83:@25519.4]
  assign buffer_10_601 = $signed(_T_72865); // @[Modules.scala 68:83:@25520.4]
  assign _T_72867 = $signed(buffer_10_420) + $signed(buffer_7_421); // @[Modules.scala 68:83:@25522.4]
  assign _T_72868 = _T_72867[10:0]; // @[Modules.scala 68:83:@25523.4]
  assign buffer_10_602 = $signed(_T_72868); // @[Modules.scala 68:83:@25524.4]
  assign _T_72870 = $signed(buffer_4_422) + $signed(buffer_3_423); // @[Modules.scala 68:83:@25526.4]
  assign _T_72871 = _T_72870[10:0]; // @[Modules.scala 68:83:@25527.4]
  assign buffer_10_603 = $signed(_T_72871); // @[Modules.scala 68:83:@25528.4]
  assign _T_72873 = $signed(buffer_10_424) + $signed(buffer_0_425); // @[Modules.scala 68:83:@25530.4]
  assign _T_72874 = _T_72873[10:0]; // @[Modules.scala 68:83:@25531.4]
  assign buffer_10_604 = $signed(_T_72874); // @[Modules.scala 68:83:@25532.4]
  assign _T_72876 = $signed(buffer_10_426) + $signed(buffer_10_427); // @[Modules.scala 68:83:@25534.4]
  assign _T_72877 = _T_72876[10:0]; // @[Modules.scala 68:83:@25535.4]
  assign buffer_10_605 = $signed(_T_72877); // @[Modules.scala 68:83:@25536.4]
  assign _T_72879 = $signed(buffer_4_428) + $signed(buffer_10_429); // @[Modules.scala 68:83:@25538.4]
  assign _T_72880 = _T_72879[10:0]; // @[Modules.scala 68:83:@25539.4]
  assign buffer_10_606 = $signed(_T_72880); // @[Modules.scala 68:83:@25540.4]
  assign _T_72882 = $signed(buffer_10_430) + $signed(buffer_10_431); // @[Modules.scala 68:83:@25542.4]
  assign _T_72883 = _T_72882[10:0]; // @[Modules.scala 68:83:@25543.4]
  assign buffer_10_607 = $signed(_T_72883); // @[Modules.scala 68:83:@25544.4]
  assign _T_72885 = $signed(buffer_10_432) + $signed(buffer_10_433); // @[Modules.scala 68:83:@25546.4]
  assign _T_72886 = _T_72885[10:0]; // @[Modules.scala 68:83:@25547.4]
  assign buffer_10_608 = $signed(_T_72886); // @[Modules.scala 68:83:@25548.4]
  assign _T_72888 = $signed(buffer_10_434) + $signed(buffer_10_435); // @[Modules.scala 68:83:@25550.4]
  assign _T_72889 = _T_72888[10:0]; // @[Modules.scala 68:83:@25551.4]
  assign buffer_10_609 = $signed(_T_72889); // @[Modules.scala 68:83:@25552.4]
  assign _T_72891 = $signed(buffer_10_436) + $signed(buffer_1_437); // @[Modules.scala 68:83:@25554.4]
  assign _T_72892 = _T_72891[10:0]; // @[Modules.scala 68:83:@25555.4]
  assign buffer_10_610 = $signed(_T_72892); // @[Modules.scala 68:83:@25556.4]
  assign _T_72897 = $signed(buffer_10_440) + $signed(buffer_3_441); // @[Modules.scala 68:83:@25562.4]
  assign _T_72898 = _T_72897[10:0]; // @[Modules.scala 68:83:@25563.4]
  assign buffer_10_612 = $signed(_T_72898); // @[Modules.scala 68:83:@25564.4]
  assign _T_72900 = $signed(buffer_10_442) + $signed(buffer_10_443); // @[Modules.scala 68:83:@25566.4]
  assign _T_72901 = _T_72900[10:0]; // @[Modules.scala 68:83:@25567.4]
  assign buffer_10_613 = $signed(_T_72901); // @[Modules.scala 68:83:@25568.4]
  assign _T_72903 = $signed(buffer_10_444) + $signed(buffer_0_445); // @[Modules.scala 68:83:@25570.4]
  assign _T_72904 = _T_72903[10:0]; // @[Modules.scala 68:83:@25571.4]
  assign buffer_10_614 = $signed(_T_72904); // @[Modules.scala 68:83:@25572.4]
  assign _T_72906 = $signed(buffer_0_395) + $signed(buffer_5_447); // @[Modules.scala 68:83:@25574.4]
  assign _T_72907 = _T_72906[10:0]; // @[Modules.scala 68:83:@25575.4]
  assign buffer_10_615 = $signed(_T_72907); // @[Modules.scala 68:83:@25576.4]
  assign _T_72909 = $signed(buffer_3_448) + $signed(buffer_10_449); // @[Modules.scala 68:83:@25578.4]
  assign _T_72910 = _T_72909[10:0]; // @[Modules.scala 68:83:@25579.4]
  assign buffer_10_616 = $signed(_T_72910); // @[Modules.scala 68:83:@25580.4]
  assign _T_72912 = $signed(buffer_0_395) + $signed(buffer_10_451); // @[Modules.scala 68:83:@25582.4]
  assign _T_72913 = _T_72912[10:0]; // @[Modules.scala 68:83:@25583.4]
  assign buffer_10_617 = $signed(_T_72913); // @[Modules.scala 68:83:@25584.4]
  assign _T_72918 = $signed(buffer_0_395) + $signed(buffer_3_455); // @[Modules.scala 68:83:@25590.4]
  assign _T_72919 = _T_72918[10:0]; // @[Modules.scala 68:83:@25591.4]
  assign buffer_10_619 = $signed(_T_72919); // @[Modules.scala 68:83:@25592.4]
  assign _T_72921 = $signed(buffer_3_456) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25594.4]
  assign _T_72922 = _T_72921[10:0]; // @[Modules.scala 68:83:@25595.4]
  assign buffer_10_620 = $signed(_T_72922); // @[Modules.scala 68:83:@25596.4]
  assign _T_72930 = $signed(buffer_9_462) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25606.4]
  assign _T_72931 = _T_72930[10:0]; // @[Modules.scala 68:83:@25607.4]
  assign buffer_10_623 = $signed(_T_72931); // @[Modules.scala 68:83:@25608.4]
  assign _T_72939 = $signed(buffer_5_468) + $signed(buffer_10_469); // @[Modules.scala 68:83:@25618.4]
  assign _T_72940 = _T_72939[10:0]; // @[Modules.scala 68:83:@25619.4]
  assign buffer_10_626 = $signed(_T_72940); // @[Modules.scala 68:83:@25620.4]
  assign _T_72945 = $signed(buffer_5_472) + $signed(buffer_10_473); // @[Modules.scala 68:83:@25626.4]
  assign _T_72946 = _T_72945[10:0]; // @[Modules.scala 68:83:@25627.4]
  assign buffer_10_628 = $signed(_T_72946); // @[Modules.scala 68:83:@25628.4]
  assign _T_72948 = $signed(buffer_0_395) + $signed(buffer_10_475); // @[Modules.scala 68:83:@25630.4]
  assign _T_72949 = _T_72948[10:0]; // @[Modules.scala 68:83:@25631.4]
  assign buffer_10_629 = $signed(_T_72949); // @[Modules.scala 68:83:@25632.4]
  assign _T_72957 = $signed(buffer_10_480) + $signed(buffer_5_481); // @[Modules.scala 68:83:@25642.4]
  assign _T_72958 = _T_72957[10:0]; // @[Modules.scala 68:83:@25643.4]
  assign buffer_10_632 = $signed(_T_72958); // @[Modules.scala 68:83:@25644.4]
  assign _T_72960 = $signed(buffer_4_482) + $signed(buffer_6_483); // @[Modules.scala 68:83:@25646.4]
  assign _T_72961 = _T_72960[10:0]; // @[Modules.scala 68:83:@25647.4]
  assign buffer_10_633 = $signed(_T_72961); // @[Modules.scala 68:83:@25648.4]
  assign _T_72966 = $signed(buffer_5_486) + $signed(buffer_10_487); // @[Modules.scala 68:83:@25654.4]
  assign _T_72967 = _T_72966[10:0]; // @[Modules.scala 68:83:@25655.4]
  assign buffer_10_635 = $signed(_T_72967); // @[Modules.scala 68:83:@25656.4]
  assign _T_72969 = $signed(buffer_10_488) + $signed(buffer_9_489); // @[Modules.scala 68:83:@25658.4]
  assign _T_72970 = _T_72969[10:0]; // @[Modules.scala 68:83:@25659.4]
  assign buffer_10_636 = $signed(_T_72970); // @[Modules.scala 68:83:@25660.4]
  assign _T_72972 = $signed(buffer_7_490) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25662.4]
  assign _T_72973 = _T_72972[10:0]; // @[Modules.scala 68:83:@25663.4]
  assign buffer_10_637 = $signed(_T_72973); // @[Modules.scala 68:83:@25664.4]
  assign _T_72975 = $signed(buffer_6_492) + $signed(buffer_10_493); // @[Modules.scala 68:83:@25666.4]
  assign _T_72976 = _T_72975[10:0]; // @[Modules.scala 68:83:@25667.4]
  assign buffer_10_638 = $signed(_T_72976); // @[Modules.scala 68:83:@25668.4]
  assign _T_72978 = $signed(buffer_7_494) + $signed(buffer_10_495); // @[Modules.scala 68:83:@25670.4]
  assign _T_72979 = _T_72978[10:0]; // @[Modules.scala 68:83:@25671.4]
  assign buffer_10_639 = $signed(_T_72979); // @[Modules.scala 68:83:@25672.4]
  assign _T_72981 = $signed(buffer_10_496) + $signed(buffer_3_497); // @[Modules.scala 68:83:@25674.4]
  assign _T_72982 = _T_72981[10:0]; // @[Modules.scala 68:83:@25675.4]
  assign buffer_10_640 = $signed(_T_72982); // @[Modules.scala 68:83:@25676.4]
  assign _T_72987 = $signed(buffer_0_500) + $signed(buffer_1_501); // @[Modules.scala 68:83:@25682.4]
  assign _T_72988 = _T_72987[10:0]; // @[Modules.scala 68:83:@25683.4]
  assign buffer_10_642 = $signed(_T_72988); // @[Modules.scala 68:83:@25684.4]
  assign _T_72990 = $signed(buffer_10_502) + $signed(buffer_3_503); // @[Modules.scala 68:83:@25686.4]
  assign _T_72991 = _T_72990[10:0]; // @[Modules.scala 68:83:@25687.4]
  assign buffer_10_643 = $signed(_T_72991); // @[Modules.scala 68:83:@25688.4]
  assign _T_72993 = $signed(buffer_9_504) + $signed(buffer_10_505); // @[Modules.scala 68:83:@25690.4]
  assign _T_72994 = _T_72993[10:0]; // @[Modules.scala 68:83:@25691.4]
  assign buffer_10_644 = $signed(_T_72994); // @[Modules.scala 68:83:@25692.4]
  assign _T_72996 = $signed(buffer_1_506) + $signed(buffer_10_507); // @[Modules.scala 68:83:@25694.4]
  assign _T_72997 = _T_72996[10:0]; // @[Modules.scala 68:83:@25695.4]
  assign buffer_10_645 = $signed(_T_72997); // @[Modules.scala 68:83:@25696.4]
  assign _T_72999 = $signed(buffer_3_508) + $signed(buffer_10_509); // @[Modules.scala 68:83:@25698.4]
  assign _T_73000 = _T_72999[10:0]; // @[Modules.scala 68:83:@25699.4]
  assign buffer_10_646 = $signed(_T_73000); // @[Modules.scala 68:83:@25700.4]
  assign _T_73005 = $signed(buffer_4_512) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25706.4]
  assign _T_73006 = _T_73005[10:0]; // @[Modules.scala 68:83:@25707.4]
  assign buffer_10_648 = $signed(_T_73006); // @[Modules.scala 68:83:@25708.4]
  assign _T_73008 = $signed(buffer_10_514) + $signed(buffer_10_515); // @[Modules.scala 68:83:@25710.4]
  assign _T_73009 = _T_73008[10:0]; // @[Modules.scala 68:83:@25711.4]
  assign buffer_10_649 = $signed(_T_73009); // @[Modules.scala 68:83:@25712.4]
  assign _T_73014 = $signed(buffer_4_518) + $signed(buffer_10_519); // @[Modules.scala 68:83:@25718.4]
  assign _T_73015 = _T_73014[10:0]; // @[Modules.scala 68:83:@25719.4]
  assign buffer_10_651 = $signed(_T_73015); // @[Modules.scala 68:83:@25720.4]
  assign _T_73017 = $signed(buffer_10_520) + $signed(buffer_10_521); // @[Modules.scala 68:83:@25722.4]
  assign _T_73018 = _T_73017[10:0]; // @[Modules.scala 68:83:@25723.4]
  assign buffer_10_652 = $signed(_T_73018); // @[Modules.scala 68:83:@25724.4]
  assign _T_73020 = $signed(buffer_1_522) + $signed(buffer_4_523); // @[Modules.scala 68:83:@25726.4]
  assign _T_73021 = _T_73020[10:0]; // @[Modules.scala 68:83:@25727.4]
  assign buffer_10_653 = $signed(_T_73021); // @[Modules.scala 68:83:@25728.4]
  assign _T_73026 = $signed(buffer_9_526) + $signed(buffer_10_527); // @[Modules.scala 68:83:@25734.4]
  assign _T_73027 = _T_73026[10:0]; // @[Modules.scala 68:83:@25735.4]
  assign buffer_10_655 = $signed(_T_73027); // @[Modules.scala 68:83:@25736.4]
  assign _T_73029 = $signed(buffer_7_528) + $signed(buffer_1_529); // @[Modules.scala 68:83:@25738.4]
  assign _T_73030 = _T_73029[10:0]; // @[Modules.scala 68:83:@25739.4]
  assign buffer_10_656 = $signed(_T_73030); // @[Modules.scala 68:83:@25740.4]
  assign _T_73032 = $signed(buffer_3_530) + $signed(buffer_5_531); // @[Modules.scala 68:83:@25742.4]
  assign _T_73033 = _T_73032[10:0]; // @[Modules.scala 68:83:@25743.4]
  assign buffer_10_657 = $signed(_T_73033); // @[Modules.scala 68:83:@25744.4]
  assign _T_73035 = $signed(buffer_8_532) + $signed(buffer_3_533); // @[Modules.scala 68:83:@25746.4]
  assign _T_73036 = _T_73035[10:0]; // @[Modules.scala 68:83:@25747.4]
  assign buffer_10_658 = $signed(_T_73036); // @[Modules.scala 68:83:@25748.4]
  assign _T_73038 = $signed(buffer_10_534) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25750.4]
  assign _T_73039 = _T_73038[10:0]; // @[Modules.scala 68:83:@25751.4]
  assign buffer_10_659 = $signed(_T_73039); // @[Modules.scala 68:83:@25752.4]
  assign _T_73041 = $signed(buffer_2_536) + $signed(buffer_10_537); // @[Modules.scala 68:83:@25754.4]
  assign _T_73042 = _T_73041[10:0]; // @[Modules.scala 68:83:@25755.4]
  assign buffer_10_660 = $signed(_T_73042); // @[Modules.scala 68:83:@25756.4]
  assign _T_73053 = $signed(buffer_10_544) + $signed(buffer_10_545); // @[Modules.scala 68:83:@25770.4]
  assign _T_73054 = _T_73053[10:0]; // @[Modules.scala 68:83:@25771.4]
  assign buffer_10_664 = $signed(_T_73054); // @[Modules.scala 68:83:@25772.4]
  assign _T_73059 = $signed(buffer_6_548) + $signed(buffer_8_549); // @[Modules.scala 68:83:@25778.4]
  assign _T_73060 = _T_73059[10:0]; // @[Modules.scala 68:83:@25779.4]
  assign buffer_10_666 = $signed(_T_73060); // @[Modules.scala 68:83:@25780.4]
  assign _T_73062 = $signed(buffer_2_550) + $signed(buffer_10_551); // @[Modules.scala 68:83:@25782.4]
  assign _T_73063 = _T_73062[10:0]; // @[Modules.scala 68:83:@25783.4]
  assign buffer_10_667 = $signed(_T_73063); // @[Modules.scala 68:83:@25784.4]
  assign _T_73065 = $signed(buffer_10_552) + $signed(buffer_10_553); // @[Modules.scala 68:83:@25786.4]
  assign _T_73066 = _T_73065[10:0]; // @[Modules.scala 68:83:@25787.4]
  assign buffer_10_668 = $signed(_T_73066); // @[Modules.scala 68:83:@25788.4]
  assign _T_73068 = $signed(buffer_1_554) + $signed(buffer_10_555); // @[Modules.scala 68:83:@25790.4]
  assign _T_73069 = _T_73068[10:0]; // @[Modules.scala 68:83:@25791.4]
  assign buffer_10_669 = $signed(_T_73069); // @[Modules.scala 68:83:@25792.4]
  assign _T_73080 = $signed(buffer_3_562) + $signed(buffer_10_563); // @[Modules.scala 68:83:@25806.4]
  assign _T_73081 = _T_73080[10:0]; // @[Modules.scala 68:83:@25807.4]
  assign buffer_10_673 = $signed(_T_73081); // @[Modules.scala 68:83:@25808.4]
  assign _T_73089 = $signed(buffer_10_568) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25818.4]
  assign _T_73090 = _T_73089[10:0]; // @[Modules.scala 68:83:@25819.4]
  assign buffer_10_676 = $signed(_T_73090); // @[Modules.scala 68:83:@25820.4]
  assign _T_73095 = $signed(buffer_0_395) + $signed(buffer_1_573); // @[Modules.scala 68:83:@25826.4]
  assign _T_73096 = _T_73095[10:0]; // @[Modules.scala 68:83:@25827.4]
  assign buffer_10_678 = $signed(_T_73096); // @[Modules.scala 68:83:@25828.4]
  assign _T_73098 = $signed(buffer_3_574) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25830.4]
  assign _T_73099 = _T_73098[10:0]; // @[Modules.scala 68:83:@25831.4]
  assign buffer_10_679 = $signed(_T_73099); // @[Modules.scala 68:83:@25832.4]
  assign _T_73101 = $signed(buffer_10_576) + $signed(buffer_0_395); // @[Modules.scala 68:83:@25834.4]
  assign _T_73102 = _T_73101[10:0]; // @[Modules.scala 68:83:@25835.4]
  assign buffer_10_680 = $signed(_T_73102); // @[Modules.scala 68:83:@25836.4]
  assign _T_73107 = $signed(buffer_10_580) + $signed(buffer_10_581); // @[Modules.scala 68:83:@25842.4]
  assign _T_73108 = _T_73107[10:0]; // @[Modules.scala 68:83:@25843.4]
  assign buffer_10_682 = $signed(_T_73108); // @[Modules.scala 68:83:@25844.4]
  assign _T_73110 = $signed(buffer_10_582) + $signed(buffer_3_583); // @[Modules.scala 68:83:@25846.4]
  assign _T_73111 = _T_73110[10:0]; // @[Modules.scala 68:83:@25847.4]
  assign buffer_10_683 = $signed(_T_73111); // @[Modules.scala 68:83:@25848.4]
  assign _T_73116 = $signed(buffer_5_586) + $signed(buffer_10_587); // @[Modules.scala 68:83:@25854.4]
  assign _T_73117 = _T_73116[10:0]; // @[Modules.scala 68:83:@25855.4]
  assign buffer_10_685 = $signed(_T_73117); // @[Modules.scala 68:83:@25856.4]
  assign _T_73119 = $signed(buffer_10_588) + $signed(buffer_10_589); // @[Modules.scala 71:109:@25858.4]
  assign _T_73120 = _T_73119[10:0]; // @[Modules.scala 71:109:@25859.4]
  assign buffer_10_686 = $signed(_T_73120); // @[Modules.scala 71:109:@25860.4]
  assign _T_73122 = $signed(buffer_9_590) + $signed(buffer_10_591); // @[Modules.scala 71:109:@25862.4]
  assign _T_73123 = _T_73122[10:0]; // @[Modules.scala 71:109:@25863.4]
  assign buffer_10_687 = $signed(_T_73123); // @[Modules.scala 71:109:@25864.4]
  assign _T_73128 = $signed(buffer_10_594) + $signed(buffer_10_595); // @[Modules.scala 71:109:@25870.4]
  assign _T_73129 = _T_73128[10:0]; // @[Modules.scala 71:109:@25871.4]
  assign buffer_10_689 = $signed(_T_73129); // @[Modules.scala 71:109:@25872.4]
  assign _T_73134 = $signed(buffer_10_598) + $signed(buffer_1_599); // @[Modules.scala 71:109:@25878.4]
  assign _T_73135 = _T_73134[10:0]; // @[Modules.scala 71:109:@25879.4]
  assign buffer_10_691 = $signed(_T_73135); // @[Modules.scala 71:109:@25880.4]
  assign _T_73137 = $signed(buffer_1_600) + $signed(buffer_10_601); // @[Modules.scala 71:109:@25882.4]
  assign _T_73138 = _T_73137[10:0]; // @[Modules.scala 71:109:@25883.4]
  assign buffer_10_692 = $signed(_T_73138); // @[Modules.scala 71:109:@25884.4]
  assign _T_73140 = $signed(buffer_10_602) + $signed(buffer_10_603); // @[Modules.scala 71:109:@25886.4]
  assign _T_73141 = _T_73140[10:0]; // @[Modules.scala 71:109:@25887.4]
  assign buffer_10_693 = $signed(_T_73141); // @[Modules.scala 71:109:@25888.4]
  assign _T_73143 = $signed(buffer_10_604) + $signed(buffer_10_605); // @[Modules.scala 71:109:@25890.4]
  assign _T_73144 = _T_73143[10:0]; // @[Modules.scala 71:109:@25891.4]
  assign buffer_10_694 = $signed(_T_73144); // @[Modules.scala 71:109:@25892.4]
  assign _T_73146 = $signed(buffer_10_606) + $signed(buffer_10_607); // @[Modules.scala 71:109:@25894.4]
  assign _T_73147 = _T_73146[10:0]; // @[Modules.scala 71:109:@25895.4]
  assign buffer_10_695 = $signed(_T_73147); // @[Modules.scala 71:109:@25896.4]
  assign _T_73149 = $signed(buffer_10_608) + $signed(buffer_10_609); // @[Modules.scala 71:109:@25898.4]
  assign _T_73150 = _T_73149[10:0]; // @[Modules.scala 71:109:@25899.4]
  assign buffer_10_696 = $signed(_T_73150); // @[Modules.scala 71:109:@25900.4]
  assign _T_73152 = $signed(buffer_10_610) + $signed(buffer_0_593); // @[Modules.scala 71:109:@25902.4]
  assign _T_73153 = _T_73152[10:0]; // @[Modules.scala 71:109:@25903.4]
  assign buffer_10_697 = $signed(_T_73153); // @[Modules.scala 71:109:@25904.4]
  assign _T_73155 = $signed(buffer_10_612) + $signed(buffer_10_613); // @[Modules.scala 71:109:@25906.4]
  assign _T_73156 = _T_73155[10:0]; // @[Modules.scala 71:109:@25907.4]
  assign buffer_10_698 = $signed(_T_73156); // @[Modules.scala 71:109:@25908.4]
  assign _T_73158 = $signed(buffer_10_614) + $signed(buffer_10_615); // @[Modules.scala 71:109:@25910.4]
  assign _T_73159 = _T_73158[10:0]; // @[Modules.scala 71:109:@25911.4]
  assign buffer_10_699 = $signed(_T_73159); // @[Modules.scala 71:109:@25912.4]
  assign _T_73161 = $signed(buffer_10_616) + $signed(buffer_10_617); // @[Modules.scala 71:109:@25914.4]
  assign _T_73162 = _T_73161[10:0]; // @[Modules.scala 71:109:@25915.4]
  assign buffer_10_700 = $signed(_T_73162); // @[Modules.scala 71:109:@25916.4]
  assign _T_73164 = $signed(buffer_0_593) + $signed(buffer_10_619); // @[Modules.scala 71:109:@25918.4]
  assign _T_73165 = _T_73164[10:0]; // @[Modules.scala 71:109:@25919.4]
  assign buffer_10_701 = $signed(_T_73165); // @[Modules.scala 71:109:@25920.4]
  assign _T_73167 = $signed(buffer_10_620) + $signed(buffer_0_593); // @[Modules.scala 71:109:@25922.4]
  assign _T_73168 = _T_73167[10:0]; // @[Modules.scala 71:109:@25923.4]
  assign buffer_10_702 = $signed(_T_73168); // @[Modules.scala 71:109:@25924.4]
  assign _T_73170 = $signed(buffer_0_593) + $signed(buffer_10_623); // @[Modules.scala 71:109:@25926.4]
  assign _T_73171 = _T_73170[10:0]; // @[Modules.scala 71:109:@25927.4]
  assign buffer_10_703 = $signed(_T_73171); // @[Modules.scala 71:109:@25928.4]
  assign _T_73173 = $signed(buffer_5_624) + $signed(buffer_0_593); // @[Modules.scala 71:109:@25930.4]
  assign _T_73174 = _T_73173[10:0]; // @[Modules.scala 71:109:@25931.4]
  assign buffer_10_704 = $signed(_T_73174); // @[Modules.scala 71:109:@25932.4]
  assign _T_73176 = $signed(buffer_10_626) + $signed(buffer_0_593); // @[Modules.scala 71:109:@25934.4]
  assign _T_73177 = _T_73176[10:0]; // @[Modules.scala 71:109:@25935.4]
  assign buffer_10_705 = $signed(_T_73177); // @[Modules.scala 71:109:@25936.4]
  assign _T_73179 = $signed(buffer_10_628) + $signed(buffer_10_629); // @[Modules.scala 71:109:@25938.4]
  assign _T_73180 = _T_73179[10:0]; // @[Modules.scala 71:109:@25939.4]
  assign buffer_10_706 = $signed(_T_73180); // @[Modules.scala 71:109:@25940.4]
  assign _T_73185 = $signed(buffer_10_632) + $signed(buffer_10_633); // @[Modules.scala 71:109:@25946.4]
  assign _T_73186 = _T_73185[10:0]; // @[Modules.scala 71:109:@25947.4]
  assign buffer_10_708 = $signed(_T_73186); // @[Modules.scala 71:109:@25948.4]
  assign _T_73188 = $signed(buffer_0_593) + $signed(buffer_10_635); // @[Modules.scala 71:109:@25950.4]
  assign _T_73189 = _T_73188[10:0]; // @[Modules.scala 71:109:@25951.4]
  assign buffer_10_709 = $signed(_T_73189); // @[Modules.scala 71:109:@25952.4]
  assign _T_73191 = $signed(buffer_10_636) + $signed(buffer_10_637); // @[Modules.scala 71:109:@25954.4]
  assign _T_73192 = _T_73191[10:0]; // @[Modules.scala 71:109:@25955.4]
  assign buffer_10_710 = $signed(_T_73192); // @[Modules.scala 71:109:@25956.4]
  assign _T_73194 = $signed(buffer_10_638) + $signed(buffer_10_639); // @[Modules.scala 71:109:@25958.4]
  assign _T_73195 = _T_73194[10:0]; // @[Modules.scala 71:109:@25959.4]
  assign buffer_10_711 = $signed(_T_73195); // @[Modules.scala 71:109:@25960.4]
  assign _T_73197 = $signed(buffer_10_640) + $signed(buffer_0_593); // @[Modules.scala 71:109:@25962.4]
  assign _T_73198 = _T_73197[10:0]; // @[Modules.scala 71:109:@25963.4]
  assign buffer_10_712 = $signed(_T_73198); // @[Modules.scala 71:109:@25964.4]
  assign _T_73200 = $signed(buffer_10_642) + $signed(buffer_10_643); // @[Modules.scala 71:109:@25966.4]
  assign _T_73201 = _T_73200[10:0]; // @[Modules.scala 71:109:@25967.4]
  assign buffer_10_713 = $signed(_T_73201); // @[Modules.scala 71:109:@25968.4]
  assign _T_73203 = $signed(buffer_10_644) + $signed(buffer_10_645); // @[Modules.scala 71:109:@25970.4]
  assign _T_73204 = _T_73203[10:0]; // @[Modules.scala 71:109:@25971.4]
  assign buffer_10_714 = $signed(_T_73204); // @[Modules.scala 71:109:@25972.4]
  assign _T_73206 = $signed(buffer_10_646) + $signed(buffer_4_647); // @[Modules.scala 71:109:@25974.4]
  assign _T_73207 = _T_73206[10:0]; // @[Modules.scala 71:109:@25975.4]
  assign buffer_10_715 = $signed(_T_73207); // @[Modules.scala 71:109:@25976.4]
  assign _T_73209 = $signed(buffer_10_648) + $signed(buffer_10_649); // @[Modules.scala 71:109:@25978.4]
  assign _T_73210 = _T_73209[10:0]; // @[Modules.scala 71:109:@25979.4]
  assign buffer_10_716 = $signed(_T_73210); // @[Modules.scala 71:109:@25980.4]
  assign _T_73212 = $signed(buffer_3_650) + $signed(buffer_10_651); // @[Modules.scala 71:109:@25982.4]
  assign _T_73213 = _T_73212[10:0]; // @[Modules.scala 71:109:@25983.4]
  assign buffer_10_717 = $signed(_T_73213); // @[Modules.scala 71:109:@25984.4]
  assign _T_73215 = $signed(buffer_10_652) + $signed(buffer_10_653); // @[Modules.scala 71:109:@25986.4]
  assign _T_73216 = _T_73215[10:0]; // @[Modules.scala 71:109:@25987.4]
  assign buffer_10_718 = $signed(_T_73216); // @[Modules.scala 71:109:@25988.4]
  assign _T_73218 = $signed(buffer_8_654) + $signed(buffer_10_655); // @[Modules.scala 71:109:@25990.4]
  assign _T_73219 = _T_73218[10:0]; // @[Modules.scala 71:109:@25991.4]
  assign buffer_10_719 = $signed(_T_73219); // @[Modules.scala 71:109:@25992.4]
  assign _T_73221 = $signed(buffer_10_656) + $signed(buffer_10_657); // @[Modules.scala 71:109:@25994.4]
  assign _T_73222 = _T_73221[10:0]; // @[Modules.scala 71:109:@25995.4]
  assign buffer_10_720 = $signed(_T_73222); // @[Modules.scala 71:109:@25996.4]
  assign _T_73224 = $signed(buffer_10_658) + $signed(buffer_10_659); // @[Modules.scala 71:109:@25998.4]
  assign _T_73225 = _T_73224[10:0]; // @[Modules.scala 71:109:@25999.4]
  assign buffer_10_721 = $signed(_T_73225); // @[Modules.scala 71:109:@26000.4]
  assign _T_73227 = $signed(buffer_10_660) + $signed(buffer_3_661); // @[Modules.scala 71:109:@26002.4]
  assign _T_73228 = _T_73227[10:0]; // @[Modules.scala 71:109:@26003.4]
  assign buffer_10_722 = $signed(_T_73228); // @[Modules.scala 71:109:@26004.4]
  assign _T_73230 = $signed(buffer_4_662) + $signed(buffer_1_663); // @[Modules.scala 71:109:@26006.4]
  assign _T_73231 = _T_73230[10:0]; // @[Modules.scala 71:109:@26007.4]
  assign buffer_10_723 = $signed(_T_73231); // @[Modules.scala 71:109:@26008.4]
  assign _T_73233 = $signed(buffer_10_664) + $signed(buffer_5_665); // @[Modules.scala 71:109:@26010.4]
  assign _T_73234 = _T_73233[10:0]; // @[Modules.scala 71:109:@26011.4]
  assign buffer_10_724 = $signed(_T_73234); // @[Modules.scala 71:109:@26012.4]
  assign _T_73236 = $signed(buffer_10_666) + $signed(buffer_10_667); // @[Modules.scala 71:109:@26014.4]
  assign _T_73237 = _T_73236[10:0]; // @[Modules.scala 71:109:@26015.4]
  assign buffer_10_725 = $signed(_T_73237); // @[Modules.scala 71:109:@26016.4]
  assign _T_73239 = $signed(buffer_10_668) + $signed(buffer_10_669); // @[Modules.scala 71:109:@26018.4]
  assign _T_73240 = _T_73239[10:0]; // @[Modules.scala 71:109:@26019.4]
  assign buffer_10_726 = $signed(_T_73240); // @[Modules.scala 71:109:@26020.4]
  assign _T_73242 = $signed(buffer_0_593) + $signed(buffer_8_671); // @[Modules.scala 71:109:@26022.4]
  assign _T_73243 = _T_73242[10:0]; // @[Modules.scala 71:109:@26023.4]
  assign buffer_10_727 = $signed(_T_73243); // @[Modules.scala 71:109:@26024.4]
  assign _T_73245 = $signed(buffer_1_672) + $signed(buffer_10_673); // @[Modules.scala 71:109:@26026.4]
  assign _T_73246 = _T_73245[10:0]; // @[Modules.scala 71:109:@26027.4]
  assign buffer_10_728 = $signed(_T_73246); // @[Modules.scala 71:109:@26028.4]
  assign _T_73248 = $signed(buffer_0_593) + $signed(buffer_9_675); // @[Modules.scala 71:109:@26030.4]
  assign _T_73249 = _T_73248[10:0]; // @[Modules.scala 71:109:@26031.4]
  assign buffer_10_729 = $signed(_T_73249); // @[Modules.scala 71:109:@26032.4]
  assign _T_73251 = $signed(buffer_10_676) + $signed(buffer_0_593); // @[Modules.scala 71:109:@26034.4]
  assign _T_73252 = _T_73251[10:0]; // @[Modules.scala 71:109:@26035.4]
  assign buffer_10_730 = $signed(_T_73252); // @[Modules.scala 71:109:@26036.4]
  assign _T_73254 = $signed(buffer_10_678) + $signed(buffer_10_679); // @[Modules.scala 71:109:@26038.4]
  assign _T_73255 = _T_73254[10:0]; // @[Modules.scala 71:109:@26039.4]
  assign buffer_10_731 = $signed(_T_73255); // @[Modules.scala 71:109:@26040.4]
  assign _T_73257 = $signed(buffer_10_680) + $signed(buffer_0_593); // @[Modules.scala 71:109:@26042.4]
  assign _T_73258 = _T_73257[10:0]; // @[Modules.scala 71:109:@26043.4]
  assign buffer_10_732 = $signed(_T_73258); // @[Modules.scala 71:109:@26044.4]
  assign _T_73260 = $signed(buffer_10_682) + $signed(buffer_10_683); // @[Modules.scala 71:109:@26046.4]
  assign _T_73261 = _T_73260[10:0]; // @[Modules.scala 71:109:@26047.4]
  assign buffer_10_733 = $signed(_T_73261); // @[Modules.scala 71:109:@26048.4]
  assign _T_73263 = $signed(buffer_9_684) + $signed(buffer_10_685); // @[Modules.scala 71:109:@26050.4]
  assign _T_73264 = _T_73263[10:0]; // @[Modules.scala 71:109:@26051.4]
  assign buffer_10_734 = $signed(_T_73264); // @[Modules.scala 71:109:@26052.4]
  assign _T_73266 = $signed(buffer_10_686) + $signed(buffer_10_687); // @[Modules.scala 78:156:@26055.4]
  assign _T_73267 = _T_73266[10:0]; // @[Modules.scala 78:156:@26056.4]
  assign buffer_10_736 = $signed(_T_73267); // @[Modules.scala 78:156:@26057.4]
  assign _T_73269 = $signed(buffer_10_736) + $signed(buffer_9_688); // @[Modules.scala 78:156:@26059.4]
  assign _T_73270 = _T_73269[10:0]; // @[Modules.scala 78:156:@26060.4]
  assign buffer_10_737 = $signed(_T_73270); // @[Modules.scala 78:156:@26061.4]
  assign _T_73272 = $signed(buffer_10_737) + $signed(buffer_10_689); // @[Modules.scala 78:156:@26063.4]
  assign _T_73273 = _T_73272[10:0]; // @[Modules.scala 78:156:@26064.4]
  assign buffer_10_738 = $signed(_T_73273); // @[Modules.scala 78:156:@26065.4]
  assign _T_73275 = $signed(buffer_10_738) + $signed(buffer_1_690); // @[Modules.scala 78:156:@26067.4]
  assign _T_73276 = _T_73275[10:0]; // @[Modules.scala 78:156:@26068.4]
  assign buffer_10_739 = $signed(_T_73276); // @[Modules.scala 78:156:@26069.4]
  assign _T_73278 = $signed(buffer_10_739) + $signed(buffer_10_691); // @[Modules.scala 78:156:@26071.4]
  assign _T_73279 = _T_73278[10:0]; // @[Modules.scala 78:156:@26072.4]
  assign buffer_10_740 = $signed(_T_73279); // @[Modules.scala 78:156:@26073.4]
  assign _T_73281 = $signed(buffer_10_740) + $signed(buffer_10_692); // @[Modules.scala 78:156:@26075.4]
  assign _T_73282 = _T_73281[10:0]; // @[Modules.scala 78:156:@26076.4]
  assign buffer_10_741 = $signed(_T_73282); // @[Modules.scala 78:156:@26077.4]
  assign _T_73284 = $signed(buffer_10_741) + $signed(buffer_10_693); // @[Modules.scala 78:156:@26079.4]
  assign _T_73285 = _T_73284[10:0]; // @[Modules.scala 78:156:@26080.4]
  assign buffer_10_742 = $signed(_T_73285); // @[Modules.scala 78:156:@26081.4]
  assign _T_73287 = $signed(buffer_10_742) + $signed(buffer_10_694); // @[Modules.scala 78:156:@26083.4]
  assign _T_73288 = _T_73287[10:0]; // @[Modules.scala 78:156:@26084.4]
  assign buffer_10_743 = $signed(_T_73288); // @[Modules.scala 78:156:@26085.4]
  assign _T_73290 = $signed(buffer_10_743) + $signed(buffer_10_695); // @[Modules.scala 78:156:@26087.4]
  assign _T_73291 = _T_73290[10:0]; // @[Modules.scala 78:156:@26088.4]
  assign buffer_10_744 = $signed(_T_73291); // @[Modules.scala 78:156:@26089.4]
  assign _T_73293 = $signed(buffer_10_744) + $signed(buffer_10_696); // @[Modules.scala 78:156:@26091.4]
  assign _T_73294 = _T_73293[10:0]; // @[Modules.scala 78:156:@26092.4]
  assign buffer_10_745 = $signed(_T_73294); // @[Modules.scala 78:156:@26093.4]
  assign _T_73296 = $signed(buffer_10_745) + $signed(buffer_10_697); // @[Modules.scala 78:156:@26095.4]
  assign _T_73297 = _T_73296[10:0]; // @[Modules.scala 78:156:@26096.4]
  assign buffer_10_746 = $signed(_T_73297); // @[Modules.scala 78:156:@26097.4]
  assign _T_73299 = $signed(buffer_10_746) + $signed(buffer_10_698); // @[Modules.scala 78:156:@26099.4]
  assign _T_73300 = _T_73299[10:0]; // @[Modules.scala 78:156:@26100.4]
  assign buffer_10_747 = $signed(_T_73300); // @[Modules.scala 78:156:@26101.4]
  assign _T_73302 = $signed(buffer_10_747) + $signed(buffer_10_699); // @[Modules.scala 78:156:@26103.4]
  assign _T_73303 = _T_73302[10:0]; // @[Modules.scala 78:156:@26104.4]
  assign buffer_10_748 = $signed(_T_73303); // @[Modules.scala 78:156:@26105.4]
  assign _T_73305 = $signed(buffer_10_748) + $signed(buffer_10_700); // @[Modules.scala 78:156:@26107.4]
  assign _T_73306 = _T_73305[10:0]; // @[Modules.scala 78:156:@26108.4]
  assign buffer_10_749 = $signed(_T_73306); // @[Modules.scala 78:156:@26109.4]
  assign _T_73308 = $signed(buffer_10_749) + $signed(buffer_10_701); // @[Modules.scala 78:156:@26111.4]
  assign _T_73309 = _T_73308[10:0]; // @[Modules.scala 78:156:@26112.4]
  assign buffer_10_750 = $signed(_T_73309); // @[Modules.scala 78:156:@26113.4]
  assign _T_73311 = $signed(buffer_10_750) + $signed(buffer_10_702); // @[Modules.scala 78:156:@26115.4]
  assign _T_73312 = _T_73311[10:0]; // @[Modules.scala 78:156:@26116.4]
  assign buffer_10_751 = $signed(_T_73312); // @[Modules.scala 78:156:@26117.4]
  assign _T_73314 = $signed(buffer_10_751) + $signed(buffer_10_703); // @[Modules.scala 78:156:@26119.4]
  assign _T_73315 = _T_73314[10:0]; // @[Modules.scala 78:156:@26120.4]
  assign buffer_10_752 = $signed(_T_73315); // @[Modules.scala 78:156:@26121.4]
  assign _T_73317 = $signed(buffer_10_752) + $signed(buffer_10_704); // @[Modules.scala 78:156:@26123.4]
  assign _T_73318 = _T_73317[10:0]; // @[Modules.scala 78:156:@26124.4]
  assign buffer_10_753 = $signed(_T_73318); // @[Modules.scala 78:156:@26125.4]
  assign _T_73320 = $signed(buffer_10_753) + $signed(buffer_10_705); // @[Modules.scala 78:156:@26127.4]
  assign _T_73321 = _T_73320[10:0]; // @[Modules.scala 78:156:@26128.4]
  assign buffer_10_754 = $signed(_T_73321); // @[Modules.scala 78:156:@26129.4]
  assign _T_73323 = $signed(buffer_10_754) + $signed(buffer_10_706); // @[Modules.scala 78:156:@26131.4]
  assign _T_73324 = _T_73323[10:0]; // @[Modules.scala 78:156:@26132.4]
  assign buffer_10_755 = $signed(_T_73324); // @[Modules.scala 78:156:@26133.4]
  assign _T_73326 = $signed(buffer_10_755) + $signed(buffer_9_707); // @[Modules.scala 78:156:@26135.4]
  assign _T_73327 = _T_73326[10:0]; // @[Modules.scala 78:156:@26136.4]
  assign buffer_10_756 = $signed(_T_73327); // @[Modules.scala 78:156:@26137.4]
  assign _T_73329 = $signed(buffer_10_756) + $signed(buffer_10_708); // @[Modules.scala 78:156:@26139.4]
  assign _T_73330 = _T_73329[10:0]; // @[Modules.scala 78:156:@26140.4]
  assign buffer_10_757 = $signed(_T_73330); // @[Modules.scala 78:156:@26141.4]
  assign _T_73332 = $signed(buffer_10_757) + $signed(buffer_10_709); // @[Modules.scala 78:156:@26143.4]
  assign _T_73333 = _T_73332[10:0]; // @[Modules.scala 78:156:@26144.4]
  assign buffer_10_758 = $signed(_T_73333); // @[Modules.scala 78:156:@26145.4]
  assign _T_73335 = $signed(buffer_10_758) + $signed(buffer_10_710); // @[Modules.scala 78:156:@26147.4]
  assign _T_73336 = _T_73335[10:0]; // @[Modules.scala 78:156:@26148.4]
  assign buffer_10_759 = $signed(_T_73336); // @[Modules.scala 78:156:@26149.4]
  assign _T_73338 = $signed(buffer_10_759) + $signed(buffer_10_711); // @[Modules.scala 78:156:@26151.4]
  assign _T_73339 = _T_73338[10:0]; // @[Modules.scala 78:156:@26152.4]
  assign buffer_10_760 = $signed(_T_73339); // @[Modules.scala 78:156:@26153.4]
  assign _T_73341 = $signed(buffer_10_760) + $signed(buffer_10_712); // @[Modules.scala 78:156:@26155.4]
  assign _T_73342 = _T_73341[10:0]; // @[Modules.scala 78:156:@26156.4]
  assign buffer_10_761 = $signed(_T_73342); // @[Modules.scala 78:156:@26157.4]
  assign _T_73344 = $signed(buffer_10_761) + $signed(buffer_10_713); // @[Modules.scala 78:156:@26159.4]
  assign _T_73345 = _T_73344[10:0]; // @[Modules.scala 78:156:@26160.4]
  assign buffer_10_762 = $signed(_T_73345); // @[Modules.scala 78:156:@26161.4]
  assign _T_73347 = $signed(buffer_10_762) + $signed(buffer_10_714); // @[Modules.scala 78:156:@26163.4]
  assign _T_73348 = _T_73347[10:0]; // @[Modules.scala 78:156:@26164.4]
  assign buffer_10_763 = $signed(_T_73348); // @[Modules.scala 78:156:@26165.4]
  assign _T_73350 = $signed(buffer_10_763) + $signed(buffer_10_715); // @[Modules.scala 78:156:@26167.4]
  assign _T_73351 = _T_73350[10:0]; // @[Modules.scala 78:156:@26168.4]
  assign buffer_10_764 = $signed(_T_73351); // @[Modules.scala 78:156:@26169.4]
  assign _T_73353 = $signed(buffer_10_764) + $signed(buffer_10_716); // @[Modules.scala 78:156:@26171.4]
  assign _T_73354 = _T_73353[10:0]; // @[Modules.scala 78:156:@26172.4]
  assign buffer_10_765 = $signed(_T_73354); // @[Modules.scala 78:156:@26173.4]
  assign _T_73356 = $signed(buffer_10_765) + $signed(buffer_10_717); // @[Modules.scala 78:156:@26175.4]
  assign _T_73357 = _T_73356[10:0]; // @[Modules.scala 78:156:@26176.4]
  assign buffer_10_766 = $signed(_T_73357); // @[Modules.scala 78:156:@26177.4]
  assign _T_73359 = $signed(buffer_10_766) + $signed(buffer_10_718); // @[Modules.scala 78:156:@26179.4]
  assign _T_73360 = _T_73359[10:0]; // @[Modules.scala 78:156:@26180.4]
  assign buffer_10_767 = $signed(_T_73360); // @[Modules.scala 78:156:@26181.4]
  assign _T_73362 = $signed(buffer_10_767) + $signed(buffer_10_719); // @[Modules.scala 78:156:@26183.4]
  assign _T_73363 = _T_73362[10:0]; // @[Modules.scala 78:156:@26184.4]
  assign buffer_10_768 = $signed(_T_73363); // @[Modules.scala 78:156:@26185.4]
  assign _T_73365 = $signed(buffer_10_768) + $signed(buffer_10_720); // @[Modules.scala 78:156:@26187.4]
  assign _T_73366 = _T_73365[10:0]; // @[Modules.scala 78:156:@26188.4]
  assign buffer_10_769 = $signed(_T_73366); // @[Modules.scala 78:156:@26189.4]
  assign _T_73368 = $signed(buffer_10_769) + $signed(buffer_10_721); // @[Modules.scala 78:156:@26191.4]
  assign _T_73369 = _T_73368[10:0]; // @[Modules.scala 78:156:@26192.4]
  assign buffer_10_770 = $signed(_T_73369); // @[Modules.scala 78:156:@26193.4]
  assign _T_73371 = $signed(buffer_10_770) + $signed(buffer_10_722); // @[Modules.scala 78:156:@26195.4]
  assign _T_73372 = _T_73371[10:0]; // @[Modules.scala 78:156:@26196.4]
  assign buffer_10_771 = $signed(_T_73372); // @[Modules.scala 78:156:@26197.4]
  assign _T_73374 = $signed(buffer_10_771) + $signed(buffer_10_723); // @[Modules.scala 78:156:@26199.4]
  assign _T_73375 = _T_73374[10:0]; // @[Modules.scala 78:156:@26200.4]
  assign buffer_10_772 = $signed(_T_73375); // @[Modules.scala 78:156:@26201.4]
  assign _T_73377 = $signed(buffer_10_772) + $signed(buffer_10_724); // @[Modules.scala 78:156:@26203.4]
  assign _T_73378 = _T_73377[10:0]; // @[Modules.scala 78:156:@26204.4]
  assign buffer_10_773 = $signed(_T_73378); // @[Modules.scala 78:156:@26205.4]
  assign _T_73380 = $signed(buffer_10_773) + $signed(buffer_10_725); // @[Modules.scala 78:156:@26207.4]
  assign _T_73381 = _T_73380[10:0]; // @[Modules.scala 78:156:@26208.4]
  assign buffer_10_774 = $signed(_T_73381); // @[Modules.scala 78:156:@26209.4]
  assign _T_73383 = $signed(buffer_10_774) + $signed(buffer_10_726); // @[Modules.scala 78:156:@26211.4]
  assign _T_73384 = _T_73383[10:0]; // @[Modules.scala 78:156:@26212.4]
  assign buffer_10_775 = $signed(_T_73384); // @[Modules.scala 78:156:@26213.4]
  assign _T_73386 = $signed(buffer_10_775) + $signed(buffer_10_727); // @[Modules.scala 78:156:@26215.4]
  assign _T_73387 = _T_73386[10:0]; // @[Modules.scala 78:156:@26216.4]
  assign buffer_10_776 = $signed(_T_73387); // @[Modules.scala 78:156:@26217.4]
  assign _T_73389 = $signed(buffer_10_776) + $signed(buffer_10_728); // @[Modules.scala 78:156:@26219.4]
  assign _T_73390 = _T_73389[10:0]; // @[Modules.scala 78:156:@26220.4]
  assign buffer_10_777 = $signed(_T_73390); // @[Modules.scala 78:156:@26221.4]
  assign _T_73392 = $signed(buffer_10_777) + $signed(buffer_10_729); // @[Modules.scala 78:156:@26223.4]
  assign _T_73393 = _T_73392[10:0]; // @[Modules.scala 78:156:@26224.4]
  assign buffer_10_778 = $signed(_T_73393); // @[Modules.scala 78:156:@26225.4]
  assign _T_73395 = $signed(buffer_10_778) + $signed(buffer_10_730); // @[Modules.scala 78:156:@26227.4]
  assign _T_73396 = _T_73395[10:0]; // @[Modules.scala 78:156:@26228.4]
  assign buffer_10_779 = $signed(_T_73396); // @[Modules.scala 78:156:@26229.4]
  assign _T_73398 = $signed(buffer_10_779) + $signed(buffer_10_731); // @[Modules.scala 78:156:@26231.4]
  assign _T_73399 = _T_73398[10:0]; // @[Modules.scala 78:156:@26232.4]
  assign buffer_10_780 = $signed(_T_73399); // @[Modules.scala 78:156:@26233.4]
  assign _T_73401 = $signed(buffer_10_780) + $signed(buffer_10_732); // @[Modules.scala 78:156:@26235.4]
  assign _T_73402 = _T_73401[10:0]; // @[Modules.scala 78:156:@26236.4]
  assign buffer_10_781 = $signed(_T_73402); // @[Modules.scala 78:156:@26237.4]
  assign _T_73404 = $signed(buffer_10_781) + $signed(buffer_10_733); // @[Modules.scala 78:156:@26239.4]
  assign _T_73405 = _T_73404[10:0]; // @[Modules.scala 78:156:@26240.4]
  assign buffer_10_782 = $signed(_T_73405); // @[Modules.scala 78:156:@26241.4]
  assign _T_73407 = $signed(buffer_10_782) + $signed(buffer_10_734); // @[Modules.scala 78:156:@26243.4]
  assign _T_73408 = _T_73407[10:0]; // @[Modules.scala 78:156:@26244.4]
  assign buffer_10_783 = $signed(_T_73408); // @[Modules.scala 78:156:@26245.4]
  assign _T_73466 = $signed(io_in_86) + $signed(io_in_87); // @[Modules.scala 37:46:@26333.4]
  assign _T_73467 = _T_73466[4:0]; // @[Modules.scala 37:46:@26334.4]
  assign _T_73468 = $signed(_T_73467); // @[Modules.scala 37:46:@26335.4]
  assign _T_73916 = $signed(buffer_0_8) + $signed(buffer_1_9); // @[Modules.scala 65:57:@26968.4]
  assign _T_73917 = _T_73916[10:0]; // @[Modules.scala 65:57:@26969.4]
  assign buffer_11_396 = $signed(_T_73917); // @[Modules.scala 65:57:@26970.4]
  assign _T_73925 = $signed(buffer_3_14) + $signed(buffer_1_15); // @[Modules.scala 65:57:@26980.4]
  assign _T_73926 = _T_73925[10:0]; // @[Modules.scala 65:57:@26981.4]
  assign buffer_11_399 = $signed(_T_73926); // @[Modules.scala 65:57:@26982.4]
  assign buffer_11_19 = {{6{io_in_39[4]}},io_in_39}; // @[Modules.scala 32:22:@8.4]
  assign _T_73931 = $signed(11'sh0) + $signed(buffer_11_19); // @[Modules.scala 65:57:@26988.4]
  assign _T_73932 = _T_73931[10:0]; // @[Modules.scala 65:57:@26989.4]
  assign buffer_11_401 = $signed(_T_73932); // @[Modules.scala 65:57:@26990.4]
  assign buffer_11_22 = {{6{io_in_44[4]}},io_in_44}; // @[Modules.scala 32:22:@8.4]
  assign buffer_11_23 = {{6{io_in_47[4]}},io_in_47}; // @[Modules.scala 32:22:@8.4]
  assign _T_73937 = $signed(buffer_11_22) + $signed(buffer_11_23); // @[Modules.scala 65:57:@26996.4]
  assign _T_73938 = _T_73937[10:0]; // @[Modules.scala 65:57:@26997.4]
  assign buffer_11_403 = $signed(_T_73938); // @[Modules.scala 65:57:@26998.4]
  assign _T_73943 = $signed(buffer_3_26) + $signed(buffer_1_27); // @[Modules.scala 65:57:@27004.4]
  assign _T_73944 = _T_73943[10:0]; // @[Modules.scala 65:57:@27005.4]
  assign buffer_11_405 = $signed(_T_73944); // @[Modules.scala 65:57:@27006.4]
  assign _T_73946 = $signed(11'sh0) + $signed(buffer_2_29); // @[Modules.scala 65:57:@27008.4]
  assign _T_73947 = _T_73946[10:0]; // @[Modules.scala 65:57:@27009.4]
  assign buffer_11_406 = $signed(_T_73947); // @[Modules.scala 65:57:@27010.4]
  assign _T_73955 = $signed(11'sh0) + $signed(buffer_1_35); // @[Modules.scala 65:57:@27020.4]
  assign _T_73956 = _T_73955[10:0]; // @[Modules.scala 65:57:@27021.4]
  assign buffer_11_409 = $signed(_T_73956); // @[Modules.scala 65:57:@27022.4]
  assign buffer_11_43 = {{6{_T_73468[4]}},_T_73468}; // @[Modules.scala 32:22:@8.4]
  assign _T_73967 = $signed(11'sh0) + $signed(buffer_11_43); // @[Modules.scala 65:57:@27036.4]
  assign _T_73968 = _T_73967[10:0]; // @[Modules.scala 65:57:@27037.4]
  assign buffer_11_413 = $signed(_T_73968); // @[Modules.scala 65:57:@27038.4]
  assign _T_73970 = $signed(buffer_2_44) + $signed(11'sh0); // @[Modules.scala 65:57:@27040.4]
  assign _T_73971 = _T_73970[10:0]; // @[Modules.scala 65:57:@27041.4]
  assign buffer_11_414 = $signed(_T_73971); // @[Modules.scala 65:57:@27042.4]
  assign _T_74006 = $signed(buffer_0_68) + $signed(buffer_3_69); // @[Modules.scala 65:57:@27088.4]
  assign _T_74007 = _T_74006[10:0]; // @[Modules.scala 65:57:@27089.4]
  assign buffer_11_426 = $signed(_T_74007); // @[Modules.scala 65:57:@27090.4]
  assign _T_74009 = $signed(buffer_0_70) + $signed(buffer_2_71); // @[Modules.scala 65:57:@27092.4]
  assign _T_74010 = _T_74009[10:0]; // @[Modules.scala 65:57:@27093.4]
  assign buffer_11_427 = $signed(_T_74010); // @[Modules.scala 65:57:@27094.4]
  assign _T_74027 = $signed(buffer_5_82) + $signed(buffer_1_83); // @[Modules.scala 65:57:@27116.4]
  assign _T_74028 = _T_74027[10:0]; // @[Modules.scala 65:57:@27117.4]
  assign buffer_11_433 = $signed(_T_74028); // @[Modules.scala 65:57:@27118.4]
  assign buffer_11_90 = {{6{io_in_181[4]}},io_in_181}; // @[Modules.scala 32:22:@8.4]
  assign _T_74039 = $signed(buffer_11_90) + $signed(buffer_1_91); // @[Modules.scala 65:57:@27132.4]
  assign _T_74040 = _T_74039[10:0]; // @[Modules.scala 65:57:@27133.4]
  assign buffer_11_437 = $signed(_T_74040); // @[Modules.scala 65:57:@27134.4]
  assign _T_74042 = $signed(buffer_3_92) + $signed(buffer_0_93); // @[Modules.scala 65:57:@27136.4]
  assign _T_74043 = _T_74042[10:0]; // @[Modules.scala 65:57:@27137.4]
  assign buffer_11_438 = $signed(_T_74043); // @[Modules.scala 65:57:@27138.4]
  assign _T_74045 = $signed(buffer_1_94) + $signed(buffer_2_95); // @[Modules.scala 65:57:@27140.4]
  assign _T_74046 = _T_74045[10:0]; // @[Modules.scala 65:57:@27141.4]
  assign buffer_11_439 = $signed(_T_74046); // @[Modules.scala 65:57:@27142.4]
  assign buffer_11_105 = {{6{io_in_211[4]}},io_in_211}; // @[Modules.scala 32:22:@8.4]
  assign _T_74060 = $signed(buffer_0_104) + $signed(buffer_11_105); // @[Modules.scala 65:57:@27160.4]
  assign _T_74061 = _T_74060[10:0]; // @[Modules.scala 65:57:@27161.4]
  assign buffer_11_444 = $signed(_T_74061); // @[Modules.scala 65:57:@27162.4]
  assign _T_74063 = $signed(11'sh0) + $signed(buffer_6_107); // @[Modules.scala 65:57:@27164.4]
  assign _T_74064 = _T_74063[10:0]; // @[Modules.scala 65:57:@27165.4]
  assign buffer_11_445 = $signed(_T_74064); // @[Modules.scala 65:57:@27166.4]
  assign buffer_11_112 = {{6{io_in_224[4]}},io_in_224}; // @[Modules.scala 32:22:@8.4]
  assign _T_74072 = $signed(buffer_11_112) + $signed(11'sh0); // @[Modules.scala 65:57:@27176.4]
  assign _T_74073 = _T_74072[10:0]; // @[Modules.scala 65:57:@27177.4]
  assign buffer_11_448 = $signed(_T_74073); // @[Modules.scala 65:57:@27178.4]
  assign _T_74078 = $signed(11'sh0) + $signed(buffer_7_117); // @[Modules.scala 65:57:@27184.4]
  assign _T_74079 = _T_74078[10:0]; // @[Modules.scala 65:57:@27185.4]
  assign buffer_11_450 = $signed(_T_74079); // @[Modules.scala 65:57:@27186.4]
  assign buffer_11_119 = {{6{io_in_239[4]}},io_in_239}; // @[Modules.scala 32:22:@8.4]
  assign _T_74081 = $signed(buffer_3_118) + $signed(buffer_11_119); // @[Modules.scala 65:57:@27188.4]
  assign _T_74082 = _T_74081[10:0]; // @[Modules.scala 65:57:@27189.4]
  assign buffer_11_451 = $signed(_T_74082); // @[Modules.scala 65:57:@27190.4]
  assign _T_74084 = $signed(buffer_6_120) + $signed(buffer_4_121); // @[Modules.scala 65:57:@27192.4]
  assign _T_74085 = _T_74084[10:0]; // @[Modules.scala 65:57:@27193.4]
  assign buffer_11_452 = $signed(_T_74085); // @[Modules.scala 65:57:@27194.4]
  assign _T_74087 = $signed(buffer_9_122) + $signed(buffer_3_123); // @[Modules.scala 65:57:@27196.4]
  assign _T_74088 = _T_74087[10:0]; // @[Modules.scala 65:57:@27197.4]
  assign buffer_11_453 = $signed(_T_74088); // @[Modules.scala 65:57:@27198.4]
  assign _T_74096 = $signed(11'sh0) + $signed(buffer_4_129); // @[Modules.scala 65:57:@27208.4]
  assign _T_74097 = _T_74096[10:0]; // @[Modules.scala 65:57:@27209.4]
  assign buffer_11_456 = $signed(_T_74097); // @[Modules.scala 65:57:@27210.4]
  assign _T_74102 = $signed(buffer_5_132) + $signed(11'sh0); // @[Modules.scala 65:57:@27216.4]
  assign _T_74103 = _T_74102[10:0]; // @[Modules.scala 65:57:@27217.4]
  assign buffer_11_458 = $signed(_T_74103); // @[Modules.scala 65:57:@27218.4]
  assign buffer_11_135 = {{6{io_in_271[4]}},io_in_271}; // @[Modules.scala 32:22:@8.4]
  assign _T_74105 = $signed(11'sh0) + $signed(buffer_11_135); // @[Modules.scala 65:57:@27220.4]
  assign _T_74106 = _T_74105[10:0]; // @[Modules.scala 65:57:@27221.4]
  assign buffer_11_459 = $signed(_T_74106); // @[Modules.scala 65:57:@27222.4]
  assign _T_74114 = $signed(buffer_3_140) + $signed(11'sh0); // @[Modules.scala 65:57:@27232.4]
  assign _T_74115 = _T_74114[10:0]; // @[Modules.scala 65:57:@27233.4]
  assign buffer_11_462 = $signed(_T_74115); // @[Modules.scala 65:57:@27234.4]
  assign _T_74117 = $signed(11'sh0) + $signed(buffer_7_143); // @[Modules.scala 65:57:@27236.4]
  assign _T_74118 = _T_74117[10:0]; // @[Modules.scala 65:57:@27237.4]
  assign buffer_11_463 = $signed(_T_74118); // @[Modules.scala 65:57:@27238.4]
  assign _T_74138 = $signed(buffer_6_156) + $signed(buffer_2_157); // @[Modules.scala 65:57:@27264.4]
  assign _T_74139 = _T_74138[10:0]; // @[Modules.scala 65:57:@27265.4]
  assign buffer_11_470 = $signed(_T_74139); // @[Modules.scala 65:57:@27266.4]
  assign _T_74144 = $signed(buffer_1_160) + $signed(buffer_5_161); // @[Modules.scala 65:57:@27272.4]
  assign _T_74145 = _T_74144[10:0]; // @[Modules.scala 65:57:@27273.4]
  assign buffer_11_472 = $signed(_T_74145); // @[Modules.scala 65:57:@27274.4]
  assign _T_74174 = $signed(buffer_1_180) + $signed(buffer_8_181); // @[Modules.scala 65:57:@27312.4]
  assign _T_74175 = _T_74174[10:0]; // @[Modules.scala 65:57:@27313.4]
  assign buffer_11_482 = $signed(_T_74175); // @[Modules.scala 65:57:@27314.4]
  assign buffer_11_185 = {{6{io_in_371[4]}},io_in_371}; // @[Modules.scala 32:22:@8.4]
  assign _T_74180 = $signed(11'sh0) + $signed(buffer_11_185); // @[Modules.scala 65:57:@27320.4]
  assign _T_74181 = _T_74180[10:0]; // @[Modules.scala 65:57:@27321.4]
  assign buffer_11_484 = $signed(_T_74181); // @[Modules.scala 65:57:@27322.4]
  assign buffer_11_186 = {{6{io_in_373[4]}},io_in_373}; // @[Modules.scala 32:22:@8.4]
  assign _T_74183 = $signed(buffer_11_186) + $signed(11'sh0); // @[Modules.scala 65:57:@27324.4]
  assign _T_74184 = _T_74183[10:0]; // @[Modules.scala 65:57:@27325.4]
  assign buffer_11_485 = $signed(_T_74184); // @[Modules.scala 65:57:@27326.4]
  assign _T_74195 = $signed(buffer_5_194) + $signed(buffer_4_195); // @[Modules.scala 65:57:@27340.4]
  assign _T_74196 = _T_74195[10:0]; // @[Modules.scala 65:57:@27341.4]
  assign buffer_11_489 = $signed(_T_74196); // @[Modules.scala 65:57:@27342.4]
  assign _T_74204 = $signed(11'sh0) + $signed(buffer_3_201); // @[Modules.scala 65:57:@27352.4]
  assign _T_74205 = _T_74204[10:0]; // @[Modules.scala 65:57:@27353.4]
  assign buffer_11_492 = $signed(_T_74205); // @[Modules.scala 65:57:@27354.4]
  assign _T_74219 = $signed(buffer_3_210) + $signed(buffer_1_211); // @[Modules.scala 65:57:@27372.4]
  assign _T_74220 = _T_74219[10:0]; // @[Modules.scala 65:57:@27373.4]
  assign buffer_11_497 = $signed(_T_74220); // @[Modules.scala 65:57:@27374.4]
  assign buffer_11_214 = {{6{io_in_429[4]}},io_in_429}; // @[Modules.scala 32:22:@8.4]
  assign _T_74225 = $signed(buffer_11_214) + $signed(11'sh0); // @[Modules.scala 65:57:@27380.4]
  assign _T_74226 = _T_74225[10:0]; // @[Modules.scala 65:57:@27381.4]
  assign buffer_11_499 = $signed(_T_74226); // @[Modules.scala 65:57:@27382.4]
  assign buffer_11_217 = {{6{io_in_434[4]}},io_in_434}; // @[Modules.scala 32:22:@8.4]
  assign _T_74228 = $signed(buffer_0_216) + $signed(buffer_11_217); // @[Modules.scala 65:57:@27384.4]
  assign _T_74229 = _T_74228[10:0]; // @[Modules.scala 65:57:@27385.4]
  assign buffer_11_500 = $signed(_T_74229); // @[Modules.scala 65:57:@27386.4]
  assign buffer_11_225 = {{6{io_in_450[4]}},io_in_450}; // @[Modules.scala 32:22:@8.4]
  assign _T_74240 = $signed(buffer_1_224) + $signed(buffer_11_225); // @[Modules.scala 65:57:@27400.4]
  assign _T_74241 = _T_74240[10:0]; // @[Modules.scala 65:57:@27401.4]
  assign buffer_11_504 = $signed(_T_74241); // @[Modules.scala 65:57:@27402.4]
  assign _T_74246 = $signed(buffer_1_228) + $signed(11'sh0); // @[Modules.scala 65:57:@27408.4]
  assign _T_74247 = _T_74246[10:0]; // @[Modules.scala 65:57:@27409.4]
  assign buffer_11_506 = $signed(_T_74247); // @[Modules.scala 65:57:@27410.4]
  assign buffer_11_235 = {{6{io_in_471[4]}},io_in_471}; // @[Modules.scala 32:22:@8.4]
  assign _T_74255 = $signed(11'sh0) + $signed(buffer_11_235); // @[Modules.scala 65:57:@27420.4]
  assign _T_74256 = _T_74255[10:0]; // @[Modules.scala 65:57:@27421.4]
  assign buffer_11_509 = $signed(_T_74256); // @[Modules.scala 65:57:@27422.4]
  assign _T_74261 = $signed(buffer_1_238) + $signed(11'sh0); // @[Modules.scala 65:57:@27428.4]
  assign _T_74262 = _T_74261[10:0]; // @[Modules.scala 65:57:@27429.4]
  assign buffer_11_511 = $signed(_T_74262); // @[Modules.scala 65:57:@27430.4]
  assign buffer_11_240 = {{6{io_in_481[4]}},io_in_481}; // @[Modules.scala 32:22:@8.4]
  assign _T_74264 = $signed(buffer_11_240) + $signed(buffer_3_241); // @[Modules.scala 65:57:@27432.4]
  assign _T_74265 = _T_74264[10:0]; // @[Modules.scala 65:57:@27433.4]
  assign buffer_11_512 = $signed(_T_74265); // @[Modules.scala 65:57:@27434.4]
  assign buffer_11_249 = {{6{io_in_499[4]}},io_in_499}; // @[Modules.scala 32:22:@8.4]
  assign _T_74276 = $signed(11'sh0) + $signed(buffer_11_249); // @[Modules.scala 65:57:@27448.4]
  assign _T_74277 = _T_74276[10:0]; // @[Modules.scala 65:57:@27449.4]
  assign buffer_11_516 = $signed(_T_74277); // @[Modules.scala 65:57:@27450.4]
  assign _T_74288 = $signed(buffer_0_256) + $signed(buffer_4_257); // @[Modules.scala 65:57:@27464.4]
  assign _T_74289 = _T_74288[10:0]; // @[Modules.scala 65:57:@27465.4]
  assign buffer_11_520 = $signed(_T_74289); // @[Modules.scala 65:57:@27466.4]
  assign buffer_11_258 = {{6{io_in_517[4]}},io_in_517}; // @[Modules.scala 32:22:@8.4]
  assign _T_74291 = $signed(buffer_11_258) + $signed(11'sh0); // @[Modules.scala 65:57:@27468.4]
  assign _T_74292 = _T_74291[10:0]; // @[Modules.scala 65:57:@27469.4]
  assign buffer_11_521 = $signed(_T_74292); // @[Modules.scala 65:57:@27470.4]
  assign _T_74297 = $signed(buffer_7_262) + $signed(buffer_1_263); // @[Modules.scala 65:57:@27476.4]
  assign _T_74298 = _T_74297[10:0]; // @[Modules.scala 65:57:@27477.4]
  assign buffer_11_523 = $signed(_T_74298); // @[Modules.scala 65:57:@27478.4]
  assign _T_74309 = $signed(buffer_1_270) + $signed(buffer_0_271); // @[Modules.scala 65:57:@27492.4]
  assign _T_74310 = _T_74309[10:0]; // @[Modules.scala 65:57:@27493.4]
  assign buffer_11_527 = $signed(_T_74310); // @[Modules.scala 65:57:@27494.4]
  assign _T_74312 = $signed(buffer_1_272) + $signed(11'sh0); // @[Modules.scala 65:57:@27496.4]
  assign _T_74313 = _T_74312[10:0]; // @[Modules.scala 65:57:@27497.4]
  assign buffer_11_528 = $signed(_T_74313); // @[Modules.scala 65:57:@27498.4]
  assign _T_74318 = $signed(11'sh0) + $signed(buffer_3_277); // @[Modules.scala 65:57:@27504.4]
  assign _T_74319 = _T_74318[10:0]; // @[Modules.scala 65:57:@27505.4]
  assign buffer_11_530 = $signed(_T_74319); // @[Modules.scala 65:57:@27506.4]
  assign buffer_11_281 = {{6{io_in_562[4]}},io_in_562}; // @[Modules.scala 32:22:@8.4]
  assign _T_74324 = $signed(11'sh0) + $signed(buffer_11_281); // @[Modules.scala 65:57:@27512.4]
  assign _T_74325 = _T_74324[10:0]; // @[Modules.scala 65:57:@27513.4]
  assign buffer_11_532 = $signed(_T_74325); // @[Modules.scala 65:57:@27514.4]
  assign _T_74333 = $signed(buffer_3_286) + $signed(11'sh0); // @[Modules.scala 65:57:@27524.4]
  assign _T_74334 = _T_74333[10:0]; // @[Modules.scala 65:57:@27525.4]
  assign buffer_11_535 = $signed(_T_74334); // @[Modules.scala 65:57:@27526.4]
  assign _T_74339 = $signed(11'sh0) + $signed(buffer_3_291); // @[Modules.scala 65:57:@27532.4]
  assign _T_74340 = _T_74339[10:0]; // @[Modules.scala 65:57:@27533.4]
  assign buffer_11_537 = $signed(_T_74340); // @[Modules.scala 65:57:@27534.4]
  assign _T_74348 = $signed(11'sh0) + $signed(buffer_3_297); // @[Modules.scala 65:57:@27544.4]
  assign _T_74349 = _T_74348[10:0]; // @[Modules.scala 65:57:@27545.4]
  assign buffer_11_540 = $signed(_T_74349); // @[Modules.scala 65:57:@27546.4]
  assign _T_74357 = $signed(buffer_0_302) + $signed(buffer_8_303); // @[Modules.scala 65:57:@27556.4]
  assign _T_74358 = _T_74357[10:0]; // @[Modules.scala 65:57:@27557.4]
  assign buffer_11_543 = $signed(_T_74358); // @[Modules.scala 65:57:@27558.4]
  assign buffer_11_310 = {{6{io_in_621[4]}},io_in_621}; // @[Modules.scala 32:22:@8.4]
  assign _T_74369 = $signed(buffer_11_310) + $signed(buffer_7_311); // @[Modules.scala 65:57:@27572.4]
  assign _T_74370 = _T_74369[10:0]; // @[Modules.scala 65:57:@27573.4]
  assign buffer_11_547 = $signed(_T_74370); // @[Modules.scala 65:57:@27574.4]
  assign _T_74372 = $signed(11'sh0) + $signed(buffer_3_313); // @[Modules.scala 65:57:@27576.4]
  assign _T_74373 = _T_74372[10:0]; // @[Modules.scala 65:57:@27577.4]
  assign buffer_11_548 = $signed(_T_74373); // @[Modules.scala 65:57:@27578.4]
  assign _T_74384 = $signed(11'sh0) + $signed(buffer_3_321); // @[Modules.scala 65:57:@27592.4]
  assign _T_74385 = _T_74384[10:0]; // @[Modules.scala 65:57:@27593.4]
  assign buffer_11_552 = $signed(_T_74385); // @[Modules.scala 65:57:@27594.4]
  assign _T_74393 = $signed(11'sh0) + $signed(buffer_8_327); // @[Modules.scala 65:57:@27604.4]
  assign _T_74394 = _T_74393[10:0]; // @[Modules.scala 65:57:@27605.4]
  assign buffer_11_555 = $signed(_T_74394); // @[Modules.scala 65:57:@27606.4]
  assign _T_74423 = $signed(buffer_0_346) + $signed(11'sh0); // @[Modules.scala 65:57:@27644.4]
  assign _T_74424 = _T_74423[10:0]; // @[Modules.scala 65:57:@27645.4]
  assign buffer_11_565 = $signed(_T_74424); // @[Modules.scala 65:57:@27646.4]
  assign _T_74429 = $signed(buffer_5_350) + $signed(buffer_1_351); // @[Modules.scala 65:57:@27652.4]
  assign _T_74430 = _T_74429[10:0]; // @[Modules.scala 65:57:@27653.4]
  assign buffer_11_567 = $signed(_T_74430); // @[Modules.scala 65:57:@27654.4]
  assign buffer_11_361 = {{6{io_in_723[4]}},io_in_723}; // @[Modules.scala 32:22:@8.4]
  assign _T_74444 = $signed(11'sh0) + $signed(buffer_11_361); // @[Modules.scala 65:57:@27672.4]
  assign _T_74445 = _T_74444[10:0]; // @[Modules.scala 65:57:@27673.4]
  assign buffer_11_572 = $signed(_T_74445); // @[Modules.scala 65:57:@27674.4]
  assign _T_74471 = $signed(11'sh0) + $signed(buffer_9_379); // @[Modules.scala 65:57:@27708.4]
  assign _T_74472 = _T_74471[10:0]; // @[Modules.scala 65:57:@27709.4]
  assign buffer_11_581 = $signed(_T_74472); // @[Modules.scala 65:57:@27710.4]
  assign _T_74492 = $signed(buffer_3_392) + $signed(buffer_6_393); // @[Modules.scala 68:83:@27736.4]
  assign _T_74493 = _T_74492[10:0]; // @[Modules.scala 68:83:@27737.4]
  assign buffer_11_588 = $signed(_T_74493); // @[Modules.scala 68:83:@27738.4]
  assign _T_74495 = $signed(buffer_10_394) + $signed(buffer_1_395); // @[Modules.scala 68:83:@27740.4]
  assign _T_74496 = _T_74495[10:0]; // @[Modules.scala 68:83:@27741.4]
  assign buffer_11_589 = $signed(_T_74496); // @[Modules.scala 68:83:@27742.4]
  assign _T_74498 = $signed(buffer_11_396) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27744.4]
  assign _T_74499 = _T_74498[10:0]; // @[Modules.scala 68:83:@27745.4]
  assign buffer_11_590 = $signed(_T_74499); // @[Modules.scala 68:83:@27746.4]
  assign _T_74501 = $signed(buffer_0_398) + $signed(buffer_11_399); // @[Modules.scala 68:83:@27748.4]
  assign _T_74502 = _T_74501[10:0]; // @[Modules.scala 68:83:@27749.4]
  assign buffer_11_591 = $signed(_T_74502); // @[Modules.scala 68:83:@27750.4]
  assign _T_74504 = $signed(buffer_1_400) + $signed(buffer_11_401); // @[Modules.scala 68:83:@27752.4]
  assign _T_74505 = _T_74504[10:0]; // @[Modules.scala 68:83:@27753.4]
  assign buffer_11_592 = $signed(_T_74505); // @[Modules.scala 68:83:@27754.4]
  assign _T_74507 = $signed(buffer_2_402) + $signed(buffer_11_403); // @[Modules.scala 68:83:@27756.4]
  assign _T_74508 = _T_74507[10:0]; // @[Modules.scala 68:83:@27757.4]
  assign buffer_11_593 = $signed(_T_74508); // @[Modules.scala 68:83:@27758.4]
  assign _T_74510 = $signed(buffer_1_404) + $signed(buffer_11_405); // @[Modules.scala 68:83:@27760.4]
  assign _T_74511 = _T_74510[10:0]; // @[Modules.scala 68:83:@27761.4]
  assign buffer_11_594 = $signed(_T_74511); // @[Modules.scala 68:83:@27762.4]
  assign _T_74513 = $signed(buffer_11_406) + $signed(buffer_1_407); // @[Modules.scala 68:83:@27764.4]
  assign _T_74514 = _T_74513[10:0]; // @[Modules.scala 68:83:@27765.4]
  assign buffer_11_595 = $signed(_T_74514); // @[Modules.scala 68:83:@27766.4]
  assign _T_74516 = $signed(buffer_0_395) + $signed(buffer_11_409); // @[Modules.scala 68:83:@27768.4]
  assign _T_74517 = _T_74516[10:0]; // @[Modules.scala 68:83:@27769.4]
  assign buffer_11_596 = $signed(_T_74517); // @[Modules.scala 68:83:@27770.4]
  assign _T_74522 = $signed(buffer_0_412) + $signed(buffer_11_413); // @[Modules.scala 68:83:@27776.4]
  assign _T_74523 = _T_74522[10:0]; // @[Modules.scala 68:83:@27777.4]
  assign buffer_11_598 = $signed(_T_74523); // @[Modules.scala 68:83:@27778.4]
  assign _T_74525 = $signed(buffer_11_414) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27780.4]
  assign _T_74526 = _T_74525[10:0]; // @[Modules.scala 68:83:@27781.4]
  assign buffer_11_599 = $signed(_T_74526); // @[Modules.scala 68:83:@27782.4]
  assign _T_74537 = $signed(buffer_0_395) + $signed(buffer_7_423); // @[Modules.scala 68:83:@27796.4]
  assign _T_74538 = _T_74537[10:0]; // @[Modules.scala 68:83:@27797.4]
  assign buffer_11_603 = $signed(_T_74538); // @[Modules.scala 68:83:@27798.4]
  assign _T_74540 = $signed(buffer_0_395) + $signed(buffer_7_425); // @[Modules.scala 68:83:@27800.4]
  assign _T_74541 = _T_74540[10:0]; // @[Modules.scala 68:83:@27801.4]
  assign buffer_11_604 = $signed(_T_74541); // @[Modules.scala 68:83:@27802.4]
  assign _T_74543 = $signed(buffer_11_426) + $signed(buffer_11_427); // @[Modules.scala 68:83:@27804.4]
  assign _T_74544 = _T_74543[10:0]; // @[Modules.scala 68:83:@27805.4]
  assign buffer_11_605 = $signed(_T_74544); // @[Modules.scala 68:83:@27806.4]
  assign _T_74549 = $signed(buffer_10_430) + $signed(buffer_4_431); // @[Modules.scala 68:83:@27812.4]
  assign _T_74550 = _T_74549[10:0]; // @[Modules.scala 68:83:@27813.4]
  assign buffer_11_607 = $signed(_T_74550); // @[Modules.scala 68:83:@27814.4]
  assign _T_74552 = $signed(buffer_2_432) + $signed(buffer_11_433); // @[Modules.scala 68:83:@27816.4]
  assign _T_74553 = _T_74552[10:0]; // @[Modules.scala 68:83:@27817.4]
  assign buffer_11_608 = $signed(_T_74553); // @[Modules.scala 68:83:@27818.4]
  assign _T_74555 = $signed(buffer_4_434) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27820.4]
  assign _T_74556 = _T_74555[10:0]; // @[Modules.scala 68:83:@27821.4]
  assign buffer_11_609 = $signed(_T_74556); // @[Modules.scala 68:83:@27822.4]
  assign _T_74558 = $signed(buffer_0_395) + $signed(buffer_11_437); // @[Modules.scala 68:83:@27824.4]
  assign _T_74559 = _T_74558[10:0]; // @[Modules.scala 68:83:@27825.4]
  assign buffer_11_610 = $signed(_T_74559); // @[Modules.scala 68:83:@27826.4]
  assign _T_74561 = $signed(buffer_11_438) + $signed(buffer_11_439); // @[Modules.scala 68:83:@27828.4]
  assign _T_74562 = _T_74561[10:0]; // @[Modules.scala 68:83:@27829.4]
  assign buffer_11_611 = $signed(_T_74562); // @[Modules.scala 68:83:@27830.4]
  assign _T_74564 = $signed(buffer_2_440) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27832.4]
  assign _T_74565 = _T_74564[10:0]; // @[Modules.scala 68:83:@27833.4]
  assign buffer_11_612 = $signed(_T_74565); // @[Modules.scala 68:83:@27834.4]
  assign _T_74567 = $signed(buffer_0_395) + $signed(buffer_1_443); // @[Modules.scala 68:83:@27836.4]
  assign _T_74568 = _T_74567[10:0]; // @[Modules.scala 68:83:@27837.4]
  assign buffer_11_613 = $signed(_T_74568); // @[Modules.scala 68:83:@27838.4]
  assign _T_74570 = $signed(buffer_11_444) + $signed(buffer_11_445); // @[Modules.scala 68:83:@27840.4]
  assign _T_74571 = _T_74570[10:0]; // @[Modules.scala 68:83:@27841.4]
  assign buffer_11_614 = $signed(_T_74571); // @[Modules.scala 68:83:@27842.4]
  assign _T_74576 = $signed(buffer_11_448) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27848.4]
  assign _T_74577 = _T_74576[10:0]; // @[Modules.scala 68:83:@27849.4]
  assign buffer_11_616 = $signed(_T_74577); // @[Modules.scala 68:83:@27850.4]
  assign _T_74579 = $signed(buffer_11_450) + $signed(buffer_11_451); // @[Modules.scala 68:83:@27852.4]
  assign _T_74580 = _T_74579[10:0]; // @[Modules.scala 68:83:@27853.4]
  assign buffer_11_617 = $signed(_T_74580); // @[Modules.scala 68:83:@27854.4]
  assign _T_74582 = $signed(buffer_11_452) + $signed(buffer_11_453); // @[Modules.scala 68:83:@27856.4]
  assign _T_74583 = _T_74582[10:0]; // @[Modules.scala 68:83:@27857.4]
  assign buffer_11_618 = $signed(_T_74583); // @[Modules.scala 68:83:@27858.4]
  assign _T_74585 = $signed(buffer_1_454) + $signed(buffer_8_455); // @[Modules.scala 68:83:@27860.4]
  assign _T_74586 = _T_74585[10:0]; // @[Modules.scala 68:83:@27861.4]
  assign buffer_11_619 = $signed(_T_74586); // @[Modules.scala 68:83:@27862.4]
  assign _T_74588 = $signed(buffer_11_456) + $signed(buffer_6_457); // @[Modules.scala 68:83:@27864.4]
  assign _T_74589 = _T_74588[10:0]; // @[Modules.scala 68:83:@27865.4]
  assign buffer_11_620 = $signed(_T_74589); // @[Modules.scala 68:83:@27866.4]
  assign _T_74591 = $signed(buffer_11_458) + $signed(buffer_11_459); // @[Modules.scala 68:83:@27868.4]
  assign _T_74592 = _T_74591[10:0]; // @[Modules.scala 68:83:@27869.4]
  assign buffer_11_621 = $signed(_T_74592); // @[Modules.scala 68:83:@27870.4]
  assign _T_74597 = $signed(buffer_11_462) + $signed(buffer_11_463); // @[Modules.scala 68:83:@27876.4]
  assign _T_74598 = _T_74597[10:0]; // @[Modules.scala 68:83:@27877.4]
  assign buffer_11_623 = $signed(_T_74598); // @[Modules.scala 68:83:@27878.4]
  assign _T_74600 = $signed(buffer_2_464) + $signed(buffer_1_465); // @[Modules.scala 68:83:@27880.4]
  assign _T_74601 = _T_74600[10:0]; // @[Modules.scala 68:83:@27881.4]
  assign buffer_11_624 = $signed(_T_74601); // @[Modules.scala 68:83:@27882.4]
  assign _T_74609 = $signed(buffer_11_470) + $signed(buffer_0_471); // @[Modules.scala 68:83:@27892.4]
  assign _T_74610 = _T_74609[10:0]; // @[Modules.scala 68:83:@27893.4]
  assign buffer_11_627 = $signed(_T_74610); // @[Modules.scala 68:83:@27894.4]
  assign _T_74612 = $signed(buffer_11_472) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27896.4]
  assign _T_74613 = _T_74612[10:0]; // @[Modules.scala 68:83:@27897.4]
  assign buffer_11_628 = $signed(_T_74613); // @[Modules.scala 68:83:@27898.4]
  assign _T_74624 = $signed(buffer_8_480) + $signed(buffer_1_481); // @[Modules.scala 68:83:@27912.4]
  assign _T_74625 = _T_74624[10:0]; // @[Modules.scala 68:83:@27913.4]
  assign buffer_11_632 = $signed(_T_74625); // @[Modules.scala 68:83:@27914.4]
  assign _T_74627 = $signed(buffer_11_482) + $signed(buffer_4_483); // @[Modules.scala 68:83:@27916.4]
  assign _T_74628 = _T_74627[10:0]; // @[Modules.scala 68:83:@27917.4]
  assign buffer_11_633 = $signed(_T_74628); // @[Modules.scala 68:83:@27918.4]
  assign _T_74630 = $signed(buffer_11_484) + $signed(buffer_11_485); // @[Modules.scala 68:83:@27920.4]
  assign _T_74631 = _T_74630[10:0]; // @[Modules.scala 68:83:@27921.4]
  assign buffer_11_634 = $signed(_T_74631); // @[Modules.scala 68:83:@27922.4]
  assign _T_74633 = $signed(buffer_5_486) + $signed(buffer_7_487); // @[Modules.scala 68:83:@27924.4]
  assign _T_74634 = _T_74633[10:0]; // @[Modules.scala 68:83:@27925.4]
  assign buffer_11_635 = $signed(_T_74634); // @[Modules.scala 68:83:@27926.4]
  assign _T_74636 = $signed(buffer_8_488) + $signed(buffer_11_489); // @[Modules.scala 68:83:@27928.4]
  assign _T_74637 = _T_74636[10:0]; // @[Modules.scala 68:83:@27929.4]
  assign buffer_11_636 = $signed(_T_74637); // @[Modules.scala 68:83:@27930.4]
  assign _T_74642 = $signed(buffer_11_492) + $signed(buffer_0_493); // @[Modules.scala 68:83:@27936.4]
  assign _T_74643 = _T_74642[10:0]; // @[Modules.scala 68:83:@27937.4]
  assign buffer_11_638 = $signed(_T_74643); // @[Modules.scala 68:83:@27938.4]
  assign _T_74648 = $signed(buffer_0_395) + $signed(buffer_11_497); // @[Modules.scala 68:83:@27944.4]
  assign _T_74649 = _T_74648[10:0]; // @[Modules.scala 68:83:@27945.4]
  assign buffer_11_640 = $signed(_T_74649); // @[Modules.scala 68:83:@27946.4]
  assign _T_74651 = $signed(buffer_0_395) + $signed(buffer_11_499); // @[Modules.scala 68:83:@27948.4]
  assign _T_74652 = _T_74651[10:0]; // @[Modules.scala 68:83:@27949.4]
  assign buffer_11_641 = $signed(_T_74652); // @[Modules.scala 68:83:@27950.4]
  assign _T_74654 = $signed(buffer_11_500) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27952.4]
  assign _T_74655 = _T_74654[10:0]; // @[Modules.scala 68:83:@27953.4]
  assign buffer_11_642 = $signed(_T_74655); // @[Modules.scala 68:83:@27954.4]
  assign _T_74660 = $signed(buffer_11_504) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27960.4]
  assign _T_74661 = _T_74660[10:0]; // @[Modules.scala 68:83:@27961.4]
  assign buffer_11_644 = $signed(_T_74661); // @[Modules.scala 68:83:@27962.4]
  assign _T_74663 = $signed(buffer_11_506) + $signed(buffer_5_507); // @[Modules.scala 68:83:@27964.4]
  assign _T_74664 = _T_74663[10:0]; // @[Modules.scala 68:83:@27965.4]
  assign buffer_11_645 = $signed(_T_74664); // @[Modules.scala 68:83:@27966.4]
  assign _T_74666 = $signed(buffer_0_395) + $signed(buffer_11_509); // @[Modules.scala 68:83:@27968.4]
  assign _T_74667 = _T_74666[10:0]; // @[Modules.scala 68:83:@27969.4]
  assign buffer_11_646 = $signed(_T_74667); // @[Modules.scala 68:83:@27970.4]
  assign _T_74669 = $signed(buffer_0_395) + $signed(buffer_11_511); // @[Modules.scala 68:83:@27972.4]
  assign _T_74670 = _T_74669[10:0]; // @[Modules.scala 68:83:@27973.4]
  assign buffer_11_647 = $signed(_T_74670); // @[Modules.scala 68:83:@27974.4]
  assign _T_74672 = $signed(buffer_11_512) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27976.4]
  assign _T_74673 = _T_74672[10:0]; // @[Modules.scala 68:83:@27977.4]
  assign buffer_11_648 = $signed(_T_74673); // @[Modules.scala 68:83:@27978.4]
  assign _T_74675 = $signed(buffer_9_514) + $signed(buffer_5_515); // @[Modules.scala 68:83:@27980.4]
  assign _T_74676 = _T_74675[10:0]; // @[Modules.scala 68:83:@27981.4]
  assign buffer_11_649 = $signed(_T_74676); // @[Modules.scala 68:83:@27982.4]
  assign _T_74678 = $signed(buffer_11_516) + $signed(buffer_0_395); // @[Modules.scala 68:83:@27984.4]
  assign _T_74679 = _T_74678[10:0]; // @[Modules.scala 68:83:@27985.4]
  assign buffer_11_650 = $signed(_T_74679); // @[Modules.scala 68:83:@27986.4]
  assign _T_74681 = $signed(buffer_0_395) + $signed(buffer_8_519); // @[Modules.scala 68:83:@27988.4]
  assign _T_74682 = _T_74681[10:0]; // @[Modules.scala 68:83:@27989.4]
  assign buffer_11_651 = $signed(_T_74682); // @[Modules.scala 68:83:@27990.4]
  assign _T_74684 = $signed(buffer_11_520) + $signed(buffer_11_521); // @[Modules.scala 68:83:@27992.4]
  assign _T_74685 = _T_74684[10:0]; // @[Modules.scala 68:83:@27993.4]
  assign buffer_11_652 = $signed(_T_74685); // @[Modules.scala 68:83:@27994.4]
  assign _T_74687 = $signed(buffer_0_395) + $signed(buffer_11_523); // @[Modules.scala 68:83:@27996.4]
  assign _T_74688 = _T_74687[10:0]; // @[Modules.scala 68:83:@27997.4]
  assign buffer_11_653 = $signed(_T_74688); // @[Modules.scala 68:83:@27998.4]
  assign _T_74693 = $signed(buffer_0_395) + $signed(buffer_11_527); // @[Modules.scala 68:83:@28004.4]
  assign _T_74694 = _T_74693[10:0]; // @[Modules.scala 68:83:@28005.4]
  assign buffer_11_655 = $signed(_T_74694); // @[Modules.scala 68:83:@28006.4]
  assign _T_74696 = $signed(buffer_11_528) + $signed(buffer_0_395); // @[Modules.scala 68:83:@28008.4]
  assign _T_74697 = _T_74696[10:0]; // @[Modules.scala 68:83:@28009.4]
  assign buffer_11_656 = $signed(_T_74697); // @[Modules.scala 68:83:@28010.4]
  assign _T_74699 = $signed(buffer_11_530) + $signed(buffer_2_531); // @[Modules.scala 68:83:@28012.4]
  assign _T_74700 = _T_74699[10:0]; // @[Modules.scala 68:83:@28013.4]
  assign buffer_11_657 = $signed(_T_74700); // @[Modules.scala 68:83:@28014.4]
  assign _T_74702 = $signed(buffer_11_532) + $signed(buffer_7_533); // @[Modules.scala 68:83:@28016.4]
  assign _T_74703 = _T_74702[10:0]; // @[Modules.scala 68:83:@28017.4]
  assign buffer_11_658 = $signed(_T_74703); // @[Modules.scala 68:83:@28018.4]
  assign _T_74705 = $signed(buffer_1_534) + $signed(buffer_11_535); // @[Modules.scala 68:83:@28020.4]
  assign _T_74706 = _T_74705[10:0]; // @[Modules.scala 68:83:@28021.4]
  assign buffer_11_659 = $signed(_T_74706); // @[Modules.scala 68:83:@28022.4]
  assign _T_74708 = $signed(buffer_0_395) + $signed(buffer_11_537); // @[Modules.scala 68:83:@28024.4]
  assign _T_74709 = _T_74708[10:0]; // @[Modules.scala 68:83:@28025.4]
  assign buffer_11_660 = $signed(_T_74709); // @[Modules.scala 68:83:@28026.4]
  assign _T_74711 = $signed(buffer_1_538) + $signed(buffer_0_395); // @[Modules.scala 68:83:@28028.4]
  assign _T_74712 = _T_74711[10:0]; // @[Modules.scala 68:83:@28029.4]
  assign buffer_11_661 = $signed(_T_74712); // @[Modules.scala 68:83:@28030.4]
  assign _T_74714 = $signed(buffer_11_540) + $signed(buffer_4_541); // @[Modules.scala 68:83:@28032.4]
  assign _T_74715 = _T_74714[10:0]; // @[Modules.scala 68:83:@28033.4]
  assign buffer_11_662 = $signed(_T_74715); // @[Modules.scala 68:83:@28034.4]
  assign _T_74717 = $signed(buffer_2_542) + $signed(buffer_11_543); // @[Modules.scala 68:83:@28036.4]
  assign _T_74718 = _T_74717[10:0]; // @[Modules.scala 68:83:@28037.4]
  assign buffer_11_663 = $signed(_T_74718); // @[Modules.scala 68:83:@28038.4]
  assign _T_74720 = $signed(buffer_2_544) + $signed(buffer_0_395); // @[Modules.scala 68:83:@28040.4]
  assign _T_74721 = _T_74720[10:0]; // @[Modules.scala 68:83:@28041.4]
  assign buffer_11_664 = $signed(_T_74721); // @[Modules.scala 68:83:@28042.4]
  assign _T_74723 = $signed(buffer_0_395) + $signed(buffer_11_547); // @[Modules.scala 68:83:@28044.4]
  assign _T_74724 = _T_74723[10:0]; // @[Modules.scala 68:83:@28045.4]
  assign buffer_11_665 = $signed(_T_74724); // @[Modules.scala 68:83:@28046.4]
  assign _T_74726 = $signed(buffer_11_548) + $signed(buffer_1_549); // @[Modules.scala 68:83:@28048.4]
  assign _T_74727 = _T_74726[10:0]; // @[Modules.scala 68:83:@28049.4]
  assign buffer_11_666 = $signed(_T_74727); // @[Modules.scala 68:83:@28050.4]
  assign _T_74732 = $signed(buffer_11_552) + $signed(buffer_7_553); // @[Modules.scala 68:83:@28056.4]
  assign _T_74733 = _T_74732[10:0]; // @[Modules.scala 68:83:@28057.4]
  assign buffer_11_668 = $signed(_T_74733); // @[Modules.scala 68:83:@28058.4]
  assign _T_74735 = $signed(buffer_0_395) + $signed(buffer_11_555); // @[Modules.scala 68:83:@28060.4]
  assign _T_74736 = _T_74735[10:0]; // @[Modules.scala 68:83:@28061.4]
  assign buffer_11_669 = $signed(_T_74736); // @[Modules.scala 68:83:@28062.4]
  assign _T_74738 = $signed(buffer_1_556) + $signed(buffer_2_557); // @[Modules.scala 68:83:@28064.4]
  assign _T_74739 = _T_74738[10:0]; // @[Modules.scala 68:83:@28065.4]
  assign buffer_11_670 = $signed(_T_74739); // @[Modules.scala 68:83:@28066.4]
  assign _T_74741 = $signed(buffer_4_558) + $signed(buffer_2_559); // @[Modules.scala 68:83:@28068.4]
  assign _T_74742 = _T_74741[10:0]; // @[Modules.scala 68:83:@28069.4]
  assign buffer_11_671 = $signed(_T_74742); // @[Modules.scala 68:83:@28070.4]
  assign _T_74750 = $signed(buffer_0_564) + $signed(buffer_11_565); // @[Modules.scala 68:83:@28080.4]
  assign _T_74751 = _T_74750[10:0]; // @[Modules.scala 68:83:@28081.4]
  assign buffer_11_674 = $signed(_T_74751); // @[Modules.scala 68:83:@28082.4]
  assign _T_74753 = $signed(buffer_0_395) + $signed(buffer_11_567); // @[Modules.scala 68:83:@28084.4]
  assign _T_74754 = _T_74753[10:0]; // @[Modules.scala 68:83:@28085.4]
  assign buffer_11_675 = $signed(_T_74754); // @[Modules.scala 68:83:@28086.4]
  assign _T_74762 = $signed(buffer_11_572) + $signed(buffer_0_573); // @[Modules.scala 68:83:@28096.4]
  assign _T_74763 = _T_74762[10:0]; // @[Modules.scala 68:83:@28097.4]
  assign buffer_11_678 = $signed(_T_74763); // @[Modules.scala 68:83:@28098.4]
  assign _T_74774 = $signed(buffer_9_580) + $signed(buffer_11_581); // @[Modules.scala 68:83:@28112.4]
  assign _T_74775 = _T_74774[10:0]; // @[Modules.scala 68:83:@28113.4]
  assign buffer_11_682 = $signed(_T_74775); // @[Modules.scala 68:83:@28114.4]
  assign _T_74786 = $signed(buffer_11_588) + $signed(buffer_11_589); // @[Modules.scala 71:109:@28128.4]
  assign _T_74787 = _T_74786[10:0]; // @[Modules.scala 71:109:@28129.4]
  assign buffer_11_686 = $signed(_T_74787); // @[Modules.scala 71:109:@28130.4]
  assign _T_74789 = $signed(buffer_11_590) + $signed(buffer_11_591); // @[Modules.scala 71:109:@28132.4]
  assign _T_74790 = _T_74789[10:0]; // @[Modules.scala 71:109:@28133.4]
  assign buffer_11_687 = $signed(_T_74790); // @[Modules.scala 71:109:@28134.4]
  assign _T_74792 = $signed(buffer_11_592) + $signed(buffer_11_593); // @[Modules.scala 71:109:@28136.4]
  assign _T_74793 = _T_74792[10:0]; // @[Modules.scala 71:109:@28137.4]
  assign buffer_11_688 = $signed(_T_74793); // @[Modules.scala 71:109:@28138.4]
  assign _T_74795 = $signed(buffer_11_594) + $signed(buffer_11_595); // @[Modules.scala 71:109:@28140.4]
  assign _T_74796 = _T_74795[10:0]; // @[Modules.scala 71:109:@28141.4]
  assign buffer_11_689 = $signed(_T_74796); // @[Modules.scala 71:109:@28142.4]
  assign _T_74798 = $signed(buffer_11_596) + $signed(buffer_0_593); // @[Modules.scala 71:109:@28144.4]
  assign _T_74799 = _T_74798[10:0]; // @[Modules.scala 71:109:@28145.4]
  assign buffer_11_690 = $signed(_T_74799); // @[Modules.scala 71:109:@28146.4]
  assign _T_74801 = $signed(buffer_11_598) + $signed(buffer_11_599); // @[Modules.scala 71:109:@28148.4]
  assign _T_74802 = _T_74801[10:0]; // @[Modules.scala 71:109:@28149.4]
  assign buffer_11_691 = $signed(_T_74802); // @[Modules.scala 71:109:@28150.4]
  assign _T_74807 = $signed(buffer_6_602) + $signed(buffer_11_603); // @[Modules.scala 71:109:@28156.4]
  assign _T_74808 = _T_74807[10:0]; // @[Modules.scala 71:109:@28157.4]
  assign buffer_11_693 = $signed(_T_74808); // @[Modules.scala 71:109:@28158.4]
  assign _T_74810 = $signed(buffer_11_604) + $signed(buffer_11_605); // @[Modules.scala 71:109:@28160.4]
  assign _T_74811 = _T_74810[10:0]; // @[Modules.scala 71:109:@28161.4]
  assign buffer_11_694 = $signed(_T_74811); // @[Modules.scala 71:109:@28162.4]
  assign _T_74813 = $signed(buffer_0_593) + $signed(buffer_11_607); // @[Modules.scala 71:109:@28164.4]
  assign _T_74814 = _T_74813[10:0]; // @[Modules.scala 71:109:@28165.4]
  assign buffer_11_695 = $signed(_T_74814); // @[Modules.scala 71:109:@28166.4]
  assign _T_74816 = $signed(buffer_11_608) + $signed(buffer_11_609); // @[Modules.scala 71:109:@28168.4]
  assign _T_74817 = _T_74816[10:0]; // @[Modules.scala 71:109:@28169.4]
  assign buffer_11_696 = $signed(_T_74817); // @[Modules.scala 71:109:@28170.4]
  assign _T_74819 = $signed(buffer_11_610) + $signed(buffer_11_611); // @[Modules.scala 71:109:@28172.4]
  assign _T_74820 = _T_74819[10:0]; // @[Modules.scala 71:109:@28173.4]
  assign buffer_11_697 = $signed(_T_74820); // @[Modules.scala 71:109:@28174.4]
  assign _T_74822 = $signed(buffer_11_612) + $signed(buffer_11_613); // @[Modules.scala 71:109:@28176.4]
  assign _T_74823 = _T_74822[10:0]; // @[Modules.scala 71:109:@28177.4]
  assign buffer_11_698 = $signed(_T_74823); // @[Modules.scala 71:109:@28178.4]
  assign _T_74825 = $signed(buffer_11_614) + $signed(buffer_7_615); // @[Modules.scala 71:109:@28180.4]
  assign _T_74826 = _T_74825[10:0]; // @[Modules.scala 71:109:@28181.4]
  assign buffer_11_699 = $signed(_T_74826); // @[Modules.scala 71:109:@28182.4]
  assign _T_74828 = $signed(buffer_11_616) + $signed(buffer_11_617); // @[Modules.scala 71:109:@28184.4]
  assign _T_74829 = _T_74828[10:0]; // @[Modules.scala 71:109:@28185.4]
  assign buffer_11_700 = $signed(_T_74829); // @[Modules.scala 71:109:@28186.4]
  assign _T_74831 = $signed(buffer_11_618) + $signed(buffer_11_619); // @[Modules.scala 71:109:@28188.4]
  assign _T_74832 = _T_74831[10:0]; // @[Modules.scala 71:109:@28189.4]
  assign buffer_11_701 = $signed(_T_74832); // @[Modules.scala 71:109:@28190.4]
  assign _T_74834 = $signed(buffer_11_620) + $signed(buffer_11_621); // @[Modules.scala 71:109:@28192.4]
  assign _T_74835 = _T_74834[10:0]; // @[Modules.scala 71:109:@28193.4]
  assign buffer_11_702 = $signed(_T_74835); // @[Modules.scala 71:109:@28194.4]
  assign _T_74837 = $signed(buffer_7_622) + $signed(buffer_11_623); // @[Modules.scala 71:109:@28196.4]
  assign _T_74838 = _T_74837[10:0]; // @[Modules.scala 71:109:@28197.4]
  assign buffer_11_703 = $signed(_T_74838); // @[Modules.scala 71:109:@28198.4]
  assign _T_74840 = $signed(buffer_11_624) + $signed(buffer_9_625); // @[Modules.scala 71:109:@28200.4]
  assign _T_74841 = _T_74840[10:0]; // @[Modules.scala 71:109:@28201.4]
  assign buffer_11_704 = $signed(_T_74841); // @[Modules.scala 71:109:@28202.4]
  assign _T_74843 = $signed(buffer_1_626) + $signed(buffer_11_627); // @[Modules.scala 71:109:@28204.4]
  assign _T_74844 = _T_74843[10:0]; // @[Modules.scala 71:109:@28205.4]
  assign buffer_11_705 = $signed(_T_74844); // @[Modules.scala 71:109:@28206.4]
  assign _T_74846 = $signed(buffer_11_628) + $signed(buffer_1_629); // @[Modules.scala 71:109:@28208.4]
  assign _T_74847 = _T_74846[10:0]; // @[Modules.scala 71:109:@28209.4]
  assign buffer_11_706 = $signed(_T_74847); // @[Modules.scala 71:109:@28210.4]
  assign _T_74852 = $signed(buffer_11_632) + $signed(buffer_11_633); // @[Modules.scala 71:109:@28216.4]
  assign _T_74853 = _T_74852[10:0]; // @[Modules.scala 71:109:@28217.4]
  assign buffer_11_708 = $signed(_T_74853); // @[Modules.scala 71:109:@28218.4]
  assign _T_74855 = $signed(buffer_11_634) + $signed(buffer_11_635); // @[Modules.scala 71:109:@28220.4]
  assign _T_74856 = _T_74855[10:0]; // @[Modules.scala 71:109:@28221.4]
  assign buffer_11_709 = $signed(_T_74856); // @[Modules.scala 71:109:@28222.4]
  assign _T_74858 = $signed(buffer_11_636) + $signed(buffer_3_637); // @[Modules.scala 71:109:@28224.4]
  assign _T_74859 = _T_74858[10:0]; // @[Modules.scala 71:109:@28225.4]
  assign buffer_11_710 = $signed(_T_74859); // @[Modules.scala 71:109:@28226.4]
  assign _T_74861 = $signed(buffer_11_638) + $signed(buffer_0_593); // @[Modules.scala 71:109:@28228.4]
  assign _T_74862 = _T_74861[10:0]; // @[Modules.scala 71:109:@28229.4]
  assign buffer_11_711 = $signed(_T_74862); // @[Modules.scala 71:109:@28230.4]
  assign _T_74864 = $signed(buffer_11_640) + $signed(buffer_11_641); // @[Modules.scala 71:109:@28232.4]
  assign _T_74865 = _T_74864[10:0]; // @[Modules.scala 71:109:@28233.4]
  assign buffer_11_712 = $signed(_T_74865); // @[Modules.scala 71:109:@28234.4]
  assign _T_74867 = $signed(buffer_11_642) + $signed(buffer_0_593); // @[Modules.scala 71:109:@28236.4]
  assign _T_74868 = _T_74867[10:0]; // @[Modules.scala 71:109:@28237.4]
  assign buffer_11_713 = $signed(_T_74868); // @[Modules.scala 71:109:@28238.4]
  assign _T_74870 = $signed(buffer_11_644) + $signed(buffer_11_645); // @[Modules.scala 71:109:@28240.4]
  assign _T_74871 = _T_74870[10:0]; // @[Modules.scala 71:109:@28241.4]
  assign buffer_11_714 = $signed(_T_74871); // @[Modules.scala 71:109:@28242.4]
  assign _T_74873 = $signed(buffer_11_646) + $signed(buffer_11_647); // @[Modules.scala 71:109:@28244.4]
  assign _T_74874 = _T_74873[10:0]; // @[Modules.scala 71:109:@28245.4]
  assign buffer_11_715 = $signed(_T_74874); // @[Modules.scala 71:109:@28246.4]
  assign _T_74876 = $signed(buffer_11_648) + $signed(buffer_11_649); // @[Modules.scala 71:109:@28248.4]
  assign _T_74877 = _T_74876[10:0]; // @[Modules.scala 71:109:@28249.4]
  assign buffer_11_716 = $signed(_T_74877); // @[Modules.scala 71:109:@28250.4]
  assign _T_74879 = $signed(buffer_11_650) + $signed(buffer_11_651); // @[Modules.scala 71:109:@28252.4]
  assign _T_74880 = _T_74879[10:0]; // @[Modules.scala 71:109:@28253.4]
  assign buffer_11_717 = $signed(_T_74880); // @[Modules.scala 71:109:@28254.4]
  assign _T_74882 = $signed(buffer_11_652) + $signed(buffer_11_653); // @[Modules.scala 71:109:@28256.4]
  assign _T_74883 = _T_74882[10:0]; // @[Modules.scala 71:109:@28257.4]
  assign buffer_11_718 = $signed(_T_74883); // @[Modules.scala 71:109:@28258.4]
  assign _T_74885 = $signed(buffer_0_593) + $signed(buffer_11_655); // @[Modules.scala 71:109:@28260.4]
  assign _T_74886 = _T_74885[10:0]; // @[Modules.scala 71:109:@28261.4]
  assign buffer_11_719 = $signed(_T_74886); // @[Modules.scala 71:109:@28262.4]
  assign _T_74888 = $signed(buffer_11_656) + $signed(buffer_11_657); // @[Modules.scala 71:109:@28264.4]
  assign _T_74889 = _T_74888[10:0]; // @[Modules.scala 71:109:@28265.4]
  assign buffer_11_720 = $signed(_T_74889); // @[Modules.scala 71:109:@28266.4]
  assign _T_74891 = $signed(buffer_11_658) + $signed(buffer_11_659); // @[Modules.scala 71:109:@28268.4]
  assign _T_74892 = _T_74891[10:0]; // @[Modules.scala 71:109:@28269.4]
  assign buffer_11_721 = $signed(_T_74892); // @[Modules.scala 71:109:@28270.4]
  assign _T_74894 = $signed(buffer_11_660) + $signed(buffer_11_661); // @[Modules.scala 71:109:@28272.4]
  assign _T_74895 = _T_74894[10:0]; // @[Modules.scala 71:109:@28273.4]
  assign buffer_11_722 = $signed(_T_74895); // @[Modules.scala 71:109:@28274.4]
  assign _T_74897 = $signed(buffer_11_662) + $signed(buffer_11_663); // @[Modules.scala 71:109:@28276.4]
  assign _T_74898 = _T_74897[10:0]; // @[Modules.scala 71:109:@28277.4]
  assign buffer_11_723 = $signed(_T_74898); // @[Modules.scala 71:109:@28278.4]
  assign _T_74900 = $signed(buffer_11_664) + $signed(buffer_11_665); // @[Modules.scala 71:109:@28280.4]
  assign _T_74901 = _T_74900[10:0]; // @[Modules.scala 71:109:@28281.4]
  assign buffer_11_724 = $signed(_T_74901); // @[Modules.scala 71:109:@28282.4]
  assign _T_74903 = $signed(buffer_11_666) + $signed(buffer_2_667); // @[Modules.scala 71:109:@28284.4]
  assign _T_74904 = _T_74903[10:0]; // @[Modules.scala 71:109:@28285.4]
  assign buffer_11_725 = $signed(_T_74904); // @[Modules.scala 71:109:@28286.4]
  assign _T_74906 = $signed(buffer_11_668) + $signed(buffer_11_669); // @[Modules.scala 71:109:@28288.4]
  assign _T_74907 = _T_74906[10:0]; // @[Modules.scala 71:109:@28289.4]
  assign buffer_11_726 = $signed(_T_74907); // @[Modules.scala 71:109:@28290.4]
  assign _T_74909 = $signed(buffer_11_670) + $signed(buffer_11_671); // @[Modules.scala 71:109:@28292.4]
  assign _T_74910 = _T_74909[10:0]; // @[Modules.scala 71:109:@28293.4]
  assign buffer_11_727 = $signed(_T_74910); // @[Modules.scala 71:109:@28294.4]
  assign _T_74912 = $signed(buffer_0_593) + $signed(buffer_7_673); // @[Modules.scala 71:109:@28296.4]
  assign _T_74913 = _T_74912[10:0]; // @[Modules.scala 71:109:@28297.4]
  assign buffer_11_728 = $signed(_T_74913); // @[Modules.scala 71:109:@28298.4]
  assign _T_74915 = $signed(buffer_11_674) + $signed(buffer_11_675); // @[Modules.scala 71:109:@28300.4]
  assign _T_74916 = _T_74915[10:0]; // @[Modules.scala 71:109:@28301.4]
  assign buffer_11_729 = $signed(_T_74916); // @[Modules.scala 71:109:@28302.4]
  assign _T_74921 = $signed(buffer_11_678) + $signed(buffer_10_679); // @[Modules.scala 71:109:@28308.4]
  assign _T_74922 = _T_74921[10:0]; // @[Modules.scala 71:109:@28309.4]
  assign buffer_11_731 = $signed(_T_74922); // @[Modules.scala 71:109:@28310.4]
  assign _T_74927 = $signed(buffer_11_682) + $signed(buffer_0_593); // @[Modules.scala 71:109:@28316.4]
  assign _T_74928 = _T_74927[10:0]; // @[Modules.scala 71:109:@28317.4]
  assign buffer_11_733 = $signed(_T_74928); // @[Modules.scala 71:109:@28318.4]
  assign _T_74933 = $signed(buffer_11_686) + $signed(buffer_11_687); // @[Modules.scala 78:156:@28325.4]
  assign _T_74934 = _T_74933[10:0]; // @[Modules.scala 78:156:@28326.4]
  assign buffer_11_736 = $signed(_T_74934); // @[Modules.scala 78:156:@28327.4]
  assign _T_74936 = $signed(buffer_11_736) + $signed(buffer_11_688); // @[Modules.scala 78:156:@28329.4]
  assign _T_74937 = _T_74936[10:0]; // @[Modules.scala 78:156:@28330.4]
  assign buffer_11_737 = $signed(_T_74937); // @[Modules.scala 78:156:@28331.4]
  assign _T_74939 = $signed(buffer_11_737) + $signed(buffer_11_689); // @[Modules.scala 78:156:@28333.4]
  assign _T_74940 = _T_74939[10:0]; // @[Modules.scala 78:156:@28334.4]
  assign buffer_11_738 = $signed(_T_74940); // @[Modules.scala 78:156:@28335.4]
  assign _T_74942 = $signed(buffer_11_738) + $signed(buffer_11_690); // @[Modules.scala 78:156:@28337.4]
  assign _T_74943 = _T_74942[10:0]; // @[Modules.scala 78:156:@28338.4]
  assign buffer_11_739 = $signed(_T_74943); // @[Modules.scala 78:156:@28339.4]
  assign _T_74945 = $signed(buffer_11_739) + $signed(buffer_11_691); // @[Modules.scala 78:156:@28341.4]
  assign _T_74946 = _T_74945[10:0]; // @[Modules.scala 78:156:@28342.4]
  assign buffer_11_740 = $signed(_T_74946); // @[Modules.scala 78:156:@28343.4]
  assign _T_74948 = $signed(buffer_11_740) + $signed(buffer_8_692); // @[Modules.scala 78:156:@28345.4]
  assign _T_74949 = _T_74948[10:0]; // @[Modules.scala 78:156:@28346.4]
  assign buffer_11_741 = $signed(_T_74949); // @[Modules.scala 78:156:@28347.4]
  assign _T_74951 = $signed(buffer_11_741) + $signed(buffer_11_693); // @[Modules.scala 78:156:@28349.4]
  assign _T_74952 = _T_74951[10:0]; // @[Modules.scala 78:156:@28350.4]
  assign buffer_11_742 = $signed(_T_74952); // @[Modules.scala 78:156:@28351.4]
  assign _T_74954 = $signed(buffer_11_742) + $signed(buffer_11_694); // @[Modules.scala 78:156:@28353.4]
  assign _T_74955 = _T_74954[10:0]; // @[Modules.scala 78:156:@28354.4]
  assign buffer_11_743 = $signed(_T_74955); // @[Modules.scala 78:156:@28355.4]
  assign _T_74957 = $signed(buffer_11_743) + $signed(buffer_11_695); // @[Modules.scala 78:156:@28357.4]
  assign _T_74958 = _T_74957[10:0]; // @[Modules.scala 78:156:@28358.4]
  assign buffer_11_744 = $signed(_T_74958); // @[Modules.scala 78:156:@28359.4]
  assign _T_74960 = $signed(buffer_11_744) + $signed(buffer_11_696); // @[Modules.scala 78:156:@28361.4]
  assign _T_74961 = _T_74960[10:0]; // @[Modules.scala 78:156:@28362.4]
  assign buffer_11_745 = $signed(_T_74961); // @[Modules.scala 78:156:@28363.4]
  assign _T_74963 = $signed(buffer_11_745) + $signed(buffer_11_697); // @[Modules.scala 78:156:@28365.4]
  assign _T_74964 = _T_74963[10:0]; // @[Modules.scala 78:156:@28366.4]
  assign buffer_11_746 = $signed(_T_74964); // @[Modules.scala 78:156:@28367.4]
  assign _T_74966 = $signed(buffer_11_746) + $signed(buffer_11_698); // @[Modules.scala 78:156:@28369.4]
  assign _T_74967 = _T_74966[10:0]; // @[Modules.scala 78:156:@28370.4]
  assign buffer_11_747 = $signed(_T_74967); // @[Modules.scala 78:156:@28371.4]
  assign _T_74969 = $signed(buffer_11_747) + $signed(buffer_11_699); // @[Modules.scala 78:156:@28373.4]
  assign _T_74970 = _T_74969[10:0]; // @[Modules.scala 78:156:@28374.4]
  assign buffer_11_748 = $signed(_T_74970); // @[Modules.scala 78:156:@28375.4]
  assign _T_74972 = $signed(buffer_11_748) + $signed(buffer_11_700); // @[Modules.scala 78:156:@28377.4]
  assign _T_74973 = _T_74972[10:0]; // @[Modules.scala 78:156:@28378.4]
  assign buffer_11_749 = $signed(_T_74973); // @[Modules.scala 78:156:@28379.4]
  assign _T_74975 = $signed(buffer_11_749) + $signed(buffer_11_701); // @[Modules.scala 78:156:@28381.4]
  assign _T_74976 = _T_74975[10:0]; // @[Modules.scala 78:156:@28382.4]
  assign buffer_11_750 = $signed(_T_74976); // @[Modules.scala 78:156:@28383.4]
  assign _T_74978 = $signed(buffer_11_750) + $signed(buffer_11_702); // @[Modules.scala 78:156:@28385.4]
  assign _T_74979 = _T_74978[10:0]; // @[Modules.scala 78:156:@28386.4]
  assign buffer_11_751 = $signed(_T_74979); // @[Modules.scala 78:156:@28387.4]
  assign _T_74981 = $signed(buffer_11_751) + $signed(buffer_11_703); // @[Modules.scala 78:156:@28389.4]
  assign _T_74982 = _T_74981[10:0]; // @[Modules.scala 78:156:@28390.4]
  assign buffer_11_752 = $signed(_T_74982); // @[Modules.scala 78:156:@28391.4]
  assign _T_74984 = $signed(buffer_11_752) + $signed(buffer_11_704); // @[Modules.scala 78:156:@28393.4]
  assign _T_74985 = _T_74984[10:0]; // @[Modules.scala 78:156:@28394.4]
  assign buffer_11_753 = $signed(_T_74985); // @[Modules.scala 78:156:@28395.4]
  assign _T_74987 = $signed(buffer_11_753) + $signed(buffer_11_705); // @[Modules.scala 78:156:@28397.4]
  assign _T_74988 = _T_74987[10:0]; // @[Modules.scala 78:156:@28398.4]
  assign buffer_11_754 = $signed(_T_74988); // @[Modules.scala 78:156:@28399.4]
  assign _T_74990 = $signed(buffer_11_754) + $signed(buffer_11_706); // @[Modules.scala 78:156:@28401.4]
  assign _T_74991 = _T_74990[10:0]; // @[Modules.scala 78:156:@28402.4]
  assign buffer_11_755 = $signed(_T_74991); // @[Modules.scala 78:156:@28403.4]
  assign _T_74993 = $signed(buffer_11_755) + $signed(buffer_0_707); // @[Modules.scala 78:156:@28405.4]
  assign _T_74994 = _T_74993[10:0]; // @[Modules.scala 78:156:@28406.4]
  assign buffer_11_756 = $signed(_T_74994); // @[Modules.scala 78:156:@28407.4]
  assign _T_74996 = $signed(buffer_11_756) + $signed(buffer_11_708); // @[Modules.scala 78:156:@28409.4]
  assign _T_74997 = _T_74996[10:0]; // @[Modules.scala 78:156:@28410.4]
  assign buffer_11_757 = $signed(_T_74997); // @[Modules.scala 78:156:@28411.4]
  assign _T_74999 = $signed(buffer_11_757) + $signed(buffer_11_709); // @[Modules.scala 78:156:@28413.4]
  assign _T_75000 = _T_74999[10:0]; // @[Modules.scala 78:156:@28414.4]
  assign buffer_11_758 = $signed(_T_75000); // @[Modules.scala 78:156:@28415.4]
  assign _T_75002 = $signed(buffer_11_758) + $signed(buffer_11_710); // @[Modules.scala 78:156:@28417.4]
  assign _T_75003 = _T_75002[10:0]; // @[Modules.scala 78:156:@28418.4]
  assign buffer_11_759 = $signed(_T_75003); // @[Modules.scala 78:156:@28419.4]
  assign _T_75005 = $signed(buffer_11_759) + $signed(buffer_11_711); // @[Modules.scala 78:156:@28421.4]
  assign _T_75006 = _T_75005[10:0]; // @[Modules.scala 78:156:@28422.4]
  assign buffer_11_760 = $signed(_T_75006); // @[Modules.scala 78:156:@28423.4]
  assign _T_75008 = $signed(buffer_11_760) + $signed(buffer_11_712); // @[Modules.scala 78:156:@28425.4]
  assign _T_75009 = _T_75008[10:0]; // @[Modules.scala 78:156:@28426.4]
  assign buffer_11_761 = $signed(_T_75009); // @[Modules.scala 78:156:@28427.4]
  assign _T_75011 = $signed(buffer_11_761) + $signed(buffer_11_713); // @[Modules.scala 78:156:@28429.4]
  assign _T_75012 = _T_75011[10:0]; // @[Modules.scala 78:156:@28430.4]
  assign buffer_11_762 = $signed(_T_75012); // @[Modules.scala 78:156:@28431.4]
  assign _T_75014 = $signed(buffer_11_762) + $signed(buffer_11_714); // @[Modules.scala 78:156:@28433.4]
  assign _T_75015 = _T_75014[10:0]; // @[Modules.scala 78:156:@28434.4]
  assign buffer_11_763 = $signed(_T_75015); // @[Modules.scala 78:156:@28435.4]
  assign _T_75017 = $signed(buffer_11_763) + $signed(buffer_11_715); // @[Modules.scala 78:156:@28437.4]
  assign _T_75018 = _T_75017[10:0]; // @[Modules.scala 78:156:@28438.4]
  assign buffer_11_764 = $signed(_T_75018); // @[Modules.scala 78:156:@28439.4]
  assign _T_75020 = $signed(buffer_11_764) + $signed(buffer_11_716); // @[Modules.scala 78:156:@28441.4]
  assign _T_75021 = _T_75020[10:0]; // @[Modules.scala 78:156:@28442.4]
  assign buffer_11_765 = $signed(_T_75021); // @[Modules.scala 78:156:@28443.4]
  assign _T_75023 = $signed(buffer_11_765) + $signed(buffer_11_717); // @[Modules.scala 78:156:@28445.4]
  assign _T_75024 = _T_75023[10:0]; // @[Modules.scala 78:156:@28446.4]
  assign buffer_11_766 = $signed(_T_75024); // @[Modules.scala 78:156:@28447.4]
  assign _T_75026 = $signed(buffer_11_766) + $signed(buffer_11_718); // @[Modules.scala 78:156:@28449.4]
  assign _T_75027 = _T_75026[10:0]; // @[Modules.scala 78:156:@28450.4]
  assign buffer_11_767 = $signed(_T_75027); // @[Modules.scala 78:156:@28451.4]
  assign _T_75029 = $signed(buffer_11_767) + $signed(buffer_11_719); // @[Modules.scala 78:156:@28453.4]
  assign _T_75030 = _T_75029[10:0]; // @[Modules.scala 78:156:@28454.4]
  assign buffer_11_768 = $signed(_T_75030); // @[Modules.scala 78:156:@28455.4]
  assign _T_75032 = $signed(buffer_11_768) + $signed(buffer_11_720); // @[Modules.scala 78:156:@28457.4]
  assign _T_75033 = _T_75032[10:0]; // @[Modules.scala 78:156:@28458.4]
  assign buffer_11_769 = $signed(_T_75033); // @[Modules.scala 78:156:@28459.4]
  assign _T_75035 = $signed(buffer_11_769) + $signed(buffer_11_721); // @[Modules.scala 78:156:@28461.4]
  assign _T_75036 = _T_75035[10:0]; // @[Modules.scala 78:156:@28462.4]
  assign buffer_11_770 = $signed(_T_75036); // @[Modules.scala 78:156:@28463.4]
  assign _T_75038 = $signed(buffer_11_770) + $signed(buffer_11_722); // @[Modules.scala 78:156:@28465.4]
  assign _T_75039 = _T_75038[10:0]; // @[Modules.scala 78:156:@28466.4]
  assign buffer_11_771 = $signed(_T_75039); // @[Modules.scala 78:156:@28467.4]
  assign _T_75041 = $signed(buffer_11_771) + $signed(buffer_11_723); // @[Modules.scala 78:156:@28469.4]
  assign _T_75042 = _T_75041[10:0]; // @[Modules.scala 78:156:@28470.4]
  assign buffer_11_772 = $signed(_T_75042); // @[Modules.scala 78:156:@28471.4]
  assign _T_75044 = $signed(buffer_11_772) + $signed(buffer_11_724); // @[Modules.scala 78:156:@28473.4]
  assign _T_75045 = _T_75044[10:0]; // @[Modules.scala 78:156:@28474.4]
  assign buffer_11_773 = $signed(_T_75045); // @[Modules.scala 78:156:@28475.4]
  assign _T_75047 = $signed(buffer_11_773) + $signed(buffer_11_725); // @[Modules.scala 78:156:@28477.4]
  assign _T_75048 = _T_75047[10:0]; // @[Modules.scala 78:156:@28478.4]
  assign buffer_11_774 = $signed(_T_75048); // @[Modules.scala 78:156:@28479.4]
  assign _T_75050 = $signed(buffer_11_774) + $signed(buffer_11_726); // @[Modules.scala 78:156:@28481.4]
  assign _T_75051 = _T_75050[10:0]; // @[Modules.scala 78:156:@28482.4]
  assign buffer_11_775 = $signed(_T_75051); // @[Modules.scala 78:156:@28483.4]
  assign _T_75053 = $signed(buffer_11_775) + $signed(buffer_11_727); // @[Modules.scala 78:156:@28485.4]
  assign _T_75054 = _T_75053[10:0]; // @[Modules.scala 78:156:@28486.4]
  assign buffer_11_776 = $signed(_T_75054); // @[Modules.scala 78:156:@28487.4]
  assign _T_75056 = $signed(buffer_11_776) + $signed(buffer_11_728); // @[Modules.scala 78:156:@28489.4]
  assign _T_75057 = _T_75056[10:0]; // @[Modules.scala 78:156:@28490.4]
  assign buffer_11_777 = $signed(_T_75057); // @[Modules.scala 78:156:@28491.4]
  assign _T_75059 = $signed(buffer_11_777) + $signed(buffer_11_729); // @[Modules.scala 78:156:@28493.4]
  assign _T_75060 = _T_75059[10:0]; // @[Modules.scala 78:156:@28494.4]
  assign buffer_11_778 = $signed(_T_75060); // @[Modules.scala 78:156:@28495.4]
  assign _T_75062 = $signed(buffer_11_778) + $signed(buffer_0_701); // @[Modules.scala 78:156:@28497.4]
  assign _T_75063 = _T_75062[10:0]; // @[Modules.scala 78:156:@28498.4]
  assign buffer_11_779 = $signed(_T_75063); // @[Modules.scala 78:156:@28499.4]
  assign _T_75065 = $signed(buffer_11_779) + $signed(buffer_11_731); // @[Modules.scala 78:156:@28501.4]
  assign _T_75066 = _T_75065[10:0]; // @[Modules.scala 78:156:@28502.4]
  assign buffer_11_780 = $signed(_T_75066); // @[Modules.scala 78:156:@28503.4]
  assign _T_75068 = $signed(buffer_11_780) + $signed(buffer_0_701); // @[Modules.scala 78:156:@28505.4]
  assign _T_75069 = _T_75068[10:0]; // @[Modules.scala 78:156:@28506.4]
  assign buffer_11_781 = $signed(_T_75069); // @[Modules.scala 78:156:@28507.4]
  assign _T_75071 = $signed(buffer_11_781) + $signed(buffer_11_733); // @[Modules.scala 78:156:@28509.4]
  assign _T_75072 = _T_75071[10:0]; // @[Modules.scala 78:156:@28510.4]
  assign buffer_11_782 = $signed(_T_75072); // @[Modules.scala 78:156:@28511.4]
  assign _T_75074 = $signed(buffer_11_782) + $signed(buffer_2_734); // @[Modules.scala 78:156:@28513.4]
  assign _T_75075 = _T_75074[10:0]; // @[Modules.scala 78:156:@28514.4]
  assign buffer_11_783 = $signed(_T_75075); // @[Modules.scala 78:156:@28515.4]
  assign _T_75490 = $signed(io_in_560) + $signed(io_in_561); // @[Modules.scala 37:46:@29119.4]
  assign _T_75491 = _T_75490[4:0]; // @[Modules.scala 37:46:@29120.4]
  assign _T_75492 = $signed(_T_75491); // @[Modules.scala 37:46:@29121.4]
  assign _T_75665 = $signed(buffer_7_0) + $signed(buffer_4_1); // @[Modules.scala 65:57:@29366.4]
  assign _T_75666 = _T_75665[10:0]; // @[Modules.scala 65:57:@29367.4]
  assign buffer_12_392 = $signed(_T_75666); // @[Modules.scala 65:57:@29368.4]
  assign buffer_12_7 = {{6{io_in_14[4]}},io_in_14}; // @[Modules.scala 32:22:@8.4]
  assign _T_75674 = $signed(buffer_1_6) + $signed(buffer_12_7); // @[Modules.scala 65:57:@29378.4]
  assign _T_75675 = _T_75674[10:0]; // @[Modules.scala 65:57:@29379.4]
  assign buffer_12_395 = $signed(_T_75675); // @[Modules.scala 65:57:@29380.4]
  assign _T_75677 = $signed(buffer_7_8) + $signed(buffer_1_9); // @[Modules.scala 65:57:@29382.4]
  assign _T_75678 = _T_75677[10:0]; // @[Modules.scala 65:57:@29383.4]
  assign buffer_12_396 = $signed(_T_75678); // @[Modules.scala 65:57:@29384.4]
  assign _T_75680 = $signed(11'sh0) + $signed(buffer_1_11); // @[Modules.scala 65:57:@29386.4]
  assign _T_75681 = _T_75680[10:0]; // @[Modules.scala 65:57:@29387.4]
  assign buffer_12_397 = $signed(_T_75681); // @[Modules.scala 65:57:@29388.4]
  assign _T_75683 = $signed(buffer_0_12) + $signed(11'sh0); // @[Modules.scala 65:57:@29390.4]
  assign _T_75684 = _T_75683[10:0]; // @[Modules.scala 65:57:@29391.4]
  assign buffer_12_398 = $signed(_T_75684); // @[Modules.scala 65:57:@29392.4]
  assign _T_75686 = $signed(buffer_1_14) + $signed(buffer_2_15); // @[Modules.scala 65:57:@29394.4]
  assign _T_75687 = _T_75686[10:0]; // @[Modules.scala 65:57:@29395.4]
  assign buffer_12_399 = $signed(_T_75687); // @[Modules.scala 65:57:@29396.4]
  assign _T_75746 = $signed(buffer_1_54) + $signed(buffer_3_55); // @[Modules.scala 65:57:@29474.4]
  assign _T_75747 = _T_75746[10:0]; // @[Modules.scala 65:57:@29475.4]
  assign buffer_12_419 = $signed(_T_75747); // @[Modules.scala 65:57:@29476.4]
  assign _T_75752 = $signed(11'sh0) + $signed(buffer_4_59); // @[Modules.scala 65:57:@29482.4]
  assign _T_75753 = _T_75752[10:0]; // @[Modules.scala 65:57:@29483.4]
  assign buffer_12_421 = $signed(_T_75753); // @[Modules.scala 65:57:@29484.4]
  assign _T_75758 = $signed(buffer_8_62) + $signed(11'sh0); // @[Modules.scala 65:57:@29490.4]
  assign _T_75759 = _T_75758[10:0]; // @[Modules.scala 65:57:@29491.4]
  assign buffer_12_423 = $signed(_T_75759); // @[Modules.scala 65:57:@29492.4]
  assign _T_75764 = $signed(buffer_5_66) + $signed(buffer_3_67); // @[Modules.scala 65:57:@29498.4]
  assign _T_75765 = _T_75764[10:0]; // @[Modules.scala 65:57:@29499.4]
  assign buffer_12_425 = $signed(_T_75765); // @[Modules.scala 65:57:@29500.4]
  assign _T_75767 = $signed(11'sh0) + $signed(buffer_1_69); // @[Modules.scala 65:57:@29502.4]
  assign _T_75768 = _T_75767[10:0]; // @[Modules.scala 65:57:@29503.4]
  assign buffer_12_426 = $signed(_T_75768); // @[Modules.scala 65:57:@29504.4]
  assign _T_75773 = $signed(buffer_0_72) + $signed(11'sh0); // @[Modules.scala 65:57:@29510.4]
  assign _T_75774 = _T_75773[10:0]; // @[Modules.scala 65:57:@29511.4]
  assign buffer_12_428 = $signed(_T_75774); // @[Modules.scala 65:57:@29512.4]
  assign _T_75776 = $signed(buffer_0_74) + $signed(buffer_1_75); // @[Modules.scala 65:57:@29514.4]
  assign _T_75777 = _T_75776[10:0]; // @[Modules.scala 65:57:@29515.4]
  assign buffer_12_429 = $signed(_T_75777); // @[Modules.scala 65:57:@29516.4]
  assign _T_75782 = $signed(buffer_9_78) + $signed(buffer_3_79); // @[Modules.scala 65:57:@29522.4]
  assign _T_75783 = _T_75782[10:0]; // @[Modules.scala 65:57:@29523.4]
  assign buffer_12_431 = $signed(_T_75783); // @[Modules.scala 65:57:@29524.4]
  assign _T_75788 = $signed(11'sh0) + $signed(buffer_0_83); // @[Modules.scala 65:57:@29530.4]
  assign _T_75789 = _T_75788[10:0]; // @[Modules.scala 65:57:@29531.4]
  assign buffer_12_433 = $signed(_T_75789); // @[Modules.scala 65:57:@29532.4]
  assign _T_75803 = $signed(buffer_4_92) + $signed(buffer_3_93); // @[Modules.scala 65:57:@29550.4]
  assign _T_75804 = _T_75803[10:0]; // @[Modules.scala 65:57:@29551.4]
  assign buffer_12_438 = $signed(_T_75804); // @[Modules.scala 65:57:@29552.4]
  assign _T_75815 = $signed(11'sh0) + $signed(buffer_5_101); // @[Modules.scala 65:57:@29566.4]
  assign _T_75816 = _T_75815[10:0]; // @[Modules.scala 65:57:@29567.4]
  assign buffer_12_442 = $signed(_T_75816); // @[Modules.scala 65:57:@29568.4]
  assign _T_75818 = $signed(buffer_1_102) + $signed(buffer_0_103); // @[Modules.scala 65:57:@29570.4]
  assign _T_75819 = _T_75818[10:0]; // @[Modules.scala 65:57:@29571.4]
  assign buffer_12_443 = $signed(_T_75819); // @[Modules.scala 65:57:@29572.4]
  assign _T_75824 = $signed(buffer_1_106) + $signed(buffer_2_107); // @[Modules.scala 65:57:@29578.4]
  assign _T_75825 = _T_75824[10:0]; // @[Modules.scala 65:57:@29579.4]
  assign buffer_12_445 = $signed(_T_75825); // @[Modules.scala 65:57:@29580.4]
  assign buffer_12_113 = {{6{io_in_226[4]}},io_in_226}; // @[Modules.scala 32:22:@8.4]
  assign _T_75833 = $signed(buffer_1_112) + $signed(buffer_12_113); // @[Modules.scala 65:57:@29590.4]
  assign _T_75834 = _T_75833[10:0]; // @[Modules.scala 65:57:@29591.4]
  assign buffer_12_448 = $signed(_T_75834); // @[Modules.scala 65:57:@29592.4]
  assign _T_75839 = $signed(buffer_7_116) + $signed(buffer_3_117); // @[Modules.scala 65:57:@29598.4]
  assign _T_75840 = _T_75839[10:0]; // @[Modules.scala 65:57:@29599.4]
  assign buffer_12_450 = $signed(_T_75840); // @[Modules.scala 65:57:@29600.4]
  assign _T_75842 = $signed(11'sh0) + $signed(buffer_3_119); // @[Modules.scala 65:57:@29602.4]
  assign _T_75843 = _T_75842[10:0]; // @[Modules.scala 65:57:@29603.4]
  assign buffer_12_451 = $signed(_T_75843); // @[Modules.scala 65:57:@29604.4]
  assign _T_75854 = $signed(buffer_3_126) + $signed(buffer_8_127); // @[Modules.scala 65:57:@29618.4]
  assign _T_75855 = _T_75854[10:0]; // @[Modules.scala 65:57:@29619.4]
  assign buffer_12_455 = $signed(_T_75855); // @[Modules.scala 65:57:@29620.4]
  assign _T_75857 = $signed(buffer_4_128) + $signed(11'sh0); // @[Modules.scala 65:57:@29622.4]
  assign _T_75858 = _T_75857[10:0]; // @[Modules.scala 65:57:@29623.4]
  assign buffer_12_456 = $signed(_T_75858); // @[Modules.scala 65:57:@29624.4]
  assign _T_75860 = $signed(buffer_1_130) + $signed(buffer_0_131); // @[Modules.scala 65:57:@29626.4]
  assign _T_75861 = _T_75860[10:0]; // @[Modules.scala 65:57:@29627.4]
  assign buffer_12_457 = $signed(_T_75861); // @[Modules.scala 65:57:@29628.4]
  assign _T_75863 = $signed(buffer_3_132) + $signed(buffer_9_133); // @[Modules.scala 65:57:@29630.4]
  assign _T_75864 = _T_75863[10:0]; // @[Modules.scala 65:57:@29631.4]
  assign buffer_12_458 = $signed(_T_75864); // @[Modules.scala 65:57:@29632.4]
  assign _T_75866 = $signed(buffer_3_134) + $signed(buffer_11_135); // @[Modules.scala 65:57:@29634.4]
  assign _T_75867 = _T_75866[10:0]; // @[Modules.scala 65:57:@29635.4]
  assign buffer_12_459 = $signed(_T_75867); // @[Modules.scala 65:57:@29636.4]
  assign _T_75875 = $signed(buffer_3_140) + $signed(buffer_8_141); // @[Modules.scala 65:57:@29646.4]
  assign _T_75876 = _T_75875[10:0]; // @[Modules.scala 65:57:@29647.4]
  assign buffer_12_462 = $signed(_T_75876); // @[Modules.scala 65:57:@29648.4]
  assign _T_75887 = $signed(11'sh0) + $signed(buffer_3_149); // @[Modules.scala 65:57:@29662.4]
  assign _T_75888 = _T_75887[10:0]; // @[Modules.scala 65:57:@29663.4]
  assign buffer_12_466 = $signed(_T_75888); // @[Modules.scala 65:57:@29664.4]
  assign _T_75890 = $signed(buffer_6_150) + $signed(buffer_5_151); // @[Modules.scala 65:57:@29666.4]
  assign _T_75891 = _T_75890[10:0]; // @[Modules.scala 65:57:@29667.4]
  assign buffer_12_467 = $signed(_T_75891); // @[Modules.scala 65:57:@29668.4]
  assign buffer_12_155 = {{6{io_in_310[4]}},io_in_310}; // @[Modules.scala 32:22:@8.4]
  assign _T_75896 = $signed(buffer_10_154) + $signed(buffer_12_155); // @[Modules.scala 65:57:@29674.4]
  assign _T_75897 = _T_75896[10:0]; // @[Modules.scala 65:57:@29675.4]
  assign buffer_12_469 = $signed(_T_75897); // @[Modules.scala 65:57:@29676.4]
  assign buffer_12_163 = {{6{io_in_327[4]}},io_in_327}; // @[Modules.scala 32:22:@8.4]
  assign _T_75908 = $signed(11'sh0) + $signed(buffer_12_163); // @[Modules.scala 65:57:@29690.4]
  assign _T_75909 = _T_75908[10:0]; // @[Modules.scala 65:57:@29691.4]
  assign buffer_12_473 = $signed(_T_75909); // @[Modules.scala 65:57:@29692.4]
  assign buffer_12_164 = {{6{io_in_329[4]}},io_in_329}; // @[Modules.scala 32:22:@8.4]
  assign _T_75911 = $signed(buffer_12_164) + $signed(buffer_5_165); // @[Modules.scala 65:57:@29694.4]
  assign _T_75912 = _T_75911[10:0]; // @[Modules.scala 65:57:@29695.4]
  assign buffer_12_474 = $signed(_T_75912); // @[Modules.scala 65:57:@29696.4]
  assign buffer_12_166 = {{6{io_in_332[4]}},io_in_332}; // @[Modules.scala 32:22:@8.4]
  assign _T_75914 = $signed(buffer_12_166) + $signed(11'sh0); // @[Modules.scala 65:57:@29698.4]
  assign _T_75915 = _T_75914[10:0]; // @[Modules.scala 65:57:@29699.4]
  assign buffer_12_475 = $signed(_T_75915); // @[Modules.scala 65:57:@29700.4]
  assign _T_75917 = $signed(buffer_5_168) + $signed(buffer_3_169); // @[Modules.scala 65:57:@29702.4]
  assign _T_75918 = _T_75917[10:0]; // @[Modules.scala 65:57:@29703.4]
  assign buffer_12_476 = $signed(_T_75918); // @[Modules.scala 65:57:@29704.4]
  assign _T_75959 = $signed(11'sh0) + $signed(buffer_3_197); // @[Modules.scala 65:57:@29758.4]
  assign _T_75960 = _T_75959[10:0]; // @[Modules.scala 65:57:@29759.4]
  assign buffer_12_490 = $signed(_T_75960); // @[Modules.scala 65:57:@29760.4]
  assign _T_75962 = $signed(11'sh0) + $signed(buffer_4_199); // @[Modules.scala 65:57:@29762.4]
  assign _T_75963 = _T_75962[10:0]; // @[Modules.scala 65:57:@29763.4]
  assign buffer_12_491 = $signed(_T_75963); // @[Modules.scala 65:57:@29764.4]
  assign buffer_12_206 = {{6{io_in_413[4]}},io_in_413}; // @[Modules.scala 32:22:@8.4]
  assign _T_75974 = $signed(buffer_12_206) + $signed(buffer_0_207); // @[Modules.scala 65:57:@29778.4]
  assign _T_75975 = _T_75974[10:0]; // @[Modules.scala 65:57:@29779.4]
  assign buffer_12_495 = $signed(_T_75975); // @[Modules.scala 65:57:@29780.4]
  assign _T_75980 = $signed(buffer_3_210) + $signed(11'sh0); // @[Modules.scala 65:57:@29786.4]
  assign _T_75981 = _T_75980[10:0]; // @[Modules.scala 65:57:@29787.4]
  assign buffer_12_497 = $signed(_T_75981); // @[Modules.scala 65:57:@29788.4]
  assign _T_75995 = $signed(buffer_0_220) + $signed(buffer_1_221); // @[Modules.scala 65:57:@29806.4]
  assign _T_75996 = _T_75995[10:0]; // @[Modules.scala 65:57:@29807.4]
  assign buffer_12_502 = $signed(_T_75996); // @[Modules.scala 65:57:@29808.4]
  assign _T_76010 = $signed(buffer_0_230) + $signed(11'sh0); // @[Modules.scala 65:57:@29826.4]
  assign _T_76011 = _T_76010[10:0]; // @[Modules.scala 65:57:@29827.4]
  assign buffer_12_507 = $signed(_T_76011); // @[Modules.scala 65:57:@29828.4]
  assign _T_76016 = $signed(buffer_1_234) + $signed(11'sh0); // @[Modules.scala 65:57:@29834.4]
  assign _T_76017 = _T_76016[10:0]; // @[Modules.scala 65:57:@29835.4]
  assign buffer_12_509 = $signed(_T_76017); // @[Modules.scala 65:57:@29836.4]
  assign buffer_12_238 = {{6{io_in_476[4]}},io_in_476}; // @[Modules.scala 32:22:@8.4]
  assign _T_76022 = $signed(buffer_12_238) + $signed(11'sh0); // @[Modules.scala 65:57:@29842.4]
  assign _T_76023 = _T_76022[10:0]; // @[Modules.scala 65:57:@29843.4]
  assign buffer_12_511 = $signed(_T_76023); // @[Modules.scala 65:57:@29844.4]
  assign buffer_12_244 = {{6{io_in_488[4]}},io_in_488}; // @[Modules.scala 32:22:@8.4]
  assign buffer_12_245 = {{6{io_in_491[4]}},io_in_491}; // @[Modules.scala 32:22:@8.4]
  assign _T_76031 = $signed(buffer_12_244) + $signed(buffer_12_245); // @[Modules.scala 65:57:@29854.4]
  assign _T_76032 = _T_76031[10:0]; // @[Modules.scala 65:57:@29855.4]
  assign buffer_12_514 = $signed(_T_76032); // @[Modules.scala 65:57:@29856.4]
  assign _T_76043 = $signed(buffer_3_252) + $signed(11'sh0); // @[Modules.scala 65:57:@29870.4]
  assign _T_76044 = _T_76043[10:0]; // @[Modules.scala 65:57:@29871.4]
  assign buffer_12_518 = $signed(_T_76044); // @[Modules.scala 65:57:@29872.4]
  assign _T_76046 = $signed(buffer_8_254) + $signed(buffer_10_255); // @[Modules.scala 65:57:@29874.4]
  assign _T_76047 = _T_76046[10:0]; // @[Modules.scala 65:57:@29875.4]
  assign buffer_12_519 = $signed(_T_76047); // @[Modules.scala 65:57:@29876.4]
  assign _T_76052 = $signed(buffer_2_258) + $signed(buffer_4_259); // @[Modules.scala 65:57:@29882.4]
  assign _T_76053 = _T_76052[10:0]; // @[Modules.scala 65:57:@29883.4]
  assign buffer_12_521 = $signed(_T_76053); // @[Modules.scala 65:57:@29884.4]
  assign _T_76058 = $signed(buffer_7_262) + $signed(buffer_0_263); // @[Modules.scala 65:57:@29890.4]
  assign _T_76059 = _T_76058[10:0]; // @[Modules.scala 65:57:@29891.4]
  assign buffer_12_523 = $signed(_T_76059); // @[Modules.scala 65:57:@29892.4]
  assign _T_76064 = $signed(buffer_1_266) + $signed(11'sh0); // @[Modules.scala 65:57:@29898.4]
  assign _T_76065 = _T_76064[10:0]; // @[Modules.scala 65:57:@29899.4]
  assign buffer_12_525 = $signed(_T_76065); // @[Modules.scala 65:57:@29900.4]
  assign _T_76076 = $signed(11'sh0) + $signed(buffer_2_275); // @[Modules.scala 65:57:@29914.4]
  assign _T_76077 = _T_76076[10:0]; // @[Modules.scala 65:57:@29915.4]
  assign buffer_12_529 = $signed(_T_76077); // @[Modules.scala 65:57:@29916.4]
  assign buffer_12_280 = {{6{_T_75492[4]}},_T_75492}; // @[Modules.scala 32:22:@8.4]
  assign _T_76085 = $signed(buffer_12_280) + $signed(11'sh0); // @[Modules.scala 65:57:@29926.4]
  assign _T_76086 = _T_76085[10:0]; // @[Modules.scala 65:57:@29927.4]
  assign buffer_12_532 = $signed(_T_76086); // @[Modules.scala 65:57:@29928.4]
  assign buffer_12_288 = {{6{io_in_577[4]}},io_in_577}; // @[Modules.scala 32:22:@8.4]
  assign _T_76097 = $signed(buffer_12_288) + $signed(buffer_1_289); // @[Modules.scala 65:57:@29942.4]
  assign _T_76098 = _T_76097[10:0]; // @[Modules.scala 65:57:@29943.4]
  assign buffer_12_536 = $signed(_T_76098); // @[Modules.scala 65:57:@29944.4]
  assign _T_76106 = $signed(buffer_2_294) + $signed(buffer_1_295); // @[Modules.scala 65:57:@29954.4]
  assign _T_76107 = _T_76106[10:0]; // @[Modules.scala 65:57:@29955.4]
  assign buffer_12_539 = $signed(_T_76107); // @[Modules.scala 65:57:@29956.4]
  assign buffer_12_296 = {{6{io_in_593[4]}},io_in_593}; // @[Modules.scala 32:22:@8.4]
  assign _T_76109 = $signed(buffer_12_296) + $signed(buffer_2_297); // @[Modules.scala 65:57:@29958.4]
  assign _T_76110 = _T_76109[10:0]; // @[Modules.scala 65:57:@29959.4]
  assign buffer_12_540 = $signed(_T_76110); // @[Modules.scala 65:57:@29960.4]
  assign _T_76112 = $signed(buffer_8_298) + $signed(buffer_1_299); // @[Modules.scala 65:57:@29962.4]
  assign _T_76113 = _T_76112[10:0]; // @[Modules.scala 65:57:@29963.4]
  assign buffer_12_541 = $signed(_T_76113); // @[Modules.scala 65:57:@29964.4]
  assign buffer_12_309 = {{6{io_in_619[4]}},io_in_619}; // @[Modules.scala 32:22:@8.4]
  assign _T_76127 = $signed(buffer_2_308) + $signed(buffer_12_309); // @[Modules.scala 65:57:@29982.4]
  assign _T_76128 = _T_76127[10:0]; // @[Modules.scala 65:57:@29983.4]
  assign buffer_12_546 = $signed(_T_76128); // @[Modules.scala 65:57:@29984.4]
  assign _T_76148 = $signed(buffer_10_322) + $signed(11'sh0); // @[Modules.scala 65:57:@30010.4]
  assign _T_76149 = _T_76148[10:0]; // @[Modules.scala 65:57:@30011.4]
  assign buffer_12_553 = $signed(_T_76149); // @[Modules.scala 65:57:@30012.4]
  assign _T_76166 = $signed(buffer_0_334) + $signed(buffer_4_335); // @[Modules.scala 65:57:@30034.4]
  assign _T_76167 = _T_76166[10:0]; // @[Modules.scala 65:57:@30035.4]
  assign buffer_12_559 = $signed(_T_76167); // @[Modules.scala 65:57:@30036.4]
  assign _T_76175 = $signed(buffer_1_340) + $signed(11'sh0); // @[Modules.scala 65:57:@30046.4]
  assign _T_76176 = _T_76175[10:0]; // @[Modules.scala 65:57:@30047.4]
  assign buffer_12_562 = $signed(_T_76176); // @[Modules.scala 65:57:@30048.4]
  assign _T_76178 = $signed(buffer_1_342) + $signed(11'sh0); // @[Modules.scala 65:57:@30050.4]
  assign _T_76179 = _T_76178[10:0]; // @[Modules.scala 65:57:@30051.4]
  assign buffer_12_563 = $signed(_T_76179); // @[Modules.scala 65:57:@30052.4]
  assign _T_76187 = $signed(buffer_0_348) + $signed(buffer_4_349); // @[Modules.scala 65:57:@30062.4]
  assign _T_76188 = _T_76187[10:0]; // @[Modules.scala 65:57:@30063.4]
  assign buffer_12_566 = $signed(_T_76188); // @[Modules.scala 65:57:@30064.4]
  assign _T_76190 = $signed(buffer_0_350) + $signed(11'sh0); // @[Modules.scala 65:57:@30066.4]
  assign _T_76191 = _T_76190[10:0]; // @[Modules.scala 65:57:@30067.4]
  assign buffer_12_567 = $signed(_T_76191); // @[Modules.scala 65:57:@30068.4]
  assign _T_76211 = $signed(buffer_0_364) + $signed(buffer_3_365); // @[Modules.scala 65:57:@30094.4]
  assign _T_76212 = _T_76211[10:0]; // @[Modules.scala 65:57:@30095.4]
  assign buffer_12_574 = $signed(_T_76212); // @[Modules.scala 65:57:@30096.4]
  assign _T_76229 = $signed(11'sh0) + $signed(buffer_0_377); // @[Modules.scala 65:57:@30118.4]
  assign _T_76230 = _T_76229[10:0]; // @[Modules.scala 65:57:@30119.4]
  assign buffer_12_580 = $signed(_T_76230); // @[Modules.scala 65:57:@30120.4]
  assign _T_76232 = $signed(buffer_3_378) + $signed(buffer_8_379); // @[Modules.scala 65:57:@30122.4]
  assign _T_76233 = _T_76232[10:0]; // @[Modules.scala 65:57:@30123.4]
  assign buffer_12_581 = $signed(_T_76233); // @[Modules.scala 65:57:@30124.4]
  assign _T_76238 = $signed(buffer_8_382) + $signed(buffer_4_383); // @[Modules.scala 65:57:@30130.4]
  assign _T_76239 = _T_76238[10:0]; // @[Modules.scala 65:57:@30131.4]
  assign buffer_12_583 = $signed(_T_76239); // @[Modules.scala 65:57:@30132.4]
  assign buffer_12_388 = {{6{io_in_776[4]}},io_in_776}; // @[Modules.scala 32:22:@8.4]
  assign _T_76247 = $signed(buffer_12_388) + $signed(11'sh0); // @[Modules.scala 65:57:@30142.4]
  assign _T_76248 = _T_76247[10:0]; // @[Modules.scala 65:57:@30143.4]
  assign buffer_12_586 = $signed(_T_76248); // @[Modules.scala 65:57:@30144.4]
  assign _T_76253 = $signed(buffer_12_392) + $signed(buffer_0_395); // @[Modules.scala 68:83:@30150.4]
  assign _T_76254 = _T_76253[10:0]; // @[Modules.scala 68:83:@30151.4]
  assign buffer_12_588 = $signed(_T_76254); // @[Modules.scala 68:83:@30152.4]
  assign _T_76256 = $signed(buffer_1_394) + $signed(buffer_12_395); // @[Modules.scala 68:83:@30154.4]
  assign _T_76257 = _T_76256[10:0]; // @[Modules.scala 68:83:@30155.4]
  assign buffer_12_589 = $signed(_T_76257); // @[Modules.scala 68:83:@30156.4]
  assign _T_76259 = $signed(buffer_12_396) + $signed(buffer_12_397); // @[Modules.scala 68:83:@30158.4]
  assign _T_76260 = _T_76259[10:0]; // @[Modules.scala 68:83:@30159.4]
  assign buffer_12_590 = $signed(_T_76260); // @[Modules.scala 68:83:@30160.4]
  assign _T_76262 = $signed(buffer_12_398) + $signed(buffer_12_399); // @[Modules.scala 68:83:@30162.4]
  assign _T_76263 = _T_76262[10:0]; // @[Modules.scala 68:83:@30163.4]
  assign buffer_12_591 = $signed(_T_76263); // @[Modules.scala 68:83:@30164.4]
  assign _T_76274 = $signed(buffer_1_406) + $signed(buffer_7_407); // @[Modules.scala 68:83:@30178.4]
  assign _T_76275 = _T_76274[10:0]; // @[Modules.scala 68:83:@30179.4]
  assign buffer_12_595 = $signed(_T_76275); // @[Modules.scala 68:83:@30180.4]
  assign _T_76283 = $signed(buffer_1_412) + $signed(buffer_4_413); // @[Modules.scala 68:83:@30190.4]
  assign _T_76284 = _T_76283[10:0]; // @[Modules.scala 68:83:@30191.4]
  assign buffer_12_598 = $signed(_T_76284); // @[Modules.scala 68:83:@30192.4]
  assign _T_76292 = $signed(buffer_0_418) + $signed(buffer_12_419); // @[Modules.scala 68:83:@30202.4]
  assign _T_76293 = _T_76292[10:0]; // @[Modules.scala 68:83:@30203.4]
  assign buffer_12_601 = $signed(_T_76293); // @[Modules.scala 68:83:@30204.4]
  assign _T_76295 = $signed(buffer_0_395) + $signed(buffer_12_421); // @[Modules.scala 68:83:@30206.4]
  assign _T_76296 = _T_76295[10:0]; // @[Modules.scala 68:83:@30207.4]
  assign buffer_12_602 = $signed(_T_76296); // @[Modules.scala 68:83:@30208.4]
  assign _T_76298 = $signed(buffer_4_422) + $signed(buffer_12_423); // @[Modules.scala 68:83:@30210.4]
  assign _T_76299 = _T_76298[10:0]; // @[Modules.scala 68:83:@30211.4]
  assign buffer_12_603 = $signed(_T_76299); // @[Modules.scala 68:83:@30212.4]
  assign _T_76301 = $signed(buffer_0_395) + $signed(buffer_12_425); // @[Modules.scala 68:83:@30214.4]
  assign _T_76302 = _T_76301[10:0]; // @[Modules.scala 68:83:@30215.4]
  assign buffer_12_604 = $signed(_T_76302); // @[Modules.scala 68:83:@30216.4]
  assign _T_76304 = $signed(buffer_12_426) + $signed(buffer_0_427); // @[Modules.scala 68:83:@30218.4]
  assign _T_76305 = _T_76304[10:0]; // @[Modules.scala 68:83:@30219.4]
  assign buffer_12_605 = $signed(_T_76305); // @[Modules.scala 68:83:@30220.4]
  assign _T_76307 = $signed(buffer_12_428) + $signed(buffer_12_429); // @[Modules.scala 68:83:@30222.4]
  assign _T_76308 = _T_76307[10:0]; // @[Modules.scala 68:83:@30223.4]
  assign buffer_12_606 = $signed(_T_76308); // @[Modules.scala 68:83:@30224.4]
  assign _T_76310 = $signed(buffer_4_430) + $signed(buffer_12_431); // @[Modules.scala 68:83:@30226.4]
  assign _T_76311 = _T_76310[10:0]; // @[Modules.scala 68:83:@30227.4]
  assign buffer_12_607 = $signed(_T_76311); // @[Modules.scala 68:83:@30228.4]
  assign _T_76313 = $signed(buffer_5_432) + $signed(buffer_12_433); // @[Modules.scala 68:83:@30230.4]
  assign _T_76314 = _T_76313[10:0]; // @[Modules.scala 68:83:@30231.4]
  assign buffer_12_608 = $signed(_T_76314); // @[Modules.scala 68:83:@30232.4]
  assign _T_76319 = $signed(buffer_0_395) + $signed(buffer_5_437); // @[Modules.scala 68:83:@30238.4]
  assign _T_76320 = _T_76319[10:0]; // @[Modules.scala 68:83:@30239.4]
  assign buffer_12_610 = $signed(_T_76320); // @[Modules.scala 68:83:@30240.4]
  assign _T_76322 = $signed(buffer_12_438) + $signed(buffer_0_395); // @[Modules.scala 68:83:@30242.4]
  assign _T_76323 = _T_76322[10:0]; // @[Modules.scala 68:83:@30243.4]
  assign buffer_12_611 = $signed(_T_76323); // @[Modules.scala 68:83:@30244.4]
  assign _T_76328 = $signed(buffer_12_442) + $signed(buffer_12_443); // @[Modules.scala 68:83:@30250.4]
  assign _T_76329 = _T_76328[10:0]; // @[Modules.scala 68:83:@30251.4]
  assign buffer_12_613 = $signed(_T_76329); // @[Modules.scala 68:83:@30252.4]
  assign _T_76331 = $signed(buffer_1_444) + $signed(buffer_12_445); // @[Modules.scala 68:83:@30254.4]
  assign _T_76332 = _T_76331[10:0]; // @[Modules.scala 68:83:@30255.4]
  assign buffer_12_614 = $signed(_T_76332); // @[Modules.scala 68:83:@30256.4]
  assign _T_76337 = $signed(buffer_12_448) + $signed(buffer_7_449); // @[Modules.scala 68:83:@30262.4]
  assign _T_76338 = _T_76337[10:0]; // @[Modules.scala 68:83:@30263.4]
  assign buffer_12_616 = $signed(_T_76338); // @[Modules.scala 68:83:@30264.4]
  assign _T_76340 = $signed(buffer_12_450) + $signed(buffer_12_451); // @[Modules.scala 68:83:@30266.4]
  assign _T_76341 = _T_76340[10:0]; // @[Modules.scala 68:83:@30267.4]
  assign buffer_12_617 = $signed(_T_76341); // @[Modules.scala 68:83:@30268.4]
  assign _T_76343 = $signed(buffer_1_452) + $signed(buffer_9_453); // @[Modules.scala 68:83:@30270.4]
  assign _T_76344 = _T_76343[10:0]; // @[Modules.scala 68:83:@30271.4]
  assign buffer_12_618 = $signed(_T_76344); // @[Modules.scala 68:83:@30272.4]
  assign _T_76346 = $signed(buffer_0_395) + $signed(buffer_12_455); // @[Modules.scala 68:83:@30274.4]
  assign _T_76347 = _T_76346[10:0]; // @[Modules.scala 68:83:@30275.4]
  assign buffer_12_619 = $signed(_T_76347); // @[Modules.scala 68:83:@30276.4]
  assign _T_76349 = $signed(buffer_12_456) + $signed(buffer_12_457); // @[Modules.scala 68:83:@30278.4]
  assign _T_76350 = _T_76349[10:0]; // @[Modules.scala 68:83:@30279.4]
  assign buffer_12_620 = $signed(_T_76350); // @[Modules.scala 68:83:@30280.4]
  assign _T_76352 = $signed(buffer_12_458) + $signed(buffer_12_459); // @[Modules.scala 68:83:@30282.4]
  assign _T_76353 = _T_76352[10:0]; // @[Modules.scala 68:83:@30283.4]
  assign buffer_12_621 = $signed(_T_76353); // @[Modules.scala 68:83:@30284.4]
  assign _T_76358 = $signed(buffer_12_462) + $signed(buffer_0_395); // @[Modules.scala 68:83:@30290.4]
  assign _T_76359 = _T_76358[10:0]; // @[Modules.scala 68:83:@30291.4]
  assign buffer_12_623 = $signed(_T_76359); // @[Modules.scala 68:83:@30292.4]
  assign _T_76361 = $signed(buffer_0_395) + $signed(buffer_7_465); // @[Modules.scala 68:83:@30294.4]
  assign _T_76362 = _T_76361[10:0]; // @[Modules.scala 68:83:@30295.4]
  assign buffer_12_624 = $signed(_T_76362); // @[Modules.scala 68:83:@30296.4]
  assign _T_76364 = $signed(buffer_12_466) + $signed(buffer_12_467); // @[Modules.scala 68:83:@30298.4]
  assign _T_76365 = _T_76364[10:0]; // @[Modules.scala 68:83:@30299.4]
  assign buffer_12_625 = $signed(_T_76365); // @[Modules.scala 68:83:@30300.4]
  assign _T_76367 = $signed(buffer_0_395) + $signed(buffer_12_469); // @[Modules.scala 68:83:@30302.4]
  assign _T_76368 = _T_76367[10:0]; // @[Modules.scala 68:83:@30303.4]
  assign buffer_12_626 = $signed(_T_76368); // @[Modules.scala 68:83:@30304.4]
  assign _T_76373 = $signed(buffer_0_395) + $signed(buffer_12_473); // @[Modules.scala 68:83:@30310.4]
  assign _T_76374 = _T_76373[10:0]; // @[Modules.scala 68:83:@30311.4]
  assign buffer_12_628 = $signed(_T_76374); // @[Modules.scala 68:83:@30312.4]
  assign _T_76376 = $signed(buffer_12_474) + $signed(buffer_12_475); // @[Modules.scala 68:83:@30314.4]
  assign _T_76377 = _T_76376[10:0]; // @[Modules.scala 68:83:@30315.4]
  assign buffer_12_629 = $signed(_T_76377); // @[Modules.scala 68:83:@30316.4]
  assign _T_76379 = $signed(buffer_12_476) + $signed(buffer_0_395); // @[Modules.scala 68:83:@30318.4]
  assign _T_76380 = _T_76379[10:0]; // @[Modules.scala 68:83:@30319.4]
  assign buffer_12_630 = $signed(_T_76380); // @[Modules.scala 68:83:@30320.4]
  assign _T_76385 = $signed(buffer_0_395) + $signed(buffer_0_481); // @[Modules.scala 68:83:@30326.4]
  assign _T_76386 = _T_76385[10:0]; // @[Modules.scala 68:83:@30327.4]
  assign buffer_12_632 = $signed(_T_76386); // @[Modules.scala 68:83:@30328.4]
  assign _T_76388 = $signed(buffer_11_482) + $signed(buffer_3_483); // @[Modules.scala 68:83:@30330.4]
  assign _T_76389 = _T_76388[10:0]; // @[Modules.scala 68:83:@30331.4]
  assign buffer_12_633 = $signed(_T_76389); // @[Modules.scala 68:83:@30332.4]
  assign _T_76397 = $signed(buffer_0_488) + $signed(buffer_9_489); // @[Modules.scala 68:83:@30342.4]
  assign _T_76398 = _T_76397[10:0]; // @[Modules.scala 68:83:@30343.4]
  assign buffer_12_636 = $signed(_T_76398); // @[Modules.scala 68:83:@30344.4]
  assign _T_76400 = $signed(buffer_12_490) + $signed(buffer_12_491); // @[Modules.scala 68:83:@30346.4]
  assign _T_76401 = _T_76400[10:0]; // @[Modules.scala 68:83:@30347.4]
  assign buffer_12_637 = $signed(_T_76401); // @[Modules.scala 68:83:@30348.4]
  assign _T_76403 = $signed(buffer_4_492) + $signed(buffer_0_395); // @[Modules.scala 68:83:@30350.4]
  assign _T_76404 = _T_76403[10:0]; // @[Modules.scala 68:83:@30351.4]
  assign buffer_12_638 = $signed(_T_76404); // @[Modules.scala 68:83:@30352.4]
  assign _T_76406 = $signed(buffer_1_494) + $signed(buffer_12_495); // @[Modules.scala 68:83:@30354.4]
  assign _T_76407 = _T_76406[10:0]; // @[Modules.scala 68:83:@30355.4]
  assign buffer_12_639 = $signed(_T_76407); // @[Modules.scala 68:83:@30356.4]
  assign _T_76409 = $signed(buffer_10_496) + $signed(buffer_12_497); // @[Modules.scala 68:83:@30358.4]
  assign _T_76410 = _T_76409[10:0]; // @[Modules.scala 68:83:@30359.4]
  assign buffer_12_640 = $signed(_T_76410); // @[Modules.scala 68:83:@30360.4]
  assign _T_76418 = $signed(buffer_12_502) + $signed(buffer_3_503); // @[Modules.scala 68:83:@30370.4]
  assign _T_76419 = _T_76418[10:0]; // @[Modules.scala 68:83:@30371.4]
  assign buffer_12_643 = $signed(_T_76419); // @[Modules.scala 68:83:@30372.4]
  assign _T_76424 = $signed(buffer_0_506) + $signed(buffer_12_507); // @[Modules.scala 68:83:@30378.4]
  assign _T_76425 = _T_76424[10:0]; // @[Modules.scala 68:83:@30379.4]
  assign buffer_12_645 = $signed(_T_76425); // @[Modules.scala 68:83:@30380.4]
  assign _T_76427 = $signed(buffer_0_508) + $signed(buffer_12_509); // @[Modules.scala 68:83:@30382.4]
  assign _T_76428 = _T_76427[10:0]; // @[Modules.scala 68:83:@30383.4]
  assign buffer_12_646 = $signed(_T_76428); // @[Modules.scala 68:83:@30384.4]
  assign _T_76430 = $signed(buffer_3_510) + $signed(buffer_12_511); // @[Modules.scala 68:83:@30386.4]
  assign _T_76431 = _T_76430[10:0]; // @[Modules.scala 68:83:@30387.4]
  assign buffer_12_647 = $signed(_T_76431); // @[Modules.scala 68:83:@30388.4]
  assign _T_76433 = $signed(buffer_4_512) + $signed(buffer_0_513); // @[Modules.scala 68:83:@30390.4]
  assign _T_76434 = _T_76433[10:0]; // @[Modules.scala 68:83:@30391.4]
  assign buffer_12_648 = $signed(_T_76434); // @[Modules.scala 68:83:@30392.4]
  assign _T_76436 = $signed(buffer_12_514) + $signed(buffer_8_515); // @[Modules.scala 68:83:@30394.4]
  assign _T_76437 = _T_76436[10:0]; // @[Modules.scala 68:83:@30395.4]
  assign buffer_12_649 = $signed(_T_76437); // @[Modules.scala 68:83:@30396.4]
  assign _T_76442 = $signed(buffer_12_518) + $signed(buffer_12_519); // @[Modules.scala 68:83:@30402.4]
  assign _T_76443 = _T_76442[10:0]; // @[Modules.scala 68:83:@30403.4]
  assign buffer_12_651 = $signed(_T_76443); // @[Modules.scala 68:83:@30404.4]
  assign _T_76445 = $signed(buffer_0_520) + $signed(buffer_12_521); // @[Modules.scala 68:83:@30406.4]
  assign _T_76446 = _T_76445[10:0]; // @[Modules.scala 68:83:@30407.4]
  assign buffer_12_652 = $signed(_T_76446); // @[Modules.scala 68:83:@30408.4]
  assign _T_76448 = $signed(buffer_4_522) + $signed(buffer_12_523); // @[Modules.scala 68:83:@30410.4]
  assign _T_76449 = _T_76448[10:0]; // @[Modules.scala 68:83:@30411.4]
  assign buffer_12_653 = $signed(_T_76449); // @[Modules.scala 68:83:@30412.4]
  assign _T_76451 = $signed(buffer_3_524) + $signed(buffer_12_525); // @[Modules.scala 68:83:@30414.4]
  assign _T_76452 = _T_76451[10:0]; // @[Modules.scala 68:83:@30415.4]
  assign buffer_12_654 = $signed(_T_76452); // @[Modules.scala 68:83:@30416.4]
  assign _T_76457 = $signed(buffer_7_528) + $signed(buffer_12_529); // @[Modules.scala 68:83:@30422.4]
  assign _T_76458 = _T_76457[10:0]; // @[Modules.scala 68:83:@30423.4]
  assign buffer_12_656 = $signed(_T_76458); // @[Modules.scala 68:83:@30424.4]
  assign _T_76463 = $signed(buffer_12_532) + $signed(buffer_3_533); // @[Modules.scala 68:83:@30430.4]
  assign _T_76464 = _T_76463[10:0]; // @[Modules.scala 68:83:@30431.4]
  assign buffer_12_658 = $signed(_T_76464); // @[Modules.scala 68:83:@30432.4]
  assign _T_76469 = $signed(buffer_12_536) + $signed(buffer_4_537); // @[Modules.scala 68:83:@30438.4]
  assign _T_76470 = _T_76469[10:0]; // @[Modules.scala 68:83:@30439.4]
  assign buffer_12_660 = $signed(_T_76470); // @[Modules.scala 68:83:@30440.4]
  assign _T_76472 = $signed(buffer_3_538) + $signed(buffer_12_539); // @[Modules.scala 68:83:@30442.4]
  assign _T_76473 = _T_76472[10:0]; // @[Modules.scala 68:83:@30443.4]
  assign buffer_12_661 = $signed(_T_76473); // @[Modules.scala 68:83:@30444.4]
  assign _T_76475 = $signed(buffer_12_540) + $signed(buffer_12_541); // @[Modules.scala 68:83:@30446.4]
  assign _T_76476 = _T_76475[10:0]; // @[Modules.scala 68:83:@30447.4]
  assign buffer_12_662 = $signed(_T_76476); // @[Modules.scala 68:83:@30448.4]
  assign _T_76481 = $signed(buffer_4_544) + $signed(buffer_10_545); // @[Modules.scala 68:83:@30454.4]
  assign _T_76482 = _T_76481[10:0]; // @[Modules.scala 68:83:@30455.4]
  assign buffer_12_664 = $signed(_T_76482); // @[Modules.scala 68:83:@30456.4]
  assign _T_76484 = $signed(buffer_12_546) + $signed(buffer_3_547); // @[Modules.scala 68:83:@30458.4]
  assign _T_76485 = _T_76484[10:0]; // @[Modules.scala 68:83:@30459.4]
  assign buffer_12_665 = $signed(_T_76485); // @[Modules.scala 68:83:@30460.4]
  assign _T_76487 = $signed(buffer_8_548) + $signed(buffer_6_549); // @[Modules.scala 68:83:@30462.4]
  assign _T_76488 = _T_76487[10:0]; // @[Modules.scala 68:83:@30463.4]
  assign buffer_12_666 = $signed(_T_76488); // @[Modules.scala 68:83:@30464.4]
  assign _T_76490 = $signed(buffer_2_550) + $signed(buffer_3_551); // @[Modules.scala 68:83:@30466.4]
  assign _T_76491 = _T_76490[10:0]; // @[Modules.scala 68:83:@30467.4]
  assign buffer_12_667 = $signed(_T_76491); // @[Modules.scala 68:83:@30468.4]
  assign _T_76493 = $signed(buffer_0_552) + $signed(buffer_12_553); // @[Modules.scala 68:83:@30470.4]
  assign _T_76494 = _T_76493[10:0]; // @[Modules.scala 68:83:@30471.4]
  assign buffer_12_668 = $signed(_T_76494); // @[Modules.scala 68:83:@30472.4]
  assign _T_76496 = $signed(buffer_1_554) + $signed(buffer_8_555); // @[Modules.scala 68:83:@30474.4]
  assign _T_76497 = _T_76496[10:0]; // @[Modules.scala 68:83:@30475.4]
  assign buffer_12_669 = $signed(_T_76497); // @[Modules.scala 68:83:@30476.4]
  assign _T_76502 = $signed(buffer_5_558) + $signed(buffer_12_559); // @[Modules.scala 68:83:@30482.4]
  assign _T_76503 = _T_76502[10:0]; // @[Modules.scala 68:83:@30483.4]
  assign buffer_12_671 = $signed(_T_76503); // @[Modules.scala 68:83:@30484.4]
  assign _T_76508 = $signed(buffer_12_562) + $signed(buffer_12_563); // @[Modules.scala 68:83:@30490.4]
  assign _T_76509 = _T_76508[10:0]; // @[Modules.scala 68:83:@30491.4]
  assign buffer_12_673 = $signed(_T_76509); // @[Modules.scala 68:83:@30492.4]
  assign _T_76514 = $signed(buffer_12_566) + $signed(buffer_12_567); // @[Modules.scala 68:83:@30498.4]
  assign _T_76515 = _T_76514[10:0]; // @[Modules.scala 68:83:@30499.4]
  assign buffer_12_675 = $signed(_T_76515); // @[Modules.scala 68:83:@30500.4]
  assign _T_76526 = $signed(buffer_12_574) + $signed(buffer_0_395); // @[Modules.scala 68:83:@30514.4]
  assign _T_76527 = _T_76526[10:0]; // @[Modules.scala 68:83:@30515.4]
  assign buffer_12_679 = $signed(_T_76527); // @[Modules.scala 68:83:@30516.4]
  assign _T_76535 = $signed(buffer_12_580) + $signed(buffer_12_581); // @[Modules.scala 68:83:@30526.4]
  assign _T_76536 = _T_76535[10:0]; // @[Modules.scala 68:83:@30527.4]
  assign buffer_12_682 = $signed(_T_76536); // @[Modules.scala 68:83:@30528.4]
  assign _T_76538 = $signed(buffer_1_582) + $signed(buffer_12_583); // @[Modules.scala 68:83:@30530.4]
  assign _T_76539 = _T_76538[10:0]; // @[Modules.scala 68:83:@30531.4]
  assign buffer_12_683 = $signed(_T_76539); // @[Modules.scala 68:83:@30532.4]
  assign _T_76544 = $signed(buffer_12_586) + $signed(buffer_0_587); // @[Modules.scala 68:83:@30538.4]
  assign _T_76545 = _T_76544[10:0]; // @[Modules.scala 68:83:@30539.4]
  assign buffer_12_685 = $signed(_T_76545); // @[Modules.scala 68:83:@30540.4]
  assign _T_76547 = $signed(buffer_12_588) + $signed(buffer_12_589); // @[Modules.scala 71:109:@30542.4]
  assign _T_76548 = _T_76547[10:0]; // @[Modules.scala 71:109:@30543.4]
  assign buffer_12_686 = $signed(_T_76548); // @[Modules.scala 71:109:@30544.4]
  assign _T_76550 = $signed(buffer_12_590) + $signed(buffer_12_591); // @[Modules.scala 71:109:@30546.4]
  assign _T_76551 = _T_76550[10:0]; // @[Modules.scala 71:109:@30547.4]
  assign buffer_12_687 = $signed(_T_76551); // @[Modules.scala 71:109:@30548.4]
  assign _T_76553 = $signed(buffer_1_592) + $signed(buffer_9_593); // @[Modules.scala 71:109:@30550.4]
  assign _T_76554 = _T_76553[10:0]; // @[Modules.scala 71:109:@30551.4]
  assign buffer_12_688 = $signed(_T_76554); // @[Modules.scala 71:109:@30552.4]
  assign _T_76556 = $signed(buffer_2_594) + $signed(buffer_12_595); // @[Modules.scala 71:109:@30554.4]
  assign _T_76557 = _T_76556[10:0]; // @[Modules.scala 71:109:@30555.4]
  assign buffer_12_689 = $signed(_T_76557); // @[Modules.scala 71:109:@30556.4]
  assign _T_76562 = $signed(buffer_12_598) + $signed(buffer_1_599); // @[Modules.scala 71:109:@30562.4]
  assign _T_76563 = _T_76562[10:0]; // @[Modules.scala 71:109:@30563.4]
  assign buffer_12_691 = $signed(_T_76563); // @[Modules.scala 71:109:@30564.4]
  assign _T_76565 = $signed(buffer_1_600) + $signed(buffer_12_601); // @[Modules.scala 71:109:@30566.4]
  assign _T_76566 = _T_76565[10:0]; // @[Modules.scala 71:109:@30567.4]
  assign buffer_12_692 = $signed(_T_76566); // @[Modules.scala 71:109:@30568.4]
  assign _T_76568 = $signed(buffer_12_602) + $signed(buffer_12_603); // @[Modules.scala 71:109:@30570.4]
  assign _T_76569 = _T_76568[10:0]; // @[Modules.scala 71:109:@30571.4]
  assign buffer_12_693 = $signed(_T_76569); // @[Modules.scala 71:109:@30572.4]
  assign _T_76571 = $signed(buffer_12_604) + $signed(buffer_12_605); // @[Modules.scala 71:109:@30574.4]
  assign _T_76572 = _T_76571[10:0]; // @[Modules.scala 71:109:@30575.4]
  assign buffer_12_694 = $signed(_T_76572); // @[Modules.scala 71:109:@30576.4]
  assign _T_76574 = $signed(buffer_12_606) + $signed(buffer_12_607); // @[Modules.scala 71:109:@30578.4]
  assign _T_76575 = _T_76574[10:0]; // @[Modules.scala 71:109:@30579.4]
  assign buffer_12_695 = $signed(_T_76575); // @[Modules.scala 71:109:@30580.4]
  assign _T_76577 = $signed(buffer_12_608) + $signed(buffer_0_609); // @[Modules.scala 71:109:@30582.4]
  assign _T_76578 = _T_76577[10:0]; // @[Modules.scala 71:109:@30583.4]
  assign buffer_12_696 = $signed(_T_76578); // @[Modules.scala 71:109:@30584.4]
  assign _T_76580 = $signed(buffer_12_610) + $signed(buffer_12_611); // @[Modules.scala 71:109:@30586.4]
  assign _T_76581 = _T_76580[10:0]; // @[Modules.scala 71:109:@30587.4]
  assign buffer_12_697 = $signed(_T_76581); // @[Modules.scala 71:109:@30588.4]
  assign _T_76583 = $signed(buffer_0_612) + $signed(buffer_12_613); // @[Modules.scala 71:109:@30590.4]
  assign _T_76584 = _T_76583[10:0]; // @[Modules.scala 71:109:@30591.4]
  assign buffer_12_698 = $signed(_T_76584); // @[Modules.scala 71:109:@30592.4]
  assign _T_76586 = $signed(buffer_12_614) + $signed(buffer_0_593); // @[Modules.scala 71:109:@30594.4]
  assign _T_76587 = _T_76586[10:0]; // @[Modules.scala 71:109:@30595.4]
  assign buffer_12_699 = $signed(_T_76587); // @[Modules.scala 71:109:@30596.4]
  assign _T_76589 = $signed(buffer_12_616) + $signed(buffer_12_617); // @[Modules.scala 71:109:@30598.4]
  assign _T_76590 = _T_76589[10:0]; // @[Modules.scala 71:109:@30599.4]
  assign buffer_12_700 = $signed(_T_76590); // @[Modules.scala 71:109:@30600.4]
  assign _T_76592 = $signed(buffer_12_618) + $signed(buffer_12_619); // @[Modules.scala 71:109:@30602.4]
  assign _T_76593 = _T_76592[10:0]; // @[Modules.scala 71:109:@30603.4]
  assign buffer_12_701 = $signed(_T_76593); // @[Modules.scala 71:109:@30604.4]
  assign _T_76595 = $signed(buffer_12_620) + $signed(buffer_12_621); // @[Modules.scala 71:109:@30606.4]
  assign _T_76596 = _T_76595[10:0]; // @[Modules.scala 71:109:@30607.4]
  assign buffer_12_702 = $signed(_T_76596); // @[Modules.scala 71:109:@30608.4]
  assign _T_76598 = $signed(buffer_6_622) + $signed(buffer_12_623); // @[Modules.scala 71:109:@30610.4]
  assign _T_76599 = _T_76598[10:0]; // @[Modules.scala 71:109:@30611.4]
  assign buffer_12_703 = $signed(_T_76599); // @[Modules.scala 71:109:@30612.4]
  assign _T_76601 = $signed(buffer_12_624) + $signed(buffer_12_625); // @[Modules.scala 71:109:@30614.4]
  assign _T_76602 = _T_76601[10:0]; // @[Modules.scala 71:109:@30615.4]
  assign buffer_12_704 = $signed(_T_76602); // @[Modules.scala 71:109:@30616.4]
  assign _T_76604 = $signed(buffer_12_626) + $signed(buffer_0_593); // @[Modules.scala 71:109:@30618.4]
  assign _T_76605 = _T_76604[10:0]; // @[Modules.scala 71:109:@30619.4]
  assign buffer_12_705 = $signed(_T_76605); // @[Modules.scala 71:109:@30620.4]
  assign _T_76607 = $signed(buffer_12_628) + $signed(buffer_12_629); // @[Modules.scala 71:109:@30622.4]
  assign _T_76608 = _T_76607[10:0]; // @[Modules.scala 71:109:@30623.4]
  assign buffer_12_706 = $signed(_T_76608); // @[Modules.scala 71:109:@30624.4]
  assign _T_76610 = $signed(buffer_12_630) + $signed(buffer_0_593); // @[Modules.scala 71:109:@30626.4]
  assign _T_76611 = _T_76610[10:0]; // @[Modules.scala 71:109:@30627.4]
  assign buffer_12_707 = $signed(_T_76611); // @[Modules.scala 71:109:@30628.4]
  assign _T_76613 = $signed(buffer_12_632) + $signed(buffer_12_633); // @[Modules.scala 71:109:@30630.4]
  assign _T_76614 = _T_76613[10:0]; // @[Modules.scala 71:109:@30631.4]
  assign buffer_12_708 = $signed(_T_76614); // @[Modules.scala 71:109:@30632.4]
  assign _T_76619 = $signed(buffer_12_636) + $signed(buffer_12_637); // @[Modules.scala 71:109:@30638.4]
  assign _T_76620 = _T_76619[10:0]; // @[Modules.scala 71:109:@30639.4]
  assign buffer_12_710 = $signed(_T_76620); // @[Modules.scala 71:109:@30640.4]
  assign _T_76622 = $signed(buffer_12_638) + $signed(buffer_12_639); // @[Modules.scala 71:109:@30642.4]
  assign _T_76623 = _T_76622[10:0]; // @[Modules.scala 71:109:@30643.4]
  assign buffer_12_711 = $signed(_T_76623); // @[Modules.scala 71:109:@30644.4]
  assign _T_76625 = $signed(buffer_12_640) + $signed(buffer_0_641); // @[Modules.scala 71:109:@30646.4]
  assign _T_76626 = _T_76625[10:0]; // @[Modules.scala 71:109:@30647.4]
  assign buffer_12_712 = $signed(_T_76626); // @[Modules.scala 71:109:@30648.4]
  assign _T_76628 = $signed(buffer_1_642) + $signed(buffer_12_643); // @[Modules.scala 71:109:@30650.4]
  assign _T_76629 = _T_76628[10:0]; // @[Modules.scala 71:109:@30651.4]
  assign buffer_12_713 = $signed(_T_76629); // @[Modules.scala 71:109:@30652.4]
  assign _T_76631 = $signed(buffer_6_644) + $signed(buffer_12_645); // @[Modules.scala 71:109:@30654.4]
  assign _T_76632 = _T_76631[10:0]; // @[Modules.scala 71:109:@30655.4]
  assign buffer_12_714 = $signed(_T_76632); // @[Modules.scala 71:109:@30656.4]
  assign _T_76634 = $signed(buffer_12_646) + $signed(buffer_12_647); // @[Modules.scala 71:109:@30658.4]
  assign _T_76635 = _T_76634[10:0]; // @[Modules.scala 71:109:@30659.4]
  assign buffer_12_715 = $signed(_T_76635); // @[Modules.scala 71:109:@30660.4]
  assign _T_76637 = $signed(buffer_12_648) + $signed(buffer_12_649); // @[Modules.scala 71:109:@30662.4]
  assign _T_76638 = _T_76637[10:0]; // @[Modules.scala 71:109:@30663.4]
  assign buffer_12_716 = $signed(_T_76638); // @[Modules.scala 71:109:@30664.4]
  assign _T_76640 = $signed(buffer_3_650) + $signed(buffer_12_651); // @[Modules.scala 71:109:@30666.4]
  assign _T_76641 = _T_76640[10:0]; // @[Modules.scala 71:109:@30667.4]
  assign buffer_12_717 = $signed(_T_76641); // @[Modules.scala 71:109:@30668.4]
  assign _T_76643 = $signed(buffer_12_652) + $signed(buffer_12_653); // @[Modules.scala 71:109:@30670.4]
  assign _T_76644 = _T_76643[10:0]; // @[Modules.scala 71:109:@30671.4]
  assign buffer_12_718 = $signed(_T_76644); // @[Modules.scala 71:109:@30672.4]
  assign _T_76646 = $signed(buffer_12_654) + $signed(buffer_9_655); // @[Modules.scala 71:109:@30674.4]
  assign _T_76647 = _T_76646[10:0]; // @[Modules.scala 71:109:@30675.4]
  assign buffer_12_719 = $signed(_T_76647); // @[Modules.scala 71:109:@30676.4]
  assign _T_76649 = $signed(buffer_12_656) + $signed(buffer_3_657); // @[Modules.scala 71:109:@30678.4]
  assign _T_76650 = _T_76649[10:0]; // @[Modules.scala 71:109:@30679.4]
  assign buffer_12_720 = $signed(_T_76650); // @[Modules.scala 71:109:@30680.4]
  assign _T_76652 = $signed(buffer_12_658) + $signed(buffer_1_659); // @[Modules.scala 71:109:@30682.4]
  assign _T_76653 = _T_76652[10:0]; // @[Modules.scala 71:109:@30683.4]
  assign buffer_12_721 = $signed(_T_76653); // @[Modules.scala 71:109:@30684.4]
  assign _T_76655 = $signed(buffer_12_660) + $signed(buffer_12_661); // @[Modules.scala 71:109:@30686.4]
  assign _T_76656 = _T_76655[10:0]; // @[Modules.scala 71:109:@30687.4]
  assign buffer_12_722 = $signed(_T_76656); // @[Modules.scala 71:109:@30688.4]
  assign _T_76658 = $signed(buffer_12_662) + $signed(buffer_0_663); // @[Modules.scala 71:109:@30690.4]
  assign _T_76659 = _T_76658[10:0]; // @[Modules.scala 71:109:@30691.4]
  assign buffer_12_723 = $signed(_T_76659); // @[Modules.scala 71:109:@30692.4]
  assign _T_76661 = $signed(buffer_12_664) + $signed(buffer_12_665); // @[Modules.scala 71:109:@30694.4]
  assign _T_76662 = _T_76661[10:0]; // @[Modules.scala 71:109:@30695.4]
  assign buffer_12_724 = $signed(_T_76662); // @[Modules.scala 71:109:@30696.4]
  assign _T_76664 = $signed(buffer_12_666) + $signed(buffer_12_667); // @[Modules.scala 71:109:@30698.4]
  assign _T_76665 = _T_76664[10:0]; // @[Modules.scala 71:109:@30699.4]
  assign buffer_12_725 = $signed(_T_76665); // @[Modules.scala 71:109:@30700.4]
  assign _T_76667 = $signed(buffer_12_668) + $signed(buffer_12_669); // @[Modules.scala 71:109:@30702.4]
  assign _T_76668 = _T_76667[10:0]; // @[Modules.scala 71:109:@30703.4]
  assign buffer_12_726 = $signed(_T_76668); // @[Modules.scala 71:109:@30704.4]
  assign _T_76670 = $signed(buffer_0_593) + $signed(buffer_12_671); // @[Modules.scala 71:109:@30706.4]
  assign _T_76671 = _T_76670[10:0]; // @[Modules.scala 71:109:@30707.4]
  assign buffer_12_727 = $signed(_T_76671); // @[Modules.scala 71:109:@30708.4]
  assign _T_76673 = $signed(buffer_2_672) + $signed(buffer_12_673); // @[Modules.scala 71:109:@30710.4]
  assign _T_76674 = _T_76673[10:0]; // @[Modules.scala 71:109:@30711.4]
  assign buffer_12_728 = $signed(_T_76674); // @[Modules.scala 71:109:@30712.4]
  assign _T_76676 = $signed(buffer_0_593) + $signed(buffer_12_675); // @[Modules.scala 71:109:@30714.4]
  assign _T_76677 = _T_76676[10:0]; // @[Modules.scala 71:109:@30715.4]
  assign buffer_12_729 = $signed(_T_76677); // @[Modules.scala 71:109:@30716.4]
  assign _T_76682 = $signed(buffer_9_678) + $signed(buffer_12_679); // @[Modules.scala 71:109:@30722.4]
  assign _T_76683 = _T_76682[10:0]; // @[Modules.scala 71:109:@30723.4]
  assign buffer_12_731 = $signed(_T_76683); // @[Modules.scala 71:109:@30724.4]
  assign _T_76688 = $signed(buffer_12_682) + $signed(buffer_12_683); // @[Modules.scala 71:109:@30730.4]
  assign _T_76689 = _T_76688[10:0]; // @[Modules.scala 71:109:@30731.4]
  assign buffer_12_733 = $signed(_T_76689); // @[Modules.scala 71:109:@30732.4]
  assign _T_76691 = $signed(buffer_3_684) + $signed(buffer_12_685); // @[Modules.scala 71:109:@30734.4]
  assign _T_76692 = _T_76691[10:0]; // @[Modules.scala 71:109:@30735.4]
  assign buffer_12_734 = $signed(_T_76692); // @[Modules.scala 71:109:@30736.4]
  assign _T_76694 = $signed(buffer_12_686) + $signed(buffer_12_687); // @[Modules.scala 78:156:@30739.4]
  assign _T_76695 = _T_76694[10:0]; // @[Modules.scala 78:156:@30740.4]
  assign buffer_12_736 = $signed(_T_76695); // @[Modules.scala 78:156:@30741.4]
  assign _T_76697 = $signed(buffer_12_736) + $signed(buffer_12_688); // @[Modules.scala 78:156:@30743.4]
  assign _T_76698 = _T_76697[10:0]; // @[Modules.scala 78:156:@30744.4]
  assign buffer_12_737 = $signed(_T_76698); // @[Modules.scala 78:156:@30745.4]
  assign _T_76700 = $signed(buffer_12_737) + $signed(buffer_12_689); // @[Modules.scala 78:156:@30747.4]
  assign _T_76701 = _T_76700[10:0]; // @[Modules.scala 78:156:@30748.4]
  assign buffer_12_738 = $signed(_T_76701); // @[Modules.scala 78:156:@30749.4]
  assign _T_76703 = $signed(buffer_12_738) + $signed(buffer_1_690); // @[Modules.scala 78:156:@30751.4]
  assign _T_76704 = _T_76703[10:0]; // @[Modules.scala 78:156:@30752.4]
  assign buffer_12_739 = $signed(_T_76704); // @[Modules.scala 78:156:@30753.4]
  assign _T_76706 = $signed(buffer_12_739) + $signed(buffer_12_691); // @[Modules.scala 78:156:@30755.4]
  assign _T_76707 = _T_76706[10:0]; // @[Modules.scala 78:156:@30756.4]
  assign buffer_12_740 = $signed(_T_76707); // @[Modules.scala 78:156:@30757.4]
  assign _T_76709 = $signed(buffer_12_740) + $signed(buffer_12_692); // @[Modules.scala 78:156:@30759.4]
  assign _T_76710 = _T_76709[10:0]; // @[Modules.scala 78:156:@30760.4]
  assign buffer_12_741 = $signed(_T_76710); // @[Modules.scala 78:156:@30761.4]
  assign _T_76712 = $signed(buffer_12_741) + $signed(buffer_12_693); // @[Modules.scala 78:156:@30763.4]
  assign _T_76713 = _T_76712[10:0]; // @[Modules.scala 78:156:@30764.4]
  assign buffer_12_742 = $signed(_T_76713); // @[Modules.scala 78:156:@30765.4]
  assign _T_76715 = $signed(buffer_12_742) + $signed(buffer_12_694); // @[Modules.scala 78:156:@30767.4]
  assign _T_76716 = _T_76715[10:0]; // @[Modules.scala 78:156:@30768.4]
  assign buffer_12_743 = $signed(_T_76716); // @[Modules.scala 78:156:@30769.4]
  assign _T_76718 = $signed(buffer_12_743) + $signed(buffer_12_695); // @[Modules.scala 78:156:@30771.4]
  assign _T_76719 = _T_76718[10:0]; // @[Modules.scala 78:156:@30772.4]
  assign buffer_12_744 = $signed(_T_76719); // @[Modules.scala 78:156:@30773.4]
  assign _T_76721 = $signed(buffer_12_744) + $signed(buffer_12_696); // @[Modules.scala 78:156:@30775.4]
  assign _T_76722 = _T_76721[10:0]; // @[Modules.scala 78:156:@30776.4]
  assign buffer_12_745 = $signed(_T_76722); // @[Modules.scala 78:156:@30777.4]
  assign _T_76724 = $signed(buffer_12_745) + $signed(buffer_12_697); // @[Modules.scala 78:156:@30779.4]
  assign _T_76725 = _T_76724[10:0]; // @[Modules.scala 78:156:@30780.4]
  assign buffer_12_746 = $signed(_T_76725); // @[Modules.scala 78:156:@30781.4]
  assign _T_76727 = $signed(buffer_12_746) + $signed(buffer_12_698); // @[Modules.scala 78:156:@30783.4]
  assign _T_76728 = _T_76727[10:0]; // @[Modules.scala 78:156:@30784.4]
  assign buffer_12_747 = $signed(_T_76728); // @[Modules.scala 78:156:@30785.4]
  assign _T_76730 = $signed(buffer_12_747) + $signed(buffer_12_699); // @[Modules.scala 78:156:@30787.4]
  assign _T_76731 = _T_76730[10:0]; // @[Modules.scala 78:156:@30788.4]
  assign buffer_12_748 = $signed(_T_76731); // @[Modules.scala 78:156:@30789.4]
  assign _T_76733 = $signed(buffer_12_748) + $signed(buffer_12_700); // @[Modules.scala 78:156:@30791.4]
  assign _T_76734 = _T_76733[10:0]; // @[Modules.scala 78:156:@30792.4]
  assign buffer_12_749 = $signed(_T_76734); // @[Modules.scala 78:156:@30793.4]
  assign _T_76736 = $signed(buffer_12_749) + $signed(buffer_12_701); // @[Modules.scala 78:156:@30795.4]
  assign _T_76737 = _T_76736[10:0]; // @[Modules.scala 78:156:@30796.4]
  assign buffer_12_750 = $signed(_T_76737); // @[Modules.scala 78:156:@30797.4]
  assign _T_76739 = $signed(buffer_12_750) + $signed(buffer_12_702); // @[Modules.scala 78:156:@30799.4]
  assign _T_76740 = _T_76739[10:0]; // @[Modules.scala 78:156:@30800.4]
  assign buffer_12_751 = $signed(_T_76740); // @[Modules.scala 78:156:@30801.4]
  assign _T_76742 = $signed(buffer_12_751) + $signed(buffer_12_703); // @[Modules.scala 78:156:@30803.4]
  assign _T_76743 = _T_76742[10:0]; // @[Modules.scala 78:156:@30804.4]
  assign buffer_12_752 = $signed(_T_76743); // @[Modules.scala 78:156:@30805.4]
  assign _T_76745 = $signed(buffer_12_752) + $signed(buffer_12_704); // @[Modules.scala 78:156:@30807.4]
  assign _T_76746 = _T_76745[10:0]; // @[Modules.scala 78:156:@30808.4]
  assign buffer_12_753 = $signed(_T_76746); // @[Modules.scala 78:156:@30809.4]
  assign _T_76748 = $signed(buffer_12_753) + $signed(buffer_12_705); // @[Modules.scala 78:156:@30811.4]
  assign _T_76749 = _T_76748[10:0]; // @[Modules.scala 78:156:@30812.4]
  assign buffer_12_754 = $signed(_T_76749); // @[Modules.scala 78:156:@30813.4]
  assign _T_76751 = $signed(buffer_12_754) + $signed(buffer_12_706); // @[Modules.scala 78:156:@30815.4]
  assign _T_76752 = _T_76751[10:0]; // @[Modules.scala 78:156:@30816.4]
  assign buffer_12_755 = $signed(_T_76752); // @[Modules.scala 78:156:@30817.4]
  assign _T_76754 = $signed(buffer_12_755) + $signed(buffer_12_707); // @[Modules.scala 78:156:@30819.4]
  assign _T_76755 = _T_76754[10:0]; // @[Modules.scala 78:156:@30820.4]
  assign buffer_12_756 = $signed(_T_76755); // @[Modules.scala 78:156:@30821.4]
  assign _T_76757 = $signed(buffer_12_756) + $signed(buffer_12_708); // @[Modules.scala 78:156:@30823.4]
  assign _T_76758 = _T_76757[10:0]; // @[Modules.scala 78:156:@30824.4]
  assign buffer_12_757 = $signed(_T_76758); // @[Modules.scala 78:156:@30825.4]
  assign _T_76760 = $signed(buffer_12_757) + $signed(buffer_0_701); // @[Modules.scala 78:156:@30827.4]
  assign _T_76761 = _T_76760[10:0]; // @[Modules.scala 78:156:@30828.4]
  assign buffer_12_758 = $signed(_T_76761); // @[Modules.scala 78:156:@30829.4]
  assign _T_76763 = $signed(buffer_12_758) + $signed(buffer_12_710); // @[Modules.scala 78:156:@30831.4]
  assign _T_76764 = _T_76763[10:0]; // @[Modules.scala 78:156:@30832.4]
  assign buffer_12_759 = $signed(_T_76764); // @[Modules.scala 78:156:@30833.4]
  assign _T_76766 = $signed(buffer_12_759) + $signed(buffer_12_711); // @[Modules.scala 78:156:@30835.4]
  assign _T_76767 = _T_76766[10:0]; // @[Modules.scala 78:156:@30836.4]
  assign buffer_12_760 = $signed(_T_76767); // @[Modules.scala 78:156:@30837.4]
  assign _T_76769 = $signed(buffer_12_760) + $signed(buffer_12_712); // @[Modules.scala 78:156:@30839.4]
  assign _T_76770 = _T_76769[10:0]; // @[Modules.scala 78:156:@30840.4]
  assign buffer_12_761 = $signed(_T_76770); // @[Modules.scala 78:156:@30841.4]
  assign _T_76772 = $signed(buffer_12_761) + $signed(buffer_12_713); // @[Modules.scala 78:156:@30843.4]
  assign _T_76773 = _T_76772[10:0]; // @[Modules.scala 78:156:@30844.4]
  assign buffer_12_762 = $signed(_T_76773); // @[Modules.scala 78:156:@30845.4]
  assign _T_76775 = $signed(buffer_12_762) + $signed(buffer_12_714); // @[Modules.scala 78:156:@30847.4]
  assign _T_76776 = _T_76775[10:0]; // @[Modules.scala 78:156:@30848.4]
  assign buffer_12_763 = $signed(_T_76776); // @[Modules.scala 78:156:@30849.4]
  assign _T_76778 = $signed(buffer_12_763) + $signed(buffer_12_715); // @[Modules.scala 78:156:@30851.4]
  assign _T_76779 = _T_76778[10:0]; // @[Modules.scala 78:156:@30852.4]
  assign buffer_12_764 = $signed(_T_76779); // @[Modules.scala 78:156:@30853.4]
  assign _T_76781 = $signed(buffer_12_764) + $signed(buffer_12_716); // @[Modules.scala 78:156:@30855.4]
  assign _T_76782 = _T_76781[10:0]; // @[Modules.scala 78:156:@30856.4]
  assign buffer_12_765 = $signed(_T_76782); // @[Modules.scala 78:156:@30857.4]
  assign _T_76784 = $signed(buffer_12_765) + $signed(buffer_12_717); // @[Modules.scala 78:156:@30859.4]
  assign _T_76785 = _T_76784[10:0]; // @[Modules.scala 78:156:@30860.4]
  assign buffer_12_766 = $signed(_T_76785); // @[Modules.scala 78:156:@30861.4]
  assign _T_76787 = $signed(buffer_12_766) + $signed(buffer_12_718); // @[Modules.scala 78:156:@30863.4]
  assign _T_76788 = _T_76787[10:0]; // @[Modules.scala 78:156:@30864.4]
  assign buffer_12_767 = $signed(_T_76788); // @[Modules.scala 78:156:@30865.4]
  assign _T_76790 = $signed(buffer_12_767) + $signed(buffer_12_719); // @[Modules.scala 78:156:@30867.4]
  assign _T_76791 = _T_76790[10:0]; // @[Modules.scala 78:156:@30868.4]
  assign buffer_12_768 = $signed(_T_76791); // @[Modules.scala 78:156:@30869.4]
  assign _T_76793 = $signed(buffer_12_768) + $signed(buffer_12_720); // @[Modules.scala 78:156:@30871.4]
  assign _T_76794 = _T_76793[10:0]; // @[Modules.scala 78:156:@30872.4]
  assign buffer_12_769 = $signed(_T_76794); // @[Modules.scala 78:156:@30873.4]
  assign _T_76796 = $signed(buffer_12_769) + $signed(buffer_12_721); // @[Modules.scala 78:156:@30875.4]
  assign _T_76797 = _T_76796[10:0]; // @[Modules.scala 78:156:@30876.4]
  assign buffer_12_770 = $signed(_T_76797); // @[Modules.scala 78:156:@30877.4]
  assign _T_76799 = $signed(buffer_12_770) + $signed(buffer_12_722); // @[Modules.scala 78:156:@30879.4]
  assign _T_76800 = _T_76799[10:0]; // @[Modules.scala 78:156:@30880.4]
  assign buffer_12_771 = $signed(_T_76800); // @[Modules.scala 78:156:@30881.4]
  assign _T_76802 = $signed(buffer_12_771) + $signed(buffer_12_723); // @[Modules.scala 78:156:@30883.4]
  assign _T_76803 = _T_76802[10:0]; // @[Modules.scala 78:156:@30884.4]
  assign buffer_12_772 = $signed(_T_76803); // @[Modules.scala 78:156:@30885.4]
  assign _T_76805 = $signed(buffer_12_772) + $signed(buffer_12_724); // @[Modules.scala 78:156:@30887.4]
  assign _T_76806 = _T_76805[10:0]; // @[Modules.scala 78:156:@30888.4]
  assign buffer_12_773 = $signed(_T_76806); // @[Modules.scala 78:156:@30889.4]
  assign _T_76808 = $signed(buffer_12_773) + $signed(buffer_12_725); // @[Modules.scala 78:156:@30891.4]
  assign _T_76809 = _T_76808[10:0]; // @[Modules.scala 78:156:@30892.4]
  assign buffer_12_774 = $signed(_T_76809); // @[Modules.scala 78:156:@30893.4]
  assign _T_76811 = $signed(buffer_12_774) + $signed(buffer_12_726); // @[Modules.scala 78:156:@30895.4]
  assign _T_76812 = _T_76811[10:0]; // @[Modules.scala 78:156:@30896.4]
  assign buffer_12_775 = $signed(_T_76812); // @[Modules.scala 78:156:@30897.4]
  assign _T_76814 = $signed(buffer_12_775) + $signed(buffer_12_727); // @[Modules.scala 78:156:@30899.4]
  assign _T_76815 = _T_76814[10:0]; // @[Modules.scala 78:156:@30900.4]
  assign buffer_12_776 = $signed(_T_76815); // @[Modules.scala 78:156:@30901.4]
  assign _T_76817 = $signed(buffer_12_776) + $signed(buffer_12_728); // @[Modules.scala 78:156:@30903.4]
  assign _T_76818 = _T_76817[10:0]; // @[Modules.scala 78:156:@30904.4]
  assign buffer_12_777 = $signed(_T_76818); // @[Modules.scala 78:156:@30905.4]
  assign _T_76820 = $signed(buffer_12_777) + $signed(buffer_12_729); // @[Modules.scala 78:156:@30907.4]
  assign _T_76821 = _T_76820[10:0]; // @[Modules.scala 78:156:@30908.4]
  assign buffer_12_778 = $signed(_T_76821); // @[Modules.scala 78:156:@30909.4]
  assign _T_76823 = $signed(buffer_12_778) + $signed(buffer_0_701); // @[Modules.scala 78:156:@30911.4]
  assign _T_76824 = _T_76823[10:0]; // @[Modules.scala 78:156:@30912.4]
  assign buffer_12_779 = $signed(_T_76824); // @[Modules.scala 78:156:@30913.4]
  assign _T_76826 = $signed(buffer_12_779) + $signed(buffer_12_731); // @[Modules.scala 78:156:@30915.4]
  assign _T_76827 = _T_76826[10:0]; // @[Modules.scala 78:156:@30916.4]
  assign buffer_12_780 = $signed(_T_76827); // @[Modules.scala 78:156:@30917.4]
  assign _T_76829 = $signed(buffer_12_780) + $signed(buffer_0_701); // @[Modules.scala 78:156:@30919.4]
  assign _T_76830 = _T_76829[10:0]; // @[Modules.scala 78:156:@30920.4]
  assign buffer_12_781 = $signed(_T_76830); // @[Modules.scala 78:156:@30921.4]
  assign _T_76832 = $signed(buffer_12_781) + $signed(buffer_12_733); // @[Modules.scala 78:156:@30923.4]
  assign _T_76833 = _T_76832[10:0]; // @[Modules.scala 78:156:@30924.4]
  assign buffer_12_782 = $signed(_T_76833); // @[Modules.scala 78:156:@30925.4]
  assign _T_76835 = $signed(buffer_12_782) + $signed(buffer_12_734); // @[Modules.scala 78:156:@30927.4]
  assign _T_76836 = _T_76835[10:0]; // @[Modules.scala 78:156:@30928.4]
  assign buffer_12_783 = $signed(_T_76836); // @[Modules.scala 78:156:@30929.4]
  assign _T_77356 = $signed(buffer_7_0) + $signed(buffer_3_1); // @[Modules.scala 65:57:@31693.4]
  assign _T_77357 = _T_77356[10:0]; // @[Modules.scala 65:57:@31694.4]
  assign buffer_13_392 = $signed(_T_77357); // @[Modules.scala 65:57:@31695.4]
  assign buffer_13_6 = {{6{io_in_12[4]}},io_in_12}; // @[Modules.scala 32:22:@8.4]
  assign _T_77365 = $signed(buffer_13_6) + $signed(11'sh0); // @[Modules.scala 65:57:@31705.4]
  assign _T_77366 = _T_77365[10:0]; // @[Modules.scala 65:57:@31706.4]
  assign buffer_13_395 = $signed(_T_77366); // @[Modules.scala 65:57:@31707.4]
  assign _T_77377 = $signed(buffer_4_14) + $signed(buffer_0_15); // @[Modules.scala 65:57:@31721.4]
  assign _T_77378 = _T_77377[10:0]; // @[Modules.scala 65:57:@31722.4]
  assign buffer_13_399 = $signed(_T_77378); // @[Modules.scala 65:57:@31723.4]
  assign buffer_13_18 = {{6{io_in_36[4]}},io_in_36}; // @[Modules.scala 32:22:@8.4]
  assign _T_77383 = $signed(buffer_13_18) + $signed(11'sh0); // @[Modules.scala 65:57:@31729.4]
  assign _T_77384 = _T_77383[10:0]; // @[Modules.scala 65:57:@31730.4]
  assign buffer_13_401 = $signed(_T_77384); // @[Modules.scala 65:57:@31731.4]
  assign _T_77395 = $signed(buffer_1_26) + $signed(11'sh0); // @[Modules.scala 65:57:@31745.4]
  assign _T_77396 = _T_77395[10:0]; // @[Modules.scala 65:57:@31746.4]
  assign buffer_13_405 = $signed(_T_77396); // @[Modules.scala 65:57:@31747.4]
  assign buffer_13_35 = {{6{io_in_70[4]}},io_in_70}; // @[Modules.scala 32:22:@8.4]
  assign _T_77407 = $signed(buffer_1_34) + $signed(buffer_13_35); // @[Modules.scala 65:57:@31761.4]
  assign _T_77408 = _T_77407[10:0]; // @[Modules.scala 65:57:@31762.4]
  assign buffer_13_409 = $signed(_T_77408); // @[Modules.scala 65:57:@31763.4]
  assign _T_77410 = $signed(buffer_5_36) + $signed(buffer_1_37); // @[Modules.scala 65:57:@31765.4]
  assign _T_77411 = _T_77410[10:0]; // @[Modules.scala 65:57:@31766.4]
  assign buffer_13_410 = $signed(_T_77411); // @[Modules.scala 65:57:@31767.4]
  assign buffer_13_40 = {{6{io_in_80[4]}},io_in_80}; // @[Modules.scala 32:22:@8.4]
  assign _T_77416 = $signed(buffer_13_40) + $signed(buffer_0_41); // @[Modules.scala 65:57:@31773.4]
  assign _T_77417 = _T_77416[10:0]; // @[Modules.scala 65:57:@31774.4]
  assign buffer_13_412 = $signed(_T_77417); // @[Modules.scala 65:57:@31775.4]
  assign _T_77428 = $signed(buffer_1_48) + $signed(11'sh0); // @[Modules.scala 65:57:@31789.4]
  assign _T_77429 = _T_77428[10:0]; // @[Modules.scala 65:57:@31790.4]
  assign buffer_13_416 = $signed(_T_77429); // @[Modules.scala 65:57:@31791.4]
  assign _T_77446 = $signed(buffer_8_60) + $signed(buffer_4_61); // @[Modules.scala 65:57:@31813.4]
  assign _T_77447 = _T_77446[10:0]; // @[Modules.scala 65:57:@31814.4]
  assign buffer_13_422 = $signed(_T_77447); // @[Modules.scala 65:57:@31815.4]
  assign buffer_13_79 = {{6{io_in_158[4]}},io_in_158}; // @[Modules.scala 32:22:@8.4]
  assign _T_77473 = $signed(buffer_4_78) + $signed(buffer_13_79); // @[Modules.scala 65:57:@31849.4]
  assign _T_77474 = _T_77473[10:0]; // @[Modules.scala 65:57:@31850.4]
  assign buffer_13_431 = $signed(_T_77474); // @[Modules.scala 65:57:@31851.4]
  assign _T_77476 = $signed(buffer_4_80) + $signed(11'sh0); // @[Modules.scala 65:57:@31853.4]
  assign _T_77477 = _T_77476[10:0]; // @[Modules.scala 65:57:@31854.4]
  assign buffer_13_432 = $signed(_T_77477); // @[Modules.scala 65:57:@31855.4]
  assign buffer_13_85 = {{6{io_in_170[4]}},io_in_170}; // @[Modules.scala 32:22:@8.4]
  assign _T_77482 = $signed(11'sh0) + $signed(buffer_13_85); // @[Modules.scala 65:57:@31861.4]
  assign _T_77483 = _T_77482[10:0]; // @[Modules.scala 65:57:@31862.4]
  assign buffer_13_434 = $signed(_T_77483); // @[Modules.scala 65:57:@31863.4]
  assign buffer_13_90 = {{6{io_in_180[4]}},io_in_180}; // @[Modules.scala 32:22:@8.4]
  assign _T_77491 = $signed(buffer_13_90) + $signed(buffer_9_91); // @[Modules.scala 65:57:@31873.4]
  assign _T_77492 = _T_77491[10:0]; // @[Modules.scala 65:57:@31874.4]
  assign buffer_13_437 = $signed(_T_77492); // @[Modules.scala 65:57:@31875.4]
  assign buffer_13_93 = {{6{io_in_187[4]}},io_in_187}; // @[Modules.scala 32:22:@8.4]
  assign _T_77494 = $signed(buffer_5_92) + $signed(buffer_13_93); // @[Modules.scala 65:57:@31877.4]
  assign _T_77495 = _T_77494[10:0]; // @[Modules.scala 65:57:@31878.4]
  assign buffer_13_438 = $signed(_T_77495); // @[Modules.scala 65:57:@31879.4]
  assign _T_77497 = $signed(buffer_4_94) + $signed(buffer_0_95); // @[Modules.scala 65:57:@31881.4]
  assign _T_77498 = _T_77497[10:0]; // @[Modules.scala 65:57:@31882.4]
  assign buffer_13_439 = $signed(_T_77498); // @[Modules.scala 65:57:@31883.4]
  assign _T_77503 = $signed(11'sh0) + $signed(buffer_0_99); // @[Modules.scala 65:57:@31889.4]
  assign _T_77504 = _T_77503[10:0]; // @[Modules.scala 65:57:@31890.4]
  assign buffer_13_441 = $signed(_T_77504); // @[Modules.scala 65:57:@31891.4]
  assign _T_77506 = $signed(buffer_10_100) + $signed(11'sh0); // @[Modules.scala 65:57:@31893.4]
  assign _T_77507 = _T_77506[10:0]; // @[Modules.scala 65:57:@31894.4]
  assign buffer_13_442 = $signed(_T_77507); // @[Modules.scala 65:57:@31895.4]
  assign _T_77512 = $signed(11'sh0) + $signed(buffer_11_105); // @[Modules.scala 65:57:@31901.4]
  assign _T_77513 = _T_77512[10:0]; // @[Modules.scala 65:57:@31902.4]
  assign buffer_13_444 = $signed(_T_77513); // @[Modules.scala 65:57:@31903.4]
  assign _T_77524 = $signed(11'sh0) + $signed(buffer_12_113); // @[Modules.scala 65:57:@31917.4]
  assign _T_77525 = _T_77524[10:0]; // @[Modules.scala 65:57:@31918.4]
  assign buffer_13_448 = $signed(_T_77525); // @[Modules.scala 65:57:@31919.4]
  assign _T_77527 = $signed(11'sh0) + $signed(buffer_5_115); // @[Modules.scala 65:57:@31921.4]
  assign _T_77528 = _T_77527[10:0]; // @[Modules.scala 65:57:@31922.4]
  assign buffer_13_449 = $signed(_T_77528); // @[Modules.scala 65:57:@31923.4]
  assign buffer_13_120 = {{6{io_in_240[4]}},io_in_240}; // @[Modules.scala 32:22:@8.4]
  assign _T_77536 = $signed(buffer_13_120) + $signed(buffer_4_121); // @[Modules.scala 65:57:@31933.4]
  assign _T_77537 = _T_77536[10:0]; // @[Modules.scala 65:57:@31934.4]
  assign buffer_13_452 = $signed(_T_77537); // @[Modules.scala 65:57:@31935.4]
  assign _T_77551 = $signed(buffer_2_130) + $signed(buffer_0_131); // @[Modules.scala 65:57:@31953.4]
  assign _T_77552 = _T_77551[10:0]; // @[Modules.scala 65:57:@31954.4]
  assign buffer_13_457 = $signed(_T_77552); // @[Modules.scala 65:57:@31955.4]
  assign buffer_13_132 = {{6{io_in_264[4]}},io_in_264}; // @[Modules.scala 32:22:@8.4]
  assign _T_77554 = $signed(buffer_13_132) + $signed(11'sh0); // @[Modules.scala 65:57:@31957.4]
  assign _T_77555 = _T_77554[10:0]; // @[Modules.scala 65:57:@31958.4]
  assign buffer_13_458 = $signed(_T_77555); // @[Modules.scala 65:57:@31959.4]
  assign _T_77560 = $signed(11'sh0) + $signed(buffer_3_137); // @[Modules.scala 65:57:@31965.4]
  assign _T_77561 = _T_77560[10:0]; // @[Modules.scala 65:57:@31966.4]
  assign buffer_13_460 = $signed(_T_77561); // @[Modules.scala 65:57:@31967.4]
  assign buffer_13_145 = {{6{io_in_291[4]}},io_in_291}; // @[Modules.scala 32:22:@8.4]
  assign _T_77572 = $signed(buffer_2_144) + $signed(buffer_13_145); // @[Modules.scala 65:57:@31981.4]
  assign _T_77573 = _T_77572[10:0]; // @[Modules.scala 65:57:@31982.4]
  assign buffer_13_464 = $signed(_T_77573); // @[Modules.scala 65:57:@31983.4]
  assign _T_77578 = $signed(buffer_4_148) + $signed(buffer_3_149); // @[Modules.scala 65:57:@31989.4]
  assign _T_77579 = _T_77578[10:0]; // @[Modules.scala 65:57:@31990.4]
  assign buffer_13_466 = $signed(_T_77579); // @[Modules.scala 65:57:@31991.4]
  assign _T_77581 = $signed(buffer_5_150) + $signed(buffer_4_151); // @[Modules.scala 65:57:@31993.4]
  assign _T_77582 = _T_77581[10:0]; // @[Modules.scala 65:57:@31994.4]
  assign buffer_13_467 = $signed(_T_77582); // @[Modules.scala 65:57:@31995.4]
  assign _T_77590 = $signed(buffer_6_156) + $signed(buffer_1_157); // @[Modules.scala 65:57:@32005.4]
  assign _T_77591 = _T_77590[10:0]; // @[Modules.scala 65:57:@32006.4]
  assign buffer_13_470 = $signed(_T_77591); // @[Modules.scala 65:57:@32007.4]
  assign buffer_13_158 = {{6{io_in_316[4]}},io_in_316}; // @[Modules.scala 32:22:@8.4]
  assign _T_77593 = $signed(buffer_13_158) + $signed(buffer_0_159); // @[Modules.scala 65:57:@32009.4]
  assign _T_77594 = _T_77593[10:0]; // @[Modules.scala 65:57:@32010.4]
  assign buffer_13_471 = $signed(_T_77594); // @[Modules.scala 65:57:@32011.4]
  assign _T_77599 = $signed(11'sh0) + $signed(buffer_5_163); // @[Modules.scala 65:57:@32017.4]
  assign _T_77600 = _T_77599[10:0]; // @[Modules.scala 65:57:@32018.4]
  assign buffer_13_473 = $signed(_T_77600); // @[Modules.scala 65:57:@32019.4]
  assign _T_77608 = $signed(buffer_3_168) + $signed(11'sh0); // @[Modules.scala 65:57:@32029.4]
  assign _T_77609 = _T_77608[10:0]; // @[Modules.scala 65:57:@32030.4]
  assign buffer_13_476 = $signed(_T_77609); // @[Modules.scala 65:57:@32031.4]
  assign buffer_13_171 = {{6{io_in_342[4]}},io_in_342}; // @[Modules.scala 32:22:@8.4]
  assign _T_77611 = $signed(buffer_0_170) + $signed(buffer_13_171); // @[Modules.scala 65:57:@32033.4]
  assign _T_77612 = _T_77611[10:0]; // @[Modules.scala 65:57:@32034.4]
  assign buffer_13_477 = $signed(_T_77612); // @[Modules.scala 65:57:@32035.4]
  assign buffer_13_172 = {{6{io_in_345[4]}},io_in_345}; // @[Modules.scala 32:22:@8.4]
  assign _T_77614 = $signed(buffer_13_172) + $signed(11'sh0); // @[Modules.scala 65:57:@32037.4]
  assign _T_77615 = _T_77614[10:0]; // @[Modules.scala 65:57:@32038.4]
  assign buffer_13_478 = $signed(_T_77615); // @[Modules.scala 65:57:@32039.4]
  assign buffer_13_174 = {{6{io_in_348[4]}},io_in_348}; // @[Modules.scala 32:22:@8.4]
  assign _T_77617 = $signed(buffer_13_174) + $signed(11'sh0); // @[Modules.scala 65:57:@32041.4]
  assign _T_77618 = _T_77617[10:0]; // @[Modules.scala 65:57:@32042.4]
  assign buffer_13_479 = $signed(_T_77618); // @[Modules.scala 65:57:@32043.4]
  assign buffer_13_176 = {{6{io_in_353[4]}},io_in_353}; // @[Modules.scala 32:22:@8.4]
  assign _T_77620 = $signed(buffer_13_176) + $signed(buffer_5_177); // @[Modules.scala 65:57:@32045.4]
  assign _T_77621 = _T_77620[10:0]; // @[Modules.scala 65:57:@32046.4]
  assign buffer_13_480 = $signed(_T_77621); // @[Modules.scala 65:57:@32047.4]
  assign _T_77629 = $signed(buffer_7_182) + $signed(11'sh0); // @[Modules.scala 65:57:@32057.4]
  assign _T_77630 = _T_77629[10:0]; // @[Modules.scala 65:57:@32058.4]
  assign buffer_13_483 = $signed(_T_77630); // @[Modules.scala 65:57:@32059.4]
  assign _T_77635 = $signed(11'sh0) + $signed(buffer_0_187); // @[Modules.scala 65:57:@32065.4]
  assign _T_77636 = _T_77635[10:0]; // @[Modules.scala 65:57:@32066.4]
  assign buffer_13_485 = $signed(_T_77636); // @[Modules.scala 65:57:@32067.4]
  assign _T_77641 = $signed(buffer_4_190) + $signed(buffer_0_191); // @[Modules.scala 65:57:@32073.4]
  assign _T_77642 = _T_77641[10:0]; // @[Modules.scala 65:57:@32074.4]
  assign buffer_13_487 = $signed(_T_77642); // @[Modules.scala 65:57:@32075.4]
  assign _T_77644 = $signed(buffer_2_192) + $signed(buffer_0_193); // @[Modules.scala 65:57:@32077.4]
  assign _T_77645 = _T_77644[10:0]; // @[Modules.scala 65:57:@32078.4]
  assign buffer_13_488 = $signed(_T_77645); // @[Modules.scala 65:57:@32079.4]
  assign _T_77659 = $signed(buffer_1_202) + $signed(buffer_0_203); // @[Modules.scala 65:57:@32097.4]
  assign _T_77660 = _T_77659[10:0]; // @[Modules.scala 65:57:@32098.4]
  assign buffer_13_493 = $signed(_T_77660); // @[Modules.scala 65:57:@32099.4]
  assign _T_77662 = $signed(buffer_8_204) + $signed(11'sh0); // @[Modules.scala 65:57:@32101.4]
  assign _T_77663 = _T_77662[10:0]; // @[Modules.scala 65:57:@32102.4]
  assign buffer_13_494 = $signed(_T_77663); // @[Modules.scala 65:57:@32103.4]
  assign _T_77701 = $signed(buffer_2_230) + $signed(11'sh0); // @[Modules.scala 65:57:@32153.4]
  assign _T_77702 = _T_77701[10:0]; // @[Modules.scala 65:57:@32154.4]
  assign buffer_13_507 = $signed(_T_77702); // @[Modules.scala 65:57:@32155.4]
  assign _T_77704 = $signed(buffer_5_232) + $signed(buffer_1_233); // @[Modules.scala 65:57:@32157.4]
  assign _T_77705 = _T_77704[10:0]; // @[Modules.scala 65:57:@32158.4]
  assign buffer_13_508 = $signed(_T_77705); // @[Modules.scala 65:57:@32159.4]
  assign _T_77707 = $signed(buffer_0_234) + $signed(buffer_11_235); // @[Modules.scala 65:57:@32161.4]
  assign _T_77708 = _T_77707[10:0]; // @[Modules.scala 65:57:@32162.4]
  assign buffer_13_509 = $signed(_T_77708); // @[Modules.scala 65:57:@32163.4]
  assign _T_77716 = $signed(buffer_11_240) + $signed(buffer_0_241); // @[Modules.scala 65:57:@32173.4]
  assign _T_77717 = _T_77716[10:0]; // @[Modules.scala 65:57:@32174.4]
  assign buffer_13_512 = $signed(_T_77717); // @[Modules.scala 65:57:@32175.4]
  assign _T_77725 = $signed(11'sh0) + $signed(buffer_0_247); // @[Modules.scala 65:57:@32185.4]
  assign _T_77726 = _T_77725[10:0]; // @[Modules.scala 65:57:@32186.4]
  assign buffer_13_515 = $signed(_T_77726); // @[Modules.scala 65:57:@32187.4]
  assign buffer_13_248 = {{6{io_in_496[4]}},io_in_496}; // @[Modules.scala 32:22:@8.4]
  assign _T_77728 = $signed(buffer_13_248) + $signed(buffer_11_249); // @[Modules.scala 65:57:@32189.4]
  assign _T_77729 = _T_77728[10:0]; // @[Modules.scala 65:57:@32190.4]
  assign buffer_13_516 = $signed(_T_77729); // @[Modules.scala 65:57:@32191.4]
  assign _T_77746 = $signed(buffer_4_260) + $signed(buffer_0_261); // @[Modules.scala 65:57:@32213.4]
  assign _T_77747 = _T_77746[10:0]; // @[Modules.scala 65:57:@32214.4]
  assign buffer_13_522 = $signed(_T_77747); // @[Modules.scala 65:57:@32215.4]
  assign _T_77749 = $signed(11'sh0) + $signed(buffer_0_263); // @[Modules.scala 65:57:@32217.4]
  assign _T_77750 = _T_77749[10:0]; // @[Modules.scala 65:57:@32218.4]
  assign buffer_13_523 = $signed(_T_77750); // @[Modules.scala 65:57:@32219.4]
  assign buffer_13_265 = {{6{io_in_530[4]}},io_in_530}; // @[Modules.scala 32:22:@8.4]
  assign _T_77752 = $signed(buffer_0_264) + $signed(buffer_13_265); // @[Modules.scala 65:57:@32221.4]
  assign _T_77753 = _T_77752[10:0]; // @[Modules.scala 65:57:@32222.4]
  assign buffer_13_524 = $signed(_T_77753); // @[Modules.scala 65:57:@32223.4]
  assign _T_77758 = $signed(11'sh0) + $signed(buffer_5_269); // @[Modules.scala 65:57:@32229.4]
  assign _T_77759 = _T_77758[10:0]; // @[Modules.scala 65:57:@32230.4]
  assign buffer_13_526 = $signed(_T_77759); // @[Modules.scala 65:57:@32231.4]
  assign _T_77764 = $signed(buffer_4_272) + $signed(buffer_1_273); // @[Modules.scala 65:57:@32237.4]
  assign _T_77765 = _T_77764[10:0]; // @[Modules.scala 65:57:@32238.4]
  assign buffer_13_528 = $signed(_T_77765); // @[Modules.scala 65:57:@32239.4]
  assign _T_77776 = $signed(buffer_1_280) + $signed(11'sh0); // @[Modules.scala 65:57:@32253.4]
  assign _T_77777 = _T_77776[10:0]; // @[Modules.scala 65:57:@32254.4]
  assign buffer_13_532 = $signed(_T_77777); // @[Modules.scala 65:57:@32255.4]
  assign buffer_13_282 = {{6{io_in_565[4]}},io_in_565}; // @[Modules.scala 32:22:@8.4]
  assign _T_77779 = $signed(buffer_13_282) + $signed(buffer_9_283); // @[Modules.scala 65:57:@32257.4]
  assign _T_77780 = _T_77779[10:0]; // @[Modules.scala 65:57:@32258.4]
  assign buffer_13_533 = $signed(_T_77780); // @[Modules.scala 65:57:@32259.4]
  assign _T_77791 = $signed(buffer_5_290) + $signed(buffer_3_291); // @[Modules.scala 65:57:@32273.4]
  assign _T_77792 = _T_77791[10:0]; // @[Modules.scala 65:57:@32274.4]
  assign buffer_13_537 = $signed(_T_77792); // @[Modules.scala 65:57:@32275.4]
  assign _T_77794 = $signed(buffer_0_292) + $signed(11'sh0); // @[Modules.scala 65:57:@32277.4]
  assign _T_77795 = _T_77794[10:0]; // @[Modules.scala 65:57:@32278.4]
  assign buffer_13_538 = $signed(_T_77795); // @[Modules.scala 65:57:@32279.4]
  assign _T_77800 = $signed(buffer_12_296) + $signed(11'sh0); // @[Modules.scala 65:57:@32285.4]
  assign _T_77801 = _T_77800[10:0]; // @[Modules.scala 65:57:@32286.4]
  assign buffer_13_540 = $signed(_T_77801); // @[Modules.scala 65:57:@32287.4]
  assign buffer_13_309 = {{6{io_in_618[4]}},io_in_618}; // @[Modules.scala 32:22:@8.4]
  assign _T_77818 = $signed(buffer_2_308) + $signed(buffer_13_309); // @[Modules.scala 65:57:@32309.4]
  assign _T_77819 = _T_77818[10:0]; // @[Modules.scala 65:57:@32310.4]
  assign buffer_13_546 = $signed(_T_77819); // @[Modules.scala 65:57:@32311.4]
  assign _T_77821 = $signed(11'sh0) + $signed(buffer_4_311); // @[Modules.scala 65:57:@32313.4]
  assign _T_77822 = _T_77821[10:0]; // @[Modules.scala 65:57:@32314.4]
  assign buffer_13_547 = $signed(_T_77822); // @[Modules.scala 65:57:@32315.4]
  assign _T_77824 = $signed(buffer_2_312) + $signed(buffer_3_313); // @[Modules.scala 65:57:@32317.4]
  assign _T_77825 = _T_77824[10:0]; // @[Modules.scala 65:57:@32318.4]
  assign buffer_13_548 = $signed(_T_77825); // @[Modules.scala 65:57:@32319.4]
  assign _T_77827 = $signed(buffer_1_314) + $signed(11'sh0); // @[Modules.scala 65:57:@32321.4]
  assign _T_77828 = _T_77827[10:0]; // @[Modules.scala 65:57:@32322.4]
  assign buffer_13_549 = $signed(_T_77828); // @[Modules.scala 65:57:@32323.4]
  assign _T_77830 = $signed(buffer_3_316) + $signed(buffer_1_317); // @[Modules.scala 65:57:@32325.4]
  assign _T_77831 = _T_77830[10:0]; // @[Modules.scala 65:57:@32326.4]
  assign buffer_13_550 = $signed(_T_77831); // @[Modules.scala 65:57:@32327.4]
  assign _T_77836 = $signed(buffer_0_320) + $signed(11'sh0); // @[Modules.scala 65:57:@32333.4]
  assign _T_77837 = _T_77836[10:0]; // @[Modules.scala 65:57:@32334.4]
  assign buffer_13_552 = $signed(_T_77837); // @[Modules.scala 65:57:@32335.4]
  assign buffer_13_329 = {{6{io_in_659[4]}},io_in_659}; // @[Modules.scala 32:22:@8.4]
  assign _T_77848 = $signed(buffer_1_328) + $signed(buffer_13_329); // @[Modules.scala 65:57:@32349.4]
  assign _T_77849 = _T_77848[10:0]; // @[Modules.scala 65:57:@32350.4]
  assign buffer_13_556 = $signed(_T_77849); // @[Modules.scala 65:57:@32351.4]
  assign _T_77860 = $signed(buffer_3_336) + $signed(11'sh0); // @[Modules.scala 65:57:@32365.4]
  assign _T_77861 = _T_77860[10:0]; // @[Modules.scala 65:57:@32366.4]
  assign buffer_13_560 = $signed(_T_77861); // @[Modules.scala 65:57:@32367.4]
  assign _T_77869 = $signed(11'sh0) + $signed(buffer_3_343); // @[Modules.scala 65:57:@32377.4]
  assign _T_77870 = _T_77869[10:0]; // @[Modules.scala 65:57:@32378.4]
  assign buffer_13_563 = $signed(_T_77870); // @[Modules.scala 65:57:@32379.4]
  assign _T_77881 = $signed(buffer_1_350) + $signed(buffer_0_351); // @[Modules.scala 65:57:@32393.4]
  assign _T_77882 = _T_77881[10:0]; // @[Modules.scala 65:57:@32394.4]
  assign buffer_13_567 = $signed(_T_77882); // @[Modules.scala 65:57:@32395.4]
  assign _T_77902 = $signed(11'sh0) + $signed(buffer_2_365); // @[Modules.scala 65:57:@32421.4]
  assign _T_77903 = _T_77902[10:0]; // @[Modules.scala 65:57:@32422.4]
  assign buffer_13_574 = $signed(_T_77903); // @[Modules.scala 65:57:@32423.4]
  assign _T_77923 = $signed(11'sh0) + $signed(buffer_8_379); // @[Modules.scala 65:57:@32449.4]
  assign _T_77924 = _T_77923[10:0]; // @[Modules.scala 65:57:@32450.4]
  assign buffer_13_581 = $signed(_T_77924); // @[Modules.scala 65:57:@32451.4]
  assign buffer_13_391 = {{6{io_in_782[4]}},io_in_782}; // @[Modules.scala 32:22:@8.4]
  assign _T_77941 = $signed(11'sh0) + $signed(buffer_13_391); // @[Modules.scala 65:57:@32473.4]
  assign _T_77942 = _T_77941[10:0]; // @[Modules.scala 65:57:@32474.4]
  assign buffer_13_587 = $signed(_T_77942); // @[Modules.scala 65:57:@32475.4]
  assign _T_77944 = $signed(buffer_13_392) + $signed(buffer_0_393); // @[Modules.scala 68:83:@32477.4]
  assign _T_77945 = _T_77944[10:0]; // @[Modules.scala 68:83:@32478.4]
  assign buffer_13_588 = $signed(_T_77945); // @[Modules.scala 68:83:@32479.4]
  assign _T_77947 = $signed(buffer_4_394) + $signed(buffer_13_395); // @[Modules.scala 68:83:@32481.4]
  assign _T_77948 = _T_77947[10:0]; // @[Modules.scala 68:83:@32482.4]
  assign buffer_13_589 = $signed(_T_77948); // @[Modules.scala 68:83:@32483.4]
  assign _T_77950 = $signed(buffer_2_396) + $signed(buffer_3_397); // @[Modules.scala 68:83:@32485.4]
  assign _T_77951 = _T_77950[10:0]; // @[Modules.scala 68:83:@32486.4]
  assign buffer_13_590 = $signed(_T_77951); // @[Modules.scala 68:83:@32487.4]
  assign _T_77953 = $signed(buffer_0_395) + $signed(buffer_13_399); // @[Modules.scala 68:83:@32489.4]
  assign _T_77954 = _T_77953[10:0]; // @[Modules.scala 68:83:@32490.4]
  assign buffer_13_591 = $signed(_T_77954); // @[Modules.scala 68:83:@32491.4]
  assign _T_77956 = $signed(buffer_1_400) + $signed(buffer_13_401); // @[Modules.scala 68:83:@32493.4]
  assign _T_77957 = _T_77956[10:0]; // @[Modules.scala 68:83:@32494.4]
  assign buffer_13_592 = $signed(_T_77957); // @[Modules.scala 68:83:@32495.4]
  assign _T_77959 = $signed(buffer_4_402) + $signed(buffer_3_403); // @[Modules.scala 68:83:@32497.4]
  assign _T_77960 = _T_77959[10:0]; // @[Modules.scala 68:83:@32498.4]
  assign buffer_13_593 = $signed(_T_77960); // @[Modules.scala 68:83:@32499.4]
  assign _T_77962 = $signed(buffer_0_395) + $signed(buffer_13_405); // @[Modules.scala 68:83:@32501.4]
  assign _T_77963 = _T_77962[10:0]; // @[Modules.scala 68:83:@32502.4]
  assign buffer_13_594 = $signed(_T_77963); // @[Modules.scala 68:83:@32503.4]
  assign _T_77965 = $signed(buffer_1_406) + $signed(buffer_10_407); // @[Modules.scala 68:83:@32505.4]
  assign _T_77966 = _T_77965[10:0]; // @[Modules.scala 68:83:@32506.4]
  assign buffer_13_595 = $signed(_T_77966); // @[Modules.scala 68:83:@32507.4]
  assign _T_77968 = $signed(buffer_1_408) + $signed(buffer_13_409); // @[Modules.scala 68:83:@32509.4]
  assign _T_77969 = _T_77968[10:0]; // @[Modules.scala 68:83:@32510.4]
  assign buffer_13_596 = $signed(_T_77969); // @[Modules.scala 68:83:@32511.4]
  assign _T_77971 = $signed(buffer_13_410) + $signed(buffer_1_411); // @[Modules.scala 68:83:@32513.4]
  assign _T_77972 = _T_77971[10:0]; // @[Modules.scala 68:83:@32514.4]
  assign buffer_13_597 = $signed(_T_77972); // @[Modules.scala 68:83:@32515.4]
  assign _T_77974 = $signed(buffer_13_412) + $signed(buffer_5_413); // @[Modules.scala 68:83:@32517.4]
  assign _T_77975 = _T_77974[10:0]; // @[Modules.scala 68:83:@32518.4]
  assign buffer_13_598 = $signed(_T_77975); // @[Modules.scala 68:83:@32519.4]
  assign _T_77980 = $signed(buffer_13_416) + $signed(buffer_0_417); // @[Modules.scala 68:83:@32525.4]
  assign _T_77981 = _T_77980[10:0]; // @[Modules.scala 68:83:@32526.4]
  assign buffer_13_600 = $signed(_T_77981); // @[Modules.scala 68:83:@32527.4]
  assign _T_77986 = $signed(buffer_0_420) + $signed(buffer_4_421); // @[Modules.scala 68:83:@32533.4]
  assign _T_77987 = _T_77986[10:0]; // @[Modules.scala 68:83:@32534.4]
  assign buffer_13_602 = $signed(_T_77987); // @[Modules.scala 68:83:@32535.4]
  assign _T_77989 = $signed(buffer_13_422) + $signed(buffer_12_423); // @[Modules.scala 68:83:@32537.4]
  assign _T_77990 = _T_77989[10:0]; // @[Modules.scala 68:83:@32538.4]
  assign buffer_13_603 = $signed(_T_77990); // @[Modules.scala 68:83:@32539.4]
  assign _T_77995 = $signed(buffer_10_426) + $signed(buffer_4_427); // @[Modules.scala 68:83:@32545.4]
  assign _T_77996 = _T_77995[10:0]; // @[Modules.scala 68:83:@32546.4]
  assign buffer_13_605 = $signed(_T_77996); // @[Modules.scala 68:83:@32547.4]
  assign _T_77998 = $signed(buffer_7_428) + $signed(buffer_3_429); // @[Modules.scala 68:83:@32549.4]
  assign _T_77999 = _T_77998[10:0]; // @[Modules.scala 68:83:@32550.4]
  assign buffer_13_606 = $signed(_T_77999); // @[Modules.scala 68:83:@32551.4]
  assign _T_78001 = $signed(buffer_4_430) + $signed(buffer_13_431); // @[Modules.scala 68:83:@32553.4]
  assign _T_78002 = _T_78001[10:0]; // @[Modules.scala 68:83:@32554.4]
  assign buffer_13_607 = $signed(_T_78002); // @[Modules.scala 68:83:@32555.4]
  assign _T_78004 = $signed(buffer_13_432) + $signed(buffer_12_433); // @[Modules.scala 68:83:@32557.4]
  assign _T_78005 = _T_78004[10:0]; // @[Modules.scala 68:83:@32558.4]
  assign buffer_13_608 = $signed(_T_78005); // @[Modules.scala 68:83:@32559.4]
  assign _T_78007 = $signed(buffer_13_434) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32561.4]
  assign _T_78008 = _T_78007[10:0]; // @[Modules.scala 68:83:@32562.4]
  assign buffer_13_609 = $signed(_T_78008); // @[Modules.scala 68:83:@32563.4]
  assign _T_78010 = $signed(buffer_0_395) + $signed(buffer_13_437); // @[Modules.scala 68:83:@32565.4]
  assign _T_78011 = _T_78010[10:0]; // @[Modules.scala 68:83:@32566.4]
  assign buffer_13_610 = $signed(_T_78011); // @[Modules.scala 68:83:@32567.4]
  assign _T_78013 = $signed(buffer_13_438) + $signed(buffer_13_439); // @[Modules.scala 68:83:@32569.4]
  assign _T_78014 = _T_78013[10:0]; // @[Modules.scala 68:83:@32570.4]
  assign buffer_13_611 = $signed(_T_78014); // @[Modules.scala 68:83:@32571.4]
  assign _T_78016 = $signed(buffer_0_395) + $signed(buffer_13_441); // @[Modules.scala 68:83:@32573.4]
  assign _T_78017 = _T_78016[10:0]; // @[Modules.scala 68:83:@32574.4]
  assign buffer_13_612 = $signed(_T_78017); // @[Modules.scala 68:83:@32575.4]
  assign _T_78019 = $signed(buffer_13_442) + $signed(buffer_9_443); // @[Modules.scala 68:83:@32577.4]
  assign _T_78020 = _T_78019[10:0]; // @[Modules.scala 68:83:@32578.4]
  assign buffer_13_613 = $signed(_T_78020); // @[Modules.scala 68:83:@32579.4]
  assign _T_78022 = $signed(buffer_13_444) + $signed(buffer_11_445); // @[Modules.scala 68:83:@32581.4]
  assign _T_78023 = _T_78022[10:0]; // @[Modules.scala 68:83:@32582.4]
  assign buffer_13_614 = $signed(_T_78023); // @[Modules.scala 68:83:@32583.4]
  assign _T_78025 = $signed(buffer_3_446) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32585.4]
  assign _T_78026 = _T_78025[10:0]; // @[Modules.scala 68:83:@32586.4]
  assign buffer_13_615 = $signed(_T_78026); // @[Modules.scala 68:83:@32587.4]
  assign _T_78028 = $signed(buffer_13_448) + $signed(buffer_13_449); // @[Modules.scala 68:83:@32589.4]
  assign _T_78029 = _T_78028[10:0]; // @[Modules.scala 68:83:@32590.4]
  assign buffer_13_616 = $signed(_T_78029); // @[Modules.scala 68:83:@32591.4]
  assign _T_78031 = $signed(buffer_4_450) + $signed(buffer_0_451); // @[Modules.scala 68:83:@32593.4]
  assign _T_78032 = _T_78031[10:0]; // @[Modules.scala 68:83:@32594.4]
  assign buffer_13_617 = $signed(_T_78032); // @[Modules.scala 68:83:@32595.4]
  assign _T_78034 = $signed(buffer_13_452) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32597.4]
  assign _T_78035 = _T_78034[10:0]; // @[Modules.scala 68:83:@32598.4]
  assign buffer_13_618 = $signed(_T_78035); // @[Modules.scala 68:83:@32599.4]
  assign _T_78040 = $signed(buffer_0_395) + $signed(buffer_13_457); // @[Modules.scala 68:83:@32605.4]
  assign _T_78041 = _T_78040[10:0]; // @[Modules.scala 68:83:@32606.4]
  assign buffer_13_620 = $signed(_T_78041); // @[Modules.scala 68:83:@32607.4]
  assign _T_78043 = $signed(buffer_13_458) + $signed(buffer_7_459); // @[Modules.scala 68:83:@32609.4]
  assign _T_78044 = _T_78043[10:0]; // @[Modules.scala 68:83:@32610.4]
  assign buffer_13_621 = $signed(_T_78044); // @[Modules.scala 68:83:@32611.4]
  assign _T_78046 = $signed(buffer_13_460) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32613.4]
  assign _T_78047 = _T_78046[10:0]; // @[Modules.scala 68:83:@32614.4]
  assign buffer_13_622 = $signed(_T_78047); // @[Modules.scala 68:83:@32615.4]
  assign _T_78049 = $signed(buffer_0_395) + $signed(buffer_11_463); // @[Modules.scala 68:83:@32617.4]
  assign _T_78050 = _T_78049[10:0]; // @[Modules.scala 68:83:@32618.4]
  assign buffer_13_623 = $signed(_T_78050); // @[Modules.scala 68:83:@32619.4]
  assign _T_78052 = $signed(buffer_13_464) + $signed(buffer_7_465); // @[Modules.scala 68:83:@32621.4]
  assign _T_78053 = _T_78052[10:0]; // @[Modules.scala 68:83:@32622.4]
  assign buffer_13_624 = $signed(_T_78053); // @[Modules.scala 68:83:@32623.4]
  assign _T_78055 = $signed(buffer_13_466) + $signed(buffer_13_467); // @[Modules.scala 68:83:@32625.4]
  assign _T_78056 = _T_78055[10:0]; // @[Modules.scala 68:83:@32626.4]
  assign buffer_13_625 = $signed(_T_78056); // @[Modules.scala 68:83:@32627.4]
  assign _T_78061 = $signed(buffer_13_470) + $signed(buffer_13_471); // @[Modules.scala 68:83:@32633.4]
  assign _T_78062 = _T_78061[10:0]; // @[Modules.scala 68:83:@32634.4]
  assign buffer_13_627 = $signed(_T_78062); // @[Modules.scala 68:83:@32635.4]
  assign _T_78064 = $signed(buffer_4_472) + $signed(buffer_13_473); // @[Modules.scala 68:83:@32637.4]
  assign _T_78065 = _T_78064[10:0]; // @[Modules.scala 68:83:@32638.4]
  assign buffer_13_628 = $signed(_T_78065); // @[Modules.scala 68:83:@32639.4]
  assign _T_78067 = $signed(buffer_5_474) + $signed(buffer_12_475); // @[Modules.scala 68:83:@32641.4]
  assign _T_78068 = _T_78067[10:0]; // @[Modules.scala 68:83:@32642.4]
  assign buffer_13_629 = $signed(_T_78068); // @[Modules.scala 68:83:@32643.4]
  assign _T_78070 = $signed(buffer_13_476) + $signed(buffer_13_477); // @[Modules.scala 68:83:@32645.4]
  assign _T_78071 = _T_78070[10:0]; // @[Modules.scala 68:83:@32646.4]
  assign buffer_13_630 = $signed(_T_78071); // @[Modules.scala 68:83:@32647.4]
  assign _T_78073 = $signed(buffer_13_478) + $signed(buffer_13_479); // @[Modules.scala 68:83:@32649.4]
  assign _T_78074 = _T_78073[10:0]; // @[Modules.scala 68:83:@32650.4]
  assign buffer_13_631 = $signed(_T_78074); // @[Modules.scala 68:83:@32651.4]
  assign _T_78076 = $signed(buffer_13_480) + $signed(buffer_0_481); // @[Modules.scala 68:83:@32653.4]
  assign _T_78077 = _T_78076[10:0]; // @[Modules.scala 68:83:@32654.4]
  assign buffer_13_632 = $signed(_T_78077); // @[Modules.scala 68:83:@32655.4]
  assign _T_78079 = $signed(buffer_4_482) + $signed(buffer_13_483); // @[Modules.scala 68:83:@32657.4]
  assign _T_78080 = _T_78079[10:0]; // @[Modules.scala 68:83:@32658.4]
  assign buffer_13_633 = $signed(_T_78080); // @[Modules.scala 68:83:@32659.4]
  assign _T_78082 = $signed(buffer_11_484) + $signed(buffer_13_485); // @[Modules.scala 68:83:@32661.4]
  assign _T_78083 = _T_78082[10:0]; // @[Modules.scala 68:83:@32662.4]
  assign buffer_13_634 = $signed(_T_78083); // @[Modules.scala 68:83:@32663.4]
  assign _T_78085 = $signed(buffer_0_395) + $signed(buffer_13_487); // @[Modules.scala 68:83:@32665.4]
  assign _T_78086 = _T_78085[10:0]; // @[Modules.scala 68:83:@32666.4]
  assign buffer_13_635 = $signed(_T_78086); // @[Modules.scala 68:83:@32667.4]
  assign _T_78088 = $signed(buffer_13_488) + $signed(buffer_9_489); // @[Modules.scala 68:83:@32669.4]
  assign _T_78089 = _T_78088[10:0]; // @[Modules.scala 68:83:@32670.4]
  assign buffer_13_636 = $signed(_T_78089); // @[Modules.scala 68:83:@32671.4]
  assign _T_78091 = $signed(buffer_12_490) + $signed(buffer_1_491); // @[Modules.scala 68:83:@32673.4]
  assign _T_78092 = _T_78091[10:0]; // @[Modules.scala 68:83:@32674.4]
  assign buffer_13_637 = $signed(_T_78092); // @[Modules.scala 68:83:@32675.4]
  assign _T_78094 = $signed(buffer_0_492) + $signed(buffer_13_493); // @[Modules.scala 68:83:@32677.4]
  assign _T_78095 = _T_78094[10:0]; // @[Modules.scala 68:83:@32678.4]
  assign buffer_13_638 = $signed(_T_78095); // @[Modules.scala 68:83:@32679.4]
  assign _T_78097 = $signed(buffer_13_494) + $signed(buffer_0_495); // @[Modules.scala 68:83:@32681.4]
  assign _T_78098 = _T_78097[10:0]; // @[Modules.scala 68:83:@32682.4]
  assign buffer_13_639 = $signed(_T_78098); // @[Modules.scala 68:83:@32683.4]
  assign _T_78100 = $signed(buffer_10_496) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32685.4]
  assign _T_78101 = _T_78100[10:0]; // @[Modules.scala 68:83:@32686.4]
  assign buffer_13_640 = $signed(_T_78101); // @[Modules.scala 68:83:@32687.4]
  assign _T_78103 = $signed(buffer_7_498) + $signed(buffer_0_499); // @[Modules.scala 68:83:@32689.4]
  assign _T_78104 = _T_78103[10:0]; // @[Modules.scala 68:83:@32690.4]
  assign buffer_13_641 = $signed(_T_78104); // @[Modules.scala 68:83:@32691.4]
  assign _T_78106 = $signed(buffer_11_500) + $signed(buffer_5_501); // @[Modules.scala 68:83:@32693.4]
  assign _T_78107 = _T_78106[10:0]; // @[Modules.scala 68:83:@32694.4]
  assign buffer_13_642 = $signed(_T_78107); // @[Modules.scala 68:83:@32695.4]
  assign _T_78109 = $signed(buffer_2_502) + $signed(buffer_3_503); // @[Modules.scala 68:83:@32697.4]
  assign _T_78110 = _T_78109[10:0]; // @[Modules.scala 68:83:@32698.4]
  assign buffer_13_643 = $signed(_T_78110); // @[Modules.scala 68:83:@32699.4]
  assign _T_78112 = $signed(buffer_0_395) + $signed(buffer_0_505); // @[Modules.scala 68:83:@32701.4]
  assign _T_78113 = _T_78112[10:0]; // @[Modules.scala 68:83:@32702.4]
  assign buffer_13_644 = $signed(_T_78113); // @[Modules.scala 68:83:@32703.4]
  assign _T_78115 = $signed(buffer_0_506) + $signed(buffer_13_507); // @[Modules.scala 68:83:@32705.4]
  assign _T_78116 = _T_78115[10:0]; // @[Modules.scala 68:83:@32706.4]
  assign buffer_13_645 = $signed(_T_78116); // @[Modules.scala 68:83:@32707.4]
  assign _T_78118 = $signed(buffer_13_508) + $signed(buffer_13_509); // @[Modules.scala 68:83:@32709.4]
  assign _T_78119 = _T_78118[10:0]; // @[Modules.scala 68:83:@32710.4]
  assign buffer_13_646 = $signed(_T_78119); // @[Modules.scala 68:83:@32711.4]
  assign _T_78124 = $signed(buffer_13_512) + $signed(buffer_0_513); // @[Modules.scala 68:83:@32717.4]
  assign _T_78125 = _T_78124[10:0]; // @[Modules.scala 68:83:@32718.4]
  assign buffer_13_648 = $signed(_T_78125); // @[Modules.scala 68:83:@32719.4]
  assign _T_78127 = $signed(buffer_2_514) + $signed(buffer_13_515); // @[Modules.scala 68:83:@32721.4]
  assign _T_78128 = _T_78127[10:0]; // @[Modules.scala 68:83:@32722.4]
  assign buffer_13_649 = $signed(_T_78128); // @[Modules.scala 68:83:@32723.4]
  assign _T_78130 = $signed(buffer_13_516) + $signed(buffer_3_517); // @[Modules.scala 68:83:@32725.4]
  assign _T_78131 = _T_78130[10:0]; // @[Modules.scala 68:83:@32726.4]
  assign buffer_13_650 = $signed(_T_78131); // @[Modules.scala 68:83:@32727.4]
  assign _T_78139 = $signed(buffer_13_522) + $signed(buffer_13_523); // @[Modules.scala 68:83:@32737.4]
  assign _T_78140 = _T_78139[10:0]; // @[Modules.scala 68:83:@32738.4]
  assign buffer_13_653 = $signed(_T_78140); // @[Modules.scala 68:83:@32739.4]
  assign _T_78142 = $signed(buffer_13_524) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32741.4]
  assign _T_78143 = _T_78142[10:0]; // @[Modules.scala 68:83:@32742.4]
  assign buffer_13_654 = $signed(_T_78143); // @[Modules.scala 68:83:@32743.4]
  assign _T_78145 = $signed(buffer_13_526) + $signed(buffer_1_527); // @[Modules.scala 68:83:@32745.4]
  assign _T_78146 = _T_78145[10:0]; // @[Modules.scala 68:83:@32746.4]
  assign buffer_13_655 = $signed(_T_78146); // @[Modules.scala 68:83:@32747.4]
  assign _T_78148 = $signed(buffer_13_528) + $signed(buffer_7_529); // @[Modules.scala 68:83:@32749.4]
  assign _T_78149 = _T_78148[10:0]; // @[Modules.scala 68:83:@32750.4]
  assign buffer_13_656 = $signed(_T_78149); // @[Modules.scala 68:83:@32751.4]
  assign _T_78154 = $signed(buffer_13_532) + $signed(buffer_13_533); // @[Modules.scala 68:83:@32757.4]
  assign _T_78155 = _T_78154[10:0]; // @[Modules.scala 68:83:@32758.4]
  assign buffer_13_658 = $signed(_T_78155); // @[Modules.scala 68:83:@32759.4]
  assign _T_78160 = $signed(buffer_5_536) + $signed(buffer_13_537); // @[Modules.scala 68:83:@32765.4]
  assign _T_78161 = _T_78160[10:0]; // @[Modules.scala 68:83:@32766.4]
  assign buffer_13_660 = $signed(_T_78161); // @[Modules.scala 68:83:@32767.4]
  assign _T_78163 = $signed(buffer_13_538) + $signed(buffer_6_539); // @[Modules.scala 68:83:@32769.4]
  assign _T_78164 = _T_78163[10:0]; // @[Modules.scala 68:83:@32770.4]
  assign buffer_13_661 = $signed(_T_78164); // @[Modules.scala 68:83:@32771.4]
  assign _T_78166 = $signed(buffer_13_540) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32773.4]
  assign _T_78167 = _T_78166[10:0]; // @[Modules.scala 68:83:@32774.4]
  assign buffer_13_662 = $signed(_T_78167); // @[Modules.scala 68:83:@32775.4]
  assign _T_78175 = $signed(buffer_13_546) + $signed(buffer_13_547); // @[Modules.scala 68:83:@32785.4]
  assign _T_78176 = _T_78175[10:0]; // @[Modules.scala 68:83:@32786.4]
  assign buffer_13_665 = $signed(_T_78176); // @[Modules.scala 68:83:@32787.4]
  assign _T_78178 = $signed(buffer_13_548) + $signed(buffer_13_549); // @[Modules.scala 68:83:@32789.4]
  assign _T_78179 = _T_78178[10:0]; // @[Modules.scala 68:83:@32790.4]
  assign buffer_13_666 = $signed(_T_78179); // @[Modules.scala 68:83:@32791.4]
  assign _T_78181 = $signed(buffer_13_550) + $signed(buffer_3_551); // @[Modules.scala 68:83:@32793.4]
  assign _T_78182 = _T_78181[10:0]; // @[Modules.scala 68:83:@32794.4]
  assign buffer_13_667 = $signed(_T_78182); // @[Modules.scala 68:83:@32795.4]
  assign _T_78184 = $signed(buffer_13_552) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32797.4]
  assign _T_78185 = _T_78184[10:0]; // @[Modules.scala 68:83:@32798.4]
  assign buffer_13_668 = $signed(_T_78185); // @[Modules.scala 68:83:@32799.4]
  assign _T_78190 = $signed(buffer_13_556) + $signed(buffer_1_557); // @[Modules.scala 68:83:@32805.4]
  assign _T_78191 = _T_78190[10:0]; // @[Modules.scala 68:83:@32806.4]
  assign buffer_13_670 = $signed(_T_78191); // @[Modules.scala 68:83:@32807.4]
  assign _T_78196 = $signed(buffer_13_560) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32813.4]
  assign _T_78197 = _T_78196[10:0]; // @[Modules.scala 68:83:@32814.4]
  assign buffer_13_672 = $signed(_T_78197); // @[Modules.scala 68:83:@32815.4]
  assign _T_78199 = $signed(buffer_0_395) + $signed(buffer_13_563); // @[Modules.scala 68:83:@32817.4]
  assign _T_78200 = _T_78199[10:0]; // @[Modules.scala 68:83:@32818.4]
  assign buffer_13_673 = $signed(_T_78200); // @[Modules.scala 68:83:@32819.4]
  assign _T_78205 = $signed(buffer_0_566) + $signed(buffer_13_567); // @[Modules.scala 68:83:@32825.4]
  assign _T_78206 = _T_78205[10:0]; // @[Modules.scala 68:83:@32826.4]
  assign buffer_13_675 = $signed(_T_78206); // @[Modules.scala 68:83:@32827.4]
  assign _T_78217 = $signed(buffer_13_574) + $signed(buffer_0_395); // @[Modules.scala 68:83:@32841.4]
  assign _T_78218 = _T_78217[10:0]; // @[Modules.scala 68:83:@32842.4]
  assign buffer_13_679 = $signed(_T_78218); // @[Modules.scala 68:83:@32843.4]
  assign _T_78226 = $signed(buffer_7_580) + $signed(buffer_13_581); // @[Modules.scala 68:83:@32853.4]
  assign _T_78227 = _T_78226[10:0]; // @[Modules.scala 68:83:@32854.4]
  assign buffer_13_682 = $signed(_T_78227); // @[Modules.scala 68:83:@32855.4]
  assign _T_78235 = $signed(buffer_0_395) + $signed(buffer_13_587); // @[Modules.scala 68:83:@32865.4]
  assign _T_78236 = _T_78235[10:0]; // @[Modules.scala 68:83:@32866.4]
  assign buffer_13_685 = $signed(_T_78236); // @[Modules.scala 68:83:@32867.4]
  assign _T_78238 = $signed(buffer_13_588) + $signed(buffer_13_589); // @[Modules.scala 71:109:@32869.4]
  assign _T_78239 = _T_78238[10:0]; // @[Modules.scala 71:109:@32870.4]
  assign buffer_13_686 = $signed(_T_78239); // @[Modules.scala 71:109:@32871.4]
  assign _T_78241 = $signed(buffer_13_590) + $signed(buffer_13_591); // @[Modules.scala 71:109:@32873.4]
  assign _T_78242 = _T_78241[10:0]; // @[Modules.scala 71:109:@32874.4]
  assign buffer_13_687 = $signed(_T_78242); // @[Modules.scala 71:109:@32875.4]
  assign _T_78244 = $signed(buffer_13_592) + $signed(buffer_13_593); // @[Modules.scala 71:109:@32877.4]
  assign _T_78245 = _T_78244[10:0]; // @[Modules.scala 71:109:@32878.4]
  assign buffer_13_688 = $signed(_T_78245); // @[Modules.scala 71:109:@32879.4]
  assign _T_78247 = $signed(buffer_13_594) + $signed(buffer_13_595); // @[Modules.scala 71:109:@32881.4]
  assign _T_78248 = _T_78247[10:0]; // @[Modules.scala 71:109:@32882.4]
  assign buffer_13_689 = $signed(_T_78248); // @[Modules.scala 71:109:@32883.4]
  assign _T_78250 = $signed(buffer_13_596) + $signed(buffer_13_597); // @[Modules.scala 71:109:@32885.4]
  assign _T_78251 = _T_78250[10:0]; // @[Modules.scala 71:109:@32886.4]
  assign buffer_13_690 = $signed(_T_78251); // @[Modules.scala 71:109:@32887.4]
  assign _T_78253 = $signed(buffer_13_598) + $signed(buffer_0_599); // @[Modules.scala 71:109:@32889.4]
  assign _T_78254 = _T_78253[10:0]; // @[Modules.scala 71:109:@32890.4]
  assign buffer_13_691 = $signed(_T_78254); // @[Modules.scala 71:109:@32891.4]
  assign _T_78256 = $signed(buffer_13_600) + $signed(buffer_1_601); // @[Modules.scala 71:109:@32893.4]
  assign _T_78257 = _T_78256[10:0]; // @[Modules.scala 71:109:@32894.4]
  assign buffer_13_692 = $signed(_T_78257); // @[Modules.scala 71:109:@32895.4]
  assign _T_78259 = $signed(buffer_13_602) + $signed(buffer_13_603); // @[Modules.scala 71:109:@32897.4]
  assign _T_78260 = _T_78259[10:0]; // @[Modules.scala 71:109:@32898.4]
  assign buffer_13_693 = $signed(_T_78260); // @[Modules.scala 71:109:@32899.4]
  assign _T_78262 = $signed(buffer_0_593) + $signed(buffer_13_605); // @[Modules.scala 71:109:@32901.4]
  assign _T_78263 = _T_78262[10:0]; // @[Modules.scala 71:109:@32902.4]
  assign buffer_13_694 = $signed(_T_78263); // @[Modules.scala 71:109:@32903.4]
  assign _T_78265 = $signed(buffer_13_606) + $signed(buffer_13_607); // @[Modules.scala 71:109:@32905.4]
  assign _T_78266 = _T_78265[10:0]; // @[Modules.scala 71:109:@32906.4]
  assign buffer_13_695 = $signed(_T_78266); // @[Modules.scala 71:109:@32907.4]
  assign _T_78268 = $signed(buffer_13_608) + $signed(buffer_13_609); // @[Modules.scala 71:109:@32909.4]
  assign _T_78269 = _T_78268[10:0]; // @[Modules.scala 71:109:@32910.4]
  assign buffer_13_696 = $signed(_T_78269); // @[Modules.scala 71:109:@32911.4]
  assign _T_78271 = $signed(buffer_13_610) + $signed(buffer_13_611); // @[Modules.scala 71:109:@32913.4]
  assign _T_78272 = _T_78271[10:0]; // @[Modules.scala 71:109:@32914.4]
  assign buffer_13_697 = $signed(_T_78272); // @[Modules.scala 71:109:@32915.4]
  assign _T_78274 = $signed(buffer_13_612) + $signed(buffer_13_613); // @[Modules.scala 71:109:@32917.4]
  assign _T_78275 = _T_78274[10:0]; // @[Modules.scala 71:109:@32918.4]
  assign buffer_13_698 = $signed(_T_78275); // @[Modules.scala 71:109:@32919.4]
  assign _T_78277 = $signed(buffer_13_614) + $signed(buffer_13_615); // @[Modules.scala 71:109:@32921.4]
  assign _T_78278 = _T_78277[10:0]; // @[Modules.scala 71:109:@32922.4]
  assign buffer_13_699 = $signed(_T_78278); // @[Modules.scala 71:109:@32923.4]
  assign _T_78280 = $signed(buffer_13_616) + $signed(buffer_13_617); // @[Modules.scala 71:109:@32925.4]
  assign _T_78281 = _T_78280[10:0]; // @[Modules.scala 71:109:@32926.4]
  assign buffer_13_700 = $signed(_T_78281); // @[Modules.scala 71:109:@32927.4]
  assign _T_78283 = $signed(buffer_13_618) + $signed(buffer_0_593); // @[Modules.scala 71:109:@32929.4]
  assign _T_78284 = _T_78283[10:0]; // @[Modules.scala 71:109:@32930.4]
  assign buffer_13_701 = $signed(_T_78284); // @[Modules.scala 71:109:@32931.4]
  assign _T_78286 = $signed(buffer_13_620) + $signed(buffer_13_621); // @[Modules.scala 71:109:@32933.4]
  assign _T_78287 = _T_78286[10:0]; // @[Modules.scala 71:109:@32934.4]
  assign buffer_13_702 = $signed(_T_78287); // @[Modules.scala 71:109:@32935.4]
  assign _T_78289 = $signed(buffer_13_622) + $signed(buffer_13_623); // @[Modules.scala 71:109:@32937.4]
  assign _T_78290 = _T_78289[10:0]; // @[Modules.scala 71:109:@32938.4]
  assign buffer_13_703 = $signed(_T_78290); // @[Modules.scala 71:109:@32939.4]
  assign _T_78292 = $signed(buffer_13_624) + $signed(buffer_13_625); // @[Modules.scala 71:109:@32941.4]
  assign _T_78293 = _T_78292[10:0]; // @[Modules.scala 71:109:@32942.4]
  assign buffer_13_704 = $signed(_T_78293); // @[Modules.scala 71:109:@32943.4]
  assign _T_78295 = $signed(buffer_0_593) + $signed(buffer_13_627); // @[Modules.scala 71:109:@32945.4]
  assign _T_78296 = _T_78295[10:0]; // @[Modules.scala 71:109:@32946.4]
  assign buffer_13_705 = $signed(_T_78296); // @[Modules.scala 71:109:@32947.4]
  assign _T_78298 = $signed(buffer_13_628) + $signed(buffer_13_629); // @[Modules.scala 71:109:@32949.4]
  assign _T_78299 = _T_78298[10:0]; // @[Modules.scala 71:109:@32950.4]
  assign buffer_13_706 = $signed(_T_78299); // @[Modules.scala 71:109:@32951.4]
  assign _T_78301 = $signed(buffer_13_630) + $signed(buffer_13_631); // @[Modules.scala 71:109:@32953.4]
  assign _T_78302 = _T_78301[10:0]; // @[Modules.scala 71:109:@32954.4]
  assign buffer_13_707 = $signed(_T_78302); // @[Modules.scala 71:109:@32955.4]
  assign _T_78304 = $signed(buffer_13_632) + $signed(buffer_13_633); // @[Modules.scala 71:109:@32957.4]
  assign _T_78305 = _T_78304[10:0]; // @[Modules.scala 71:109:@32958.4]
  assign buffer_13_708 = $signed(_T_78305); // @[Modules.scala 71:109:@32959.4]
  assign _T_78307 = $signed(buffer_13_634) + $signed(buffer_13_635); // @[Modules.scala 71:109:@32961.4]
  assign _T_78308 = _T_78307[10:0]; // @[Modules.scala 71:109:@32962.4]
  assign buffer_13_709 = $signed(_T_78308); // @[Modules.scala 71:109:@32963.4]
  assign _T_78310 = $signed(buffer_13_636) + $signed(buffer_13_637); // @[Modules.scala 71:109:@32965.4]
  assign _T_78311 = _T_78310[10:0]; // @[Modules.scala 71:109:@32966.4]
  assign buffer_13_710 = $signed(_T_78311); // @[Modules.scala 71:109:@32967.4]
  assign _T_78313 = $signed(buffer_13_638) + $signed(buffer_13_639); // @[Modules.scala 71:109:@32969.4]
  assign _T_78314 = _T_78313[10:0]; // @[Modules.scala 71:109:@32970.4]
  assign buffer_13_711 = $signed(_T_78314); // @[Modules.scala 71:109:@32971.4]
  assign _T_78316 = $signed(buffer_13_640) + $signed(buffer_13_641); // @[Modules.scala 71:109:@32973.4]
  assign _T_78317 = _T_78316[10:0]; // @[Modules.scala 71:109:@32974.4]
  assign buffer_13_712 = $signed(_T_78317); // @[Modules.scala 71:109:@32975.4]
  assign _T_78319 = $signed(buffer_13_642) + $signed(buffer_13_643); // @[Modules.scala 71:109:@32977.4]
  assign _T_78320 = _T_78319[10:0]; // @[Modules.scala 71:109:@32978.4]
  assign buffer_13_713 = $signed(_T_78320); // @[Modules.scala 71:109:@32979.4]
  assign _T_78322 = $signed(buffer_13_644) + $signed(buffer_13_645); // @[Modules.scala 71:109:@32981.4]
  assign _T_78323 = _T_78322[10:0]; // @[Modules.scala 71:109:@32982.4]
  assign buffer_13_714 = $signed(_T_78323); // @[Modules.scala 71:109:@32983.4]
  assign _T_78325 = $signed(buffer_13_646) + $signed(buffer_7_647); // @[Modules.scala 71:109:@32985.4]
  assign _T_78326 = _T_78325[10:0]; // @[Modules.scala 71:109:@32986.4]
  assign buffer_13_715 = $signed(_T_78326); // @[Modules.scala 71:109:@32987.4]
  assign _T_78328 = $signed(buffer_13_648) + $signed(buffer_13_649); // @[Modules.scala 71:109:@32989.4]
  assign _T_78329 = _T_78328[10:0]; // @[Modules.scala 71:109:@32990.4]
  assign buffer_13_716 = $signed(_T_78329); // @[Modules.scala 71:109:@32991.4]
  assign _T_78331 = $signed(buffer_13_650) + $signed(buffer_11_651); // @[Modules.scala 71:109:@32993.4]
  assign _T_78332 = _T_78331[10:0]; // @[Modules.scala 71:109:@32994.4]
  assign buffer_13_717 = $signed(_T_78332); // @[Modules.scala 71:109:@32995.4]
  assign _T_78334 = $signed(buffer_7_652) + $signed(buffer_13_653); // @[Modules.scala 71:109:@32997.4]
  assign _T_78335 = _T_78334[10:0]; // @[Modules.scala 71:109:@32998.4]
  assign buffer_13_718 = $signed(_T_78335); // @[Modules.scala 71:109:@32999.4]
  assign _T_78337 = $signed(buffer_13_654) + $signed(buffer_13_655); // @[Modules.scala 71:109:@33001.4]
  assign _T_78338 = _T_78337[10:0]; // @[Modules.scala 71:109:@33002.4]
  assign buffer_13_719 = $signed(_T_78338); // @[Modules.scala 71:109:@33003.4]
  assign _T_78340 = $signed(buffer_13_656) + $signed(buffer_3_657); // @[Modules.scala 71:109:@33005.4]
  assign _T_78341 = _T_78340[10:0]; // @[Modules.scala 71:109:@33006.4]
  assign buffer_13_720 = $signed(_T_78341); // @[Modules.scala 71:109:@33007.4]
  assign _T_78343 = $signed(buffer_13_658) + $signed(buffer_9_659); // @[Modules.scala 71:109:@33009.4]
  assign _T_78344 = _T_78343[10:0]; // @[Modules.scala 71:109:@33010.4]
  assign buffer_13_721 = $signed(_T_78344); // @[Modules.scala 71:109:@33011.4]
  assign _T_78346 = $signed(buffer_13_660) + $signed(buffer_13_661); // @[Modules.scala 71:109:@33013.4]
  assign _T_78347 = _T_78346[10:0]; // @[Modules.scala 71:109:@33014.4]
  assign buffer_13_722 = $signed(_T_78347); // @[Modules.scala 71:109:@33015.4]
  assign _T_78349 = $signed(buffer_13_662) + $signed(buffer_7_663); // @[Modules.scala 71:109:@33017.4]
  assign _T_78350 = _T_78349[10:0]; // @[Modules.scala 71:109:@33018.4]
  assign buffer_13_723 = $signed(_T_78350); // @[Modules.scala 71:109:@33019.4]
  assign _T_78352 = $signed(buffer_3_664) + $signed(buffer_13_665); // @[Modules.scala 71:109:@33021.4]
  assign _T_78353 = _T_78352[10:0]; // @[Modules.scala 71:109:@33022.4]
  assign buffer_13_724 = $signed(_T_78353); // @[Modules.scala 71:109:@33023.4]
  assign _T_78355 = $signed(buffer_13_666) + $signed(buffer_13_667); // @[Modules.scala 71:109:@33025.4]
  assign _T_78356 = _T_78355[10:0]; // @[Modules.scala 71:109:@33026.4]
  assign buffer_13_725 = $signed(_T_78356); // @[Modules.scala 71:109:@33027.4]
  assign _T_78358 = $signed(buffer_13_668) + $signed(buffer_0_593); // @[Modules.scala 71:109:@33029.4]
  assign _T_78359 = _T_78358[10:0]; // @[Modules.scala 71:109:@33030.4]
  assign buffer_13_726 = $signed(_T_78359); // @[Modules.scala 71:109:@33031.4]
  assign _T_78361 = $signed(buffer_13_670) + $signed(buffer_0_671); // @[Modules.scala 71:109:@33033.4]
  assign _T_78362 = _T_78361[10:0]; // @[Modules.scala 71:109:@33034.4]
  assign buffer_13_727 = $signed(_T_78362); // @[Modules.scala 71:109:@33035.4]
  assign _T_78364 = $signed(buffer_13_672) + $signed(buffer_13_673); // @[Modules.scala 71:109:@33037.4]
  assign _T_78365 = _T_78364[10:0]; // @[Modules.scala 71:109:@33038.4]
  assign buffer_13_728 = $signed(_T_78365); // @[Modules.scala 71:109:@33039.4]
  assign _T_78367 = $signed(buffer_0_674) + $signed(buffer_13_675); // @[Modules.scala 71:109:@33041.4]
  assign _T_78368 = _T_78367[10:0]; // @[Modules.scala 71:109:@33042.4]
  assign buffer_13_729 = $signed(_T_78368); // @[Modules.scala 71:109:@33043.4]
  assign _T_78373 = $signed(buffer_0_593) + $signed(buffer_13_679); // @[Modules.scala 71:109:@33049.4]
  assign _T_78374 = _T_78373[10:0]; // @[Modules.scala 71:109:@33050.4]
  assign buffer_13_731 = $signed(_T_78374); // @[Modules.scala 71:109:@33051.4]
  assign _T_78379 = $signed(buffer_13_682) + $signed(buffer_0_593); // @[Modules.scala 71:109:@33057.4]
  assign _T_78380 = _T_78379[10:0]; // @[Modules.scala 71:109:@33058.4]
  assign buffer_13_733 = $signed(_T_78380); // @[Modules.scala 71:109:@33059.4]
  assign _T_78382 = $signed(buffer_0_593) + $signed(buffer_13_685); // @[Modules.scala 71:109:@33061.4]
  assign _T_78383 = _T_78382[10:0]; // @[Modules.scala 71:109:@33062.4]
  assign buffer_13_734 = $signed(_T_78383); // @[Modules.scala 71:109:@33063.4]
  assign _T_78385 = $signed(buffer_13_686) + $signed(buffer_13_687); // @[Modules.scala 78:156:@33066.4]
  assign _T_78386 = _T_78385[10:0]; // @[Modules.scala 78:156:@33067.4]
  assign buffer_13_736 = $signed(_T_78386); // @[Modules.scala 78:156:@33068.4]
  assign _T_78388 = $signed(buffer_13_736) + $signed(buffer_13_688); // @[Modules.scala 78:156:@33070.4]
  assign _T_78389 = _T_78388[10:0]; // @[Modules.scala 78:156:@33071.4]
  assign buffer_13_737 = $signed(_T_78389); // @[Modules.scala 78:156:@33072.4]
  assign _T_78391 = $signed(buffer_13_737) + $signed(buffer_13_689); // @[Modules.scala 78:156:@33074.4]
  assign _T_78392 = _T_78391[10:0]; // @[Modules.scala 78:156:@33075.4]
  assign buffer_13_738 = $signed(_T_78392); // @[Modules.scala 78:156:@33076.4]
  assign _T_78394 = $signed(buffer_13_738) + $signed(buffer_13_690); // @[Modules.scala 78:156:@33078.4]
  assign _T_78395 = _T_78394[10:0]; // @[Modules.scala 78:156:@33079.4]
  assign buffer_13_739 = $signed(_T_78395); // @[Modules.scala 78:156:@33080.4]
  assign _T_78397 = $signed(buffer_13_739) + $signed(buffer_13_691); // @[Modules.scala 78:156:@33082.4]
  assign _T_78398 = _T_78397[10:0]; // @[Modules.scala 78:156:@33083.4]
  assign buffer_13_740 = $signed(_T_78398); // @[Modules.scala 78:156:@33084.4]
  assign _T_78400 = $signed(buffer_13_740) + $signed(buffer_13_692); // @[Modules.scala 78:156:@33086.4]
  assign _T_78401 = _T_78400[10:0]; // @[Modules.scala 78:156:@33087.4]
  assign buffer_13_741 = $signed(_T_78401); // @[Modules.scala 78:156:@33088.4]
  assign _T_78403 = $signed(buffer_13_741) + $signed(buffer_13_693); // @[Modules.scala 78:156:@33090.4]
  assign _T_78404 = _T_78403[10:0]; // @[Modules.scala 78:156:@33091.4]
  assign buffer_13_742 = $signed(_T_78404); // @[Modules.scala 78:156:@33092.4]
  assign _T_78406 = $signed(buffer_13_742) + $signed(buffer_13_694); // @[Modules.scala 78:156:@33094.4]
  assign _T_78407 = _T_78406[10:0]; // @[Modules.scala 78:156:@33095.4]
  assign buffer_13_743 = $signed(_T_78407); // @[Modules.scala 78:156:@33096.4]
  assign _T_78409 = $signed(buffer_13_743) + $signed(buffer_13_695); // @[Modules.scala 78:156:@33098.4]
  assign _T_78410 = _T_78409[10:0]; // @[Modules.scala 78:156:@33099.4]
  assign buffer_13_744 = $signed(_T_78410); // @[Modules.scala 78:156:@33100.4]
  assign _T_78412 = $signed(buffer_13_744) + $signed(buffer_13_696); // @[Modules.scala 78:156:@33102.4]
  assign _T_78413 = _T_78412[10:0]; // @[Modules.scala 78:156:@33103.4]
  assign buffer_13_745 = $signed(_T_78413); // @[Modules.scala 78:156:@33104.4]
  assign _T_78415 = $signed(buffer_13_745) + $signed(buffer_13_697); // @[Modules.scala 78:156:@33106.4]
  assign _T_78416 = _T_78415[10:0]; // @[Modules.scala 78:156:@33107.4]
  assign buffer_13_746 = $signed(_T_78416); // @[Modules.scala 78:156:@33108.4]
  assign _T_78418 = $signed(buffer_13_746) + $signed(buffer_13_698); // @[Modules.scala 78:156:@33110.4]
  assign _T_78419 = _T_78418[10:0]; // @[Modules.scala 78:156:@33111.4]
  assign buffer_13_747 = $signed(_T_78419); // @[Modules.scala 78:156:@33112.4]
  assign _T_78421 = $signed(buffer_13_747) + $signed(buffer_13_699); // @[Modules.scala 78:156:@33114.4]
  assign _T_78422 = _T_78421[10:0]; // @[Modules.scala 78:156:@33115.4]
  assign buffer_13_748 = $signed(_T_78422); // @[Modules.scala 78:156:@33116.4]
  assign _T_78424 = $signed(buffer_13_748) + $signed(buffer_13_700); // @[Modules.scala 78:156:@33118.4]
  assign _T_78425 = _T_78424[10:0]; // @[Modules.scala 78:156:@33119.4]
  assign buffer_13_749 = $signed(_T_78425); // @[Modules.scala 78:156:@33120.4]
  assign _T_78427 = $signed(buffer_13_749) + $signed(buffer_13_701); // @[Modules.scala 78:156:@33122.4]
  assign _T_78428 = _T_78427[10:0]; // @[Modules.scala 78:156:@33123.4]
  assign buffer_13_750 = $signed(_T_78428); // @[Modules.scala 78:156:@33124.4]
  assign _T_78430 = $signed(buffer_13_750) + $signed(buffer_13_702); // @[Modules.scala 78:156:@33126.4]
  assign _T_78431 = _T_78430[10:0]; // @[Modules.scala 78:156:@33127.4]
  assign buffer_13_751 = $signed(_T_78431); // @[Modules.scala 78:156:@33128.4]
  assign _T_78433 = $signed(buffer_13_751) + $signed(buffer_13_703); // @[Modules.scala 78:156:@33130.4]
  assign _T_78434 = _T_78433[10:0]; // @[Modules.scala 78:156:@33131.4]
  assign buffer_13_752 = $signed(_T_78434); // @[Modules.scala 78:156:@33132.4]
  assign _T_78436 = $signed(buffer_13_752) + $signed(buffer_13_704); // @[Modules.scala 78:156:@33134.4]
  assign _T_78437 = _T_78436[10:0]; // @[Modules.scala 78:156:@33135.4]
  assign buffer_13_753 = $signed(_T_78437); // @[Modules.scala 78:156:@33136.4]
  assign _T_78439 = $signed(buffer_13_753) + $signed(buffer_13_705); // @[Modules.scala 78:156:@33138.4]
  assign _T_78440 = _T_78439[10:0]; // @[Modules.scala 78:156:@33139.4]
  assign buffer_13_754 = $signed(_T_78440); // @[Modules.scala 78:156:@33140.4]
  assign _T_78442 = $signed(buffer_13_754) + $signed(buffer_13_706); // @[Modules.scala 78:156:@33142.4]
  assign _T_78443 = _T_78442[10:0]; // @[Modules.scala 78:156:@33143.4]
  assign buffer_13_755 = $signed(_T_78443); // @[Modules.scala 78:156:@33144.4]
  assign _T_78445 = $signed(buffer_13_755) + $signed(buffer_13_707); // @[Modules.scala 78:156:@33146.4]
  assign _T_78446 = _T_78445[10:0]; // @[Modules.scala 78:156:@33147.4]
  assign buffer_13_756 = $signed(_T_78446); // @[Modules.scala 78:156:@33148.4]
  assign _T_78448 = $signed(buffer_13_756) + $signed(buffer_13_708); // @[Modules.scala 78:156:@33150.4]
  assign _T_78449 = _T_78448[10:0]; // @[Modules.scala 78:156:@33151.4]
  assign buffer_13_757 = $signed(_T_78449); // @[Modules.scala 78:156:@33152.4]
  assign _T_78451 = $signed(buffer_13_757) + $signed(buffer_13_709); // @[Modules.scala 78:156:@33154.4]
  assign _T_78452 = _T_78451[10:0]; // @[Modules.scala 78:156:@33155.4]
  assign buffer_13_758 = $signed(_T_78452); // @[Modules.scala 78:156:@33156.4]
  assign _T_78454 = $signed(buffer_13_758) + $signed(buffer_13_710); // @[Modules.scala 78:156:@33158.4]
  assign _T_78455 = _T_78454[10:0]; // @[Modules.scala 78:156:@33159.4]
  assign buffer_13_759 = $signed(_T_78455); // @[Modules.scala 78:156:@33160.4]
  assign _T_78457 = $signed(buffer_13_759) + $signed(buffer_13_711); // @[Modules.scala 78:156:@33162.4]
  assign _T_78458 = _T_78457[10:0]; // @[Modules.scala 78:156:@33163.4]
  assign buffer_13_760 = $signed(_T_78458); // @[Modules.scala 78:156:@33164.4]
  assign _T_78460 = $signed(buffer_13_760) + $signed(buffer_13_712); // @[Modules.scala 78:156:@33166.4]
  assign _T_78461 = _T_78460[10:0]; // @[Modules.scala 78:156:@33167.4]
  assign buffer_13_761 = $signed(_T_78461); // @[Modules.scala 78:156:@33168.4]
  assign _T_78463 = $signed(buffer_13_761) + $signed(buffer_13_713); // @[Modules.scala 78:156:@33170.4]
  assign _T_78464 = _T_78463[10:0]; // @[Modules.scala 78:156:@33171.4]
  assign buffer_13_762 = $signed(_T_78464); // @[Modules.scala 78:156:@33172.4]
  assign _T_78466 = $signed(buffer_13_762) + $signed(buffer_13_714); // @[Modules.scala 78:156:@33174.4]
  assign _T_78467 = _T_78466[10:0]; // @[Modules.scala 78:156:@33175.4]
  assign buffer_13_763 = $signed(_T_78467); // @[Modules.scala 78:156:@33176.4]
  assign _T_78469 = $signed(buffer_13_763) + $signed(buffer_13_715); // @[Modules.scala 78:156:@33178.4]
  assign _T_78470 = _T_78469[10:0]; // @[Modules.scala 78:156:@33179.4]
  assign buffer_13_764 = $signed(_T_78470); // @[Modules.scala 78:156:@33180.4]
  assign _T_78472 = $signed(buffer_13_764) + $signed(buffer_13_716); // @[Modules.scala 78:156:@33182.4]
  assign _T_78473 = _T_78472[10:0]; // @[Modules.scala 78:156:@33183.4]
  assign buffer_13_765 = $signed(_T_78473); // @[Modules.scala 78:156:@33184.4]
  assign _T_78475 = $signed(buffer_13_765) + $signed(buffer_13_717); // @[Modules.scala 78:156:@33186.4]
  assign _T_78476 = _T_78475[10:0]; // @[Modules.scala 78:156:@33187.4]
  assign buffer_13_766 = $signed(_T_78476); // @[Modules.scala 78:156:@33188.4]
  assign _T_78478 = $signed(buffer_13_766) + $signed(buffer_13_718); // @[Modules.scala 78:156:@33190.4]
  assign _T_78479 = _T_78478[10:0]; // @[Modules.scala 78:156:@33191.4]
  assign buffer_13_767 = $signed(_T_78479); // @[Modules.scala 78:156:@33192.4]
  assign _T_78481 = $signed(buffer_13_767) + $signed(buffer_13_719); // @[Modules.scala 78:156:@33194.4]
  assign _T_78482 = _T_78481[10:0]; // @[Modules.scala 78:156:@33195.4]
  assign buffer_13_768 = $signed(_T_78482); // @[Modules.scala 78:156:@33196.4]
  assign _T_78484 = $signed(buffer_13_768) + $signed(buffer_13_720); // @[Modules.scala 78:156:@33198.4]
  assign _T_78485 = _T_78484[10:0]; // @[Modules.scala 78:156:@33199.4]
  assign buffer_13_769 = $signed(_T_78485); // @[Modules.scala 78:156:@33200.4]
  assign _T_78487 = $signed(buffer_13_769) + $signed(buffer_13_721); // @[Modules.scala 78:156:@33202.4]
  assign _T_78488 = _T_78487[10:0]; // @[Modules.scala 78:156:@33203.4]
  assign buffer_13_770 = $signed(_T_78488); // @[Modules.scala 78:156:@33204.4]
  assign _T_78490 = $signed(buffer_13_770) + $signed(buffer_13_722); // @[Modules.scala 78:156:@33206.4]
  assign _T_78491 = _T_78490[10:0]; // @[Modules.scala 78:156:@33207.4]
  assign buffer_13_771 = $signed(_T_78491); // @[Modules.scala 78:156:@33208.4]
  assign _T_78493 = $signed(buffer_13_771) + $signed(buffer_13_723); // @[Modules.scala 78:156:@33210.4]
  assign _T_78494 = _T_78493[10:0]; // @[Modules.scala 78:156:@33211.4]
  assign buffer_13_772 = $signed(_T_78494); // @[Modules.scala 78:156:@33212.4]
  assign _T_78496 = $signed(buffer_13_772) + $signed(buffer_13_724); // @[Modules.scala 78:156:@33214.4]
  assign _T_78497 = _T_78496[10:0]; // @[Modules.scala 78:156:@33215.4]
  assign buffer_13_773 = $signed(_T_78497); // @[Modules.scala 78:156:@33216.4]
  assign _T_78499 = $signed(buffer_13_773) + $signed(buffer_13_725); // @[Modules.scala 78:156:@33218.4]
  assign _T_78500 = _T_78499[10:0]; // @[Modules.scala 78:156:@33219.4]
  assign buffer_13_774 = $signed(_T_78500); // @[Modules.scala 78:156:@33220.4]
  assign _T_78502 = $signed(buffer_13_774) + $signed(buffer_13_726); // @[Modules.scala 78:156:@33222.4]
  assign _T_78503 = _T_78502[10:0]; // @[Modules.scala 78:156:@33223.4]
  assign buffer_13_775 = $signed(_T_78503); // @[Modules.scala 78:156:@33224.4]
  assign _T_78505 = $signed(buffer_13_775) + $signed(buffer_13_727); // @[Modules.scala 78:156:@33226.4]
  assign _T_78506 = _T_78505[10:0]; // @[Modules.scala 78:156:@33227.4]
  assign buffer_13_776 = $signed(_T_78506); // @[Modules.scala 78:156:@33228.4]
  assign _T_78508 = $signed(buffer_13_776) + $signed(buffer_13_728); // @[Modules.scala 78:156:@33230.4]
  assign _T_78509 = _T_78508[10:0]; // @[Modules.scala 78:156:@33231.4]
  assign buffer_13_777 = $signed(_T_78509); // @[Modules.scala 78:156:@33232.4]
  assign _T_78511 = $signed(buffer_13_777) + $signed(buffer_13_729); // @[Modules.scala 78:156:@33234.4]
  assign _T_78512 = _T_78511[10:0]; // @[Modules.scala 78:156:@33235.4]
  assign buffer_13_778 = $signed(_T_78512); // @[Modules.scala 78:156:@33236.4]
  assign _T_78514 = $signed(buffer_13_778) + $signed(buffer_0_701); // @[Modules.scala 78:156:@33238.4]
  assign _T_78515 = _T_78514[10:0]; // @[Modules.scala 78:156:@33239.4]
  assign buffer_13_779 = $signed(_T_78515); // @[Modules.scala 78:156:@33240.4]
  assign _T_78517 = $signed(buffer_13_779) + $signed(buffer_13_731); // @[Modules.scala 78:156:@33242.4]
  assign _T_78518 = _T_78517[10:0]; // @[Modules.scala 78:156:@33243.4]
  assign buffer_13_780 = $signed(_T_78518); // @[Modules.scala 78:156:@33244.4]
  assign _T_78520 = $signed(buffer_13_780) + $signed(buffer_0_701); // @[Modules.scala 78:156:@33246.4]
  assign _T_78521 = _T_78520[10:0]; // @[Modules.scala 78:156:@33247.4]
  assign buffer_13_781 = $signed(_T_78521); // @[Modules.scala 78:156:@33248.4]
  assign _T_78523 = $signed(buffer_13_781) + $signed(buffer_13_733); // @[Modules.scala 78:156:@33250.4]
  assign _T_78524 = _T_78523[10:0]; // @[Modules.scala 78:156:@33251.4]
  assign buffer_13_782 = $signed(_T_78524); // @[Modules.scala 78:156:@33252.4]
  assign _T_78526 = $signed(buffer_13_782) + $signed(buffer_13_734); // @[Modules.scala 78:156:@33254.4]
  assign _T_78527 = _T_78526[10:0]; // @[Modules.scala 78:156:@33255.4]
  assign buffer_13_783 = $signed(_T_78527); // @[Modules.scala 78:156:@33256.4]
  assign _T_79137 = $signed(buffer_0_0) + $signed(buffer_3_1); // @[Modules.scala 65:57:@34137.4]
  assign _T_79138 = _T_79137[10:0]; // @[Modules.scala 65:57:@34138.4]
  assign buffer_14_392 = $signed(_T_79138); // @[Modules.scala 65:57:@34139.4]
  assign _T_79143 = $signed(buffer_0_4) + $signed(buffer_4_5); // @[Modules.scala 65:57:@34145.4]
  assign _T_79144 = _T_79143[10:0]; // @[Modules.scala 65:57:@34146.4]
  assign buffer_14_394 = $signed(_T_79144); // @[Modules.scala 65:57:@34147.4]
  assign _T_79158 = $signed(buffer_3_14) + $signed(buffer_2_15); // @[Modules.scala 65:57:@34165.4]
  assign _T_79159 = _T_79158[10:0]; // @[Modules.scala 65:57:@34166.4]
  assign buffer_14_399 = $signed(_T_79159); // @[Modules.scala 65:57:@34167.4]
  assign _T_79167 = $signed(11'sh0) + $signed(buffer_1_21); // @[Modules.scala 65:57:@34177.4]
  assign _T_79168 = _T_79167[10:0]; // @[Modules.scala 65:57:@34178.4]
  assign buffer_14_402 = $signed(_T_79168); // @[Modules.scala 65:57:@34179.4]
  assign _T_79176 = $signed(buffer_1_26) + $signed(buffer_7_27); // @[Modules.scala 65:57:@34189.4]
  assign _T_79177 = _T_79176[10:0]; // @[Modules.scala 65:57:@34190.4]
  assign buffer_14_405 = $signed(_T_79177); // @[Modules.scala 65:57:@34191.4]
  assign buffer_14_30 = {{6{io_in_60[4]}},io_in_60}; // @[Modules.scala 32:22:@8.4]
  assign _T_79182 = $signed(buffer_14_30) + $signed(buffer_1_31); // @[Modules.scala 65:57:@34197.4]
  assign _T_79183 = _T_79182[10:0]; // @[Modules.scala 65:57:@34198.4]
  assign buffer_14_407 = $signed(_T_79183); // @[Modules.scala 65:57:@34199.4]
  assign _T_79200 = $signed(buffer_5_42) + $signed(buffer_1_43); // @[Modules.scala 65:57:@34221.4]
  assign _T_79201 = _T_79200[10:0]; // @[Modules.scala 65:57:@34222.4]
  assign buffer_14_413 = $signed(_T_79201); // @[Modules.scala 65:57:@34223.4]
  assign buffer_14_45 = {{6{io_in_91[4]}},io_in_91}; // @[Modules.scala 32:22:@8.4]
  assign _T_79203 = $signed(buffer_2_44) + $signed(buffer_14_45); // @[Modules.scala 65:57:@34225.4]
  assign _T_79204 = _T_79203[10:0]; // @[Modules.scala 65:57:@34226.4]
  assign buffer_14_414 = $signed(_T_79204); // @[Modules.scala 65:57:@34227.4]
  assign buffer_14_48 = {{6{io_in_96[4]}},io_in_96}; // @[Modules.scala 32:22:@8.4]
  assign _T_79209 = $signed(buffer_14_48) + $signed(11'sh0); // @[Modules.scala 65:57:@34233.4]
  assign _T_79210 = _T_79209[10:0]; // @[Modules.scala 65:57:@34234.4]
  assign buffer_14_416 = $signed(_T_79210); // @[Modules.scala 65:57:@34235.4]
  assign _T_79221 = $signed(buffer_3_56) + $signed(11'sh0); // @[Modules.scala 65:57:@34249.4]
  assign _T_79222 = _T_79221[10:0]; // @[Modules.scala 65:57:@34250.4]
  assign buffer_14_420 = $signed(_T_79222); // @[Modules.scala 65:57:@34251.4]
  assign _T_79230 = $signed(buffer_3_62) + $signed(11'sh0); // @[Modules.scala 65:57:@34261.4]
  assign _T_79231 = _T_79230[10:0]; // @[Modules.scala 65:57:@34262.4]
  assign buffer_14_423 = $signed(_T_79231); // @[Modules.scala 65:57:@34263.4]
  assign _T_79242 = $signed(11'sh0) + $signed(buffer_5_71); // @[Modules.scala 65:57:@34277.4]
  assign _T_79243 = _T_79242[10:0]; // @[Modules.scala 65:57:@34278.4]
  assign buffer_14_427 = $signed(_T_79243); // @[Modules.scala 65:57:@34279.4]
  assign buffer_14_88 = {{6{io_in_177[4]}},io_in_177}; // @[Modules.scala 32:22:@8.4]
  assign _T_79269 = $signed(buffer_14_88) + $signed(11'sh0); // @[Modules.scala 65:57:@34313.4]
  assign _T_79270 = _T_79269[10:0]; // @[Modules.scala 65:57:@34314.4]
  assign buffer_14_436 = $signed(_T_79270); // @[Modules.scala 65:57:@34315.4]
  assign _T_79275 = $signed(buffer_5_92) + $signed(buffer_0_93); // @[Modules.scala 65:57:@34321.4]
  assign _T_79276 = _T_79275[10:0]; // @[Modules.scala 65:57:@34322.4]
  assign buffer_14_438 = $signed(_T_79276); // @[Modules.scala 65:57:@34323.4]
  assign _T_79278 = $signed(buffer_4_94) + $signed(11'sh0); // @[Modules.scala 65:57:@34325.4]
  assign _T_79279 = _T_79278[10:0]; // @[Modules.scala 65:57:@34326.4]
  assign buffer_14_439 = $signed(_T_79279); // @[Modules.scala 65:57:@34327.4]
  assign _T_79317 = $signed(buffer_1_120) + $signed(buffer_6_121); // @[Modules.scala 65:57:@34377.4]
  assign _T_79318 = _T_79317[10:0]; // @[Modules.scala 65:57:@34378.4]
  assign buffer_14_452 = $signed(_T_79318); // @[Modules.scala 65:57:@34379.4]
  assign buffer_14_134 = {{6{io_in_269[4]}},io_in_269}; // @[Modules.scala 32:22:@8.4]
  assign _T_79338 = $signed(buffer_14_134) + $signed(buffer_3_135); // @[Modules.scala 65:57:@34405.4]
  assign _T_79339 = _T_79338[10:0]; // @[Modules.scala 65:57:@34406.4]
  assign buffer_14_459 = $signed(_T_79339); // @[Modules.scala 65:57:@34407.4]
  assign _T_79341 = $signed(buffer_5_136) + $signed(buffer_1_137); // @[Modules.scala 65:57:@34409.4]
  assign _T_79342 = _T_79341[10:0]; // @[Modules.scala 65:57:@34410.4]
  assign buffer_14_460 = $signed(_T_79342); // @[Modules.scala 65:57:@34411.4]
  assign _T_79344 = $signed(buffer_1_138) + $signed(buffer_5_139); // @[Modules.scala 65:57:@34413.4]
  assign _T_79345 = _T_79344[10:0]; // @[Modules.scala 65:57:@34414.4]
  assign buffer_14_461 = $signed(_T_79345); // @[Modules.scala 65:57:@34415.4]
  assign buffer_14_164 = {{6{io_in_328[4]}},io_in_328}; // @[Modules.scala 32:22:@8.4]
  assign _T_79383 = $signed(buffer_14_164) + $signed(buffer_5_165); // @[Modules.scala 65:57:@34465.4]
  assign _T_79384 = _T_79383[10:0]; // @[Modules.scala 65:57:@34466.4]
  assign buffer_14_474 = $signed(_T_79384); // @[Modules.scala 65:57:@34467.4]
  assign _T_79392 = $signed(buffer_0_170) + $signed(11'sh0); // @[Modules.scala 65:57:@34477.4]
  assign _T_79393 = _T_79392[10:0]; // @[Modules.scala 65:57:@34478.4]
  assign buffer_14_477 = $signed(_T_79393); // @[Modules.scala 65:57:@34479.4]
  assign buffer_14_173 = {{6{io_in_346[4]}},io_in_346}; // @[Modules.scala 32:22:@8.4]
  assign _T_79395 = $signed(11'sh0) + $signed(buffer_14_173); // @[Modules.scala 65:57:@34481.4]
  assign _T_79396 = _T_79395[10:0]; // @[Modules.scala 65:57:@34482.4]
  assign buffer_14_478 = $signed(_T_79396); // @[Modules.scala 65:57:@34483.4]
  assign buffer_14_180 = {{6{io_in_360[4]}},io_in_360}; // @[Modules.scala 32:22:@8.4]
  assign _T_79407 = $signed(buffer_14_180) + $signed(buffer_2_181); // @[Modules.scala 65:57:@34497.4]
  assign _T_79408 = _T_79407[10:0]; // @[Modules.scala 65:57:@34498.4]
  assign buffer_14_482 = $signed(_T_79408); // @[Modules.scala 65:57:@34499.4]
  assign _T_79413 = $signed(buffer_1_184) + $signed(buffer_11_185); // @[Modules.scala 65:57:@34505.4]
  assign _T_79414 = _T_79413[10:0]; // @[Modules.scala 65:57:@34506.4]
  assign buffer_14_484 = $signed(_T_79414); // @[Modules.scala 65:57:@34507.4]
  assign _T_79416 = $signed(buffer_11_186) + $signed(buffer_3_187); // @[Modules.scala 65:57:@34509.4]
  assign _T_79417 = _T_79416[10:0]; // @[Modules.scala 65:57:@34510.4]
  assign buffer_14_485 = $signed(_T_79417); // @[Modules.scala 65:57:@34511.4]
  assign _T_79425 = $signed(buffer_0_192) + $signed(11'sh0); // @[Modules.scala 65:57:@34521.4]
  assign _T_79426 = _T_79425[10:0]; // @[Modules.scala 65:57:@34522.4]
  assign buffer_14_488 = $signed(_T_79426); // @[Modules.scala 65:57:@34523.4]
  assign _T_79449 = $signed(11'sh0) + $signed(buffer_4_209); // @[Modules.scala 65:57:@34553.4]
  assign _T_79450 = _T_79449[10:0]; // @[Modules.scala 65:57:@34554.4]
  assign buffer_14_496 = $signed(_T_79450); // @[Modules.scala 65:57:@34555.4]
  assign buffer_14_215 = {{6{io_in_430[4]}},io_in_430}; // @[Modules.scala 32:22:@8.4]
  assign _T_79458 = $signed(buffer_0_214) + $signed(buffer_14_215); // @[Modules.scala 65:57:@34565.4]
  assign _T_79459 = _T_79458[10:0]; // @[Modules.scala 65:57:@34566.4]
  assign buffer_14_499 = $signed(_T_79459); // @[Modules.scala 65:57:@34567.4]
  assign buffer_14_216 = {{6{io_in_433[4]}},io_in_433}; // @[Modules.scala 32:22:@8.4]
  assign _T_79461 = $signed(buffer_14_216) + $signed(11'sh0); // @[Modules.scala 65:57:@34569.4]
  assign _T_79462 = _T_79461[10:0]; // @[Modules.scala 65:57:@34570.4]
  assign buffer_14_500 = $signed(_T_79462); // @[Modules.scala 65:57:@34571.4]
  assign _T_79464 = $signed(buffer_4_218) + $signed(11'sh0); // @[Modules.scala 65:57:@34573.4]
  assign _T_79465 = _T_79464[10:0]; // @[Modules.scala 65:57:@34574.4]
  assign buffer_14_501 = $signed(_T_79465); // @[Modules.scala 65:57:@34575.4]
  assign _T_79485 = $signed(11'sh0) + $signed(buffer_6_233); // @[Modules.scala 65:57:@34601.4]
  assign _T_79486 = _T_79485[10:0]; // @[Modules.scala 65:57:@34602.4]
  assign buffer_14_508 = $signed(_T_79486); // @[Modules.scala 65:57:@34603.4]
  assign _T_79488 = $signed(11'sh0) + $signed(buffer_6_235); // @[Modules.scala 65:57:@34605.4]
  assign _T_79489 = _T_79488[10:0]; // @[Modules.scala 65:57:@34606.4]
  assign buffer_14_509 = $signed(_T_79489); // @[Modules.scala 65:57:@34607.4]
  assign _T_79491 = $signed(11'sh0) + $signed(buffer_3_237); // @[Modules.scala 65:57:@34609.4]
  assign _T_79492 = _T_79491[10:0]; // @[Modules.scala 65:57:@34610.4]
  assign buffer_14_510 = $signed(_T_79492); // @[Modules.scala 65:57:@34611.4]
  assign _T_79494 = $signed(buffer_12_238) + $signed(buffer_1_239); // @[Modules.scala 65:57:@34613.4]
  assign _T_79495 = _T_79494[10:0]; // @[Modules.scala 65:57:@34614.4]
  assign buffer_14_511 = $signed(_T_79495); // @[Modules.scala 65:57:@34615.4]
  assign _T_79503 = $signed(buffer_12_244) + $signed(11'sh0); // @[Modules.scala 65:57:@34625.4]
  assign _T_79504 = _T_79503[10:0]; // @[Modules.scala 65:57:@34626.4]
  assign buffer_14_514 = $signed(_T_79504); // @[Modules.scala 65:57:@34627.4]
  assign _T_79509 = $signed(buffer_13_248) + $signed(buffer_0_249); // @[Modules.scala 65:57:@34633.4]
  assign _T_79510 = _T_79509[10:0]; // @[Modules.scala 65:57:@34634.4]
  assign buffer_14_516 = $signed(_T_79510); // @[Modules.scala 65:57:@34635.4]
  assign _T_79515 = $signed(buffer_3_252) + $signed(buffer_0_253); // @[Modules.scala 65:57:@34641.4]
  assign _T_79516 = _T_79515[10:0]; // @[Modules.scala 65:57:@34642.4]
  assign buffer_14_518 = $signed(_T_79516); // @[Modules.scala 65:57:@34643.4]
  assign _T_79524 = $signed(11'sh0) + $signed(buffer_4_259); // @[Modules.scala 65:57:@34653.4]
  assign _T_79525 = _T_79524[10:0]; // @[Modules.scala 65:57:@34654.4]
  assign buffer_14_521 = $signed(_T_79525); // @[Modules.scala 65:57:@34655.4]
  assign _T_79536 = $signed(buffer_0_266) + $signed(buffer_1_267); // @[Modules.scala 65:57:@34669.4]
  assign _T_79537 = _T_79536[10:0]; // @[Modules.scala 65:57:@34670.4]
  assign buffer_14_525 = $signed(_T_79537); // @[Modules.scala 65:57:@34671.4]
  assign _T_79542 = $signed(buffer_1_270) + $signed(11'sh0); // @[Modules.scala 65:57:@34677.4]
  assign _T_79543 = _T_79542[10:0]; // @[Modules.scala 65:57:@34678.4]
  assign buffer_14_527 = $signed(_T_79543); // @[Modules.scala 65:57:@34679.4]
  assign _T_79557 = $signed(buffer_12_280) + $signed(buffer_1_281); // @[Modules.scala 65:57:@34697.4]
  assign _T_79558 = _T_79557[10:0]; // @[Modules.scala 65:57:@34698.4]
  assign buffer_14_532 = $signed(_T_79558); // @[Modules.scala 65:57:@34699.4]
  assign buffer_14_284 = {{6{io_in_568[4]}},io_in_568}; // @[Modules.scala 32:22:@8.4]
  assign _T_79563 = $signed(buffer_14_284) + $signed(11'sh0); // @[Modules.scala 65:57:@34705.4]
  assign _T_79564 = _T_79563[10:0]; // @[Modules.scala 65:57:@34706.4]
  assign buffer_14_534 = $signed(_T_79564); // @[Modules.scala 65:57:@34707.4]
  assign _T_79569 = $signed(buffer_12_288) + $signed(buffer_5_289); // @[Modules.scala 65:57:@34713.4]
  assign _T_79570 = _T_79569[10:0]; // @[Modules.scala 65:57:@34714.4]
  assign buffer_14_536 = $signed(_T_79570); // @[Modules.scala 65:57:@34715.4]
  assign _T_79578 = $signed(buffer_6_294) + $signed(buffer_1_295); // @[Modules.scala 65:57:@34725.4]
  assign _T_79579 = _T_79578[10:0]; // @[Modules.scala 65:57:@34726.4]
  assign buffer_14_539 = $signed(_T_79579); // @[Modules.scala 65:57:@34727.4]
  assign _T_79590 = $signed(11'sh0) + $signed(buffer_0_303); // @[Modules.scala 65:57:@34741.4]
  assign _T_79591 = _T_79590[10:0]; // @[Modules.scala 65:57:@34742.4]
  assign buffer_14_543 = $signed(_T_79591); // @[Modules.scala 65:57:@34743.4]
  assign _T_79599 = $signed(buffer_2_308) + $signed(buffer_0_309); // @[Modules.scala 65:57:@34753.4]
  assign _T_79600 = _T_79599[10:0]; // @[Modules.scala 65:57:@34754.4]
  assign buffer_14_546 = $signed(_T_79600); // @[Modules.scala 65:57:@34755.4]
  assign _T_79602 = $signed(buffer_1_310) + $signed(buffer_4_311); // @[Modules.scala 65:57:@34757.4]
  assign _T_79603 = _T_79602[10:0]; // @[Modules.scala 65:57:@34758.4]
  assign buffer_14_547 = $signed(_T_79603); // @[Modules.scala 65:57:@34759.4]
  assign _T_79617 = $signed(buffer_5_320) + $signed(11'sh0); // @[Modules.scala 65:57:@34777.4]
  assign _T_79618 = _T_79617[10:0]; // @[Modules.scala 65:57:@34778.4]
  assign buffer_14_552 = $signed(_T_79618); // @[Modules.scala 65:57:@34779.4]
  assign _T_79626 = $signed(11'sh0) + $signed(buffer_1_327); // @[Modules.scala 65:57:@34789.4]
  assign _T_79627 = _T_79626[10:0]; // @[Modules.scala 65:57:@34790.4]
  assign buffer_14_555 = $signed(_T_79627); // @[Modules.scala 65:57:@34791.4]
  assign _T_79659 = $signed(buffer_1_348) + $signed(buffer_0_349); // @[Modules.scala 65:57:@34833.4]
  assign _T_79660 = _T_79659[10:0]; // @[Modules.scala 65:57:@34834.4]
  assign buffer_14_566 = $signed(_T_79660); // @[Modules.scala 65:57:@34835.4]
  assign _T_79665 = $signed(buffer_5_352) + $signed(buffer_10_353); // @[Modules.scala 65:57:@34841.4]
  assign _T_79666 = _T_79665[10:0]; // @[Modules.scala 65:57:@34842.4]
  assign buffer_14_568 = $signed(_T_79666); // @[Modules.scala 65:57:@34843.4]
  assign buffer_14_354 = {{6{io_in_709[4]}},io_in_709}; // @[Modules.scala 32:22:@8.4]
  assign _T_79668 = $signed(buffer_14_354) + $signed(buffer_0_355); // @[Modules.scala 65:57:@34845.4]
  assign _T_79669 = _T_79668[10:0]; // @[Modules.scala 65:57:@34846.4]
  assign buffer_14_569 = $signed(_T_79669); // @[Modules.scala 65:57:@34847.4]
  assign _T_79671 = $signed(buffer_9_356) + $signed(buffer_0_357); // @[Modules.scala 65:57:@34849.4]
  assign _T_79672 = _T_79671[10:0]; // @[Modules.scala 65:57:@34850.4]
  assign buffer_14_570 = $signed(_T_79672); // @[Modules.scala 65:57:@34851.4]
  assign buffer_14_363 = {{6{io_in_727[4]}},io_in_727}; // @[Modules.scala 32:22:@8.4]
  assign _T_79680 = $signed(buffer_1_362) + $signed(buffer_14_363); // @[Modules.scala 65:57:@34861.4]
  assign _T_79681 = _T_79680[10:0]; // @[Modules.scala 65:57:@34862.4]
  assign buffer_14_573 = $signed(_T_79681); // @[Modules.scala 65:57:@34863.4]
  assign _T_79683 = $signed(buffer_9_364) + $signed(buffer_0_365); // @[Modules.scala 65:57:@34865.4]
  assign _T_79684 = _T_79683[10:0]; // @[Modules.scala 65:57:@34866.4]
  assign buffer_14_574 = $signed(_T_79684); // @[Modules.scala 65:57:@34867.4]
  assign buffer_14_367 = {{6{io_in_735[4]}},io_in_735}; // @[Modules.scala 32:22:@8.4]
  assign _T_79686 = $signed(buffer_0_366) + $signed(buffer_14_367); // @[Modules.scala 65:57:@34869.4]
  assign _T_79687 = _T_79686[10:0]; // @[Modules.scala 65:57:@34870.4]
  assign buffer_14_575 = $signed(_T_79687); // @[Modules.scala 65:57:@34871.4]
  assign buffer_14_368 = {{6{io_in_736[4]}},io_in_736}; // @[Modules.scala 32:22:@8.4]
  assign buffer_14_369 = {{6{io_in_738[4]}},io_in_738}; // @[Modules.scala 32:22:@8.4]
  assign _T_79689 = $signed(buffer_14_368) + $signed(buffer_14_369); // @[Modules.scala 65:57:@34873.4]
  assign _T_79690 = _T_79689[10:0]; // @[Modules.scala 65:57:@34874.4]
  assign buffer_14_576 = $signed(_T_79690); // @[Modules.scala 65:57:@34875.4]
  assign _T_79692 = $signed(buffer_0_370) + $signed(buffer_5_371); // @[Modules.scala 65:57:@34877.4]
  assign _T_79693 = _T_79692[10:0]; // @[Modules.scala 65:57:@34878.4]
  assign buffer_14_577 = $signed(_T_79693); // @[Modules.scala 65:57:@34879.4]
  assign _T_79722 = $signed(buffer_0_390) + $signed(11'sh0); // @[Modules.scala 65:57:@34917.4]
  assign _T_79723 = _T_79722[10:0]; // @[Modules.scala 65:57:@34918.4]
  assign buffer_14_587 = $signed(_T_79723); // @[Modules.scala 65:57:@34919.4]
  assign _T_79725 = $signed(buffer_14_392) + $signed(buffer_7_393); // @[Modules.scala 68:83:@34921.4]
  assign _T_79726 = _T_79725[10:0]; // @[Modules.scala 68:83:@34922.4]
  assign buffer_14_588 = $signed(_T_79726); // @[Modules.scala 68:83:@34923.4]
  assign _T_79728 = $signed(buffer_14_394) + $signed(buffer_0_395); // @[Modules.scala 68:83:@34925.4]
  assign _T_79729 = _T_79728[10:0]; // @[Modules.scala 68:83:@34926.4]
  assign buffer_14_589 = $signed(_T_79729); // @[Modules.scala 68:83:@34927.4]
  assign _T_79731 = $signed(buffer_2_396) + $signed(buffer_7_397); // @[Modules.scala 68:83:@34929.4]
  assign _T_79732 = _T_79731[10:0]; // @[Modules.scala 68:83:@34930.4]
  assign buffer_14_590 = $signed(_T_79732); // @[Modules.scala 68:83:@34931.4]
  assign _T_79734 = $signed(buffer_3_398) + $signed(buffer_14_399); // @[Modules.scala 68:83:@34933.4]
  assign _T_79735 = _T_79734[10:0]; // @[Modules.scala 68:83:@34934.4]
  assign buffer_14_591 = $signed(_T_79735); // @[Modules.scala 68:83:@34935.4]
  assign _T_79737 = $signed(buffer_2_400) + $signed(buffer_0_395); // @[Modules.scala 68:83:@34937.4]
  assign _T_79738 = _T_79737[10:0]; // @[Modules.scala 68:83:@34938.4]
  assign buffer_14_592 = $signed(_T_79738); // @[Modules.scala 68:83:@34939.4]
  assign _T_79740 = $signed(buffer_14_402) + $signed(buffer_4_403); // @[Modules.scala 68:83:@34941.4]
  assign _T_79741 = _T_79740[10:0]; // @[Modules.scala 68:83:@34942.4]
  assign buffer_14_593 = $signed(_T_79741); // @[Modules.scala 68:83:@34943.4]
  assign _T_79743 = $signed(buffer_0_395) + $signed(buffer_14_405); // @[Modules.scala 68:83:@34945.4]
  assign _T_79744 = _T_79743[10:0]; // @[Modules.scala 68:83:@34946.4]
  assign buffer_14_594 = $signed(_T_79744); // @[Modules.scala 68:83:@34947.4]
  assign _T_79746 = $signed(buffer_11_406) + $signed(buffer_14_407); // @[Modules.scala 68:83:@34949.4]
  assign _T_79747 = _T_79746[10:0]; // @[Modules.scala 68:83:@34950.4]
  assign buffer_14_595 = $signed(_T_79747); // @[Modules.scala 68:83:@34951.4]
  assign _T_79755 = $signed(buffer_3_412) + $signed(buffer_14_413); // @[Modules.scala 68:83:@34961.4]
  assign _T_79756 = _T_79755[10:0]; // @[Modules.scala 68:83:@34962.4]
  assign buffer_14_598 = $signed(_T_79756); // @[Modules.scala 68:83:@34963.4]
  assign _T_79758 = $signed(buffer_14_414) + $signed(buffer_1_415); // @[Modules.scala 68:83:@34965.4]
  assign _T_79759 = _T_79758[10:0]; // @[Modules.scala 68:83:@34966.4]
  assign buffer_14_599 = $signed(_T_79759); // @[Modules.scala 68:83:@34967.4]
  assign _T_79761 = $signed(buffer_14_416) + $signed(buffer_0_395); // @[Modules.scala 68:83:@34969.4]
  assign _T_79762 = _T_79761[10:0]; // @[Modules.scala 68:83:@34970.4]
  assign buffer_14_600 = $signed(_T_79762); // @[Modules.scala 68:83:@34971.4]
  assign _T_79764 = $signed(buffer_0_395) + $signed(buffer_6_419); // @[Modules.scala 68:83:@34973.4]
  assign _T_79765 = _T_79764[10:0]; // @[Modules.scala 68:83:@34974.4]
  assign buffer_14_601 = $signed(_T_79765); // @[Modules.scala 68:83:@34975.4]
  assign _T_79767 = $signed(buffer_14_420) + $signed(buffer_5_421); // @[Modules.scala 68:83:@34977.4]
  assign _T_79768 = _T_79767[10:0]; // @[Modules.scala 68:83:@34978.4]
  assign buffer_14_602 = $signed(_T_79768); // @[Modules.scala 68:83:@34979.4]
  assign _T_79770 = $signed(buffer_3_422) + $signed(buffer_14_423); // @[Modules.scala 68:83:@34981.4]
  assign _T_79771 = _T_79770[10:0]; // @[Modules.scala 68:83:@34982.4]
  assign buffer_14_603 = $signed(_T_79771); // @[Modules.scala 68:83:@34983.4]
  assign _T_79773 = $signed(buffer_2_424) + $signed(buffer_0_395); // @[Modules.scala 68:83:@34985.4]
  assign _T_79774 = _T_79773[10:0]; // @[Modules.scala 68:83:@34986.4]
  assign buffer_14_604 = $signed(_T_79774); // @[Modules.scala 68:83:@34987.4]
  assign _T_79776 = $signed(buffer_10_426) + $signed(buffer_14_427); // @[Modules.scala 68:83:@34989.4]
  assign _T_79777 = _T_79776[10:0]; // @[Modules.scala 68:83:@34990.4]
  assign buffer_14_605 = $signed(_T_79777); // @[Modules.scala 68:83:@34991.4]
  assign _T_79779 = $signed(buffer_0_428) + $signed(buffer_3_429); // @[Modules.scala 68:83:@34993.4]
  assign _T_79780 = _T_79779[10:0]; // @[Modules.scala 68:83:@34994.4]
  assign buffer_14_606 = $signed(_T_79780); // @[Modules.scala 68:83:@34995.4]
  assign _T_79785 = $signed(buffer_0_395) + $signed(buffer_5_433); // @[Modules.scala 68:83:@35001.4]
  assign _T_79786 = _T_79785[10:0]; // @[Modules.scala 68:83:@35002.4]
  assign buffer_14_608 = $signed(_T_79786); // @[Modules.scala 68:83:@35003.4]
  assign _T_79788 = $signed(buffer_1_434) + $signed(buffer_0_395); // @[Modules.scala 68:83:@35005.4]
  assign _T_79789 = _T_79788[10:0]; // @[Modules.scala 68:83:@35006.4]
  assign buffer_14_609 = $signed(_T_79789); // @[Modules.scala 68:83:@35007.4]
  assign _T_79791 = $signed(buffer_14_436) + $signed(buffer_5_437); // @[Modules.scala 68:83:@35009.4]
  assign _T_79792 = _T_79791[10:0]; // @[Modules.scala 68:83:@35010.4]
  assign buffer_14_610 = $signed(_T_79792); // @[Modules.scala 68:83:@35011.4]
  assign _T_79794 = $signed(buffer_14_438) + $signed(buffer_14_439); // @[Modules.scala 68:83:@35013.4]
  assign _T_79795 = _T_79794[10:0]; // @[Modules.scala 68:83:@35014.4]
  assign buffer_14_611 = $signed(_T_79795); // @[Modules.scala 68:83:@35015.4]
  assign _T_79800 = $signed(buffer_0_395) + $signed(buffer_5_443); // @[Modules.scala 68:83:@35021.4]
  assign _T_79801 = _T_79800[10:0]; // @[Modules.scala 68:83:@35022.4]
  assign buffer_14_613 = $signed(_T_79801); // @[Modules.scala 68:83:@35023.4]
  assign _T_79803 = $signed(buffer_5_444) + $signed(buffer_3_445); // @[Modules.scala 68:83:@35025.4]
  assign _T_79804 = _T_79803[10:0]; // @[Modules.scala 68:83:@35026.4]
  assign buffer_14_614 = $signed(_T_79804); // @[Modules.scala 68:83:@35027.4]
  assign _T_79806 = $signed(buffer_1_446) + $signed(buffer_2_447); // @[Modules.scala 68:83:@35029.4]
  assign _T_79807 = _T_79806[10:0]; // @[Modules.scala 68:83:@35030.4]
  assign buffer_14_615 = $signed(_T_79807); // @[Modules.scala 68:83:@35031.4]
  assign _T_79812 = $signed(buffer_0_395) + $signed(buffer_3_451); // @[Modules.scala 68:83:@35037.4]
  assign _T_79813 = _T_79812[10:0]; // @[Modules.scala 68:83:@35038.4]
  assign buffer_14_617 = $signed(_T_79813); // @[Modules.scala 68:83:@35039.4]
  assign _T_79815 = $signed(buffer_14_452) + $signed(buffer_4_453); // @[Modules.scala 68:83:@35041.4]
  assign _T_79816 = _T_79815[10:0]; // @[Modules.scala 68:83:@35042.4]
  assign buffer_14_618 = $signed(_T_79816); // @[Modules.scala 68:83:@35043.4]
  assign _T_79824 = $signed(buffer_11_458) + $signed(buffer_14_459); // @[Modules.scala 68:83:@35053.4]
  assign _T_79825 = _T_79824[10:0]; // @[Modules.scala 68:83:@35054.4]
  assign buffer_14_621 = $signed(_T_79825); // @[Modules.scala 68:83:@35055.4]
  assign _T_79827 = $signed(buffer_14_460) + $signed(buffer_14_461); // @[Modules.scala 68:83:@35057.4]
  assign _T_79828 = _T_79827[10:0]; // @[Modules.scala 68:83:@35058.4]
  assign buffer_14_622 = $signed(_T_79828); // @[Modules.scala 68:83:@35059.4]
  assign _T_79833 = $signed(buffer_2_464) + $signed(buffer_7_465); // @[Modules.scala 68:83:@35065.4]
  assign _T_79834 = _T_79833[10:0]; // @[Modules.scala 68:83:@35066.4]
  assign buffer_14_624 = $signed(_T_79834); // @[Modules.scala 68:83:@35067.4]
  assign _T_79836 = $signed(buffer_12_466) + $signed(buffer_9_467); // @[Modules.scala 68:83:@35069.4]
  assign _T_79837 = _T_79836[10:0]; // @[Modules.scala 68:83:@35070.4]
  assign buffer_14_625 = $signed(_T_79837); // @[Modules.scala 68:83:@35071.4]
  assign _T_79845 = $signed(buffer_4_472) + $signed(buffer_12_473); // @[Modules.scala 68:83:@35081.4]
  assign _T_79846 = _T_79845[10:0]; // @[Modules.scala 68:83:@35082.4]
  assign buffer_14_628 = $signed(_T_79846); // @[Modules.scala 68:83:@35083.4]
  assign _T_79848 = $signed(buffer_14_474) + $signed(buffer_1_475); // @[Modules.scala 68:83:@35085.4]
  assign _T_79849 = _T_79848[10:0]; // @[Modules.scala 68:83:@35086.4]
  assign buffer_14_629 = $signed(_T_79849); // @[Modules.scala 68:83:@35087.4]
  assign _T_79851 = $signed(buffer_0_395) + $signed(buffer_14_477); // @[Modules.scala 68:83:@35089.4]
  assign _T_79852 = _T_79851[10:0]; // @[Modules.scala 68:83:@35090.4]
  assign buffer_14_630 = $signed(_T_79852); // @[Modules.scala 68:83:@35091.4]
  assign _T_79854 = $signed(buffer_14_478) + $signed(buffer_0_479); // @[Modules.scala 68:83:@35093.4]
  assign _T_79855 = _T_79854[10:0]; // @[Modules.scala 68:83:@35094.4]
  assign buffer_14_631 = $signed(_T_79855); // @[Modules.scala 68:83:@35095.4]
  assign _T_79860 = $signed(buffer_14_482) + $signed(buffer_4_483); // @[Modules.scala 68:83:@35101.4]
  assign _T_79861 = _T_79860[10:0]; // @[Modules.scala 68:83:@35102.4]
  assign buffer_14_633 = $signed(_T_79861); // @[Modules.scala 68:83:@35103.4]
  assign _T_79863 = $signed(buffer_14_484) + $signed(buffer_14_485); // @[Modules.scala 68:83:@35105.4]
  assign _T_79864 = _T_79863[10:0]; // @[Modules.scala 68:83:@35106.4]
  assign buffer_14_634 = $signed(_T_79864); // @[Modules.scala 68:83:@35107.4]
  assign _T_79866 = $signed(buffer_8_486) + $signed(buffer_4_487); // @[Modules.scala 68:83:@35109.4]
  assign _T_79867 = _T_79866[10:0]; // @[Modules.scala 68:83:@35110.4]
  assign buffer_14_635 = $signed(_T_79867); // @[Modules.scala 68:83:@35111.4]
  assign _T_79869 = $signed(buffer_14_488) + $signed(buffer_3_489); // @[Modules.scala 68:83:@35113.4]
  assign _T_79870 = _T_79869[10:0]; // @[Modules.scala 68:83:@35114.4]
  assign buffer_14_636 = $signed(_T_79870); // @[Modules.scala 68:83:@35115.4]
  assign _T_79875 = $signed(buffer_4_492) + $signed(buffer_0_493); // @[Modules.scala 68:83:@35121.4]
  assign _T_79876 = _T_79875[10:0]; // @[Modules.scala 68:83:@35122.4]
  assign buffer_14_638 = $signed(_T_79876); // @[Modules.scala 68:83:@35123.4]
  assign _T_79878 = $signed(buffer_13_494) + $signed(buffer_0_395); // @[Modules.scala 68:83:@35125.4]
  assign _T_79879 = _T_79878[10:0]; // @[Modules.scala 68:83:@35126.4]
  assign buffer_14_639 = $signed(_T_79879); // @[Modules.scala 68:83:@35127.4]
  assign _T_79881 = $signed(buffer_14_496) + $signed(buffer_0_395); // @[Modules.scala 68:83:@35129.4]
  assign _T_79882 = _T_79881[10:0]; // @[Modules.scala 68:83:@35130.4]
  assign buffer_14_640 = $signed(_T_79882); // @[Modules.scala 68:83:@35131.4]
  assign _T_79884 = $signed(buffer_3_498) + $signed(buffer_14_499); // @[Modules.scala 68:83:@35133.4]
  assign _T_79885 = _T_79884[10:0]; // @[Modules.scala 68:83:@35134.4]
  assign buffer_14_641 = $signed(_T_79885); // @[Modules.scala 68:83:@35135.4]
  assign _T_79887 = $signed(buffer_14_500) + $signed(buffer_14_501); // @[Modules.scala 68:83:@35137.4]
  assign _T_79888 = _T_79887[10:0]; // @[Modules.scala 68:83:@35138.4]
  assign buffer_14_642 = $signed(_T_79888); // @[Modules.scala 68:83:@35139.4]
  assign _T_79890 = $signed(buffer_0_395) + $signed(buffer_8_503); // @[Modules.scala 68:83:@35141.4]
  assign _T_79891 = _T_79890[10:0]; // @[Modules.scala 68:83:@35142.4]
  assign buffer_14_643 = $signed(_T_79891); // @[Modules.scala 68:83:@35143.4]
  assign _T_79893 = $signed(buffer_1_504) + $signed(buffer_5_505); // @[Modules.scala 68:83:@35145.4]
  assign _T_79894 = _T_79893[10:0]; // @[Modules.scala 68:83:@35146.4]
  assign buffer_14_644 = $signed(_T_79894); // @[Modules.scala 68:83:@35147.4]
  assign _T_79899 = $signed(buffer_14_508) + $signed(buffer_14_509); // @[Modules.scala 68:83:@35153.4]
  assign _T_79900 = _T_79899[10:0]; // @[Modules.scala 68:83:@35154.4]
  assign buffer_14_646 = $signed(_T_79900); // @[Modules.scala 68:83:@35155.4]
  assign _T_79902 = $signed(buffer_14_510) + $signed(buffer_14_511); // @[Modules.scala 68:83:@35157.4]
  assign _T_79903 = _T_79902[10:0]; // @[Modules.scala 68:83:@35158.4]
  assign buffer_14_647 = $signed(_T_79903); // @[Modules.scala 68:83:@35159.4]
  assign _T_79908 = $signed(buffer_14_514) + $signed(buffer_10_515); // @[Modules.scala 68:83:@35165.4]
  assign _T_79909 = _T_79908[10:0]; // @[Modules.scala 68:83:@35166.4]
  assign buffer_14_649 = $signed(_T_79909); // @[Modules.scala 68:83:@35167.4]
  assign _T_79911 = $signed(buffer_14_516) + $signed(buffer_3_517); // @[Modules.scala 68:83:@35169.4]
  assign _T_79912 = _T_79911[10:0]; // @[Modules.scala 68:83:@35170.4]
  assign buffer_14_650 = $signed(_T_79912); // @[Modules.scala 68:83:@35171.4]
  assign _T_79914 = $signed(buffer_14_518) + $signed(buffer_3_519); // @[Modules.scala 68:83:@35173.4]
  assign _T_79915 = _T_79914[10:0]; // @[Modules.scala 68:83:@35174.4]
  assign buffer_14_651 = $signed(_T_79915); // @[Modules.scala 68:83:@35175.4]
  assign _T_79917 = $signed(buffer_10_520) + $signed(buffer_14_521); // @[Modules.scala 68:83:@35177.4]
  assign _T_79918 = _T_79917[10:0]; // @[Modules.scala 68:83:@35178.4]
  assign buffer_14_652 = $signed(_T_79918); // @[Modules.scala 68:83:@35179.4]
  assign _T_79920 = $signed(buffer_7_522) + $signed(buffer_4_523); // @[Modules.scala 68:83:@35181.4]
  assign _T_79921 = _T_79920[10:0]; // @[Modules.scala 68:83:@35182.4]
  assign buffer_14_653 = $signed(_T_79921); // @[Modules.scala 68:83:@35183.4]
  assign _T_79923 = $signed(buffer_13_524) + $signed(buffer_14_525); // @[Modules.scala 68:83:@35185.4]
  assign _T_79924 = _T_79923[10:0]; // @[Modules.scala 68:83:@35186.4]
  assign buffer_14_654 = $signed(_T_79924); // @[Modules.scala 68:83:@35187.4]
  assign _T_79926 = $signed(buffer_1_526) + $signed(buffer_14_527); // @[Modules.scala 68:83:@35189.4]
  assign _T_79927 = _T_79926[10:0]; // @[Modules.scala 68:83:@35190.4]
  assign buffer_14_655 = $signed(_T_79927); // @[Modules.scala 68:83:@35191.4]
  assign _T_79929 = $signed(buffer_0_395) + $signed(buffer_1_529); // @[Modules.scala 68:83:@35193.4]
  assign _T_79930 = _T_79929[10:0]; // @[Modules.scala 68:83:@35194.4]
  assign buffer_14_656 = $signed(_T_79930); // @[Modules.scala 68:83:@35195.4]
  assign _T_79935 = $signed(buffer_14_532) + $signed(buffer_3_533); // @[Modules.scala 68:83:@35201.4]
  assign _T_79936 = _T_79935[10:0]; // @[Modules.scala 68:83:@35202.4]
  assign buffer_14_658 = $signed(_T_79936); // @[Modules.scala 68:83:@35203.4]
  assign _T_79938 = $signed(buffer_14_534) + $signed(buffer_0_395); // @[Modules.scala 68:83:@35205.4]
  assign _T_79939 = _T_79938[10:0]; // @[Modules.scala 68:83:@35206.4]
  assign buffer_14_659 = $signed(_T_79939); // @[Modules.scala 68:83:@35207.4]
  assign _T_79941 = $signed(buffer_14_536) + $signed(buffer_4_537); // @[Modules.scala 68:83:@35209.4]
  assign _T_79942 = _T_79941[10:0]; // @[Modules.scala 68:83:@35210.4]
  assign buffer_14_660 = $signed(_T_79942); // @[Modules.scala 68:83:@35211.4]
  assign _T_79944 = $signed(buffer_13_538) + $signed(buffer_14_539); // @[Modules.scala 68:83:@35213.4]
  assign _T_79945 = _T_79944[10:0]; // @[Modules.scala 68:83:@35214.4]
  assign buffer_14_661 = $signed(_T_79945); // @[Modules.scala 68:83:@35215.4]
  assign _T_79947 = $signed(buffer_3_540) + $signed(buffer_5_541); // @[Modules.scala 68:83:@35217.4]
  assign _T_79948 = _T_79947[10:0]; // @[Modules.scala 68:83:@35218.4]
  assign buffer_14_662 = $signed(_T_79948); // @[Modules.scala 68:83:@35219.4]
  assign _T_79950 = $signed(buffer_0_395) + $signed(buffer_14_543); // @[Modules.scala 68:83:@35221.4]
  assign _T_79951 = _T_79950[10:0]; // @[Modules.scala 68:83:@35222.4]
  assign buffer_14_663 = $signed(_T_79951); // @[Modules.scala 68:83:@35223.4]
  assign _T_79956 = $signed(buffer_14_546) + $signed(buffer_14_547); // @[Modules.scala 68:83:@35229.4]
  assign _T_79957 = _T_79956[10:0]; // @[Modules.scala 68:83:@35230.4]
  assign buffer_14_665 = $signed(_T_79957); // @[Modules.scala 68:83:@35231.4]
  assign _T_79965 = $signed(buffer_14_552) + $signed(buffer_1_553); // @[Modules.scala 68:83:@35241.4]
  assign _T_79966 = _T_79965[10:0]; // @[Modules.scala 68:83:@35242.4]
  assign buffer_14_668 = $signed(_T_79966); // @[Modules.scala 68:83:@35243.4]
  assign _T_79968 = $signed(buffer_4_554) + $signed(buffer_14_555); // @[Modules.scala 68:83:@35245.4]
  assign _T_79969 = _T_79968[10:0]; // @[Modules.scala 68:83:@35246.4]
  assign buffer_14_669 = $signed(_T_79969); // @[Modules.scala 68:83:@35247.4]
  assign _T_79977 = $signed(buffer_1_560) + $signed(buffer_8_561); // @[Modules.scala 68:83:@35257.4]
  assign _T_79978 = _T_79977[10:0]; // @[Modules.scala 68:83:@35258.4]
  assign buffer_14_672 = $signed(_T_79978); // @[Modules.scala 68:83:@35259.4]
  assign _T_79980 = $signed(buffer_5_562) + $signed(buffer_4_563); // @[Modules.scala 68:83:@35261.4]
  assign _T_79981 = _T_79980[10:0]; // @[Modules.scala 68:83:@35262.4]
  assign buffer_14_673 = $signed(_T_79981); // @[Modules.scala 68:83:@35263.4]
  assign _T_79986 = $signed(buffer_14_566) + $signed(buffer_2_567); // @[Modules.scala 68:83:@35269.4]
  assign _T_79987 = _T_79986[10:0]; // @[Modules.scala 68:83:@35270.4]
  assign buffer_14_675 = $signed(_T_79987); // @[Modules.scala 68:83:@35271.4]
  assign _T_79989 = $signed(buffer_14_568) + $signed(buffer_14_569); // @[Modules.scala 68:83:@35273.4]
  assign _T_79990 = _T_79989[10:0]; // @[Modules.scala 68:83:@35274.4]
  assign buffer_14_676 = $signed(_T_79990); // @[Modules.scala 68:83:@35275.4]
  assign _T_79992 = $signed(buffer_14_570) + $signed(buffer_0_571); // @[Modules.scala 68:83:@35277.4]
  assign _T_79993 = _T_79992[10:0]; // @[Modules.scala 68:83:@35278.4]
  assign buffer_14_677 = $signed(_T_79993); // @[Modules.scala 68:83:@35279.4]
  assign _T_79995 = $signed(buffer_0_572) + $signed(buffer_14_573); // @[Modules.scala 68:83:@35281.4]
  assign _T_79996 = _T_79995[10:0]; // @[Modules.scala 68:83:@35282.4]
  assign buffer_14_678 = $signed(_T_79996); // @[Modules.scala 68:83:@35283.4]
  assign _T_79998 = $signed(buffer_14_574) + $signed(buffer_14_575); // @[Modules.scala 68:83:@35285.4]
  assign _T_79999 = _T_79998[10:0]; // @[Modules.scala 68:83:@35286.4]
  assign buffer_14_679 = $signed(_T_79999); // @[Modules.scala 68:83:@35287.4]
  assign _T_80001 = $signed(buffer_14_576) + $signed(buffer_14_577); // @[Modules.scala 68:83:@35289.4]
  assign _T_80002 = _T_80001[10:0]; // @[Modules.scala 68:83:@35290.4]
  assign buffer_14_680 = $signed(_T_80002); // @[Modules.scala 68:83:@35291.4]
  assign _T_80004 = $signed(buffer_3_578) + $signed(buffer_9_579); // @[Modules.scala 68:83:@35293.4]
  assign _T_80005 = _T_80004[10:0]; // @[Modules.scala 68:83:@35294.4]
  assign buffer_14_681 = $signed(_T_80005); // @[Modules.scala 68:83:@35295.4]
  assign _T_80007 = $signed(buffer_12_580) + $signed(buffer_10_581); // @[Modules.scala 68:83:@35297.4]
  assign _T_80008 = _T_80007[10:0]; // @[Modules.scala 68:83:@35298.4]
  assign buffer_14_682 = $signed(_T_80008); // @[Modules.scala 68:83:@35299.4]
  assign _T_80010 = $signed(buffer_1_582) + $signed(buffer_5_583); // @[Modules.scala 68:83:@35301.4]
  assign _T_80011 = _T_80010[10:0]; // @[Modules.scala 68:83:@35302.4]
  assign buffer_14_683 = $signed(_T_80011); // @[Modules.scala 68:83:@35303.4]
  assign _T_80016 = $signed(buffer_0_395) + $signed(buffer_14_587); // @[Modules.scala 68:83:@35309.4]
  assign _T_80017 = _T_80016[10:0]; // @[Modules.scala 68:83:@35310.4]
  assign buffer_14_685 = $signed(_T_80017); // @[Modules.scala 68:83:@35311.4]
  assign _T_80019 = $signed(buffer_14_588) + $signed(buffer_14_589); // @[Modules.scala 71:109:@35313.4]
  assign _T_80020 = _T_80019[10:0]; // @[Modules.scala 71:109:@35314.4]
  assign buffer_14_686 = $signed(_T_80020); // @[Modules.scala 71:109:@35315.4]
  assign _T_80022 = $signed(buffer_14_590) + $signed(buffer_14_591); // @[Modules.scala 71:109:@35317.4]
  assign _T_80023 = _T_80022[10:0]; // @[Modules.scala 71:109:@35318.4]
  assign buffer_14_687 = $signed(_T_80023); // @[Modules.scala 71:109:@35319.4]
  assign _T_80025 = $signed(buffer_14_592) + $signed(buffer_14_593); // @[Modules.scala 71:109:@35321.4]
  assign _T_80026 = _T_80025[10:0]; // @[Modules.scala 71:109:@35322.4]
  assign buffer_14_688 = $signed(_T_80026); // @[Modules.scala 71:109:@35323.4]
  assign _T_80028 = $signed(buffer_14_594) + $signed(buffer_14_595); // @[Modules.scala 71:109:@35325.4]
  assign _T_80029 = _T_80028[10:0]; // @[Modules.scala 71:109:@35326.4]
  assign buffer_14_689 = $signed(_T_80029); // @[Modules.scala 71:109:@35327.4]
  assign _T_80034 = $signed(buffer_14_598) + $signed(buffer_14_599); // @[Modules.scala 71:109:@35333.4]
  assign _T_80035 = _T_80034[10:0]; // @[Modules.scala 71:109:@35334.4]
  assign buffer_14_691 = $signed(_T_80035); // @[Modules.scala 71:109:@35335.4]
  assign _T_80037 = $signed(buffer_14_600) + $signed(buffer_14_601); // @[Modules.scala 71:109:@35337.4]
  assign _T_80038 = _T_80037[10:0]; // @[Modules.scala 71:109:@35338.4]
  assign buffer_14_692 = $signed(_T_80038); // @[Modules.scala 71:109:@35339.4]
  assign _T_80040 = $signed(buffer_14_602) + $signed(buffer_14_603); // @[Modules.scala 71:109:@35341.4]
  assign _T_80041 = _T_80040[10:0]; // @[Modules.scala 71:109:@35342.4]
  assign buffer_14_693 = $signed(_T_80041); // @[Modules.scala 71:109:@35343.4]
  assign _T_80043 = $signed(buffer_14_604) + $signed(buffer_14_605); // @[Modules.scala 71:109:@35345.4]
  assign _T_80044 = _T_80043[10:0]; // @[Modules.scala 71:109:@35346.4]
  assign buffer_14_694 = $signed(_T_80044); // @[Modules.scala 71:109:@35347.4]
  assign _T_80046 = $signed(buffer_14_606) + $signed(buffer_4_607); // @[Modules.scala 71:109:@35349.4]
  assign _T_80047 = _T_80046[10:0]; // @[Modules.scala 71:109:@35350.4]
  assign buffer_14_695 = $signed(_T_80047); // @[Modules.scala 71:109:@35351.4]
  assign _T_80049 = $signed(buffer_14_608) + $signed(buffer_14_609); // @[Modules.scala 71:109:@35353.4]
  assign _T_80050 = _T_80049[10:0]; // @[Modules.scala 71:109:@35354.4]
  assign buffer_14_696 = $signed(_T_80050); // @[Modules.scala 71:109:@35355.4]
  assign _T_80052 = $signed(buffer_14_610) + $signed(buffer_14_611); // @[Modules.scala 71:109:@35357.4]
  assign _T_80053 = _T_80052[10:0]; // @[Modules.scala 71:109:@35358.4]
  assign buffer_14_697 = $signed(_T_80053); // @[Modules.scala 71:109:@35359.4]
  assign _T_80055 = $signed(buffer_4_612) + $signed(buffer_14_613); // @[Modules.scala 71:109:@35361.4]
  assign _T_80056 = _T_80055[10:0]; // @[Modules.scala 71:109:@35362.4]
  assign buffer_14_698 = $signed(_T_80056); // @[Modules.scala 71:109:@35363.4]
  assign _T_80058 = $signed(buffer_14_614) + $signed(buffer_14_615); // @[Modules.scala 71:109:@35365.4]
  assign _T_80059 = _T_80058[10:0]; // @[Modules.scala 71:109:@35366.4]
  assign buffer_14_699 = $signed(_T_80059); // @[Modules.scala 71:109:@35367.4]
  assign _T_80061 = $signed(buffer_11_616) + $signed(buffer_14_617); // @[Modules.scala 71:109:@35369.4]
  assign _T_80062 = _T_80061[10:0]; // @[Modules.scala 71:109:@35370.4]
  assign buffer_14_700 = $signed(_T_80062); // @[Modules.scala 71:109:@35371.4]
  assign _T_80064 = $signed(buffer_14_618) + $signed(buffer_2_619); // @[Modules.scala 71:109:@35373.4]
  assign _T_80065 = _T_80064[10:0]; // @[Modules.scala 71:109:@35374.4]
  assign buffer_14_701 = $signed(_T_80065); // @[Modules.scala 71:109:@35375.4]
  assign _T_80067 = $signed(buffer_0_620) + $signed(buffer_14_621); // @[Modules.scala 71:109:@35377.4]
  assign _T_80068 = _T_80067[10:0]; // @[Modules.scala 71:109:@35378.4]
  assign buffer_14_702 = $signed(_T_80068); // @[Modules.scala 71:109:@35379.4]
  assign _T_80070 = $signed(buffer_14_622) + $signed(buffer_0_593); // @[Modules.scala 71:109:@35381.4]
  assign _T_80071 = _T_80070[10:0]; // @[Modules.scala 71:109:@35382.4]
  assign buffer_14_703 = $signed(_T_80071); // @[Modules.scala 71:109:@35383.4]
  assign _T_80073 = $signed(buffer_14_624) + $signed(buffer_14_625); // @[Modules.scala 71:109:@35385.4]
  assign _T_80074 = _T_80073[10:0]; // @[Modules.scala 71:109:@35386.4]
  assign buffer_14_704 = $signed(_T_80074); // @[Modules.scala 71:109:@35387.4]
  assign _T_80076 = $signed(buffer_1_626) + $signed(buffer_2_627); // @[Modules.scala 71:109:@35389.4]
  assign _T_80077 = _T_80076[10:0]; // @[Modules.scala 71:109:@35390.4]
  assign buffer_14_705 = $signed(_T_80077); // @[Modules.scala 71:109:@35391.4]
  assign _T_80079 = $signed(buffer_14_628) + $signed(buffer_14_629); // @[Modules.scala 71:109:@35393.4]
  assign _T_80080 = _T_80079[10:0]; // @[Modules.scala 71:109:@35394.4]
  assign buffer_14_706 = $signed(_T_80080); // @[Modules.scala 71:109:@35395.4]
  assign _T_80082 = $signed(buffer_14_630) + $signed(buffer_14_631); // @[Modules.scala 71:109:@35397.4]
  assign _T_80083 = _T_80082[10:0]; // @[Modules.scala 71:109:@35398.4]
  assign buffer_14_707 = $signed(_T_80083); // @[Modules.scala 71:109:@35399.4]
  assign _T_80085 = $signed(buffer_13_632) + $signed(buffer_14_633); // @[Modules.scala 71:109:@35401.4]
  assign _T_80086 = _T_80085[10:0]; // @[Modules.scala 71:109:@35402.4]
  assign buffer_14_708 = $signed(_T_80086); // @[Modules.scala 71:109:@35403.4]
  assign _T_80088 = $signed(buffer_14_634) + $signed(buffer_14_635); // @[Modules.scala 71:109:@35405.4]
  assign _T_80089 = _T_80088[10:0]; // @[Modules.scala 71:109:@35406.4]
  assign buffer_14_709 = $signed(_T_80089); // @[Modules.scala 71:109:@35407.4]
  assign _T_80091 = $signed(buffer_14_636) + $signed(buffer_0_593); // @[Modules.scala 71:109:@35409.4]
  assign _T_80092 = _T_80091[10:0]; // @[Modules.scala 71:109:@35410.4]
  assign buffer_14_710 = $signed(_T_80092); // @[Modules.scala 71:109:@35411.4]
  assign _T_80094 = $signed(buffer_14_638) + $signed(buffer_14_639); // @[Modules.scala 71:109:@35413.4]
  assign _T_80095 = _T_80094[10:0]; // @[Modules.scala 71:109:@35414.4]
  assign buffer_14_711 = $signed(_T_80095); // @[Modules.scala 71:109:@35415.4]
  assign _T_80097 = $signed(buffer_14_640) + $signed(buffer_14_641); // @[Modules.scala 71:109:@35417.4]
  assign _T_80098 = _T_80097[10:0]; // @[Modules.scala 71:109:@35418.4]
  assign buffer_14_712 = $signed(_T_80098); // @[Modules.scala 71:109:@35419.4]
  assign _T_80100 = $signed(buffer_14_642) + $signed(buffer_14_643); // @[Modules.scala 71:109:@35421.4]
  assign _T_80101 = _T_80100[10:0]; // @[Modules.scala 71:109:@35422.4]
  assign buffer_14_713 = $signed(_T_80101); // @[Modules.scala 71:109:@35423.4]
  assign _T_80103 = $signed(buffer_14_644) + $signed(buffer_12_645); // @[Modules.scala 71:109:@35425.4]
  assign _T_80104 = _T_80103[10:0]; // @[Modules.scala 71:109:@35426.4]
  assign buffer_14_714 = $signed(_T_80104); // @[Modules.scala 71:109:@35427.4]
  assign _T_80106 = $signed(buffer_14_646) + $signed(buffer_14_647); // @[Modules.scala 71:109:@35429.4]
  assign _T_80107 = _T_80106[10:0]; // @[Modules.scala 71:109:@35430.4]
  assign buffer_14_715 = $signed(_T_80107); // @[Modules.scala 71:109:@35431.4]
  assign _T_80109 = $signed(buffer_8_648) + $signed(buffer_14_649); // @[Modules.scala 71:109:@35433.4]
  assign _T_80110 = _T_80109[10:0]; // @[Modules.scala 71:109:@35434.4]
  assign buffer_14_716 = $signed(_T_80110); // @[Modules.scala 71:109:@35435.4]
  assign _T_80112 = $signed(buffer_14_650) + $signed(buffer_14_651); // @[Modules.scala 71:109:@35437.4]
  assign _T_80113 = _T_80112[10:0]; // @[Modules.scala 71:109:@35438.4]
  assign buffer_14_717 = $signed(_T_80113); // @[Modules.scala 71:109:@35439.4]
  assign _T_80115 = $signed(buffer_14_652) + $signed(buffer_14_653); // @[Modules.scala 71:109:@35441.4]
  assign _T_80116 = _T_80115[10:0]; // @[Modules.scala 71:109:@35442.4]
  assign buffer_14_718 = $signed(_T_80116); // @[Modules.scala 71:109:@35443.4]
  assign _T_80118 = $signed(buffer_14_654) + $signed(buffer_14_655); // @[Modules.scala 71:109:@35445.4]
  assign _T_80119 = _T_80118[10:0]; // @[Modules.scala 71:109:@35446.4]
  assign buffer_14_719 = $signed(_T_80119); // @[Modules.scala 71:109:@35447.4]
  assign _T_80121 = $signed(buffer_14_656) + $signed(buffer_3_657); // @[Modules.scala 71:109:@35449.4]
  assign _T_80122 = _T_80121[10:0]; // @[Modules.scala 71:109:@35450.4]
  assign buffer_14_720 = $signed(_T_80122); // @[Modules.scala 71:109:@35451.4]
  assign _T_80124 = $signed(buffer_14_658) + $signed(buffer_14_659); // @[Modules.scala 71:109:@35453.4]
  assign _T_80125 = _T_80124[10:0]; // @[Modules.scala 71:109:@35454.4]
  assign buffer_14_721 = $signed(_T_80125); // @[Modules.scala 71:109:@35455.4]
  assign _T_80127 = $signed(buffer_14_660) + $signed(buffer_14_661); // @[Modules.scala 71:109:@35457.4]
  assign _T_80128 = _T_80127[10:0]; // @[Modules.scala 71:109:@35458.4]
  assign buffer_14_722 = $signed(_T_80128); // @[Modules.scala 71:109:@35459.4]
  assign _T_80130 = $signed(buffer_14_662) + $signed(buffer_14_663); // @[Modules.scala 71:109:@35461.4]
  assign _T_80131 = _T_80130[10:0]; // @[Modules.scala 71:109:@35462.4]
  assign buffer_14_723 = $signed(_T_80131); // @[Modules.scala 71:109:@35463.4]
  assign _T_80133 = $signed(buffer_12_664) + $signed(buffer_14_665); // @[Modules.scala 71:109:@35465.4]
  assign _T_80134 = _T_80133[10:0]; // @[Modules.scala 71:109:@35466.4]
  assign buffer_14_724 = $signed(_T_80134); // @[Modules.scala 71:109:@35467.4]
  assign _T_80136 = $signed(buffer_1_666) + $signed(buffer_4_667); // @[Modules.scala 71:109:@35469.4]
  assign _T_80137 = _T_80136[10:0]; // @[Modules.scala 71:109:@35470.4]
  assign buffer_14_725 = $signed(_T_80137); // @[Modules.scala 71:109:@35471.4]
  assign _T_80139 = $signed(buffer_14_668) + $signed(buffer_14_669); // @[Modules.scala 71:109:@35473.4]
  assign _T_80140 = _T_80139[10:0]; // @[Modules.scala 71:109:@35474.4]
  assign buffer_14_726 = $signed(_T_80140); // @[Modules.scala 71:109:@35475.4]
  assign _T_80142 = $signed(buffer_11_670) + $signed(buffer_0_671); // @[Modules.scala 71:109:@35477.4]
  assign _T_80143 = _T_80142[10:0]; // @[Modules.scala 71:109:@35478.4]
  assign buffer_14_727 = $signed(_T_80143); // @[Modules.scala 71:109:@35479.4]
  assign _T_80145 = $signed(buffer_14_672) + $signed(buffer_14_673); // @[Modules.scala 71:109:@35481.4]
  assign _T_80146 = _T_80145[10:0]; // @[Modules.scala 71:109:@35482.4]
  assign buffer_14_728 = $signed(_T_80146); // @[Modules.scala 71:109:@35483.4]
  assign _T_80148 = $signed(buffer_0_674) + $signed(buffer_14_675); // @[Modules.scala 71:109:@35485.4]
  assign _T_80149 = _T_80148[10:0]; // @[Modules.scala 71:109:@35486.4]
  assign buffer_14_729 = $signed(_T_80149); // @[Modules.scala 71:109:@35487.4]
  assign _T_80151 = $signed(buffer_14_676) + $signed(buffer_14_677); // @[Modules.scala 71:109:@35489.4]
  assign _T_80152 = _T_80151[10:0]; // @[Modules.scala 71:109:@35490.4]
  assign buffer_14_730 = $signed(_T_80152); // @[Modules.scala 71:109:@35491.4]
  assign _T_80154 = $signed(buffer_14_678) + $signed(buffer_14_679); // @[Modules.scala 71:109:@35493.4]
  assign _T_80155 = _T_80154[10:0]; // @[Modules.scala 71:109:@35494.4]
  assign buffer_14_731 = $signed(_T_80155); // @[Modules.scala 71:109:@35495.4]
  assign _T_80157 = $signed(buffer_14_680) + $signed(buffer_14_681); // @[Modules.scala 71:109:@35497.4]
  assign _T_80158 = _T_80157[10:0]; // @[Modules.scala 71:109:@35498.4]
  assign buffer_14_732 = $signed(_T_80158); // @[Modules.scala 71:109:@35499.4]
  assign _T_80160 = $signed(buffer_14_682) + $signed(buffer_14_683); // @[Modules.scala 71:109:@35501.4]
  assign _T_80161 = _T_80160[10:0]; // @[Modules.scala 71:109:@35502.4]
  assign buffer_14_733 = $signed(_T_80161); // @[Modules.scala 71:109:@35503.4]
  assign _T_80163 = $signed(buffer_0_593) + $signed(buffer_14_685); // @[Modules.scala 71:109:@35505.4]
  assign _T_80164 = _T_80163[10:0]; // @[Modules.scala 71:109:@35506.4]
  assign buffer_14_734 = $signed(_T_80164); // @[Modules.scala 71:109:@35507.4]
  assign _T_80166 = $signed(buffer_14_686) + $signed(buffer_14_687); // @[Modules.scala 78:156:@35510.4]
  assign _T_80167 = _T_80166[10:0]; // @[Modules.scala 78:156:@35511.4]
  assign buffer_14_736 = $signed(_T_80167); // @[Modules.scala 78:156:@35512.4]
  assign _T_80169 = $signed(buffer_14_736) + $signed(buffer_14_688); // @[Modules.scala 78:156:@35514.4]
  assign _T_80170 = _T_80169[10:0]; // @[Modules.scala 78:156:@35515.4]
  assign buffer_14_737 = $signed(_T_80170); // @[Modules.scala 78:156:@35516.4]
  assign _T_80172 = $signed(buffer_14_737) + $signed(buffer_14_689); // @[Modules.scala 78:156:@35518.4]
  assign _T_80173 = _T_80172[10:0]; // @[Modules.scala 78:156:@35519.4]
  assign buffer_14_738 = $signed(_T_80173); // @[Modules.scala 78:156:@35520.4]
  assign _T_80175 = $signed(buffer_14_738) + $signed(buffer_0_701); // @[Modules.scala 78:156:@35522.4]
  assign _T_80176 = _T_80175[10:0]; // @[Modules.scala 78:156:@35523.4]
  assign buffer_14_739 = $signed(_T_80176); // @[Modules.scala 78:156:@35524.4]
  assign _T_80178 = $signed(buffer_14_739) + $signed(buffer_14_691); // @[Modules.scala 78:156:@35526.4]
  assign _T_80179 = _T_80178[10:0]; // @[Modules.scala 78:156:@35527.4]
  assign buffer_14_740 = $signed(_T_80179); // @[Modules.scala 78:156:@35528.4]
  assign _T_80181 = $signed(buffer_14_740) + $signed(buffer_14_692); // @[Modules.scala 78:156:@35530.4]
  assign _T_80182 = _T_80181[10:0]; // @[Modules.scala 78:156:@35531.4]
  assign buffer_14_741 = $signed(_T_80182); // @[Modules.scala 78:156:@35532.4]
  assign _T_80184 = $signed(buffer_14_741) + $signed(buffer_14_693); // @[Modules.scala 78:156:@35534.4]
  assign _T_80185 = _T_80184[10:0]; // @[Modules.scala 78:156:@35535.4]
  assign buffer_14_742 = $signed(_T_80185); // @[Modules.scala 78:156:@35536.4]
  assign _T_80187 = $signed(buffer_14_742) + $signed(buffer_14_694); // @[Modules.scala 78:156:@35538.4]
  assign _T_80188 = _T_80187[10:0]; // @[Modules.scala 78:156:@35539.4]
  assign buffer_14_743 = $signed(_T_80188); // @[Modules.scala 78:156:@35540.4]
  assign _T_80190 = $signed(buffer_14_743) + $signed(buffer_14_695); // @[Modules.scala 78:156:@35542.4]
  assign _T_80191 = _T_80190[10:0]; // @[Modules.scala 78:156:@35543.4]
  assign buffer_14_744 = $signed(_T_80191); // @[Modules.scala 78:156:@35544.4]
  assign _T_80193 = $signed(buffer_14_744) + $signed(buffer_14_696); // @[Modules.scala 78:156:@35546.4]
  assign _T_80194 = _T_80193[10:0]; // @[Modules.scala 78:156:@35547.4]
  assign buffer_14_745 = $signed(_T_80194); // @[Modules.scala 78:156:@35548.4]
  assign _T_80196 = $signed(buffer_14_745) + $signed(buffer_14_697); // @[Modules.scala 78:156:@35550.4]
  assign _T_80197 = _T_80196[10:0]; // @[Modules.scala 78:156:@35551.4]
  assign buffer_14_746 = $signed(_T_80197); // @[Modules.scala 78:156:@35552.4]
  assign _T_80199 = $signed(buffer_14_746) + $signed(buffer_14_698); // @[Modules.scala 78:156:@35554.4]
  assign _T_80200 = _T_80199[10:0]; // @[Modules.scala 78:156:@35555.4]
  assign buffer_14_747 = $signed(_T_80200); // @[Modules.scala 78:156:@35556.4]
  assign _T_80202 = $signed(buffer_14_747) + $signed(buffer_14_699); // @[Modules.scala 78:156:@35558.4]
  assign _T_80203 = _T_80202[10:0]; // @[Modules.scala 78:156:@35559.4]
  assign buffer_14_748 = $signed(_T_80203); // @[Modules.scala 78:156:@35560.4]
  assign _T_80205 = $signed(buffer_14_748) + $signed(buffer_14_700); // @[Modules.scala 78:156:@35562.4]
  assign _T_80206 = _T_80205[10:0]; // @[Modules.scala 78:156:@35563.4]
  assign buffer_14_749 = $signed(_T_80206); // @[Modules.scala 78:156:@35564.4]
  assign _T_80208 = $signed(buffer_14_749) + $signed(buffer_14_701); // @[Modules.scala 78:156:@35566.4]
  assign _T_80209 = _T_80208[10:0]; // @[Modules.scala 78:156:@35567.4]
  assign buffer_14_750 = $signed(_T_80209); // @[Modules.scala 78:156:@35568.4]
  assign _T_80211 = $signed(buffer_14_750) + $signed(buffer_14_702); // @[Modules.scala 78:156:@35570.4]
  assign _T_80212 = _T_80211[10:0]; // @[Modules.scala 78:156:@35571.4]
  assign buffer_14_751 = $signed(_T_80212); // @[Modules.scala 78:156:@35572.4]
  assign _T_80214 = $signed(buffer_14_751) + $signed(buffer_14_703); // @[Modules.scala 78:156:@35574.4]
  assign _T_80215 = _T_80214[10:0]; // @[Modules.scala 78:156:@35575.4]
  assign buffer_14_752 = $signed(_T_80215); // @[Modules.scala 78:156:@35576.4]
  assign _T_80217 = $signed(buffer_14_752) + $signed(buffer_14_704); // @[Modules.scala 78:156:@35578.4]
  assign _T_80218 = _T_80217[10:0]; // @[Modules.scala 78:156:@35579.4]
  assign buffer_14_753 = $signed(_T_80218); // @[Modules.scala 78:156:@35580.4]
  assign _T_80220 = $signed(buffer_14_753) + $signed(buffer_14_705); // @[Modules.scala 78:156:@35582.4]
  assign _T_80221 = _T_80220[10:0]; // @[Modules.scala 78:156:@35583.4]
  assign buffer_14_754 = $signed(_T_80221); // @[Modules.scala 78:156:@35584.4]
  assign _T_80223 = $signed(buffer_14_754) + $signed(buffer_14_706); // @[Modules.scala 78:156:@35586.4]
  assign _T_80224 = _T_80223[10:0]; // @[Modules.scala 78:156:@35587.4]
  assign buffer_14_755 = $signed(_T_80224); // @[Modules.scala 78:156:@35588.4]
  assign _T_80226 = $signed(buffer_14_755) + $signed(buffer_14_707); // @[Modules.scala 78:156:@35590.4]
  assign _T_80227 = _T_80226[10:0]; // @[Modules.scala 78:156:@35591.4]
  assign buffer_14_756 = $signed(_T_80227); // @[Modules.scala 78:156:@35592.4]
  assign _T_80229 = $signed(buffer_14_756) + $signed(buffer_14_708); // @[Modules.scala 78:156:@35594.4]
  assign _T_80230 = _T_80229[10:0]; // @[Modules.scala 78:156:@35595.4]
  assign buffer_14_757 = $signed(_T_80230); // @[Modules.scala 78:156:@35596.4]
  assign _T_80232 = $signed(buffer_14_757) + $signed(buffer_14_709); // @[Modules.scala 78:156:@35598.4]
  assign _T_80233 = _T_80232[10:0]; // @[Modules.scala 78:156:@35599.4]
  assign buffer_14_758 = $signed(_T_80233); // @[Modules.scala 78:156:@35600.4]
  assign _T_80235 = $signed(buffer_14_758) + $signed(buffer_14_710); // @[Modules.scala 78:156:@35602.4]
  assign _T_80236 = _T_80235[10:0]; // @[Modules.scala 78:156:@35603.4]
  assign buffer_14_759 = $signed(_T_80236); // @[Modules.scala 78:156:@35604.4]
  assign _T_80238 = $signed(buffer_14_759) + $signed(buffer_14_711); // @[Modules.scala 78:156:@35606.4]
  assign _T_80239 = _T_80238[10:0]; // @[Modules.scala 78:156:@35607.4]
  assign buffer_14_760 = $signed(_T_80239); // @[Modules.scala 78:156:@35608.4]
  assign _T_80241 = $signed(buffer_14_760) + $signed(buffer_14_712); // @[Modules.scala 78:156:@35610.4]
  assign _T_80242 = _T_80241[10:0]; // @[Modules.scala 78:156:@35611.4]
  assign buffer_14_761 = $signed(_T_80242); // @[Modules.scala 78:156:@35612.4]
  assign _T_80244 = $signed(buffer_14_761) + $signed(buffer_14_713); // @[Modules.scala 78:156:@35614.4]
  assign _T_80245 = _T_80244[10:0]; // @[Modules.scala 78:156:@35615.4]
  assign buffer_14_762 = $signed(_T_80245); // @[Modules.scala 78:156:@35616.4]
  assign _T_80247 = $signed(buffer_14_762) + $signed(buffer_14_714); // @[Modules.scala 78:156:@35618.4]
  assign _T_80248 = _T_80247[10:0]; // @[Modules.scala 78:156:@35619.4]
  assign buffer_14_763 = $signed(_T_80248); // @[Modules.scala 78:156:@35620.4]
  assign _T_80250 = $signed(buffer_14_763) + $signed(buffer_14_715); // @[Modules.scala 78:156:@35622.4]
  assign _T_80251 = _T_80250[10:0]; // @[Modules.scala 78:156:@35623.4]
  assign buffer_14_764 = $signed(_T_80251); // @[Modules.scala 78:156:@35624.4]
  assign _T_80253 = $signed(buffer_14_764) + $signed(buffer_14_716); // @[Modules.scala 78:156:@35626.4]
  assign _T_80254 = _T_80253[10:0]; // @[Modules.scala 78:156:@35627.4]
  assign buffer_14_765 = $signed(_T_80254); // @[Modules.scala 78:156:@35628.4]
  assign _T_80256 = $signed(buffer_14_765) + $signed(buffer_14_717); // @[Modules.scala 78:156:@35630.4]
  assign _T_80257 = _T_80256[10:0]; // @[Modules.scala 78:156:@35631.4]
  assign buffer_14_766 = $signed(_T_80257); // @[Modules.scala 78:156:@35632.4]
  assign _T_80259 = $signed(buffer_14_766) + $signed(buffer_14_718); // @[Modules.scala 78:156:@35634.4]
  assign _T_80260 = _T_80259[10:0]; // @[Modules.scala 78:156:@35635.4]
  assign buffer_14_767 = $signed(_T_80260); // @[Modules.scala 78:156:@35636.4]
  assign _T_80262 = $signed(buffer_14_767) + $signed(buffer_14_719); // @[Modules.scala 78:156:@35638.4]
  assign _T_80263 = _T_80262[10:0]; // @[Modules.scala 78:156:@35639.4]
  assign buffer_14_768 = $signed(_T_80263); // @[Modules.scala 78:156:@35640.4]
  assign _T_80265 = $signed(buffer_14_768) + $signed(buffer_14_720); // @[Modules.scala 78:156:@35642.4]
  assign _T_80266 = _T_80265[10:0]; // @[Modules.scala 78:156:@35643.4]
  assign buffer_14_769 = $signed(_T_80266); // @[Modules.scala 78:156:@35644.4]
  assign _T_80268 = $signed(buffer_14_769) + $signed(buffer_14_721); // @[Modules.scala 78:156:@35646.4]
  assign _T_80269 = _T_80268[10:0]; // @[Modules.scala 78:156:@35647.4]
  assign buffer_14_770 = $signed(_T_80269); // @[Modules.scala 78:156:@35648.4]
  assign _T_80271 = $signed(buffer_14_770) + $signed(buffer_14_722); // @[Modules.scala 78:156:@35650.4]
  assign _T_80272 = _T_80271[10:0]; // @[Modules.scala 78:156:@35651.4]
  assign buffer_14_771 = $signed(_T_80272); // @[Modules.scala 78:156:@35652.4]
  assign _T_80274 = $signed(buffer_14_771) + $signed(buffer_14_723); // @[Modules.scala 78:156:@35654.4]
  assign _T_80275 = _T_80274[10:0]; // @[Modules.scala 78:156:@35655.4]
  assign buffer_14_772 = $signed(_T_80275); // @[Modules.scala 78:156:@35656.4]
  assign _T_80277 = $signed(buffer_14_772) + $signed(buffer_14_724); // @[Modules.scala 78:156:@35658.4]
  assign _T_80278 = _T_80277[10:0]; // @[Modules.scala 78:156:@35659.4]
  assign buffer_14_773 = $signed(_T_80278); // @[Modules.scala 78:156:@35660.4]
  assign _T_80280 = $signed(buffer_14_773) + $signed(buffer_14_725); // @[Modules.scala 78:156:@35662.4]
  assign _T_80281 = _T_80280[10:0]; // @[Modules.scala 78:156:@35663.4]
  assign buffer_14_774 = $signed(_T_80281); // @[Modules.scala 78:156:@35664.4]
  assign _T_80283 = $signed(buffer_14_774) + $signed(buffer_14_726); // @[Modules.scala 78:156:@35666.4]
  assign _T_80284 = _T_80283[10:0]; // @[Modules.scala 78:156:@35667.4]
  assign buffer_14_775 = $signed(_T_80284); // @[Modules.scala 78:156:@35668.4]
  assign _T_80286 = $signed(buffer_14_775) + $signed(buffer_14_727); // @[Modules.scala 78:156:@35670.4]
  assign _T_80287 = _T_80286[10:0]; // @[Modules.scala 78:156:@35671.4]
  assign buffer_14_776 = $signed(_T_80287); // @[Modules.scala 78:156:@35672.4]
  assign _T_80289 = $signed(buffer_14_776) + $signed(buffer_14_728); // @[Modules.scala 78:156:@35674.4]
  assign _T_80290 = _T_80289[10:0]; // @[Modules.scala 78:156:@35675.4]
  assign buffer_14_777 = $signed(_T_80290); // @[Modules.scala 78:156:@35676.4]
  assign _T_80292 = $signed(buffer_14_777) + $signed(buffer_14_729); // @[Modules.scala 78:156:@35678.4]
  assign _T_80293 = _T_80292[10:0]; // @[Modules.scala 78:156:@35679.4]
  assign buffer_14_778 = $signed(_T_80293); // @[Modules.scala 78:156:@35680.4]
  assign _T_80295 = $signed(buffer_14_778) + $signed(buffer_14_730); // @[Modules.scala 78:156:@35682.4]
  assign _T_80296 = _T_80295[10:0]; // @[Modules.scala 78:156:@35683.4]
  assign buffer_14_779 = $signed(_T_80296); // @[Modules.scala 78:156:@35684.4]
  assign _T_80298 = $signed(buffer_14_779) + $signed(buffer_14_731); // @[Modules.scala 78:156:@35686.4]
  assign _T_80299 = _T_80298[10:0]; // @[Modules.scala 78:156:@35687.4]
  assign buffer_14_780 = $signed(_T_80299); // @[Modules.scala 78:156:@35688.4]
  assign _T_80301 = $signed(buffer_14_780) + $signed(buffer_14_732); // @[Modules.scala 78:156:@35690.4]
  assign _T_80302 = _T_80301[10:0]; // @[Modules.scala 78:156:@35691.4]
  assign buffer_14_781 = $signed(_T_80302); // @[Modules.scala 78:156:@35692.4]
  assign _T_80304 = $signed(buffer_14_781) + $signed(buffer_14_733); // @[Modules.scala 78:156:@35694.4]
  assign _T_80305 = _T_80304[10:0]; // @[Modules.scala 78:156:@35695.4]
  assign buffer_14_782 = $signed(_T_80305); // @[Modules.scala 78:156:@35696.4]
  assign _T_80307 = $signed(buffer_14_782) + $signed(buffer_14_734); // @[Modules.scala 78:156:@35698.4]
  assign _T_80308 = _T_80307[10:0]; // @[Modules.scala 78:156:@35699.4]
  assign buffer_14_783 = $signed(_T_80308); // @[Modules.scala 78:156:@35700.4]
  assign _T_80589 = $signed(io_in_366) + $signed(io_in_367); // @[Modules.scala 37:46:@36108.4]
  assign _T_80590 = _T_80589[4:0]; // @[Modules.scala 37:46:@36109.4]
  assign _T_80591 = $signed(_T_80590); // @[Modules.scala 37:46:@36110.4]
  assign _T_80926 = $signed(buffer_1_6) + $signed(11'sh0); // @[Modules.scala 65:57:@36599.4]
  assign _T_80927 = _T_80926[10:0]; // @[Modules.scala 65:57:@36600.4]
  assign buffer_15_395 = $signed(_T_80927); // @[Modules.scala 65:57:@36601.4]
  assign _T_80929 = $signed(buffer_0_8) + $signed(buffer_9_9); // @[Modules.scala 65:57:@36603.4]
  assign _T_80930 = _T_80929[10:0]; // @[Modules.scala 65:57:@36604.4]
  assign buffer_15_396 = $signed(_T_80930); // @[Modules.scala 65:57:@36605.4]
  assign _T_80932 = $signed(buffer_5_10) + $signed(buffer_1_11); // @[Modules.scala 65:57:@36607.4]
  assign _T_80933 = _T_80932[10:0]; // @[Modules.scala 65:57:@36608.4]
  assign buffer_15_397 = $signed(_T_80933); // @[Modules.scala 65:57:@36609.4]
  assign _T_80935 = $signed(buffer_0_12) + $signed(buffer_4_13); // @[Modules.scala 65:57:@36611.4]
  assign _T_80936 = _T_80935[10:0]; // @[Modules.scala 65:57:@36612.4]
  assign buffer_15_398 = $signed(_T_80936); // @[Modules.scala 65:57:@36613.4]
  assign _T_80944 = $signed(11'sh0) + $signed(buffer_1_19); // @[Modules.scala 65:57:@36623.4]
  assign _T_80945 = _T_80944[10:0]; // @[Modules.scala 65:57:@36624.4]
  assign buffer_15_401 = $signed(_T_80945); // @[Modules.scala 65:57:@36625.4]
  assign _T_80950 = $signed(buffer_4_22) + $signed(buffer_11_23); // @[Modules.scala 65:57:@36631.4]
  assign _T_80951 = _T_80950[10:0]; // @[Modules.scala 65:57:@36632.4]
  assign buffer_15_403 = $signed(_T_80951); // @[Modules.scala 65:57:@36633.4]
  assign buffer_15_24 = {{6{io_in_48[4]}},io_in_48}; // @[Modules.scala 32:22:@8.4]
  assign _T_80953 = $signed(buffer_15_24) + $signed(buffer_1_25); // @[Modules.scala 65:57:@36635.4]
  assign _T_80954 = _T_80953[10:0]; // @[Modules.scala 65:57:@36636.4]
  assign buffer_15_404 = $signed(_T_80954); // @[Modules.scala 65:57:@36637.4]
  assign buffer_15_38 = {{6{io_in_77[4]}},io_in_77}; // @[Modules.scala 32:22:@8.4]
  assign _T_80974 = $signed(buffer_15_38) + $signed(buffer_0_39); // @[Modules.scala 65:57:@36663.4]
  assign _T_80975 = _T_80974[10:0]; // @[Modules.scala 65:57:@36664.4]
  assign buffer_15_411 = $signed(_T_80975); // @[Modules.scala 65:57:@36665.4]
  assign _T_80980 = $signed(buffer_1_42) + $signed(buffer_11_43); // @[Modules.scala 65:57:@36671.4]
  assign _T_80981 = _T_80980[10:0]; // @[Modules.scala 65:57:@36672.4]
  assign buffer_15_413 = $signed(_T_80981); // @[Modules.scala 65:57:@36673.4]
  assign _T_80983 = $signed(11'sh0) + $signed(buffer_14_45); // @[Modules.scala 65:57:@36675.4]
  assign _T_80984 = _T_80983[10:0]; // @[Modules.scala 65:57:@36676.4]
  assign buffer_15_414 = $signed(_T_80984); // @[Modules.scala 65:57:@36677.4]
  assign _T_81007 = $signed(buffer_8_60) + $signed(11'sh0); // @[Modules.scala 65:57:@36707.4]
  assign _T_81008 = _T_81007[10:0]; // @[Modules.scala 65:57:@36708.4]
  assign buffer_15_422 = $signed(_T_81008); // @[Modules.scala 65:57:@36709.4]
  assign _T_81013 = $signed(buffer_1_64) + $signed(buffer_0_65); // @[Modules.scala 65:57:@36715.4]
  assign _T_81014 = _T_81013[10:0]; // @[Modules.scala 65:57:@36716.4]
  assign buffer_15_424 = $signed(_T_81014); // @[Modules.scala 65:57:@36717.4]
  assign _T_81022 = $signed(11'sh0) + $signed(buffer_1_71); // @[Modules.scala 65:57:@36727.4]
  assign _T_81023 = _T_81022[10:0]; // @[Modules.scala 65:57:@36728.4]
  assign buffer_15_427 = $signed(_T_81023); // @[Modules.scala 65:57:@36729.4]
  assign _T_81031 = $signed(buffer_3_76) + $signed(buffer_10_77); // @[Modules.scala 65:57:@36739.4]
  assign _T_81032 = _T_81031[10:0]; // @[Modules.scala 65:57:@36740.4]
  assign buffer_15_430 = $signed(_T_81032); // @[Modules.scala 65:57:@36741.4]
  assign _T_81034 = $signed(11'sh0) + $signed(buffer_3_79); // @[Modules.scala 65:57:@36743.4]
  assign _T_81035 = _T_81034[10:0]; // @[Modules.scala 65:57:@36744.4]
  assign buffer_15_431 = $signed(_T_81035); // @[Modules.scala 65:57:@36745.4]
  assign _T_81043 = $signed(11'sh0) + $signed(buffer_9_85); // @[Modules.scala 65:57:@36755.4]
  assign _T_81044 = _T_81043[10:0]; // @[Modules.scala 65:57:@36756.4]
  assign buffer_15_434 = $signed(_T_81044); // @[Modules.scala 65:57:@36757.4]
  assign _T_81046 = $signed(11'sh0) + $signed(buffer_1_87); // @[Modules.scala 65:57:@36759.4]
  assign _T_81047 = _T_81046[10:0]; // @[Modules.scala 65:57:@36760.4]
  assign buffer_15_435 = $signed(_T_81047); // @[Modules.scala 65:57:@36761.4]
  assign _T_81049 = $signed(buffer_10_88) + $signed(buffer_1_89); // @[Modules.scala 65:57:@36763.4]
  assign _T_81050 = _T_81049[10:0]; // @[Modules.scala 65:57:@36764.4]
  assign buffer_15_436 = $signed(_T_81050); // @[Modules.scala 65:57:@36765.4]
  assign _T_81064 = $signed(buffer_0_98) + $signed(buffer_3_99); // @[Modules.scala 65:57:@36783.4]
  assign _T_81065 = _T_81064[10:0]; // @[Modules.scala 65:57:@36784.4]
  assign buffer_15_441 = $signed(_T_81065); // @[Modules.scala 65:57:@36785.4]
  assign _T_81067 = $signed(11'sh0) + $signed(buffer_1_101); // @[Modules.scala 65:57:@36787.4]
  assign _T_81068 = _T_81067[10:0]; // @[Modules.scala 65:57:@36788.4]
  assign buffer_15_442 = $signed(_T_81068); // @[Modules.scala 65:57:@36789.4]
  assign _T_81076 = $signed(11'sh0) + $signed(buffer_2_107); // @[Modules.scala 65:57:@36799.4]
  assign _T_81077 = _T_81076[10:0]; // @[Modules.scala 65:57:@36800.4]
  assign buffer_15_445 = $signed(_T_81077); // @[Modules.scala 65:57:@36801.4]
  assign _T_81091 = $signed(11'sh0) + $signed(buffer_3_117); // @[Modules.scala 65:57:@36819.4]
  assign _T_81092 = _T_81091[10:0]; // @[Modules.scala 65:57:@36820.4]
  assign buffer_15_450 = $signed(_T_81092); // @[Modules.scala 65:57:@36821.4]
  assign buffer_15_129 = {{6{io_in_259[4]}},io_in_259}; // @[Modules.scala 32:22:@8.4]
  assign _T_81109 = $signed(buffer_3_128) + $signed(buffer_15_129); // @[Modules.scala 65:57:@36843.4]
  assign _T_81110 = _T_81109[10:0]; // @[Modules.scala 65:57:@36844.4]
  assign buffer_15_456 = $signed(_T_81110); // @[Modules.scala 65:57:@36845.4]
  assign _T_81130 = $signed(buffer_7_142) + $signed(buffer_2_143); // @[Modules.scala 65:57:@36871.4]
  assign _T_81131 = _T_81130[10:0]; // @[Modules.scala 65:57:@36872.4]
  assign buffer_15_463 = $signed(_T_81131); // @[Modules.scala 65:57:@36873.4]
  assign _T_81142 = $signed(buffer_5_150) + $signed(11'sh0); // @[Modules.scala 65:57:@36887.4]
  assign _T_81143 = _T_81142[10:0]; // @[Modules.scala 65:57:@36888.4]
  assign buffer_15_467 = $signed(_T_81143); // @[Modules.scala 65:57:@36889.4]
  assign _T_81151 = $signed(buffer_9_156) + $signed(buffer_2_157); // @[Modules.scala 65:57:@36899.4]
  assign _T_81152 = _T_81151[10:0]; // @[Modules.scala 65:57:@36900.4]
  assign buffer_15_470 = $signed(_T_81152); // @[Modules.scala 65:57:@36901.4]
  assign _T_81154 = $signed(buffer_13_158) + $signed(11'sh0); // @[Modules.scala 65:57:@36903.4]
  assign _T_81155 = _T_81154[10:0]; // @[Modules.scala 65:57:@36904.4]
  assign buffer_15_471 = $signed(_T_81155); // @[Modules.scala 65:57:@36905.4]
  assign _T_81160 = $signed(buffer_0_162) + $signed(buffer_5_163); // @[Modules.scala 65:57:@36911.4]
  assign _T_81161 = _T_81160[10:0]; // @[Modules.scala 65:57:@36912.4]
  assign buffer_15_473 = $signed(_T_81161); // @[Modules.scala 65:57:@36913.4]
  assign _T_81169 = $signed(buffer_5_168) + $signed(buffer_6_169); // @[Modules.scala 65:57:@36923.4]
  assign _T_81170 = _T_81169[10:0]; // @[Modules.scala 65:57:@36924.4]
  assign buffer_15_476 = $signed(_T_81170); // @[Modules.scala 65:57:@36925.4]
  assign _T_81187 = $signed(buffer_14_180) + $signed(buffer_0_181); // @[Modules.scala 65:57:@36947.4]
  assign _T_81188 = _T_81187[10:0]; // @[Modules.scala 65:57:@36948.4]
  assign buffer_15_482 = $signed(_T_81188); // @[Modules.scala 65:57:@36949.4]
  assign buffer_15_183 = {{6{_T_80591[4]}},_T_80591}; // @[Modules.scala 32:22:@8.4]
  assign _T_81190 = $signed(buffer_3_182) + $signed(buffer_15_183); // @[Modules.scala 65:57:@36951.4]
  assign _T_81191 = _T_81190[10:0]; // @[Modules.scala 65:57:@36952.4]
  assign buffer_15_483 = $signed(_T_81191); // @[Modules.scala 65:57:@36953.4]
  assign _T_81193 = $signed(buffer_0_184) + $signed(11'sh0); // @[Modules.scala 65:57:@36955.4]
  assign _T_81194 = _T_81193[10:0]; // @[Modules.scala 65:57:@36956.4]
  assign buffer_15_484 = $signed(_T_81194); // @[Modules.scala 65:57:@36957.4]
  assign _T_81223 = $signed(11'sh0) + $signed(buffer_2_205); // @[Modules.scala 65:57:@36995.4]
  assign _T_81224 = _T_81223[10:0]; // @[Modules.scala 65:57:@36996.4]
  assign buffer_15_494 = $signed(_T_81224); // @[Modules.scala 65:57:@36997.4]
  assign _T_81244 = $signed(11'sh0) + $signed(buffer_6_219); // @[Modules.scala 65:57:@37023.4]
  assign _T_81245 = _T_81244[10:0]; // @[Modules.scala 65:57:@37024.4]
  assign buffer_15_501 = $signed(_T_81245); // @[Modules.scala 65:57:@37025.4]
  assign _T_81259 = $signed(buffer_0_228) + $signed(buffer_1_229); // @[Modules.scala 65:57:@37043.4]
  assign _T_81260 = _T_81259[10:0]; // @[Modules.scala 65:57:@37044.4]
  assign buffer_15_506 = $signed(_T_81260); // @[Modules.scala 65:57:@37045.4]
  assign _T_81262 = $signed(11'sh0) + $signed(buffer_4_231); // @[Modules.scala 65:57:@37047.4]
  assign _T_81263 = _T_81262[10:0]; // @[Modules.scala 65:57:@37048.4]
  assign buffer_15_507 = $signed(_T_81263); // @[Modules.scala 65:57:@37049.4]
  assign _T_81286 = $signed(buffer_0_246) + $signed(buffer_1_247); // @[Modules.scala 65:57:@37079.4]
  assign _T_81287 = _T_81286[10:0]; // @[Modules.scala 65:57:@37080.4]
  assign buffer_15_515 = $signed(_T_81287); // @[Modules.scala 65:57:@37081.4]
  assign buffer_15_249 = {{6{io_in_498[4]}},io_in_498}; // @[Modules.scala 32:22:@8.4]
  assign _T_81289 = $signed(buffer_13_248) + $signed(buffer_15_249); // @[Modules.scala 65:57:@37083.4]
  assign _T_81290 = _T_81289[10:0]; // @[Modules.scala 65:57:@37084.4]
  assign buffer_15_516 = $signed(_T_81290); // @[Modules.scala 65:57:@37085.4]
  assign _T_81310 = $signed(11'sh0) + $signed(buffer_7_263); // @[Modules.scala 65:57:@37111.4]
  assign _T_81311 = _T_81310[10:0]; // @[Modules.scala 65:57:@37112.4]
  assign buffer_15_523 = $signed(_T_81311); // @[Modules.scala 65:57:@37113.4]
  assign _T_81325 = $signed(buffer_1_272) + $signed(buffer_3_273); // @[Modules.scala 65:57:@37131.4]
  assign _T_81326 = _T_81325[10:0]; // @[Modules.scala 65:57:@37132.4]
  assign buffer_15_528 = $signed(_T_81326); // @[Modules.scala 65:57:@37133.4]
  assign _T_81328 = $signed(buffer_2_274) + $signed(buffer_0_275); // @[Modules.scala 65:57:@37135.4]
  assign _T_81329 = _T_81328[10:0]; // @[Modules.scala 65:57:@37136.4]
  assign buffer_15_529 = $signed(_T_81329); // @[Modules.scala 65:57:@37137.4]
  assign _T_81343 = $signed(11'sh0) + $signed(buffer_1_285); // @[Modules.scala 65:57:@37155.4]
  assign _T_81344 = _T_81343[10:0]; // @[Modules.scala 65:57:@37156.4]
  assign buffer_15_534 = $signed(_T_81344); // @[Modules.scala 65:57:@37157.4]
  assign buffer_15_287 = {{6{io_in_574[4]}},io_in_574}; // @[Modules.scala 32:22:@8.4]
  assign _T_81346 = $signed(buffer_1_286) + $signed(buffer_15_287); // @[Modules.scala 65:57:@37159.4]
  assign _T_81347 = _T_81346[10:0]; // @[Modules.scala 65:57:@37160.4]
  assign buffer_15_535 = $signed(_T_81347); // @[Modules.scala 65:57:@37161.4]
  assign _T_81349 = $signed(buffer_0_288) + $signed(buffer_5_289); // @[Modules.scala 65:57:@37163.4]
  assign _T_81350 = _T_81349[10:0]; // @[Modules.scala 65:57:@37164.4]
  assign buffer_15_536 = $signed(_T_81350); // @[Modules.scala 65:57:@37165.4]
  assign _T_81358 = $signed(buffer_2_294) + $signed(11'sh0); // @[Modules.scala 65:57:@37175.4]
  assign _T_81359 = _T_81358[10:0]; // @[Modules.scala 65:57:@37176.4]
  assign buffer_15_539 = $signed(_T_81359); // @[Modules.scala 65:57:@37177.4]
  assign _T_81364 = $signed(11'sh0) + $signed(buffer_7_299); // @[Modules.scala 65:57:@37183.4]
  assign _T_81365 = _T_81364[10:0]; // @[Modules.scala 65:57:@37184.4]
  assign buffer_15_541 = $signed(_T_81365); // @[Modules.scala 65:57:@37185.4]
  assign _T_81367 = $signed(buffer_2_300) + $signed(buffer_0_301); // @[Modules.scala 65:57:@37187.4]
  assign _T_81368 = _T_81367[10:0]; // @[Modules.scala 65:57:@37188.4]
  assign buffer_15_542 = $signed(_T_81368); // @[Modules.scala 65:57:@37189.4]
  assign _T_81370 = $signed(buffer_5_302) + $signed(buffer_8_303); // @[Modules.scala 65:57:@37191.4]
  assign _T_81371 = _T_81370[10:0]; // @[Modules.scala 65:57:@37192.4]
  assign buffer_15_543 = $signed(_T_81371); // @[Modules.scala 65:57:@37193.4]
  assign _T_81373 = $signed(11'sh0) + $signed(buffer_3_305); // @[Modules.scala 65:57:@37195.4]
  assign _T_81374 = _T_81373[10:0]; // @[Modules.scala 65:57:@37196.4]
  assign buffer_15_544 = $signed(_T_81374); // @[Modules.scala 65:57:@37197.4]
  assign buffer_15_308 = {{6{io_in_616[4]}},io_in_616}; // @[Modules.scala 32:22:@8.4]
  assign _T_81379 = $signed(buffer_15_308) + $signed(11'sh0); // @[Modules.scala 65:57:@37203.4]
  assign _T_81380 = _T_81379[10:0]; // @[Modules.scala 65:57:@37204.4]
  assign buffer_15_546 = $signed(_T_81380); // @[Modules.scala 65:57:@37205.4]
  assign _T_81382 = $signed(buffer_11_310) + $signed(11'sh0); // @[Modules.scala 65:57:@37207.4]
  assign _T_81383 = _T_81382[10:0]; // @[Modules.scala 65:57:@37208.4]
  assign buffer_15_547 = $signed(_T_81383); // @[Modules.scala 65:57:@37209.4]
  assign _T_81388 = $signed(11'sh0) + $signed(buffer_1_315); // @[Modules.scala 65:57:@37215.4]
  assign _T_81389 = _T_81388[10:0]; // @[Modules.scala 65:57:@37216.4]
  assign buffer_15_549 = $signed(_T_81389); // @[Modules.scala 65:57:@37217.4]
  assign _T_81397 = $signed(buffer_0_320) + $signed(buffer_1_321); // @[Modules.scala 65:57:@37227.4]
  assign _T_81398 = _T_81397[10:0]; // @[Modules.scala 65:57:@37228.4]
  assign buffer_15_552 = $signed(_T_81398); // @[Modules.scala 65:57:@37229.4]
  assign _T_81400 = $signed(buffer_0_322) + $signed(11'sh0); // @[Modules.scala 65:57:@37231.4]
  assign _T_81401 = _T_81400[10:0]; // @[Modules.scala 65:57:@37232.4]
  assign buffer_15_553 = $signed(_T_81401); // @[Modules.scala 65:57:@37233.4]
  assign _T_81403 = $signed(11'sh0) + $signed(buffer_3_325); // @[Modules.scala 65:57:@37235.4]
  assign _T_81404 = _T_81403[10:0]; // @[Modules.scala 65:57:@37236.4]
  assign buffer_15_554 = $signed(_T_81404); // @[Modules.scala 65:57:@37237.4]
  assign buffer_15_338 = {{6{io_in_677[4]}},io_in_677}; // @[Modules.scala 32:22:@8.4]
  assign _T_81424 = $signed(buffer_15_338) + $signed(11'sh0); // @[Modules.scala 65:57:@37263.4]
  assign _T_81425 = _T_81424[10:0]; // @[Modules.scala 65:57:@37264.4]
  assign buffer_15_561 = $signed(_T_81425); // @[Modules.scala 65:57:@37265.4]
  assign _T_81427 = $signed(11'sh0) + $signed(buffer_1_341); // @[Modules.scala 65:57:@37267.4]
  assign _T_81428 = _T_81427[10:0]; // @[Modules.scala 65:57:@37268.4]
  assign buffer_15_562 = $signed(_T_81428); // @[Modules.scala 65:57:@37269.4]
  assign _T_81442 = $signed(buffer_1_350) + $signed(11'sh0); // @[Modules.scala 65:57:@37287.4]
  assign _T_81443 = _T_81442[10:0]; // @[Modules.scala 65:57:@37288.4]
  assign buffer_15_567 = $signed(_T_81443); // @[Modules.scala 65:57:@37289.4]
  assign _T_81445 = $signed(buffer_0_352) + $signed(11'sh0); // @[Modules.scala 65:57:@37291.4]
  assign _T_81446 = _T_81445[10:0]; // @[Modules.scala 65:57:@37292.4]
  assign buffer_15_568 = $signed(_T_81446); // @[Modules.scala 65:57:@37293.4]
  assign buffer_15_356 = {{6{io_in_713[4]}},io_in_713}; // @[Modules.scala 32:22:@8.4]
  assign _T_81451 = $signed(buffer_15_356) + $signed(11'sh0); // @[Modules.scala 65:57:@37299.4]
  assign _T_81452 = _T_81451[10:0]; // @[Modules.scala 65:57:@37300.4]
  assign buffer_15_570 = $signed(_T_81452); // @[Modules.scala 65:57:@37301.4]
  assign buffer_15_366 = {{6{io_in_733[4]}},io_in_733}; // @[Modules.scala 32:22:@8.4]
  assign _T_81466 = $signed(buffer_15_366) + $signed(buffer_0_367); // @[Modules.scala 65:57:@37319.4]
  assign _T_81467 = _T_81466[10:0]; // @[Modules.scala 65:57:@37320.4]
  assign buffer_15_575 = $signed(_T_81467); // @[Modules.scala 65:57:@37321.4]
  assign buffer_15_389 = {{6{io_in_778[4]}},io_in_778}; // @[Modules.scala 32:22:@8.4]
  assign _T_81499 = $signed(buffer_0_388) + $signed(buffer_15_389); // @[Modules.scala 65:57:@37363.4]
  assign _T_81500 = _T_81499[10:0]; // @[Modules.scala 65:57:@37364.4]
  assign buffer_15_586 = $signed(_T_81500); // @[Modules.scala 65:57:@37365.4]
  assign _T_81505 = $signed(buffer_14_392) + $signed(buffer_0_393); // @[Modules.scala 68:83:@37371.4]
  assign _T_81506 = _T_81505[10:0]; // @[Modules.scala 68:83:@37372.4]
  assign buffer_15_588 = $signed(_T_81506); // @[Modules.scala 68:83:@37373.4]
  assign _T_81508 = $signed(buffer_8_394) + $signed(buffer_15_395); // @[Modules.scala 68:83:@37375.4]
  assign _T_81509 = _T_81508[10:0]; // @[Modules.scala 68:83:@37376.4]
  assign buffer_15_589 = $signed(_T_81509); // @[Modules.scala 68:83:@37377.4]
  assign _T_81511 = $signed(buffer_15_396) + $signed(buffer_15_397); // @[Modules.scala 68:83:@37379.4]
  assign _T_81512 = _T_81511[10:0]; // @[Modules.scala 68:83:@37380.4]
  assign buffer_15_590 = $signed(_T_81512); // @[Modules.scala 68:83:@37381.4]
  assign _T_81514 = $signed(buffer_15_398) + $signed(buffer_12_399); // @[Modules.scala 68:83:@37383.4]
  assign _T_81515 = _T_81514[10:0]; // @[Modules.scala 68:83:@37384.4]
  assign buffer_15_591 = $signed(_T_81515); // @[Modules.scala 68:83:@37385.4]
  assign _T_81517 = $signed(buffer_2_400) + $signed(buffer_15_401); // @[Modules.scala 68:83:@37387.4]
  assign _T_81518 = _T_81517[10:0]; // @[Modules.scala 68:83:@37388.4]
  assign buffer_15_592 = $signed(_T_81518); // @[Modules.scala 68:83:@37389.4]
  assign _T_81520 = $signed(buffer_1_402) + $signed(buffer_15_403); // @[Modules.scala 68:83:@37391.4]
  assign _T_81521 = _T_81520[10:0]; // @[Modules.scala 68:83:@37392.4]
  assign buffer_15_593 = $signed(_T_81521); // @[Modules.scala 68:83:@37393.4]
  assign _T_81523 = $signed(buffer_15_404) + $signed(buffer_0_395); // @[Modules.scala 68:83:@37395.4]
  assign _T_81524 = _T_81523[10:0]; // @[Modules.scala 68:83:@37396.4]
  assign buffer_15_594 = $signed(_T_81524); // @[Modules.scala 68:83:@37397.4]
  assign _T_81526 = $signed(buffer_5_406) + $signed(buffer_1_407); // @[Modules.scala 68:83:@37399.4]
  assign _T_81527 = _T_81526[10:0]; // @[Modules.scala 68:83:@37400.4]
  assign buffer_15_595 = $signed(_T_81527); // @[Modules.scala 68:83:@37401.4]
  assign _T_81532 = $signed(buffer_1_410) + $signed(buffer_15_411); // @[Modules.scala 68:83:@37407.4]
  assign _T_81533 = _T_81532[10:0]; // @[Modules.scala 68:83:@37408.4]
  assign buffer_15_597 = $signed(_T_81533); // @[Modules.scala 68:83:@37409.4]
  assign _T_81535 = $signed(buffer_3_412) + $signed(buffer_15_413); // @[Modules.scala 68:83:@37411.4]
  assign _T_81536 = _T_81535[10:0]; // @[Modules.scala 68:83:@37412.4]
  assign buffer_15_598 = $signed(_T_81536); // @[Modules.scala 68:83:@37413.4]
  assign _T_81538 = $signed(buffer_15_414) + $signed(buffer_1_415); // @[Modules.scala 68:83:@37415.4]
  assign _T_81539 = _T_81538[10:0]; // @[Modules.scala 68:83:@37416.4]
  assign buffer_15_599 = $signed(_T_81539); // @[Modules.scala 68:83:@37417.4]
  assign _T_81547 = $signed(buffer_0_420) + $signed(buffer_12_421); // @[Modules.scala 68:83:@37427.4]
  assign _T_81548 = _T_81547[10:0]; // @[Modules.scala 68:83:@37428.4]
  assign buffer_15_602 = $signed(_T_81548); // @[Modules.scala 68:83:@37429.4]
  assign _T_81550 = $signed(buffer_15_422) + $signed(buffer_14_423); // @[Modules.scala 68:83:@37431.4]
  assign _T_81551 = _T_81550[10:0]; // @[Modules.scala 68:83:@37432.4]
  assign buffer_15_603 = $signed(_T_81551); // @[Modules.scala 68:83:@37433.4]
  assign _T_81553 = $signed(buffer_15_424) + $signed(buffer_0_425); // @[Modules.scala 68:83:@37435.4]
  assign _T_81554 = _T_81553[10:0]; // @[Modules.scala 68:83:@37436.4]
  assign buffer_15_604 = $signed(_T_81554); // @[Modules.scala 68:83:@37437.4]
  assign _T_81556 = $signed(buffer_12_426) + $signed(buffer_15_427); // @[Modules.scala 68:83:@37439.4]
  assign _T_81557 = _T_81556[10:0]; // @[Modules.scala 68:83:@37440.4]
  assign buffer_15_605 = $signed(_T_81557); // @[Modules.scala 68:83:@37441.4]
  assign _T_81559 = $signed(buffer_0_395) + $signed(buffer_0_429); // @[Modules.scala 68:83:@37443.4]
  assign _T_81560 = _T_81559[10:0]; // @[Modules.scala 68:83:@37444.4]
  assign buffer_15_606 = $signed(_T_81560); // @[Modules.scala 68:83:@37445.4]
  assign _T_81562 = $signed(buffer_15_430) + $signed(buffer_15_431); // @[Modules.scala 68:83:@37447.4]
  assign _T_81563 = _T_81562[10:0]; // @[Modules.scala 68:83:@37448.4]
  assign buffer_15_607 = $signed(_T_81563); // @[Modules.scala 68:83:@37449.4]
  assign _T_81565 = $signed(buffer_5_432) + $signed(buffer_0_395); // @[Modules.scala 68:83:@37451.4]
  assign _T_81566 = _T_81565[10:0]; // @[Modules.scala 68:83:@37452.4]
  assign buffer_15_608 = $signed(_T_81566); // @[Modules.scala 68:83:@37453.4]
  assign _T_81568 = $signed(buffer_15_434) + $signed(buffer_15_435); // @[Modules.scala 68:83:@37455.4]
  assign _T_81569 = _T_81568[10:0]; // @[Modules.scala 68:83:@37456.4]
  assign buffer_15_609 = $signed(_T_81569); // @[Modules.scala 68:83:@37457.4]
  assign _T_81571 = $signed(buffer_15_436) + $signed(buffer_1_437); // @[Modules.scala 68:83:@37459.4]
  assign _T_81572 = _T_81571[10:0]; // @[Modules.scala 68:83:@37460.4]
  assign buffer_15_610 = $signed(_T_81572); // @[Modules.scala 68:83:@37461.4]
  assign _T_81574 = $signed(buffer_4_438) + $signed(buffer_6_439); // @[Modules.scala 68:83:@37463.4]
  assign _T_81575 = _T_81574[10:0]; // @[Modules.scala 68:83:@37464.4]
  assign buffer_15_611 = $signed(_T_81575); // @[Modules.scala 68:83:@37465.4]
  assign _T_81577 = $signed(buffer_0_395) + $signed(buffer_15_441); // @[Modules.scala 68:83:@37467.4]
  assign _T_81578 = _T_81577[10:0]; // @[Modules.scala 68:83:@37468.4]
  assign buffer_15_612 = $signed(_T_81578); // @[Modules.scala 68:83:@37469.4]
  assign _T_81580 = $signed(buffer_15_442) + $signed(buffer_1_443); // @[Modules.scala 68:83:@37471.4]
  assign _T_81581 = _T_81580[10:0]; // @[Modules.scala 68:83:@37472.4]
  assign buffer_15_613 = $signed(_T_81581); // @[Modules.scala 68:83:@37473.4]
  assign _T_81583 = $signed(buffer_6_444) + $signed(buffer_15_445); // @[Modules.scala 68:83:@37475.4]
  assign _T_81584 = _T_81583[10:0]; // @[Modules.scala 68:83:@37476.4]
  assign buffer_15_614 = $signed(_T_81584); // @[Modules.scala 68:83:@37477.4]
  assign _T_81586 = $signed(buffer_9_446) + $signed(buffer_0_395); // @[Modules.scala 68:83:@37479.4]
  assign _T_81587 = _T_81586[10:0]; // @[Modules.scala 68:83:@37480.4]
  assign buffer_15_615 = $signed(_T_81587); // @[Modules.scala 68:83:@37481.4]
  assign _T_81589 = $signed(buffer_3_448) + $signed(buffer_13_449); // @[Modules.scala 68:83:@37483.4]
  assign _T_81590 = _T_81589[10:0]; // @[Modules.scala 68:83:@37484.4]
  assign buffer_15_616 = $signed(_T_81590); // @[Modules.scala 68:83:@37485.4]
  assign _T_81592 = $signed(buffer_15_450) + $signed(buffer_12_451); // @[Modules.scala 68:83:@37487.4]
  assign _T_81593 = _T_81592[10:0]; // @[Modules.scala 68:83:@37488.4]
  assign buffer_15_617 = $signed(_T_81593); // @[Modules.scala 68:83:@37489.4]
  assign _T_81595 = $signed(buffer_6_452) + $signed(buffer_9_453); // @[Modules.scala 68:83:@37491.4]
  assign _T_81596 = _T_81595[10:0]; // @[Modules.scala 68:83:@37492.4]
  assign buffer_15_618 = $signed(_T_81596); // @[Modules.scala 68:83:@37493.4]
  assign _T_81601 = $signed(buffer_15_456) + $signed(buffer_12_457); // @[Modules.scala 68:83:@37499.4]
  assign _T_81602 = _T_81601[10:0]; // @[Modules.scala 68:83:@37500.4]
  assign buffer_15_620 = $signed(_T_81602); // @[Modules.scala 68:83:@37501.4]
  assign _T_81604 = $signed(buffer_5_458) + $signed(buffer_3_459); // @[Modules.scala 68:83:@37503.4]
  assign _T_81605 = _T_81604[10:0]; // @[Modules.scala 68:83:@37504.4]
  assign buffer_15_621 = $signed(_T_81605); // @[Modules.scala 68:83:@37505.4]
  assign _T_81610 = $signed(buffer_3_462) + $signed(buffer_15_463); // @[Modules.scala 68:83:@37511.4]
  assign _T_81611 = _T_81610[10:0]; // @[Modules.scala 68:83:@37512.4]
  assign buffer_15_623 = $signed(_T_81611); // @[Modules.scala 68:83:@37513.4]
  assign _T_81616 = $signed(buffer_3_466) + $signed(buffer_15_467); // @[Modules.scala 68:83:@37519.4]
  assign _T_81617 = _T_81616[10:0]; // @[Modules.scala 68:83:@37520.4]
  assign buffer_15_625 = $signed(_T_81617); // @[Modules.scala 68:83:@37521.4]
  assign _T_81619 = $signed(buffer_0_395) + $signed(buffer_10_469); // @[Modules.scala 68:83:@37523.4]
  assign _T_81620 = _T_81619[10:0]; // @[Modules.scala 68:83:@37524.4]
  assign buffer_15_626 = $signed(_T_81620); // @[Modules.scala 68:83:@37525.4]
  assign _T_81622 = $signed(buffer_15_470) + $signed(buffer_15_471); // @[Modules.scala 68:83:@37527.4]
  assign _T_81623 = _T_81622[10:0]; // @[Modules.scala 68:83:@37528.4]
  assign buffer_15_627 = $signed(_T_81623); // @[Modules.scala 68:83:@37529.4]
  assign _T_81625 = $signed(buffer_0_395) + $signed(buffer_15_473); // @[Modules.scala 68:83:@37531.4]
  assign _T_81626 = _T_81625[10:0]; // @[Modules.scala 68:83:@37532.4]
  assign buffer_15_628 = $signed(_T_81626); // @[Modules.scala 68:83:@37533.4]
  assign _T_81628 = $signed(buffer_5_474) + $signed(buffer_0_395); // @[Modules.scala 68:83:@37535.4]
  assign _T_81629 = _T_81628[10:0]; // @[Modules.scala 68:83:@37536.4]
  assign buffer_15_629 = $signed(_T_81629); // @[Modules.scala 68:83:@37537.4]
  assign _T_81631 = $signed(buffer_15_476) + $signed(buffer_6_477); // @[Modules.scala 68:83:@37539.4]
  assign _T_81632 = _T_81631[10:0]; // @[Modules.scala 68:83:@37540.4]
  assign buffer_15_630 = $signed(_T_81632); // @[Modules.scala 68:83:@37541.4]
  assign _T_81637 = $signed(buffer_9_480) + $signed(buffer_0_481); // @[Modules.scala 68:83:@37547.4]
  assign _T_81638 = _T_81637[10:0]; // @[Modules.scala 68:83:@37548.4]
  assign buffer_15_632 = $signed(_T_81638); // @[Modules.scala 68:83:@37549.4]
  assign _T_81640 = $signed(buffer_15_482) + $signed(buffer_15_483); // @[Modules.scala 68:83:@37551.4]
  assign _T_81641 = _T_81640[10:0]; // @[Modules.scala 68:83:@37552.4]
  assign buffer_15_633 = $signed(_T_81641); // @[Modules.scala 68:83:@37553.4]
  assign _T_81643 = $signed(buffer_15_484) + $signed(buffer_0_395); // @[Modules.scala 68:83:@37555.4]
  assign _T_81644 = _T_81643[10:0]; // @[Modules.scala 68:83:@37556.4]
  assign buffer_15_634 = $signed(_T_81644); // @[Modules.scala 68:83:@37557.4]
  assign _T_81649 = $signed(buffer_4_488) + $signed(buffer_9_489); // @[Modules.scala 68:83:@37563.4]
  assign _T_81650 = _T_81649[10:0]; // @[Modules.scala 68:83:@37564.4]
  assign buffer_15_636 = $signed(_T_81650); // @[Modules.scala 68:83:@37565.4]
  assign _T_81658 = $signed(buffer_15_494) + $signed(buffer_0_495); // @[Modules.scala 68:83:@37575.4]
  assign _T_81659 = _T_81658[10:0]; // @[Modules.scala 68:83:@37576.4]
  assign buffer_15_639 = $signed(_T_81659); // @[Modules.scala 68:83:@37577.4]
  assign _T_81661 = $signed(buffer_10_496) + $signed(buffer_7_497); // @[Modules.scala 68:83:@37579.4]
  assign _T_81662 = _T_81661[10:0]; // @[Modules.scala 68:83:@37580.4]
  assign buffer_15_640 = $signed(_T_81662); // @[Modules.scala 68:83:@37581.4]
  assign _T_81667 = $signed(buffer_0_395) + $signed(buffer_15_501); // @[Modules.scala 68:83:@37587.4]
  assign _T_81668 = _T_81667[10:0]; // @[Modules.scala 68:83:@37588.4]
  assign buffer_15_642 = $signed(_T_81668); // @[Modules.scala 68:83:@37589.4]
  assign _T_81670 = $signed(buffer_1_502) + $signed(buffer_3_503); // @[Modules.scala 68:83:@37591.4]
  assign _T_81671 = _T_81670[10:0]; // @[Modules.scala 68:83:@37592.4]
  assign buffer_15_643 = $signed(_T_81671); // @[Modules.scala 68:83:@37593.4]
  assign _T_81676 = $signed(buffer_15_506) + $signed(buffer_15_507); // @[Modules.scala 68:83:@37599.4]
  assign _T_81677 = _T_81676[10:0]; // @[Modules.scala 68:83:@37600.4]
  assign buffer_15_645 = $signed(_T_81677); // @[Modules.scala 68:83:@37601.4]
  assign _T_81679 = $signed(buffer_0_508) + $signed(buffer_10_509); // @[Modules.scala 68:83:@37603.4]
  assign _T_81680 = _T_81679[10:0]; // @[Modules.scala 68:83:@37604.4]
  assign buffer_15_646 = $signed(_T_81680); // @[Modules.scala 68:83:@37605.4]
  assign _T_81688 = $signed(buffer_2_514) + $signed(buffer_15_515); // @[Modules.scala 68:83:@37615.4]
  assign _T_81689 = _T_81688[10:0]; // @[Modules.scala 68:83:@37616.4]
  assign buffer_15_649 = $signed(_T_81689); // @[Modules.scala 68:83:@37617.4]
  assign _T_81691 = $signed(buffer_15_516) + $signed(buffer_3_517); // @[Modules.scala 68:83:@37619.4]
  assign _T_81692 = _T_81691[10:0]; // @[Modules.scala 68:83:@37620.4]
  assign buffer_15_650 = $signed(_T_81692); // @[Modules.scala 68:83:@37621.4]
  assign _T_81694 = $signed(buffer_12_518) + $signed(buffer_8_519); // @[Modules.scala 68:83:@37623.4]
  assign _T_81695 = _T_81694[10:0]; // @[Modules.scala 68:83:@37624.4]
  assign buffer_15_651 = $signed(_T_81695); // @[Modules.scala 68:83:@37625.4]
  assign _T_81697 = $signed(buffer_0_520) + $signed(buffer_2_521); // @[Modules.scala 68:83:@37627.4]
  assign _T_81698 = _T_81697[10:0]; // @[Modules.scala 68:83:@37628.4]
  assign buffer_15_652 = $signed(_T_81698); // @[Modules.scala 68:83:@37629.4]
  assign _T_81700 = $signed(buffer_5_522) + $signed(buffer_15_523); // @[Modules.scala 68:83:@37631.4]
  assign _T_81701 = _T_81700[10:0]; // @[Modules.scala 68:83:@37632.4]
  assign buffer_15_653 = $signed(_T_81701); // @[Modules.scala 68:83:@37633.4]
  assign _T_81706 = $signed(buffer_0_395) + $signed(buffer_1_527); // @[Modules.scala 68:83:@37639.4]
  assign _T_81707 = _T_81706[10:0]; // @[Modules.scala 68:83:@37640.4]
  assign buffer_15_655 = $signed(_T_81707); // @[Modules.scala 68:83:@37641.4]
  assign _T_81709 = $signed(buffer_15_528) + $signed(buffer_15_529); // @[Modules.scala 68:83:@37643.4]
  assign _T_81710 = _T_81709[10:0]; // @[Modules.scala 68:83:@37644.4]
  assign buffer_15_656 = $signed(_T_81710); // @[Modules.scala 68:83:@37645.4]
  assign _T_81718 = $signed(buffer_15_534) + $signed(buffer_15_535); // @[Modules.scala 68:83:@37655.4]
  assign _T_81719 = _T_81718[10:0]; // @[Modules.scala 68:83:@37656.4]
  assign buffer_15_659 = $signed(_T_81719); // @[Modules.scala 68:83:@37657.4]
  assign _T_81721 = $signed(buffer_15_536) + $signed(buffer_10_537); // @[Modules.scala 68:83:@37659.4]
  assign _T_81722 = _T_81721[10:0]; // @[Modules.scala 68:83:@37660.4]
  assign buffer_15_660 = $signed(_T_81722); // @[Modules.scala 68:83:@37661.4]
  assign _T_81724 = $signed(buffer_8_538) + $signed(buffer_15_539); // @[Modules.scala 68:83:@37663.4]
  assign _T_81725 = _T_81724[10:0]; // @[Modules.scala 68:83:@37664.4]
  assign buffer_15_661 = $signed(_T_81725); // @[Modules.scala 68:83:@37665.4]
  assign _T_81727 = $signed(buffer_11_540) + $signed(buffer_15_541); // @[Modules.scala 68:83:@37667.4]
  assign _T_81728 = _T_81727[10:0]; // @[Modules.scala 68:83:@37668.4]
  assign buffer_15_662 = $signed(_T_81728); // @[Modules.scala 68:83:@37669.4]
  assign _T_81730 = $signed(buffer_15_542) + $signed(buffer_15_543); // @[Modules.scala 68:83:@37671.4]
  assign _T_81731 = _T_81730[10:0]; // @[Modules.scala 68:83:@37672.4]
  assign buffer_15_663 = $signed(_T_81731); // @[Modules.scala 68:83:@37673.4]
  assign _T_81733 = $signed(buffer_15_544) + $signed(buffer_10_545); // @[Modules.scala 68:83:@37675.4]
  assign _T_81734 = _T_81733[10:0]; // @[Modules.scala 68:83:@37676.4]
  assign buffer_15_664 = $signed(_T_81734); // @[Modules.scala 68:83:@37677.4]
  assign _T_81736 = $signed(buffer_15_546) + $signed(buffer_15_547); // @[Modules.scala 68:83:@37679.4]
  assign _T_81737 = _T_81736[10:0]; // @[Modules.scala 68:83:@37680.4]
  assign buffer_15_665 = $signed(_T_81737); // @[Modules.scala 68:83:@37681.4]
  assign _T_81739 = $signed(buffer_8_548) + $signed(buffer_15_549); // @[Modules.scala 68:83:@37683.4]
  assign _T_81740 = _T_81739[10:0]; // @[Modules.scala 68:83:@37684.4]
  assign buffer_15_666 = $signed(_T_81740); // @[Modules.scala 68:83:@37685.4]
  assign _T_81745 = $signed(buffer_15_552) + $signed(buffer_15_553); // @[Modules.scala 68:83:@37691.4]
  assign _T_81746 = _T_81745[10:0]; // @[Modules.scala 68:83:@37692.4]
  assign buffer_15_668 = $signed(_T_81746); // @[Modules.scala 68:83:@37693.4]
  assign _T_81748 = $signed(buffer_15_554) + $signed(buffer_8_555); // @[Modules.scala 68:83:@37695.4]
  assign _T_81749 = _T_81748[10:0]; // @[Modules.scala 68:83:@37696.4]
  assign buffer_15_669 = $signed(_T_81749); // @[Modules.scala 68:83:@37697.4]
  assign _T_81754 = $signed(buffer_5_558) + $signed(buffer_3_559); // @[Modules.scala 68:83:@37703.4]
  assign _T_81755 = _T_81754[10:0]; // @[Modules.scala 68:83:@37704.4]
  assign buffer_15_671 = $signed(_T_81755); // @[Modules.scala 68:83:@37705.4]
  assign _T_81757 = $signed(buffer_6_560) + $signed(buffer_15_561); // @[Modules.scala 68:83:@37707.4]
  assign _T_81758 = _T_81757[10:0]; // @[Modules.scala 68:83:@37708.4]
  assign buffer_15_672 = $signed(_T_81758); // @[Modules.scala 68:83:@37709.4]
  assign _T_81760 = $signed(buffer_15_562) + $signed(buffer_3_563); // @[Modules.scala 68:83:@37711.4]
  assign _T_81761 = _T_81760[10:0]; // @[Modules.scala 68:83:@37712.4]
  assign buffer_15_673 = $signed(_T_81761); // @[Modules.scala 68:83:@37713.4]
  assign _T_81766 = $signed(buffer_12_566) + $signed(buffer_15_567); // @[Modules.scala 68:83:@37719.4]
  assign _T_81767 = _T_81766[10:0]; // @[Modules.scala 68:83:@37720.4]
  assign buffer_15_675 = $signed(_T_81767); // @[Modules.scala 68:83:@37721.4]
  assign _T_81769 = $signed(buffer_15_568) + $signed(buffer_6_569); // @[Modules.scala 68:83:@37723.4]
  assign _T_81770 = _T_81769[10:0]; // @[Modules.scala 68:83:@37724.4]
  assign buffer_15_676 = $signed(_T_81770); // @[Modules.scala 68:83:@37725.4]
  assign _T_81772 = $signed(buffer_15_570) + $signed(buffer_1_571); // @[Modules.scala 68:83:@37727.4]
  assign _T_81773 = _T_81772[10:0]; // @[Modules.scala 68:83:@37728.4]
  assign buffer_15_677 = $signed(_T_81773); // @[Modules.scala 68:83:@37729.4]
  assign _T_81778 = $signed(buffer_3_574) + $signed(buffer_15_575); // @[Modules.scala 68:83:@37735.4]
  assign _T_81779 = _T_81778[10:0]; // @[Modules.scala 68:83:@37736.4]
  assign buffer_15_679 = $signed(_T_81779); // @[Modules.scala 68:83:@37737.4]
  assign _T_81796 = $signed(buffer_15_586) + $signed(buffer_13_587); // @[Modules.scala 68:83:@37759.4]
  assign _T_81797 = _T_81796[10:0]; // @[Modules.scala 68:83:@37760.4]
  assign buffer_15_685 = $signed(_T_81797); // @[Modules.scala 68:83:@37761.4]
  assign _T_81799 = $signed(buffer_15_588) + $signed(buffer_15_589); // @[Modules.scala 71:109:@37763.4]
  assign _T_81800 = _T_81799[10:0]; // @[Modules.scala 71:109:@37764.4]
  assign buffer_15_686 = $signed(_T_81800); // @[Modules.scala 71:109:@37765.4]
  assign _T_81802 = $signed(buffer_15_590) + $signed(buffer_15_591); // @[Modules.scala 71:109:@37767.4]
  assign _T_81803 = _T_81802[10:0]; // @[Modules.scala 71:109:@37768.4]
  assign buffer_15_687 = $signed(_T_81803); // @[Modules.scala 71:109:@37769.4]
  assign _T_81805 = $signed(buffer_15_592) + $signed(buffer_15_593); // @[Modules.scala 71:109:@37771.4]
  assign _T_81806 = _T_81805[10:0]; // @[Modules.scala 71:109:@37772.4]
  assign buffer_15_688 = $signed(_T_81806); // @[Modules.scala 71:109:@37773.4]
  assign _T_81808 = $signed(buffer_15_594) + $signed(buffer_15_595); // @[Modules.scala 71:109:@37775.4]
  assign _T_81809 = _T_81808[10:0]; // @[Modules.scala 71:109:@37776.4]
  assign buffer_15_689 = $signed(_T_81809); // @[Modules.scala 71:109:@37777.4]
  assign _T_81811 = $signed(buffer_1_596) + $signed(buffer_15_597); // @[Modules.scala 71:109:@37779.4]
  assign _T_81812 = _T_81811[10:0]; // @[Modules.scala 71:109:@37780.4]
  assign buffer_15_690 = $signed(_T_81812); // @[Modules.scala 71:109:@37781.4]
  assign _T_81814 = $signed(buffer_15_598) + $signed(buffer_15_599); // @[Modules.scala 71:109:@37783.4]
  assign _T_81815 = _T_81814[10:0]; // @[Modules.scala 71:109:@37784.4]
  assign buffer_15_691 = $signed(_T_81815); // @[Modules.scala 71:109:@37785.4]
  assign _T_81820 = $signed(buffer_15_602) + $signed(buffer_15_603); // @[Modules.scala 71:109:@37791.4]
  assign _T_81821 = _T_81820[10:0]; // @[Modules.scala 71:109:@37792.4]
  assign buffer_15_693 = $signed(_T_81821); // @[Modules.scala 71:109:@37793.4]
  assign _T_81823 = $signed(buffer_15_604) + $signed(buffer_15_605); // @[Modules.scala 71:109:@37795.4]
  assign _T_81824 = _T_81823[10:0]; // @[Modules.scala 71:109:@37796.4]
  assign buffer_15_694 = $signed(_T_81824); // @[Modules.scala 71:109:@37797.4]
  assign _T_81826 = $signed(buffer_15_606) + $signed(buffer_15_607); // @[Modules.scala 71:109:@37799.4]
  assign _T_81827 = _T_81826[10:0]; // @[Modules.scala 71:109:@37800.4]
  assign buffer_15_695 = $signed(_T_81827); // @[Modules.scala 71:109:@37801.4]
  assign _T_81829 = $signed(buffer_15_608) + $signed(buffer_15_609); // @[Modules.scala 71:109:@37803.4]
  assign _T_81830 = _T_81829[10:0]; // @[Modules.scala 71:109:@37804.4]
  assign buffer_15_696 = $signed(_T_81830); // @[Modules.scala 71:109:@37805.4]
  assign _T_81832 = $signed(buffer_15_610) + $signed(buffer_15_611); // @[Modules.scala 71:109:@37807.4]
  assign _T_81833 = _T_81832[10:0]; // @[Modules.scala 71:109:@37808.4]
  assign buffer_15_697 = $signed(_T_81833); // @[Modules.scala 71:109:@37809.4]
  assign _T_81835 = $signed(buffer_15_612) + $signed(buffer_15_613); // @[Modules.scala 71:109:@37811.4]
  assign _T_81836 = _T_81835[10:0]; // @[Modules.scala 71:109:@37812.4]
  assign buffer_15_698 = $signed(_T_81836); // @[Modules.scala 71:109:@37813.4]
  assign _T_81838 = $signed(buffer_15_614) + $signed(buffer_15_615); // @[Modules.scala 71:109:@37815.4]
  assign _T_81839 = _T_81838[10:0]; // @[Modules.scala 71:109:@37816.4]
  assign buffer_15_699 = $signed(_T_81839); // @[Modules.scala 71:109:@37817.4]
  assign _T_81841 = $signed(buffer_15_616) + $signed(buffer_15_617); // @[Modules.scala 71:109:@37819.4]
  assign _T_81842 = _T_81841[10:0]; // @[Modules.scala 71:109:@37820.4]
  assign buffer_15_700 = $signed(_T_81842); // @[Modules.scala 71:109:@37821.4]
  assign _T_81844 = $signed(buffer_15_618) + $signed(buffer_10_619); // @[Modules.scala 71:109:@37823.4]
  assign _T_81845 = _T_81844[10:0]; // @[Modules.scala 71:109:@37824.4]
  assign buffer_15_701 = $signed(_T_81845); // @[Modules.scala 71:109:@37825.4]
  assign _T_81847 = $signed(buffer_15_620) + $signed(buffer_15_621); // @[Modules.scala 71:109:@37827.4]
  assign _T_81848 = _T_81847[10:0]; // @[Modules.scala 71:109:@37828.4]
  assign buffer_15_702 = $signed(_T_81848); // @[Modules.scala 71:109:@37829.4]
  assign _T_81850 = $signed(buffer_0_593) + $signed(buffer_15_623); // @[Modules.scala 71:109:@37831.4]
  assign _T_81851 = _T_81850[10:0]; // @[Modules.scala 71:109:@37832.4]
  assign buffer_15_703 = $signed(_T_81851); // @[Modules.scala 71:109:@37833.4]
  assign _T_81853 = $signed(buffer_5_624) + $signed(buffer_15_625); // @[Modules.scala 71:109:@37835.4]
  assign _T_81854 = _T_81853[10:0]; // @[Modules.scala 71:109:@37836.4]
  assign buffer_15_704 = $signed(_T_81854); // @[Modules.scala 71:109:@37837.4]
  assign _T_81856 = $signed(buffer_15_626) + $signed(buffer_15_627); // @[Modules.scala 71:109:@37839.4]
  assign _T_81857 = _T_81856[10:0]; // @[Modules.scala 71:109:@37840.4]
  assign buffer_15_705 = $signed(_T_81857); // @[Modules.scala 71:109:@37841.4]
  assign _T_81859 = $signed(buffer_15_628) + $signed(buffer_15_629); // @[Modules.scala 71:109:@37843.4]
  assign _T_81860 = _T_81859[10:0]; // @[Modules.scala 71:109:@37844.4]
  assign buffer_15_706 = $signed(_T_81860); // @[Modules.scala 71:109:@37845.4]
  assign _T_81862 = $signed(buffer_15_630) + $signed(buffer_0_593); // @[Modules.scala 71:109:@37847.4]
  assign _T_81863 = _T_81862[10:0]; // @[Modules.scala 71:109:@37848.4]
  assign buffer_15_707 = $signed(_T_81863); // @[Modules.scala 71:109:@37849.4]
  assign _T_81865 = $signed(buffer_15_632) + $signed(buffer_15_633); // @[Modules.scala 71:109:@37851.4]
  assign _T_81866 = _T_81865[10:0]; // @[Modules.scala 71:109:@37852.4]
  assign buffer_15_708 = $signed(_T_81866); // @[Modules.scala 71:109:@37853.4]
  assign _T_81868 = $signed(buffer_15_634) + $signed(buffer_0_593); // @[Modules.scala 71:109:@37855.4]
  assign _T_81869 = _T_81868[10:0]; // @[Modules.scala 71:109:@37856.4]
  assign buffer_15_709 = $signed(_T_81869); // @[Modules.scala 71:109:@37857.4]
  assign _T_81871 = $signed(buffer_15_636) + $signed(buffer_8_637); // @[Modules.scala 71:109:@37859.4]
  assign _T_81872 = _T_81871[10:0]; // @[Modules.scala 71:109:@37860.4]
  assign buffer_15_710 = $signed(_T_81872); // @[Modules.scala 71:109:@37861.4]
  assign _T_81874 = $signed(buffer_0_593) + $signed(buffer_15_639); // @[Modules.scala 71:109:@37863.4]
  assign _T_81875 = _T_81874[10:0]; // @[Modules.scala 71:109:@37864.4]
  assign buffer_15_711 = $signed(_T_81875); // @[Modules.scala 71:109:@37865.4]
  assign _T_81877 = $signed(buffer_15_640) + $signed(buffer_8_641); // @[Modules.scala 71:109:@37867.4]
  assign _T_81878 = _T_81877[10:0]; // @[Modules.scala 71:109:@37868.4]
  assign buffer_15_712 = $signed(_T_81878); // @[Modules.scala 71:109:@37869.4]
  assign _T_81880 = $signed(buffer_15_642) + $signed(buffer_15_643); // @[Modules.scala 71:109:@37871.4]
  assign _T_81881 = _T_81880[10:0]; // @[Modules.scala 71:109:@37872.4]
  assign buffer_15_713 = $signed(_T_81881); // @[Modules.scala 71:109:@37873.4]
  assign _T_81883 = $signed(buffer_8_644) + $signed(buffer_15_645); // @[Modules.scala 71:109:@37875.4]
  assign _T_81884 = _T_81883[10:0]; // @[Modules.scala 71:109:@37876.4]
  assign buffer_15_714 = $signed(_T_81884); // @[Modules.scala 71:109:@37877.4]
  assign _T_81886 = $signed(buffer_15_646) + $signed(buffer_7_647); // @[Modules.scala 71:109:@37879.4]
  assign _T_81887 = _T_81886[10:0]; // @[Modules.scala 71:109:@37880.4]
  assign buffer_15_715 = $signed(_T_81887); // @[Modules.scala 71:109:@37881.4]
  assign _T_81889 = $signed(buffer_12_648) + $signed(buffer_15_649); // @[Modules.scala 71:109:@37883.4]
  assign _T_81890 = _T_81889[10:0]; // @[Modules.scala 71:109:@37884.4]
  assign buffer_15_716 = $signed(_T_81890); // @[Modules.scala 71:109:@37885.4]
  assign _T_81892 = $signed(buffer_15_650) + $signed(buffer_15_651); // @[Modules.scala 71:109:@37887.4]
  assign _T_81893 = _T_81892[10:0]; // @[Modules.scala 71:109:@37888.4]
  assign buffer_15_717 = $signed(_T_81893); // @[Modules.scala 71:109:@37889.4]
  assign _T_81895 = $signed(buffer_15_652) + $signed(buffer_15_653); // @[Modules.scala 71:109:@37891.4]
  assign _T_81896 = _T_81895[10:0]; // @[Modules.scala 71:109:@37892.4]
  assign buffer_15_718 = $signed(_T_81896); // @[Modules.scala 71:109:@37893.4]
  assign _T_81898 = $signed(buffer_12_654) + $signed(buffer_15_655); // @[Modules.scala 71:109:@37895.4]
  assign _T_81899 = _T_81898[10:0]; // @[Modules.scala 71:109:@37896.4]
  assign buffer_15_719 = $signed(_T_81899); // @[Modules.scala 71:109:@37897.4]
  assign _T_81901 = $signed(buffer_15_656) + $signed(buffer_8_657); // @[Modules.scala 71:109:@37899.4]
  assign _T_81902 = _T_81901[10:0]; // @[Modules.scala 71:109:@37900.4]
  assign buffer_15_720 = $signed(_T_81902); // @[Modules.scala 71:109:@37901.4]
  assign _T_81904 = $signed(buffer_2_658) + $signed(buffer_15_659); // @[Modules.scala 71:109:@37903.4]
  assign _T_81905 = _T_81904[10:0]; // @[Modules.scala 71:109:@37904.4]
  assign buffer_15_721 = $signed(_T_81905); // @[Modules.scala 71:109:@37905.4]
  assign _T_81907 = $signed(buffer_15_660) + $signed(buffer_15_661); // @[Modules.scala 71:109:@37907.4]
  assign _T_81908 = _T_81907[10:0]; // @[Modules.scala 71:109:@37908.4]
  assign buffer_15_722 = $signed(_T_81908); // @[Modules.scala 71:109:@37909.4]
  assign _T_81910 = $signed(buffer_15_662) + $signed(buffer_15_663); // @[Modules.scala 71:109:@37911.4]
  assign _T_81911 = _T_81910[10:0]; // @[Modules.scala 71:109:@37912.4]
  assign buffer_15_723 = $signed(_T_81911); // @[Modules.scala 71:109:@37913.4]
  assign _T_81913 = $signed(buffer_15_664) + $signed(buffer_15_665); // @[Modules.scala 71:109:@37915.4]
  assign _T_81914 = _T_81913[10:0]; // @[Modules.scala 71:109:@37916.4]
  assign buffer_15_724 = $signed(_T_81914); // @[Modules.scala 71:109:@37917.4]
  assign _T_81916 = $signed(buffer_15_666) + $signed(buffer_3_667); // @[Modules.scala 71:109:@37919.4]
  assign _T_81917 = _T_81916[10:0]; // @[Modules.scala 71:109:@37920.4]
  assign buffer_15_725 = $signed(_T_81917); // @[Modules.scala 71:109:@37921.4]
  assign _T_81919 = $signed(buffer_15_668) + $signed(buffer_15_669); // @[Modules.scala 71:109:@37923.4]
  assign _T_81920 = _T_81919[10:0]; // @[Modules.scala 71:109:@37924.4]
  assign buffer_15_726 = $signed(_T_81920); // @[Modules.scala 71:109:@37925.4]
  assign _T_81922 = $signed(buffer_0_670) + $signed(buffer_15_671); // @[Modules.scala 71:109:@37927.4]
  assign _T_81923 = _T_81922[10:0]; // @[Modules.scala 71:109:@37928.4]
  assign buffer_15_727 = $signed(_T_81923); // @[Modules.scala 71:109:@37929.4]
  assign _T_81925 = $signed(buffer_15_672) + $signed(buffer_15_673); // @[Modules.scala 71:109:@37931.4]
  assign _T_81926 = _T_81925[10:0]; // @[Modules.scala 71:109:@37932.4]
  assign buffer_15_728 = $signed(_T_81926); // @[Modules.scala 71:109:@37933.4]
  assign _T_81928 = $signed(buffer_0_593) + $signed(buffer_15_675); // @[Modules.scala 71:109:@37935.4]
  assign _T_81929 = _T_81928[10:0]; // @[Modules.scala 71:109:@37936.4]
  assign buffer_15_729 = $signed(_T_81929); // @[Modules.scala 71:109:@37937.4]
  assign _T_81931 = $signed(buffer_15_676) + $signed(buffer_15_677); // @[Modules.scala 71:109:@37939.4]
  assign _T_81932 = _T_81931[10:0]; // @[Modules.scala 71:109:@37940.4]
  assign buffer_15_730 = $signed(_T_81932); // @[Modules.scala 71:109:@37941.4]
  assign _T_81934 = $signed(buffer_9_678) + $signed(buffer_15_679); // @[Modules.scala 71:109:@37943.4]
  assign _T_81935 = _T_81934[10:0]; // @[Modules.scala 71:109:@37944.4]
  assign buffer_15_731 = $signed(_T_81935); // @[Modules.scala 71:109:@37945.4]
  assign _T_81937 = $signed(buffer_5_680) + $signed(buffer_3_681); // @[Modules.scala 71:109:@37947.4]
  assign _T_81938 = _T_81937[10:0]; // @[Modules.scala 71:109:@37948.4]
  assign buffer_15_732 = $signed(_T_81938); // @[Modules.scala 71:109:@37949.4]
  assign _T_81940 = $signed(buffer_8_682) + $signed(buffer_10_683); // @[Modules.scala 71:109:@37951.4]
  assign _T_81941 = _T_81940[10:0]; // @[Modules.scala 71:109:@37952.4]
  assign buffer_15_733 = $signed(_T_81941); // @[Modules.scala 71:109:@37953.4]
  assign _T_81943 = $signed(buffer_3_684) + $signed(buffer_15_685); // @[Modules.scala 71:109:@37955.4]
  assign _T_81944 = _T_81943[10:0]; // @[Modules.scala 71:109:@37956.4]
  assign buffer_15_734 = $signed(_T_81944); // @[Modules.scala 71:109:@37957.4]
  assign _T_81946 = $signed(buffer_15_686) + $signed(buffer_15_687); // @[Modules.scala 78:156:@37960.4]
  assign _T_81947 = _T_81946[10:0]; // @[Modules.scala 78:156:@37961.4]
  assign buffer_15_736 = $signed(_T_81947); // @[Modules.scala 78:156:@37962.4]
  assign _T_81949 = $signed(buffer_15_736) + $signed(buffer_15_688); // @[Modules.scala 78:156:@37964.4]
  assign _T_81950 = _T_81949[10:0]; // @[Modules.scala 78:156:@37965.4]
  assign buffer_15_737 = $signed(_T_81950); // @[Modules.scala 78:156:@37966.4]
  assign _T_81952 = $signed(buffer_15_737) + $signed(buffer_15_689); // @[Modules.scala 78:156:@37968.4]
  assign _T_81953 = _T_81952[10:0]; // @[Modules.scala 78:156:@37969.4]
  assign buffer_15_738 = $signed(_T_81953); // @[Modules.scala 78:156:@37970.4]
  assign _T_81955 = $signed(buffer_15_738) + $signed(buffer_15_690); // @[Modules.scala 78:156:@37972.4]
  assign _T_81956 = _T_81955[10:0]; // @[Modules.scala 78:156:@37973.4]
  assign buffer_15_739 = $signed(_T_81956); // @[Modules.scala 78:156:@37974.4]
  assign _T_81958 = $signed(buffer_15_739) + $signed(buffer_15_691); // @[Modules.scala 78:156:@37976.4]
  assign _T_81959 = _T_81958[10:0]; // @[Modules.scala 78:156:@37977.4]
  assign buffer_15_740 = $signed(_T_81959); // @[Modules.scala 78:156:@37978.4]
  assign _T_81961 = $signed(buffer_15_740) + $signed(buffer_12_692); // @[Modules.scala 78:156:@37980.4]
  assign _T_81962 = _T_81961[10:0]; // @[Modules.scala 78:156:@37981.4]
  assign buffer_15_741 = $signed(_T_81962); // @[Modules.scala 78:156:@37982.4]
  assign _T_81964 = $signed(buffer_15_741) + $signed(buffer_15_693); // @[Modules.scala 78:156:@37984.4]
  assign _T_81965 = _T_81964[10:0]; // @[Modules.scala 78:156:@37985.4]
  assign buffer_15_742 = $signed(_T_81965); // @[Modules.scala 78:156:@37986.4]
  assign _T_81967 = $signed(buffer_15_742) + $signed(buffer_15_694); // @[Modules.scala 78:156:@37988.4]
  assign _T_81968 = _T_81967[10:0]; // @[Modules.scala 78:156:@37989.4]
  assign buffer_15_743 = $signed(_T_81968); // @[Modules.scala 78:156:@37990.4]
  assign _T_81970 = $signed(buffer_15_743) + $signed(buffer_15_695); // @[Modules.scala 78:156:@37992.4]
  assign _T_81971 = _T_81970[10:0]; // @[Modules.scala 78:156:@37993.4]
  assign buffer_15_744 = $signed(_T_81971); // @[Modules.scala 78:156:@37994.4]
  assign _T_81973 = $signed(buffer_15_744) + $signed(buffer_15_696); // @[Modules.scala 78:156:@37996.4]
  assign _T_81974 = _T_81973[10:0]; // @[Modules.scala 78:156:@37997.4]
  assign buffer_15_745 = $signed(_T_81974); // @[Modules.scala 78:156:@37998.4]
  assign _T_81976 = $signed(buffer_15_745) + $signed(buffer_15_697); // @[Modules.scala 78:156:@38000.4]
  assign _T_81977 = _T_81976[10:0]; // @[Modules.scala 78:156:@38001.4]
  assign buffer_15_746 = $signed(_T_81977); // @[Modules.scala 78:156:@38002.4]
  assign _T_81979 = $signed(buffer_15_746) + $signed(buffer_15_698); // @[Modules.scala 78:156:@38004.4]
  assign _T_81980 = _T_81979[10:0]; // @[Modules.scala 78:156:@38005.4]
  assign buffer_15_747 = $signed(_T_81980); // @[Modules.scala 78:156:@38006.4]
  assign _T_81982 = $signed(buffer_15_747) + $signed(buffer_15_699); // @[Modules.scala 78:156:@38008.4]
  assign _T_81983 = _T_81982[10:0]; // @[Modules.scala 78:156:@38009.4]
  assign buffer_15_748 = $signed(_T_81983); // @[Modules.scala 78:156:@38010.4]
  assign _T_81985 = $signed(buffer_15_748) + $signed(buffer_15_700); // @[Modules.scala 78:156:@38012.4]
  assign _T_81986 = _T_81985[10:0]; // @[Modules.scala 78:156:@38013.4]
  assign buffer_15_749 = $signed(_T_81986); // @[Modules.scala 78:156:@38014.4]
  assign _T_81988 = $signed(buffer_15_749) + $signed(buffer_15_701); // @[Modules.scala 78:156:@38016.4]
  assign _T_81989 = _T_81988[10:0]; // @[Modules.scala 78:156:@38017.4]
  assign buffer_15_750 = $signed(_T_81989); // @[Modules.scala 78:156:@38018.4]
  assign _T_81991 = $signed(buffer_15_750) + $signed(buffer_15_702); // @[Modules.scala 78:156:@38020.4]
  assign _T_81992 = _T_81991[10:0]; // @[Modules.scala 78:156:@38021.4]
  assign buffer_15_751 = $signed(_T_81992); // @[Modules.scala 78:156:@38022.4]
  assign _T_81994 = $signed(buffer_15_751) + $signed(buffer_15_703); // @[Modules.scala 78:156:@38024.4]
  assign _T_81995 = _T_81994[10:0]; // @[Modules.scala 78:156:@38025.4]
  assign buffer_15_752 = $signed(_T_81995); // @[Modules.scala 78:156:@38026.4]
  assign _T_81997 = $signed(buffer_15_752) + $signed(buffer_15_704); // @[Modules.scala 78:156:@38028.4]
  assign _T_81998 = _T_81997[10:0]; // @[Modules.scala 78:156:@38029.4]
  assign buffer_15_753 = $signed(_T_81998); // @[Modules.scala 78:156:@38030.4]
  assign _T_82000 = $signed(buffer_15_753) + $signed(buffer_15_705); // @[Modules.scala 78:156:@38032.4]
  assign _T_82001 = _T_82000[10:0]; // @[Modules.scala 78:156:@38033.4]
  assign buffer_15_754 = $signed(_T_82001); // @[Modules.scala 78:156:@38034.4]
  assign _T_82003 = $signed(buffer_15_754) + $signed(buffer_15_706); // @[Modules.scala 78:156:@38036.4]
  assign _T_82004 = _T_82003[10:0]; // @[Modules.scala 78:156:@38037.4]
  assign buffer_15_755 = $signed(_T_82004); // @[Modules.scala 78:156:@38038.4]
  assign _T_82006 = $signed(buffer_15_755) + $signed(buffer_15_707); // @[Modules.scala 78:156:@38040.4]
  assign _T_82007 = _T_82006[10:0]; // @[Modules.scala 78:156:@38041.4]
  assign buffer_15_756 = $signed(_T_82007); // @[Modules.scala 78:156:@38042.4]
  assign _T_82009 = $signed(buffer_15_756) + $signed(buffer_15_708); // @[Modules.scala 78:156:@38044.4]
  assign _T_82010 = _T_82009[10:0]; // @[Modules.scala 78:156:@38045.4]
  assign buffer_15_757 = $signed(_T_82010); // @[Modules.scala 78:156:@38046.4]
  assign _T_82012 = $signed(buffer_15_757) + $signed(buffer_15_709); // @[Modules.scala 78:156:@38048.4]
  assign _T_82013 = _T_82012[10:0]; // @[Modules.scala 78:156:@38049.4]
  assign buffer_15_758 = $signed(_T_82013); // @[Modules.scala 78:156:@38050.4]
  assign _T_82015 = $signed(buffer_15_758) + $signed(buffer_15_710); // @[Modules.scala 78:156:@38052.4]
  assign _T_82016 = _T_82015[10:0]; // @[Modules.scala 78:156:@38053.4]
  assign buffer_15_759 = $signed(_T_82016); // @[Modules.scala 78:156:@38054.4]
  assign _T_82018 = $signed(buffer_15_759) + $signed(buffer_15_711); // @[Modules.scala 78:156:@38056.4]
  assign _T_82019 = _T_82018[10:0]; // @[Modules.scala 78:156:@38057.4]
  assign buffer_15_760 = $signed(_T_82019); // @[Modules.scala 78:156:@38058.4]
  assign _T_82021 = $signed(buffer_15_760) + $signed(buffer_15_712); // @[Modules.scala 78:156:@38060.4]
  assign _T_82022 = _T_82021[10:0]; // @[Modules.scala 78:156:@38061.4]
  assign buffer_15_761 = $signed(_T_82022); // @[Modules.scala 78:156:@38062.4]
  assign _T_82024 = $signed(buffer_15_761) + $signed(buffer_15_713); // @[Modules.scala 78:156:@38064.4]
  assign _T_82025 = _T_82024[10:0]; // @[Modules.scala 78:156:@38065.4]
  assign buffer_15_762 = $signed(_T_82025); // @[Modules.scala 78:156:@38066.4]
  assign _T_82027 = $signed(buffer_15_762) + $signed(buffer_15_714); // @[Modules.scala 78:156:@38068.4]
  assign _T_82028 = _T_82027[10:0]; // @[Modules.scala 78:156:@38069.4]
  assign buffer_15_763 = $signed(_T_82028); // @[Modules.scala 78:156:@38070.4]
  assign _T_82030 = $signed(buffer_15_763) + $signed(buffer_15_715); // @[Modules.scala 78:156:@38072.4]
  assign _T_82031 = _T_82030[10:0]; // @[Modules.scala 78:156:@38073.4]
  assign buffer_15_764 = $signed(_T_82031); // @[Modules.scala 78:156:@38074.4]
  assign _T_82033 = $signed(buffer_15_764) + $signed(buffer_15_716); // @[Modules.scala 78:156:@38076.4]
  assign _T_82034 = _T_82033[10:0]; // @[Modules.scala 78:156:@38077.4]
  assign buffer_15_765 = $signed(_T_82034); // @[Modules.scala 78:156:@38078.4]
  assign _T_82036 = $signed(buffer_15_765) + $signed(buffer_15_717); // @[Modules.scala 78:156:@38080.4]
  assign _T_82037 = _T_82036[10:0]; // @[Modules.scala 78:156:@38081.4]
  assign buffer_15_766 = $signed(_T_82037); // @[Modules.scala 78:156:@38082.4]
  assign _T_82039 = $signed(buffer_15_766) + $signed(buffer_15_718); // @[Modules.scala 78:156:@38084.4]
  assign _T_82040 = _T_82039[10:0]; // @[Modules.scala 78:156:@38085.4]
  assign buffer_15_767 = $signed(_T_82040); // @[Modules.scala 78:156:@38086.4]
  assign _T_82042 = $signed(buffer_15_767) + $signed(buffer_15_719); // @[Modules.scala 78:156:@38088.4]
  assign _T_82043 = _T_82042[10:0]; // @[Modules.scala 78:156:@38089.4]
  assign buffer_15_768 = $signed(_T_82043); // @[Modules.scala 78:156:@38090.4]
  assign _T_82045 = $signed(buffer_15_768) + $signed(buffer_15_720); // @[Modules.scala 78:156:@38092.4]
  assign _T_82046 = _T_82045[10:0]; // @[Modules.scala 78:156:@38093.4]
  assign buffer_15_769 = $signed(_T_82046); // @[Modules.scala 78:156:@38094.4]
  assign _T_82048 = $signed(buffer_15_769) + $signed(buffer_15_721); // @[Modules.scala 78:156:@38096.4]
  assign _T_82049 = _T_82048[10:0]; // @[Modules.scala 78:156:@38097.4]
  assign buffer_15_770 = $signed(_T_82049); // @[Modules.scala 78:156:@38098.4]
  assign _T_82051 = $signed(buffer_15_770) + $signed(buffer_15_722); // @[Modules.scala 78:156:@38100.4]
  assign _T_82052 = _T_82051[10:0]; // @[Modules.scala 78:156:@38101.4]
  assign buffer_15_771 = $signed(_T_82052); // @[Modules.scala 78:156:@38102.4]
  assign _T_82054 = $signed(buffer_15_771) + $signed(buffer_15_723); // @[Modules.scala 78:156:@38104.4]
  assign _T_82055 = _T_82054[10:0]; // @[Modules.scala 78:156:@38105.4]
  assign buffer_15_772 = $signed(_T_82055); // @[Modules.scala 78:156:@38106.4]
  assign _T_82057 = $signed(buffer_15_772) + $signed(buffer_15_724); // @[Modules.scala 78:156:@38108.4]
  assign _T_82058 = _T_82057[10:0]; // @[Modules.scala 78:156:@38109.4]
  assign buffer_15_773 = $signed(_T_82058); // @[Modules.scala 78:156:@38110.4]
  assign _T_82060 = $signed(buffer_15_773) + $signed(buffer_15_725); // @[Modules.scala 78:156:@38112.4]
  assign _T_82061 = _T_82060[10:0]; // @[Modules.scala 78:156:@38113.4]
  assign buffer_15_774 = $signed(_T_82061); // @[Modules.scala 78:156:@38114.4]
  assign _T_82063 = $signed(buffer_15_774) + $signed(buffer_15_726); // @[Modules.scala 78:156:@38116.4]
  assign _T_82064 = _T_82063[10:0]; // @[Modules.scala 78:156:@38117.4]
  assign buffer_15_775 = $signed(_T_82064); // @[Modules.scala 78:156:@38118.4]
  assign _T_82066 = $signed(buffer_15_775) + $signed(buffer_15_727); // @[Modules.scala 78:156:@38120.4]
  assign _T_82067 = _T_82066[10:0]; // @[Modules.scala 78:156:@38121.4]
  assign buffer_15_776 = $signed(_T_82067); // @[Modules.scala 78:156:@38122.4]
  assign _T_82069 = $signed(buffer_15_776) + $signed(buffer_15_728); // @[Modules.scala 78:156:@38124.4]
  assign _T_82070 = _T_82069[10:0]; // @[Modules.scala 78:156:@38125.4]
  assign buffer_15_777 = $signed(_T_82070); // @[Modules.scala 78:156:@38126.4]
  assign _T_82072 = $signed(buffer_15_777) + $signed(buffer_15_729); // @[Modules.scala 78:156:@38128.4]
  assign _T_82073 = _T_82072[10:0]; // @[Modules.scala 78:156:@38129.4]
  assign buffer_15_778 = $signed(_T_82073); // @[Modules.scala 78:156:@38130.4]
  assign _T_82075 = $signed(buffer_15_778) + $signed(buffer_15_730); // @[Modules.scala 78:156:@38132.4]
  assign _T_82076 = _T_82075[10:0]; // @[Modules.scala 78:156:@38133.4]
  assign buffer_15_779 = $signed(_T_82076); // @[Modules.scala 78:156:@38134.4]
  assign _T_82078 = $signed(buffer_15_779) + $signed(buffer_15_731); // @[Modules.scala 78:156:@38136.4]
  assign _T_82079 = _T_82078[10:0]; // @[Modules.scala 78:156:@38137.4]
  assign buffer_15_780 = $signed(_T_82079); // @[Modules.scala 78:156:@38138.4]
  assign _T_82081 = $signed(buffer_15_780) + $signed(buffer_15_732); // @[Modules.scala 78:156:@38140.4]
  assign _T_82082 = _T_82081[10:0]; // @[Modules.scala 78:156:@38141.4]
  assign buffer_15_781 = $signed(_T_82082); // @[Modules.scala 78:156:@38142.4]
  assign _T_82084 = $signed(buffer_15_781) + $signed(buffer_15_733); // @[Modules.scala 78:156:@38144.4]
  assign _T_82085 = _T_82084[10:0]; // @[Modules.scala 78:156:@38145.4]
  assign buffer_15_782 = $signed(_T_82085); // @[Modules.scala 78:156:@38146.4]
  assign _T_82087 = $signed(buffer_15_782) + $signed(buffer_15_734); // @[Modules.scala 78:156:@38148.4]
  assign _T_82088 = _T_82087[10:0]; // @[Modules.scala 78:156:@38149.4]
  assign buffer_15_783 = $signed(_T_82088); // @[Modules.scala 78:156:@38150.4]
  assign io_out_0 = buffer_0_783;
  assign io_out_1 = buffer_1_783;
  assign io_out_2 = buffer_2_783;
  assign io_out_3 = buffer_3_783;
  assign io_out_4 = buffer_4_783;
  assign io_out_5 = buffer_5_783;
  assign io_out_6 = buffer_6_783;
  assign io_out_7 = buffer_7_783;
  assign io_out_8 = buffer_8_783;
  assign io_out_9 = buffer_9_783;
  assign io_out_10 = buffer_10_783;
  assign io_out_11 = buffer_11_783;
  assign io_out_12 = buffer_12_783;
  assign io_out_13 = buffer_13_783;
  assign io_out_14 = buffer_14_783;
  assign io_out_15 = buffer_15_783;
endmodule
module ShifBatchNorm( // @[:@38154.2]
  input  [10:0] io_in_0, // @[:@38157.4]
  input  [10:0] io_in_1, // @[:@38157.4]
  input  [10:0] io_in_2, // @[:@38157.4]
  input  [10:0] io_in_3, // @[:@38157.4]
  input  [10:0] io_in_4, // @[:@38157.4]
  input  [10:0] io_in_5, // @[:@38157.4]
  input  [10:0] io_in_6, // @[:@38157.4]
  input  [10:0] io_in_7, // @[:@38157.4]
  input  [10:0] io_in_8, // @[:@38157.4]
  input  [10:0] io_in_9, // @[:@38157.4]
  input  [10:0] io_in_10, // @[:@38157.4]
  input  [10:0] io_in_11, // @[:@38157.4]
  input  [10:0] io_in_12, // @[:@38157.4]
  input  [10:0] io_in_13, // @[:@38157.4]
  input  [10:0] io_in_14, // @[:@38157.4]
  input  [10:0] io_in_15, // @[:@38157.4]
  output [10:0] io_out_0, // @[:@38157.4]
  output [10:0] io_out_1, // @[:@38157.4]
  output [10:0] io_out_2, // @[:@38157.4]
  output [10:0] io_out_3, // @[:@38157.4]
  output [10:0] io_out_4, // @[:@38157.4]
  output [10:0] io_out_5, // @[:@38157.4]
  output [10:0] io_out_6, // @[:@38157.4]
  output [10:0] io_out_7, // @[:@38157.4]
  output [10:0] io_out_8, // @[:@38157.4]
  output [10:0] io_out_9, // @[:@38157.4]
  output [10:0] io_out_10, // @[:@38157.4]
  output [10:0] io_out_11, // @[:@38157.4]
  output [10:0] io_out_12, // @[:@38157.4]
  output [10:0] io_out_13, // @[:@38157.4]
  output [10:0] io_out_14, // @[:@38157.4]
  output [10:0] io_out_15 // @[:@38157.4]
);
  wire [11:0] _T_108; // @[Modules.scala 132:28:@38162.4]
  wire [10:0] _T_109; // @[Modules.scala 132:28:@38163.4]
  wire [10:0] c_x_0; // @[Modules.scala 132:28:@38164.4]
  wire [25:0] _GEN_0; // @[Modules.scala 137:32:@38166.4]
  wire [25:0] _T_112; // @[Modules.scala 137:32:@38166.4]
  wire [10:0] _GEN_1; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_0; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_2; // @[Modules.scala 139:37:@38168.4]
  wire [25:0] _T_114; // @[Modules.scala 139:37:@38168.4]
  wire [10:0] _GEN_3; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_0; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_116; // @[Modules.scala 140:38:@38170.4]
  wire [10:0] _T_117; // @[Modules.scala 140:38:@38171.4]
  wire [10:0] _T_118; // @[Modules.scala 140:38:@38172.4]
  wire [11:0] _T_120; // @[Modules.scala 132:28:@38174.4]
  wire [10:0] _T_121; // @[Modules.scala 132:28:@38175.4]
  wire [10:0] c_x_1; // @[Modules.scala 132:28:@38176.4]
  wire [25:0] _GEN_4; // @[Modules.scala 137:32:@38178.4]
  wire [25:0] _T_124; // @[Modules.scala 137:32:@38178.4]
  wire [10:0] _GEN_5; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_1; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_6; // @[Modules.scala 139:37:@38180.4]
  wire [25:0] _T_126; // @[Modules.scala 139:37:@38180.4]
  wire [10:0] _GEN_7; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_1; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_128; // @[Modules.scala 140:38:@38182.4]
  wire [10:0] _T_129; // @[Modules.scala 140:38:@38183.4]
  wire [10:0] _T_130; // @[Modules.scala 140:38:@38184.4]
  wire [11:0] _T_132; // @[Modules.scala 132:28:@38186.4]
  wire [10:0] _T_133; // @[Modules.scala 132:28:@38187.4]
  wire [10:0] c_x_2; // @[Modules.scala 132:28:@38188.4]
  wire [25:0] _GEN_8; // @[Modules.scala 137:32:@38190.4]
  wire [25:0] _T_136; // @[Modules.scala 137:32:@38190.4]
  wire [10:0] _GEN_9; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_2; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_10; // @[Modules.scala 139:37:@38192.4]
  wire [25:0] _T_138; // @[Modules.scala 139:37:@38192.4]
  wire [10:0] _GEN_11; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_2; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_140; // @[Modules.scala 140:38:@38194.4]
  wire [10:0] _T_141; // @[Modules.scala 140:38:@38195.4]
  wire [10:0] _T_142; // @[Modules.scala 140:38:@38196.4]
  wire [11:0] _T_144; // @[Modules.scala 132:28:@38198.4]
  wire [10:0] _T_145; // @[Modules.scala 132:28:@38199.4]
  wire [10:0] c_x_3; // @[Modules.scala 132:28:@38200.4]
  wire [25:0] _GEN_12; // @[Modules.scala 137:32:@38202.4]
  wire [25:0] _T_148; // @[Modules.scala 137:32:@38202.4]
  wire [10:0] _GEN_13; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_3; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_14; // @[Modules.scala 139:37:@38204.4]
  wire [25:0] _T_150; // @[Modules.scala 139:37:@38204.4]
  wire [10:0] _GEN_15; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_3; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_152; // @[Modules.scala 140:38:@38206.4]
  wire [10:0] _T_153; // @[Modules.scala 140:38:@38207.4]
  wire [10:0] _T_154; // @[Modules.scala 140:38:@38208.4]
  wire [11:0] _T_156; // @[Modules.scala 132:28:@38210.4]
  wire [10:0] _T_157; // @[Modules.scala 132:28:@38211.4]
  wire [10:0] c_x_4; // @[Modules.scala 132:28:@38212.4]
  wire [25:0] _GEN_16; // @[Modules.scala 137:32:@38214.4]
  wire [25:0] _T_160; // @[Modules.scala 137:32:@38214.4]
  wire [10:0] _GEN_17; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_4; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_18; // @[Modules.scala 139:37:@38216.4]
  wire [25:0] _T_162; // @[Modules.scala 139:37:@38216.4]
  wire [10:0] _GEN_19; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_4; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_164; // @[Modules.scala 140:38:@38218.4]
  wire [10:0] _T_165; // @[Modules.scala 140:38:@38219.4]
  wire [10:0] _T_166; // @[Modules.scala 140:38:@38220.4]
  wire [11:0] _T_168; // @[Modules.scala 132:28:@38222.4]
  wire [10:0] _T_169; // @[Modules.scala 132:28:@38223.4]
  wire [10:0] c_x_5; // @[Modules.scala 132:28:@38224.4]
  wire [25:0] _GEN_20; // @[Modules.scala 137:32:@38226.4]
  wire [25:0] _T_172; // @[Modules.scala 137:32:@38226.4]
  wire [10:0] _GEN_21; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_5; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_22; // @[Modules.scala 139:37:@38228.4]
  wire [25:0] _T_174; // @[Modules.scala 139:37:@38228.4]
  wire [10:0] _GEN_23; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_5; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_176; // @[Modules.scala 140:38:@38230.4]
  wire [10:0] _T_177; // @[Modules.scala 140:38:@38231.4]
  wire [10:0] _T_178; // @[Modules.scala 140:38:@38232.4]
  wire [11:0] _T_180; // @[Modules.scala 132:28:@38234.4]
  wire [10:0] _T_181; // @[Modules.scala 132:28:@38235.4]
  wire [10:0] c_x_6; // @[Modules.scala 132:28:@38236.4]
  wire [25:0] _GEN_24; // @[Modules.scala 137:32:@38238.4]
  wire [25:0] _T_184; // @[Modules.scala 137:32:@38238.4]
  wire [10:0] _GEN_25; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_6; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_26; // @[Modules.scala 139:37:@38240.4]
  wire [25:0] _T_186; // @[Modules.scala 139:37:@38240.4]
  wire [10:0] _GEN_27; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_6; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_188; // @[Modules.scala 140:38:@38242.4]
  wire [10:0] _T_189; // @[Modules.scala 140:38:@38243.4]
  wire [10:0] _T_190; // @[Modules.scala 140:38:@38244.4]
  wire [11:0] _T_192; // @[Modules.scala 132:28:@38246.4]
  wire [10:0] _T_193; // @[Modules.scala 132:28:@38247.4]
  wire [10:0] c_x_7; // @[Modules.scala 132:28:@38248.4]
  wire [25:0] _GEN_28; // @[Modules.scala 137:32:@38250.4]
  wire [25:0] _T_196; // @[Modules.scala 137:32:@38250.4]
  wire [10:0] _GEN_29; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_7; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_30; // @[Modules.scala 139:37:@38252.4]
  wire [25:0] _T_198; // @[Modules.scala 139:37:@38252.4]
  wire [10:0] _GEN_31; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_7; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_200; // @[Modules.scala 140:38:@38254.4]
  wire [10:0] _T_201; // @[Modules.scala 140:38:@38255.4]
  wire [10:0] _T_202; // @[Modules.scala 140:38:@38256.4]
  wire [11:0] _T_204; // @[Modules.scala 132:28:@38258.4]
  wire [10:0] _T_205; // @[Modules.scala 132:28:@38259.4]
  wire [10:0] c_x_8; // @[Modules.scala 132:28:@38260.4]
  wire [25:0] _GEN_32; // @[Modules.scala 137:32:@38262.4]
  wire [25:0] _T_208; // @[Modules.scala 137:32:@38262.4]
  wire [10:0] _GEN_33; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_8; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_34; // @[Modules.scala 139:37:@38264.4]
  wire [25:0] _T_210; // @[Modules.scala 139:37:@38264.4]
  wire [10:0] _GEN_35; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_8; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_212; // @[Modules.scala 140:38:@38266.4]
  wire [10:0] _T_213; // @[Modules.scala 140:38:@38267.4]
  wire [10:0] _T_214; // @[Modules.scala 140:38:@38268.4]
  wire [11:0] _T_216; // @[Modules.scala 132:28:@38270.4]
  wire [10:0] _T_217; // @[Modules.scala 132:28:@38271.4]
  wire [10:0] c_x_9; // @[Modules.scala 132:28:@38272.4]
  wire [25:0] _GEN_36; // @[Modules.scala 137:32:@38274.4]
  wire [25:0] _T_220; // @[Modules.scala 137:32:@38274.4]
  wire [10:0] _GEN_37; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_9; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_38; // @[Modules.scala 139:37:@38276.4]
  wire [25:0] _T_222; // @[Modules.scala 139:37:@38276.4]
  wire [10:0] _GEN_39; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_9; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_224; // @[Modules.scala 140:38:@38278.4]
  wire [10:0] _T_225; // @[Modules.scala 140:38:@38279.4]
  wire [10:0] _T_226; // @[Modules.scala 140:38:@38280.4]
  wire [11:0] _T_228; // @[Modules.scala 132:28:@38282.4]
  wire [10:0] _T_229; // @[Modules.scala 132:28:@38283.4]
  wire [10:0] c_x_10; // @[Modules.scala 132:28:@38284.4]
  wire [25:0] _GEN_40; // @[Modules.scala 137:32:@38286.4]
  wire [25:0] _T_232; // @[Modules.scala 137:32:@38286.4]
  wire [10:0] _GEN_41; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_10; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_42; // @[Modules.scala 139:37:@38288.4]
  wire [25:0] _T_234; // @[Modules.scala 139:37:@38288.4]
  wire [10:0] _GEN_43; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_10; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_236; // @[Modules.scala 140:38:@38290.4]
  wire [10:0] _T_237; // @[Modules.scala 140:38:@38291.4]
  wire [10:0] _T_238; // @[Modules.scala 140:38:@38292.4]
  wire [11:0] _T_240; // @[Modules.scala 132:28:@38294.4]
  wire [10:0] _T_241; // @[Modules.scala 132:28:@38295.4]
  wire [10:0] c_x_11; // @[Modules.scala 132:28:@38296.4]
  wire [25:0] _GEN_44; // @[Modules.scala 137:32:@38298.4]
  wire [25:0] _T_244; // @[Modules.scala 137:32:@38298.4]
  wire [10:0] _GEN_45; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_11; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_46; // @[Modules.scala 139:37:@38300.4]
  wire [25:0] _T_246; // @[Modules.scala 139:37:@38300.4]
  wire [10:0] _GEN_47; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_11; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_248; // @[Modules.scala 140:38:@38302.4]
  wire [10:0] _T_249; // @[Modules.scala 140:38:@38303.4]
  wire [10:0] _T_250; // @[Modules.scala 140:38:@38304.4]
  wire [11:0] _T_252; // @[Modules.scala 132:28:@38306.4]
  wire [10:0] _T_253; // @[Modules.scala 132:28:@38307.4]
  wire [10:0] c_x_12; // @[Modules.scala 132:28:@38308.4]
  wire [25:0] _GEN_48; // @[Modules.scala 137:32:@38310.4]
  wire [25:0] _T_256; // @[Modules.scala 137:32:@38310.4]
  wire [10:0] _GEN_49; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_12; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_50; // @[Modules.scala 139:37:@38312.4]
  wire [25:0] _T_258; // @[Modules.scala 139:37:@38312.4]
  wire [10:0] _GEN_51; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_12; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_260; // @[Modules.scala 140:38:@38314.4]
  wire [10:0] _T_261; // @[Modules.scala 140:38:@38315.4]
  wire [10:0] _T_262; // @[Modules.scala 140:38:@38316.4]
  wire [11:0] _T_264; // @[Modules.scala 132:28:@38318.4]
  wire [10:0] _T_265; // @[Modules.scala 132:28:@38319.4]
  wire [10:0] c_x_13; // @[Modules.scala 132:28:@38320.4]
  wire [25:0] _GEN_52; // @[Modules.scala 137:32:@38322.4]
  wire [25:0] _T_268; // @[Modules.scala 137:32:@38322.4]
  wire [10:0] _GEN_53; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_13; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_54; // @[Modules.scala 139:37:@38324.4]
  wire [25:0] _T_270; // @[Modules.scala 139:37:@38324.4]
  wire [10:0] _GEN_55; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_13; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_272; // @[Modules.scala 140:38:@38326.4]
  wire [10:0] _T_273; // @[Modules.scala 140:38:@38327.4]
  wire [10:0] _T_274; // @[Modules.scala 140:38:@38328.4]
  wire [11:0] _T_276; // @[Modules.scala 132:28:@38330.4]
  wire [10:0] _T_277; // @[Modules.scala 132:28:@38331.4]
  wire [10:0] c_x_14; // @[Modules.scala 132:28:@38332.4]
  wire [25:0] _GEN_56; // @[Modules.scala 137:32:@38334.4]
  wire [25:0] _T_280; // @[Modules.scala 137:32:@38334.4]
  wire [10:0] _GEN_57; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_14; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_58; // @[Modules.scala 139:37:@38336.4]
  wire [25:0] _T_282; // @[Modules.scala 139:37:@38336.4]
  wire [10:0] _GEN_59; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_14; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_284; // @[Modules.scala 140:38:@38338.4]
  wire [10:0] _T_285; // @[Modules.scala 140:38:@38339.4]
  wire [10:0] _T_286; // @[Modules.scala 140:38:@38340.4]
  wire [11:0] _T_288; // @[Modules.scala 132:28:@38342.4]
  wire [10:0] _T_289; // @[Modules.scala 132:28:@38343.4]
  wire [10:0] c_x_15; // @[Modules.scala 132:28:@38344.4]
  wire [25:0] _GEN_60; // @[Modules.scala 137:32:@38346.4]
  wire [25:0] _T_292; // @[Modules.scala 137:32:@38346.4]
  wire [10:0] _GEN_61; // @[Modules.scala 129:21:@38160.4]
  wire [10:0] x_hat_15; // @[Modules.scala 129:21:@38160.4]
  wire [25:0] _GEN_62; // @[Modules.scala 139:37:@38348.4]
  wire [25:0] _T_294; // @[Modules.scala 139:37:@38348.4]
  wire [10:0] _GEN_63; // @[Modules.scala 130:28:@38161.4]
  wire [10:0] normed_x_hat_15; // @[Modules.scala 130:28:@38161.4]
  wire [11:0] _T_296; // @[Modules.scala 140:38:@38350.4]
  wire [10:0] _T_297; // @[Modules.scala 140:38:@38351.4]
  wire [10:0] _T_298; // @[Modules.scala 140:38:@38352.4]
  assign _T_108 = $signed(io_in_0) - $signed(11'sh49); // @[Modules.scala 132:28:@38162.4]
  assign _T_109 = _T_108[10:0]; // @[Modules.scala 132:28:@38163.4]
  assign c_x_0 = $signed(_T_109); // @[Modules.scala 132:28:@38164.4]
  assign _GEN_0 = {{15{c_x_0[10]}},c_x_0}; // @[Modules.scala 137:32:@38166.4]
  assign _T_112 = $signed(_GEN_0) << 4'h4; // @[Modules.scala 137:32:@38166.4]
  assign _GEN_1 = _T_112[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_0 = $signed(_GEN_1); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_2 = {{15{x_hat_0[10]}},x_hat_0}; // @[Modules.scala 139:37:@38168.4]
  assign _T_114 = $signed(_GEN_2) << 4'h2; // @[Modules.scala 139:37:@38168.4]
  assign _GEN_3 = _T_114[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_0 = $signed(_GEN_3); // @[Modules.scala 130:28:@38161.4]
  assign _T_116 = $signed(normed_x_hat_0) + $signed(-11'shf); // @[Modules.scala 140:38:@38170.4]
  assign _T_117 = _T_116[10:0]; // @[Modules.scala 140:38:@38171.4]
  assign _T_118 = $signed(_T_117); // @[Modules.scala 140:38:@38172.4]
  assign _T_120 = $signed(io_in_1) - $signed(-11'sh2f); // @[Modules.scala 132:28:@38174.4]
  assign _T_121 = _T_120[10:0]; // @[Modules.scala 132:28:@38175.4]
  assign c_x_1 = $signed(_T_121); // @[Modules.scala 132:28:@38176.4]
  assign _GEN_4 = {{15{c_x_1[10]}},c_x_1}; // @[Modules.scala 137:32:@38178.4]
  assign _T_124 = $signed(_GEN_4) << 4'h4; // @[Modules.scala 137:32:@38178.4]
  assign _GEN_5 = _T_124[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_1 = $signed(_GEN_5); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_6 = {{15{x_hat_1[10]}},x_hat_1}; // @[Modules.scala 139:37:@38180.4]
  assign _T_126 = $signed(_GEN_6) << 4'h2; // @[Modules.scala 139:37:@38180.4]
  assign _GEN_7 = _T_126[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_1 = $signed(_GEN_7); // @[Modules.scala 130:28:@38161.4]
  assign _T_128 = $signed(normed_x_hat_1) + $signed(-11'sh5); // @[Modules.scala 140:38:@38182.4]
  assign _T_129 = _T_128[10:0]; // @[Modules.scala 140:38:@38183.4]
  assign _T_130 = $signed(_T_129); // @[Modules.scala 140:38:@38184.4]
  assign _T_132 = $signed(io_in_2) - $signed(11'sh4a); // @[Modules.scala 132:28:@38186.4]
  assign _T_133 = _T_132[10:0]; // @[Modules.scala 132:28:@38187.4]
  assign c_x_2 = $signed(_T_133); // @[Modules.scala 132:28:@38188.4]
  assign _GEN_8 = {{15{c_x_2[10]}},c_x_2}; // @[Modules.scala 137:32:@38190.4]
  assign _T_136 = $signed(_GEN_8) << 4'h4; // @[Modules.scala 137:32:@38190.4]
  assign _GEN_9 = _T_136[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_2 = $signed(_GEN_9); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_10 = {{15{x_hat_2[10]}},x_hat_2}; // @[Modules.scala 139:37:@38192.4]
  assign _T_138 = $signed(_GEN_10) << 4'h2; // @[Modules.scala 139:37:@38192.4]
  assign _GEN_11 = _T_138[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_2 = $signed(_GEN_11); // @[Modules.scala 130:28:@38161.4]
  assign _T_140 = $signed(normed_x_hat_2) + $signed(-11'sh2); // @[Modules.scala 140:38:@38194.4]
  assign _T_141 = _T_140[10:0]; // @[Modules.scala 140:38:@38195.4]
  assign _T_142 = $signed(_T_141); // @[Modules.scala 140:38:@38196.4]
  assign _T_144 = $signed(io_in_3) - $signed(-11'sh90); // @[Modules.scala 132:28:@38198.4]
  assign _T_145 = _T_144[10:0]; // @[Modules.scala 132:28:@38199.4]
  assign c_x_3 = $signed(_T_145); // @[Modules.scala 132:28:@38200.4]
  assign _GEN_12 = {{15{c_x_3[10]}},c_x_3}; // @[Modules.scala 137:32:@38202.4]
  assign _T_148 = $signed(_GEN_12) << 4'h4; // @[Modules.scala 137:32:@38202.4]
  assign _GEN_13 = _T_148[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_3 = $signed(_GEN_13); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_14 = {{15{x_hat_3[10]}},x_hat_3}; // @[Modules.scala 139:37:@38204.4]
  assign _T_150 = $signed(_GEN_14) << 4'h2; // @[Modules.scala 139:37:@38204.4]
  assign _GEN_15 = _T_150[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_3 = $signed(_GEN_15); // @[Modules.scala 130:28:@38161.4]
  assign _T_152 = $signed(normed_x_hat_3) + $signed(11'sh0); // @[Modules.scala 140:38:@38206.4]
  assign _T_153 = _T_152[10:0]; // @[Modules.scala 140:38:@38207.4]
  assign _T_154 = $signed(_T_153); // @[Modules.scala 140:38:@38208.4]
  assign _T_156 = $signed(io_in_4) - $signed(-11'shc); // @[Modules.scala 132:28:@38210.4]
  assign _T_157 = _T_156[10:0]; // @[Modules.scala 132:28:@38211.4]
  assign c_x_4 = $signed(_T_157); // @[Modules.scala 132:28:@38212.4]
  assign _GEN_16 = {{15{c_x_4[10]}},c_x_4}; // @[Modules.scala 137:32:@38214.4]
  assign _T_160 = $signed(_GEN_16) << 4'h4; // @[Modules.scala 137:32:@38214.4]
  assign _GEN_17 = _T_160[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_4 = $signed(_GEN_17); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_18 = {{15{x_hat_4[10]}},x_hat_4}; // @[Modules.scala 139:37:@38216.4]
  assign _T_162 = $signed(_GEN_18) << 4'h2; // @[Modules.scala 139:37:@38216.4]
  assign _GEN_19 = _T_162[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_4 = $signed(_GEN_19); // @[Modules.scala 130:28:@38161.4]
  assign _T_164 = $signed(normed_x_hat_4) + $signed(11'sh11); // @[Modules.scala 140:38:@38218.4]
  assign _T_165 = _T_164[10:0]; // @[Modules.scala 140:38:@38219.4]
  assign _T_166 = $signed(_T_165); // @[Modules.scala 140:38:@38220.4]
  assign _T_168 = $signed(io_in_5) - $signed(11'shc); // @[Modules.scala 132:28:@38222.4]
  assign _T_169 = _T_168[10:0]; // @[Modules.scala 132:28:@38223.4]
  assign c_x_5 = $signed(_T_169); // @[Modules.scala 132:28:@38224.4]
  assign _GEN_20 = {{15{c_x_5[10]}},c_x_5}; // @[Modules.scala 137:32:@38226.4]
  assign _T_172 = $signed(_GEN_20) << 4'h4; // @[Modules.scala 137:32:@38226.4]
  assign _GEN_21 = _T_172[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_5 = $signed(_GEN_21); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_22 = {{15{x_hat_5[10]}},x_hat_5}; // @[Modules.scala 139:37:@38228.4]
  assign _T_174 = $signed(_GEN_22) << 4'h2; // @[Modules.scala 139:37:@38228.4]
  assign _GEN_23 = _T_174[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_5 = $signed(_GEN_23); // @[Modules.scala 130:28:@38161.4]
  assign _T_176 = $signed(normed_x_hat_5) + $signed(11'sh3); // @[Modules.scala 140:38:@38230.4]
  assign _T_177 = _T_176[10:0]; // @[Modules.scala 140:38:@38231.4]
  assign _T_178 = $signed(_T_177); // @[Modules.scala 140:38:@38232.4]
  assign _T_180 = $signed(io_in_6) - $signed(11'sh7d); // @[Modules.scala 132:28:@38234.4]
  assign _T_181 = _T_180[10:0]; // @[Modules.scala 132:28:@38235.4]
  assign c_x_6 = $signed(_T_181); // @[Modules.scala 132:28:@38236.4]
  assign _GEN_24 = {{15{c_x_6[10]}},c_x_6}; // @[Modules.scala 137:32:@38238.4]
  assign _T_184 = $signed(_GEN_24) << 4'h4; // @[Modules.scala 137:32:@38238.4]
  assign _GEN_25 = _T_184[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_6 = $signed(_GEN_25); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_26 = {{15{x_hat_6[10]}},x_hat_6}; // @[Modules.scala 139:37:@38240.4]
  assign _T_186 = $signed(_GEN_26) << 4'h2; // @[Modules.scala 139:37:@38240.4]
  assign _GEN_27 = _T_186[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_6 = $signed(_GEN_27); // @[Modules.scala 130:28:@38161.4]
  assign _T_188 = $signed(normed_x_hat_6) + $signed(-11'sh11); // @[Modules.scala 140:38:@38242.4]
  assign _T_189 = _T_188[10:0]; // @[Modules.scala 140:38:@38243.4]
  assign _T_190 = $signed(_T_189); // @[Modules.scala 140:38:@38244.4]
  assign _T_192 = $signed(io_in_7) - $signed(11'sh3); // @[Modules.scala 132:28:@38246.4]
  assign _T_193 = _T_192[10:0]; // @[Modules.scala 132:28:@38247.4]
  assign c_x_7 = $signed(_T_193); // @[Modules.scala 132:28:@38248.4]
  assign _GEN_28 = {{15{c_x_7[10]}},c_x_7}; // @[Modules.scala 137:32:@38250.4]
  assign _T_196 = $signed(_GEN_28) << 4'h4; // @[Modules.scala 137:32:@38250.4]
  assign _GEN_29 = _T_196[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_7 = $signed(_GEN_29); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_30 = {{15{x_hat_7[10]}},x_hat_7}; // @[Modules.scala 139:37:@38252.4]
  assign _T_198 = $signed(_GEN_30) << 4'h1; // @[Modules.scala 139:37:@38252.4]
  assign _GEN_31 = _T_198[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_7 = $signed(_GEN_31); // @[Modules.scala 130:28:@38161.4]
  assign _T_200 = $signed(normed_x_hat_7) + $signed(11'sh1); // @[Modules.scala 140:38:@38254.4]
  assign _T_201 = _T_200[10:0]; // @[Modules.scala 140:38:@38255.4]
  assign _T_202 = $signed(_T_201); // @[Modules.scala 140:38:@38256.4]
  assign _T_204 = $signed(io_in_8) - $signed(-11'sh5); // @[Modules.scala 132:28:@38258.4]
  assign _T_205 = _T_204[10:0]; // @[Modules.scala 132:28:@38259.4]
  assign c_x_8 = $signed(_T_205); // @[Modules.scala 132:28:@38260.4]
  assign _GEN_32 = {{15{c_x_8[10]}},c_x_8}; // @[Modules.scala 137:32:@38262.4]
  assign _T_208 = $signed(_GEN_32) << 4'h4; // @[Modules.scala 137:32:@38262.4]
  assign _GEN_33 = _T_208[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_8 = $signed(_GEN_33); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_34 = {{15{x_hat_8[10]}},x_hat_8}; // @[Modules.scala 139:37:@38264.4]
  assign _T_210 = $signed(_GEN_34) << 4'h2; // @[Modules.scala 139:37:@38264.4]
  assign _GEN_35 = _T_210[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_8 = $signed(_GEN_35); // @[Modules.scala 130:28:@38161.4]
  assign _T_212 = $signed(normed_x_hat_8) + $signed(-11'sh6); // @[Modules.scala 140:38:@38266.4]
  assign _T_213 = _T_212[10:0]; // @[Modules.scala 140:38:@38267.4]
  assign _T_214 = $signed(_T_213); // @[Modules.scala 140:38:@38268.4]
  assign _T_216 = $signed(io_in_9) - $signed(-11'sh3d); // @[Modules.scala 132:28:@38270.4]
  assign _T_217 = _T_216[10:0]; // @[Modules.scala 132:28:@38271.4]
  assign c_x_9 = $signed(_T_217); // @[Modules.scala 132:28:@38272.4]
  assign _GEN_36 = {{15{c_x_9[10]}},c_x_9}; // @[Modules.scala 137:32:@38274.4]
  assign _T_220 = $signed(_GEN_36) << 4'h4; // @[Modules.scala 137:32:@38274.4]
  assign _GEN_37 = _T_220[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_9 = $signed(_GEN_37); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_38 = {{15{x_hat_9[10]}},x_hat_9}; // @[Modules.scala 139:37:@38276.4]
  assign _T_222 = $signed(_GEN_38) << 4'h1; // @[Modules.scala 139:37:@38276.4]
  assign _GEN_39 = _T_222[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_9 = $signed(_GEN_39); // @[Modules.scala 130:28:@38161.4]
  assign _T_224 = $signed(normed_x_hat_9) + $signed(11'sh1); // @[Modules.scala 140:38:@38278.4]
  assign _T_225 = _T_224[10:0]; // @[Modules.scala 140:38:@38279.4]
  assign _T_226 = $signed(_T_225); // @[Modules.scala 140:38:@38280.4]
  assign _T_228 = $signed(io_in_10) - $signed(-11'shaf); // @[Modules.scala 132:28:@38282.4]
  assign _T_229 = _T_228[10:0]; // @[Modules.scala 132:28:@38283.4]
  assign c_x_10 = $signed(_T_229); // @[Modules.scala 132:28:@38284.4]
  assign _GEN_40 = {{15{c_x_10[10]}},c_x_10}; // @[Modules.scala 137:32:@38286.4]
  assign _T_232 = $signed(_GEN_40) << 4'h4; // @[Modules.scala 137:32:@38286.4]
  assign _GEN_41 = _T_232[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_10 = $signed(_GEN_41); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_42 = {{15{x_hat_10[10]}},x_hat_10}; // @[Modules.scala 139:37:@38288.4]
  assign _T_234 = $signed(_GEN_42) << 4'h2; // @[Modules.scala 139:37:@38288.4]
  assign _GEN_43 = _T_234[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_10 = $signed(_GEN_43); // @[Modules.scala 130:28:@38161.4]
  assign _T_236 = $signed(normed_x_hat_10) + $signed(-11'sh6); // @[Modules.scala 140:38:@38290.4]
  assign _T_237 = _T_236[10:0]; // @[Modules.scala 140:38:@38291.4]
  assign _T_238 = $signed(_T_237); // @[Modules.scala 140:38:@38292.4]
  assign _T_240 = $signed(io_in_11) - $signed(11'sh75); // @[Modules.scala 132:28:@38294.4]
  assign _T_241 = _T_240[10:0]; // @[Modules.scala 132:28:@38295.4]
  assign c_x_11 = $signed(_T_241); // @[Modules.scala 132:28:@38296.4]
  assign _GEN_44 = {{15{c_x_11[10]}},c_x_11}; // @[Modules.scala 137:32:@38298.4]
  assign _T_244 = $signed(_GEN_44) << 4'h4; // @[Modules.scala 137:32:@38298.4]
  assign _GEN_45 = _T_244[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_11 = $signed(_GEN_45); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_46 = {{15{x_hat_11[10]}},x_hat_11}; // @[Modules.scala 139:37:@38300.4]
  assign _T_246 = $signed(_GEN_46) << 4'h1; // @[Modules.scala 139:37:@38300.4]
  assign _GEN_47 = _T_246[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_11 = $signed(_GEN_47); // @[Modules.scala 130:28:@38161.4]
  assign _T_248 = $signed(normed_x_hat_11) + $signed(-11'sh9); // @[Modules.scala 140:38:@38302.4]
  assign _T_249 = _T_248[10:0]; // @[Modules.scala 140:38:@38303.4]
  assign _T_250 = $signed(_T_249); // @[Modules.scala 140:38:@38304.4]
  assign _T_252 = $signed(io_in_12) - $signed(-11'sh32); // @[Modules.scala 132:28:@38306.4]
  assign _T_253 = _T_252[10:0]; // @[Modules.scala 132:28:@38307.4]
  assign c_x_12 = $signed(_T_253); // @[Modules.scala 132:28:@38308.4]
  assign _GEN_48 = {{15{c_x_12[10]}},c_x_12}; // @[Modules.scala 137:32:@38310.4]
  assign _T_256 = $signed(_GEN_48) << 4'h4; // @[Modules.scala 137:32:@38310.4]
  assign _GEN_49 = _T_256[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_12 = $signed(_GEN_49); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_50 = {{15{x_hat_12[10]}},x_hat_12}; // @[Modules.scala 139:37:@38312.4]
  assign _T_258 = $signed(_GEN_50) << 4'h2; // @[Modules.scala 139:37:@38312.4]
  assign _GEN_51 = _T_258[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_12 = $signed(_GEN_51); // @[Modules.scala 130:28:@38161.4]
  assign _T_260 = $signed(normed_x_hat_12) + $signed(-11'sh9); // @[Modules.scala 140:38:@38314.4]
  assign _T_261 = _T_260[10:0]; // @[Modules.scala 140:38:@38315.4]
  assign _T_262 = $signed(_T_261); // @[Modules.scala 140:38:@38316.4]
  assign _T_264 = $signed(io_in_13) - $signed(11'sh77); // @[Modules.scala 132:28:@38318.4]
  assign _T_265 = _T_264[10:0]; // @[Modules.scala 132:28:@38319.4]
  assign c_x_13 = $signed(_T_265); // @[Modules.scala 132:28:@38320.4]
  assign _GEN_52 = {{15{c_x_13[10]}},c_x_13}; // @[Modules.scala 137:32:@38322.4]
  assign _T_268 = $signed(_GEN_52) << 4'h4; // @[Modules.scala 137:32:@38322.4]
  assign _GEN_53 = _T_268[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_13 = $signed(_GEN_53); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_54 = {{15{x_hat_13[10]}},x_hat_13}; // @[Modules.scala 139:37:@38324.4]
  assign _T_270 = $signed(_GEN_54) << 4'h1; // @[Modules.scala 139:37:@38324.4]
  assign _GEN_55 = _T_270[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_13 = $signed(_GEN_55); // @[Modules.scala 130:28:@38161.4]
  assign _T_272 = $signed(normed_x_hat_13) + $signed(11'sh5); // @[Modules.scala 140:38:@38326.4]
  assign _T_273 = _T_272[10:0]; // @[Modules.scala 140:38:@38327.4]
  assign _T_274 = $signed(_T_273); // @[Modules.scala 140:38:@38328.4]
  assign _T_276 = $signed(io_in_14) - $signed(11'sh19); // @[Modules.scala 132:28:@38330.4]
  assign _T_277 = _T_276[10:0]; // @[Modules.scala 132:28:@38331.4]
  assign c_x_14 = $signed(_T_277); // @[Modules.scala 132:28:@38332.4]
  assign _GEN_56 = {{15{c_x_14[10]}},c_x_14}; // @[Modules.scala 137:32:@38334.4]
  assign _T_280 = $signed(_GEN_56) << 4'h4; // @[Modules.scala 137:32:@38334.4]
  assign _GEN_57 = _T_280[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_14 = $signed(_GEN_57); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_58 = {{15{x_hat_14[10]}},x_hat_14}; // @[Modules.scala 139:37:@38336.4]
  assign _T_282 = $signed(_GEN_58) << 4'h2; // @[Modules.scala 139:37:@38336.4]
  assign _GEN_59 = _T_282[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_14 = $signed(_GEN_59); // @[Modules.scala 130:28:@38161.4]
  assign _T_284 = $signed(normed_x_hat_14) + $signed(11'sh7); // @[Modules.scala 140:38:@38338.4]
  assign _T_285 = _T_284[10:0]; // @[Modules.scala 140:38:@38339.4]
  assign _T_286 = $signed(_T_285); // @[Modules.scala 140:38:@38340.4]
  assign _T_288 = $signed(io_in_15) - $signed(-11'sh64); // @[Modules.scala 132:28:@38342.4]
  assign _T_289 = _T_288[10:0]; // @[Modules.scala 132:28:@38343.4]
  assign c_x_15 = $signed(_T_289); // @[Modules.scala 132:28:@38344.4]
  assign _GEN_60 = {{15{c_x_15[10]}},c_x_15}; // @[Modules.scala 137:32:@38346.4]
  assign _T_292 = $signed(_GEN_60) << 4'h4; // @[Modules.scala 137:32:@38346.4]
  assign _GEN_61 = _T_292[10:0]; // @[Modules.scala 129:21:@38160.4]
  assign x_hat_15 = $signed(_GEN_61); // @[Modules.scala 129:21:@38160.4]
  assign _GEN_62 = {{15{x_hat_15[10]}},x_hat_15}; // @[Modules.scala 139:37:@38348.4]
  assign _T_294 = $signed(_GEN_62) << 4'h1; // @[Modules.scala 139:37:@38348.4]
  assign _GEN_63 = _T_294[10:0]; // @[Modules.scala 130:28:@38161.4]
  assign normed_x_hat_15 = $signed(_GEN_63); // @[Modules.scala 130:28:@38161.4]
  assign _T_296 = $signed(normed_x_hat_15) + $signed(11'sh4); // @[Modules.scala 140:38:@38350.4]
  assign _T_297 = _T_296[10:0]; // @[Modules.scala 140:38:@38351.4]
  assign _T_298 = $signed(_T_297); // @[Modules.scala 140:38:@38352.4]
  assign io_out_0 = _T_118;
  assign io_out_1 = _T_130;
  assign io_out_2 = _T_142;
  assign io_out_3 = _T_154;
  assign io_out_4 = _T_166;
  assign io_out_5 = _T_178;
  assign io_out_6 = _T_190;
  assign io_out_7 = _T_202;
  assign io_out_8 = _T_214;
  assign io_out_9 = _T_226;
  assign io_out_10 = _T_238;
  assign io_out_11 = _T_250;
  assign io_out_12 = _T_262;
  assign io_out_13 = _T_274;
  assign io_out_14 = _T_286;
  assign io_out_15 = _T_298;
endmodule
module Binarize( // @[:@38355.2]
  input  [10:0] io_in_0, // @[:@38358.4]
  input  [10:0] io_in_1, // @[:@38358.4]
  input  [10:0] io_in_2, // @[:@38358.4]
  input  [10:0] io_in_3, // @[:@38358.4]
  input  [10:0] io_in_4, // @[:@38358.4]
  input  [10:0] io_in_5, // @[:@38358.4]
  input  [10:0] io_in_6, // @[:@38358.4]
  input  [10:0] io_in_7, // @[:@38358.4]
  input  [10:0] io_in_8, // @[:@38358.4]
  input  [10:0] io_in_9, // @[:@38358.4]
  input  [10:0] io_in_10, // @[:@38358.4]
  input  [10:0] io_in_11, // @[:@38358.4]
  input  [10:0] io_in_12, // @[:@38358.4]
  input  [10:0] io_in_13, // @[:@38358.4]
  input  [10:0] io_in_14, // @[:@38358.4]
  input  [10:0] io_in_15, // @[:@38358.4]
  output [1:0]  io_out_0, // @[:@38358.4]
  output [1:0]  io_out_1, // @[:@38358.4]
  output [1:0]  io_out_2, // @[:@38358.4]
  output [1:0]  io_out_3, // @[:@38358.4]
  output [1:0]  io_out_4, // @[:@38358.4]
  output [1:0]  io_out_5, // @[:@38358.4]
  output [1:0]  io_out_6, // @[:@38358.4]
  output [1:0]  io_out_7, // @[:@38358.4]
  output [1:0]  io_out_8, // @[:@38358.4]
  output [1:0]  io_out_9, // @[:@38358.4]
  output [1:0]  io_out_10, // @[:@38358.4]
  output [1:0]  io_out_11, // @[:@38358.4]
  output [1:0]  io_out_12, // @[:@38358.4]
  output [1:0]  io_out_13, // @[:@38358.4]
  output [1:0]  io_out_14, // @[:@38358.4]
  output [1:0]  io_out_15 // @[:@38358.4]
);
  wire  _T_45; // @[Modules.scala 151:24:@38360.4]
  wire [1:0] _GEN_0; // @[Modules.scala 151:32:@38361.4]
  wire  _T_49; // @[Modules.scala 151:24:@38367.4]
  wire [1:0] _GEN_1; // @[Modules.scala 151:32:@38368.4]
  wire  _T_53; // @[Modules.scala 151:24:@38374.4]
  wire [1:0] _GEN_2; // @[Modules.scala 151:32:@38375.4]
  wire  _T_57; // @[Modules.scala 151:24:@38381.4]
  wire [1:0] _GEN_3; // @[Modules.scala 151:32:@38382.4]
  wire  _T_61; // @[Modules.scala 151:24:@38388.4]
  wire [1:0] _GEN_4; // @[Modules.scala 151:32:@38389.4]
  wire  _T_65; // @[Modules.scala 151:24:@38395.4]
  wire [1:0] _GEN_5; // @[Modules.scala 151:32:@38396.4]
  wire  _T_69; // @[Modules.scala 151:24:@38402.4]
  wire [1:0] _GEN_6; // @[Modules.scala 151:32:@38403.4]
  wire  _T_73; // @[Modules.scala 151:24:@38409.4]
  wire [1:0] _GEN_7; // @[Modules.scala 151:32:@38410.4]
  wire  _T_77; // @[Modules.scala 151:24:@38416.4]
  wire [1:0] _GEN_8; // @[Modules.scala 151:32:@38417.4]
  wire  _T_81; // @[Modules.scala 151:24:@38423.4]
  wire [1:0] _GEN_9; // @[Modules.scala 151:32:@38424.4]
  wire  _T_85; // @[Modules.scala 151:24:@38430.4]
  wire [1:0] _GEN_10; // @[Modules.scala 151:32:@38431.4]
  wire  _T_89; // @[Modules.scala 151:24:@38437.4]
  wire [1:0] _GEN_11; // @[Modules.scala 151:32:@38438.4]
  wire  _T_93; // @[Modules.scala 151:24:@38444.4]
  wire [1:0] _GEN_12; // @[Modules.scala 151:32:@38445.4]
  wire  _T_97; // @[Modules.scala 151:24:@38451.4]
  wire [1:0] _GEN_13; // @[Modules.scala 151:32:@38452.4]
  wire  _T_101; // @[Modules.scala 151:24:@38458.4]
  wire [1:0] _GEN_14; // @[Modules.scala 151:32:@38459.4]
  wire  _T_105; // @[Modules.scala 151:24:@38465.4]
  wire [1:0] _GEN_15; // @[Modules.scala 151:32:@38466.4]
  assign _T_45 = $signed(io_in_0) >= $signed(11'sh0); // @[Modules.scala 151:24:@38360.4]
  assign _GEN_0 = _T_45 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38361.4]
  assign _T_49 = $signed(io_in_1) >= $signed(11'sh0); // @[Modules.scala 151:24:@38367.4]
  assign _GEN_1 = _T_49 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38368.4]
  assign _T_53 = $signed(io_in_2) >= $signed(11'sh0); // @[Modules.scala 151:24:@38374.4]
  assign _GEN_2 = _T_53 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38375.4]
  assign _T_57 = $signed(io_in_3) >= $signed(11'sh0); // @[Modules.scala 151:24:@38381.4]
  assign _GEN_3 = _T_57 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38382.4]
  assign _T_61 = $signed(io_in_4) >= $signed(11'sh0); // @[Modules.scala 151:24:@38388.4]
  assign _GEN_4 = _T_61 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38389.4]
  assign _T_65 = $signed(io_in_5) >= $signed(11'sh0); // @[Modules.scala 151:24:@38395.4]
  assign _GEN_5 = _T_65 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38396.4]
  assign _T_69 = $signed(io_in_6) >= $signed(11'sh0); // @[Modules.scala 151:24:@38402.4]
  assign _GEN_6 = _T_69 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38403.4]
  assign _T_73 = $signed(io_in_7) >= $signed(11'sh0); // @[Modules.scala 151:24:@38409.4]
  assign _GEN_7 = _T_73 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38410.4]
  assign _T_77 = $signed(io_in_8) >= $signed(11'sh0); // @[Modules.scala 151:24:@38416.4]
  assign _GEN_8 = _T_77 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38417.4]
  assign _T_81 = $signed(io_in_9) >= $signed(11'sh0); // @[Modules.scala 151:24:@38423.4]
  assign _GEN_9 = _T_81 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38424.4]
  assign _T_85 = $signed(io_in_10) >= $signed(11'sh0); // @[Modules.scala 151:24:@38430.4]
  assign _GEN_10 = _T_85 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38431.4]
  assign _T_89 = $signed(io_in_11) >= $signed(11'sh0); // @[Modules.scala 151:24:@38437.4]
  assign _GEN_11 = _T_89 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38438.4]
  assign _T_93 = $signed(io_in_12) >= $signed(11'sh0); // @[Modules.scala 151:24:@38444.4]
  assign _GEN_12 = _T_93 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38445.4]
  assign _T_97 = $signed(io_in_13) >= $signed(11'sh0); // @[Modules.scala 151:24:@38451.4]
  assign _GEN_13 = _T_97 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38452.4]
  assign _T_101 = $signed(io_in_14) >= $signed(11'sh0); // @[Modules.scala 151:24:@38458.4]
  assign _GEN_14 = _T_101 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38459.4]
  assign _T_105 = $signed(io_in_15) >= $signed(11'sh0); // @[Modules.scala 151:24:@38465.4]
  assign _GEN_15 = _T_105 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@38466.4]
  assign io_out_0 = _GEN_0;
  assign io_out_1 = _GEN_1;
  assign io_out_2 = _GEN_2;
  assign io_out_3 = _GEN_3;
  assign io_out_4 = _GEN_4;
  assign io_out_5 = _GEN_5;
  assign io_out_6 = _GEN_6;
  assign io_out_7 = _GEN_7;
  assign io_out_8 = _GEN_8;
  assign io_out_9 = _GEN_9;
  assign io_out_10 = _GEN_10;
  assign io_out_11 = _GEN_11;
  assign io_out_12 = _GEN_12;
  assign io_out_13 = _GEN_13;
  assign io_out_14 = _GEN_14;
  assign io_out_15 = _GEN_15;
endmodule
module Linear( // @[:@38473.2]
  input  [1:0] io_in_0, // @[:@38476.4]
  input  [1:0] io_in_1, // @[:@38476.4]
  input  [1:0] io_in_2, // @[:@38476.4]
  input  [1:0] io_in_3, // @[:@38476.4]
  input  [1:0] io_in_4, // @[:@38476.4]
  input  [1:0] io_in_5, // @[:@38476.4]
  input  [1:0] io_in_6, // @[:@38476.4]
  input  [1:0] io_in_7, // @[:@38476.4]
  input  [1:0] io_in_8, // @[:@38476.4]
  input  [1:0] io_in_9, // @[:@38476.4]
  input  [1:0] io_in_10, // @[:@38476.4]
  input  [1:0] io_in_11, // @[:@38476.4]
  input  [1:0] io_in_12, // @[:@38476.4]
  input  [1:0] io_in_13, // @[:@38476.4]
  input  [1:0] io_in_14, // @[:@38476.4]
  input  [1:0] io_in_15, // @[:@38476.4]
  output [7:0] io_out_0, // @[:@38476.4]
  output [7:0] io_out_1, // @[:@38476.4]
  output [7:0] io_out_2, // @[:@38476.4]
  output [7:0] io_out_3, // @[:@38476.4]
  output [7:0] io_out_4, // @[:@38476.4]
  output [7:0] io_out_5, // @[:@38476.4]
  output [7:0] io_out_6, // @[:@38476.4]
  output [7:0] io_out_7, // @[:@38476.4]
  output [7:0] io_out_8, // @[:@38476.4]
  output [7:0] io_out_9, // @[:@38476.4]
  output [7:0] io_out_10, // @[:@38476.4]
  output [7:0] io_out_11, // @[:@38476.4]
  output [7:0] io_out_12, // @[:@38476.4]
  output [7:0] io_out_13, // @[:@38476.4]
  output [7:0] io_out_14, // @[:@38476.4]
  output [7:0] io_out_15 // @[:@38476.4]
);
  wire [7:0] _GEN_0; // @[Modules.scala 108:54:@38481.4]
  wire [8:0] _T_1275; // @[Modules.scala 108:54:@38481.4]
  wire [7:0] _T_1276; // @[Modules.scala 108:54:@38482.4]
  wire [7:0] buffer_0_2; // @[Modules.scala 108:54:@38483.4]
  wire [7:0] _GEN_1; // @[Modules.scala 108:54:@38487.4]
  wire [8:0] _T_1278; // @[Modules.scala 108:54:@38487.4]
  wire [7:0] _T_1279; // @[Modules.scala 108:54:@38488.4]
  wire [7:0] buffer_0_5; // @[Modules.scala 108:54:@38489.4]
  wire [7:0] _GEN_2; // @[Modules.scala 108:54:@38491.4]
  wire [8:0] _T_1281; // @[Modules.scala 108:54:@38491.4]
  wire [7:0] _T_1282; // @[Modules.scala 108:54:@38492.4]
  wire [7:0] buffer_0_6; // @[Modules.scala 108:54:@38493.4]
  wire [7:0] _GEN_3; // @[Modules.scala 108:54:@38495.4]
  wire [8:0] _T_1284; // @[Modules.scala 108:54:@38495.4]
  wire [7:0] _T_1285; // @[Modules.scala 108:54:@38496.4]
  wire [7:0] buffer_0_7; // @[Modules.scala 108:54:@38497.4]
  wire [7:0] _GEN_4; // @[Modules.scala 108:54:@38502.4]
  wire [8:0] _T_1287; // @[Modules.scala 108:54:@38502.4]
  wire [7:0] _T_1288; // @[Modules.scala 108:54:@38503.4]
  wire [7:0] buffer_0_11; // @[Modules.scala 108:54:@38504.4]
  wire [7:0] buffer_1_0; // @[Modules.scala 91:22:@38478.4]
  wire [7:0] _GEN_5; // @[Modules.scala 108:54:@38512.4]
  wire [8:0] _T_1290; // @[Modules.scala 108:54:@38512.4]
  wire [7:0] _T_1291; // @[Modules.scala 108:54:@38513.4]
  wire [7:0] buffer_1_1; // @[Modules.scala 108:54:@38514.4]
  wire [8:0] _T_1293; // @[Modules.scala 108:54:@38516.4]
  wire [7:0] _T_1294; // @[Modules.scala 108:54:@38517.4]
  wire [7:0] buffer_1_2; // @[Modules.scala 108:54:@38518.4]
  wire [7:0] _GEN_7; // @[Modules.scala 108:54:@38521.4]
  wire [8:0] _T_1296; // @[Modules.scala 108:54:@38521.4]
  wire [7:0] _T_1297; // @[Modules.scala 108:54:@38522.4]
  wire [7:0] buffer_1_4; // @[Modules.scala 108:54:@38523.4]
  wire [8:0] _T_1299; // @[Modules.scala 108:54:@38526.4]
  wire [7:0] _T_1300; // @[Modules.scala 108:54:@38527.4]
  wire [7:0] buffer_1_6; // @[Modules.scala 108:54:@38528.4]
  wire [7:0] _GEN_9; // @[Modules.scala 108:54:@38535.4]
  wire [8:0] _T_1302; // @[Modules.scala 108:54:@38535.4]
  wire [7:0] _T_1303; // @[Modules.scala 108:54:@38536.4]
  wire [7:0] buffer_1_12; // @[Modules.scala 108:54:@38537.4]
  wire [7:0] _GEN_10; // @[Modules.scala 108:54:@38539.4]
  wire [8:0] _T_1305; // @[Modules.scala 108:54:@38539.4]
  wire [7:0] _T_1306; // @[Modules.scala 108:54:@38540.4]
  wire [7:0] buffer_1_13; // @[Modules.scala 108:54:@38541.4]
  wire [7:0] _GEN_11; // @[Modules.scala 108:54:@38544.4]
  wire [8:0] _T_1308; // @[Modules.scala 108:54:@38544.4]
  wire [7:0] _T_1309; // @[Modules.scala 108:54:@38545.4]
  wire [7:0] buffer_1_15; // @[Modules.scala 108:54:@38546.4]
  wire [8:0] _T_1311; // @[Modules.scala 108:54:@38551.4]
  wire [7:0] _T_1312; // @[Modules.scala 108:54:@38552.4]
  wire [7:0] buffer_2_2; // @[Modules.scala 108:54:@38553.4]
  wire [8:0] _T_1314; // @[Modules.scala 108:54:@38556.4]
  wire [7:0] _T_1315; // @[Modules.scala 108:54:@38557.4]
  wire [7:0] buffer_2_4; // @[Modules.scala 108:54:@38558.4]
  wire [8:0] _T_1317; // @[Modules.scala 108:54:@38562.4]
  wire [7:0] _T_1318; // @[Modules.scala 108:54:@38563.4]
  wire [7:0] buffer_2_7; // @[Modules.scala 108:54:@38564.4]
  wire [7:0] _GEN_15; // @[Modules.scala 108:54:@38566.4]
  wire [8:0] _T_1320; // @[Modules.scala 108:54:@38566.4]
  wire [7:0] _T_1321; // @[Modules.scala 108:54:@38567.4]
  wire [7:0] buffer_2_8; // @[Modules.scala 108:54:@38568.4]
  wire [7:0] _GEN_16; // @[Modules.scala 108:54:@38570.4]
  wire [8:0] _T_1323; // @[Modules.scala 108:54:@38570.4]
  wire [7:0] _T_1324; // @[Modules.scala 108:54:@38571.4]
  wire [7:0] buffer_2_9; // @[Modules.scala 108:54:@38572.4]
  wire [7:0] _GEN_17; // @[Modules.scala 108:54:@38574.4]
  wire [8:0] _T_1326; // @[Modules.scala 108:54:@38574.4]
  wire [7:0] _T_1327; // @[Modules.scala 108:54:@38575.4]
  wire [7:0] buffer_2_10; // @[Modules.scala 108:54:@38576.4]
  wire [8:0] _T_1329; // @[Modules.scala 108:54:@38578.4]
  wire [7:0] _T_1330; // @[Modules.scala 108:54:@38579.4]
  wire [7:0] buffer_2_11; // @[Modules.scala 108:54:@38580.4]
  wire [8:0] _T_1332; // @[Modules.scala 108:54:@38582.4]
  wire [7:0] _T_1333; // @[Modules.scala 108:54:@38583.4]
  wire [7:0] buffer_2_12; // @[Modules.scala 108:54:@38584.4]
  wire [8:0] _T_1335; // @[Modules.scala 108:54:@38586.4]
  wire [7:0] _T_1336; // @[Modules.scala 108:54:@38587.4]
  wire [7:0] buffer_2_13; // @[Modules.scala 108:54:@38588.4]
  wire [8:0] _T_1338; // @[Modules.scala 108:54:@38591.4]
  wire [7:0] _T_1339; // @[Modules.scala 108:54:@38592.4]
  wire [7:0] buffer_2_15; // @[Modules.scala 108:54:@38593.4]
  wire [7:0] _GEN_22; // @[Modules.scala 108:54:@38599.4]
  wire [8:0] _T_1342; // @[Modules.scala 108:54:@38599.4]
  wire [7:0] _T_1343; // @[Modules.scala 108:54:@38600.4]
  wire [7:0] buffer_3_3; // @[Modules.scala 108:54:@38601.4]
  wire [8:0] _T_1345; // @[Modules.scala 108:54:@38604.4]
  wire [7:0] _T_1346; // @[Modules.scala 108:54:@38605.4]
  wire [7:0] buffer_3_5; // @[Modules.scala 108:54:@38606.4]
  wire [8:0] _T_1348; // @[Modules.scala 108:54:@38609.4]
  wire [7:0] _T_1349; // @[Modules.scala 108:54:@38610.4]
  wire [7:0] buffer_3_7; // @[Modules.scala 108:54:@38611.4]
  wire [8:0] _T_1351; // @[Modules.scala 108:54:@38613.4]
  wire [7:0] _T_1352; // @[Modules.scala 108:54:@38614.4]
  wire [7:0] buffer_3_8; // @[Modules.scala 108:54:@38615.4]
  wire [8:0] _T_1354; // @[Modules.scala 108:54:@38617.4]
  wire [7:0] _T_1355; // @[Modules.scala 108:54:@38618.4]
  wire [7:0] buffer_3_9; // @[Modules.scala 108:54:@38619.4]
  wire [8:0] _T_1357; // @[Modules.scala 108:54:@38621.4]
  wire [7:0] _T_1358; // @[Modules.scala 108:54:@38622.4]
  wire [7:0] buffer_3_10; // @[Modules.scala 108:54:@38623.4]
  wire [8:0] _T_1360; // @[Modules.scala 108:54:@38626.4]
  wire [7:0] _T_1361; // @[Modules.scala 108:54:@38627.4]
  wire [7:0] buffer_3_12; // @[Modules.scala 108:54:@38628.4]
  wire [8:0] _T_1363; // @[Modules.scala 108:54:@38632.4]
  wire [7:0] _T_1364; // @[Modules.scala 108:54:@38633.4]
  wire [7:0] buffer_3_15; // @[Modules.scala 108:54:@38634.4]
  wire [8:0] _T_1378; // @[Modules.scala 108:54:@38656.4]
  wire [7:0] _T_1379; // @[Modules.scala 108:54:@38657.4]
  wire [7:0] buffer_4_7; // @[Modules.scala 108:54:@38658.4]
  wire [8:0] _T_1381; // @[Modules.scala 108:54:@38660.4]
  wire [7:0] _T_1382; // @[Modules.scala 108:54:@38661.4]
  wire [7:0] buffer_4_8; // @[Modules.scala 108:54:@38662.4]
  wire [8:0] _T_1384; // @[Modules.scala 108:54:@38665.4]
  wire [7:0] _T_1385; // @[Modules.scala 108:54:@38666.4]
  wire [7:0] buffer_4_10; // @[Modules.scala 108:54:@38667.4]
  wire [8:0] _T_1387; // @[Modules.scala 108:54:@38669.4]
  wire [7:0] _T_1388; // @[Modules.scala 108:54:@38670.4]
  wire [7:0] buffer_4_11; // @[Modules.scala 108:54:@38671.4]
  wire [8:0] _T_1391; // @[Modules.scala 108:54:@38679.4]
  wire [7:0] _T_1392; // @[Modules.scala 108:54:@38680.4]
  wire [7:0] buffer_5_1; // @[Modules.scala 108:54:@38681.4]
  wire [8:0] _T_1394; // @[Modules.scala 108:54:@38683.4]
  wire [7:0] _T_1395; // @[Modules.scala 108:54:@38684.4]
  wire [7:0] buffer_5_2; // @[Modules.scala 108:54:@38685.4]
  wire [8:0] _T_1397; // @[Modules.scala 108:54:@38688.4]
  wire [7:0] _T_1398; // @[Modules.scala 108:54:@38689.4]
  wire [7:0] buffer_5_4; // @[Modules.scala 108:54:@38690.4]
  wire [8:0] _T_1400; // @[Modules.scala 108:54:@38694.4]
  wire [7:0] _T_1401; // @[Modules.scala 108:54:@38695.4]
  wire [7:0] buffer_5_7; // @[Modules.scala 108:54:@38696.4]
  wire [8:0] _T_1403; // @[Modules.scala 108:54:@38699.4]
  wire [7:0] _T_1404; // @[Modules.scala 108:54:@38700.4]
  wire [7:0] buffer_5_9; // @[Modules.scala 108:54:@38701.4]
  wire [8:0] _T_1406; // @[Modules.scala 108:54:@38703.4]
  wire [7:0] _T_1407; // @[Modules.scala 108:54:@38704.4]
  wire [7:0] buffer_5_10; // @[Modules.scala 108:54:@38705.4]
  wire [8:0] _T_1409; // @[Modules.scala 108:54:@38707.4]
  wire [7:0] _T_1410; // @[Modules.scala 108:54:@38708.4]
  wire [7:0] buffer_5_11; // @[Modules.scala 108:54:@38709.4]
  wire [8:0] _T_1415; // @[Modules.scala 108:54:@38724.4]
  wire [7:0] _T_1416; // @[Modules.scala 108:54:@38725.4]
  wire [7:0] buffer_6_5; // @[Modules.scala 108:54:@38726.4]
  wire [8:0] _T_1418; // @[Modules.scala 108:54:@38729.4]
  wire [7:0] _T_1419; // @[Modules.scala 108:54:@38730.4]
  wire [7:0] buffer_6_7; // @[Modules.scala 108:54:@38731.4]
  wire [8:0] _T_1421; // @[Modules.scala 108:54:@38733.4]
  wire [7:0] _T_1422; // @[Modules.scala 108:54:@38734.4]
  wire [7:0] buffer_6_8; // @[Modules.scala 108:54:@38735.4]
  wire [8:0] _T_1424; // @[Modules.scala 108:54:@38739.4]
  wire [7:0] _T_1425; // @[Modules.scala 108:54:@38740.4]
  wire [7:0] buffer_6_11; // @[Modules.scala 108:54:@38741.4]
  wire [8:0] _T_1427; // @[Modules.scala 108:54:@38744.4]
  wire [7:0] _T_1428; // @[Modules.scala 108:54:@38745.4]
  wire [7:0] buffer_6_13; // @[Modules.scala 108:54:@38746.4]
  wire [7:0] _GEN_51; // @[Modules.scala 108:54:@38748.4]
  wire [8:0] _T_1430; // @[Modules.scala 108:54:@38748.4]
  wire [7:0] _T_1431; // @[Modules.scala 108:54:@38749.4]
  wire [7:0] buffer_6_14; // @[Modules.scala 108:54:@38750.4]
  wire [8:0] _T_1433; // @[Modules.scala 108:54:@38757.4]
  wire [7:0] _T_1434; // @[Modules.scala 108:54:@38758.4]
  wire [7:0] buffer_7_3; // @[Modules.scala 108:54:@38759.4]
  wire [8:0] _T_1436; // @[Modules.scala 108:54:@38762.4]
  wire [7:0] _T_1437; // @[Modules.scala 108:54:@38763.4]
  wire [7:0] buffer_7_5; // @[Modules.scala 108:54:@38764.4]
  wire [8:0] _T_1439; // @[Modules.scala 108:54:@38766.4]
  wire [7:0] _T_1440; // @[Modules.scala 108:54:@38767.4]
  wire [7:0] buffer_7_6; // @[Modules.scala 108:54:@38768.4]
  wire [8:0] _T_1442; // @[Modules.scala 108:54:@38771.4]
  wire [7:0] _T_1443; // @[Modules.scala 108:54:@38772.4]
  wire [7:0] buffer_7_8; // @[Modules.scala 108:54:@38773.4]
  wire [8:0] _T_1445; // @[Modules.scala 108:54:@38775.4]
  wire [7:0] _T_1446; // @[Modules.scala 108:54:@38776.4]
  wire [7:0] buffer_7_9; // @[Modules.scala 108:54:@38777.4]
  wire [8:0] _T_1448; // @[Modules.scala 108:54:@38779.4]
  wire [7:0] _T_1449; // @[Modules.scala 108:54:@38780.4]
  wire [7:0] buffer_7_10; // @[Modules.scala 108:54:@38781.4]
  wire [8:0] _T_1451; // @[Modules.scala 108:54:@38787.4]
  wire [7:0] _T_1452; // @[Modules.scala 108:54:@38788.4]
  wire [7:0] buffer_7_15; // @[Modules.scala 108:54:@38789.4]
  wire [8:0] _T_1460; // @[Modules.scala 108:54:@38804.4]
  wire [7:0] _T_1461; // @[Modules.scala 108:54:@38805.4]
  wire [7:0] buffer_8_6; // @[Modules.scala 108:54:@38806.4]
  wire [8:0] _T_1463; // @[Modules.scala 108:54:@38808.4]
  wire [7:0] _T_1464; // @[Modules.scala 108:54:@38809.4]
  wire [7:0] buffer_8_7; // @[Modules.scala 108:54:@38810.4]
  wire [8:0] _T_1466; // @[Modules.scala 108:54:@38812.4]
  wire [7:0] _T_1467; // @[Modules.scala 108:54:@38813.4]
  wire [7:0] buffer_8_8; // @[Modules.scala 108:54:@38814.4]
  wire [8:0] _T_1469; // @[Modules.scala 108:54:@38817.4]
  wire [7:0] _T_1470; // @[Modules.scala 108:54:@38818.4]
  wire [7:0] buffer_8_10; // @[Modules.scala 108:54:@38819.4]
  wire [8:0] _T_1472; // @[Modules.scala 108:54:@38822.4]
  wire [7:0] _T_1473; // @[Modules.scala 108:54:@38823.4]
  wire [7:0] buffer_8_12; // @[Modules.scala 108:54:@38824.4]
  wire [8:0] _T_1475; // @[Modules.scala 108:54:@38826.4]
  wire [7:0] _T_1476; // @[Modules.scala 108:54:@38827.4]
  wire [7:0] buffer_8_13; // @[Modules.scala 108:54:@38828.4]
  wire [8:0] _T_1478; // @[Modules.scala 108:54:@38831.4]
  wire [7:0] _T_1479; // @[Modules.scala 108:54:@38832.4]
  wire [7:0] buffer_8_15; // @[Modules.scala 108:54:@38833.4]
  wire [8:0] _T_1487; // @[Modules.scala 108:54:@38845.4]
  wire [7:0] _T_1488; // @[Modules.scala 108:54:@38846.4]
  wire [7:0] buffer_9_3; // @[Modules.scala 108:54:@38847.4]
  wire [8:0] _T_1490; // @[Modules.scala 108:54:@38849.4]
  wire [7:0] _T_1491; // @[Modules.scala 108:54:@38850.4]
  wire [7:0] buffer_9_4; // @[Modules.scala 108:54:@38851.4]
  wire [8:0] _T_1493; // @[Modules.scala 108:54:@38854.4]
  wire [7:0] _T_1494; // @[Modules.scala 108:54:@38855.4]
  wire [7:0] buffer_9_6; // @[Modules.scala 108:54:@38856.4]
  wire [8:0] _T_1496; // @[Modules.scala 108:54:@38859.4]
  wire [7:0] _T_1497; // @[Modules.scala 108:54:@38860.4]
  wire [7:0] buffer_9_8; // @[Modules.scala 108:54:@38861.4]
  wire [8:0] _T_1499; // @[Modules.scala 108:54:@38868.4]
  wire [7:0] _T_1500; // @[Modules.scala 108:54:@38869.4]
  wire [7:0] buffer_9_14; // @[Modules.scala 108:54:@38870.4]
  wire [8:0] _T_1509; // @[Modules.scala 108:54:@38883.4]
  wire [7:0] _T_1510; // @[Modules.scala 108:54:@38884.4]
  wire [7:0] buffer_10_3; // @[Modules.scala 108:54:@38885.4]
  wire [8:0] _T_1512; // @[Modules.scala 108:54:@38893.4]
  wire [7:0] _T_1513; // @[Modules.scala 108:54:@38894.4]
  wire [7:0] buffer_10_10; // @[Modules.scala 108:54:@38895.4]
  wire [8:0] _T_1515; // @[Modules.scala 108:54:@38897.4]
  wire [7:0] _T_1516; // @[Modules.scala 108:54:@38898.4]
  wire [7:0] buffer_10_11; // @[Modules.scala 108:54:@38899.4]
  wire [8:0] _T_1518; // @[Modules.scala 108:54:@38901.4]
  wire [7:0] _T_1519; // @[Modules.scala 108:54:@38902.4]
  wire [7:0] buffer_10_12; // @[Modules.scala 108:54:@38903.4]
  wire [8:0] _T_1521; // @[Modules.scala 108:54:@38907.4]
  wire [7:0] _T_1522; // @[Modules.scala 108:54:@38908.4]
  wire [7:0] buffer_10_15; // @[Modules.scala 108:54:@38909.4]
  wire [8:0] _T_1528; // @[Modules.scala 108:54:@38919.4]
  wire [7:0] _T_1529; // @[Modules.scala 108:54:@38920.4]
  wire [7:0] buffer_11_4; // @[Modules.scala 108:54:@38921.4]
  wire [8:0] _T_1531; // @[Modules.scala 108:54:@38924.4]
  wire [7:0] _T_1532; // @[Modules.scala 108:54:@38925.4]
  wire [7:0] buffer_11_6; // @[Modules.scala 108:54:@38926.4]
  wire [8:0] _T_1534; // @[Modules.scala 108:54:@38929.4]
  wire [7:0] _T_1535; // @[Modules.scala 108:54:@38930.4]
  wire [7:0] buffer_11_8; // @[Modules.scala 108:54:@38931.4]
  wire [8:0] _T_1537; // @[Modules.scala 108:54:@38936.4]
  wire [7:0] _T_1538; // @[Modules.scala 108:54:@38937.4]
  wire [7:0] buffer_11_12; // @[Modules.scala 108:54:@38938.4]
  wire [8:0] _T_1540; // @[Modules.scala 108:54:@38940.4]
  wire [7:0] _T_1541; // @[Modules.scala 108:54:@38941.4]
  wire [7:0] buffer_11_13; // @[Modules.scala 108:54:@38942.4]
  wire [8:0] _T_1543; // @[Modules.scala 108:54:@38945.4]
  wire [7:0] _T_1544; // @[Modules.scala 108:54:@38946.4]
  wire [7:0] buffer_11_15; // @[Modules.scala 108:54:@38947.4]
  wire [8:0] _T_1549; // @[Modules.scala 108:54:@38956.4]
  wire [7:0] _T_1550; // @[Modules.scala 108:54:@38957.4]
  wire [7:0] buffer_12_3; // @[Modules.scala 108:54:@38958.4]
  wire [8:0] _T_1552; // @[Modules.scala 108:54:@38960.4]
  wire [7:0] _T_1553; // @[Modules.scala 108:54:@38961.4]
  wire [7:0] buffer_12_4; // @[Modules.scala 108:54:@38962.4]
  wire [8:0] _T_1555; // @[Modules.scala 108:54:@38966.4]
  wire [7:0] _T_1556; // @[Modules.scala 108:54:@38967.4]
  wire [7:0] buffer_12_7; // @[Modules.scala 108:54:@38968.4]
  wire [8:0] _T_1558; // @[Modules.scala 108:54:@38971.4]
  wire [7:0] _T_1559; // @[Modules.scala 108:54:@38972.4]
  wire [7:0] buffer_12_9; // @[Modules.scala 108:54:@38973.4]
  wire [8:0] _T_1561; // @[Modules.scala 108:54:@38975.4]
  wire [7:0] _T_1562; // @[Modules.scala 108:54:@38976.4]
  wire [7:0] buffer_12_10; // @[Modules.scala 108:54:@38977.4]
  wire [8:0] _T_1564; // @[Modules.scala 108:54:@38980.4]
  wire [7:0] _T_1565; // @[Modules.scala 108:54:@38981.4]
  wire [7:0] buffer_12_12; // @[Modules.scala 108:54:@38982.4]
  wire [8:0] _T_1567; // @[Modules.scala 108:54:@38984.4]
  wire [7:0] _T_1568; // @[Modules.scala 108:54:@38985.4]
  wire [7:0] buffer_12_13; // @[Modules.scala 108:54:@38986.4]
  wire [8:0] _T_1570; // @[Modules.scala 108:54:@38988.4]
  wire [7:0] _T_1571; // @[Modules.scala 108:54:@38989.4]
  wire [7:0] buffer_12_14; // @[Modules.scala 108:54:@38990.4]
  wire [8:0] _T_1573; // @[Modules.scala 108:54:@38992.4]
  wire [7:0] _T_1574; // @[Modules.scala 108:54:@38993.4]
  wire [7:0] buffer_12_15; // @[Modules.scala 108:54:@38994.4]
  wire [8:0] _T_1588; // @[Modules.scala 108:54:@39016.4]
  wire [7:0] _T_1589; // @[Modules.scala 108:54:@39017.4]
  wire [7:0] buffer_13_7; // @[Modules.scala 108:54:@39018.4]
  wire [8:0] _T_1591; // @[Modules.scala 108:54:@39020.4]
  wire [7:0] _T_1592; // @[Modules.scala 108:54:@39021.4]
  wire [7:0] buffer_13_8; // @[Modules.scala 108:54:@39022.4]
  wire [8:0] _T_1594; // @[Modules.scala 108:54:@39026.4]
  wire [7:0] _T_1595; // @[Modules.scala 108:54:@39027.4]
  wire [7:0] buffer_13_11; // @[Modules.scala 108:54:@39028.4]
  wire [8:0] _T_1597; // @[Modules.scala 108:54:@39030.4]
  wire [7:0] _T_1598; // @[Modules.scala 108:54:@39031.4]
  wire [7:0] buffer_13_12; // @[Modules.scala 108:54:@39032.4]
  wire [8:0] _T_1600; // @[Modules.scala 108:54:@39034.4]
  wire [7:0] _T_1601; // @[Modules.scala 108:54:@39035.4]
  wire [7:0] buffer_13_13; // @[Modules.scala 108:54:@39036.4]
  wire [8:0] _T_1603; // @[Modules.scala 108:54:@39039.4]
  wire [7:0] _T_1604; // @[Modules.scala 108:54:@39040.4]
  wire [7:0] buffer_13_15; // @[Modules.scala 108:54:@39041.4]
  wire [8:0] _T_1612; // @[Modules.scala 108:54:@39055.4]
  wire [7:0] _T_1613; // @[Modules.scala 108:54:@39056.4]
  wire [7:0] buffer_14_5; // @[Modules.scala 108:54:@39057.4]
  wire [8:0] _T_1615; // @[Modules.scala 108:54:@39059.4]
  wire [7:0] _T_1616; // @[Modules.scala 108:54:@39060.4]
  wire [7:0] buffer_14_6; // @[Modules.scala 108:54:@39061.4]
  wire [8:0] _T_1618; // @[Modules.scala 108:54:@39063.4]
  wire [7:0] _T_1619; // @[Modules.scala 108:54:@39064.4]
  wire [7:0] buffer_14_7; // @[Modules.scala 108:54:@39065.4]
  wire [8:0] _T_1621; // @[Modules.scala 108:54:@39068.4]
  wire [7:0] _T_1622; // @[Modules.scala 108:54:@39069.4]
  wire [7:0] buffer_14_9; // @[Modules.scala 108:54:@39070.4]
  wire [8:0] _T_1624; // @[Modules.scala 108:54:@39074.4]
  wire [7:0] _T_1625; // @[Modules.scala 108:54:@39075.4]
  wire [7:0] buffer_14_12; // @[Modules.scala 108:54:@39076.4]
  wire [8:0] _T_1627; // @[Modules.scala 108:54:@39078.4]
  wire [7:0] _T_1628; // @[Modules.scala 108:54:@39079.4]
  wire [7:0] buffer_14_13; // @[Modules.scala 108:54:@39080.4]
  wire [8:0] _T_1630; // @[Modules.scala 108:54:@39082.4]
  wire [7:0] _T_1631; // @[Modules.scala 108:54:@39083.4]
  wire [7:0] buffer_14_14; // @[Modules.scala 108:54:@39084.4]
  wire [8:0] _T_1639; // @[Modules.scala 108:54:@39100.4]
  wire [7:0] _T_1640; // @[Modules.scala 108:54:@39101.4]
  wire [7:0] buffer_15_6; // @[Modules.scala 108:54:@39102.4]
  wire [8:0] _T_1642; // @[Modules.scala 108:54:@39109.4]
  wire [7:0] _T_1643; // @[Modules.scala 108:54:@39110.4]
  wire [7:0] buffer_15_12; // @[Modules.scala 108:54:@39111.4]
  wire [8:0] _T_1645; // @[Modules.scala 108:54:@39113.4]
  wire [7:0] _T_1646; // @[Modules.scala 108:54:@39114.4]
  wire [7:0] buffer_15_13; // @[Modules.scala 108:54:@39115.4]
  wire [8:0] _T_1648; // @[Modules.scala 108:54:@39118.4]
  wire [7:0] _T_1649; // @[Modules.scala 108:54:@39119.4]
  wire [7:0] buffer_15_15; // @[Modules.scala 108:54:@39120.4]
  assign _GEN_0 = {{6{io_in_2[1]}},io_in_2}; // @[Modules.scala 108:54:@38481.4]
  assign _T_1275 = $signed(8'sh0) + $signed(_GEN_0); // @[Modules.scala 108:54:@38481.4]
  assign _T_1276 = _T_1275[7:0]; // @[Modules.scala 108:54:@38482.4]
  assign buffer_0_2 = $signed(_T_1276); // @[Modules.scala 108:54:@38483.4]
  assign _GEN_1 = {{6{io_in_5[1]}},io_in_5}; // @[Modules.scala 108:54:@38487.4]
  assign _T_1278 = $signed(buffer_0_2) + $signed(_GEN_1); // @[Modules.scala 108:54:@38487.4]
  assign _T_1279 = _T_1278[7:0]; // @[Modules.scala 108:54:@38488.4]
  assign buffer_0_5 = $signed(_T_1279); // @[Modules.scala 108:54:@38489.4]
  assign _GEN_2 = {{6{io_in_6[1]}},io_in_6}; // @[Modules.scala 108:54:@38491.4]
  assign _T_1281 = $signed(buffer_0_5) + $signed(_GEN_2); // @[Modules.scala 108:54:@38491.4]
  assign _T_1282 = _T_1281[7:0]; // @[Modules.scala 108:54:@38492.4]
  assign buffer_0_6 = $signed(_T_1282); // @[Modules.scala 108:54:@38493.4]
  assign _GEN_3 = {{6{io_in_7[1]}},io_in_7}; // @[Modules.scala 108:54:@38495.4]
  assign _T_1284 = $signed(buffer_0_6) + $signed(_GEN_3); // @[Modules.scala 108:54:@38495.4]
  assign _T_1285 = _T_1284[7:0]; // @[Modules.scala 108:54:@38496.4]
  assign buffer_0_7 = $signed(_T_1285); // @[Modules.scala 108:54:@38497.4]
  assign _GEN_4 = {{6{io_in_11[1]}},io_in_11}; // @[Modules.scala 108:54:@38502.4]
  assign _T_1287 = $signed(buffer_0_7) + $signed(_GEN_4); // @[Modules.scala 108:54:@38502.4]
  assign _T_1288 = _T_1287[7:0]; // @[Modules.scala 108:54:@38503.4]
  assign buffer_0_11 = $signed(_T_1288); // @[Modules.scala 108:54:@38504.4]
  assign buffer_1_0 = {{6{io_in_0[1]}},io_in_0}; // @[Modules.scala 91:22:@38478.4]
  assign _GEN_5 = {{6{io_in_1[1]}},io_in_1}; // @[Modules.scala 108:54:@38512.4]
  assign _T_1290 = $signed(buffer_1_0) + $signed(_GEN_5); // @[Modules.scala 108:54:@38512.4]
  assign _T_1291 = _T_1290[7:0]; // @[Modules.scala 108:54:@38513.4]
  assign buffer_1_1 = $signed(_T_1291); // @[Modules.scala 108:54:@38514.4]
  assign _T_1293 = $signed(buffer_1_1) + $signed(_GEN_0); // @[Modules.scala 108:54:@38516.4]
  assign _T_1294 = _T_1293[7:0]; // @[Modules.scala 108:54:@38517.4]
  assign buffer_1_2 = $signed(_T_1294); // @[Modules.scala 108:54:@38518.4]
  assign _GEN_7 = {{6{io_in_4[1]}},io_in_4}; // @[Modules.scala 108:54:@38521.4]
  assign _T_1296 = $signed(buffer_1_2) + $signed(_GEN_7); // @[Modules.scala 108:54:@38521.4]
  assign _T_1297 = _T_1296[7:0]; // @[Modules.scala 108:54:@38522.4]
  assign buffer_1_4 = $signed(_T_1297); // @[Modules.scala 108:54:@38523.4]
  assign _T_1299 = $signed(buffer_1_4) + $signed(_GEN_2); // @[Modules.scala 108:54:@38526.4]
  assign _T_1300 = _T_1299[7:0]; // @[Modules.scala 108:54:@38527.4]
  assign buffer_1_6 = $signed(_T_1300); // @[Modules.scala 108:54:@38528.4]
  assign _GEN_9 = {{6{io_in_12[1]}},io_in_12}; // @[Modules.scala 108:54:@38535.4]
  assign _T_1302 = $signed(buffer_1_6) + $signed(_GEN_9); // @[Modules.scala 108:54:@38535.4]
  assign _T_1303 = _T_1302[7:0]; // @[Modules.scala 108:54:@38536.4]
  assign buffer_1_12 = $signed(_T_1303); // @[Modules.scala 108:54:@38537.4]
  assign _GEN_10 = {{6{io_in_13[1]}},io_in_13}; // @[Modules.scala 108:54:@38539.4]
  assign _T_1305 = $signed(buffer_1_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@38539.4]
  assign _T_1306 = _T_1305[7:0]; // @[Modules.scala 108:54:@38540.4]
  assign buffer_1_13 = $signed(_T_1306); // @[Modules.scala 108:54:@38541.4]
  assign _GEN_11 = {{6{io_in_15[1]}},io_in_15}; // @[Modules.scala 108:54:@38544.4]
  assign _T_1308 = $signed(buffer_1_13) + $signed(_GEN_11); // @[Modules.scala 108:54:@38544.4]
  assign _T_1309 = _T_1308[7:0]; // @[Modules.scala 108:54:@38545.4]
  assign buffer_1_15 = $signed(_T_1309); // @[Modules.scala 108:54:@38546.4]
  assign _T_1311 = $signed(buffer_1_0) + $signed(_GEN_0); // @[Modules.scala 108:54:@38551.4]
  assign _T_1312 = _T_1311[7:0]; // @[Modules.scala 108:54:@38552.4]
  assign buffer_2_2 = $signed(_T_1312); // @[Modules.scala 108:54:@38553.4]
  assign _T_1314 = $signed(buffer_2_2) + $signed(_GEN_7); // @[Modules.scala 108:54:@38556.4]
  assign _T_1315 = _T_1314[7:0]; // @[Modules.scala 108:54:@38557.4]
  assign buffer_2_4 = $signed(_T_1315); // @[Modules.scala 108:54:@38558.4]
  assign _T_1317 = $signed(buffer_2_4) + $signed(_GEN_3); // @[Modules.scala 108:54:@38562.4]
  assign _T_1318 = _T_1317[7:0]; // @[Modules.scala 108:54:@38563.4]
  assign buffer_2_7 = $signed(_T_1318); // @[Modules.scala 108:54:@38564.4]
  assign _GEN_15 = {{6{io_in_8[1]}},io_in_8}; // @[Modules.scala 108:54:@38566.4]
  assign _T_1320 = $signed(buffer_2_7) + $signed(_GEN_15); // @[Modules.scala 108:54:@38566.4]
  assign _T_1321 = _T_1320[7:0]; // @[Modules.scala 108:54:@38567.4]
  assign buffer_2_8 = $signed(_T_1321); // @[Modules.scala 108:54:@38568.4]
  assign _GEN_16 = {{6{io_in_9[1]}},io_in_9}; // @[Modules.scala 108:54:@38570.4]
  assign _T_1323 = $signed(buffer_2_8) + $signed(_GEN_16); // @[Modules.scala 108:54:@38570.4]
  assign _T_1324 = _T_1323[7:0]; // @[Modules.scala 108:54:@38571.4]
  assign buffer_2_9 = $signed(_T_1324); // @[Modules.scala 108:54:@38572.4]
  assign _GEN_17 = {{6{io_in_10[1]}},io_in_10}; // @[Modules.scala 108:54:@38574.4]
  assign _T_1326 = $signed(buffer_2_9) + $signed(_GEN_17); // @[Modules.scala 108:54:@38574.4]
  assign _T_1327 = _T_1326[7:0]; // @[Modules.scala 108:54:@38575.4]
  assign buffer_2_10 = $signed(_T_1327); // @[Modules.scala 108:54:@38576.4]
  assign _T_1329 = $signed(buffer_2_10) + $signed(_GEN_4); // @[Modules.scala 108:54:@38578.4]
  assign _T_1330 = _T_1329[7:0]; // @[Modules.scala 108:54:@38579.4]
  assign buffer_2_11 = $signed(_T_1330); // @[Modules.scala 108:54:@38580.4]
  assign _T_1332 = $signed(buffer_2_11) + $signed(_GEN_9); // @[Modules.scala 108:54:@38582.4]
  assign _T_1333 = _T_1332[7:0]; // @[Modules.scala 108:54:@38583.4]
  assign buffer_2_12 = $signed(_T_1333); // @[Modules.scala 108:54:@38584.4]
  assign _T_1335 = $signed(buffer_2_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@38586.4]
  assign _T_1336 = _T_1335[7:0]; // @[Modules.scala 108:54:@38587.4]
  assign buffer_2_13 = $signed(_T_1336); // @[Modules.scala 108:54:@38588.4]
  assign _T_1338 = $signed(buffer_2_13) + $signed(_GEN_11); // @[Modules.scala 108:54:@38591.4]
  assign _T_1339 = _T_1338[7:0]; // @[Modules.scala 108:54:@38592.4]
  assign buffer_2_15 = $signed(_T_1339); // @[Modules.scala 108:54:@38593.4]
  assign _GEN_22 = {{6{io_in_3[1]}},io_in_3}; // @[Modules.scala 108:54:@38599.4]
  assign _T_1342 = $signed(8'sh0) + $signed(_GEN_22); // @[Modules.scala 108:54:@38599.4]
  assign _T_1343 = _T_1342[7:0]; // @[Modules.scala 108:54:@38600.4]
  assign buffer_3_3 = $signed(_T_1343); // @[Modules.scala 108:54:@38601.4]
  assign _T_1345 = $signed(buffer_3_3) + $signed(_GEN_1); // @[Modules.scala 108:54:@38604.4]
  assign _T_1346 = _T_1345[7:0]; // @[Modules.scala 108:54:@38605.4]
  assign buffer_3_5 = $signed(_T_1346); // @[Modules.scala 108:54:@38606.4]
  assign _T_1348 = $signed(buffer_3_5) + $signed(_GEN_3); // @[Modules.scala 108:54:@38609.4]
  assign _T_1349 = _T_1348[7:0]; // @[Modules.scala 108:54:@38610.4]
  assign buffer_3_7 = $signed(_T_1349); // @[Modules.scala 108:54:@38611.4]
  assign _T_1351 = $signed(buffer_3_7) + $signed(_GEN_15); // @[Modules.scala 108:54:@38613.4]
  assign _T_1352 = _T_1351[7:0]; // @[Modules.scala 108:54:@38614.4]
  assign buffer_3_8 = $signed(_T_1352); // @[Modules.scala 108:54:@38615.4]
  assign _T_1354 = $signed(buffer_3_8) + $signed(_GEN_16); // @[Modules.scala 108:54:@38617.4]
  assign _T_1355 = _T_1354[7:0]; // @[Modules.scala 108:54:@38618.4]
  assign buffer_3_9 = $signed(_T_1355); // @[Modules.scala 108:54:@38619.4]
  assign _T_1357 = $signed(buffer_3_9) + $signed(_GEN_17); // @[Modules.scala 108:54:@38621.4]
  assign _T_1358 = _T_1357[7:0]; // @[Modules.scala 108:54:@38622.4]
  assign buffer_3_10 = $signed(_T_1358); // @[Modules.scala 108:54:@38623.4]
  assign _T_1360 = $signed(buffer_3_10) + $signed(_GEN_9); // @[Modules.scala 108:54:@38626.4]
  assign _T_1361 = _T_1360[7:0]; // @[Modules.scala 108:54:@38627.4]
  assign buffer_3_12 = $signed(_T_1361); // @[Modules.scala 108:54:@38628.4]
  assign _T_1363 = $signed(buffer_3_12) + $signed(_GEN_11); // @[Modules.scala 108:54:@38632.4]
  assign _T_1364 = _T_1363[7:0]; // @[Modules.scala 108:54:@38633.4]
  assign buffer_3_15 = $signed(_T_1364); // @[Modules.scala 108:54:@38634.4]
  assign _T_1378 = $signed(buffer_1_6) + $signed(_GEN_3); // @[Modules.scala 108:54:@38656.4]
  assign _T_1379 = _T_1378[7:0]; // @[Modules.scala 108:54:@38657.4]
  assign buffer_4_7 = $signed(_T_1379); // @[Modules.scala 108:54:@38658.4]
  assign _T_1381 = $signed(buffer_4_7) + $signed(_GEN_15); // @[Modules.scala 108:54:@38660.4]
  assign _T_1382 = _T_1381[7:0]; // @[Modules.scala 108:54:@38661.4]
  assign buffer_4_8 = $signed(_T_1382); // @[Modules.scala 108:54:@38662.4]
  assign _T_1384 = $signed(buffer_4_8) + $signed(_GEN_17); // @[Modules.scala 108:54:@38665.4]
  assign _T_1385 = _T_1384[7:0]; // @[Modules.scala 108:54:@38666.4]
  assign buffer_4_10 = $signed(_T_1385); // @[Modules.scala 108:54:@38667.4]
  assign _T_1387 = $signed(buffer_4_10) + $signed(_GEN_4); // @[Modules.scala 108:54:@38669.4]
  assign _T_1388 = _T_1387[7:0]; // @[Modules.scala 108:54:@38670.4]
  assign buffer_4_11 = $signed(_T_1388); // @[Modules.scala 108:54:@38671.4]
  assign _T_1391 = $signed(8'sh0) + $signed(_GEN_5); // @[Modules.scala 108:54:@38679.4]
  assign _T_1392 = _T_1391[7:0]; // @[Modules.scala 108:54:@38680.4]
  assign buffer_5_1 = $signed(_T_1392); // @[Modules.scala 108:54:@38681.4]
  assign _T_1394 = $signed(buffer_5_1) + $signed(_GEN_0); // @[Modules.scala 108:54:@38683.4]
  assign _T_1395 = _T_1394[7:0]; // @[Modules.scala 108:54:@38684.4]
  assign buffer_5_2 = $signed(_T_1395); // @[Modules.scala 108:54:@38685.4]
  assign _T_1397 = $signed(buffer_5_2) + $signed(_GEN_7); // @[Modules.scala 108:54:@38688.4]
  assign _T_1398 = _T_1397[7:0]; // @[Modules.scala 108:54:@38689.4]
  assign buffer_5_4 = $signed(_T_1398); // @[Modules.scala 108:54:@38690.4]
  assign _T_1400 = $signed(buffer_5_4) + $signed(_GEN_3); // @[Modules.scala 108:54:@38694.4]
  assign _T_1401 = _T_1400[7:0]; // @[Modules.scala 108:54:@38695.4]
  assign buffer_5_7 = $signed(_T_1401); // @[Modules.scala 108:54:@38696.4]
  assign _T_1403 = $signed(buffer_5_7) + $signed(_GEN_16); // @[Modules.scala 108:54:@38699.4]
  assign _T_1404 = _T_1403[7:0]; // @[Modules.scala 108:54:@38700.4]
  assign buffer_5_9 = $signed(_T_1404); // @[Modules.scala 108:54:@38701.4]
  assign _T_1406 = $signed(buffer_5_9) + $signed(_GEN_17); // @[Modules.scala 108:54:@38703.4]
  assign _T_1407 = _T_1406[7:0]; // @[Modules.scala 108:54:@38704.4]
  assign buffer_5_10 = $signed(_T_1407); // @[Modules.scala 108:54:@38705.4]
  assign _T_1409 = $signed(buffer_5_10) + $signed(_GEN_4); // @[Modules.scala 108:54:@38707.4]
  assign _T_1410 = _T_1409[7:0]; // @[Modules.scala 108:54:@38708.4]
  assign buffer_5_11 = $signed(_T_1410); // @[Modules.scala 108:54:@38709.4]
  assign _T_1415 = $signed(buffer_2_2) + $signed(_GEN_1); // @[Modules.scala 108:54:@38724.4]
  assign _T_1416 = _T_1415[7:0]; // @[Modules.scala 108:54:@38725.4]
  assign buffer_6_5 = $signed(_T_1416); // @[Modules.scala 108:54:@38726.4]
  assign _T_1418 = $signed(buffer_6_5) + $signed(_GEN_3); // @[Modules.scala 108:54:@38729.4]
  assign _T_1419 = _T_1418[7:0]; // @[Modules.scala 108:54:@38730.4]
  assign buffer_6_7 = $signed(_T_1419); // @[Modules.scala 108:54:@38731.4]
  assign _T_1421 = $signed(buffer_6_7) + $signed(_GEN_15); // @[Modules.scala 108:54:@38733.4]
  assign _T_1422 = _T_1421[7:0]; // @[Modules.scala 108:54:@38734.4]
  assign buffer_6_8 = $signed(_T_1422); // @[Modules.scala 108:54:@38735.4]
  assign _T_1424 = $signed(buffer_6_8) + $signed(_GEN_4); // @[Modules.scala 108:54:@38739.4]
  assign _T_1425 = _T_1424[7:0]; // @[Modules.scala 108:54:@38740.4]
  assign buffer_6_11 = $signed(_T_1425); // @[Modules.scala 108:54:@38741.4]
  assign _T_1427 = $signed(buffer_6_11) + $signed(_GEN_10); // @[Modules.scala 108:54:@38744.4]
  assign _T_1428 = _T_1427[7:0]; // @[Modules.scala 108:54:@38745.4]
  assign buffer_6_13 = $signed(_T_1428); // @[Modules.scala 108:54:@38746.4]
  assign _GEN_51 = {{6{io_in_14[1]}},io_in_14}; // @[Modules.scala 108:54:@38748.4]
  assign _T_1430 = $signed(buffer_6_13) + $signed(_GEN_51); // @[Modules.scala 108:54:@38748.4]
  assign _T_1431 = _T_1430[7:0]; // @[Modules.scala 108:54:@38749.4]
  assign buffer_6_14 = $signed(_T_1431); // @[Modules.scala 108:54:@38750.4]
  assign _T_1433 = $signed(buffer_1_0) + $signed(_GEN_22); // @[Modules.scala 108:54:@38757.4]
  assign _T_1434 = _T_1433[7:0]; // @[Modules.scala 108:54:@38758.4]
  assign buffer_7_3 = $signed(_T_1434); // @[Modules.scala 108:54:@38759.4]
  assign _T_1436 = $signed(buffer_7_3) + $signed(_GEN_1); // @[Modules.scala 108:54:@38762.4]
  assign _T_1437 = _T_1436[7:0]; // @[Modules.scala 108:54:@38763.4]
  assign buffer_7_5 = $signed(_T_1437); // @[Modules.scala 108:54:@38764.4]
  assign _T_1439 = $signed(buffer_7_5) + $signed(_GEN_2); // @[Modules.scala 108:54:@38766.4]
  assign _T_1440 = _T_1439[7:0]; // @[Modules.scala 108:54:@38767.4]
  assign buffer_7_6 = $signed(_T_1440); // @[Modules.scala 108:54:@38768.4]
  assign _T_1442 = $signed(buffer_7_6) + $signed(_GEN_15); // @[Modules.scala 108:54:@38771.4]
  assign _T_1443 = _T_1442[7:0]; // @[Modules.scala 108:54:@38772.4]
  assign buffer_7_8 = $signed(_T_1443); // @[Modules.scala 108:54:@38773.4]
  assign _T_1445 = $signed(buffer_7_8) + $signed(_GEN_16); // @[Modules.scala 108:54:@38775.4]
  assign _T_1446 = _T_1445[7:0]; // @[Modules.scala 108:54:@38776.4]
  assign buffer_7_9 = $signed(_T_1446); // @[Modules.scala 108:54:@38777.4]
  assign _T_1448 = $signed(buffer_7_9) + $signed(_GEN_17); // @[Modules.scala 108:54:@38779.4]
  assign _T_1449 = _T_1448[7:0]; // @[Modules.scala 108:54:@38780.4]
  assign buffer_7_10 = $signed(_T_1449); // @[Modules.scala 108:54:@38781.4]
  assign _T_1451 = $signed(buffer_7_10) + $signed(_GEN_11); // @[Modules.scala 108:54:@38787.4]
  assign _T_1452 = _T_1451[7:0]; // @[Modules.scala 108:54:@38788.4]
  assign buffer_7_15 = $signed(_T_1452); // @[Modules.scala 108:54:@38789.4]
  assign _T_1460 = $signed(buffer_6_5) + $signed(_GEN_2); // @[Modules.scala 108:54:@38804.4]
  assign _T_1461 = _T_1460[7:0]; // @[Modules.scala 108:54:@38805.4]
  assign buffer_8_6 = $signed(_T_1461); // @[Modules.scala 108:54:@38806.4]
  assign _T_1463 = $signed(buffer_8_6) + $signed(_GEN_3); // @[Modules.scala 108:54:@38808.4]
  assign _T_1464 = _T_1463[7:0]; // @[Modules.scala 108:54:@38809.4]
  assign buffer_8_7 = $signed(_T_1464); // @[Modules.scala 108:54:@38810.4]
  assign _T_1466 = $signed(buffer_8_7) + $signed(_GEN_15); // @[Modules.scala 108:54:@38812.4]
  assign _T_1467 = _T_1466[7:0]; // @[Modules.scala 108:54:@38813.4]
  assign buffer_8_8 = $signed(_T_1467); // @[Modules.scala 108:54:@38814.4]
  assign _T_1469 = $signed(buffer_8_8) + $signed(_GEN_17); // @[Modules.scala 108:54:@38817.4]
  assign _T_1470 = _T_1469[7:0]; // @[Modules.scala 108:54:@38818.4]
  assign buffer_8_10 = $signed(_T_1470); // @[Modules.scala 108:54:@38819.4]
  assign _T_1472 = $signed(buffer_8_10) + $signed(_GEN_9); // @[Modules.scala 108:54:@38822.4]
  assign _T_1473 = _T_1472[7:0]; // @[Modules.scala 108:54:@38823.4]
  assign buffer_8_12 = $signed(_T_1473); // @[Modules.scala 108:54:@38824.4]
  assign _T_1475 = $signed(buffer_8_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@38826.4]
  assign _T_1476 = _T_1475[7:0]; // @[Modules.scala 108:54:@38827.4]
  assign buffer_8_13 = $signed(_T_1476); // @[Modules.scala 108:54:@38828.4]
  assign _T_1478 = $signed(buffer_8_13) + $signed(_GEN_11); // @[Modules.scala 108:54:@38831.4]
  assign _T_1479 = _T_1478[7:0]; // @[Modules.scala 108:54:@38832.4]
  assign buffer_8_15 = $signed(_T_1479); // @[Modules.scala 108:54:@38833.4]
  assign _T_1487 = $signed(buffer_1_2) + $signed(_GEN_22); // @[Modules.scala 108:54:@38845.4]
  assign _T_1488 = _T_1487[7:0]; // @[Modules.scala 108:54:@38846.4]
  assign buffer_9_3 = $signed(_T_1488); // @[Modules.scala 108:54:@38847.4]
  assign _T_1490 = $signed(buffer_9_3) + $signed(_GEN_7); // @[Modules.scala 108:54:@38849.4]
  assign _T_1491 = _T_1490[7:0]; // @[Modules.scala 108:54:@38850.4]
  assign buffer_9_4 = $signed(_T_1491); // @[Modules.scala 108:54:@38851.4]
  assign _T_1493 = $signed(buffer_9_4) + $signed(_GEN_2); // @[Modules.scala 108:54:@38854.4]
  assign _T_1494 = _T_1493[7:0]; // @[Modules.scala 108:54:@38855.4]
  assign buffer_9_6 = $signed(_T_1494); // @[Modules.scala 108:54:@38856.4]
  assign _T_1496 = $signed(buffer_9_6) + $signed(_GEN_15); // @[Modules.scala 108:54:@38859.4]
  assign _T_1497 = _T_1496[7:0]; // @[Modules.scala 108:54:@38860.4]
  assign buffer_9_8 = $signed(_T_1497); // @[Modules.scala 108:54:@38861.4]
  assign _T_1499 = $signed(buffer_9_8) + $signed(_GEN_51); // @[Modules.scala 108:54:@38868.4]
  assign _T_1500 = _T_1499[7:0]; // @[Modules.scala 108:54:@38869.4]
  assign buffer_9_14 = $signed(_T_1500); // @[Modules.scala 108:54:@38870.4]
  assign _T_1509 = $signed(buffer_5_2) + $signed(_GEN_22); // @[Modules.scala 108:54:@38883.4]
  assign _T_1510 = _T_1509[7:0]; // @[Modules.scala 108:54:@38884.4]
  assign buffer_10_3 = $signed(_T_1510); // @[Modules.scala 108:54:@38885.4]
  assign _T_1512 = $signed(buffer_10_3) + $signed(_GEN_17); // @[Modules.scala 108:54:@38893.4]
  assign _T_1513 = _T_1512[7:0]; // @[Modules.scala 108:54:@38894.4]
  assign buffer_10_10 = $signed(_T_1513); // @[Modules.scala 108:54:@38895.4]
  assign _T_1515 = $signed(buffer_10_10) + $signed(_GEN_4); // @[Modules.scala 108:54:@38897.4]
  assign _T_1516 = _T_1515[7:0]; // @[Modules.scala 108:54:@38898.4]
  assign buffer_10_11 = $signed(_T_1516); // @[Modules.scala 108:54:@38899.4]
  assign _T_1518 = $signed(buffer_10_11) + $signed(_GEN_9); // @[Modules.scala 108:54:@38901.4]
  assign _T_1519 = _T_1518[7:0]; // @[Modules.scala 108:54:@38902.4]
  assign buffer_10_12 = $signed(_T_1519); // @[Modules.scala 108:54:@38903.4]
  assign _T_1521 = $signed(buffer_10_12) + $signed(_GEN_11); // @[Modules.scala 108:54:@38907.4]
  assign _T_1522 = _T_1521[7:0]; // @[Modules.scala 108:54:@38908.4]
  assign buffer_10_15 = $signed(_T_1522); // @[Modules.scala 108:54:@38909.4]
  assign _T_1528 = $signed(buffer_3_3) + $signed(_GEN_7); // @[Modules.scala 108:54:@38919.4]
  assign _T_1529 = _T_1528[7:0]; // @[Modules.scala 108:54:@38920.4]
  assign buffer_11_4 = $signed(_T_1529); // @[Modules.scala 108:54:@38921.4]
  assign _T_1531 = $signed(buffer_11_4) + $signed(_GEN_2); // @[Modules.scala 108:54:@38924.4]
  assign _T_1532 = _T_1531[7:0]; // @[Modules.scala 108:54:@38925.4]
  assign buffer_11_6 = $signed(_T_1532); // @[Modules.scala 108:54:@38926.4]
  assign _T_1534 = $signed(buffer_11_6) + $signed(_GEN_15); // @[Modules.scala 108:54:@38929.4]
  assign _T_1535 = _T_1534[7:0]; // @[Modules.scala 108:54:@38930.4]
  assign buffer_11_8 = $signed(_T_1535); // @[Modules.scala 108:54:@38931.4]
  assign _T_1537 = $signed(buffer_11_8) + $signed(_GEN_9); // @[Modules.scala 108:54:@38936.4]
  assign _T_1538 = _T_1537[7:0]; // @[Modules.scala 108:54:@38937.4]
  assign buffer_11_12 = $signed(_T_1538); // @[Modules.scala 108:54:@38938.4]
  assign _T_1540 = $signed(buffer_11_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@38940.4]
  assign _T_1541 = _T_1540[7:0]; // @[Modules.scala 108:54:@38941.4]
  assign buffer_11_13 = $signed(_T_1541); // @[Modules.scala 108:54:@38942.4]
  assign _T_1543 = $signed(buffer_11_13) + $signed(_GEN_11); // @[Modules.scala 108:54:@38945.4]
  assign _T_1544 = _T_1543[7:0]; // @[Modules.scala 108:54:@38946.4]
  assign buffer_11_15 = $signed(_T_1544); // @[Modules.scala 108:54:@38947.4]
  assign _T_1549 = $signed(buffer_1_1) + $signed(_GEN_22); // @[Modules.scala 108:54:@38956.4]
  assign _T_1550 = _T_1549[7:0]; // @[Modules.scala 108:54:@38957.4]
  assign buffer_12_3 = $signed(_T_1550); // @[Modules.scala 108:54:@38958.4]
  assign _T_1552 = $signed(buffer_12_3) + $signed(_GEN_7); // @[Modules.scala 108:54:@38960.4]
  assign _T_1553 = _T_1552[7:0]; // @[Modules.scala 108:54:@38961.4]
  assign buffer_12_4 = $signed(_T_1553); // @[Modules.scala 108:54:@38962.4]
  assign _T_1555 = $signed(buffer_12_4) + $signed(_GEN_3); // @[Modules.scala 108:54:@38966.4]
  assign _T_1556 = _T_1555[7:0]; // @[Modules.scala 108:54:@38967.4]
  assign buffer_12_7 = $signed(_T_1556); // @[Modules.scala 108:54:@38968.4]
  assign _T_1558 = $signed(buffer_12_7) + $signed(_GEN_16); // @[Modules.scala 108:54:@38971.4]
  assign _T_1559 = _T_1558[7:0]; // @[Modules.scala 108:54:@38972.4]
  assign buffer_12_9 = $signed(_T_1559); // @[Modules.scala 108:54:@38973.4]
  assign _T_1561 = $signed(buffer_12_9) + $signed(_GEN_17); // @[Modules.scala 108:54:@38975.4]
  assign _T_1562 = _T_1561[7:0]; // @[Modules.scala 108:54:@38976.4]
  assign buffer_12_10 = $signed(_T_1562); // @[Modules.scala 108:54:@38977.4]
  assign _T_1564 = $signed(buffer_12_10) + $signed(_GEN_9); // @[Modules.scala 108:54:@38980.4]
  assign _T_1565 = _T_1564[7:0]; // @[Modules.scala 108:54:@38981.4]
  assign buffer_12_12 = $signed(_T_1565); // @[Modules.scala 108:54:@38982.4]
  assign _T_1567 = $signed(buffer_12_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@38984.4]
  assign _T_1568 = _T_1567[7:0]; // @[Modules.scala 108:54:@38985.4]
  assign buffer_12_13 = $signed(_T_1568); // @[Modules.scala 108:54:@38986.4]
  assign _T_1570 = $signed(buffer_12_13) + $signed(_GEN_51); // @[Modules.scala 108:54:@38988.4]
  assign _T_1571 = _T_1570[7:0]; // @[Modules.scala 108:54:@38989.4]
  assign buffer_12_14 = $signed(_T_1571); // @[Modules.scala 108:54:@38990.4]
  assign _T_1573 = $signed(buffer_12_14) + $signed(_GEN_11); // @[Modules.scala 108:54:@38992.4]
  assign _T_1574 = _T_1573[7:0]; // @[Modules.scala 108:54:@38993.4]
  assign buffer_12_15 = $signed(_T_1574); // @[Modules.scala 108:54:@38994.4]
  assign _T_1588 = $signed(buffer_9_4) + $signed(_GEN_3); // @[Modules.scala 108:54:@39016.4]
  assign _T_1589 = _T_1588[7:0]; // @[Modules.scala 108:54:@39017.4]
  assign buffer_13_7 = $signed(_T_1589); // @[Modules.scala 108:54:@39018.4]
  assign _T_1591 = $signed(buffer_13_7) + $signed(_GEN_15); // @[Modules.scala 108:54:@39020.4]
  assign _T_1592 = _T_1591[7:0]; // @[Modules.scala 108:54:@39021.4]
  assign buffer_13_8 = $signed(_T_1592); // @[Modules.scala 108:54:@39022.4]
  assign _T_1594 = $signed(buffer_13_8) + $signed(_GEN_4); // @[Modules.scala 108:54:@39026.4]
  assign _T_1595 = _T_1594[7:0]; // @[Modules.scala 108:54:@39027.4]
  assign buffer_13_11 = $signed(_T_1595); // @[Modules.scala 108:54:@39028.4]
  assign _T_1597 = $signed(buffer_13_11) + $signed(_GEN_9); // @[Modules.scala 108:54:@39030.4]
  assign _T_1598 = _T_1597[7:0]; // @[Modules.scala 108:54:@39031.4]
  assign buffer_13_12 = $signed(_T_1598); // @[Modules.scala 108:54:@39032.4]
  assign _T_1600 = $signed(buffer_13_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@39034.4]
  assign _T_1601 = _T_1600[7:0]; // @[Modules.scala 108:54:@39035.4]
  assign buffer_13_13 = $signed(_T_1601); // @[Modules.scala 108:54:@39036.4]
  assign _T_1603 = $signed(buffer_13_13) + $signed(_GEN_11); // @[Modules.scala 108:54:@39039.4]
  assign _T_1604 = _T_1603[7:0]; // @[Modules.scala 108:54:@39040.4]
  assign buffer_13_15 = $signed(_T_1604); // @[Modules.scala 108:54:@39041.4]
  assign _T_1612 = $signed(buffer_2_4) + $signed(_GEN_1); // @[Modules.scala 108:54:@39055.4]
  assign _T_1613 = _T_1612[7:0]; // @[Modules.scala 108:54:@39056.4]
  assign buffer_14_5 = $signed(_T_1613); // @[Modules.scala 108:54:@39057.4]
  assign _T_1615 = $signed(buffer_14_5) + $signed(_GEN_2); // @[Modules.scala 108:54:@39059.4]
  assign _T_1616 = _T_1615[7:0]; // @[Modules.scala 108:54:@39060.4]
  assign buffer_14_6 = $signed(_T_1616); // @[Modules.scala 108:54:@39061.4]
  assign _T_1618 = $signed(buffer_14_6) + $signed(_GEN_3); // @[Modules.scala 108:54:@39063.4]
  assign _T_1619 = _T_1618[7:0]; // @[Modules.scala 108:54:@39064.4]
  assign buffer_14_7 = $signed(_T_1619); // @[Modules.scala 108:54:@39065.4]
  assign _T_1621 = $signed(buffer_14_7) + $signed(_GEN_16); // @[Modules.scala 108:54:@39068.4]
  assign _T_1622 = _T_1621[7:0]; // @[Modules.scala 108:54:@39069.4]
  assign buffer_14_9 = $signed(_T_1622); // @[Modules.scala 108:54:@39070.4]
  assign _T_1624 = $signed(buffer_14_9) + $signed(_GEN_9); // @[Modules.scala 108:54:@39074.4]
  assign _T_1625 = _T_1624[7:0]; // @[Modules.scala 108:54:@39075.4]
  assign buffer_14_12 = $signed(_T_1625); // @[Modules.scala 108:54:@39076.4]
  assign _T_1627 = $signed(buffer_14_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@39078.4]
  assign _T_1628 = _T_1627[7:0]; // @[Modules.scala 108:54:@39079.4]
  assign buffer_14_13 = $signed(_T_1628); // @[Modules.scala 108:54:@39080.4]
  assign _T_1630 = $signed(buffer_14_13) + $signed(_GEN_51); // @[Modules.scala 108:54:@39082.4]
  assign _T_1631 = _T_1630[7:0]; // @[Modules.scala 108:54:@39083.4]
  assign buffer_14_14 = $signed(_T_1631); // @[Modules.scala 108:54:@39084.4]
  assign _T_1639 = $signed(buffer_1_2) + $signed(_GEN_2); // @[Modules.scala 108:54:@39100.4]
  assign _T_1640 = _T_1639[7:0]; // @[Modules.scala 108:54:@39101.4]
  assign buffer_15_6 = $signed(_T_1640); // @[Modules.scala 108:54:@39102.4]
  assign _T_1642 = $signed(buffer_15_6) + $signed(_GEN_9); // @[Modules.scala 108:54:@39109.4]
  assign _T_1643 = _T_1642[7:0]; // @[Modules.scala 108:54:@39110.4]
  assign buffer_15_12 = $signed(_T_1643); // @[Modules.scala 108:54:@39111.4]
  assign _T_1645 = $signed(buffer_15_12) + $signed(_GEN_10); // @[Modules.scala 108:54:@39113.4]
  assign _T_1646 = _T_1645[7:0]; // @[Modules.scala 108:54:@39114.4]
  assign buffer_15_13 = $signed(_T_1646); // @[Modules.scala 108:54:@39115.4]
  assign _T_1648 = $signed(buffer_15_13) + $signed(_GEN_11); // @[Modules.scala 108:54:@39118.4]
  assign _T_1649 = _T_1648[7:0]; // @[Modules.scala 108:54:@39119.4]
  assign buffer_15_15 = $signed(_T_1649); // @[Modules.scala 108:54:@39120.4]
  assign io_out_0 = buffer_0_11;
  assign io_out_1 = buffer_1_15;
  assign io_out_2 = buffer_2_15;
  assign io_out_3 = buffer_3_15;
  assign io_out_4 = buffer_4_11;
  assign io_out_5 = buffer_5_11;
  assign io_out_6 = buffer_6_14;
  assign io_out_7 = buffer_7_15;
  assign io_out_8 = buffer_8_15;
  assign io_out_9 = buffer_9_14;
  assign io_out_10 = buffer_10_15;
  assign io_out_11 = buffer_11_15;
  assign io_out_12 = buffer_12_15;
  assign io_out_13 = buffer_13_15;
  assign io_out_14 = buffer_14_14;
  assign io_out_15 = buffer_15_15;
endmodule
module ShifBatchNorm_1( // @[:@39124.2]
  input  [7:0] io_in_0, // @[:@39127.4]
  input  [7:0] io_in_1, // @[:@39127.4]
  input  [7:0] io_in_2, // @[:@39127.4]
  input  [7:0] io_in_3, // @[:@39127.4]
  input  [7:0] io_in_4, // @[:@39127.4]
  input  [7:0] io_in_5, // @[:@39127.4]
  input  [7:0] io_in_6, // @[:@39127.4]
  input  [7:0] io_in_7, // @[:@39127.4]
  input  [7:0] io_in_8, // @[:@39127.4]
  input  [7:0] io_in_9, // @[:@39127.4]
  input  [7:0] io_in_10, // @[:@39127.4]
  input  [7:0] io_in_11, // @[:@39127.4]
  input  [7:0] io_in_12, // @[:@39127.4]
  input  [7:0] io_in_13, // @[:@39127.4]
  input  [7:0] io_in_14, // @[:@39127.4]
  input  [7:0] io_in_15, // @[:@39127.4]
  output [7:0] io_out_0, // @[:@39127.4]
  output [7:0] io_out_1, // @[:@39127.4]
  output [7:0] io_out_2, // @[:@39127.4]
  output [7:0] io_out_3, // @[:@39127.4]
  output [7:0] io_out_4, // @[:@39127.4]
  output [7:0] io_out_5, // @[:@39127.4]
  output [7:0] io_out_6, // @[:@39127.4]
  output [7:0] io_out_7, // @[:@39127.4]
  output [7:0] io_out_8, // @[:@39127.4]
  output [7:0] io_out_9, // @[:@39127.4]
  output [7:0] io_out_10, // @[:@39127.4]
  output [7:0] io_out_11, // @[:@39127.4]
  output [7:0] io_out_12, // @[:@39127.4]
  output [7:0] io_out_13, // @[:@39127.4]
  output [7:0] io_out_14, // @[:@39127.4]
  output [7:0] io_out_15 // @[:@39127.4]
);
  wire [8:0] _T_108; // @[Modules.scala 132:28:@39132.4]
  wire [7:0] _T_109; // @[Modules.scala 132:28:@39133.4]
  wire [7:0] c_x_0; // @[Modules.scala 132:28:@39134.4]
  wire [22:0] _GEN_0; // @[Modules.scala 137:32:@39136.4]
  wire [22:0] _T_112; // @[Modules.scala 137:32:@39136.4]
  wire [7:0] _GEN_1; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_0; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_2; // @[Modules.scala 139:37:@39138.4]
  wire [22:0] _T_114; // @[Modules.scala 139:37:@39138.4]
  wire [7:0] _GEN_3; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_0; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_116; // @[Modules.scala 140:38:@39140.4]
  wire [7:0] _T_117; // @[Modules.scala 140:38:@39141.4]
  wire [7:0] _T_118; // @[Modules.scala 140:38:@39142.4]
  wire [8:0] _T_120; // @[Modules.scala 132:28:@39144.4]
  wire [7:0] _T_121; // @[Modules.scala 132:28:@39145.4]
  wire [7:0] c_x_1; // @[Modules.scala 132:28:@39146.4]
  wire [22:0] _GEN_4; // @[Modules.scala 137:32:@39148.4]
  wire [22:0] _T_124; // @[Modules.scala 137:32:@39148.4]
  wire [7:0] _GEN_5; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_1; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_6; // @[Modules.scala 139:37:@39150.4]
  wire [22:0] _T_126; // @[Modules.scala 139:37:@39150.4]
  wire [7:0] _GEN_7; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_1; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_128; // @[Modules.scala 140:38:@39152.4]
  wire [7:0] _T_129; // @[Modules.scala 140:38:@39153.4]
  wire [7:0] _T_130; // @[Modules.scala 140:38:@39154.4]
  wire [8:0] _T_132; // @[Modules.scala 132:28:@39156.4]
  wire [7:0] _T_133; // @[Modules.scala 132:28:@39157.4]
  wire [7:0] c_x_2; // @[Modules.scala 132:28:@39158.4]
  wire [22:0] _GEN_8; // @[Modules.scala 137:32:@39160.4]
  wire [22:0] _T_136; // @[Modules.scala 137:32:@39160.4]
  wire [7:0] _GEN_9; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_2; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_10; // @[Modules.scala 139:37:@39162.4]
  wire [22:0] _T_138; // @[Modules.scala 139:37:@39162.4]
  wire [7:0] _GEN_11; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_2; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_140; // @[Modules.scala 140:38:@39164.4]
  wire [7:0] _T_141; // @[Modules.scala 140:38:@39165.4]
  wire [7:0] _T_142; // @[Modules.scala 140:38:@39166.4]
  wire [8:0] _T_144; // @[Modules.scala 132:28:@39168.4]
  wire [7:0] _T_145; // @[Modules.scala 132:28:@39169.4]
  wire [7:0] c_x_3; // @[Modules.scala 132:28:@39170.4]
  wire [22:0] _GEN_12; // @[Modules.scala 137:32:@39172.4]
  wire [22:0] _T_148; // @[Modules.scala 137:32:@39172.4]
  wire [7:0] _GEN_13; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_3; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_14; // @[Modules.scala 139:37:@39174.4]
  wire [22:0] _T_150; // @[Modules.scala 139:37:@39174.4]
  wire [7:0] _GEN_15; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_3; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_152; // @[Modules.scala 140:38:@39176.4]
  wire [7:0] _T_153; // @[Modules.scala 140:38:@39177.4]
  wire [7:0] _T_154; // @[Modules.scala 140:38:@39178.4]
  wire [8:0] _T_156; // @[Modules.scala 132:28:@39180.4]
  wire [7:0] _T_157; // @[Modules.scala 132:28:@39181.4]
  wire [7:0] c_x_4; // @[Modules.scala 132:28:@39182.4]
  wire [22:0] _GEN_16; // @[Modules.scala 137:32:@39184.4]
  wire [22:0] _T_160; // @[Modules.scala 137:32:@39184.4]
  wire [7:0] _GEN_17; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_4; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_18; // @[Modules.scala 139:37:@39186.4]
  wire [22:0] _T_162; // @[Modules.scala 139:37:@39186.4]
  wire [7:0] _GEN_19; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_4; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_164; // @[Modules.scala 140:38:@39188.4]
  wire [7:0] _T_165; // @[Modules.scala 140:38:@39189.4]
  wire [7:0] _T_166; // @[Modules.scala 140:38:@39190.4]
  wire [8:0] _T_168; // @[Modules.scala 132:28:@39192.4]
  wire [7:0] _T_169; // @[Modules.scala 132:28:@39193.4]
  wire [7:0] c_x_5; // @[Modules.scala 132:28:@39194.4]
  wire [22:0] _GEN_20; // @[Modules.scala 137:32:@39196.4]
  wire [22:0] _T_172; // @[Modules.scala 137:32:@39196.4]
  wire [7:0] _GEN_21; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_5; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_22; // @[Modules.scala 139:37:@39198.4]
  wire [22:0] _T_174; // @[Modules.scala 139:37:@39198.4]
  wire [7:0] _GEN_23; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_5; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_176; // @[Modules.scala 140:38:@39200.4]
  wire [7:0] _T_177; // @[Modules.scala 140:38:@39201.4]
  wire [7:0] _T_178; // @[Modules.scala 140:38:@39202.4]
  wire [8:0] _T_180; // @[Modules.scala 132:28:@39204.4]
  wire [7:0] _T_181; // @[Modules.scala 132:28:@39205.4]
  wire [7:0] c_x_6; // @[Modules.scala 132:28:@39206.4]
  wire [22:0] _GEN_24; // @[Modules.scala 137:32:@39208.4]
  wire [22:0] _T_184; // @[Modules.scala 137:32:@39208.4]
  wire [7:0] _GEN_25; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_6; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_26; // @[Modules.scala 139:37:@39210.4]
  wire [22:0] _T_186; // @[Modules.scala 139:37:@39210.4]
  wire [7:0] _GEN_27; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_6; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_188; // @[Modules.scala 140:38:@39212.4]
  wire [7:0] _T_189; // @[Modules.scala 140:38:@39213.4]
  wire [7:0] _T_190; // @[Modules.scala 140:38:@39214.4]
  wire [8:0] _T_192; // @[Modules.scala 132:28:@39216.4]
  wire [7:0] _T_193; // @[Modules.scala 132:28:@39217.4]
  wire [7:0] c_x_7; // @[Modules.scala 132:28:@39218.4]
  wire [22:0] _GEN_28; // @[Modules.scala 137:32:@39220.4]
  wire [22:0] _T_196; // @[Modules.scala 137:32:@39220.4]
  wire [7:0] _GEN_29; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_7; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_30; // @[Modules.scala 139:37:@39222.4]
  wire [22:0] _T_198; // @[Modules.scala 139:37:@39222.4]
  wire [7:0] _GEN_31; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_7; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_200; // @[Modules.scala 140:38:@39224.4]
  wire [7:0] _T_201; // @[Modules.scala 140:38:@39225.4]
  wire [7:0] _T_202; // @[Modules.scala 140:38:@39226.4]
  wire [8:0] _T_204; // @[Modules.scala 132:28:@39228.4]
  wire [7:0] _T_205; // @[Modules.scala 132:28:@39229.4]
  wire [7:0] c_x_8; // @[Modules.scala 132:28:@39230.4]
  wire [22:0] _GEN_32; // @[Modules.scala 137:32:@39232.4]
  wire [22:0] _T_208; // @[Modules.scala 137:32:@39232.4]
  wire [7:0] _GEN_33; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_8; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_34; // @[Modules.scala 139:37:@39234.4]
  wire [22:0] _T_210; // @[Modules.scala 139:37:@39234.4]
  wire [7:0] _GEN_35; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_8; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_212; // @[Modules.scala 140:38:@39236.4]
  wire [7:0] _T_213; // @[Modules.scala 140:38:@39237.4]
  wire [7:0] _T_214; // @[Modules.scala 140:38:@39238.4]
  wire [8:0] _T_216; // @[Modules.scala 132:28:@39240.4]
  wire [7:0] _T_217; // @[Modules.scala 132:28:@39241.4]
  wire [7:0] c_x_9; // @[Modules.scala 132:28:@39242.4]
  wire [22:0] _GEN_36; // @[Modules.scala 137:32:@39244.4]
  wire [22:0] _T_220; // @[Modules.scala 137:32:@39244.4]
  wire [7:0] _GEN_37; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_9; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_38; // @[Modules.scala 139:37:@39246.4]
  wire [22:0] _T_222; // @[Modules.scala 139:37:@39246.4]
  wire [7:0] _GEN_39; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_9; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_224; // @[Modules.scala 140:38:@39248.4]
  wire [7:0] _T_225; // @[Modules.scala 140:38:@39249.4]
  wire [7:0] _T_226; // @[Modules.scala 140:38:@39250.4]
  wire [8:0] _T_228; // @[Modules.scala 132:28:@39252.4]
  wire [7:0] _T_229; // @[Modules.scala 132:28:@39253.4]
  wire [7:0] c_x_10; // @[Modules.scala 132:28:@39254.4]
  wire [22:0] _GEN_40; // @[Modules.scala 137:32:@39256.4]
  wire [22:0] _T_232; // @[Modules.scala 137:32:@39256.4]
  wire [7:0] _GEN_41; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_10; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_42; // @[Modules.scala 139:37:@39258.4]
  wire [22:0] _T_234; // @[Modules.scala 139:37:@39258.4]
  wire [7:0] _GEN_43; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_10; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_236; // @[Modules.scala 140:38:@39260.4]
  wire [7:0] _T_237; // @[Modules.scala 140:38:@39261.4]
  wire [7:0] _T_238; // @[Modules.scala 140:38:@39262.4]
  wire [8:0] _T_240; // @[Modules.scala 132:28:@39264.4]
  wire [7:0] _T_241; // @[Modules.scala 132:28:@39265.4]
  wire [7:0] c_x_11; // @[Modules.scala 132:28:@39266.4]
  wire [22:0] _GEN_44; // @[Modules.scala 137:32:@39268.4]
  wire [22:0] _T_244; // @[Modules.scala 137:32:@39268.4]
  wire [7:0] _GEN_45; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_11; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_46; // @[Modules.scala 139:37:@39270.4]
  wire [22:0] _T_246; // @[Modules.scala 139:37:@39270.4]
  wire [7:0] _GEN_47; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_11; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_248; // @[Modules.scala 140:38:@39272.4]
  wire [7:0] _T_249; // @[Modules.scala 140:38:@39273.4]
  wire [7:0] _T_250; // @[Modules.scala 140:38:@39274.4]
  wire [8:0] _T_252; // @[Modules.scala 132:28:@39276.4]
  wire [7:0] _T_253; // @[Modules.scala 132:28:@39277.4]
  wire [7:0] c_x_12; // @[Modules.scala 132:28:@39278.4]
  wire [22:0] _GEN_48; // @[Modules.scala 137:32:@39280.4]
  wire [22:0] _T_256; // @[Modules.scala 137:32:@39280.4]
  wire [7:0] _GEN_49; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_12; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_50; // @[Modules.scala 139:37:@39282.4]
  wire [22:0] _T_258; // @[Modules.scala 139:37:@39282.4]
  wire [7:0] _GEN_51; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_12; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_260; // @[Modules.scala 140:38:@39284.4]
  wire [7:0] _T_261; // @[Modules.scala 140:38:@39285.4]
  wire [7:0] _T_262; // @[Modules.scala 140:38:@39286.4]
  wire [8:0] _T_264; // @[Modules.scala 132:28:@39288.4]
  wire [7:0] _T_265; // @[Modules.scala 132:28:@39289.4]
  wire [7:0] c_x_13; // @[Modules.scala 132:28:@39290.4]
  wire [22:0] _GEN_52; // @[Modules.scala 137:32:@39292.4]
  wire [22:0] _T_268; // @[Modules.scala 137:32:@39292.4]
  wire [7:0] _GEN_53; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_13; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_54; // @[Modules.scala 139:37:@39294.4]
  wire [22:0] _T_270; // @[Modules.scala 139:37:@39294.4]
  wire [7:0] _GEN_55; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_13; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_272; // @[Modules.scala 140:38:@39296.4]
  wire [7:0] _T_273; // @[Modules.scala 140:38:@39297.4]
  wire [7:0] _T_274; // @[Modules.scala 140:38:@39298.4]
  wire [8:0] _T_276; // @[Modules.scala 132:28:@39300.4]
  wire [7:0] _T_277; // @[Modules.scala 132:28:@39301.4]
  wire [7:0] c_x_14; // @[Modules.scala 132:28:@39302.4]
  wire [22:0] _GEN_56; // @[Modules.scala 137:32:@39304.4]
  wire [22:0] _T_280; // @[Modules.scala 137:32:@39304.4]
  wire [7:0] _GEN_57; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_14; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_58; // @[Modules.scala 139:37:@39306.4]
  wire [22:0] _T_282; // @[Modules.scala 139:37:@39306.4]
  wire [7:0] _GEN_59; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_14; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_284; // @[Modules.scala 140:38:@39308.4]
  wire [7:0] _T_285; // @[Modules.scala 140:38:@39309.4]
  wire [7:0] _T_286; // @[Modules.scala 140:38:@39310.4]
  wire [8:0] _T_288; // @[Modules.scala 132:28:@39312.4]
  wire [7:0] _T_289; // @[Modules.scala 132:28:@39313.4]
  wire [7:0] c_x_15; // @[Modules.scala 132:28:@39314.4]
  wire [22:0] _GEN_60; // @[Modules.scala 137:32:@39316.4]
  wire [22:0] _T_292; // @[Modules.scala 137:32:@39316.4]
  wire [7:0] _GEN_61; // @[Modules.scala 129:21:@39130.4]
  wire [7:0] x_hat_15; // @[Modules.scala 129:21:@39130.4]
  wire [22:0] _GEN_62; // @[Modules.scala 139:37:@39318.4]
  wire [22:0] _T_294; // @[Modules.scala 139:37:@39318.4]
  wire [7:0] _GEN_63; // @[Modules.scala 130:28:@39131.4]
  wire [7:0] normed_x_hat_15; // @[Modules.scala 130:28:@39131.4]
  wire [8:0] _T_296; // @[Modules.scala 140:38:@39320.4]
  wire [7:0] _T_297; // @[Modules.scala 140:38:@39321.4]
  wire [7:0] _T_298; // @[Modules.scala 140:38:@39322.4]
  assign _T_108 = $signed(io_in_0) - $signed(8'sh0); // @[Modules.scala 132:28:@39132.4]
  assign _T_109 = _T_108[7:0]; // @[Modules.scala 132:28:@39133.4]
  assign c_x_0 = $signed(_T_109); // @[Modules.scala 132:28:@39134.4]
  assign _GEN_0 = {{15{c_x_0[7]}},c_x_0}; // @[Modules.scala 137:32:@39136.4]
  assign _T_112 = $signed(_GEN_0) << 4'h2; // @[Modules.scala 137:32:@39136.4]
  assign _GEN_1 = _T_112[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_0 = $signed(_GEN_1); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_2 = {{15{x_hat_0[7]}},x_hat_0}; // @[Modules.scala 139:37:@39138.4]
  assign _T_114 = $signed(_GEN_2) << 4'h1; // @[Modules.scala 139:37:@39138.4]
  assign _GEN_3 = _T_114[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_0 = $signed(_GEN_3); // @[Modules.scala 130:28:@39131.4]
  assign _T_116 = $signed(normed_x_hat_0) + $signed(8'sh0); // @[Modules.scala 140:38:@39140.4]
  assign _T_117 = _T_116[7:0]; // @[Modules.scala 140:38:@39141.4]
  assign _T_118 = $signed(_T_117); // @[Modules.scala 140:38:@39142.4]
  assign _T_120 = $signed(io_in_1) - $signed(-8'sh1); // @[Modules.scala 132:28:@39144.4]
  assign _T_121 = _T_120[7:0]; // @[Modules.scala 132:28:@39145.4]
  assign c_x_1 = $signed(_T_121); // @[Modules.scala 132:28:@39146.4]
  assign _GEN_4 = {{15{c_x_1[7]}},c_x_1}; // @[Modules.scala 137:32:@39148.4]
  assign _T_124 = $signed(_GEN_4) << 4'h3; // @[Modules.scala 137:32:@39148.4]
  assign _GEN_5 = _T_124[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_1 = $signed(_GEN_5); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_6 = {{15{x_hat_1[7]}},x_hat_1}; // @[Modules.scala 139:37:@39150.4]
  assign _T_126 = $signed(_GEN_6) << 4'h1; // @[Modules.scala 139:37:@39150.4]
  assign _GEN_7 = _T_126[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_1 = $signed(_GEN_7); // @[Modules.scala 130:28:@39131.4]
  assign _T_128 = $signed(normed_x_hat_1) + $signed(8'sh0); // @[Modules.scala 140:38:@39152.4]
  assign _T_129 = _T_128[7:0]; // @[Modules.scala 140:38:@39153.4]
  assign _T_130 = $signed(_T_129); // @[Modules.scala 140:38:@39154.4]
  assign _T_132 = $signed(io_in_2) - $signed(8'sh0); // @[Modules.scala 132:28:@39156.4]
  assign _T_133 = _T_132[7:0]; // @[Modules.scala 132:28:@39157.4]
  assign c_x_2 = $signed(_T_133); // @[Modules.scala 132:28:@39158.4]
  assign _GEN_8 = {{15{c_x_2[7]}},c_x_2}; // @[Modules.scala 137:32:@39160.4]
  assign _T_136 = $signed(_GEN_8) << 4'h3; // @[Modules.scala 137:32:@39160.4]
  assign _GEN_9 = _T_136[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_2 = $signed(_GEN_9); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_10 = {{15{x_hat_2[7]}},x_hat_2}; // @[Modules.scala 139:37:@39162.4]
  assign _T_138 = $signed(_GEN_10) << 4'h1; // @[Modules.scala 139:37:@39162.4]
  assign _GEN_11 = _T_138[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_2 = $signed(_GEN_11); // @[Modules.scala 130:28:@39131.4]
  assign _T_140 = $signed(normed_x_hat_2) + $signed(8'sh0); // @[Modules.scala 140:38:@39164.4]
  assign _T_141 = _T_140[7:0]; // @[Modules.scala 140:38:@39165.4]
  assign _T_142 = $signed(_T_141); // @[Modules.scala 140:38:@39166.4]
  assign _T_144 = $signed(io_in_3) - $signed(8'sh1); // @[Modules.scala 132:28:@39168.4]
  assign _T_145 = _T_144[7:0]; // @[Modules.scala 132:28:@39169.4]
  assign c_x_3 = $signed(_T_145); // @[Modules.scala 132:28:@39170.4]
  assign _GEN_12 = {{15{c_x_3[7]}},c_x_3}; // @[Modules.scala 137:32:@39172.4]
  assign _T_148 = $signed(_GEN_12) << 4'h2; // @[Modules.scala 137:32:@39172.4]
  assign _GEN_13 = _T_148[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_3 = $signed(_GEN_13); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_14 = {{15{x_hat_3[7]}},x_hat_3}; // @[Modules.scala 139:37:@39174.4]
  assign _T_150 = $signed(_GEN_14) << 4'h1; // @[Modules.scala 139:37:@39174.4]
  assign _GEN_15 = _T_150[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_3 = $signed(_GEN_15); // @[Modules.scala 130:28:@39131.4]
  assign _T_152 = $signed(normed_x_hat_3) + $signed(8'sh0); // @[Modules.scala 140:38:@39176.4]
  assign _T_153 = _T_152[7:0]; // @[Modules.scala 140:38:@39177.4]
  assign _T_154 = $signed(_T_153); // @[Modules.scala 140:38:@39178.4]
  assign _T_156 = $signed(io_in_4) - $signed(-8'sh1); // @[Modules.scala 132:28:@39180.4]
  assign _T_157 = _T_156[7:0]; // @[Modules.scala 132:28:@39181.4]
  assign c_x_4 = $signed(_T_157); // @[Modules.scala 132:28:@39182.4]
  assign _GEN_16 = {{15{c_x_4[7]}},c_x_4}; // @[Modules.scala 137:32:@39184.4]
  assign _T_160 = $signed(_GEN_16) << 4'h2; // @[Modules.scala 137:32:@39184.4]
  assign _GEN_17 = _T_160[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_4 = $signed(_GEN_17); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_18 = {{15{x_hat_4[7]}},x_hat_4}; // @[Modules.scala 139:37:@39186.4]
  assign _T_162 = $signed(_GEN_18) << 4'h1; // @[Modules.scala 139:37:@39186.4]
  assign _GEN_19 = _T_162[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_4 = $signed(_GEN_19); // @[Modules.scala 130:28:@39131.4]
  assign _T_164 = $signed(normed_x_hat_4) + $signed(8'sh0); // @[Modules.scala 140:38:@39188.4]
  assign _T_165 = _T_164[7:0]; // @[Modules.scala 140:38:@39189.4]
  assign _T_166 = $signed(_T_165); // @[Modules.scala 140:38:@39190.4]
  assign _T_168 = $signed(io_in_5) - $signed(8'sh1); // @[Modules.scala 132:28:@39192.4]
  assign _T_169 = _T_168[7:0]; // @[Modules.scala 132:28:@39193.4]
  assign c_x_5 = $signed(_T_169); // @[Modules.scala 132:28:@39194.4]
  assign _GEN_20 = {{15{c_x_5[7]}},c_x_5}; // @[Modules.scala 137:32:@39196.4]
  assign _T_172 = $signed(_GEN_20) << 4'h2; // @[Modules.scala 137:32:@39196.4]
  assign _GEN_21 = _T_172[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_5 = $signed(_GEN_21); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_22 = {{15{x_hat_5[7]}},x_hat_5}; // @[Modules.scala 139:37:@39198.4]
  assign _T_174 = $signed(_GEN_22) << 4'h1; // @[Modules.scala 139:37:@39198.4]
  assign _GEN_23 = _T_174[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_5 = $signed(_GEN_23); // @[Modules.scala 130:28:@39131.4]
  assign _T_176 = $signed(normed_x_hat_5) + $signed(8'sh0); // @[Modules.scala 140:38:@39200.4]
  assign _T_177 = _T_176[7:0]; // @[Modules.scala 140:38:@39201.4]
  assign _T_178 = $signed(_T_177); // @[Modules.scala 140:38:@39202.4]
  assign _T_180 = $signed(io_in_6) - $signed(8'sh0); // @[Modules.scala 132:28:@39204.4]
  assign _T_181 = _T_180[7:0]; // @[Modules.scala 132:28:@39205.4]
  assign c_x_6 = $signed(_T_181); // @[Modules.scala 132:28:@39206.4]
  assign _GEN_24 = {{15{c_x_6[7]}},c_x_6}; // @[Modules.scala 137:32:@39208.4]
  assign _T_184 = $signed(_GEN_24) << 4'h2; // @[Modules.scala 137:32:@39208.4]
  assign _GEN_25 = _T_184[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_6 = $signed(_GEN_25); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_26 = {{15{x_hat_6[7]}},x_hat_6}; // @[Modules.scala 139:37:@39210.4]
  assign _T_186 = $signed(_GEN_26) << 4'h1; // @[Modules.scala 139:37:@39210.4]
  assign _GEN_27 = _T_186[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_6 = $signed(_GEN_27); // @[Modules.scala 130:28:@39131.4]
  assign _T_188 = $signed(normed_x_hat_6) + $signed(8'sh0); // @[Modules.scala 140:38:@39212.4]
  assign _T_189 = _T_188[7:0]; // @[Modules.scala 140:38:@39213.4]
  assign _T_190 = $signed(_T_189); // @[Modules.scala 140:38:@39214.4]
  assign _T_192 = $signed(io_in_7) - $signed(-8'sh1); // @[Modules.scala 132:28:@39216.4]
  assign _T_193 = _T_192[7:0]; // @[Modules.scala 132:28:@39217.4]
  assign c_x_7 = $signed(_T_193); // @[Modules.scala 132:28:@39218.4]
  assign _GEN_28 = {{15{c_x_7[7]}},c_x_7}; // @[Modules.scala 137:32:@39220.4]
  assign _T_196 = $signed(_GEN_28) << 4'h2; // @[Modules.scala 137:32:@39220.4]
  assign _GEN_29 = _T_196[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_7 = $signed(_GEN_29); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_30 = {{15{x_hat_7[7]}},x_hat_7}; // @[Modules.scala 139:37:@39222.4]
  assign _T_198 = $signed(_GEN_30) << 4'h1; // @[Modules.scala 139:37:@39222.4]
  assign _GEN_31 = _T_198[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_7 = $signed(_GEN_31); // @[Modules.scala 130:28:@39131.4]
  assign _T_200 = $signed(normed_x_hat_7) + $signed(8'sh0); // @[Modules.scala 140:38:@39224.4]
  assign _T_201 = _T_200[7:0]; // @[Modules.scala 140:38:@39225.4]
  assign _T_202 = $signed(_T_201); // @[Modules.scala 140:38:@39226.4]
  assign _T_204 = $signed(io_in_8) - $signed(-8'sh1); // @[Modules.scala 132:28:@39228.4]
  assign _T_205 = _T_204[7:0]; // @[Modules.scala 132:28:@39229.4]
  assign c_x_8 = $signed(_T_205); // @[Modules.scala 132:28:@39230.4]
  assign _GEN_32 = {{15{c_x_8[7]}},c_x_8}; // @[Modules.scala 137:32:@39232.4]
  assign _T_208 = $signed(_GEN_32) << 4'h2; // @[Modules.scala 137:32:@39232.4]
  assign _GEN_33 = _T_208[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_8 = $signed(_GEN_33); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_34 = {{15{x_hat_8[7]}},x_hat_8}; // @[Modules.scala 139:37:@39234.4]
  assign _T_210 = $signed(_GEN_34) << 4'h1; // @[Modules.scala 139:37:@39234.4]
  assign _GEN_35 = _T_210[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_8 = $signed(_GEN_35); // @[Modules.scala 130:28:@39131.4]
  assign _T_212 = $signed(normed_x_hat_8) + $signed(8'sh0); // @[Modules.scala 140:38:@39236.4]
  assign _T_213 = _T_212[7:0]; // @[Modules.scala 140:38:@39237.4]
  assign _T_214 = $signed(_T_213); // @[Modules.scala 140:38:@39238.4]
  assign _T_216 = $signed(io_in_9) - $signed(8'sh0); // @[Modules.scala 132:28:@39240.4]
  assign _T_217 = _T_216[7:0]; // @[Modules.scala 132:28:@39241.4]
  assign c_x_9 = $signed(_T_217); // @[Modules.scala 132:28:@39242.4]
  assign _GEN_36 = {{15{c_x_9[7]}},c_x_9}; // @[Modules.scala 137:32:@39244.4]
  assign _T_220 = $signed(_GEN_36) << 4'h2; // @[Modules.scala 137:32:@39244.4]
  assign _GEN_37 = _T_220[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_9 = $signed(_GEN_37); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_38 = {{15{x_hat_9[7]}},x_hat_9}; // @[Modules.scala 139:37:@39246.4]
  assign _T_222 = $signed(_GEN_38) << 4'h1; // @[Modules.scala 139:37:@39246.4]
  assign _GEN_39 = _T_222[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_9 = $signed(_GEN_39); // @[Modules.scala 130:28:@39131.4]
  assign _T_224 = $signed(normed_x_hat_9) + $signed(8'sh0); // @[Modules.scala 140:38:@39248.4]
  assign _T_225 = _T_224[7:0]; // @[Modules.scala 140:38:@39249.4]
  assign _T_226 = $signed(_T_225); // @[Modules.scala 140:38:@39250.4]
  assign _T_228 = $signed(io_in_10) - $signed(-8'sh1); // @[Modules.scala 132:28:@39252.4]
  assign _T_229 = _T_228[7:0]; // @[Modules.scala 132:28:@39253.4]
  assign c_x_10 = $signed(_T_229); // @[Modules.scala 132:28:@39254.4]
  assign _GEN_40 = {{15{c_x_10[7]}},c_x_10}; // @[Modules.scala 137:32:@39256.4]
  assign _T_232 = $signed(_GEN_40) << 4'h2; // @[Modules.scala 137:32:@39256.4]
  assign _GEN_41 = _T_232[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_10 = $signed(_GEN_41); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_42 = {{15{x_hat_10[7]}},x_hat_10}; // @[Modules.scala 139:37:@39258.4]
  assign _T_234 = $signed(_GEN_42) << 4'h0; // @[Modules.scala 139:37:@39258.4]
  assign _GEN_43 = _T_234[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_10 = $signed(_GEN_43); // @[Modules.scala 130:28:@39131.4]
  assign _T_236 = $signed(normed_x_hat_10) + $signed(8'sh0); // @[Modules.scala 140:38:@39260.4]
  assign _T_237 = _T_236[7:0]; // @[Modules.scala 140:38:@39261.4]
  assign _T_238 = $signed(_T_237); // @[Modules.scala 140:38:@39262.4]
  assign _T_240 = $signed(io_in_11) - $signed(8'sh0); // @[Modules.scala 132:28:@39264.4]
  assign _T_241 = _T_240[7:0]; // @[Modules.scala 132:28:@39265.4]
  assign c_x_11 = $signed(_T_241); // @[Modules.scala 132:28:@39266.4]
  assign _GEN_44 = {{15{c_x_11[7]}},c_x_11}; // @[Modules.scala 137:32:@39268.4]
  assign _T_244 = $signed(_GEN_44) << 4'h2; // @[Modules.scala 137:32:@39268.4]
  assign _GEN_45 = _T_244[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_11 = $signed(_GEN_45); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_46 = {{15{x_hat_11[7]}},x_hat_11}; // @[Modules.scala 139:37:@39270.4]
  assign _T_246 = $signed(_GEN_46) << 4'h1; // @[Modules.scala 139:37:@39270.4]
  assign _GEN_47 = _T_246[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_11 = $signed(_GEN_47); // @[Modules.scala 130:28:@39131.4]
  assign _T_248 = $signed(normed_x_hat_11) + $signed(8'sh0); // @[Modules.scala 140:38:@39272.4]
  assign _T_249 = _T_248[7:0]; // @[Modules.scala 140:38:@39273.4]
  assign _T_250 = $signed(_T_249); // @[Modules.scala 140:38:@39274.4]
  assign _T_252 = $signed(io_in_12) - $signed(8'sh0); // @[Modules.scala 132:28:@39276.4]
  assign _T_253 = _T_252[7:0]; // @[Modules.scala 132:28:@39277.4]
  assign c_x_12 = $signed(_T_253); // @[Modules.scala 132:28:@39278.4]
  assign _GEN_48 = {{15{c_x_12[7]}},c_x_12}; // @[Modules.scala 137:32:@39280.4]
  assign _T_256 = $signed(_GEN_48) << 4'h3; // @[Modules.scala 137:32:@39280.4]
  assign _GEN_49 = _T_256[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_12 = $signed(_GEN_49); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_50 = {{15{x_hat_12[7]}},x_hat_12}; // @[Modules.scala 139:37:@39282.4]
  assign _T_258 = $signed(_GEN_50) << 4'h1; // @[Modules.scala 139:37:@39282.4]
  assign _GEN_51 = _T_258[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_12 = $signed(_GEN_51); // @[Modules.scala 130:28:@39131.4]
  assign _T_260 = $signed(normed_x_hat_12) + $signed(8'sh1); // @[Modules.scala 140:38:@39284.4]
  assign _T_261 = _T_260[7:0]; // @[Modules.scala 140:38:@39285.4]
  assign _T_262 = $signed(_T_261); // @[Modules.scala 140:38:@39286.4]
  assign _T_264 = $signed(io_in_13) - $signed(8'sh0); // @[Modules.scala 132:28:@39288.4]
  assign _T_265 = _T_264[7:0]; // @[Modules.scala 132:28:@39289.4]
  assign c_x_13 = $signed(_T_265); // @[Modules.scala 132:28:@39290.4]
  assign _GEN_52 = {{15{c_x_13[7]}},c_x_13}; // @[Modules.scala 137:32:@39292.4]
  assign _T_268 = $signed(_GEN_52) << 4'h2; // @[Modules.scala 137:32:@39292.4]
  assign _GEN_53 = _T_268[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_13 = $signed(_GEN_53); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_54 = {{15{x_hat_13[7]}},x_hat_13}; // @[Modules.scala 139:37:@39294.4]
  assign _T_270 = $signed(_GEN_54) << 4'h1; // @[Modules.scala 139:37:@39294.4]
  assign _GEN_55 = _T_270[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_13 = $signed(_GEN_55); // @[Modules.scala 130:28:@39131.4]
  assign _T_272 = $signed(normed_x_hat_13) + $signed(8'sh0); // @[Modules.scala 140:38:@39296.4]
  assign _T_273 = _T_272[7:0]; // @[Modules.scala 140:38:@39297.4]
  assign _T_274 = $signed(_T_273); // @[Modules.scala 140:38:@39298.4]
  assign _T_276 = $signed(io_in_14) - $signed(8'sh1); // @[Modules.scala 132:28:@39300.4]
  assign _T_277 = _T_276[7:0]; // @[Modules.scala 132:28:@39301.4]
  assign c_x_14 = $signed(_T_277); // @[Modules.scala 132:28:@39302.4]
  assign _GEN_56 = {{15{c_x_14[7]}},c_x_14}; // @[Modules.scala 137:32:@39304.4]
  assign _T_280 = $signed(_GEN_56) << 4'h2; // @[Modules.scala 137:32:@39304.4]
  assign _GEN_57 = _T_280[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_14 = $signed(_GEN_57); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_58 = {{15{x_hat_14[7]}},x_hat_14}; // @[Modules.scala 139:37:@39306.4]
  assign _T_282 = $signed(_GEN_58) << 4'h1; // @[Modules.scala 139:37:@39306.4]
  assign _GEN_59 = _T_282[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_14 = $signed(_GEN_59); // @[Modules.scala 130:28:@39131.4]
  assign _T_284 = $signed(normed_x_hat_14) + $signed(8'sh0); // @[Modules.scala 140:38:@39308.4]
  assign _T_285 = _T_284[7:0]; // @[Modules.scala 140:38:@39309.4]
  assign _T_286 = $signed(_T_285); // @[Modules.scala 140:38:@39310.4]
  assign _T_288 = $signed(io_in_15) - $signed(-8'sh1); // @[Modules.scala 132:28:@39312.4]
  assign _T_289 = _T_288[7:0]; // @[Modules.scala 132:28:@39313.4]
  assign c_x_15 = $signed(_T_289); // @[Modules.scala 132:28:@39314.4]
  assign _GEN_60 = {{15{c_x_15[7]}},c_x_15}; // @[Modules.scala 137:32:@39316.4]
  assign _T_292 = $signed(_GEN_60) << 4'h3; // @[Modules.scala 137:32:@39316.4]
  assign _GEN_61 = _T_292[7:0]; // @[Modules.scala 129:21:@39130.4]
  assign x_hat_15 = $signed(_GEN_61); // @[Modules.scala 129:21:@39130.4]
  assign _GEN_62 = {{15{x_hat_15[7]}},x_hat_15}; // @[Modules.scala 139:37:@39318.4]
  assign _T_294 = $signed(_GEN_62) << 4'h1; // @[Modules.scala 139:37:@39318.4]
  assign _GEN_63 = _T_294[7:0]; // @[Modules.scala 130:28:@39131.4]
  assign normed_x_hat_15 = $signed(_GEN_63); // @[Modules.scala 130:28:@39131.4]
  assign _T_296 = $signed(normed_x_hat_15) + $signed(8'sh0); // @[Modules.scala 140:38:@39320.4]
  assign _T_297 = _T_296[7:0]; // @[Modules.scala 140:38:@39321.4]
  assign _T_298 = $signed(_T_297); // @[Modules.scala 140:38:@39322.4]
  assign io_out_0 = _T_118;
  assign io_out_1 = _T_130;
  assign io_out_2 = _T_142;
  assign io_out_3 = _T_154;
  assign io_out_4 = _T_166;
  assign io_out_5 = _T_178;
  assign io_out_6 = _T_190;
  assign io_out_7 = _T_202;
  assign io_out_8 = _T_214;
  assign io_out_9 = _T_226;
  assign io_out_10 = _T_238;
  assign io_out_11 = _T_250;
  assign io_out_12 = _T_262;
  assign io_out_13 = _T_274;
  assign io_out_14 = _T_286;
  assign io_out_15 = _T_298;
endmodule
module Binarize_1( // @[:@39325.2]
  input  [7:0] io_in_0, // @[:@39328.4]
  input  [7:0] io_in_1, // @[:@39328.4]
  input  [7:0] io_in_2, // @[:@39328.4]
  input  [7:0] io_in_3, // @[:@39328.4]
  input  [7:0] io_in_4, // @[:@39328.4]
  input  [7:0] io_in_5, // @[:@39328.4]
  input  [7:0] io_in_6, // @[:@39328.4]
  input  [7:0] io_in_7, // @[:@39328.4]
  input  [7:0] io_in_8, // @[:@39328.4]
  input  [7:0] io_in_9, // @[:@39328.4]
  input  [7:0] io_in_10, // @[:@39328.4]
  input  [7:0] io_in_11, // @[:@39328.4]
  input  [7:0] io_in_12, // @[:@39328.4]
  input  [7:0] io_in_13, // @[:@39328.4]
  input  [7:0] io_in_14, // @[:@39328.4]
  input  [7:0] io_in_15, // @[:@39328.4]
  output [1:0] io_out_0, // @[:@39328.4]
  output [1:0] io_out_1, // @[:@39328.4]
  output [1:0] io_out_2, // @[:@39328.4]
  output [1:0] io_out_3, // @[:@39328.4]
  output [1:0] io_out_4, // @[:@39328.4]
  output [1:0] io_out_5, // @[:@39328.4]
  output [1:0] io_out_6, // @[:@39328.4]
  output [1:0] io_out_7, // @[:@39328.4]
  output [1:0] io_out_8, // @[:@39328.4]
  output [1:0] io_out_9, // @[:@39328.4]
  output [1:0] io_out_10, // @[:@39328.4]
  output [1:0] io_out_11, // @[:@39328.4]
  output [1:0] io_out_12, // @[:@39328.4]
  output [1:0] io_out_13, // @[:@39328.4]
  output [1:0] io_out_14, // @[:@39328.4]
  output [1:0] io_out_15 // @[:@39328.4]
);
  wire  _T_45; // @[Modules.scala 151:24:@39330.4]
  wire [1:0] _GEN_0; // @[Modules.scala 151:32:@39331.4]
  wire  _T_49; // @[Modules.scala 151:24:@39337.4]
  wire [1:0] _GEN_1; // @[Modules.scala 151:32:@39338.4]
  wire  _T_53; // @[Modules.scala 151:24:@39344.4]
  wire [1:0] _GEN_2; // @[Modules.scala 151:32:@39345.4]
  wire  _T_57; // @[Modules.scala 151:24:@39351.4]
  wire [1:0] _GEN_3; // @[Modules.scala 151:32:@39352.4]
  wire  _T_61; // @[Modules.scala 151:24:@39358.4]
  wire [1:0] _GEN_4; // @[Modules.scala 151:32:@39359.4]
  wire  _T_65; // @[Modules.scala 151:24:@39365.4]
  wire [1:0] _GEN_5; // @[Modules.scala 151:32:@39366.4]
  wire  _T_69; // @[Modules.scala 151:24:@39372.4]
  wire [1:0] _GEN_6; // @[Modules.scala 151:32:@39373.4]
  wire  _T_73; // @[Modules.scala 151:24:@39379.4]
  wire [1:0] _GEN_7; // @[Modules.scala 151:32:@39380.4]
  wire  _T_77; // @[Modules.scala 151:24:@39386.4]
  wire [1:0] _GEN_8; // @[Modules.scala 151:32:@39387.4]
  wire  _T_81; // @[Modules.scala 151:24:@39393.4]
  wire [1:0] _GEN_9; // @[Modules.scala 151:32:@39394.4]
  wire  _T_85; // @[Modules.scala 151:24:@39400.4]
  wire [1:0] _GEN_10; // @[Modules.scala 151:32:@39401.4]
  wire  _T_89; // @[Modules.scala 151:24:@39407.4]
  wire [1:0] _GEN_11; // @[Modules.scala 151:32:@39408.4]
  wire  _T_93; // @[Modules.scala 151:24:@39414.4]
  wire [1:0] _GEN_12; // @[Modules.scala 151:32:@39415.4]
  wire  _T_97; // @[Modules.scala 151:24:@39421.4]
  wire [1:0] _GEN_13; // @[Modules.scala 151:32:@39422.4]
  wire  _T_101; // @[Modules.scala 151:24:@39428.4]
  wire [1:0] _GEN_14; // @[Modules.scala 151:32:@39429.4]
  wire  _T_105; // @[Modules.scala 151:24:@39435.4]
  wire [1:0] _GEN_15; // @[Modules.scala 151:32:@39436.4]
  assign _T_45 = $signed(io_in_0) >= $signed(8'sh0); // @[Modules.scala 151:24:@39330.4]
  assign _GEN_0 = _T_45 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39331.4]
  assign _T_49 = $signed(io_in_1) >= $signed(8'sh0); // @[Modules.scala 151:24:@39337.4]
  assign _GEN_1 = _T_49 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39338.4]
  assign _T_53 = $signed(io_in_2) >= $signed(8'sh0); // @[Modules.scala 151:24:@39344.4]
  assign _GEN_2 = _T_53 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39345.4]
  assign _T_57 = $signed(io_in_3) >= $signed(8'sh0); // @[Modules.scala 151:24:@39351.4]
  assign _GEN_3 = _T_57 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39352.4]
  assign _T_61 = $signed(io_in_4) >= $signed(8'sh0); // @[Modules.scala 151:24:@39358.4]
  assign _GEN_4 = _T_61 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39359.4]
  assign _T_65 = $signed(io_in_5) >= $signed(8'sh0); // @[Modules.scala 151:24:@39365.4]
  assign _GEN_5 = _T_65 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39366.4]
  assign _T_69 = $signed(io_in_6) >= $signed(8'sh0); // @[Modules.scala 151:24:@39372.4]
  assign _GEN_6 = _T_69 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39373.4]
  assign _T_73 = $signed(io_in_7) >= $signed(8'sh0); // @[Modules.scala 151:24:@39379.4]
  assign _GEN_7 = _T_73 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39380.4]
  assign _T_77 = $signed(io_in_8) >= $signed(8'sh0); // @[Modules.scala 151:24:@39386.4]
  assign _GEN_8 = _T_77 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39387.4]
  assign _T_81 = $signed(io_in_9) >= $signed(8'sh0); // @[Modules.scala 151:24:@39393.4]
  assign _GEN_9 = _T_81 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39394.4]
  assign _T_85 = $signed(io_in_10) >= $signed(8'sh0); // @[Modules.scala 151:24:@39400.4]
  assign _GEN_10 = _T_85 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39401.4]
  assign _T_89 = $signed(io_in_11) >= $signed(8'sh0); // @[Modules.scala 151:24:@39407.4]
  assign _GEN_11 = _T_89 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39408.4]
  assign _T_93 = $signed(io_in_12) >= $signed(8'sh0); // @[Modules.scala 151:24:@39414.4]
  assign _GEN_12 = _T_93 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39415.4]
  assign _T_97 = $signed(io_in_13) >= $signed(8'sh0); // @[Modules.scala 151:24:@39421.4]
  assign _GEN_13 = _T_97 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39422.4]
  assign _T_101 = $signed(io_in_14) >= $signed(8'sh0); // @[Modules.scala 151:24:@39428.4]
  assign _GEN_14 = _T_101 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39429.4]
  assign _T_105 = $signed(io_in_15) >= $signed(8'sh0); // @[Modules.scala 151:24:@39435.4]
  assign _GEN_15 = _T_105 ? $signed(2'sh1) : $signed(-2'sh1); // @[Modules.scala 151:32:@39436.4]
  assign io_out_0 = _GEN_0;
  assign io_out_1 = _GEN_1;
  assign io_out_2 = _GEN_2;
  assign io_out_3 = _GEN_3;
  assign io_out_4 = _GEN_4;
  assign io_out_5 = _GEN_5;
  assign io_out_6 = _GEN_6;
  assign io_out_7 = _GEN_7;
  assign io_out_8 = _GEN_8;
  assign io_out_9 = _GEN_9;
  assign io_out_10 = _GEN_10;
  assign io_out_11 = _GEN_11;
  assign io_out_12 = _GEN_12;
  assign io_out_13 = _GEN_13;
  assign io_out_14 = _GEN_14;
  assign io_out_15 = _GEN_15;
endmodule
module Linear_1( // @[:@39443.2]
  input  [1:0] io_in_0, // @[:@39446.4]
  input  [1:0] io_in_1, // @[:@39446.4]
  input  [1:0] io_in_2, // @[:@39446.4]
  input  [1:0] io_in_3, // @[:@39446.4]
  input  [1:0] io_in_4, // @[:@39446.4]
  input  [1:0] io_in_5, // @[:@39446.4]
  input  [1:0] io_in_6, // @[:@39446.4]
  input  [1:0] io_in_7, // @[:@39446.4]
  input  [1:0] io_in_8, // @[:@39446.4]
  input  [1:0] io_in_9, // @[:@39446.4]
  input  [1:0] io_in_10, // @[:@39446.4]
  input  [1:0] io_in_11, // @[:@39446.4]
  input  [1:0] io_in_12, // @[:@39446.4]
  input  [1:0] io_in_13, // @[:@39446.4]
  input  [1:0] io_in_14, // @[:@39446.4]
  input  [1:0] io_in_15, // @[:@39446.4]
  output [7:0] io_out_0, // @[:@39446.4]
  output [7:0] io_out_1, // @[:@39446.4]
  output [7:0] io_out_2, // @[:@39446.4]
  output [7:0] io_out_3, // @[:@39446.4]
  output [7:0] io_out_4, // @[:@39446.4]
  output [7:0] io_out_5, // @[:@39446.4]
  output [7:0] io_out_6, // @[:@39446.4]
  output [7:0] io_out_7, // @[:@39446.4]
  output [7:0] io_out_8, // @[:@39446.4]
  output [7:0] io_out_9 // @[:@39446.4]
);
  wire [7:0] _GEN_0; // @[Modules.scala 108:54:@39450.4]
  wire [8:0] _T_837; // @[Modules.scala 108:54:@39450.4]
  wire [7:0] _T_838; // @[Modules.scala 108:54:@39451.4]
  wire [7:0] buffer_0_1; // @[Modules.scala 108:54:@39452.4]
  wire [7:0] _GEN_1; // @[Modules.scala 108:54:@39461.4]
  wire [8:0] _T_840; // @[Modules.scala 108:54:@39461.4]
  wire [7:0] _T_841; // @[Modules.scala 108:54:@39462.4]
  wire [7:0] buffer_0_9; // @[Modules.scala 108:54:@39463.4]
  wire [7:0] _GEN_2; // @[Modules.scala 108:54:@39465.4]
  wire [8:0] _T_843; // @[Modules.scala 108:54:@39465.4]
  wire [7:0] _T_844; // @[Modules.scala 108:54:@39466.4]
  wire [7:0] buffer_0_10; // @[Modules.scala 108:54:@39467.4]
  wire [7:0] _GEN_3; // @[Modules.scala 108:54:@39469.4]
  wire [8:0] _T_846; // @[Modules.scala 108:54:@39469.4]
  wire [7:0] _T_847; // @[Modules.scala 108:54:@39470.4]
  wire [7:0] buffer_0_11; // @[Modules.scala 108:54:@39471.4]
  wire [7:0] _GEN_4; // @[Modules.scala 108:54:@39473.4]
  wire [8:0] _T_849; // @[Modules.scala 108:54:@39473.4]
  wire [7:0] _T_850; // @[Modules.scala 108:54:@39474.4]
  wire [7:0] buffer_0_12; // @[Modules.scala 108:54:@39475.4]
  wire [7:0] _GEN_5; // @[Modules.scala 108:54:@39477.4]
  wire [8:0] _T_852; // @[Modules.scala 108:54:@39477.4]
  wire [7:0] _T_853; // @[Modules.scala 108:54:@39478.4]
  wire [7:0] buffer_0_13; // @[Modules.scala 108:54:@39479.4]
  wire [7:0] _GEN_6; // @[Modules.scala 108:54:@39482.4]
  wire [8:0] _T_855; // @[Modules.scala 108:54:@39482.4]
  wire [7:0] _T_856; // @[Modules.scala 108:54:@39483.4]
  wire [7:0] buffer_0_15; // @[Modules.scala 108:54:@39484.4]
  wire [7:0] buffer_1_0; // @[Modules.scala 91:22:@39448.4]
  wire [7:0] _GEN_7; // @[Modules.scala 108:54:@39489.4]
  wire [8:0] _T_858; // @[Modules.scala 108:54:@39489.4]
  wire [7:0] _T_859; // @[Modules.scala 108:54:@39490.4]
  wire [7:0] buffer_1_2; // @[Modules.scala 108:54:@39491.4]
  wire [7:0] _GEN_8; // @[Modules.scala 108:54:@39493.4]
  wire [8:0] _T_861; // @[Modules.scala 108:54:@39493.4]
  wire [7:0] _T_862; // @[Modules.scala 108:54:@39494.4]
  wire [7:0] buffer_1_3; // @[Modules.scala 108:54:@39495.4]
  wire [7:0] _GEN_9; // @[Modules.scala 108:54:@39497.4]
  wire [8:0] _T_864; // @[Modules.scala 108:54:@39497.4]
  wire [7:0] _T_865; // @[Modules.scala 108:54:@39498.4]
  wire [7:0] buffer_1_4; // @[Modules.scala 108:54:@39499.4]
  wire [7:0] _GEN_10; // @[Modules.scala 108:54:@39501.4]
  wire [8:0] _T_867; // @[Modules.scala 108:54:@39501.4]
  wire [7:0] _T_868; // @[Modules.scala 108:54:@39502.4]
  wire [7:0] buffer_1_5; // @[Modules.scala 108:54:@39503.4]
  wire [7:0] _GEN_11; // @[Modules.scala 108:54:@39505.4]
  wire [8:0] _T_870; // @[Modules.scala 108:54:@39505.4]
  wire [7:0] _T_871; // @[Modules.scala 108:54:@39506.4]
  wire [7:0] buffer_1_6; // @[Modules.scala 108:54:@39507.4]
  wire [7:0] _GEN_12; // @[Modules.scala 108:54:@39509.4]
  wire [8:0] _T_873; // @[Modules.scala 108:54:@39509.4]
  wire [7:0] _T_874; // @[Modules.scala 108:54:@39510.4]
  wire [7:0] buffer_1_7; // @[Modules.scala 108:54:@39511.4]
  wire [7:0] _GEN_13; // @[Modules.scala 108:54:@39513.4]
  wire [8:0] _T_876; // @[Modules.scala 108:54:@39513.4]
  wire [7:0] _T_877; // @[Modules.scala 108:54:@39514.4]
  wire [7:0] buffer_1_8; // @[Modules.scala 108:54:@39515.4]
  wire [8:0] _T_879; // @[Modules.scala 108:54:@39518.4]
  wire [7:0] _T_880; // @[Modules.scala 108:54:@39519.4]
  wire [7:0] buffer_1_10; // @[Modules.scala 108:54:@39520.4]
  wire [8:0] _T_883; // @[Modules.scala 108:54:@39530.4]
  wire [7:0] _T_884; // @[Modules.scala 108:54:@39531.4]
  wire [7:0] buffer_2_2; // @[Modules.scala 108:54:@39532.4]
  wire [8:0] _T_886; // @[Modules.scala 108:54:@39534.4]
  wire [7:0] _T_887; // @[Modules.scala 108:54:@39535.4]
  wire [7:0] buffer_2_3; // @[Modules.scala 108:54:@39536.4]
  wire [8:0] _T_889; // @[Modules.scala 108:54:@39541.4]
  wire [7:0] _T_890; // @[Modules.scala 108:54:@39542.4]
  wire [7:0] buffer_2_7; // @[Modules.scala 108:54:@39543.4]
  wire [8:0] _T_892; // @[Modules.scala 108:54:@39545.4]
  wire [7:0] _T_893; // @[Modules.scala 108:54:@39546.4]
  wire [7:0] buffer_2_8; // @[Modules.scala 108:54:@39547.4]
  wire [8:0] _T_895; // @[Modules.scala 108:54:@39551.4]
  wire [7:0] _T_896; // @[Modules.scala 108:54:@39552.4]
  wire [7:0] buffer_2_11; // @[Modules.scala 108:54:@39553.4]
  wire [8:0] _T_898; // @[Modules.scala 108:54:@39555.4]
  wire [7:0] _T_899; // @[Modules.scala 108:54:@39556.4]
  wire [7:0] buffer_2_12; // @[Modules.scala 108:54:@39557.4]
  wire [8:0] _T_901; // @[Modules.scala 108:54:@39559.4]
  wire [7:0] _T_902; // @[Modules.scala 108:54:@39560.4]
  wire [7:0] buffer_2_13; // @[Modules.scala 108:54:@39561.4]
  wire [7:0] _GEN_22; // @[Modules.scala 108:54:@39563.4]
  wire [8:0] _T_904; // @[Modules.scala 108:54:@39563.4]
  wire [7:0] _T_905; // @[Modules.scala 108:54:@39564.4]
  wire [7:0] buffer_2_14; // @[Modules.scala 108:54:@39565.4]
  wire [8:0] _T_908; // @[Modules.scala 108:54:@39572.4]
  wire [7:0] _T_909; // @[Modules.scala 108:54:@39573.4]
  wire [7:0] buffer_3_3; // @[Modules.scala 108:54:@39574.4]
  wire [8:0] _T_911; // @[Modules.scala 108:54:@39576.4]
  wire [7:0] _T_912; // @[Modules.scala 108:54:@39577.4]
  wire [7:0] buffer_3_4; // @[Modules.scala 108:54:@39578.4]
  wire [8:0] _T_914; // @[Modules.scala 108:54:@39580.4]
  wire [7:0] _T_915; // @[Modules.scala 108:54:@39581.4]
  wire [7:0] buffer_3_5; // @[Modules.scala 108:54:@39582.4]
  wire [8:0] _T_917; // @[Modules.scala 108:54:@39585.4]
  wire [7:0] _T_918; // @[Modules.scala 108:54:@39586.4]
  wire [7:0] buffer_3_7; // @[Modules.scala 108:54:@39587.4]
  wire [8:0] _T_920; // @[Modules.scala 108:54:@39590.4]
  wire [7:0] _T_921; // @[Modules.scala 108:54:@39591.4]
  wire [7:0] buffer_3_9; // @[Modules.scala 108:54:@39592.4]
  wire [8:0] _T_923; // @[Modules.scala 108:54:@39596.4]
  wire [7:0] _T_924; // @[Modules.scala 108:54:@39597.4]
  wire [7:0] buffer_3_12; // @[Modules.scala 108:54:@39598.4]
  wire [8:0] _T_926; // @[Modules.scala 108:54:@39601.4]
  wire [7:0] _T_927; // @[Modules.scala 108:54:@39602.4]
  wire [7:0] buffer_3_14; // @[Modules.scala 108:54:@39603.4]
  wire [8:0] _T_929; // @[Modules.scala 108:54:@39608.4]
  wire [7:0] _T_930; // @[Modules.scala 108:54:@39609.4]
  wire [7:0] buffer_4_1; // @[Modules.scala 108:54:@39610.4]
  wire [8:0] _T_932; // @[Modules.scala 108:54:@39612.4]
  wire [7:0] _T_933; // @[Modules.scala 108:54:@39613.4]
  wire [7:0] buffer_4_2; // @[Modules.scala 108:54:@39614.4]
  wire [8:0] _T_935; // @[Modules.scala 108:54:@39617.4]
  wire [7:0] _T_936; // @[Modules.scala 108:54:@39618.4]
  wire [7:0] buffer_4_4; // @[Modules.scala 108:54:@39619.4]
  wire [8:0] _T_938; // @[Modules.scala 108:54:@39621.4]
  wire [7:0] _T_939; // @[Modules.scala 108:54:@39622.4]
  wire [7:0] buffer_4_5; // @[Modules.scala 108:54:@39623.4]
  wire [8:0] _T_941; // @[Modules.scala 108:54:@39625.4]
  wire [7:0] _T_942; // @[Modules.scala 108:54:@39626.4]
  wire [7:0] buffer_4_6; // @[Modules.scala 108:54:@39627.4]
  wire [8:0] _T_944; // @[Modules.scala 108:54:@39630.4]
  wire [7:0] _T_945; // @[Modules.scala 108:54:@39631.4]
  wire [7:0] buffer_4_8; // @[Modules.scala 108:54:@39632.4]
  wire [8:0] _T_947; // @[Modules.scala 108:54:@39634.4]
  wire [7:0] _T_948; // @[Modules.scala 108:54:@39635.4]
  wire [7:0] buffer_4_9; // @[Modules.scala 108:54:@39636.4]
  wire [8:0] _T_950; // @[Modules.scala 108:54:@39639.4]
  wire [7:0] _T_951; // @[Modules.scala 108:54:@39640.4]
  wire [7:0] buffer_4_11; // @[Modules.scala 108:54:@39641.4]
  wire [8:0] _T_953; // @[Modules.scala 108:54:@39644.4]
  wire [7:0] _T_954; // @[Modules.scala 108:54:@39645.4]
  wire [7:0] buffer_4_13; // @[Modules.scala 108:54:@39646.4]
  wire [8:0] _T_956; // @[Modules.scala 108:54:@39648.4]
  wire [7:0] _T_957; // @[Modules.scala 108:54:@39649.4]
  wire [7:0] buffer_4_14; // @[Modules.scala 108:54:@39650.4]
  wire [8:0] _T_959; // @[Modules.scala 108:54:@39652.4]
  wire [7:0] _T_960; // @[Modules.scala 108:54:@39653.4]
  wire [7:0] buffer_4_15; // @[Modules.scala 108:54:@39654.4]
  wire [8:0] _T_965; // @[Modules.scala 108:54:@39664.4]
  wire [7:0] _T_966; // @[Modules.scala 108:54:@39665.4]
  wire [7:0] buffer_5_4; // @[Modules.scala 108:54:@39666.4]
  wire [8:0] _T_968; // @[Modules.scala 108:54:@39668.4]
  wire [7:0] _T_969; // @[Modules.scala 108:54:@39669.4]
  wire [7:0] buffer_5_5; // @[Modules.scala 108:54:@39670.4]
  wire [8:0] _T_971; // @[Modules.scala 108:54:@39672.4]
  wire [7:0] _T_972; // @[Modules.scala 108:54:@39673.4]
  wire [7:0] buffer_5_6; // @[Modules.scala 108:54:@39674.4]
  wire [8:0] _T_974; // @[Modules.scala 108:54:@39678.4]
  wire [7:0] _T_975; // @[Modules.scala 108:54:@39679.4]
  wire [7:0] buffer_5_9; // @[Modules.scala 108:54:@39680.4]
  wire [8:0] _T_977; // @[Modules.scala 108:54:@39682.4]
  wire [7:0] _T_978; // @[Modules.scala 108:54:@39683.4]
  wire [7:0] buffer_5_10; // @[Modules.scala 108:54:@39684.4]
  wire [8:0] _T_980; // @[Modules.scala 108:54:@39687.4]
  wire [7:0] _T_981; // @[Modules.scala 108:54:@39688.4]
  wire [7:0] buffer_5_12; // @[Modules.scala 108:54:@39689.4]
  wire [8:0] _T_983; // @[Modules.scala 108:54:@39691.4]
  wire [7:0] _T_984; // @[Modules.scala 108:54:@39692.4]
  wire [7:0] buffer_5_13; // @[Modules.scala 108:54:@39693.4]
  wire [8:0] _T_990; // @[Modules.scala 108:54:@39703.4]
  wire [7:0] _T_991; // @[Modules.scala 108:54:@39704.4]
  wire [7:0] buffer_6_2; // @[Modules.scala 108:54:@39705.4]
  wire [8:0] _T_993; // @[Modules.scala 108:54:@39708.4]
  wire [7:0] _T_994; // @[Modules.scala 108:54:@39709.4]
  wire [7:0] buffer_6_4; // @[Modules.scala 108:54:@39710.4]
  wire [8:0] _T_996; // @[Modules.scala 108:54:@39712.4]
  wire [7:0] _T_997; // @[Modules.scala 108:54:@39713.4]
  wire [7:0] buffer_6_5; // @[Modules.scala 108:54:@39714.4]
  wire [8:0] _T_999; // @[Modules.scala 108:54:@39718.4]
  wire [7:0] _T_1000; // @[Modules.scala 108:54:@39719.4]
  wire [7:0] buffer_6_8; // @[Modules.scala 108:54:@39720.4]
  wire [8:0] _T_1002; // @[Modules.scala 108:54:@39723.4]
  wire [7:0] _T_1003; // @[Modules.scala 108:54:@39724.4]
  wire [7:0] buffer_6_10; // @[Modules.scala 108:54:@39725.4]
  wire [8:0] _T_1005; // @[Modules.scala 108:54:@39728.4]
  wire [7:0] _T_1006; // @[Modules.scala 108:54:@39729.4]
  wire [7:0] buffer_6_12; // @[Modules.scala 108:54:@39730.4]
  wire [8:0] _T_1008; // @[Modules.scala 108:54:@39732.4]
  wire [7:0] _T_1009; // @[Modules.scala 108:54:@39733.4]
  wire [7:0] buffer_6_13; // @[Modules.scala 108:54:@39734.4]
  wire [8:0] _T_1011; // @[Modules.scala 108:54:@39736.4]
  wire [7:0] _T_1012; // @[Modules.scala 108:54:@39737.4]
  wire [7:0] buffer_6_14; // @[Modules.scala 108:54:@39738.4]
  wire [8:0] _T_1014; // @[Modules.scala 108:54:@39740.4]
  wire [7:0] _T_1015; // @[Modules.scala 108:54:@39741.4]
  wire [7:0] buffer_6_15; // @[Modules.scala 108:54:@39742.4]
  wire [8:0] _T_1020; // @[Modules.scala 108:54:@39751.4]
  wire [7:0] _T_1021; // @[Modules.scala 108:54:@39752.4]
  wire [7:0] buffer_7_3; // @[Modules.scala 108:54:@39753.4]
  wire [8:0] _T_1023; // @[Modules.scala 108:54:@39758.4]
  wire [7:0] _T_1024; // @[Modules.scala 108:54:@39759.4]
  wire [7:0] buffer_7_7; // @[Modules.scala 108:54:@39760.4]
  wire [8:0] _T_1026; // @[Modules.scala 108:54:@39762.4]
  wire [7:0] _T_1027; // @[Modules.scala 108:54:@39763.4]
  wire [7:0] buffer_7_8; // @[Modules.scala 108:54:@39764.4]
  wire [8:0] _T_1029; // @[Modules.scala 108:54:@39766.4]
  wire [7:0] _T_1030; // @[Modules.scala 108:54:@39767.4]
  wire [7:0] buffer_7_9; // @[Modules.scala 108:54:@39768.4]
  wire [8:0] _T_1032; // @[Modules.scala 108:54:@39770.4]
  wire [7:0] _T_1033; // @[Modules.scala 108:54:@39771.4]
  wire [7:0] buffer_7_10; // @[Modules.scala 108:54:@39772.4]
  wire [8:0] _T_1035; // @[Modules.scala 108:54:@39774.4]
  wire [7:0] _T_1036; // @[Modules.scala 108:54:@39775.4]
  wire [7:0] buffer_7_11; // @[Modules.scala 108:54:@39776.4]
  wire [8:0] _T_1038; // @[Modules.scala 108:54:@39781.4]
  wire [7:0] _T_1039; // @[Modules.scala 108:54:@39782.4]
  wire [7:0] buffer_7_15; // @[Modules.scala 108:54:@39783.4]
  wire [8:0] _T_1044; // @[Modules.scala 108:54:@39794.4]
  wire [7:0] _T_1045; // @[Modules.scala 108:54:@39795.4]
  wire [7:0] buffer_8_5; // @[Modules.scala 108:54:@39796.4]
  wire [8:0] _T_1047; // @[Modules.scala 108:54:@39798.4]
  wire [7:0] _T_1048; // @[Modules.scala 108:54:@39799.4]
  wire [7:0] buffer_8_6; // @[Modules.scala 108:54:@39800.4]
  wire [8:0] _T_1050; // @[Modules.scala 108:54:@39807.4]
  wire [7:0] _T_1051; // @[Modules.scala 108:54:@39808.4]
  wire [7:0] buffer_8_12; // @[Modules.scala 108:54:@39809.4]
  wire [8:0] _T_1053; // @[Modules.scala 108:54:@39812.4]
  wire [7:0] _T_1054; // @[Modules.scala 108:54:@39813.4]
  wire [7:0] buffer_8_14; // @[Modules.scala 108:54:@39814.4]
  wire [8:0] _T_1059; // @[Modules.scala 108:54:@39827.4]
  wire [7:0] _T_1060; // @[Modules.scala 108:54:@39828.4]
  wire [7:0] buffer_9_6; // @[Modules.scala 108:54:@39829.4]
  wire [8:0] _T_1062; // @[Modules.scala 108:54:@39831.4]
  wire [7:0] _T_1063; // @[Modules.scala 108:54:@39832.4]
  wire [7:0] buffer_9_7; // @[Modules.scala 108:54:@39833.4]
  wire [8:0] _T_1065; // @[Modules.scala 108:54:@39835.4]
  wire [7:0] _T_1066; // @[Modules.scala 108:54:@39836.4]
  wire [7:0] buffer_9_8; // @[Modules.scala 108:54:@39837.4]
  wire [8:0] _T_1068; // @[Modules.scala 108:54:@39839.4]
  wire [7:0] _T_1069; // @[Modules.scala 108:54:@39840.4]
  wire [7:0] buffer_9_9; // @[Modules.scala 108:54:@39841.4]
  wire [8:0] _T_1071; // @[Modules.scala 108:54:@39847.4]
  wire [7:0] _T_1072; // @[Modules.scala 108:54:@39848.4]
  wire [7:0] buffer_9_14; // @[Modules.scala 108:54:@39849.4]
  wire [8:0] _T_1074; // @[Modules.scala 108:54:@39851.4]
  wire [7:0] _T_1075; // @[Modules.scala 108:54:@39852.4]
  wire [7:0] buffer_9_15; // @[Modules.scala 108:54:@39853.4]
  assign _GEN_0 = {{6{io_in_1[1]}},io_in_1}; // @[Modules.scala 108:54:@39450.4]
  assign _T_837 = $signed(8'sh0) + $signed(_GEN_0); // @[Modules.scala 108:54:@39450.4]
  assign _T_838 = _T_837[7:0]; // @[Modules.scala 108:54:@39451.4]
  assign buffer_0_1 = $signed(_T_838); // @[Modules.scala 108:54:@39452.4]
  assign _GEN_1 = {{6{io_in_9[1]}},io_in_9}; // @[Modules.scala 108:54:@39461.4]
  assign _T_840 = $signed(buffer_0_1) + $signed(_GEN_1); // @[Modules.scala 108:54:@39461.4]
  assign _T_841 = _T_840[7:0]; // @[Modules.scala 108:54:@39462.4]
  assign buffer_0_9 = $signed(_T_841); // @[Modules.scala 108:54:@39463.4]
  assign _GEN_2 = {{6{io_in_10[1]}},io_in_10}; // @[Modules.scala 108:54:@39465.4]
  assign _T_843 = $signed(buffer_0_9) + $signed(_GEN_2); // @[Modules.scala 108:54:@39465.4]
  assign _T_844 = _T_843[7:0]; // @[Modules.scala 108:54:@39466.4]
  assign buffer_0_10 = $signed(_T_844); // @[Modules.scala 108:54:@39467.4]
  assign _GEN_3 = {{6{io_in_11[1]}},io_in_11}; // @[Modules.scala 108:54:@39469.4]
  assign _T_846 = $signed(buffer_0_10) + $signed(_GEN_3); // @[Modules.scala 108:54:@39469.4]
  assign _T_847 = _T_846[7:0]; // @[Modules.scala 108:54:@39470.4]
  assign buffer_0_11 = $signed(_T_847); // @[Modules.scala 108:54:@39471.4]
  assign _GEN_4 = {{6{io_in_12[1]}},io_in_12}; // @[Modules.scala 108:54:@39473.4]
  assign _T_849 = $signed(buffer_0_11) + $signed(_GEN_4); // @[Modules.scala 108:54:@39473.4]
  assign _T_850 = _T_849[7:0]; // @[Modules.scala 108:54:@39474.4]
  assign buffer_0_12 = $signed(_T_850); // @[Modules.scala 108:54:@39475.4]
  assign _GEN_5 = {{6{io_in_13[1]}},io_in_13}; // @[Modules.scala 108:54:@39477.4]
  assign _T_852 = $signed(buffer_0_12) + $signed(_GEN_5); // @[Modules.scala 108:54:@39477.4]
  assign _T_853 = _T_852[7:0]; // @[Modules.scala 108:54:@39478.4]
  assign buffer_0_13 = $signed(_T_853); // @[Modules.scala 108:54:@39479.4]
  assign _GEN_6 = {{6{io_in_15[1]}},io_in_15}; // @[Modules.scala 108:54:@39482.4]
  assign _T_855 = $signed(buffer_0_13) + $signed(_GEN_6); // @[Modules.scala 108:54:@39482.4]
  assign _T_856 = _T_855[7:0]; // @[Modules.scala 108:54:@39483.4]
  assign buffer_0_15 = $signed(_T_856); // @[Modules.scala 108:54:@39484.4]
  assign buffer_1_0 = {{6{io_in_0[1]}},io_in_0}; // @[Modules.scala 91:22:@39448.4]
  assign _GEN_7 = {{6{io_in_2[1]}},io_in_2}; // @[Modules.scala 108:54:@39489.4]
  assign _T_858 = $signed(buffer_1_0) + $signed(_GEN_7); // @[Modules.scala 108:54:@39489.4]
  assign _T_859 = _T_858[7:0]; // @[Modules.scala 108:54:@39490.4]
  assign buffer_1_2 = $signed(_T_859); // @[Modules.scala 108:54:@39491.4]
  assign _GEN_8 = {{6{io_in_3[1]}},io_in_3}; // @[Modules.scala 108:54:@39493.4]
  assign _T_861 = $signed(buffer_1_2) + $signed(_GEN_8); // @[Modules.scala 108:54:@39493.4]
  assign _T_862 = _T_861[7:0]; // @[Modules.scala 108:54:@39494.4]
  assign buffer_1_3 = $signed(_T_862); // @[Modules.scala 108:54:@39495.4]
  assign _GEN_9 = {{6{io_in_4[1]}},io_in_4}; // @[Modules.scala 108:54:@39497.4]
  assign _T_864 = $signed(buffer_1_3) + $signed(_GEN_9); // @[Modules.scala 108:54:@39497.4]
  assign _T_865 = _T_864[7:0]; // @[Modules.scala 108:54:@39498.4]
  assign buffer_1_4 = $signed(_T_865); // @[Modules.scala 108:54:@39499.4]
  assign _GEN_10 = {{6{io_in_5[1]}},io_in_5}; // @[Modules.scala 108:54:@39501.4]
  assign _T_867 = $signed(buffer_1_4) + $signed(_GEN_10); // @[Modules.scala 108:54:@39501.4]
  assign _T_868 = _T_867[7:0]; // @[Modules.scala 108:54:@39502.4]
  assign buffer_1_5 = $signed(_T_868); // @[Modules.scala 108:54:@39503.4]
  assign _GEN_11 = {{6{io_in_6[1]}},io_in_6}; // @[Modules.scala 108:54:@39505.4]
  assign _T_870 = $signed(buffer_1_5) + $signed(_GEN_11); // @[Modules.scala 108:54:@39505.4]
  assign _T_871 = _T_870[7:0]; // @[Modules.scala 108:54:@39506.4]
  assign buffer_1_6 = $signed(_T_871); // @[Modules.scala 108:54:@39507.4]
  assign _GEN_12 = {{6{io_in_7[1]}},io_in_7}; // @[Modules.scala 108:54:@39509.4]
  assign _T_873 = $signed(buffer_1_6) + $signed(_GEN_12); // @[Modules.scala 108:54:@39509.4]
  assign _T_874 = _T_873[7:0]; // @[Modules.scala 108:54:@39510.4]
  assign buffer_1_7 = $signed(_T_874); // @[Modules.scala 108:54:@39511.4]
  assign _GEN_13 = {{6{io_in_8[1]}},io_in_8}; // @[Modules.scala 108:54:@39513.4]
  assign _T_876 = $signed(buffer_1_7) + $signed(_GEN_13); // @[Modules.scala 108:54:@39513.4]
  assign _T_877 = _T_876[7:0]; // @[Modules.scala 108:54:@39514.4]
  assign buffer_1_8 = $signed(_T_877); // @[Modules.scala 108:54:@39515.4]
  assign _T_879 = $signed(buffer_1_8) + $signed(_GEN_2); // @[Modules.scala 108:54:@39518.4]
  assign _T_880 = _T_879[7:0]; // @[Modules.scala 108:54:@39519.4]
  assign buffer_1_10 = $signed(_T_880); // @[Modules.scala 108:54:@39520.4]
  assign _T_883 = $signed(8'sh0) + $signed(_GEN_7); // @[Modules.scala 108:54:@39530.4]
  assign _T_884 = _T_883[7:0]; // @[Modules.scala 108:54:@39531.4]
  assign buffer_2_2 = $signed(_T_884); // @[Modules.scala 108:54:@39532.4]
  assign _T_886 = $signed(buffer_2_2) + $signed(_GEN_8); // @[Modules.scala 108:54:@39534.4]
  assign _T_887 = _T_886[7:0]; // @[Modules.scala 108:54:@39535.4]
  assign buffer_2_3 = $signed(_T_887); // @[Modules.scala 108:54:@39536.4]
  assign _T_889 = $signed(buffer_2_3) + $signed(_GEN_12); // @[Modules.scala 108:54:@39541.4]
  assign _T_890 = _T_889[7:0]; // @[Modules.scala 108:54:@39542.4]
  assign buffer_2_7 = $signed(_T_890); // @[Modules.scala 108:54:@39543.4]
  assign _T_892 = $signed(buffer_2_7) + $signed(_GEN_13); // @[Modules.scala 108:54:@39545.4]
  assign _T_893 = _T_892[7:0]; // @[Modules.scala 108:54:@39546.4]
  assign buffer_2_8 = $signed(_T_893); // @[Modules.scala 108:54:@39547.4]
  assign _T_895 = $signed(buffer_2_8) + $signed(_GEN_3); // @[Modules.scala 108:54:@39551.4]
  assign _T_896 = _T_895[7:0]; // @[Modules.scala 108:54:@39552.4]
  assign buffer_2_11 = $signed(_T_896); // @[Modules.scala 108:54:@39553.4]
  assign _T_898 = $signed(buffer_2_11) + $signed(_GEN_4); // @[Modules.scala 108:54:@39555.4]
  assign _T_899 = _T_898[7:0]; // @[Modules.scala 108:54:@39556.4]
  assign buffer_2_12 = $signed(_T_899); // @[Modules.scala 108:54:@39557.4]
  assign _T_901 = $signed(buffer_2_12) + $signed(_GEN_5); // @[Modules.scala 108:54:@39559.4]
  assign _T_902 = _T_901[7:0]; // @[Modules.scala 108:54:@39560.4]
  assign buffer_2_13 = $signed(_T_902); // @[Modules.scala 108:54:@39561.4]
  assign _GEN_22 = {{6{io_in_14[1]}},io_in_14}; // @[Modules.scala 108:54:@39563.4]
  assign _T_904 = $signed(buffer_2_13) + $signed(_GEN_22); // @[Modules.scala 108:54:@39563.4]
  assign _T_905 = _T_904[7:0]; // @[Modules.scala 108:54:@39564.4]
  assign buffer_2_14 = $signed(_T_905); // @[Modules.scala 108:54:@39565.4]
  assign _T_908 = $signed(8'sh0) + $signed(_GEN_8); // @[Modules.scala 108:54:@39572.4]
  assign _T_909 = _T_908[7:0]; // @[Modules.scala 108:54:@39573.4]
  assign buffer_3_3 = $signed(_T_909); // @[Modules.scala 108:54:@39574.4]
  assign _T_911 = $signed(buffer_3_3) + $signed(_GEN_9); // @[Modules.scala 108:54:@39576.4]
  assign _T_912 = _T_911[7:0]; // @[Modules.scala 108:54:@39577.4]
  assign buffer_3_4 = $signed(_T_912); // @[Modules.scala 108:54:@39578.4]
  assign _T_914 = $signed(buffer_3_4) + $signed(_GEN_10); // @[Modules.scala 108:54:@39580.4]
  assign _T_915 = _T_914[7:0]; // @[Modules.scala 108:54:@39581.4]
  assign buffer_3_5 = $signed(_T_915); // @[Modules.scala 108:54:@39582.4]
  assign _T_917 = $signed(buffer_3_5) + $signed(_GEN_12); // @[Modules.scala 108:54:@39585.4]
  assign _T_918 = _T_917[7:0]; // @[Modules.scala 108:54:@39586.4]
  assign buffer_3_7 = $signed(_T_918); // @[Modules.scala 108:54:@39587.4]
  assign _T_920 = $signed(buffer_3_7) + $signed(_GEN_1); // @[Modules.scala 108:54:@39590.4]
  assign _T_921 = _T_920[7:0]; // @[Modules.scala 108:54:@39591.4]
  assign buffer_3_9 = $signed(_T_921); // @[Modules.scala 108:54:@39592.4]
  assign _T_923 = $signed(buffer_3_9) + $signed(_GEN_4); // @[Modules.scala 108:54:@39596.4]
  assign _T_924 = _T_923[7:0]; // @[Modules.scala 108:54:@39597.4]
  assign buffer_3_12 = $signed(_T_924); // @[Modules.scala 108:54:@39598.4]
  assign _T_926 = $signed(buffer_3_12) + $signed(_GEN_22); // @[Modules.scala 108:54:@39601.4]
  assign _T_927 = _T_926[7:0]; // @[Modules.scala 108:54:@39602.4]
  assign buffer_3_14 = $signed(_T_927); // @[Modules.scala 108:54:@39603.4]
  assign _T_929 = $signed(buffer_1_0) + $signed(_GEN_0); // @[Modules.scala 108:54:@39608.4]
  assign _T_930 = _T_929[7:0]; // @[Modules.scala 108:54:@39609.4]
  assign buffer_4_1 = $signed(_T_930); // @[Modules.scala 108:54:@39610.4]
  assign _T_932 = $signed(buffer_4_1) + $signed(_GEN_7); // @[Modules.scala 108:54:@39612.4]
  assign _T_933 = _T_932[7:0]; // @[Modules.scala 108:54:@39613.4]
  assign buffer_4_2 = $signed(_T_933); // @[Modules.scala 108:54:@39614.4]
  assign _T_935 = $signed(buffer_4_2) + $signed(_GEN_9); // @[Modules.scala 108:54:@39617.4]
  assign _T_936 = _T_935[7:0]; // @[Modules.scala 108:54:@39618.4]
  assign buffer_4_4 = $signed(_T_936); // @[Modules.scala 108:54:@39619.4]
  assign _T_938 = $signed(buffer_4_4) + $signed(_GEN_10); // @[Modules.scala 108:54:@39621.4]
  assign _T_939 = _T_938[7:0]; // @[Modules.scala 108:54:@39622.4]
  assign buffer_4_5 = $signed(_T_939); // @[Modules.scala 108:54:@39623.4]
  assign _T_941 = $signed(buffer_4_5) + $signed(_GEN_11); // @[Modules.scala 108:54:@39625.4]
  assign _T_942 = _T_941[7:0]; // @[Modules.scala 108:54:@39626.4]
  assign buffer_4_6 = $signed(_T_942); // @[Modules.scala 108:54:@39627.4]
  assign _T_944 = $signed(buffer_4_6) + $signed(_GEN_13); // @[Modules.scala 108:54:@39630.4]
  assign _T_945 = _T_944[7:0]; // @[Modules.scala 108:54:@39631.4]
  assign buffer_4_8 = $signed(_T_945); // @[Modules.scala 108:54:@39632.4]
  assign _T_947 = $signed(buffer_4_8) + $signed(_GEN_1); // @[Modules.scala 108:54:@39634.4]
  assign _T_948 = _T_947[7:0]; // @[Modules.scala 108:54:@39635.4]
  assign buffer_4_9 = $signed(_T_948); // @[Modules.scala 108:54:@39636.4]
  assign _T_950 = $signed(buffer_4_9) + $signed(_GEN_3); // @[Modules.scala 108:54:@39639.4]
  assign _T_951 = _T_950[7:0]; // @[Modules.scala 108:54:@39640.4]
  assign buffer_4_11 = $signed(_T_951); // @[Modules.scala 108:54:@39641.4]
  assign _T_953 = $signed(buffer_4_11) + $signed(_GEN_5); // @[Modules.scala 108:54:@39644.4]
  assign _T_954 = _T_953[7:0]; // @[Modules.scala 108:54:@39645.4]
  assign buffer_4_13 = $signed(_T_954); // @[Modules.scala 108:54:@39646.4]
  assign _T_956 = $signed(buffer_4_13) + $signed(_GEN_22); // @[Modules.scala 108:54:@39648.4]
  assign _T_957 = _T_956[7:0]; // @[Modules.scala 108:54:@39649.4]
  assign buffer_4_14 = $signed(_T_957); // @[Modules.scala 108:54:@39650.4]
  assign _T_959 = $signed(buffer_4_14) + $signed(_GEN_6); // @[Modules.scala 108:54:@39652.4]
  assign _T_960 = _T_959[7:0]; // @[Modules.scala 108:54:@39653.4]
  assign buffer_4_15 = $signed(_T_960); // @[Modules.scala 108:54:@39654.4]
  assign _T_965 = $signed(buffer_4_1) + $signed(_GEN_9); // @[Modules.scala 108:54:@39664.4]
  assign _T_966 = _T_965[7:0]; // @[Modules.scala 108:54:@39665.4]
  assign buffer_5_4 = $signed(_T_966); // @[Modules.scala 108:54:@39666.4]
  assign _T_968 = $signed(buffer_5_4) + $signed(_GEN_10); // @[Modules.scala 108:54:@39668.4]
  assign _T_969 = _T_968[7:0]; // @[Modules.scala 108:54:@39669.4]
  assign buffer_5_5 = $signed(_T_969); // @[Modules.scala 108:54:@39670.4]
  assign _T_971 = $signed(buffer_5_5) + $signed(_GEN_11); // @[Modules.scala 108:54:@39672.4]
  assign _T_972 = _T_971[7:0]; // @[Modules.scala 108:54:@39673.4]
  assign buffer_5_6 = $signed(_T_972); // @[Modules.scala 108:54:@39674.4]
  assign _T_974 = $signed(buffer_5_6) + $signed(_GEN_1); // @[Modules.scala 108:54:@39678.4]
  assign _T_975 = _T_974[7:0]; // @[Modules.scala 108:54:@39679.4]
  assign buffer_5_9 = $signed(_T_975); // @[Modules.scala 108:54:@39680.4]
  assign _T_977 = $signed(buffer_5_9) + $signed(_GEN_2); // @[Modules.scala 108:54:@39682.4]
  assign _T_978 = _T_977[7:0]; // @[Modules.scala 108:54:@39683.4]
  assign buffer_5_10 = $signed(_T_978); // @[Modules.scala 108:54:@39684.4]
  assign _T_980 = $signed(buffer_5_10) + $signed(_GEN_4); // @[Modules.scala 108:54:@39687.4]
  assign _T_981 = _T_980[7:0]; // @[Modules.scala 108:54:@39688.4]
  assign buffer_5_12 = $signed(_T_981); // @[Modules.scala 108:54:@39689.4]
  assign _T_983 = $signed(buffer_5_12) + $signed(_GEN_5); // @[Modules.scala 108:54:@39691.4]
  assign _T_984 = _T_983[7:0]; // @[Modules.scala 108:54:@39692.4]
  assign buffer_5_13 = $signed(_T_984); // @[Modules.scala 108:54:@39693.4]
  assign _T_990 = $signed(buffer_0_1) + $signed(_GEN_7); // @[Modules.scala 108:54:@39703.4]
  assign _T_991 = _T_990[7:0]; // @[Modules.scala 108:54:@39704.4]
  assign buffer_6_2 = $signed(_T_991); // @[Modules.scala 108:54:@39705.4]
  assign _T_993 = $signed(buffer_6_2) + $signed(_GEN_9); // @[Modules.scala 108:54:@39708.4]
  assign _T_994 = _T_993[7:0]; // @[Modules.scala 108:54:@39709.4]
  assign buffer_6_4 = $signed(_T_994); // @[Modules.scala 108:54:@39710.4]
  assign _T_996 = $signed(buffer_6_4) + $signed(_GEN_10); // @[Modules.scala 108:54:@39712.4]
  assign _T_997 = _T_996[7:0]; // @[Modules.scala 108:54:@39713.4]
  assign buffer_6_5 = $signed(_T_997); // @[Modules.scala 108:54:@39714.4]
  assign _T_999 = $signed(buffer_6_5) + $signed(_GEN_13); // @[Modules.scala 108:54:@39718.4]
  assign _T_1000 = _T_999[7:0]; // @[Modules.scala 108:54:@39719.4]
  assign buffer_6_8 = $signed(_T_1000); // @[Modules.scala 108:54:@39720.4]
  assign _T_1002 = $signed(buffer_6_8) + $signed(_GEN_2); // @[Modules.scala 108:54:@39723.4]
  assign _T_1003 = _T_1002[7:0]; // @[Modules.scala 108:54:@39724.4]
  assign buffer_6_10 = $signed(_T_1003); // @[Modules.scala 108:54:@39725.4]
  assign _T_1005 = $signed(buffer_6_10) + $signed(_GEN_4); // @[Modules.scala 108:54:@39728.4]
  assign _T_1006 = _T_1005[7:0]; // @[Modules.scala 108:54:@39729.4]
  assign buffer_6_12 = $signed(_T_1006); // @[Modules.scala 108:54:@39730.4]
  assign _T_1008 = $signed(buffer_6_12) + $signed(_GEN_5); // @[Modules.scala 108:54:@39732.4]
  assign _T_1009 = _T_1008[7:0]; // @[Modules.scala 108:54:@39733.4]
  assign buffer_6_13 = $signed(_T_1009); // @[Modules.scala 108:54:@39734.4]
  assign _T_1011 = $signed(buffer_6_13) + $signed(_GEN_22); // @[Modules.scala 108:54:@39736.4]
  assign _T_1012 = _T_1011[7:0]; // @[Modules.scala 108:54:@39737.4]
  assign buffer_6_14 = $signed(_T_1012); // @[Modules.scala 108:54:@39738.4]
  assign _T_1014 = $signed(buffer_6_14) + $signed(_GEN_6); // @[Modules.scala 108:54:@39740.4]
  assign _T_1015 = _T_1014[7:0]; // @[Modules.scala 108:54:@39741.4]
  assign buffer_6_15 = $signed(_T_1015); // @[Modules.scala 108:54:@39742.4]
  assign _T_1020 = $signed(buffer_4_1) + $signed(_GEN_8); // @[Modules.scala 108:54:@39751.4]
  assign _T_1021 = _T_1020[7:0]; // @[Modules.scala 108:54:@39752.4]
  assign buffer_7_3 = $signed(_T_1021); // @[Modules.scala 108:54:@39753.4]
  assign _T_1023 = $signed(buffer_7_3) + $signed(_GEN_12); // @[Modules.scala 108:54:@39758.4]
  assign _T_1024 = _T_1023[7:0]; // @[Modules.scala 108:54:@39759.4]
  assign buffer_7_7 = $signed(_T_1024); // @[Modules.scala 108:54:@39760.4]
  assign _T_1026 = $signed(buffer_7_7) + $signed(_GEN_13); // @[Modules.scala 108:54:@39762.4]
  assign _T_1027 = _T_1026[7:0]; // @[Modules.scala 108:54:@39763.4]
  assign buffer_7_8 = $signed(_T_1027); // @[Modules.scala 108:54:@39764.4]
  assign _T_1029 = $signed(buffer_7_8) + $signed(_GEN_1); // @[Modules.scala 108:54:@39766.4]
  assign _T_1030 = _T_1029[7:0]; // @[Modules.scala 108:54:@39767.4]
  assign buffer_7_9 = $signed(_T_1030); // @[Modules.scala 108:54:@39768.4]
  assign _T_1032 = $signed(buffer_7_9) + $signed(_GEN_2); // @[Modules.scala 108:54:@39770.4]
  assign _T_1033 = _T_1032[7:0]; // @[Modules.scala 108:54:@39771.4]
  assign buffer_7_10 = $signed(_T_1033); // @[Modules.scala 108:54:@39772.4]
  assign _T_1035 = $signed(buffer_7_10) + $signed(_GEN_3); // @[Modules.scala 108:54:@39774.4]
  assign _T_1036 = _T_1035[7:0]; // @[Modules.scala 108:54:@39775.4]
  assign buffer_7_11 = $signed(_T_1036); // @[Modules.scala 108:54:@39776.4]
  assign _T_1038 = $signed(buffer_7_11) + $signed(_GEN_6); // @[Modules.scala 108:54:@39781.4]
  assign _T_1039 = _T_1038[7:0]; // @[Modules.scala 108:54:@39782.4]
  assign buffer_7_15 = $signed(_T_1039); // @[Modules.scala 108:54:@39783.4]
  assign _T_1044 = $signed(buffer_1_2) + $signed(_GEN_10); // @[Modules.scala 108:54:@39794.4]
  assign _T_1045 = _T_1044[7:0]; // @[Modules.scala 108:54:@39795.4]
  assign buffer_8_5 = $signed(_T_1045); // @[Modules.scala 108:54:@39796.4]
  assign _T_1047 = $signed(buffer_8_5) + $signed(_GEN_11); // @[Modules.scala 108:54:@39798.4]
  assign _T_1048 = _T_1047[7:0]; // @[Modules.scala 108:54:@39799.4]
  assign buffer_8_6 = $signed(_T_1048); // @[Modules.scala 108:54:@39800.4]
  assign _T_1050 = $signed(buffer_8_6) + $signed(_GEN_4); // @[Modules.scala 108:54:@39807.4]
  assign _T_1051 = _T_1050[7:0]; // @[Modules.scala 108:54:@39808.4]
  assign buffer_8_12 = $signed(_T_1051); // @[Modules.scala 108:54:@39809.4]
  assign _T_1053 = $signed(buffer_8_12) + $signed(_GEN_22); // @[Modules.scala 108:54:@39812.4]
  assign _T_1054 = _T_1053[7:0]; // @[Modules.scala 108:54:@39813.4]
  assign buffer_8_14 = $signed(_T_1054); // @[Modules.scala 108:54:@39814.4]
  assign _T_1059 = $signed(buffer_4_1) + $signed(_GEN_11); // @[Modules.scala 108:54:@39827.4]
  assign _T_1060 = _T_1059[7:0]; // @[Modules.scala 108:54:@39828.4]
  assign buffer_9_6 = $signed(_T_1060); // @[Modules.scala 108:54:@39829.4]
  assign _T_1062 = $signed(buffer_9_6) + $signed(_GEN_12); // @[Modules.scala 108:54:@39831.4]
  assign _T_1063 = _T_1062[7:0]; // @[Modules.scala 108:54:@39832.4]
  assign buffer_9_7 = $signed(_T_1063); // @[Modules.scala 108:54:@39833.4]
  assign _T_1065 = $signed(buffer_9_7) + $signed(_GEN_13); // @[Modules.scala 108:54:@39835.4]
  assign _T_1066 = _T_1065[7:0]; // @[Modules.scala 108:54:@39836.4]
  assign buffer_9_8 = $signed(_T_1066); // @[Modules.scala 108:54:@39837.4]
  assign _T_1068 = $signed(buffer_9_8) + $signed(_GEN_1); // @[Modules.scala 108:54:@39839.4]
  assign _T_1069 = _T_1068[7:0]; // @[Modules.scala 108:54:@39840.4]
  assign buffer_9_9 = $signed(_T_1069); // @[Modules.scala 108:54:@39841.4]
  assign _T_1071 = $signed(buffer_9_9) + $signed(_GEN_22); // @[Modules.scala 108:54:@39847.4]
  assign _T_1072 = _T_1071[7:0]; // @[Modules.scala 108:54:@39848.4]
  assign buffer_9_14 = $signed(_T_1072); // @[Modules.scala 108:54:@39849.4]
  assign _T_1074 = $signed(buffer_9_14) + $signed(_GEN_6); // @[Modules.scala 108:54:@39851.4]
  assign _T_1075 = _T_1074[7:0]; // @[Modules.scala 108:54:@39852.4]
  assign buffer_9_15 = $signed(_T_1075); // @[Modules.scala 108:54:@39853.4]
  assign io_out_0 = buffer_0_15;
  assign io_out_1 = buffer_1_10;
  assign io_out_2 = buffer_2_14;
  assign io_out_3 = buffer_3_14;
  assign io_out_4 = buffer_4_15;
  assign io_out_5 = buffer_5_13;
  assign io_out_6 = buffer_6_15;
  assign io_out_7 = buffer_7_15;
  assign io_out_8 = buffer_8_14;
  assign io_out_9 = buffer_9_15;
endmodule
module ShifBatchNorm_2( // @[:@39857.2]
  input  [7:0] io_in_0, // @[:@39860.4]
  input  [7:0] io_in_1, // @[:@39860.4]
  input  [7:0] io_in_2, // @[:@39860.4]
  input  [7:0] io_in_3, // @[:@39860.4]
  input  [7:0] io_in_4, // @[:@39860.4]
  input  [7:0] io_in_5, // @[:@39860.4]
  input  [7:0] io_in_6, // @[:@39860.4]
  input  [7:0] io_in_7, // @[:@39860.4]
  input  [7:0] io_in_8, // @[:@39860.4]
  input  [7:0] io_in_9, // @[:@39860.4]
  output [7:0] io_out_0, // @[:@39860.4]
  output [7:0] io_out_1, // @[:@39860.4]
  output [7:0] io_out_2, // @[:@39860.4]
  output [7:0] io_out_3, // @[:@39860.4]
  output [7:0] io_out_4, // @[:@39860.4]
  output [7:0] io_out_5, // @[:@39860.4]
  output [7:0] io_out_6, // @[:@39860.4]
  output [7:0] io_out_7, // @[:@39860.4]
  output [7:0] io_out_8, // @[:@39860.4]
  output [7:0] io_out_9 // @[:@39860.4]
);
  wire [8:0] _T_78; // @[Modules.scala 132:28:@39865.4]
  wire [7:0] _T_79; // @[Modules.scala 132:28:@39866.4]
  wire [7:0] c_x_0; // @[Modules.scala 132:28:@39867.4]
  wire [22:0] _GEN_0; // @[Modules.scala 137:32:@39869.4]
  wire [22:0] _T_82; // @[Modules.scala 137:32:@39869.4]
  wire [7:0] _GEN_1; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_0; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_2; // @[Modules.scala 139:37:@39871.4]
  wire [22:0] _T_84; // @[Modules.scala 139:37:@39871.4]
  wire [7:0] _GEN_3; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_0; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_86; // @[Modules.scala 140:38:@39873.4]
  wire [7:0] _T_87; // @[Modules.scala 140:38:@39874.4]
  wire [7:0] _T_88; // @[Modules.scala 140:38:@39875.4]
  wire [8:0] _T_90; // @[Modules.scala 132:28:@39877.4]
  wire [7:0] _T_91; // @[Modules.scala 132:28:@39878.4]
  wire [7:0] c_x_1; // @[Modules.scala 132:28:@39879.4]
  wire [22:0] _GEN_4; // @[Modules.scala 137:32:@39881.4]
  wire [22:0] _T_94; // @[Modules.scala 137:32:@39881.4]
  wire [7:0] _GEN_5; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_1; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_6; // @[Modules.scala 139:37:@39883.4]
  wire [22:0] _T_96; // @[Modules.scala 139:37:@39883.4]
  wire [7:0] _GEN_7; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_1; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_98; // @[Modules.scala 140:38:@39885.4]
  wire [7:0] _T_99; // @[Modules.scala 140:38:@39886.4]
  wire [7:0] _T_100; // @[Modules.scala 140:38:@39887.4]
  wire [8:0] _T_102; // @[Modules.scala 132:28:@39889.4]
  wire [7:0] _T_103; // @[Modules.scala 132:28:@39890.4]
  wire [7:0] c_x_2; // @[Modules.scala 132:28:@39891.4]
  wire [22:0] _GEN_8; // @[Modules.scala 137:32:@39893.4]
  wire [22:0] _T_106; // @[Modules.scala 137:32:@39893.4]
  wire [7:0] _GEN_9; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_2; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_10; // @[Modules.scala 139:37:@39895.4]
  wire [22:0] _T_108; // @[Modules.scala 139:37:@39895.4]
  wire [7:0] _GEN_11; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_2; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_110; // @[Modules.scala 140:38:@39897.4]
  wire [7:0] _T_111; // @[Modules.scala 140:38:@39898.4]
  wire [7:0] _T_112; // @[Modules.scala 140:38:@39899.4]
  wire [8:0] _T_114; // @[Modules.scala 132:28:@39901.4]
  wire [7:0] _T_115; // @[Modules.scala 132:28:@39902.4]
  wire [7:0] c_x_3; // @[Modules.scala 132:28:@39903.4]
  wire [22:0] _GEN_12; // @[Modules.scala 137:32:@39905.4]
  wire [22:0] _T_118; // @[Modules.scala 137:32:@39905.4]
  wire [7:0] _GEN_13; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_3; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_14; // @[Modules.scala 139:37:@39907.4]
  wire [22:0] _T_120; // @[Modules.scala 139:37:@39907.4]
  wire [7:0] _GEN_15; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_3; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_122; // @[Modules.scala 140:38:@39909.4]
  wire [7:0] _T_123; // @[Modules.scala 140:38:@39910.4]
  wire [7:0] _T_124; // @[Modules.scala 140:38:@39911.4]
  wire [8:0] _T_126; // @[Modules.scala 132:28:@39913.4]
  wire [7:0] _T_127; // @[Modules.scala 132:28:@39914.4]
  wire [7:0] c_x_4; // @[Modules.scala 132:28:@39915.4]
  wire [22:0] _GEN_16; // @[Modules.scala 137:32:@39917.4]
  wire [22:0] _T_130; // @[Modules.scala 137:32:@39917.4]
  wire [7:0] _GEN_17; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_4; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_18; // @[Modules.scala 139:37:@39919.4]
  wire [22:0] _T_132; // @[Modules.scala 139:37:@39919.4]
  wire [7:0] _GEN_19; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_4; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_134; // @[Modules.scala 140:38:@39921.4]
  wire [7:0] _T_135; // @[Modules.scala 140:38:@39922.4]
  wire [7:0] _T_136; // @[Modules.scala 140:38:@39923.4]
  wire [8:0] _T_138; // @[Modules.scala 132:28:@39925.4]
  wire [7:0] _T_139; // @[Modules.scala 132:28:@39926.4]
  wire [7:0] c_x_5; // @[Modules.scala 132:28:@39927.4]
  wire [22:0] _GEN_20; // @[Modules.scala 137:32:@39929.4]
  wire [22:0] _T_142; // @[Modules.scala 137:32:@39929.4]
  wire [7:0] _GEN_21; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_5; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_22; // @[Modules.scala 139:37:@39931.4]
  wire [22:0] _T_144; // @[Modules.scala 139:37:@39931.4]
  wire [7:0] _GEN_23; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_5; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_146; // @[Modules.scala 140:38:@39933.4]
  wire [7:0] _T_147; // @[Modules.scala 140:38:@39934.4]
  wire [7:0] _T_148; // @[Modules.scala 140:38:@39935.4]
  wire [8:0] _T_150; // @[Modules.scala 132:28:@39937.4]
  wire [7:0] _T_151; // @[Modules.scala 132:28:@39938.4]
  wire [7:0] c_x_6; // @[Modules.scala 132:28:@39939.4]
  wire [22:0] _GEN_24; // @[Modules.scala 137:32:@39941.4]
  wire [22:0] _T_154; // @[Modules.scala 137:32:@39941.4]
  wire [7:0] _GEN_25; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_6; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_26; // @[Modules.scala 139:37:@39943.4]
  wire [22:0] _T_156; // @[Modules.scala 139:37:@39943.4]
  wire [7:0] _GEN_27; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_6; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_158; // @[Modules.scala 140:38:@39945.4]
  wire [7:0] _T_159; // @[Modules.scala 140:38:@39946.4]
  wire [7:0] _T_160; // @[Modules.scala 140:38:@39947.4]
  wire [8:0] _T_162; // @[Modules.scala 132:28:@39949.4]
  wire [7:0] _T_163; // @[Modules.scala 132:28:@39950.4]
  wire [7:0] c_x_7; // @[Modules.scala 132:28:@39951.4]
  wire [22:0] _GEN_28; // @[Modules.scala 137:32:@39953.4]
  wire [22:0] _T_166; // @[Modules.scala 137:32:@39953.4]
  wire [7:0] _GEN_29; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_7; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_30; // @[Modules.scala 139:37:@39955.4]
  wire [22:0] _T_168; // @[Modules.scala 139:37:@39955.4]
  wire [7:0] _GEN_31; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_7; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_170; // @[Modules.scala 140:38:@39957.4]
  wire [7:0] _T_171; // @[Modules.scala 140:38:@39958.4]
  wire [7:0] _T_172; // @[Modules.scala 140:38:@39959.4]
  wire [8:0] _T_174; // @[Modules.scala 132:28:@39961.4]
  wire [7:0] _T_175; // @[Modules.scala 132:28:@39962.4]
  wire [7:0] c_x_8; // @[Modules.scala 132:28:@39963.4]
  wire [22:0] _GEN_32; // @[Modules.scala 137:32:@39965.4]
  wire [22:0] _T_178; // @[Modules.scala 137:32:@39965.4]
  wire [7:0] _GEN_33; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_8; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_34; // @[Modules.scala 139:37:@39967.4]
  wire [22:0] _T_180; // @[Modules.scala 139:37:@39967.4]
  wire [7:0] _GEN_35; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_8; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_182; // @[Modules.scala 140:38:@39969.4]
  wire [7:0] _T_183; // @[Modules.scala 140:38:@39970.4]
  wire [7:0] _T_184; // @[Modules.scala 140:38:@39971.4]
  wire [8:0] _T_186; // @[Modules.scala 132:28:@39973.4]
  wire [7:0] _T_187; // @[Modules.scala 132:28:@39974.4]
  wire [7:0] c_x_9; // @[Modules.scala 132:28:@39975.4]
  wire [22:0] _GEN_36; // @[Modules.scala 137:32:@39977.4]
  wire [22:0] _T_190; // @[Modules.scala 137:32:@39977.4]
  wire [7:0] _GEN_37; // @[Modules.scala 129:21:@39863.4]
  wire [7:0] x_hat_9; // @[Modules.scala 129:21:@39863.4]
  wire [22:0] _GEN_38; // @[Modules.scala 139:37:@39979.4]
  wire [22:0] _T_192; // @[Modules.scala 139:37:@39979.4]
  wire [7:0] _GEN_39; // @[Modules.scala 130:28:@39864.4]
  wire [7:0] normed_x_hat_9; // @[Modules.scala 130:28:@39864.4]
  wire [8:0] _T_194; // @[Modules.scala 140:38:@39981.4]
  wire [7:0] _T_195; // @[Modules.scala 140:38:@39982.4]
  wire [7:0] _T_196; // @[Modules.scala 140:38:@39983.4]
  assign _T_78 = $signed(io_in_0) - $signed(8'sh0); // @[Modules.scala 132:28:@39865.4]
  assign _T_79 = _T_78[7:0]; // @[Modules.scala 132:28:@39866.4]
  assign c_x_0 = $signed(_T_79); // @[Modules.scala 132:28:@39867.4]
  assign _GEN_0 = {{15{c_x_0[7]}},c_x_0}; // @[Modules.scala 137:32:@39869.4]
  assign _T_82 = $signed(_GEN_0) << 4'h3; // @[Modules.scala 137:32:@39869.4]
  assign _GEN_1 = _T_82[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_0 = $signed(_GEN_1); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_2 = {{15{x_hat_0[7]}},x_hat_0}; // @[Modules.scala 139:37:@39871.4]
  assign _T_84 = $signed(_GEN_2) << 4'h2; // @[Modules.scala 139:37:@39871.4]
  assign _GEN_3 = _T_84[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_0 = $signed(_GEN_3); // @[Modules.scala 130:28:@39864.4]
  assign _T_86 = $signed(normed_x_hat_0) + $signed(-8'sh1); // @[Modules.scala 140:38:@39873.4]
  assign _T_87 = _T_86[7:0]; // @[Modules.scala 140:38:@39874.4]
  assign _T_88 = $signed(_T_87); // @[Modules.scala 140:38:@39875.4]
  assign _T_90 = $signed(io_in_1) - $signed(8'sh0); // @[Modules.scala 132:28:@39877.4]
  assign _T_91 = _T_90[7:0]; // @[Modules.scala 132:28:@39878.4]
  assign c_x_1 = $signed(_T_91); // @[Modules.scala 132:28:@39879.4]
  assign _GEN_4 = {{15{c_x_1[7]}},c_x_1}; // @[Modules.scala 137:32:@39881.4]
  assign _T_94 = $signed(_GEN_4) << 4'h3; // @[Modules.scala 137:32:@39881.4]
  assign _GEN_5 = _T_94[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_1 = $signed(_GEN_5); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_6 = {{15{x_hat_1[7]}},x_hat_1}; // @[Modules.scala 139:37:@39883.4]
  assign _T_96 = $signed(_GEN_6) << 4'h2; // @[Modules.scala 139:37:@39883.4]
  assign _GEN_7 = _T_96[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_1 = $signed(_GEN_7); // @[Modules.scala 130:28:@39864.4]
  assign _T_98 = $signed(normed_x_hat_1) + $signed(-8'sh1); // @[Modules.scala 140:38:@39885.4]
  assign _T_99 = _T_98[7:0]; // @[Modules.scala 140:38:@39886.4]
  assign _T_100 = $signed(_T_99); // @[Modules.scala 140:38:@39887.4]
  assign _T_102 = $signed(io_in_2) - $signed(8'sh0); // @[Modules.scala 132:28:@39889.4]
  assign _T_103 = _T_102[7:0]; // @[Modules.scala 132:28:@39890.4]
  assign c_x_2 = $signed(_T_103); // @[Modules.scala 132:28:@39891.4]
  assign _GEN_8 = {{15{c_x_2[7]}},c_x_2}; // @[Modules.scala 137:32:@39893.4]
  assign _T_106 = $signed(_GEN_8) << 4'h2; // @[Modules.scala 137:32:@39893.4]
  assign _GEN_9 = _T_106[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_2 = $signed(_GEN_9); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_10 = {{15{x_hat_2[7]}},x_hat_2}; // @[Modules.scala 139:37:@39895.4]
  assign _T_108 = $signed(_GEN_10) << 4'h1; // @[Modules.scala 139:37:@39895.4]
  assign _GEN_11 = _T_108[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_2 = $signed(_GEN_11); // @[Modules.scala 130:28:@39864.4]
  assign _T_110 = $signed(normed_x_hat_2) + $signed(8'sh1); // @[Modules.scala 140:38:@39897.4]
  assign _T_111 = _T_110[7:0]; // @[Modules.scala 140:38:@39898.4]
  assign _T_112 = $signed(_T_111); // @[Modules.scala 140:38:@39899.4]
  assign _T_114 = $signed(io_in_3) - $signed(8'sh0); // @[Modules.scala 132:28:@39901.4]
  assign _T_115 = _T_114[7:0]; // @[Modules.scala 132:28:@39902.4]
  assign c_x_3 = $signed(_T_115); // @[Modules.scala 132:28:@39903.4]
  assign _GEN_12 = {{15{c_x_3[7]}},c_x_3}; // @[Modules.scala 137:32:@39905.4]
  assign _T_118 = $signed(_GEN_12) << 4'h2; // @[Modules.scala 137:32:@39905.4]
  assign _GEN_13 = _T_118[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_3 = $signed(_GEN_13); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_14 = {{15{x_hat_3[7]}},x_hat_3}; // @[Modules.scala 139:37:@39907.4]
  assign _T_120 = $signed(_GEN_14) << 4'h1; // @[Modules.scala 139:37:@39907.4]
  assign _GEN_15 = _T_120[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_3 = $signed(_GEN_15); // @[Modules.scala 130:28:@39864.4]
  assign _T_122 = $signed(normed_x_hat_3) + $signed(8'sh1); // @[Modules.scala 140:38:@39909.4]
  assign _T_123 = _T_122[7:0]; // @[Modules.scala 140:38:@39910.4]
  assign _T_124 = $signed(_T_123); // @[Modules.scala 140:38:@39911.4]
  assign _T_126 = $signed(io_in_4) - $signed(8'sh1); // @[Modules.scala 132:28:@39913.4]
  assign _T_127 = _T_126[7:0]; // @[Modules.scala 132:28:@39914.4]
  assign c_x_4 = $signed(_T_127); // @[Modules.scala 132:28:@39915.4]
  assign _GEN_16 = {{15{c_x_4[7]}},c_x_4}; // @[Modules.scala 137:32:@39917.4]
  assign _T_130 = $signed(_GEN_16) << 4'h3; // @[Modules.scala 137:32:@39917.4]
  assign _GEN_17 = _T_130[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_4 = $signed(_GEN_17); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_18 = {{15{x_hat_4[7]}},x_hat_4}; // @[Modules.scala 139:37:@39919.4]
  assign _T_132 = $signed(_GEN_18) << 4'h1; // @[Modules.scala 139:37:@39919.4]
  assign _GEN_19 = _T_132[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_4 = $signed(_GEN_19); // @[Modules.scala 130:28:@39864.4]
  assign _T_134 = $signed(normed_x_hat_4) + $signed(8'sh0); // @[Modules.scala 140:38:@39921.4]
  assign _T_135 = _T_134[7:0]; // @[Modules.scala 140:38:@39922.4]
  assign _T_136 = $signed(_T_135); // @[Modules.scala 140:38:@39923.4]
  assign _T_138 = $signed(io_in_5) - $signed(8'sh0); // @[Modules.scala 132:28:@39925.4]
  assign _T_139 = _T_138[7:0]; // @[Modules.scala 132:28:@39926.4]
  assign c_x_5 = $signed(_T_139); // @[Modules.scala 132:28:@39927.4]
  assign _GEN_20 = {{15{c_x_5[7]}},c_x_5}; // @[Modules.scala 137:32:@39929.4]
  assign _T_142 = $signed(_GEN_20) << 4'h2; // @[Modules.scala 137:32:@39929.4]
  assign _GEN_21 = _T_142[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_5 = $signed(_GEN_21); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_22 = {{15{x_hat_5[7]}},x_hat_5}; // @[Modules.scala 139:37:@39931.4]
  assign _T_144 = $signed(_GEN_22) << 4'h1; // @[Modules.scala 139:37:@39931.4]
  assign _GEN_23 = _T_144[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_5 = $signed(_GEN_23); // @[Modules.scala 130:28:@39864.4]
  assign _T_146 = $signed(normed_x_hat_5) + $signed(8'sh1); // @[Modules.scala 140:38:@39933.4]
  assign _T_147 = _T_146[7:0]; // @[Modules.scala 140:38:@39934.4]
  assign _T_148 = $signed(_T_147); // @[Modules.scala 140:38:@39935.4]
  assign _T_150 = $signed(io_in_6) - $signed(8'sh0); // @[Modules.scala 132:28:@39937.4]
  assign _T_151 = _T_150[7:0]; // @[Modules.scala 132:28:@39938.4]
  assign c_x_6 = $signed(_T_151); // @[Modules.scala 132:28:@39939.4]
  assign _GEN_24 = {{15{c_x_6[7]}},c_x_6}; // @[Modules.scala 137:32:@39941.4]
  assign _T_154 = $signed(_GEN_24) << 4'h2; // @[Modules.scala 137:32:@39941.4]
  assign _GEN_25 = _T_154[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_6 = $signed(_GEN_25); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_26 = {{15{x_hat_6[7]}},x_hat_6}; // @[Modules.scala 139:37:@39943.4]
  assign _T_156 = $signed(_GEN_26) << 4'h1; // @[Modules.scala 139:37:@39943.4]
  assign _GEN_27 = _T_156[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_6 = $signed(_GEN_27); // @[Modules.scala 130:28:@39864.4]
  assign _T_158 = $signed(normed_x_hat_6) + $signed(-8'sh1); // @[Modules.scala 140:38:@39945.4]
  assign _T_159 = _T_158[7:0]; // @[Modules.scala 140:38:@39946.4]
  assign _T_160 = $signed(_T_159); // @[Modules.scala 140:38:@39947.4]
  assign _T_162 = $signed(io_in_7) - $signed(8'sh1); // @[Modules.scala 132:28:@39949.4]
  assign _T_163 = _T_162[7:0]; // @[Modules.scala 132:28:@39950.4]
  assign c_x_7 = $signed(_T_163); // @[Modules.scala 132:28:@39951.4]
  assign _GEN_28 = {{15{c_x_7[7]}},c_x_7}; // @[Modules.scala 137:32:@39953.4]
  assign _T_166 = $signed(_GEN_28) << 4'h3; // @[Modules.scala 137:32:@39953.4]
  assign _GEN_29 = _T_166[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_7 = $signed(_GEN_29); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_30 = {{15{x_hat_7[7]}},x_hat_7}; // @[Modules.scala 139:37:@39955.4]
  assign _T_168 = $signed(_GEN_30) << 4'h1; // @[Modules.scala 139:37:@39955.4]
  assign _GEN_31 = _T_168[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_7 = $signed(_GEN_31); // @[Modules.scala 130:28:@39864.4]
  assign _T_170 = $signed(normed_x_hat_7) + $signed(8'sh0); // @[Modules.scala 140:38:@39957.4]
  assign _T_171 = _T_170[7:0]; // @[Modules.scala 140:38:@39958.4]
  assign _T_172 = $signed(_T_171); // @[Modules.scala 140:38:@39959.4]
  assign _T_174 = $signed(io_in_8) - $signed(8'sh0); // @[Modules.scala 132:28:@39961.4]
  assign _T_175 = _T_174[7:0]; // @[Modules.scala 132:28:@39962.4]
  assign c_x_8 = $signed(_T_175); // @[Modules.scala 132:28:@39963.4]
  assign _GEN_32 = {{15{c_x_8[7]}},c_x_8}; // @[Modules.scala 137:32:@39965.4]
  assign _T_178 = $signed(_GEN_32) << 4'h2; // @[Modules.scala 137:32:@39965.4]
  assign _GEN_33 = _T_178[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_8 = $signed(_GEN_33); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_34 = {{15{x_hat_8[7]}},x_hat_8}; // @[Modules.scala 139:37:@39967.4]
  assign _T_180 = $signed(_GEN_34) << 4'h1; // @[Modules.scala 139:37:@39967.4]
  assign _GEN_35 = _T_180[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_8 = $signed(_GEN_35); // @[Modules.scala 130:28:@39864.4]
  assign _T_182 = $signed(normed_x_hat_8) + $signed(8'sh1); // @[Modules.scala 140:38:@39969.4]
  assign _T_183 = _T_182[7:0]; // @[Modules.scala 140:38:@39970.4]
  assign _T_184 = $signed(_T_183); // @[Modules.scala 140:38:@39971.4]
  assign _T_186 = $signed(io_in_9) - $signed(8'sh1); // @[Modules.scala 132:28:@39973.4]
  assign _T_187 = _T_186[7:0]; // @[Modules.scala 132:28:@39974.4]
  assign c_x_9 = $signed(_T_187); // @[Modules.scala 132:28:@39975.4]
  assign _GEN_36 = {{15{c_x_9[7]}},c_x_9}; // @[Modules.scala 137:32:@39977.4]
  assign _T_190 = $signed(_GEN_36) << 4'h3; // @[Modules.scala 137:32:@39977.4]
  assign _GEN_37 = _T_190[7:0]; // @[Modules.scala 129:21:@39863.4]
  assign x_hat_9 = $signed(_GEN_37); // @[Modules.scala 129:21:@39863.4]
  assign _GEN_38 = {{15{x_hat_9[7]}},x_hat_9}; // @[Modules.scala 139:37:@39979.4]
  assign _T_192 = $signed(_GEN_38) << 4'h1; // @[Modules.scala 139:37:@39979.4]
  assign _GEN_39 = _T_192[7:0]; // @[Modules.scala 130:28:@39864.4]
  assign normed_x_hat_9 = $signed(_GEN_39); // @[Modules.scala 130:28:@39864.4]
  assign _T_194 = $signed(normed_x_hat_9) + $signed(8'sh0); // @[Modules.scala 140:38:@39981.4]
  assign _T_195 = _T_194[7:0]; // @[Modules.scala 140:38:@39982.4]
  assign _T_196 = $signed(_T_195); // @[Modules.scala 140:38:@39983.4]
  assign io_out_0 = _T_88;
  assign io_out_1 = _T_100;
  assign io_out_2 = _T_112;
  assign io_out_3 = _T_124;
  assign io_out_4 = _T_136;
  assign io_out_5 = _T_148;
  assign io_out_6 = _T_160;
  assign io_out_7 = _T_172;
  assign io_out_8 = _T_184;
  assign io_out_9 = _T_196;
endmodule
module MLP_p( // @[:@39986.2]
  input        clock, // @[:@39987.4]
  input        reset, // @[:@39988.4]
  input  [4:0] io_in_0, // @[:@39989.4]
  input  [4:0] io_in_1, // @[:@39989.4]
  input  [4:0] io_in_2, // @[:@39989.4]
  input  [4:0] io_in_3, // @[:@39989.4]
  input  [4:0] io_in_4, // @[:@39989.4]
  input  [4:0] io_in_5, // @[:@39989.4]
  input  [4:0] io_in_6, // @[:@39989.4]
  input  [4:0] io_in_7, // @[:@39989.4]
  input  [4:0] io_in_8, // @[:@39989.4]
  input  [4:0] io_in_9, // @[:@39989.4]
  input  [4:0] io_in_10, // @[:@39989.4]
  input  [4:0] io_in_11, // @[:@39989.4]
  input  [4:0] io_in_12, // @[:@39989.4]
  input  [4:0] io_in_13, // @[:@39989.4]
  input  [4:0] io_in_14, // @[:@39989.4]
  input  [4:0] io_in_15, // @[:@39989.4]
  input  [4:0] io_in_16, // @[:@39989.4]
  input  [4:0] io_in_17, // @[:@39989.4]
  input  [4:0] io_in_18, // @[:@39989.4]
  input  [4:0] io_in_19, // @[:@39989.4]
  input  [4:0] io_in_20, // @[:@39989.4]
  input  [4:0] io_in_21, // @[:@39989.4]
  input  [4:0] io_in_22, // @[:@39989.4]
  input  [4:0] io_in_23, // @[:@39989.4]
  input  [4:0] io_in_24, // @[:@39989.4]
  input  [4:0] io_in_25, // @[:@39989.4]
  input  [4:0] io_in_26, // @[:@39989.4]
  input  [4:0] io_in_27, // @[:@39989.4]
  input  [4:0] io_in_28, // @[:@39989.4]
  input  [4:0] io_in_29, // @[:@39989.4]
  input  [4:0] io_in_30, // @[:@39989.4]
  input  [4:0] io_in_31, // @[:@39989.4]
  input  [4:0] io_in_32, // @[:@39989.4]
  input  [4:0] io_in_33, // @[:@39989.4]
  input  [4:0] io_in_34, // @[:@39989.4]
  input  [4:0] io_in_35, // @[:@39989.4]
  input  [4:0] io_in_36, // @[:@39989.4]
  input  [4:0] io_in_37, // @[:@39989.4]
  input  [4:0] io_in_38, // @[:@39989.4]
  input  [4:0] io_in_39, // @[:@39989.4]
  input  [4:0] io_in_40, // @[:@39989.4]
  input  [4:0] io_in_41, // @[:@39989.4]
  input  [4:0] io_in_42, // @[:@39989.4]
  input  [4:0] io_in_43, // @[:@39989.4]
  input  [4:0] io_in_44, // @[:@39989.4]
  input  [4:0] io_in_45, // @[:@39989.4]
  input  [4:0] io_in_46, // @[:@39989.4]
  input  [4:0] io_in_47, // @[:@39989.4]
  input  [4:0] io_in_48, // @[:@39989.4]
  input  [4:0] io_in_49, // @[:@39989.4]
  input  [4:0] io_in_50, // @[:@39989.4]
  input  [4:0] io_in_51, // @[:@39989.4]
  input  [4:0] io_in_52, // @[:@39989.4]
  input  [4:0] io_in_53, // @[:@39989.4]
  input  [4:0] io_in_54, // @[:@39989.4]
  input  [4:0] io_in_55, // @[:@39989.4]
  input  [4:0] io_in_56, // @[:@39989.4]
  input  [4:0] io_in_57, // @[:@39989.4]
  input  [4:0] io_in_58, // @[:@39989.4]
  input  [4:0] io_in_59, // @[:@39989.4]
  input  [4:0] io_in_60, // @[:@39989.4]
  input  [4:0] io_in_61, // @[:@39989.4]
  input  [4:0] io_in_62, // @[:@39989.4]
  input  [4:0] io_in_63, // @[:@39989.4]
  input  [4:0] io_in_64, // @[:@39989.4]
  input  [4:0] io_in_65, // @[:@39989.4]
  input  [4:0] io_in_66, // @[:@39989.4]
  input  [4:0] io_in_67, // @[:@39989.4]
  input  [4:0] io_in_68, // @[:@39989.4]
  input  [4:0] io_in_69, // @[:@39989.4]
  input  [4:0] io_in_70, // @[:@39989.4]
  input  [4:0] io_in_71, // @[:@39989.4]
  input  [4:0] io_in_72, // @[:@39989.4]
  input  [4:0] io_in_73, // @[:@39989.4]
  input  [4:0] io_in_74, // @[:@39989.4]
  input  [4:0] io_in_75, // @[:@39989.4]
  input  [4:0] io_in_76, // @[:@39989.4]
  input  [4:0] io_in_77, // @[:@39989.4]
  input  [4:0] io_in_78, // @[:@39989.4]
  input  [4:0] io_in_79, // @[:@39989.4]
  input  [4:0] io_in_80, // @[:@39989.4]
  input  [4:0] io_in_81, // @[:@39989.4]
  input  [4:0] io_in_82, // @[:@39989.4]
  input  [4:0] io_in_83, // @[:@39989.4]
  input  [4:0] io_in_84, // @[:@39989.4]
  input  [4:0] io_in_85, // @[:@39989.4]
  input  [4:0] io_in_86, // @[:@39989.4]
  input  [4:0] io_in_87, // @[:@39989.4]
  input  [4:0] io_in_88, // @[:@39989.4]
  input  [4:0] io_in_89, // @[:@39989.4]
  input  [4:0] io_in_90, // @[:@39989.4]
  input  [4:0] io_in_91, // @[:@39989.4]
  input  [4:0] io_in_92, // @[:@39989.4]
  input  [4:0] io_in_93, // @[:@39989.4]
  input  [4:0] io_in_94, // @[:@39989.4]
  input  [4:0] io_in_95, // @[:@39989.4]
  input  [4:0] io_in_96, // @[:@39989.4]
  input  [4:0] io_in_97, // @[:@39989.4]
  input  [4:0] io_in_98, // @[:@39989.4]
  input  [4:0] io_in_99, // @[:@39989.4]
  input  [4:0] io_in_100, // @[:@39989.4]
  input  [4:0] io_in_101, // @[:@39989.4]
  input  [4:0] io_in_102, // @[:@39989.4]
  input  [4:0] io_in_103, // @[:@39989.4]
  input  [4:0] io_in_104, // @[:@39989.4]
  input  [4:0] io_in_105, // @[:@39989.4]
  input  [4:0] io_in_106, // @[:@39989.4]
  input  [4:0] io_in_107, // @[:@39989.4]
  input  [4:0] io_in_108, // @[:@39989.4]
  input  [4:0] io_in_109, // @[:@39989.4]
  input  [4:0] io_in_110, // @[:@39989.4]
  input  [4:0] io_in_111, // @[:@39989.4]
  input  [4:0] io_in_112, // @[:@39989.4]
  input  [4:0] io_in_113, // @[:@39989.4]
  input  [4:0] io_in_114, // @[:@39989.4]
  input  [4:0] io_in_115, // @[:@39989.4]
  input  [4:0] io_in_116, // @[:@39989.4]
  input  [4:0] io_in_117, // @[:@39989.4]
  input  [4:0] io_in_118, // @[:@39989.4]
  input  [4:0] io_in_119, // @[:@39989.4]
  input  [4:0] io_in_120, // @[:@39989.4]
  input  [4:0] io_in_121, // @[:@39989.4]
  input  [4:0] io_in_122, // @[:@39989.4]
  input  [4:0] io_in_123, // @[:@39989.4]
  input  [4:0] io_in_124, // @[:@39989.4]
  input  [4:0] io_in_125, // @[:@39989.4]
  input  [4:0] io_in_126, // @[:@39989.4]
  input  [4:0] io_in_127, // @[:@39989.4]
  input  [4:0] io_in_128, // @[:@39989.4]
  input  [4:0] io_in_129, // @[:@39989.4]
  input  [4:0] io_in_130, // @[:@39989.4]
  input  [4:0] io_in_131, // @[:@39989.4]
  input  [4:0] io_in_132, // @[:@39989.4]
  input  [4:0] io_in_133, // @[:@39989.4]
  input  [4:0] io_in_134, // @[:@39989.4]
  input  [4:0] io_in_135, // @[:@39989.4]
  input  [4:0] io_in_136, // @[:@39989.4]
  input  [4:0] io_in_137, // @[:@39989.4]
  input  [4:0] io_in_138, // @[:@39989.4]
  input  [4:0] io_in_139, // @[:@39989.4]
  input  [4:0] io_in_140, // @[:@39989.4]
  input  [4:0] io_in_141, // @[:@39989.4]
  input  [4:0] io_in_142, // @[:@39989.4]
  input  [4:0] io_in_143, // @[:@39989.4]
  input  [4:0] io_in_144, // @[:@39989.4]
  input  [4:0] io_in_145, // @[:@39989.4]
  input  [4:0] io_in_146, // @[:@39989.4]
  input  [4:0] io_in_147, // @[:@39989.4]
  input  [4:0] io_in_148, // @[:@39989.4]
  input  [4:0] io_in_149, // @[:@39989.4]
  input  [4:0] io_in_150, // @[:@39989.4]
  input  [4:0] io_in_151, // @[:@39989.4]
  input  [4:0] io_in_152, // @[:@39989.4]
  input  [4:0] io_in_153, // @[:@39989.4]
  input  [4:0] io_in_154, // @[:@39989.4]
  input  [4:0] io_in_155, // @[:@39989.4]
  input  [4:0] io_in_156, // @[:@39989.4]
  input  [4:0] io_in_157, // @[:@39989.4]
  input  [4:0] io_in_158, // @[:@39989.4]
  input  [4:0] io_in_159, // @[:@39989.4]
  input  [4:0] io_in_160, // @[:@39989.4]
  input  [4:0] io_in_161, // @[:@39989.4]
  input  [4:0] io_in_162, // @[:@39989.4]
  input  [4:0] io_in_163, // @[:@39989.4]
  input  [4:0] io_in_164, // @[:@39989.4]
  input  [4:0] io_in_165, // @[:@39989.4]
  input  [4:0] io_in_166, // @[:@39989.4]
  input  [4:0] io_in_167, // @[:@39989.4]
  input  [4:0] io_in_168, // @[:@39989.4]
  input  [4:0] io_in_169, // @[:@39989.4]
  input  [4:0] io_in_170, // @[:@39989.4]
  input  [4:0] io_in_171, // @[:@39989.4]
  input  [4:0] io_in_172, // @[:@39989.4]
  input  [4:0] io_in_173, // @[:@39989.4]
  input  [4:0] io_in_174, // @[:@39989.4]
  input  [4:0] io_in_175, // @[:@39989.4]
  input  [4:0] io_in_176, // @[:@39989.4]
  input  [4:0] io_in_177, // @[:@39989.4]
  input  [4:0] io_in_178, // @[:@39989.4]
  input  [4:0] io_in_179, // @[:@39989.4]
  input  [4:0] io_in_180, // @[:@39989.4]
  input  [4:0] io_in_181, // @[:@39989.4]
  input  [4:0] io_in_182, // @[:@39989.4]
  input  [4:0] io_in_183, // @[:@39989.4]
  input  [4:0] io_in_184, // @[:@39989.4]
  input  [4:0] io_in_185, // @[:@39989.4]
  input  [4:0] io_in_186, // @[:@39989.4]
  input  [4:0] io_in_187, // @[:@39989.4]
  input  [4:0] io_in_188, // @[:@39989.4]
  input  [4:0] io_in_189, // @[:@39989.4]
  input  [4:0] io_in_190, // @[:@39989.4]
  input  [4:0] io_in_191, // @[:@39989.4]
  input  [4:0] io_in_192, // @[:@39989.4]
  input  [4:0] io_in_193, // @[:@39989.4]
  input  [4:0] io_in_194, // @[:@39989.4]
  input  [4:0] io_in_195, // @[:@39989.4]
  input  [4:0] io_in_196, // @[:@39989.4]
  input  [4:0] io_in_197, // @[:@39989.4]
  input  [4:0] io_in_198, // @[:@39989.4]
  input  [4:0] io_in_199, // @[:@39989.4]
  input  [4:0] io_in_200, // @[:@39989.4]
  input  [4:0] io_in_201, // @[:@39989.4]
  input  [4:0] io_in_202, // @[:@39989.4]
  input  [4:0] io_in_203, // @[:@39989.4]
  input  [4:0] io_in_204, // @[:@39989.4]
  input  [4:0] io_in_205, // @[:@39989.4]
  input  [4:0] io_in_206, // @[:@39989.4]
  input  [4:0] io_in_207, // @[:@39989.4]
  input  [4:0] io_in_208, // @[:@39989.4]
  input  [4:0] io_in_209, // @[:@39989.4]
  input  [4:0] io_in_210, // @[:@39989.4]
  input  [4:0] io_in_211, // @[:@39989.4]
  input  [4:0] io_in_212, // @[:@39989.4]
  input  [4:0] io_in_213, // @[:@39989.4]
  input  [4:0] io_in_214, // @[:@39989.4]
  input  [4:0] io_in_215, // @[:@39989.4]
  input  [4:0] io_in_216, // @[:@39989.4]
  input  [4:0] io_in_217, // @[:@39989.4]
  input  [4:0] io_in_218, // @[:@39989.4]
  input  [4:0] io_in_219, // @[:@39989.4]
  input  [4:0] io_in_220, // @[:@39989.4]
  input  [4:0] io_in_221, // @[:@39989.4]
  input  [4:0] io_in_222, // @[:@39989.4]
  input  [4:0] io_in_223, // @[:@39989.4]
  input  [4:0] io_in_224, // @[:@39989.4]
  input  [4:0] io_in_225, // @[:@39989.4]
  input  [4:0] io_in_226, // @[:@39989.4]
  input  [4:0] io_in_227, // @[:@39989.4]
  input  [4:0] io_in_228, // @[:@39989.4]
  input  [4:0] io_in_229, // @[:@39989.4]
  input  [4:0] io_in_230, // @[:@39989.4]
  input  [4:0] io_in_231, // @[:@39989.4]
  input  [4:0] io_in_232, // @[:@39989.4]
  input  [4:0] io_in_233, // @[:@39989.4]
  input  [4:0] io_in_234, // @[:@39989.4]
  input  [4:0] io_in_235, // @[:@39989.4]
  input  [4:0] io_in_236, // @[:@39989.4]
  input  [4:0] io_in_237, // @[:@39989.4]
  input  [4:0] io_in_238, // @[:@39989.4]
  input  [4:0] io_in_239, // @[:@39989.4]
  input  [4:0] io_in_240, // @[:@39989.4]
  input  [4:0] io_in_241, // @[:@39989.4]
  input  [4:0] io_in_242, // @[:@39989.4]
  input  [4:0] io_in_243, // @[:@39989.4]
  input  [4:0] io_in_244, // @[:@39989.4]
  input  [4:0] io_in_245, // @[:@39989.4]
  input  [4:0] io_in_246, // @[:@39989.4]
  input  [4:0] io_in_247, // @[:@39989.4]
  input  [4:0] io_in_248, // @[:@39989.4]
  input  [4:0] io_in_249, // @[:@39989.4]
  input  [4:0] io_in_250, // @[:@39989.4]
  input  [4:0] io_in_251, // @[:@39989.4]
  input  [4:0] io_in_252, // @[:@39989.4]
  input  [4:0] io_in_253, // @[:@39989.4]
  input  [4:0] io_in_254, // @[:@39989.4]
  input  [4:0] io_in_255, // @[:@39989.4]
  input  [4:0] io_in_256, // @[:@39989.4]
  input  [4:0] io_in_257, // @[:@39989.4]
  input  [4:0] io_in_258, // @[:@39989.4]
  input  [4:0] io_in_259, // @[:@39989.4]
  input  [4:0] io_in_260, // @[:@39989.4]
  input  [4:0] io_in_261, // @[:@39989.4]
  input  [4:0] io_in_262, // @[:@39989.4]
  input  [4:0] io_in_263, // @[:@39989.4]
  input  [4:0] io_in_264, // @[:@39989.4]
  input  [4:0] io_in_265, // @[:@39989.4]
  input  [4:0] io_in_266, // @[:@39989.4]
  input  [4:0] io_in_267, // @[:@39989.4]
  input  [4:0] io_in_268, // @[:@39989.4]
  input  [4:0] io_in_269, // @[:@39989.4]
  input  [4:0] io_in_270, // @[:@39989.4]
  input  [4:0] io_in_271, // @[:@39989.4]
  input  [4:0] io_in_272, // @[:@39989.4]
  input  [4:0] io_in_273, // @[:@39989.4]
  input  [4:0] io_in_274, // @[:@39989.4]
  input  [4:0] io_in_275, // @[:@39989.4]
  input  [4:0] io_in_276, // @[:@39989.4]
  input  [4:0] io_in_277, // @[:@39989.4]
  input  [4:0] io_in_278, // @[:@39989.4]
  input  [4:0] io_in_279, // @[:@39989.4]
  input  [4:0] io_in_280, // @[:@39989.4]
  input  [4:0] io_in_281, // @[:@39989.4]
  input  [4:0] io_in_282, // @[:@39989.4]
  input  [4:0] io_in_283, // @[:@39989.4]
  input  [4:0] io_in_284, // @[:@39989.4]
  input  [4:0] io_in_285, // @[:@39989.4]
  input  [4:0] io_in_286, // @[:@39989.4]
  input  [4:0] io_in_287, // @[:@39989.4]
  input  [4:0] io_in_288, // @[:@39989.4]
  input  [4:0] io_in_289, // @[:@39989.4]
  input  [4:0] io_in_290, // @[:@39989.4]
  input  [4:0] io_in_291, // @[:@39989.4]
  input  [4:0] io_in_292, // @[:@39989.4]
  input  [4:0] io_in_293, // @[:@39989.4]
  input  [4:0] io_in_294, // @[:@39989.4]
  input  [4:0] io_in_295, // @[:@39989.4]
  input  [4:0] io_in_296, // @[:@39989.4]
  input  [4:0] io_in_297, // @[:@39989.4]
  input  [4:0] io_in_298, // @[:@39989.4]
  input  [4:0] io_in_299, // @[:@39989.4]
  input  [4:0] io_in_300, // @[:@39989.4]
  input  [4:0] io_in_301, // @[:@39989.4]
  input  [4:0] io_in_302, // @[:@39989.4]
  input  [4:0] io_in_303, // @[:@39989.4]
  input  [4:0] io_in_304, // @[:@39989.4]
  input  [4:0] io_in_305, // @[:@39989.4]
  input  [4:0] io_in_306, // @[:@39989.4]
  input  [4:0] io_in_307, // @[:@39989.4]
  input  [4:0] io_in_308, // @[:@39989.4]
  input  [4:0] io_in_309, // @[:@39989.4]
  input  [4:0] io_in_310, // @[:@39989.4]
  input  [4:0] io_in_311, // @[:@39989.4]
  input  [4:0] io_in_312, // @[:@39989.4]
  input  [4:0] io_in_313, // @[:@39989.4]
  input  [4:0] io_in_314, // @[:@39989.4]
  input  [4:0] io_in_315, // @[:@39989.4]
  input  [4:0] io_in_316, // @[:@39989.4]
  input  [4:0] io_in_317, // @[:@39989.4]
  input  [4:0] io_in_318, // @[:@39989.4]
  input  [4:0] io_in_319, // @[:@39989.4]
  input  [4:0] io_in_320, // @[:@39989.4]
  input  [4:0] io_in_321, // @[:@39989.4]
  input  [4:0] io_in_322, // @[:@39989.4]
  input  [4:0] io_in_323, // @[:@39989.4]
  input  [4:0] io_in_324, // @[:@39989.4]
  input  [4:0] io_in_325, // @[:@39989.4]
  input  [4:0] io_in_326, // @[:@39989.4]
  input  [4:0] io_in_327, // @[:@39989.4]
  input  [4:0] io_in_328, // @[:@39989.4]
  input  [4:0] io_in_329, // @[:@39989.4]
  input  [4:0] io_in_330, // @[:@39989.4]
  input  [4:0] io_in_331, // @[:@39989.4]
  input  [4:0] io_in_332, // @[:@39989.4]
  input  [4:0] io_in_333, // @[:@39989.4]
  input  [4:0] io_in_334, // @[:@39989.4]
  input  [4:0] io_in_335, // @[:@39989.4]
  input  [4:0] io_in_336, // @[:@39989.4]
  input  [4:0] io_in_337, // @[:@39989.4]
  input  [4:0] io_in_338, // @[:@39989.4]
  input  [4:0] io_in_339, // @[:@39989.4]
  input  [4:0] io_in_340, // @[:@39989.4]
  input  [4:0] io_in_341, // @[:@39989.4]
  input  [4:0] io_in_342, // @[:@39989.4]
  input  [4:0] io_in_343, // @[:@39989.4]
  input  [4:0] io_in_344, // @[:@39989.4]
  input  [4:0] io_in_345, // @[:@39989.4]
  input  [4:0] io_in_346, // @[:@39989.4]
  input  [4:0] io_in_347, // @[:@39989.4]
  input  [4:0] io_in_348, // @[:@39989.4]
  input  [4:0] io_in_349, // @[:@39989.4]
  input  [4:0] io_in_350, // @[:@39989.4]
  input  [4:0] io_in_351, // @[:@39989.4]
  input  [4:0] io_in_352, // @[:@39989.4]
  input  [4:0] io_in_353, // @[:@39989.4]
  input  [4:0] io_in_354, // @[:@39989.4]
  input  [4:0] io_in_355, // @[:@39989.4]
  input  [4:0] io_in_356, // @[:@39989.4]
  input  [4:0] io_in_357, // @[:@39989.4]
  input  [4:0] io_in_358, // @[:@39989.4]
  input  [4:0] io_in_359, // @[:@39989.4]
  input  [4:0] io_in_360, // @[:@39989.4]
  input  [4:0] io_in_361, // @[:@39989.4]
  input  [4:0] io_in_362, // @[:@39989.4]
  input  [4:0] io_in_363, // @[:@39989.4]
  input  [4:0] io_in_364, // @[:@39989.4]
  input  [4:0] io_in_365, // @[:@39989.4]
  input  [4:0] io_in_366, // @[:@39989.4]
  input  [4:0] io_in_367, // @[:@39989.4]
  input  [4:0] io_in_368, // @[:@39989.4]
  input  [4:0] io_in_369, // @[:@39989.4]
  input  [4:0] io_in_370, // @[:@39989.4]
  input  [4:0] io_in_371, // @[:@39989.4]
  input  [4:0] io_in_372, // @[:@39989.4]
  input  [4:0] io_in_373, // @[:@39989.4]
  input  [4:0] io_in_374, // @[:@39989.4]
  input  [4:0] io_in_375, // @[:@39989.4]
  input  [4:0] io_in_376, // @[:@39989.4]
  input  [4:0] io_in_377, // @[:@39989.4]
  input  [4:0] io_in_378, // @[:@39989.4]
  input  [4:0] io_in_379, // @[:@39989.4]
  input  [4:0] io_in_380, // @[:@39989.4]
  input  [4:0] io_in_381, // @[:@39989.4]
  input  [4:0] io_in_382, // @[:@39989.4]
  input  [4:0] io_in_383, // @[:@39989.4]
  input  [4:0] io_in_384, // @[:@39989.4]
  input  [4:0] io_in_385, // @[:@39989.4]
  input  [4:0] io_in_386, // @[:@39989.4]
  input  [4:0] io_in_387, // @[:@39989.4]
  input  [4:0] io_in_388, // @[:@39989.4]
  input  [4:0] io_in_389, // @[:@39989.4]
  input  [4:0] io_in_390, // @[:@39989.4]
  input  [4:0] io_in_391, // @[:@39989.4]
  input  [4:0] io_in_392, // @[:@39989.4]
  input  [4:0] io_in_393, // @[:@39989.4]
  input  [4:0] io_in_394, // @[:@39989.4]
  input  [4:0] io_in_395, // @[:@39989.4]
  input  [4:0] io_in_396, // @[:@39989.4]
  input  [4:0] io_in_397, // @[:@39989.4]
  input  [4:0] io_in_398, // @[:@39989.4]
  input  [4:0] io_in_399, // @[:@39989.4]
  input  [4:0] io_in_400, // @[:@39989.4]
  input  [4:0] io_in_401, // @[:@39989.4]
  input  [4:0] io_in_402, // @[:@39989.4]
  input  [4:0] io_in_403, // @[:@39989.4]
  input  [4:0] io_in_404, // @[:@39989.4]
  input  [4:0] io_in_405, // @[:@39989.4]
  input  [4:0] io_in_406, // @[:@39989.4]
  input  [4:0] io_in_407, // @[:@39989.4]
  input  [4:0] io_in_408, // @[:@39989.4]
  input  [4:0] io_in_409, // @[:@39989.4]
  input  [4:0] io_in_410, // @[:@39989.4]
  input  [4:0] io_in_411, // @[:@39989.4]
  input  [4:0] io_in_412, // @[:@39989.4]
  input  [4:0] io_in_413, // @[:@39989.4]
  input  [4:0] io_in_414, // @[:@39989.4]
  input  [4:0] io_in_415, // @[:@39989.4]
  input  [4:0] io_in_416, // @[:@39989.4]
  input  [4:0] io_in_417, // @[:@39989.4]
  input  [4:0] io_in_418, // @[:@39989.4]
  input  [4:0] io_in_419, // @[:@39989.4]
  input  [4:0] io_in_420, // @[:@39989.4]
  input  [4:0] io_in_421, // @[:@39989.4]
  input  [4:0] io_in_422, // @[:@39989.4]
  input  [4:0] io_in_423, // @[:@39989.4]
  input  [4:0] io_in_424, // @[:@39989.4]
  input  [4:0] io_in_425, // @[:@39989.4]
  input  [4:0] io_in_426, // @[:@39989.4]
  input  [4:0] io_in_427, // @[:@39989.4]
  input  [4:0] io_in_428, // @[:@39989.4]
  input  [4:0] io_in_429, // @[:@39989.4]
  input  [4:0] io_in_430, // @[:@39989.4]
  input  [4:0] io_in_431, // @[:@39989.4]
  input  [4:0] io_in_432, // @[:@39989.4]
  input  [4:0] io_in_433, // @[:@39989.4]
  input  [4:0] io_in_434, // @[:@39989.4]
  input  [4:0] io_in_435, // @[:@39989.4]
  input  [4:0] io_in_436, // @[:@39989.4]
  input  [4:0] io_in_437, // @[:@39989.4]
  input  [4:0] io_in_438, // @[:@39989.4]
  input  [4:0] io_in_439, // @[:@39989.4]
  input  [4:0] io_in_440, // @[:@39989.4]
  input  [4:0] io_in_441, // @[:@39989.4]
  input  [4:0] io_in_442, // @[:@39989.4]
  input  [4:0] io_in_443, // @[:@39989.4]
  input  [4:0] io_in_444, // @[:@39989.4]
  input  [4:0] io_in_445, // @[:@39989.4]
  input  [4:0] io_in_446, // @[:@39989.4]
  input  [4:0] io_in_447, // @[:@39989.4]
  input  [4:0] io_in_448, // @[:@39989.4]
  input  [4:0] io_in_449, // @[:@39989.4]
  input  [4:0] io_in_450, // @[:@39989.4]
  input  [4:0] io_in_451, // @[:@39989.4]
  input  [4:0] io_in_452, // @[:@39989.4]
  input  [4:0] io_in_453, // @[:@39989.4]
  input  [4:0] io_in_454, // @[:@39989.4]
  input  [4:0] io_in_455, // @[:@39989.4]
  input  [4:0] io_in_456, // @[:@39989.4]
  input  [4:0] io_in_457, // @[:@39989.4]
  input  [4:0] io_in_458, // @[:@39989.4]
  input  [4:0] io_in_459, // @[:@39989.4]
  input  [4:0] io_in_460, // @[:@39989.4]
  input  [4:0] io_in_461, // @[:@39989.4]
  input  [4:0] io_in_462, // @[:@39989.4]
  input  [4:0] io_in_463, // @[:@39989.4]
  input  [4:0] io_in_464, // @[:@39989.4]
  input  [4:0] io_in_465, // @[:@39989.4]
  input  [4:0] io_in_466, // @[:@39989.4]
  input  [4:0] io_in_467, // @[:@39989.4]
  input  [4:0] io_in_468, // @[:@39989.4]
  input  [4:0] io_in_469, // @[:@39989.4]
  input  [4:0] io_in_470, // @[:@39989.4]
  input  [4:0] io_in_471, // @[:@39989.4]
  input  [4:0] io_in_472, // @[:@39989.4]
  input  [4:0] io_in_473, // @[:@39989.4]
  input  [4:0] io_in_474, // @[:@39989.4]
  input  [4:0] io_in_475, // @[:@39989.4]
  input  [4:0] io_in_476, // @[:@39989.4]
  input  [4:0] io_in_477, // @[:@39989.4]
  input  [4:0] io_in_478, // @[:@39989.4]
  input  [4:0] io_in_479, // @[:@39989.4]
  input  [4:0] io_in_480, // @[:@39989.4]
  input  [4:0] io_in_481, // @[:@39989.4]
  input  [4:0] io_in_482, // @[:@39989.4]
  input  [4:0] io_in_483, // @[:@39989.4]
  input  [4:0] io_in_484, // @[:@39989.4]
  input  [4:0] io_in_485, // @[:@39989.4]
  input  [4:0] io_in_486, // @[:@39989.4]
  input  [4:0] io_in_487, // @[:@39989.4]
  input  [4:0] io_in_488, // @[:@39989.4]
  input  [4:0] io_in_489, // @[:@39989.4]
  input  [4:0] io_in_490, // @[:@39989.4]
  input  [4:0] io_in_491, // @[:@39989.4]
  input  [4:0] io_in_492, // @[:@39989.4]
  input  [4:0] io_in_493, // @[:@39989.4]
  input  [4:0] io_in_494, // @[:@39989.4]
  input  [4:0] io_in_495, // @[:@39989.4]
  input  [4:0] io_in_496, // @[:@39989.4]
  input  [4:0] io_in_497, // @[:@39989.4]
  input  [4:0] io_in_498, // @[:@39989.4]
  input  [4:0] io_in_499, // @[:@39989.4]
  input  [4:0] io_in_500, // @[:@39989.4]
  input  [4:0] io_in_501, // @[:@39989.4]
  input  [4:0] io_in_502, // @[:@39989.4]
  input  [4:0] io_in_503, // @[:@39989.4]
  input  [4:0] io_in_504, // @[:@39989.4]
  input  [4:0] io_in_505, // @[:@39989.4]
  input  [4:0] io_in_506, // @[:@39989.4]
  input  [4:0] io_in_507, // @[:@39989.4]
  input  [4:0] io_in_508, // @[:@39989.4]
  input  [4:0] io_in_509, // @[:@39989.4]
  input  [4:0] io_in_510, // @[:@39989.4]
  input  [4:0] io_in_511, // @[:@39989.4]
  input  [4:0] io_in_512, // @[:@39989.4]
  input  [4:0] io_in_513, // @[:@39989.4]
  input  [4:0] io_in_514, // @[:@39989.4]
  input  [4:0] io_in_515, // @[:@39989.4]
  input  [4:0] io_in_516, // @[:@39989.4]
  input  [4:0] io_in_517, // @[:@39989.4]
  input  [4:0] io_in_518, // @[:@39989.4]
  input  [4:0] io_in_519, // @[:@39989.4]
  input  [4:0] io_in_520, // @[:@39989.4]
  input  [4:0] io_in_521, // @[:@39989.4]
  input  [4:0] io_in_522, // @[:@39989.4]
  input  [4:0] io_in_523, // @[:@39989.4]
  input  [4:0] io_in_524, // @[:@39989.4]
  input  [4:0] io_in_525, // @[:@39989.4]
  input  [4:0] io_in_526, // @[:@39989.4]
  input  [4:0] io_in_527, // @[:@39989.4]
  input  [4:0] io_in_528, // @[:@39989.4]
  input  [4:0] io_in_529, // @[:@39989.4]
  input  [4:0] io_in_530, // @[:@39989.4]
  input  [4:0] io_in_531, // @[:@39989.4]
  input  [4:0] io_in_532, // @[:@39989.4]
  input  [4:0] io_in_533, // @[:@39989.4]
  input  [4:0] io_in_534, // @[:@39989.4]
  input  [4:0] io_in_535, // @[:@39989.4]
  input  [4:0] io_in_536, // @[:@39989.4]
  input  [4:0] io_in_537, // @[:@39989.4]
  input  [4:0] io_in_538, // @[:@39989.4]
  input  [4:0] io_in_539, // @[:@39989.4]
  input  [4:0] io_in_540, // @[:@39989.4]
  input  [4:0] io_in_541, // @[:@39989.4]
  input  [4:0] io_in_542, // @[:@39989.4]
  input  [4:0] io_in_543, // @[:@39989.4]
  input  [4:0] io_in_544, // @[:@39989.4]
  input  [4:0] io_in_545, // @[:@39989.4]
  input  [4:0] io_in_546, // @[:@39989.4]
  input  [4:0] io_in_547, // @[:@39989.4]
  input  [4:0] io_in_548, // @[:@39989.4]
  input  [4:0] io_in_549, // @[:@39989.4]
  input  [4:0] io_in_550, // @[:@39989.4]
  input  [4:0] io_in_551, // @[:@39989.4]
  input  [4:0] io_in_552, // @[:@39989.4]
  input  [4:0] io_in_553, // @[:@39989.4]
  input  [4:0] io_in_554, // @[:@39989.4]
  input  [4:0] io_in_555, // @[:@39989.4]
  input  [4:0] io_in_556, // @[:@39989.4]
  input  [4:0] io_in_557, // @[:@39989.4]
  input  [4:0] io_in_558, // @[:@39989.4]
  input  [4:0] io_in_559, // @[:@39989.4]
  input  [4:0] io_in_560, // @[:@39989.4]
  input  [4:0] io_in_561, // @[:@39989.4]
  input  [4:0] io_in_562, // @[:@39989.4]
  input  [4:0] io_in_563, // @[:@39989.4]
  input  [4:0] io_in_564, // @[:@39989.4]
  input  [4:0] io_in_565, // @[:@39989.4]
  input  [4:0] io_in_566, // @[:@39989.4]
  input  [4:0] io_in_567, // @[:@39989.4]
  input  [4:0] io_in_568, // @[:@39989.4]
  input  [4:0] io_in_569, // @[:@39989.4]
  input  [4:0] io_in_570, // @[:@39989.4]
  input  [4:0] io_in_571, // @[:@39989.4]
  input  [4:0] io_in_572, // @[:@39989.4]
  input  [4:0] io_in_573, // @[:@39989.4]
  input  [4:0] io_in_574, // @[:@39989.4]
  input  [4:0] io_in_575, // @[:@39989.4]
  input  [4:0] io_in_576, // @[:@39989.4]
  input  [4:0] io_in_577, // @[:@39989.4]
  input  [4:0] io_in_578, // @[:@39989.4]
  input  [4:0] io_in_579, // @[:@39989.4]
  input  [4:0] io_in_580, // @[:@39989.4]
  input  [4:0] io_in_581, // @[:@39989.4]
  input  [4:0] io_in_582, // @[:@39989.4]
  input  [4:0] io_in_583, // @[:@39989.4]
  input  [4:0] io_in_584, // @[:@39989.4]
  input  [4:0] io_in_585, // @[:@39989.4]
  input  [4:0] io_in_586, // @[:@39989.4]
  input  [4:0] io_in_587, // @[:@39989.4]
  input  [4:0] io_in_588, // @[:@39989.4]
  input  [4:0] io_in_589, // @[:@39989.4]
  input  [4:0] io_in_590, // @[:@39989.4]
  input  [4:0] io_in_591, // @[:@39989.4]
  input  [4:0] io_in_592, // @[:@39989.4]
  input  [4:0] io_in_593, // @[:@39989.4]
  input  [4:0] io_in_594, // @[:@39989.4]
  input  [4:0] io_in_595, // @[:@39989.4]
  input  [4:0] io_in_596, // @[:@39989.4]
  input  [4:0] io_in_597, // @[:@39989.4]
  input  [4:0] io_in_598, // @[:@39989.4]
  input  [4:0] io_in_599, // @[:@39989.4]
  input  [4:0] io_in_600, // @[:@39989.4]
  input  [4:0] io_in_601, // @[:@39989.4]
  input  [4:0] io_in_602, // @[:@39989.4]
  input  [4:0] io_in_603, // @[:@39989.4]
  input  [4:0] io_in_604, // @[:@39989.4]
  input  [4:0] io_in_605, // @[:@39989.4]
  input  [4:0] io_in_606, // @[:@39989.4]
  input  [4:0] io_in_607, // @[:@39989.4]
  input  [4:0] io_in_608, // @[:@39989.4]
  input  [4:0] io_in_609, // @[:@39989.4]
  input  [4:0] io_in_610, // @[:@39989.4]
  input  [4:0] io_in_611, // @[:@39989.4]
  input  [4:0] io_in_612, // @[:@39989.4]
  input  [4:0] io_in_613, // @[:@39989.4]
  input  [4:0] io_in_614, // @[:@39989.4]
  input  [4:0] io_in_615, // @[:@39989.4]
  input  [4:0] io_in_616, // @[:@39989.4]
  input  [4:0] io_in_617, // @[:@39989.4]
  input  [4:0] io_in_618, // @[:@39989.4]
  input  [4:0] io_in_619, // @[:@39989.4]
  input  [4:0] io_in_620, // @[:@39989.4]
  input  [4:0] io_in_621, // @[:@39989.4]
  input  [4:0] io_in_622, // @[:@39989.4]
  input  [4:0] io_in_623, // @[:@39989.4]
  input  [4:0] io_in_624, // @[:@39989.4]
  input  [4:0] io_in_625, // @[:@39989.4]
  input  [4:0] io_in_626, // @[:@39989.4]
  input  [4:0] io_in_627, // @[:@39989.4]
  input  [4:0] io_in_628, // @[:@39989.4]
  input  [4:0] io_in_629, // @[:@39989.4]
  input  [4:0] io_in_630, // @[:@39989.4]
  input  [4:0] io_in_631, // @[:@39989.4]
  input  [4:0] io_in_632, // @[:@39989.4]
  input  [4:0] io_in_633, // @[:@39989.4]
  input  [4:0] io_in_634, // @[:@39989.4]
  input  [4:0] io_in_635, // @[:@39989.4]
  input  [4:0] io_in_636, // @[:@39989.4]
  input  [4:0] io_in_637, // @[:@39989.4]
  input  [4:0] io_in_638, // @[:@39989.4]
  input  [4:0] io_in_639, // @[:@39989.4]
  input  [4:0] io_in_640, // @[:@39989.4]
  input  [4:0] io_in_641, // @[:@39989.4]
  input  [4:0] io_in_642, // @[:@39989.4]
  input  [4:0] io_in_643, // @[:@39989.4]
  input  [4:0] io_in_644, // @[:@39989.4]
  input  [4:0] io_in_645, // @[:@39989.4]
  input  [4:0] io_in_646, // @[:@39989.4]
  input  [4:0] io_in_647, // @[:@39989.4]
  input  [4:0] io_in_648, // @[:@39989.4]
  input  [4:0] io_in_649, // @[:@39989.4]
  input  [4:0] io_in_650, // @[:@39989.4]
  input  [4:0] io_in_651, // @[:@39989.4]
  input  [4:0] io_in_652, // @[:@39989.4]
  input  [4:0] io_in_653, // @[:@39989.4]
  input  [4:0] io_in_654, // @[:@39989.4]
  input  [4:0] io_in_655, // @[:@39989.4]
  input  [4:0] io_in_656, // @[:@39989.4]
  input  [4:0] io_in_657, // @[:@39989.4]
  input  [4:0] io_in_658, // @[:@39989.4]
  input  [4:0] io_in_659, // @[:@39989.4]
  input  [4:0] io_in_660, // @[:@39989.4]
  input  [4:0] io_in_661, // @[:@39989.4]
  input  [4:0] io_in_662, // @[:@39989.4]
  input  [4:0] io_in_663, // @[:@39989.4]
  input  [4:0] io_in_664, // @[:@39989.4]
  input  [4:0] io_in_665, // @[:@39989.4]
  input  [4:0] io_in_666, // @[:@39989.4]
  input  [4:0] io_in_667, // @[:@39989.4]
  input  [4:0] io_in_668, // @[:@39989.4]
  input  [4:0] io_in_669, // @[:@39989.4]
  input  [4:0] io_in_670, // @[:@39989.4]
  input  [4:0] io_in_671, // @[:@39989.4]
  input  [4:0] io_in_672, // @[:@39989.4]
  input  [4:0] io_in_673, // @[:@39989.4]
  input  [4:0] io_in_674, // @[:@39989.4]
  input  [4:0] io_in_675, // @[:@39989.4]
  input  [4:0] io_in_676, // @[:@39989.4]
  input  [4:0] io_in_677, // @[:@39989.4]
  input  [4:0] io_in_678, // @[:@39989.4]
  input  [4:0] io_in_679, // @[:@39989.4]
  input  [4:0] io_in_680, // @[:@39989.4]
  input  [4:0] io_in_681, // @[:@39989.4]
  input  [4:0] io_in_682, // @[:@39989.4]
  input  [4:0] io_in_683, // @[:@39989.4]
  input  [4:0] io_in_684, // @[:@39989.4]
  input  [4:0] io_in_685, // @[:@39989.4]
  input  [4:0] io_in_686, // @[:@39989.4]
  input  [4:0] io_in_687, // @[:@39989.4]
  input  [4:0] io_in_688, // @[:@39989.4]
  input  [4:0] io_in_689, // @[:@39989.4]
  input  [4:0] io_in_690, // @[:@39989.4]
  input  [4:0] io_in_691, // @[:@39989.4]
  input  [4:0] io_in_692, // @[:@39989.4]
  input  [4:0] io_in_693, // @[:@39989.4]
  input  [4:0] io_in_694, // @[:@39989.4]
  input  [4:0] io_in_695, // @[:@39989.4]
  input  [4:0] io_in_696, // @[:@39989.4]
  input  [4:0] io_in_697, // @[:@39989.4]
  input  [4:0] io_in_698, // @[:@39989.4]
  input  [4:0] io_in_699, // @[:@39989.4]
  input  [4:0] io_in_700, // @[:@39989.4]
  input  [4:0] io_in_701, // @[:@39989.4]
  input  [4:0] io_in_702, // @[:@39989.4]
  input  [4:0] io_in_703, // @[:@39989.4]
  input  [4:0] io_in_704, // @[:@39989.4]
  input  [4:0] io_in_705, // @[:@39989.4]
  input  [4:0] io_in_706, // @[:@39989.4]
  input  [4:0] io_in_707, // @[:@39989.4]
  input  [4:0] io_in_708, // @[:@39989.4]
  input  [4:0] io_in_709, // @[:@39989.4]
  input  [4:0] io_in_710, // @[:@39989.4]
  input  [4:0] io_in_711, // @[:@39989.4]
  input  [4:0] io_in_712, // @[:@39989.4]
  input  [4:0] io_in_713, // @[:@39989.4]
  input  [4:0] io_in_714, // @[:@39989.4]
  input  [4:0] io_in_715, // @[:@39989.4]
  input  [4:0] io_in_716, // @[:@39989.4]
  input  [4:0] io_in_717, // @[:@39989.4]
  input  [4:0] io_in_718, // @[:@39989.4]
  input  [4:0] io_in_719, // @[:@39989.4]
  input  [4:0] io_in_720, // @[:@39989.4]
  input  [4:0] io_in_721, // @[:@39989.4]
  input  [4:0] io_in_722, // @[:@39989.4]
  input  [4:0] io_in_723, // @[:@39989.4]
  input  [4:0] io_in_724, // @[:@39989.4]
  input  [4:0] io_in_725, // @[:@39989.4]
  input  [4:0] io_in_726, // @[:@39989.4]
  input  [4:0] io_in_727, // @[:@39989.4]
  input  [4:0] io_in_728, // @[:@39989.4]
  input  [4:0] io_in_729, // @[:@39989.4]
  input  [4:0] io_in_730, // @[:@39989.4]
  input  [4:0] io_in_731, // @[:@39989.4]
  input  [4:0] io_in_732, // @[:@39989.4]
  input  [4:0] io_in_733, // @[:@39989.4]
  input  [4:0] io_in_734, // @[:@39989.4]
  input  [4:0] io_in_735, // @[:@39989.4]
  input  [4:0] io_in_736, // @[:@39989.4]
  input  [4:0] io_in_737, // @[:@39989.4]
  input  [4:0] io_in_738, // @[:@39989.4]
  input  [4:0] io_in_739, // @[:@39989.4]
  input  [4:0] io_in_740, // @[:@39989.4]
  input  [4:0] io_in_741, // @[:@39989.4]
  input  [4:0] io_in_742, // @[:@39989.4]
  input  [4:0] io_in_743, // @[:@39989.4]
  input  [4:0] io_in_744, // @[:@39989.4]
  input  [4:0] io_in_745, // @[:@39989.4]
  input  [4:0] io_in_746, // @[:@39989.4]
  input  [4:0] io_in_747, // @[:@39989.4]
  input  [4:0] io_in_748, // @[:@39989.4]
  input  [4:0] io_in_749, // @[:@39989.4]
  input  [4:0] io_in_750, // @[:@39989.4]
  input  [4:0] io_in_751, // @[:@39989.4]
  input  [4:0] io_in_752, // @[:@39989.4]
  input  [4:0] io_in_753, // @[:@39989.4]
  input  [4:0] io_in_754, // @[:@39989.4]
  input  [4:0] io_in_755, // @[:@39989.4]
  input  [4:0] io_in_756, // @[:@39989.4]
  input  [4:0] io_in_757, // @[:@39989.4]
  input  [4:0] io_in_758, // @[:@39989.4]
  input  [4:0] io_in_759, // @[:@39989.4]
  input  [4:0] io_in_760, // @[:@39989.4]
  input  [4:0] io_in_761, // @[:@39989.4]
  input  [4:0] io_in_762, // @[:@39989.4]
  input  [4:0] io_in_763, // @[:@39989.4]
  input  [4:0] io_in_764, // @[:@39989.4]
  input  [4:0] io_in_765, // @[:@39989.4]
  input  [4:0] io_in_766, // @[:@39989.4]
  input  [4:0] io_in_767, // @[:@39989.4]
  input  [4:0] io_in_768, // @[:@39989.4]
  input  [4:0] io_in_769, // @[:@39989.4]
  input  [4:0] io_in_770, // @[:@39989.4]
  input  [4:0] io_in_771, // @[:@39989.4]
  input  [4:0] io_in_772, // @[:@39989.4]
  input  [4:0] io_in_773, // @[:@39989.4]
  input  [4:0] io_in_774, // @[:@39989.4]
  input  [4:0] io_in_775, // @[:@39989.4]
  input  [4:0] io_in_776, // @[:@39989.4]
  input  [4:0] io_in_777, // @[:@39989.4]
  input  [4:0] io_in_778, // @[:@39989.4]
  input  [4:0] io_in_779, // @[:@39989.4]
  input  [4:0] io_in_780, // @[:@39989.4]
  input  [4:0] io_in_781, // @[:@39989.4]
  input  [4:0] io_in_782, // @[:@39989.4]
  input  [4:0] io_in_783, // @[:@39989.4]
  output [7:0] io_out_0, // @[:@39989.4]
  output [7:0] io_out_1, // @[:@39989.4]
  output [7:0] io_out_2, // @[:@39989.4]
  output [7:0] io_out_3, // @[:@39989.4]
  output [7:0] io_out_4, // @[:@39989.4]
  output [7:0] io_out_5, // @[:@39989.4]
  output [7:0] io_out_6, // @[:@39989.4]
  output [7:0] io_out_7, // @[:@39989.4]
  output [7:0] io_out_8, // @[:@39989.4]
  output [7:0] io_out_9 // @[:@39989.4]
);
  wire [4:0] fc1_io_in_0; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_1; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_2; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_3; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_4; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_5; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_6; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_7; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_8; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_9; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_10; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_11; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_12; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_13; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_14; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_15; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_16; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_17; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_18; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_19; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_20; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_21; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_22; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_23; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_24; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_25; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_26; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_27; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_28; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_29; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_30; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_31; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_32; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_33; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_34; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_35; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_36; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_37; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_38; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_39; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_40; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_41; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_42; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_43; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_44; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_45; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_46; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_47; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_48; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_49; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_50; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_51; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_52; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_53; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_54; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_55; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_56; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_57; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_58; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_59; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_60; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_61; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_62; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_63; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_64; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_65; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_66; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_67; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_68; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_69; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_70; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_71; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_72; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_73; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_74; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_75; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_76; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_77; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_78; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_79; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_80; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_81; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_82; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_83; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_84; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_85; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_86; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_87; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_88; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_89; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_90; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_91; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_92; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_93; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_94; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_95; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_96; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_97; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_98; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_99; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_100; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_101; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_102; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_103; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_104; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_105; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_106; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_107; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_108; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_109; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_110; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_111; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_112; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_113; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_114; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_115; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_116; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_117; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_118; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_119; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_120; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_121; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_122; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_123; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_124; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_125; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_126; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_127; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_128; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_129; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_130; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_131; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_132; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_133; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_134; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_135; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_136; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_137; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_138; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_139; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_140; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_141; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_142; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_143; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_144; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_145; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_146; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_147; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_148; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_149; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_150; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_151; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_152; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_153; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_154; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_155; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_156; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_157; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_158; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_159; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_160; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_161; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_162; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_163; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_164; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_165; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_166; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_167; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_168; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_169; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_170; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_171; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_172; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_173; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_174; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_175; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_176; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_177; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_178; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_179; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_180; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_181; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_182; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_183; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_184; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_185; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_186; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_187; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_188; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_189; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_190; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_191; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_192; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_193; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_194; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_195; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_196; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_197; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_198; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_199; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_200; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_201; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_202; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_203; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_204; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_205; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_206; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_207; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_208; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_209; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_210; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_211; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_212; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_213; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_214; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_215; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_216; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_217; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_218; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_219; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_220; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_221; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_222; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_223; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_224; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_225; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_226; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_227; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_228; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_229; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_230; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_231; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_232; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_233; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_234; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_235; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_236; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_237; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_238; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_239; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_240; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_241; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_242; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_243; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_244; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_245; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_246; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_247; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_248; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_249; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_250; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_251; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_252; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_253; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_254; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_255; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_256; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_257; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_258; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_259; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_260; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_261; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_262; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_263; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_264; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_265; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_266; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_267; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_268; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_269; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_270; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_271; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_272; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_273; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_274; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_275; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_276; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_277; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_278; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_279; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_280; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_281; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_282; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_283; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_284; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_285; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_286; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_287; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_288; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_289; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_290; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_291; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_292; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_293; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_294; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_295; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_296; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_297; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_298; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_299; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_300; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_301; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_302; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_303; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_304; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_305; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_306; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_307; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_308; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_309; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_310; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_311; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_312; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_313; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_314; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_315; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_316; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_317; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_318; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_319; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_320; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_321; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_322; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_323; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_324; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_325; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_326; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_327; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_328; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_329; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_330; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_331; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_332; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_333; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_334; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_335; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_336; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_337; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_338; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_339; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_340; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_341; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_342; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_343; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_344; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_345; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_346; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_347; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_348; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_349; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_350; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_351; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_352; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_353; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_354; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_355; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_356; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_357; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_358; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_359; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_360; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_361; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_362; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_363; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_364; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_365; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_366; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_367; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_368; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_369; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_370; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_371; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_372; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_373; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_374; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_375; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_376; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_377; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_378; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_379; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_380; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_381; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_382; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_383; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_384; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_385; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_386; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_387; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_388; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_389; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_390; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_391; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_392; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_393; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_394; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_395; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_396; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_397; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_398; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_399; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_400; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_401; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_402; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_403; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_404; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_405; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_406; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_407; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_408; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_409; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_410; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_411; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_412; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_413; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_414; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_415; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_416; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_417; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_418; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_419; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_420; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_421; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_422; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_423; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_424; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_425; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_426; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_427; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_428; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_429; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_430; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_431; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_432; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_433; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_434; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_435; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_436; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_437; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_438; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_439; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_440; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_441; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_442; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_443; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_444; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_445; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_446; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_447; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_448; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_449; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_450; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_451; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_452; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_453; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_454; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_455; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_456; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_457; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_458; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_459; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_460; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_461; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_462; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_463; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_464; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_465; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_466; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_467; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_468; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_469; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_470; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_471; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_472; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_473; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_474; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_475; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_476; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_477; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_478; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_479; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_480; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_481; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_482; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_483; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_484; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_485; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_486; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_487; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_488; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_489; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_490; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_491; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_492; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_493; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_494; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_495; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_496; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_497; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_498; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_499; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_500; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_501; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_502; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_503; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_504; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_505; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_506; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_507; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_508; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_509; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_510; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_511; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_512; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_513; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_514; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_515; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_516; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_517; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_518; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_519; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_520; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_521; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_522; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_523; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_524; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_525; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_526; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_527; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_528; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_529; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_530; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_531; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_532; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_533; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_534; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_535; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_536; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_537; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_538; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_539; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_540; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_541; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_542; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_543; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_544; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_545; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_546; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_547; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_548; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_549; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_550; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_551; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_552; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_553; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_554; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_555; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_556; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_557; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_558; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_559; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_560; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_561; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_562; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_563; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_564; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_565; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_566; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_567; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_568; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_569; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_570; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_571; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_572; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_573; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_574; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_575; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_576; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_577; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_578; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_579; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_580; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_581; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_582; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_583; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_584; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_585; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_586; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_587; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_588; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_589; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_590; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_591; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_592; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_593; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_594; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_595; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_596; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_597; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_598; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_599; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_600; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_601; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_602; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_603; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_604; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_605; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_606; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_607; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_608; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_609; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_610; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_611; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_612; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_613; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_614; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_615; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_616; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_617; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_618; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_619; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_620; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_621; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_622; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_623; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_624; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_625; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_626; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_627; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_628; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_629; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_630; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_631; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_632; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_633; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_634; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_635; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_636; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_637; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_638; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_639; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_640; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_641; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_642; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_643; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_644; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_645; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_646; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_647; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_648; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_649; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_650; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_651; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_652; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_653; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_654; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_655; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_656; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_657; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_658; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_659; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_660; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_661; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_662; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_663; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_664; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_665; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_666; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_667; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_668; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_669; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_670; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_671; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_672; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_673; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_674; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_675; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_676; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_677; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_678; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_679; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_680; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_681; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_682; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_683; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_684; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_685; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_686; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_687; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_688; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_689; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_690; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_691; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_692; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_693; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_694; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_695; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_696; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_697; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_698; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_699; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_700; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_701; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_702; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_703; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_704; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_705; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_706; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_707; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_708; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_709; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_710; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_711; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_712; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_713; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_714; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_715; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_716; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_717; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_718; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_719; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_720; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_721; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_722; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_723; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_724; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_725; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_726; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_727; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_728; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_729; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_730; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_731; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_732; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_733; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_734; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_735; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_736; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_737; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_738; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_739; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_740; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_741; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_742; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_743; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_744; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_745; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_746; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_747; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_748; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_749; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_750; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_751; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_752; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_753; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_754; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_755; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_756; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_757; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_758; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_759; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_760; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_761; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_762; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_763; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_764; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_765; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_766; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_767; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_768; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_769; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_770; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_771; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_772; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_773; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_774; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_775; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_776; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_777; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_778; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_779; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_780; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_781; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_782; // @[Modules.scala 199:21:@39991.4]
  wire [4:0] fc1_io_in_783; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_0; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_1; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_2; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_3; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_4; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_5; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_6; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_7; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_8; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_9; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_10; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_11; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_12; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_13; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_14; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] fc1_io_out_15; // @[Modules.scala 199:21:@39991.4]
  wire [10:0] bn1_io_in_0; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_1; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_2; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_3; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_4; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_5; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_6; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_7; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_8; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_9; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_10; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_11; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_12; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_13; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_14; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_in_15; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_0; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_1; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_2; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_3; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_4; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_5; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_6; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_7; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_8; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_9; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_10; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_11; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_12; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_13; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_14; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bn1_io_out_15; // @[Modules.scala 200:21:@39994.4]
  wire [10:0] bi1_io_in_0; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_1; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_2; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_3; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_4; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_5; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_6; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_7; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_8; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_9; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_10; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_11; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_12; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_13; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_14; // @[Modules.scala 201:21:@39997.4]
  wire [10:0] bi1_io_in_15; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_0; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_1; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_2; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_3; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_4; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_5; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_6; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_7; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_8; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_9; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_10; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_11; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_12; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_13; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_14; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] bi1_io_out_15; // @[Modules.scala 201:21:@39997.4]
  wire [1:0] fc2_io_in_0; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_1; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_2; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_3; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_4; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_5; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_6; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_7; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_8; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_9; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_10; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_11; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_12; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_13; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_14; // @[Modules.scala 203:21:@40000.4]
  wire [1:0] fc2_io_in_15; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_0; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_1; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_2; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_3; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_4; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_5; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_6; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_7; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_8; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_9; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_10; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_11; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_12; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_13; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_14; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] fc2_io_out_15; // @[Modules.scala 203:21:@40000.4]
  wire [7:0] bn2_io_in_0; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_1; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_2; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_3; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_4; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_5; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_6; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_7; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_8; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_9; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_10; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_11; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_12; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_13; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_14; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_in_15; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_0; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_1; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_2; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_3; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_4; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_5; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_6; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_7; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_8; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_9; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_10; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_11; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_12; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_13; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_14; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bn2_io_out_15; // @[Modules.scala 204:21:@40003.4]
  wire [7:0] bi2_io_in_0; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_1; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_2; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_3; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_4; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_5; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_6; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_7; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_8; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_9; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_10; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_11; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_12; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_13; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_14; // @[Modules.scala 205:21:@40006.4]
  wire [7:0] bi2_io_in_15; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_0; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_1; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_2; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_3; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_4; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_5; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_6; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_7; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_8; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_9; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_10; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_11; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_12; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_13; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_14; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] bi2_io_out_15; // @[Modules.scala 205:21:@40006.4]
  wire [1:0] fc3_io_in_0; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_1; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_2; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_3; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_4; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_5; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_6; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_7; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_8; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_9; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_10; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_11; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_12; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_13; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_14; // @[Modules.scala 207:21:@40009.4]
  wire [1:0] fc3_io_in_15; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_0; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_1; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_2; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_3; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_4; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_5; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_6; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_7; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_8; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] fc3_io_out_9; // @[Modules.scala 207:21:@40009.4]
  wire [7:0] bn3_io_in_0; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_1; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_2; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_3; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_4; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_5; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_6; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_7; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_8; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_in_9; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_0; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_1; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_2; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_3; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_4; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_5; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_6; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_7; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_8; // @[Modules.scala 208:21:@40012.4]
  wire [7:0] bn3_io_out_9; // @[Modules.scala 208:21:@40012.4]
  Linear_p fc1 ( // @[Modules.scala 199:21:@39991.4]
    .io_in_0(fc1_io_in_0),
    .io_in_1(fc1_io_in_1),
    .io_in_2(fc1_io_in_2),
    .io_in_3(fc1_io_in_3),
    .io_in_4(fc1_io_in_4),
    .io_in_5(fc1_io_in_5),
    .io_in_6(fc1_io_in_6),
    .io_in_7(fc1_io_in_7),
    .io_in_8(fc1_io_in_8),
    .io_in_9(fc1_io_in_9),
    .io_in_10(fc1_io_in_10),
    .io_in_11(fc1_io_in_11),
    .io_in_12(fc1_io_in_12),
    .io_in_13(fc1_io_in_13),
    .io_in_14(fc1_io_in_14),
    .io_in_15(fc1_io_in_15),
    .io_in_16(fc1_io_in_16),
    .io_in_17(fc1_io_in_17),
    .io_in_18(fc1_io_in_18),
    .io_in_19(fc1_io_in_19),
    .io_in_20(fc1_io_in_20),
    .io_in_21(fc1_io_in_21),
    .io_in_22(fc1_io_in_22),
    .io_in_23(fc1_io_in_23),
    .io_in_24(fc1_io_in_24),
    .io_in_25(fc1_io_in_25),
    .io_in_26(fc1_io_in_26),
    .io_in_27(fc1_io_in_27),
    .io_in_28(fc1_io_in_28),
    .io_in_29(fc1_io_in_29),
    .io_in_30(fc1_io_in_30),
    .io_in_31(fc1_io_in_31),
    .io_in_32(fc1_io_in_32),
    .io_in_33(fc1_io_in_33),
    .io_in_34(fc1_io_in_34),
    .io_in_35(fc1_io_in_35),
    .io_in_36(fc1_io_in_36),
    .io_in_37(fc1_io_in_37),
    .io_in_38(fc1_io_in_38),
    .io_in_39(fc1_io_in_39),
    .io_in_40(fc1_io_in_40),
    .io_in_41(fc1_io_in_41),
    .io_in_42(fc1_io_in_42),
    .io_in_43(fc1_io_in_43),
    .io_in_44(fc1_io_in_44),
    .io_in_45(fc1_io_in_45),
    .io_in_46(fc1_io_in_46),
    .io_in_47(fc1_io_in_47),
    .io_in_48(fc1_io_in_48),
    .io_in_49(fc1_io_in_49),
    .io_in_50(fc1_io_in_50),
    .io_in_51(fc1_io_in_51),
    .io_in_52(fc1_io_in_52),
    .io_in_53(fc1_io_in_53),
    .io_in_54(fc1_io_in_54),
    .io_in_55(fc1_io_in_55),
    .io_in_56(fc1_io_in_56),
    .io_in_57(fc1_io_in_57),
    .io_in_58(fc1_io_in_58),
    .io_in_59(fc1_io_in_59),
    .io_in_60(fc1_io_in_60),
    .io_in_61(fc1_io_in_61),
    .io_in_62(fc1_io_in_62),
    .io_in_63(fc1_io_in_63),
    .io_in_64(fc1_io_in_64),
    .io_in_65(fc1_io_in_65),
    .io_in_66(fc1_io_in_66),
    .io_in_67(fc1_io_in_67),
    .io_in_68(fc1_io_in_68),
    .io_in_69(fc1_io_in_69),
    .io_in_70(fc1_io_in_70),
    .io_in_71(fc1_io_in_71),
    .io_in_72(fc1_io_in_72),
    .io_in_73(fc1_io_in_73),
    .io_in_74(fc1_io_in_74),
    .io_in_75(fc1_io_in_75),
    .io_in_76(fc1_io_in_76),
    .io_in_77(fc1_io_in_77),
    .io_in_78(fc1_io_in_78),
    .io_in_79(fc1_io_in_79),
    .io_in_80(fc1_io_in_80),
    .io_in_81(fc1_io_in_81),
    .io_in_82(fc1_io_in_82),
    .io_in_83(fc1_io_in_83),
    .io_in_84(fc1_io_in_84),
    .io_in_85(fc1_io_in_85),
    .io_in_86(fc1_io_in_86),
    .io_in_87(fc1_io_in_87),
    .io_in_88(fc1_io_in_88),
    .io_in_89(fc1_io_in_89),
    .io_in_90(fc1_io_in_90),
    .io_in_91(fc1_io_in_91),
    .io_in_92(fc1_io_in_92),
    .io_in_93(fc1_io_in_93),
    .io_in_94(fc1_io_in_94),
    .io_in_95(fc1_io_in_95),
    .io_in_96(fc1_io_in_96),
    .io_in_97(fc1_io_in_97),
    .io_in_98(fc1_io_in_98),
    .io_in_99(fc1_io_in_99),
    .io_in_100(fc1_io_in_100),
    .io_in_101(fc1_io_in_101),
    .io_in_102(fc1_io_in_102),
    .io_in_103(fc1_io_in_103),
    .io_in_104(fc1_io_in_104),
    .io_in_105(fc1_io_in_105),
    .io_in_106(fc1_io_in_106),
    .io_in_107(fc1_io_in_107),
    .io_in_108(fc1_io_in_108),
    .io_in_109(fc1_io_in_109),
    .io_in_110(fc1_io_in_110),
    .io_in_111(fc1_io_in_111),
    .io_in_112(fc1_io_in_112),
    .io_in_113(fc1_io_in_113),
    .io_in_114(fc1_io_in_114),
    .io_in_115(fc1_io_in_115),
    .io_in_116(fc1_io_in_116),
    .io_in_117(fc1_io_in_117),
    .io_in_118(fc1_io_in_118),
    .io_in_119(fc1_io_in_119),
    .io_in_120(fc1_io_in_120),
    .io_in_121(fc1_io_in_121),
    .io_in_122(fc1_io_in_122),
    .io_in_123(fc1_io_in_123),
    .io_in_124(fc1_io_in_124),
    .io_in_125(fc1_io_in_125),
    .io_in_126(fc1_io_in_126),
    .io_in_127(fc1_io_in_127),
    .io_in_128(fc1_io_in_128),
    .io_in_129(fc1_io_in_129),
    .io_in_130(fc1_io_in_130),
    .io_in_131(fc1_io_in_131),
    .io_in_132(fc1_io_in_132),
    .io_in_133(fc1_io_in_133),
    .io_in_134(fc1_io_in_134),
    .io_in_135(fc1_io_in_135),
    .io_in_136(fc1_io_in_136),
    .io_in_137(fc1_io_in_137),
    .io_in_138(fc1_io_in_138),
    .io_in_139(fc1_io_in_139),
    .io_in_140(fc1_io_in_140),
    .io_in_141(fc1_io_in_141),
    .io_in_142(fc1_io_in_142),
    .io_in_143(fc1_io_in_143),
    .io_in_144(fc1_io_in_144),
    .io_in_145(fc1_io_in_145),
    .io_in_146(fc1_io_in_146),
    .io_in_147(fc1_io_in_147),
    .io_in_148(fc1_io_in_148),
    .io_in_149(fc1_io_in_149),
    .io_in_150(fc1_io_in_150),
    .io_in_151(fc1_io_in_151),
    .io_in_152(fc1_io_in_152),
    .io_in_153(fc1_io_in_153),
    .io_in_154(fc1_io_in_154),
    .io_in_155(fc1_io_in_155),
    .io_in_156(fc1_io_in_156),
    .io_in_157(fc1_io_in_157),
    .io_in_158(fc1_io_in_158),
    .io_in_159(fc1_io_in_159),
    .io_in_160(fc1_io_in_160),
    .io_in_161(fc1_io_in_161),
    .io_in_162(fc1_io_in_162),
    .io_in_163(fc1_io_in_163),
    .io_in_164(fc1_io_in_164),
    .io_in_165(fc1_io_in_165),
    .io_in_166(fc1_io_in_166),
    .io_in_167(fc1_io_in_167),
    .io_in_168(fc1_io_in_168),
    .io_in_169(fc1_io_in_169),
    .io_in_170(fc1_io_in_170),
    .io_in_171(fc1_io_in_171),
    .io_in_172(fc1_io_in_172),
    .io_in_173(fc1_io_in_173),
    .io_in_174(fc1_io_in_174),
    .io_in_175(fc1_io_in_175),
    .io_in_176(fc1_io_in_176),
    .io_in_177(fc1_io_in_177),
    .io_in_178(fc1_io_in_178),
    .io_in_179(fc1_io_in_179),
    .io_in_180(fc1_io_in_180),
    .io_in_181(fc1_io_in_181),
    .io_in_182(fc1_io_in_182),
    .io_in_183(fc1_io_in_183),
    .io_in_184(fc1_io_in_184),
    .io_in_185(fc1_io_in_185),
    .io_in_186(fc1_io_in_186),
    .io_in_187(fc1_io_in_187),
    .io_in_188(fc1_io_in_188),
    .io_in_189(fc1_io_in_189),
    .io_in_190(fc1_io_in_190),
    .io_in_191(fc1_io_in_191),
    .io_in_192(fc1_io_in_192),
    .io_in_193(fc1_io_in_193),
    .io_in_194(fc1_io_in_194),
    .io_in_195(fc1_io_in_195),
    .io_in_196(fc1_io_in_196),
    .io_in_197(fc1_io_in_197),
    .io_in_198(fc1_io_in_198),
    .io_in_199(fc1_io_in_199),
    .io_in_200(fc1_io_in_200),
    .io_in_201(fc1_io_in_201),
    .io_in_202(fc1_io_in_202),
    .io_in_203(fc1_io_in_203),
    .io_in_204(fc1_io_in_204),
    .io_in_205(fc1_io_in_205),
    .io_in_206(fc1_io_in_206),
    .io_in_207(fc1_io_in_207),
    .io_in_208(fc1_io_in_208),
    .io_in_209(fc1_io_in_209),
    .io_in_210(fc1_io_in_210),
    .io_in_211(fc1_io_in_211),
    .io_in_212(fc1_io_in_212),
    .io_in_213(fc1_io_in_213),
    .io_in_214(fc1_io_in_214),
    .io_in_215(fc1_io_in_215),
    .io_in_216(fc1_io_in_216),
    .io_in_217(fc1_io_in_217),
    .io_in_218(fc1_io_in_218),
    .io_in_219(fc1_io_in_219),
    .io_in_220(fc1_io_in_220),
    .io_in_221(fc1_io_in_221),
    .io_in_222(fc1_io_in_222),
    .io_in_223(fc1_io_in_223),
    .io_in_224(fc1_io_in_224),
    .io_in_225(fc1_io_in_225),
    .io_in_226(fc1_io_in_226),
    .io_in_227(fc1_io_in_227),
    .io_in_228(fc1_io_in_228),
    .io_in_229(fc1_io_in_229),
    .io_in_230(fc1_io_in_230),
    .io_in_231(fc1_io_in_231),
    .io_in_232(fc1_io_in_232),
    .io_in_233(fc1_io_in_233),
    .io_in_234(fc1_io_in_234),
    .io_in_235(fc1_io_in_235),
    .io_in_236(fc1_io_in_236),
    .io_in_237(fc1_io_in_237),
    .io_in_238(fc1_io_in_238),
    .io_in_239(fc1_io_in_239),
    .io_in_240(fc1_io_in_240),
    .io_in_241(fc1_io_in_241),
    .io_in_242(fc1_io_in_242),
    .io_in_243(fc1_io_in_243),
    .io_in_244(fc1_io_in_244),
    .io_in_245(fc1_io_in_245),
    .io_in_246(fc1_io_in_246),
    .io_in_247(fc1_io_in_247),
    .io_in_248(fc1_io_in_248),
    .io_in_249(fc1_io_in_249),
    .io_in_250(fc1_io_in_250),
    .io_in_251(fc1_io_in_251),
    .io_in_252(fc1_io_in_252),
    .io_in_253(fc1_io_in_253),
    .io_in_254(fc1_io_in_254),
    .io_in_255(fc1_io_in_255),
    .io_in_256(fc1_io_in_256),
    .io_in_257(fc1_io_in_257),
    .io_in_258(fc1_io_in_258),
    .io_in_259(fc1_io_in_259),
    .io_in_260(fc1_io_in_260),
    .io_in_261(fc1_io_in_261),
    .io_in_262(fc1_io_in_262),
    .io_in_263(fc1_io_in_263),
    .io_in_264(fc1_io_in_264),
    .io_in_265(fc1_io_in_265),
    .io_in_266(fc1_io_in_266),
    .io_in_267(fc1_io_in_267),
    .io_in_268(fc1_io_in_268),
    .io_in_269(fc1_io_in_269),
    .io_in_270(fc1_io_in_270),
    .io_in_271(fc1_io_in_271),
    .io_in_272(fc1_io_in_272),
    .io_in_273(fc1_io_in_273),
    .io_in_274(fc1_io_in_274),
    .io_in_275(fc1_io_in_275),
    .io_in_276(fc1_io_in_276),
    .io_in_277(fc1_io_in_277),
    .io_in_278(fc1_io_in_278),
    .io_in_279(fc1_io_in_279),
    .io_in_280(fc1_io_in_280),
    .io_in_281(fc1_io_in_281),
    .io_in_282(fc1_io_in_282),
    .io_in_283(fc1_io_in_283),
    .io_in_284(fc1_io_in_284),
    .io_in_285(fc1_io_in_285),
    .io_in_286(fc1_io_in_286),
    .io_in_287(fc1_io_in_287),
    .io_in_288(fc1_io_in_288),
    .io_in_289(fc1_io_in_289),
    .io_in_290(fc1_io_in_290),
    .io_in_291(fc1_io_in_291),
    .io_in_292(fc1_io_in_292),
    .io_in_293(fc1_io_in_293),
    .io_in_294(fc1_io_in_294),
    .io_in_295(fc1_io_in_295),
    .io_in_296(fc1_io_in_296),
    .io_in_297(fc1_io_in_297),
    .io_in_298(fc1_io_in_298),
    .io_in_299(fc1_io_in_299),
    .io_in_300(fc1_io_in_300),
    .io_in_301(fc1_io_in_301),
    .io_in_302(fc1_io_in_302),
    .io_in_303(fc1_io_in_303),
    .io_in_304(fc1_io_in_304),
    .io_in_305(fc1_io_in_305),
    .io_in_306(fc1_io_in_306),
    .io_in_307(fc1_io_in_307),
    .io_in_308(fc1_io_in_308),
    .io_in_309(fc1_io_in_309),
    .io_in_310(fc1_io_in_310),
    .io_in_311(fc1_io_in_311),
    .io_in_312(fc1_io_in_312),
    .io_in_313(fc1_io_in_313),
    .io_in_314(fc1_io_in_314),
    .io_in_315(fc1_io_in_315),
    .io_in_316(fc1_io_in_316),
    .io_in_317(fc1_io_in_317),
    .io_in_318(fc1_io_in_318),
    .io_in_319(fc1_io_in_319),
    .io_in_320(fc1_io_in_320),
    .io_in_321(fc1_io_in_321),
    .io_in_322(fc1_io_in_322),
    .io_in_323(fc1_io_in_323),
    .io_in_324(fc1_io_in_324),
    .io_in_325(fc1_io_in_325),
    .io_in_326(fc1_io_in_326),
    .io_in_327(fc1_io_in_327),
    .io_in_328(fc1_io_in_328),
    .io_in_329(fc1_io_in_329),
    .io_in_330(fc1_io_in_330),
    .io_in_331(fc1_io_in_331),
    .io_in_332(fc1_io_in_332),
    .io_in_333(fc1_io_in_333),
    .io_in_334(fc1_io_in_334),
    .io_in_335(fc1_io_in_335),
    .io_in_336(fc1_io_in_336),
    .io_in_337(fc1_io_in_337),
    .io_in_338(fc1_io_in_338),
    .io_in_339(fc1_io_in_339),
    .io_in_340(fc1_io_in_340),
    .io_in_341(fc1_io_in_341),
    .io_in_342(fc1_io_in_342),
    .io_in_343(fc1_io_in_343),
    .io_in_344(fc1_io_in_344),
    .io_in_345(fc1_io_in_345),
    .io_in_346(fc1_io_in_346),
    .io_in_347(fc1_io_in_347),
    .io_in_348(fc1_io_in_348),
    .io_in_349(fc1_io_in_349),
    .io_in_350(fc1_io_in_350),
    .io_in_351(fc1_io_in_351),
    .io_in_352(fc1_io_in_352),
    .io_in_353(fc1_io_in_353),
    .io_in_354(fc1_io_in_354),
    .io_in_355(fc1_io_in_355),
    .io_in_356(fc1_io_in_356),
    .io_in_357(fc1_io_in_357),
    .io_in_358(fc1_io_in_358),
    .io_in_359(fc1_io_in_359),
    .io_in_360(fc1_io_in_360),
    .io_in_361(fc1_io_in_361),
    .io_in_362(fc1_io_in_362),
    .io_in_363(fc1_io_in_363),
    .io_in_364(fc1_io_in_364),
    .io_in_365(fc1_io_in_365),
    .io_in_366(fc1_io_in_366),
    .io_in_367(fc1_io_in_367),
    .io_in_368(fc1_io_in_368),
    .io_in_369(fc1_io_in_369),
    .io_in_370(fc1_io_in_370),
    .io_in_371(fc1_io_in_371),
    .io_in_372(fc1_io_in_372),
    .io_in_373(fc1_io_in_373),
    .io_in_374(fc1_io_in_374),
    .io_in_375(fc1_io_in_375),
    .io_in_376(fc1_io_in_376),
    .io_in_377(fc1_io_in_377),
    .io_in_378(fc1_io_in_378),
    .io_in_379(fc1_io_in_379),
    .io_in_380(fc1_io_in_380),
    .io_in_381(fc1_io_in_381),
    .io_in_382(fc1_io_in_382),
    .io_in_383(fc1_io_in_383),
    .io_in_384(fc1_io_in_384),
    .io_in_385(fc1_io_in_385),
    .io_in_386(fc1_io_in_386),
    .io_in_387(fc1_io_in_387),
    .io_in_388(fc1_io_in_388),
    .io_in_389(fc1_io_in_389),
    .io_in_390(fc1_io_in_390),
    .io_in_391(fc1_io_in_391),
    .io_in_392(fc1_io_in_392),
    .io_in_393(fc1_io_in_393),
    .io_in_394(fc1_io_in_394),
    .io_in_395(fc1_io_in_395),
    .io_in_396(fc1_io_in_396),
    .io_in_397(fc1_io_in_397),
    .io_in_398(fc1_io_in_398),
    .io_in_399(fc1_io_in_399),
    .io_in_400(fc1_io_in_400),
    .io_in_401(fc1_io_in_401),
    .io_in_402(fc1_io_in_402),
    .io_in_403(fc1_io_in_403),
    .io_in_404(fc1_io_in_404),
    .io_in_405(fc1_io_in_405),
    .io_in_406(fc1_io_in_406),
    .io_in_407(fc1_io_in_407),
    .io_in_408(fc1_io_in_408),
    .io_in_409(fc1_io_in_409),
    .io_in_410(fc1_io_in_410),
    .io_in_411(fc1_io_in_411),
    .io_in_412(fc1_io_in_412),
    .io_in_413(fc1_io_in_413),
    .io_in_414(fc1_io_in_414),
    .io_in_415(fc1_io_in_415),
    .io_in_416(fc1_io_in_416),
    .io_in_417(fc1_io_in_417),
    .io_in_418(fc1_io_in_418),
    .io_in_419(fc1_io_in_419),
    .io_in_420(fc1_io_in_420),
    .io_in_421(fc1_io_in_421),
    .io_in_422(fc1_io_in_422),
    .io_in_423(fc1_io_in_423),
    .io_in_424(fc1_io_in_424),
    .io_in_425(fc1_io_in_425),
    .io_in_426(fc1_io_in_426),
    .io_in_427(fc1_io_in_427),
    .io_in_428(fc1_io_in_428),
    .io_in_429(fc1_io_in_429),
    .io_in_430(fc1_io_in_430),
    .io_in_431(fc1_io_in_431),
    .io_in_432(fc1_io_in_432),
    .io_in_433(fc1_io_in_433),
    .io_in_434(fc1_io_in_434),
    .io_in_435(fc1_io_in_435),
    .io_in_436(fc1_io_in_436),
    .io_in_437(fc1_io_in_437),
    .io_in_438(fc1_io_in_438),
    .io_in_439(fc1_io_in_439),
    .io_in_440(fc1_io_in_440),
    .io_in_441(fc1_io_in_441),
    .io_in_442(fc1_io_in_442),
    .io_in_443(fc1_io_in_443),
    .io_in_444(fc1_io_in_444),
    .io_in_445(fc1_io_in_445),
    .io_in_446(fc1_io_in_446),
    .io_in_447(fc1_io_in_447),
    .io_in_448(fc1_io_in_448),
    .io_in_449(fc1_io_in_449),
    .io_in_450(fc1_io_in_450),
    .io_in_451(fc1_io_in_451),
    .io_in_452(fc1_io_in_452),
    .io_in_453(fc1_io_in_453),
    .io_in_454(fc1_io_in_454),
    .io_in_455(fc1_io_in_455),
    .io_in_456(fc1_io_in_456),
    .io_in_457(fc1_io_in_457),
    .io_in_458(fc1_io_in_458),
    .io_in_459(fc1_io_in_459),
    .io_in_460(fc1_io_in_460),
    .io_in_461(fc1_io_in_461),
    .io_in_462(fc1_io_in_462),
    .io_in_463(fc1_io_in_463),
    .io_in_464(fc1_io_in_464),
    .io_in_465(fc1_io_in_465),
    .io_in_466(fc1_io_in_466),
    .io_in_467(fc1_io_in_467),
    .io_in_468(fc1_io_in_468),
    .io_in_469(fc1_io_in_469),
    .io_in_470(fc1_io_in_470),
    .io_in_471(fc1_io_in_471),
    .io_in_472(fc1_io_in_472),
    .io_in_473(fc1_io_in_473),
    .io_in_474(fc1_io_in_474),
    .io_in_475(fc1_io_in_475),
    .io_in_476(fc1_io_in_476),
    .io_in_477(fc1_io_in_477),
    .io_in_478(fc1_io_in_478),
    .io_in_479(fc1_io_in_479),
    .io_in_480(fc1_io_in_480),
    .io_in_481(fc1_io_in_481),
    .io_in_482(fc1_io_in_482),
    .io_in_483(fc1_io_in_483),
    .io_in_484(fc1_io_in_484),
    .io_in_485(fc1_io_in_485),
    .io_in_486(fc1_io_in_486),
    .io_in_487(fc1_io_in_487),
    .io_in_488(fc1_io_in_488),
    .io_in_489(fc1_io_in_489),
    .io_in_490(fc1_io_in_490),
    .io_in_491(fc1_io_in_491),
    .io_in_492(fc1_io_in_492),
    .io_in_493(fc1_io_in_493),
    .io_in_494(fc1_io_in_494),
    .io_in_495(fc1_io_in_495),
    .io_in_496(fc1_io_in_496),
    .io_in_497(fc1_io_in_497),
    .io_in_498(fc1_io_in_498),
    .io_in_499(fc1_io_in_499),
    .io_in_500(fc1_io_in_500),
    .io_in_501(fc1_io_in_501),
    .io_in_502(fc1_io_in_502),
    .io_in_503(fc1_io_in_503),
    .io_in_504(fc1_io_in_504),
    .io_in_505(fc1_io_in_505),
    .io_in_506(fc1_io_in_506),
    .io_in_507(fc1_io_in_507),
    .io_in_508(fc1_io_in_508),
    .io_in_509(fc1_io_in_509),
    .io_in_510(fc1_io_in_510),
    .io_in_511(fc1_io_in_511),
    .io_in_512(fc1_io_in_512),
    .io_in_513(fc1_io_in_513),
    .io_in_514(fc1_io_in_514),
    .io_in_515(fc1_io_in_515),
    .io_in_516(fc1_io_in_516),
    .io_in_517(fc1_io_in_517),
    .io_in_518(fc1_io_in_518),
    .io_in_519(fc1_io_in_519),
    .io_in_520(fc1_io_in_520),
    .io_in_521(fc1_io_in_521),
    .io_in_522(fc1_io_in_522),
    .io_in_523(fc1_io_in_523),
    .io_in_524(fc1_io_in_524),
    .io_in_525(fc1_io_in_525),
    .io_in_526(fc1_io_in_526),
    .io_in_527(fc1_io_in_527),
    .io_in_528(fc1_io_in_528),
    .io_in_529(fc1_io_in_529),
    .io_in_530(fc1_io_in_530),
    .io_in_531(fc1_io_in_531),
    .io_in_532(fc1_io_in_532),
    .io_in_533(fc1_io_in_533),
    .io_in_534(fc1_io_in_534),
    .io_in_535(fc1_io_in_535),
    .io_in_536(fc1_io_in_536),
    .io_in_537(fc1_io_in_537),
    .io_in_538(fc1_io_in_538),
    .io_in_539(fc1_io_in_539),
    .io_in_540(fc1_io_in_540),
    .io_in_541(fc1_io_in_541),
    .io_in_542(fc1_io_in_542),
    .io_in_543(fc1_io_in_543),
    .io_in_544(fc1_io_in_544),
    .io_in_545(fc1_io_in_545),
    .io_in_546(fc1_io_in_546),
    .io_in_547(fc1_io_in_547),
    .io_in_548(fc1_io_in_548),
    .io_in_549(fc1_io_in_549),
    .io_in_550(fc1_io_in_550),
    .io_in_551(fc1_io_in_551),
    .io_in_552(fc1_io_in_552),
    .io_in_553(fc1_io_in_553),
    .io_in_554(fc1_io_in_554),
    .io_in_555(fc1_io_in_555),
    .io_in_556(fc1_io_in_556),
    .io_in_557(fc1_io_in_557),
    .io_in_558(fc1_io_in_558),
    .io_in_559(fc1_io_in_559),
    .io_in_560(fc1_io_in_560),
    .io_in_561(fc1_io_in_561),
    .io_in_562(fc1_io_in_562),
    .io_in_563(fc1_io_in_563),
    .io_in_564(fc1_io_in_564),
    .io_in_565(fc1_io_in_565),
    .io_in_566(fc1_io_in_566),
    .io_in_567(fc1_io_in_567),
    .io_in_568(fc1_io_in_568),
    .io_in_569(fc1_io_in_569),
    .io_in_570(fc1_io_in_570),
    .io_in_571(fc1_io_in_571),
    .io_in_572(fc1_io_in_572),
    .io_in_573(fc1_io_in_573),
    .io_in_574(fc1_io_in_574),
    .io_in_575(fc1_io_in_575),
    .io_in_576(fc1_io_in_576),
    .io_in_577(fc1_io_in_577),
    .io_in_578(fc1_io_in_578),
    .io_in_579(fc1_io_in_579),
    .io_in_580(fc1_io_in_580),
    .io_in_581(fc1_io_in_581),
    .io_in_582(fc1_io_in_582),
    .io_in_583(fc1_io_in_583),
    .io_in_584(fc1_io_in_584),
    .io_in_585(fc1_io_in_585),
    .io_in_586(fc1_io_in_586),
    .io_in_587(fc1_io_in_587),
    .io_in_588(fc1_io_in_588),
    .io_in_589(fc1_io_in_589),
    .io_in_590(fc1_io_in_590),
    .io_in_591(fc1_io_in_591),
    .io_in_592(fc1_io_in_592),
    .io_in_593(fc1_io_in_593),
    .io_in_594(fc1_io_in_594),
    .io_in_595(fc1_io_in_595),
    .io_in_596(fc1_io_in_596),
    .io_in_597(fc1_io_in_597),
    .io_in_598(fc1_io_in_598),
    .io_in_599(fc1_io_in_599),
    .io_in_600(fc1_io_in_600),
    .io_in_601(fc1_io_in_601),
    .io_in_602(fc1_io_in_602),
    .io_in_603(fc1_io_in_603),
    .io_in_604(fc1_io_in_604),
    .io_in_605(fc1_io_in_605),
    .io_in_606(fc1_io_in_606),
    .io_in_607(fc1_io_in_607),
    .io_in_608(fc1_io_in_608),
    .io_in_609(fc1_io_in_609),
    .io_in_610(fc1_io_in_610),
    .io_in_611(fc1_io_in_611),
    .io_in_612(fc1_io_in_612),
    .io_in_613(fc1_io_in_613),
    .io_in_614(fc1_io_in_614),
    .io_in_615(fc1_io_in_615),
    .io_in_616(fc1_io_in_616),
    .io_in_617(fc1_io_in_617),
    .io_in_618(fc1_io_in_618),
    .io_in_619(fc1_io_in_619),
    .io_in_620(fc1_io_in_620),
    .io_in_621(fc1_io_in_621),
    .io_in_622(fc1_io_in_622),
    .io_in_623(fc1_io_in_623),
    .io_in_624(fc1_io_in_624),
    .io_in_625(fc1_io_in_625),
    .io_in_626(fc1_io_in_626),
    .io_in_627(fc1_io_in_627),
    .io_in_628(fc1_io_in_628),
    .io_in_629(fc1_io_in_629),
    .io_in_630(fc1_io_in_630),
    .io_in_631(fc1_io_in_631),
    .io_in_632(fc1_io_in_632),
    .io_in_633(fc1_io_in_633),
    .io_in_634(fc1_io_in_634),
    .io_in_635(fc1_io_in_635),
    .io_in_636(fc1_io_in_636),
    .io_in_637(fc1_io_in_637),
    .io_in_638(fc1_io_in_638),
    .io_in_639(fc1_io_in_639),
    .io_in_640(fc1_io_in_640),
    .io_in_641(fc1_io_in_641),
    .io_in_642(fc1_io_in_642),
    .io_in_643(fc1_io_in_643),
    .io_in_644(fc1_io_in_644),
    .io_in_645(fc1_io_in_645),
    .io_in_646(fc1_io_in_646),
    .io_in_647(fc1_io_in_647),
    .io_in_648(fc1_io_in_648),
    .io_in_649(fc1_io_in_649),
    .io_in_650(fc1_io_in_650),
    .io_in_651(fc1_io_in_651),
    .io_in_652(fc1_io_in_652),
    .io_in_653(fc1_io_in_653),
    .io_in_654(fc1_io_in_654),
    .io_in_655(fc1_io_in_655),
    .io_in_656(fc1_io_in_656),
    .io_in_657(fc1_io_in_657),
    .io_in_658(fc1_io_in_658),
    .io_in_659(fc1_io_in_659),
    .io_in_660(fc1_io_in_660),
    .io_in_661(fc1_io_in_661),
    .io_in_662(fc1_io_in_662),
    .io_in_663(fc1_io_in_663),
    .io_in_664(fc1_io_in_664),
    .io_in_665(fc1_io_in_665),
    .io_in_666(fc1_io_in_666),
    .io_in_667(fc1_io_in_667),
    .io_in_668(fc1_io_in_668),
    .io_in_669(fc1_io_in_669),
    .io_in_670(fc1_io_in_670),
    .io_in_671(fc1_io_in_671),
    .io_in_672(fc1_io_in_672),
    .io_in_673(fc1_io_in_673),
    .io_in_674(fc1_io_in_674),
    .io_in_675(fc1_io_in_675),
    .io_in_676(fc1_io_in_676),
    .io_in_677(fc1_io_in_677),
    .io_in_678(fc1_io_in_678),
    .io_in_679(fc1_io_in_679),
    .io_in_680(fc1_io_in_680),
    .io_in_681(fc1_io_in_681),
    .io_in_682(fc1_io_in_682),
    .io_in_683(fc1_io_in_683),
    .io_in_684(fc1_io_in_684),
    .io_in_685(fc1_io_in_685),
    .io_in_686(fc1_io_in_686),
    .io_in_687(fc1_io_in_687),
    .io_in_688(fc1_io_in_688),
    .io_in_689(fc1_io_in_689),
    .io_in_690(fc1_io_in_690),
    .io_in_691(fc1_io_in_691),
    .io_in_692(fc1_io_in_692),
    .io_in_693(fc1_io_in_693),
    .io_in_694(fc1_io_in_694),
    .io_in_695(fc1_io_in_695),
    .io_in_696(fc1_io_in_696),
    .io_in_697(fc1_io_in_697),
    .io_in_698(fc1_io_in_698),
    .io_in_699(fc1_io_in_699),
    .io_in_700(fc1_io_in_700),
    .io_in_701(fc1_io_in_701),
    .io_in_702(fc1_io_in_702),
    .io_in_703(fc1_io_in_703),
    .io_in_704(fc1_io_in_704),
    .io_in_705(fc1_io_in_705),
    .io_in_706(fc1_io_in_706),
    .io_in_707(fc1_io_in_707),
    .io_in_708(fc1_io_in_708),
    .io_in_709(fc1_io_in_709),
    .io_in_710(fc1_io_in_710),
    .io_in_711(fc1_io_in_711),
    .io_in_712(fc1_io_in_712),
    .io_in_713(fc1_io_in_713),
    .io_in_714(fc1_io_in_714),
    .io_in_715(fc1_io_in_715),
    .io_in_716(fc1_io_in_716),
    .io_in_717(fc1_io_in_717),
    .io_in_718(fc1_io_in_718),
    .io_in_719(fc1_io_in_719),
    .io_in_720(fc1_io_in_720),
    .io_in_721(fc1_io_in_721),
    .io_in_722(fc1_io_in_722),
    .io_in_723(fc1_io_in_723),
    .io_in_724(fc1_io_in_724),
    .io_in_725(fc1_io_in_725),
    .io_in_726(fc1_io_in_726),
    .io_in_727(fc1_io_in_727),
    .io_in_728(fc1_io_in_728),
    .io_in_729(fc1_io_in_729),
    .io_in_730(fc1_io_in_730),
    .io_in_731(fc1_io_in_731),
    .io_in_732(fc1_io_in_732),
    .io_in_733(fc1_io_in_733),
    .io_in_734(fc1_io_in_734),
    .io_in_735(fc1_io_in_735),
    .io_in_736(fc1_io_in_736),
    .io_in_737(fc1_io_in_737),
    .io_in_738(fc1_io_in_738),
    .io_in_739(fc1_io_in_739),
    .io_in_740(fc1_io_in_740),
    .io_in_741(fc1_io_in_741),
    .io_in_742(fc1_io_in_742),
    .io_in_743(fc1_io_in_743),
    .io_in_744(fc1_io_in_744),
    .io_in_745(fc1_io_in_745),
    .io_in_746(fc1_io_in_746),
    .io_in_747(fc1_io_in_747),
    .io_in_748(fc1_io_in_748),
    .io_in_749(fc1_io_in_749),
    .io_in_750(fc1_io_in_750),
    .io_in_751(fc1_io_in_751),
    .io_in_752(fc1_io_in_752),
    .io_in_753(fc1_io_in_753),
    .io_in_754(fc1_io_in_754),
    .io_in_755(fc1_io_in_755),
    .io_in_756(fc1_io_in_756),
    .io_in_757(fc1_io_in_757),
    .io_in_758(fc1_io_in_758),
    .io_in_759(fc1_io_in_759),
    .io_in_760(fc1_io_in_760),
    .io_in_761(fc1_io_in_761),
    .io_in_762(fc1_io_in_762),
    .io_in_763(fc1_io_in_763),
    .io_in_764(fc1_io_in_764),
    .io_in_765(fc1_io_in_765),
    .io_in_766(fc1_io_in_766),
    .io_in_767(fc1_io_in_767),
    .io_in_768(fc1_io_in_768),
    .io_in_769(fc1_io_in_769),
    .io_in_770(fc1_io_in_770),
    .io_in_771(fc1_io_in_771),
    .io_in_772(fc1_io_in_772),
    .io_in_773(fc1_io_in_773),
    .io_in_774(fc1_io_in_774),
    .io_in_775(fc1_io_in_775),
    .io_in_776(fc1_io_in_776),
    .io_in_777(fc1_io_in_777),
    .io_in_778(fc1_io_in_778),
    .io_in_779(fc1_io_in_779),
    .io_in_780(fc1_io_in_780),
    .io_in_781(fc1_io_in_781),
    .io_in_782(fc1_io_in_782),
    .io_in_783(fc1_io_in_783),
    .io_out_0(fc1_io_out_0),
    .io_out_1(fc1_io_out_1),
    .io_out_2(fc1_io_out_2),
    .io_out_3(fc1_io_out_3),
    .io_out_4(fc1_io_out_4),
    .io_out_5(fc1_io_out_5),
    .io_out_6(fc1_io_out_6),
    .io_out_7(fc1_io_out_7),
    .io_out_8(fc1_io_out_8),
    .io_out_9(fc1_io_out_9),
    .io_out_10(fc1_io_out_10),
    .io_out_11(fc1_io_out_11),
    .io_out_12(fc1_io_out_12),
    .io_out_13(fc1_io_out_13),
    .io_out_14(fc1_io_out_14),
    .io_out_15(fc1_io_out_15)
  );
  ShifBatchNorm bn1 ( // @[Modules.scala 200:21:@39994.4]
    .io_in_0(bn1_io_in_0),
    .io_in_1(bn1_io_in_1),
    .io_in_2(bn1_io_in_2),
    .io_in_3(bn1_io_in_3),
    .io_in_4(bn1_io_in_4),
    .io_in_5(bn1_io_in_5),
    .io_in_6(bn1_io_in_6),
    .io_in_7(bn1_io_in_7),
    .io_in_8(bn1_io_in_8),
    .io_in_9(bn1_io_in_9),
    .io_in_10(bn1_io_in_10),
    .io_in_11(bn1_io_in_11),
    .io_in_12(bn1_io_in_12),
    .io_in_13(bn1_io_in_13),
    .io_in_14(bn1_io_in_14),
    .io_in_15(bn1_io_in_15),
    .io_out_0(bn1_io_out_0),
    .io_out_1(bn1_io_out_1),
    .io_out_2(bn1_io_out_2),
    .io_out_3(bn1_io_out_3),
    .io_out_4(bn1_io_out_4),
    .io_out_5(bn1_io_out_5),
    .io_out_6(bn1_io_out_6),
    .io_out_7(bn1_io_out_7),
    .io_out_8(bn1_io_out_8),
    .io_out_9(bn1_io_out_9),
    .io_out_10(bn1_io_out_10),
    .io_out_11(bn1_io_out_11),
    .io_out_12(bn1_io_out_12),
    .io_out_13(bn1_io_out_13),
    .io_out_14(bn1_io_out_14),
    .io_out_15(bn1_io_out_15)
  );
  Binarize bi1 ( // @[Modules.scala 201:21:@39997.4]
    .io_in_0(bi1_io_in_0),
    .io_in_1(bi1_io_in_1),
    .io_in_2(bi1_io_in_2),
    .io_in_3(bi1_io_in_3),
    .io_in_4(bi1_io_in_4),
    .io_in_5(bi1_io_in_5),
    .io_in_6(bi1_io_in_6),
    .io_in_7(bi1_io_in_7),
    .io_in_8(bi1_io_in_8),
    .io_in_9(bi1_io_in_9),
    .io_in_10(bi1_io_in_10),
    .io_in_11(bi1_io_in_11),
    .io_in_12(bi1_io_in_12),
    .io_in_13(bi1_io_in_13),
    .io_in_14(bi1_io_in_14),
    .io_in_15(bi1_io_in_15),
    .io_out_0(bi1_io_out_0),
    .io_out_1(bi1_io_out_1),
    .io_out_2(bi1_io_out_2),
    .io_out_3(bi1_io_out_3),
    .io_out_4(bi1_io_out_4),
    .io_out_5(bi1_io_out_5),
    .io_out_6(bi1_io_out_6),
    .io_out_7(bi1_io_out_7),
    .io_out_8(bi1_io_out_8),
    .io_out_9(bi1_io_out_9),
    .io_out_10(bi1_io_out_10),
    .io_out_11(bi1_io_out_11),
    .io_out_12(bi1_io_out_12),
    .io_out_13(bi1_io_out_13),
    .io_out_14(bi1_io_out_14),
    .io_out_15(bi1_io_out_15)
  );
  Linear fc2 ( // @[Modules.scala 203:21:@40000.4]
    .io_in_0(fc2_io_in_0),
    .io_in_1(fc2_io_in_1),
    .io_in_2(fc2_io_in_2),
    .io_in_3(fc2_io_in_3),
    .io_in_4(fc2_io_in_4),
    .io_in_5(fc2_io_in_5),
    .io_in_6(fc2_io_in_6),
    .io_in_7(fc2_io_in_7),
    .io_in_8(fc2_io_in_8),
    .io_in_9(fc2_io_in_9),
    .io_in_10(fc2_io_in_10),
    .io_in_11(fc2_io_in_11),
    .io_in_12(fc2_io_in_12),
    .io_in_13(fc2_io_in_13),
    .io_in_14(fc2_io_in_14),
    .io_in_15(fc2_io_in_15),
    .io_out_0(fc2_io_out_0),
    .io_out_1(fc2_io_out_1),
    .io_out_2(fc2_io_out_2),
    .io_out_3(fc2_io_out_3),
    .io_out_4(fc2_io_out_4),
    .io_out_5(fc2_io_out_5),
    .io_out_6(fc2_io_out_6),
    .io_out_7(fc2_io_out_7),
    .io_out_8(fc2_io_out_8),
    .io_out_9(fc2_io_out_9),
    .io_out_10(fc2_io_out_10),
    .io_out_11(fc2_io_out_11),
    .io_out_12(fc2_io_out_12),
    .io_out_13(fc2_io_out_13),
    .io_out_14(fc2_io_out_14),
    .io_out_15(fc2_io_out_15)
  );
  ShifBatchNorm_1 bn2 ( // @[Modules.scala 204:21:@40003.4]
    .io_in_0(bn2_io_in_0),
    .io_in_1(bn2_io_in_1),
    .io_in_2(bn2_io_in_2),
    .io_in_3(bn2_io_in_3),
    .io_in_4(bn2_io_in_4),
    .io_in_5(bn2_io_in_5),
    .io_in_6(bn2_io_in_6),
    .io_in_7(bn2_io_in_7),
    .io_in_8(bn2_io_in_8),
    .io_in_9(bn2_io_in_9),
    .io_in_10(bn2_io_in_10),
    .io_in_11(bn2_io_in_11),
    .io_in_12(bn2_io_in_12),
    .io_in_13(bn2_io_in_13),
    .io_in_14(bn2_io_in_14),
    .io_in_15(bn2_io_in_15),
    .io_out_0(bn2_io_out_0),
    .io_out_1(bn2_io_out_1),
    .io_out_2(bn2_io_out_2),
    .io_out_3(bn2_io_out_3),
    .io_out_4(bn2_io_out_4),
    .io_out_5(bn2_io_out_5),
    .io_out_6(bn2_io_out_6),
    .io_out_7(bn2_io_out_7),
    .io_out_8(bn2_io_out_8),
    .io_out_9(bn2_io_out_9),
    .io_out_10(bn2_io_out_10),
    .io_out_11(bn2_io_out_11),
    .io_out_12(bn2_io_out_12),
    .io_out_13(bn2_io_out_13),
    .io_out_14(bn2_io_out_14),
    .io_out_15(bn2_io_out_15)
  );
  Binarize_1 bi2 ( // @[Modules.scala 205:21:@40006.4]
    .io_in_0(bi2_io_in_0),
    .io_in_1(bi2_io_in_1),
    .io_in_2(bi2_io_in_2),
    .io_in_3(bi2_io_in_3),
    .io_in_4(bi2_io_in_4),
    .io_in_5(bi2_io_in_5),
    .io_in_6(bi2_io_in_6),
    .io_in_7(bi2_io_in_7),
    .io_in_8(bi2_io_in_8),
    .io_in_9(bi2_io_in_9),
    .io_in_10(bi2_io_in_10),
    .io_in_11(bi2_io_in_11),
    .io_in_12(bi2_io_in_12),
    .io_in_13(bi2_io_in_13),
    .io_in_14(bi2_io_in_14),
    .io_in_15(bi2_io_in_15),
    .io_out_0(bi2_io_out_0),
    .io_out_1(bi2_io_out_1),
    .io_out_2(bi2_io_out_2),
    .io_out_3(bi2_io_out_3),
    .io_out_4(bi2_io_out_4),
    .io_out_5(bi2_io_out_5),
    .io_out_6(bi2_io_out_6),
    .io_out_7(bi2_io_out_7),
    .io_out_8(bi2_io_out_8),
    .io_out_9(bi2_io_out_9),
    .io_out_10(bi2_io_out_10),
    .io_out_11(bi2_io_out_11),
    .io_out_12(bi2_io_out_12),
    .io_out_13(bi2_io_out_13),
    .io_out_14(bi2_io_out_14),
    .io_out_15(bi2_io_out_15)
  );
  Linear_1 fc3 ( // @[Modules.scala 207:21:@40009.4]
    .io_in_0(fc3_io_in_0),
    .io_in_1(fc3_io_in_1),
    .io_in_2(fc3_io_in_2),
    .io_in_3(fc3_io_in_3),
    .io_in_4(fc3_io_in_4),
    .io_in_5(fc3_io_in_5),
    .io_in_6(fc3_io_in_6),
    .io_in_7(fc3_io_in_7),
    .io_in_8(fc3_io_in_8),
    .io_in_9(fc3_io_in_9),
    .io_in_10(fc3_io_in_10),
    .io_in_11(fc3_io_in_11),
    .io_in_12(fc3_io_in_12),
    .io_in_13(fc3_io_in_13),
    .io_in_14(fc3_io_in_14),
    .io_in_15(fc3_io_in_15),
    .io_out_0(fc3_io_out_0),
    .io_out_1(fc3_io_out_1),
    .io_out_2(fc3_io_out_2),
    .io_out_3(fc3_io_out_3),
    .io_out_4(fc3_io_out_4),
    .io_out_5(fc3_io_out_5),
    .io_out_6(fc3_io_out_6),
    .io_out_7(fc3_io_out_7),
    .io_out_8(fc3_io_out_8),
    .io_out_9(fc3_io_out_9)
  );
  ShifBatchNorm_2 bn3 ( // @[Modules.scala 208:21:@40012.4]
    .io_in_0(bn3_io_in_0),
    .io_in_1(bn3_io_in_1),
    .io_in_2(bn3_io_in_2),
    .io_in_3(bn3_io_in_3),
    .io_in_4(bn3_io_in_4),
    .io_in_5(bn3_io_in_5),
    .io_in_6(bn3_io_in_6),
    .io_in_7(bn3_io_in_7),
    .io_in_8(bn3_io_in_8),
    .io_in_9(bn3_io_in_9),
    .io_out_0(bn3_io_out_0),
    .io_out_1(bn3_io_out_1),
    .io_out_2(bn3_io_out_2),
    .io_out_3(bn3_io_out_3),
    .io_out_4(bn3_io_out_4),
    .io_out_5(bn3_io_out_5),
    .io_out_6(bn3_io_out_6),
    .io_out_7(bn3_io_out_7),
    .io_out_8(bn3_io_out_8),
    .io_out_9(bn3_io_out_9)
  );
  assign io_out_0 = bn3_io_out_0;
  assign io_out_1 = bn3_io_out_1;
  assign io_out_2 = bn3_io_out_2;
  assign io_out_3 = bn3_io_out_3;
  assign io_out_4 = bn3_io_out_4;
  assign io_out_5 = bn3_io_out_5;
  assign io_out_6 = bn3_io_out_6;
  assign io_out_7 = bn3_io_out_7;
  assign io_out_8 = bn3_io_out_8;
  assign io_out_9 = bn3_io_out_9;
  assign fc1_io_in_0 = io_in_0;
  assign fc1_io_in_1 = io_in_1;
  assign fc1_io_in_2 = io_in_2;
  assign fc1_io_in_3 = io_in_3;
  assign fc1_io_in_4 = io_in_4;
  assign fc1_io_in_5 = io_in_5;
  assign fc1_io_in_6 = io_in_6;
  assign fc1_io_in_7 = io_in_7;
  assign fc1_io_in_8 = io_in_8;
  assign fc1_io_in_9 = io_in_9;
  assign fc1_io_in_10 = io_in_10;
  assign fc1_io_in_11 = io_in_11;
  assign fc1_io_in_12 = io_in_12;
  assign fc1_io_in_13 = io_in_13;
  assign fc1_io_in_14 = io_in_14;
  assign fc1_io_in_15 = io_in_15;
  assign fc1_io_in_16 = io_in_16;
  assign fc1_io_in_17 = io_in_17;
  assign fc1_io_in_18 = io_in_18;
  assign fc1_io_in_19 = io_in_19;
  assign fc1_io_in_20 = io_in_20;
  assign fc1_io_in_21 = io_in_21;
  assign fc1_io_in_22 = io_in_22;
  assign fc1_io_in_23 = io_in_23;
  assign fc1_io_in_24 = io_in_24;
  assign fc1_io_in_25 = io_in_25;
  assign fc1_io_in_26 = io_in_26;
  assign fc1_io_in_27 = io_in_27;
  assign fc1_io_in_28 = io_in_28;
  assign fc1_io_in_29 = io_in_29;
  assign fc1_io_in_30 = io_in_30;
  assign fc1_io_in_31 = io_in_31;
  assign fc1_io_in_32 = io_in_32;
  assign fc1_io_in_33 = io_in_33;
  assign fc1_io_in_34 = io_in_34;
  assign fc1_io_in_35 = io_in_35;
  assign fc1_io_in_36 = io_in_36;
  assign fc1_io_in_37 = io_in_37;
  assign fc1_io_in_38 = io_in_38;
  assign fc1_io_in_39 = io_in_39;
  assign fc1_io_in_40 = io_in_40;
  assign fc1_io_in_41 = io_in_41;
  assign fc1_io_in_42 = io_in_42;
  assign fc1_io_in_43 = io_in_43;
  assign fc1_io_in_44 = io_in_44;
  assign fc1_io_in_45 = io_in_45;
  assign fc1_io_in_46 = io_in_46;
  assign fc1_io_in_47 = io_in_47;
  assign fc1_io_in_48 = io_in_48;
  assign fc1_io_in_49 = io_in_49;
  assign fc1_io_in_50 = io_in_50;
  assign fc1_io_in_51 = io_in_51;
  assign fc1_io_in_52 = io_in_52;
  assign fc1_io_in_53 = io_in_53;
  assign fc1_io_in_54 = io_in_54;
  assign fc1_io_in_55 = io_in_55;
  assign fc1_io_in_56 = io_in_56;
  assign fc1_io_in_57 = io_in_57;
  assign fc1_io_in_58 = io_in_58;
  assign fc1_io_in_59 = io_in_59;
  assign fc1_io_in_60 = io_in_60;
  assign fc1_io_in_61 = io_in_61;
  assign fc1_io_in_62 = io_in_62;
  assign fc1_io_in_63 = io_in_63;
  assign fc1_io_in_64 = io_in_64;
  assign fc1_io_in_65 = io_in_65;
  assign fc1_io_in_66 = io_in_66;
  assign fc1_io_in_67 = io_in_67;
  assign fc1_io_in_68 = io_in_68;
  assign fc1_io_in_69 = io_in_69;
  assign fc1_io_in_70 = io_in_70;
  assign fc1_io_in_71 = io_in_71;
  assign fc1_io_in_72 = io_in_72;
  assign fc1_io_in_73 = io_in_73;
  assign fc1_io_in_74 = io_in_74;
  assign fc1_io_in_75 = io_in_75;
  assign fc1_io_in_76 = io_in_76;
  assign fc1_io_in_77 = io_in_77;
  assign fc1_io_in_78 = io_in_78;
  assign fc1_io_in_79 = io_in_79;
  assign fc1_io_in_80 = io_in_80;
  assign fc1_io_in_81 = io_in_81;
  assign fc1_io_in_82 = io_in_82;
  assign fc1_io_in_83 = io_in_83;
  assign fc1_io_in_84 = io_in_84;
  assign fc1_io_in_85 = io_in_85;
  assign fc1_io_in_86 = io_in_86;
  assign fc1_io_in_87 = io_in_87;
  assign fc1_io_in_88 = io_in_88;
  assign fc1_io_in_89 = io_in_89;
  assign fc1_io_in_90 = io_in_90;
  assign fc1_io_in_91 = io_in_91;
  assign fc1_io_in_92 = io_in_92;
  assign fc1_io_in_93 = io_in_93;
  assign fc1_io_in_94 = io_in_94;
  assign fc1_io_in_95 = io_in_95;
  assign fc1_io_in_96 = io_in_96;
  assign fc1_io_in_97 = io_in_97;
  assign fc1_io_in_98 = io_in_98;
  assign fc1_io_in_99 = io_in_99;
  assign fc1_io_in_100 = io_in_100;
  assign fc1_io_in_101 = io_in_101;
  assign fc1_io_in_102 = io_in_102;
  assign fc1_io_in_103 = io_in_103;
  assign fc1_io_in_104 = io_in_104;
  assign fc1_io_in_105 = io_in_105;
  assign fc1_io_in_106 = io_in_106;
  assign fc1_io_in_107 = io_in_107;
  assign fc1_io_in_108 = io_in_108;
  assign fc1_io_in_109 = io_in_109;
  assign fc1_io_in_110 = io_in_110;
  assign fc1_io_in_111 = io_in_111;
  assign fc1_io_in_112 = io_in_112;
  assign fc1_io_in_113 = io_in_113;
  assign fc1_io_in_114 = io_in_114;
  assign fc1_io_in_115 = io_in_115;
  assign fc1_io_in_116 = io_in_116;
  assign fc1_io_in_117 = io_in_117;
  assign fc1_io_in_118 = io_in_118;
  assign fc1_io_in_119 = io_in_119;
  assign fc1_io_in_120 = io_in_120;
  assign fc1_io_in_121 = io_in_121;
  assign fc1_io_in_122 = io_in_122;
  assign fc1_io_in_123 = io_in_123;
  assign fc1_io_in_124 = io_in_124;
  assign fc1_io_in_125 = io_in_125;
  assign fc1_io_in_126 = io_in_126;
  assign fc1_io_in_127 = io_in_127;
  assign fc1_io_in_128 = io_in_128;
  assign fc1_io_in_129 = io_in_129;
  assign fc1_io_in_130 = io_in_130;
  assign fc1_io_in_131 = io_in_131;
  assign fc1_io_in_132 = io_in_132;
  assign fc1_io_in_133 = io_in_133;
  assign fc1_io_in_134 = io_in_134;
  assign fc1_io_in_135 = io_in_135;
  assign fc1_io_in_136 = io_in_136;
  assign fc1_io_in_137 = io_in_137;
  assign fc1_io_in_138 = io_in_138;
  assign fc1_io_in_139 = io_in_139;
  assign fc1_io_in_140 = io_in_140;
  assign fc1_io_in_141 = io_in_141;
  assign fc1_io_in_142 = io_in_142;
  assign fc1_io_in_143 = io_in_143;
  assign fc1_io_in_144 = io_in_144;
  assign fc1_io_in_145 = io_in_145;
  assign fc1_io_in_146 = io_in_146;
  assign fc1_io_in_147 = io_in_147;
  assign fc1_io_in_148 = io_in_148;
  assign fc1_io_in_149 = io_in_149;
  assign fc1_io_in_150 = io_in_150;
  assign fc1_io_in_151 = io_in_151;
  assign fc1_io_in_152 = io_in_152;
  assign fc1_io_in_153 = io_in_153;
  assign fc1_io_in_154 = io_in_154;
  assign fc1_io_in_155 = io_in_155;
  assign fc1_io_in_156 = io_in_156;
  assign fc1_io_in_157 = io_in_157;
  assign fc1_io_in_158 = io_in_158;
  assign fc1_io_in_159 = io_in_159;
  assign fc1_io_in_160 = io_in_160;
  assign fc1_io_in_161 = io_in_161;
  assign fc1_io_in_162 = io_in_162;
  assign fc1_io_in_163 = io_in_163;
  assign fc1_io_in_164 = io_in_164;
  assign fc1_io_in_165 = io_in_165;
  assign fc1_io_in_166 = io_in_166;
  assign fc1_io_in_167 = io_in_167;
  assign fc1_io_in_168 = io_in_168;
  assign fc1_io_in_169 = io_in_169;
  assign fc1_io_in_170 = io_in_170;
  assign fc1_io_in_171 = io_in_171;
  assign fc1_io_in_172 = io_in_172;
  assign fc1_io_in_173 = io_in_173;
  assign fc1_io_in_174 = io_in_174;
  assign fc1_io_in_175 = io_in_175;
  assign fc1_io_in_176 = io_in_176;
  assign fc1_io_in_177 = io_in_177;
  assign fc1_io_in_178 = io_in_178;
  assign fc1_io_in_179 = io_in_179;
  assign fc1_io_in_180 = io_in_180;
  assign fc1_io_in_181 = io_in_181;
  assign fc1_io_in_182 = io_in_182;
  assign fc1_io_in_183 = io_in_183;
  assign fc1_io_in_184 = io_in_184;
  assign fc1_io_in_185 = io_in_185;
  assign fc1_io_in_186 = io_in_186;
  assign fc1_io_in_187 = io_in_187;
  assign fc1_io_in_188 = io_in_188;
  assign fc1_io_in_189 = io_in_189;
  assign fc1_io_in_190 = io_in_190;
  assign fc1_io_in_191 = io_in_191;
  assign fc1_io_in_192 = io_in_192;
  assign fc1_io_in_193 = io_in_193;
  assign fc1_io_in_194 = io_in_194;
  assign fc1_io_in_195 = io_in_195;
  assign fc1_io_in_196 = io_in_196;
  assign fc1_io_in_197 = io_in_197;
  assign fc1_io_in_198 = io_in_198;
  assign fc1_io_in_199 = io_in_199;
  assign fc1_io_in_200 = io_in_200;
  assign fc1_io_in_201 = io_in_201;
  assign fc1_io_in_202 = io_in_202;
  assign fc1_io_in_203 = io_in_203;
  assign fc1_io_in_204 = io_in_204;
  assign fc1_io_in_205 = io_in_205;
  assign fc1_io_in_206 = io_in_206;
  assign fc1_io_in_207 = io_in_207;
  assign fc1_io_in_208 = io_in_208;
  assign fc1_io_in_209 = io_in_209;
  assign fc1_io_in_210 = io_in_210;
  assign fc1_io_in_211 = io_in_211;
  assign fc1_io_in_212 = io_in_212;
  assign fc1_io_in_213 = io_in_213;
  assign fc1_io_in_214 = io_in_214;
  assign fc1_io_in_215 = io_in_215;
  assign fc1_io_in_216 = io_in_216;
  assign fc1_io_in_217 = io_in_217;
  assign fc1_io_in_218 = io_in_218;
  assign fc1_io_in_219 = io_in_219;
  assign fc1_io_in_220 = io_in_220;
  assign fc1_io_in_221 = io_in_221;
  assign fc1_io_in_222 = io_in_222;
  assign fc1_io_in_223 = io_in_223;
  assign fc1_io_in_224 = io_in_224;
  assign fc1_io_in_225 = io_in_225;
  assign fc1_io_in_226 = io_in_226;
  assign fc1_io_in_227 = io_in_227;
  assign fc1_io_in_228 = io_in_228;
  assign fc1_io_in_229 = io_in_229;
  assign fc1_io_in_230 = io_in_230;
  assign fc1_io_in_231 = io_in_231;
  assign fc1_io_in_232 = io_in_232;
  assign fc1_io_in_233 = io_in_233;
  assign fc1_io_in_234 = io_in_234;
  assign fc1_io_in_235 = io_in_235;
  assign fc1_io_in_236 = io_in_236;
  assign fc1_io_in_237 = io_in_237;
  assign fc1_io_in_238 = io_in_238;
  assign fc1_io_in_239 = io_in_239;
  assign fc1_io_in_240 = io_in_240;
  assign fc1_io_in_241 = io_in_241;
  assign fc1_io_in_242 = io_in_242;
  assign fc1_io_in_243 = io_in_243;
  assign fc1_io_in_244 = io_in_244;
  assign fc1_io_in_245 = io_in_245;
  assign fc1_io_in_246 = io_in_246;
  assign fc1_io_in_247 = io_in_247;
  assign fc1_io_in_248 = io_in_248;
  assign fc1_io_in_249 = io_in_249;
  assign fc1_io_in_250 = io_in_250;
  assign fc1_io_in_251 = io_in_251;
  assign fc1_io_in_252 = io_in_252;
  assign fc1_io_in_253 = io_in_253;
  assign fc1_io_in_254 = io_in_254;
  assign fc1_io_in_255 = io_in_255;
  assign fc1_io_in_256 = io_in_256;
  assign fc1_io_in_257 = io_in_257;
  assign fc1_io_in_258 = io_in_258;
  assign fc1_io_in_259 = io_in_259;
  assign fc1_io_in_260 = io_in_260;
  assign fc1_io_in_261 = io_in_261;
  assign fc1_io_in_262 = io_in_262;
  assign fc1_io_in_263 = io_in_263;
  assign fc1_io_in_264 = io_in_264;
  assign fc1_io_in_265 = io_in_265;
  assign fc1_io_in_266 = io_in_266;
  assign fc1_io_in_267 = io_in_267;
  assign fc1_io_in_268 = io_in_268;
  assign fc1_io_in_269 = io_in_269;
  assign fc1_io_in_270 = io_in_270;
  assign fc1_io_in_271 = io_in_271;
  assign fc1_io_in_272 = io_in_272;
  assign fc1_io_in_273 = io_in_273;
  assign fc1_io_in_274 = io_in_274;
  assign fc1_io_in_275 = io_in_275;
  assign fc1_io_in_276 = io_in_276;
  assign fc1_io_in_277 = io_in_277;
  assign fc1_io_in_278 = io_in_278;
  assign fc1_io_in_279 = io_in_279;
  assign fc1_io_in_280 = io_in_280;
  assign fc1_io_in_281 = io_in_281;
  assign fc1_io_in_282 = io_in_282;
  assign fc1_io_in_283 = io_in_283;
  assign fc1_io_in_284 = io_in_284;
  assign fc1_io_in_285 = io_in_285;
  assign fc1_io_in_286 = io_in_286;
  assign fc1_io_in_287 = io_in_287;
  assign fc1_io_in_288 = io_in_288;
  assign fc1_io_in_289 = io_in_289;
  assign fc1_io_in_290 = io_in_290;
  assign fc1_io_in_291 = io_in_291;
  assign fc1_io_in_292 = io_in_292;
  assign fc1_io_in_293 = io_in_293;
  assign fc1_io_in_294 = io_in_294;
  assign fc1_io_in_295 = io_in_295;
  assign fc1_io_in_296 = io_in_296;
  assign fc1_io_in_297 = io_in_297;
  assign fc1_io_in_298 = io_in_298;
  assign fc1_io_in_299 = io_in_299;
  assign fc1_io_in_300 = io_in_300;
  assign fc1_io_in_301 = io_in_301;
  assign fc1_io_in_302 = io_in_302;
  assign fc1_io_in_303 = io_in_303;
  assign fc1_io_in_304 = io_in_304;
  assign fc1_io_in_305 = io_in_305;
  assign fc1_io_in_306 = io_in_306;
  assign fc1_io_in_307 = io_in_307;
  assign fc1_io_in_308 = io_in_308;
  assign fc1_io_in_309 = io_in_309;
  assign fc1_io_in_310 = io_in_310;
  assign fc1_io_in_311 = io_in_311;
  assign fc1_io_in_312 = io_in_312;
  assign fc1_io_in_313 = io_in_313;
  assign fc1_io_in_314 = io_in_314;
  assign fc1_io_in_315 = io_in_315;
  assign fc1_io_in_316 = io_in_316;
  assign fc1_io_in_317 = io_in_317;
  assign fc1_io_in_318 = io_in_318;
  assign fc1_io_in_319 = io_in_319;
  assign fc1_io_in_320 = io_in_320;
  assign fc1_io_in_321 = io_in_321;
  assign fc1_io_in_322 = io_in_322;
  assign fc1_io_in_323 = io_in_323;
  assign fc1_io_in_324 = io_in_324;
  assign fc1_io_in_325 = io_in_325;
  assign fc1_io_in_326 = io_in_326;
  assign fc1_io_in_327 = io_in_327;
  assign fc1_io_in_328 = io_in_328;
  assign fc1_io_in_329 = io_in_329;
  assign fc1_io_in_330 = io_in_330;
  assign fc1_io_in_331 = io_in_331;
  assign fc1_io_in_332 = io_in_332;
  assign fc1_io_in_333 = io_in_333;
  assign fc1_io_in_334 = io_in_334;
  assign fc1_io_in_335 = io_in_335;
  assign fc1_io_in_336 = io_in_336;
  assign fc1_io_in_337 = io_in_337;
  assign fc1_io_in_338 = io_in_338;
  assign fc1_io_in_339 = io_in_339;
  assign fc1_io_in_340 = io_in_340;
  assign fc1_io_in_341 = io_in_341;
  assign fc1_io_in_342 = io_in_342;
  assign fc1_io_in_343 = io_in_343;
  assign fc1_io_in_344 = io_in_344;
  assign fc1_io_in_345 = io_in_345;
  assign fc1_io_in_346 = io_in_346;
  assign fc1_io_in_347 = io_in_347;
  assign fc1_io_in_348 = io_in_348;
  assign fc1_io_in_349 = io_in_349;
  assign fc1_io_in_350 = io_in_350;
  assign fc1_io_in_351 = io_in_351;
  assign fc1_io_in_352 = io_in_352;
  assign fc1_io_in_353 = io_in_353;
  assign fc1_io_in_354 = io_in_354;
  assign fc1_io_in_355 = io_in_355;
  assign fc1_io_in_356 = io_in_356;
  assign fc1_io_in_357 = io_in_357;
  assign fc1_io_in_358 = io_in_358;
  assign fc1_io_in_359 = io_in_359;
  assign fc1_io_in_360 = io_in_360;
  assign fc1_io_in_361 = io_in_361;
  assign fc1_io_in_362 = io_in_362;
  assign fc1_io_in_363 = io_in_363;
  assign fc1_io_in_364 = io_in_364;
  assign fc1_io_in_365 = io_in_365;
  assign fc1_io_in_366 = io_in_366;
  assign fc1_io_in_367 = io_in_367;
  assign fc1_io_in_368 = io_in_368;
  assign fc1_io_in_369 = io_in_369;
  assign fc1_io_in_370 = io_in_370;
  assign fc1_io_in_371 = io_in_371;
  assign fc1_io_in_372 = io_in_372;
  assign fc1_io_in_373 = io_in_373;
  assign fc1_io_in_374 = io_in_374;
  assign fc1_io_in_375 = io_in_375;
  assign fc1_io_in_376 = io_in_376;
  assign fc1_io_in_377 = io_in_377;
  assign fc1_io_in_378 = io_in_378;
  assign fc1_io_in_379 = io_in_379;
  assign fc1_io_in_380 = io_in_380;
  assign fc1_io_in_381 = io_in_381;
  assign fc1_io_in_382 = io_in_382;
  assign fc1_io_in_383 = io_in_383;
  assign fc1_io_in_384 = io_in_384;
  assign fc1_io_in_385 = io_in_385;
  assign fc1_io_in_386 = io_in_386;
  assign fc1_io_in_387 = io_in_387;
  assign fc1_io_in_388 = io_in_388;
  assign fc1_io_in_389 = io_in_389;
  assign fc1_io_in_390 = io_in_390;
  assign fc1_io_in_391 = io_in_391;
  assign fc1_io_in_392 = io_in_392;
  assign fc1_io_in_393 = io_in_393;
  assign fc1_io_in_394 = io_in_394;
  assign fc1_io_in_395 = io_in_395;
  assign fc1_io_in_396 = io_in_396;
  assign fc1_io_in_397 = io_in_397;
  assign fc1_io_in_398 = io_in_398;
  assign fc1_io_in_399 = io_in_399;
  assign fc1_io_in_400 = io_in_400;
  assign fc1_io_in_401 = io_in_401;
  assign fc1_io_in_402 = io_in_402;
  assign fc1_io_in_403 = io_in_403;
  assign fc1_io_in_404 = io_in_404;
  assign fc1_io_in_405 = io_in_405;
  assign fc1_io_in_406 = io_in_406;
  assign fc1_io_in_407 = io_in_407;
  assign fc1_io_in_408 = io_in_408;
  assign fc1_io_in_409 = io_in_409;
  assign fc1_io_in_410 = io_in_410;
  assign fc1_io_in_411 = io_in_411;
  assign fc1_io_in_412 = io_in_412;
  assign fc1_io_in_413 = io_in_413;
  assign fc1_io_in_414 = io_in_414;
  assign fc1_io_in_415 = io_in_415;
  assign fc1_io_in_416 = io_in_416;
  assign fc1_io_in_417 = io_in_417;
  assign fc1_io_in_418 = io_in_418;
  assign fc1_io_in_419 = io_in_419;
  assign fc1_io_in_420 = io_in_420;
  assign fc1_io_in_421 = io_in_421;
  assign fc1_io_in_422 = io_in_422;
  assign fc1_io_in_423 = io_in_423;
  assign fc1_io_in_424 = io_in_424;
  assign fc1_io_in_425 = io_in_425;
  assign fc1_io_in_426 = io_in_426;
  assign fc1_io_in_427 = io_in_427;
  assign fc1_io_in_428 = io_in_428;
  assign fc1_io_in_429 = io_in_429;
  assign fc1_io_in_430 = io_in_430;
  assign fc1_io_in_431 = io_in_431;
  assign fc1_io_in_432 = io_in_432;
  assign fc1_io_in_433 = io_in_433;
  assign fc1_io_in_434 = io_in_434;
  assign fc1_io_in_435 = io_in_435;
  assign fc1_io_in_436 = io_in_436;
  assign fc1_io_in_437 = io_in_437;
  assign fc1_io_in_438 = io_in_438;
  assign fc1_io_in_439 = io_in_439;
  assign fc1_io_in_440 = io_in_440;
  assign fc1_io_in_441 = io_in_441;
  assign fc1_io_in_442 = io_in_442;
  assign fc1_io_in_443 = io_in_443;
  assign fc1_io_in_444 = io_in_444;
  assign fc1_io_in_445 = io_in_445;
  assign fc1_io_in_446 = io_in_446;
  assign fc1_io_in_447 = io_in_447;
  assign fc1_io_in_448 = io_in_448;
  assign fc1_io_in_449 = io_in_449;
  assign fc1_io_in_450 = io_in_450;
  assign fc1_io_in_451 = io_in_451;
  assign fc1_io_in_452 = io_in_452;
  assign fc1_io_in_453 = io_in_453;
  assign fc1_io_in_454 = io_in_454;
  assign fc1_io_in_455 = io_in_455;
  assign fc1_io_in_456 = io_in_456;
  assign fc1_io_in_457 = io_in_457;
  assign fc1_io_in_458 = io_in_458;
  assign fc1_io_in_459 = io_in_459;
  assign fc1_io_in_460 = io_in_460;
  assign fc1_io_in_461 = io_in_461;
  assign fc1_io_in_462 = io_in_462;
  assign fc1_io_in_463 = io_in_463;
  assign fc1_io_in_464 = io_in_464;
  assign fc1_io_in_465 = io_in_465;
  assign fc1_io_in_466 = io_in_466;
  assign fc1_io_in_467 = io_in_467;
  assign fc1_io_in_468 = io_in_468;
  assign fc1_io_in_469 = io_in_469;
  assign fc1_io_in_470 = io_in_470;
  assign fc1_io_in_471 = io_in_471;
  assign fc1_io_in_472 = io_in_472;
  assign fc1_io_in_473 = io_in_473;
  assign fc1_io_in_474 = io_in_474;
  assign fc1_io_in_475 = io_in_475;
  assign fc1_io_in_476 = io_in_476;
  assign fc1_io_in_477 = io_in_477;
  assign fc1_io_in_478 = io_in_478;
  assign fc1_io_in_479 = io_in_479;
  assign fc1_io_in_480 = io_in_480;
  assign fc1_io_in_481 = io_in_481;
  assign fc1_io_in_482 = io_in_482;
  assign fc1_io_in_483 = io_in_483;
  assign fc1_io_in_484 = io_in_484;
  assign fc1_io_in_485 = io_in_485;
  assign fc1_io_in_486 = io_in_486;
  assign fc1_io_in_487 = io_in_487;
  assign fc1_io_in_488 = io_in_488;
  assign fc1_io_in_489 = io_in_489;
  assign fc1_io_in_490 = io_in_490;
  assign fc1_io_in_491 = io_in_491;
  assign fc1_io_in_492 = io_in_492;
  assign fc1_io_in_493 = io_in_493;
  assign fc1_io_in_494 = io_in_494;
  assign fc1_io_in_495 = io_in_495;
  assign fc1_io_in_496 = io_in_496;
  assign fc1_io_in_497 = io_in_497;
  assign fc1_io_in_498 = io_in_498;
  assign fc1_io_in_499 = io_in_499;
  assign fc1_io_in_500 = io_in_500;
  assign fc1_io_in_501 = io_in_501;
  assign fc1_io_in_502 = io_in_502;
  assign fc1_io_in_503 = io_in_503;
  assign fc1_io_in_504 = io_in_504;
  assign fc1_io_in_505 = io_in_505;
  assign fc1_io_in_506 = io_in_506;
  assign fc1_io_in_507 = io_in_507;
  assign fc1_io_in_508 = io_in_508;
  assign fc1_io_in_509 = io_in_509;
  assign fc1_io_in_510 = io_in_510;
  assign fc1_io_in_511 = io_in_511;
  assign fc1_io_in_512 = io_in_512;
  assign fc1_io_in_513 = io_in_513;
  assign fc1_io_in_514 = io_in_514;
  assign fc1_io_in_515 = io_in_515;
  assign fc1_io_in_516 = io_in_516;
  assign fc1_io_in_517 = io_in_517;
  assign fc1_io_in_518 = io_in_518;
  assign fc1_io_in_519 = io_in_519;
  assign fc1_io_in_520 = io_in_520;
  assign fc1_io_in_521 = io_in_521;
  assign fc1_io_in_522 = io_in_522;
  assign fc1_io_in_523 = io_in_523;
  assign fc1_io_in_524 = io_in_524;
  assign fc1_io_in_525 = io_in_525;
  assign fc1_io_in_526 = io_in_526;
  assign fc1_io_in_527 = io_in_527;
  assign fc1_io_in_528 = io_in_528;
  assign fc1_io_in_529 = io_in_529;
  assign fc1_io_in_530 = io_in_530;
  assign fc1_io_in_531 = io_in_531;
  assign fc1_io_in_532 = io_in_532;
  assign fc1_io_in_533 = io_in_533;
  assign fc1_io_in_534 = io_in_534;
  assign fc1_io_in_535 = io_in_535;
  assign fc1_io_in_536 = io_in_536;
  assign fc1_io_in_537 = io_in_537;
  assign fc1_io_in_538 = io_in_538;
  assign fc1_io_in_539 = io_in_539;
  assign fc1_io_in_540 = io_in_540;
  assign fc1_io_in_541 = io_in_541;
  assign fc1_io_in_542 = io_in_542;
  assign fc1_io_in_543 = io_in_543;
  assign fc1_io_in_544 = io_in_544;
  assign fc1_io_in_545 = io_in_545;
  assign fc1_io_in_546 = io_in_546;
  assign fc1_io_in_547 = io_in_547;
  assign fc1_io_in_548 = io_in_548;
  assign fc1_io_in_549 = io_in_549;
  assign fc1_io_in_550 = io_in_550;
  assign fc1_io_in_551 = io_in_551;
  assign fc1_io_in_552 = io_in_552;
  assign fc1_io_in_553 = io_in_553;
  assign fc1_io_in_554 = io_in_554;
  assign fc1_io_in_555 = io_in_555;
  assign fc1_io_in_556 = io_in_556;
  assign fc1_io_in_557 = io_in_557;
  assign fc1_io_in_558 = io_in_558;
  assign fc1_io_in_559 = io_in_559;
  assign fc1_io_in_560 = io_in_560;
  assign fc1_io_in_561 = io_in_561;
  assign fc1_io_in_562 = io_in_562;
  assign fc1_io_in_563 = io_in_563;
  assign fc1_io_in_564 = io_in_564;
  assign fc1_io_in_565 = io_in_565;
  assign fc1_io_in_566 = io_in_566;
  assign fc1_io_in_567 = io_in_567;
  assign fc1_io_in_568 = io_in_568;
  assign fc1_io_in_569 = io_in_569;
  assign fc1_io_in_570 = io_in_570;
  assign fc1_io_in_571 = io_in_571;
  assign fc1_io_in_572 = io_in_572;
  assign fc1_io_in_573 = io_in_573;
  assign fc1_io_in_574 = io_in_574;
  assign fc1_io_in_575 = io_in_575;
  assign fc1_io_in_576 = io_in_576;
  assign fc1_io_in_577 = io_in_577;
  assign fc1_io_in_578 = io_in_578;
  assign fc1_io_in_579 = io_in_579;
  assign fc1_io_in_580 = io_in_580;
  assign fc1_io_in_581 = io_in_581;
  assign fc1_io_in_582 = io_in_582;
  assign fc1_io_in_583 = io_in_583;
  assign fc1_io_in_584 = io_in_584;
  assign fc1_io_in_585 = io_in_585;
  assign fc1_io_in_586 = io_in_586;
  assign fc1_io_in_587 = io_in_587;
  assign fc1_io_in_588 = io_in_588;
  assign fc1_io_in_589 = io_in_589;
  assign fc1_io_in_590 = io_in_590;
  assign fc1_io_in_591 = io_in_591;
  assign fc1_io_in_592 = io_in_592;
  assign fc1_io_in_593 = io_in_593;
  assign fc1_io_in_594 = io_in_594;
  assign fc1_io_in_595 = io_in_595;
  assign fc1_io_in_596 = io_in_596;
  assign fc1_io_in_597 = io_in_597;
  assign fc1_io_in_598 = io_in_598;
  assign fc1_io_in_599 = io_in_599;
  assign fc1_io_in_600 = io_in_600;
  assign fc1_io_in_601 = io_in_601;
  assign fc1_io_in_602 = io_in_602;
  assign fc1_io_in_603 = io_in_603;
  assign fc1_io_in_604 = io_in_604;
  assign fc1_io_in_605 = io_in_605;
  assign fc1_io_in_606 = io_in_606;
  assign fc1_io_in_607 = io_in_607;
  assign fc1_io_in_608 = io_in_608;
  assign fc1_io_in_609 = io_in_609;
  assign fc1_io_in_610 = io_in_610;
  assign fc1_io_in_611 = io_in_611;
  assign fc1_io_in_612 = io_in_612;
  assign fc1_io_in_613 = io_in_613;
  assign fc1_io_in_614 = io_in_614;
  assign fc1_io_in_615 = io_in_615;
  assign fc1_io_in_616 = io_in_616;
  assign fc1_io_in_617 = io_in_617;
  assign fc1_io_in_618 = io_in_618;
  assign fc1_io_in_619 = io_in_619;
  assign fc1_io_in_620 = io_in_620;
  assign fc1_io_in_621 = io_in_621;
  assign fc1_io_in_622 = io_in_622;
  assign fc1_io_in_623 = io_in_623;
  assign fc1_io_in_624 = io_in_624;
  assign fc1_io_in_625 = io_in_625;
  assign fc1_io_in_626 = io_in_626;
  assign fc1_io_in_627 = io_in_627;
  assign fc1_io_in_628 = io_in_628;
  assign fc1_io_in_629 = io_in_629;
  assign fc1_io_in_630 = io_in_630;
  assign fc1_io_in_631 = io_in_631;
  assign fc1_io_in_632 = io_in_632;
  assign fc1_io_in_633 = io_in_633;
  assign fc1_io_in_634 = io_in_634;
  assign fc1_io_in_635 = io_in_635;
  assign fc1_io_in_636 = io_in_636;
  assign fc1_io_in_637 = io_in_637;
  assign fc1_io_in_638 = io_in_638;
  assign fc1_io_in_639 = io_in_639;
  assign fc1_io_in_640 = io_in_640;
  assign fc1_io_in_641 = io_in_641;
  assign fc1_io_in_642 = io_in_642;
  assign fc1_io_in_643 = io_in_643;
  assign fc1_io_in_644 = io_in_644;
  assign fc1_io_in_645 = io_in_645;
  assign fc1_io_in_646 = io_in_646;
  assign fc1_io_in_647 = io_in_647;
  assign fc1_io_in_648 = io_in_648;
  assign fc1_io_in_649 = io_in_649;
  assign fc1_io_in_650 = io_in_650;
  assign fc1_io_in_651 = io_in_651;
  assign fc1_io_in_652 = io_in_652;
  assign fc1_io_in_653 = io_in_653;
  assign fc1_io_in_654 = io_in_654;
  assign fc1_io_in_655 = io_in_655;
  assign fc1_io_in_656 = io_in_656;
  assign fc1_io_in_657 = io_in_657;
  assign fc1_io_in_658 = io_in_658;
  assign fc1_io_in_659 = io_in_659;
  assign fc1_io_in_660 = io_in_660;
  assign fc1_io_in_661 = io_in_661;
  assign fc1_io_in_662 = io_in_662;
  assign fc1_io_in_663 = io_in_663;
  assign fc1_io_in_664 = io_in_664;
  assign fc1_io_in_665 = io_in_665;
  assign fc1_io_in_666 = io_in_666;
  assign fc1_io_in_667 = io_in_667;
  assign fc1_io_in_668 = io_in_668;
  assign fc1_io_in_669 = io_in_669;
  assign fc1_io_in_670 = io_in_670;
  assign fc1_io_in_671 = io_in_671;
  assign fc1_io_in_672 = io_in_672;
  assign fc1_io_in_673 = io_in_673;
  assign fc1_io_in_674 = io_in_674;
  assign fc1_io_in_675 = io_in_675;
  assign fc1_io_in_676 = io_in_676;
  assign fc1_io_in_677 = io_in_677;
  assign fc1_io_in_678 = io_in_678;
  assign fc1_io_in_679 = io_in_679;
  assign fc1_io_in_680 = io_in_680;
  assign fc1_io_in_681 = io_in_681;
  assign fc1_io_in_682 = io_in_682;
  assign fc1_io_in_683 = io_in_683;
  assign fc1_io_in_684 = io_in_684;
  assign fc1_io_in_685 = io_in_685;
  assign fc1_io_in_686 = io_in_686;
  assign fc1_io_in_687 = io_in_687;
  assign fc1_io_in_688 = io_in_688;
  assign fc1_io_in_689 = io_in_689;
  assign fc1_io_in_690 = io_in_690;
  assign fc1_io_in_691 = io_in_691;
  assign fc1_io_in_692 = io_in_692;
  assign fc1_io_in_693 = io_in_693;
  assign fc1_io_in_694 = io_in_694;
  assign fc1_io_in_695 = io_in_695;
  assign fc1_io_in_696 = io_in_696;
  assign fc1_io_in_697 = io_in_697;
  assign fc1_io_in_698 = io_in_698;
  assign fc1_io_in_699 = io_in_699;
  assign fc1_io_in_700 = io_in_700;
  assign fc1_io_in_701 = io_in_701;
  assign fc1_io_in_702 = io_in_702;
  assign fc1_io_in_703 = io_in_703;
  assign fc1_io_in_704 = io_in_704;
  assign fc1_io_in_705 = io_in_705;
  assign fc1_io_in_706 = io_in_706;
  assign fc1_io_in_707 = io_in_707;
  assign fc1_io_in_708 = io_in_708;
  assign fc1_io_in_709 = io_in_709;
  assign fc1_io_in_710 = io_in_710;
  assign fc1_io_in_711 = io_in_711;
  assign fc1_io_in_712 = io_in_712;
  assign fc1_io_in_713 = io_in_713;
  assign fc1_io_in_714 = io_in_714;
  assign fc1_io_in_715 = io_in_715;
  assign fc1_io_in_716 = io_in_716;
  assign fc1_io_in_717 = io_in_717;
  assign fc1_io_in_718 = io_in_718;
  assign fc1_io_in_719 = io_in_719;
  assign fc1_io_in_720 = io_in_720;
  assign fc1_io_in_721 = io_in_721;
  assign fc1_io_in_722 = io_in_722;
  assign fc1_io_in_723 = io_in_723;
  assign fc1_io_in_724 = io_in_724;
  assign fc1_io_in_725 = io_in_725;
  assign fc1_io_in_726 = io_in_726;
  assign fc1_io_in_727 = io_in_727;
  assign fc1_io_in_728 = io_in_728;
  assign fc1_io_in_729 = io_in_729;
  assign fc1_io_in_730 = io_in_730;
  assign fc1_io_in_731 = io_in_731;
  assign fc1_io_in_732 = io_in_732;
  assign fc1_io_in_733 = io_in_733;
  assign fc1_io_in_734 = io_in_734;
  assign fc1_io_in_735 = io_in_735;
  assign fc1_io_in_736 = io_in_736;
  assign fc1_io_in_737 = io_in_737;
  assign fc1_io_in_738 = io_in_738;
  assign fc1_io_in_739 = io_in_739;
  assign fc1_io_in_740 = io_in_740;
  assign fc1_io_in_741 = io_in_741;
  assign fc1_io_in_742 = io_in_742;
  assign fc1_io_in_743 = io_in_743;
  assign fc1_io_in_744 = io_in_744;
  assign fc1_io_in_745 = io_in_745;
  assign fc1_io_in_746 = io_in_746;
  assign fc1_io_in_747 = io_in_747;
  assign fc1_io_in_748 = io_in_748;
  assign fc1_io_in_749 = io_in_749;
  assign fc1_io_in_750 = io_in_750;
  assign fc1_io_in_751 = io_in_751;
  assign fc1_io_in_752 = io_in_752;
  assign fc1_io_in_753 = io_in_753;
  assign fc1_io_in_754 = io_in_754;
  assign fc1_io_in_755 = io_in_755;
  assign fc1_io_in_756 = io_in_756;
  assign fc1_io_in_757 = io_in_757;
  assign fc1_io_in_758 = io_in_758;
  assign fc1_io_in_759 = io_in_759;
  assign fc1_io_in_760 = io_in_760;
  assign fc1_io_in_761 = io_in_761;
  assign fc1_io_in_762 = io_in_762;
  assign fc1_io_in_763 = io_in_763;
  assign fc1_io_in_764 = io_in_764;
  assign fc1_io_in_765 = io_in_765;
  assign fc1_io_in_766 = io_in_766;
  assign fc1_io_in_767 = io_in_767;
  assign fc1_io_in_768 = io_in_768;
  assign fc1_io_in_769 = io_in_769;
  assign fc1_io_in_770 = io_in_770;
  assign fc1_io_in_771 = io_in_771;
  assign fc1_io_in_772 = io_in_772;
  assign fc1_io_in_773 = io_in_773;
  assign fc1_io_in_774 = io_in_774;
  assign fc1_io_in_775 = io_in_775;
  assign fc1_io_in_776 = io_in_776;
  assign fc1_io_in_777 = io_in_777;
  assign fc1_io_in_778 = io_in_778;
  assign fc1_io_in_779 = io_in_779;
  assign fc1_io_in_780 = io_in_780;
  assign fc1_io_in_781 = io_in_781;
  assign fc1_io_in_782 = io_in_782;
  assign fc1_io_in_783 = io_in_783;
  assign bn1_io_in_0 = fc1_io_out_0;
  assign bn1_io_in_1 = fc1_io_out_1;
  assign bn1_io_in_2 = fc1_io_out_2;
  assign bn1_io_in_3 = fc1_io_out_3;
  assign bn1_io_in_4 = fc1_io_out_4;
  assign bn1_io_in_5 = fc1_io_out_5;
  assign bn1_io_in_6 = fc1_io_out_6;
  assign bn1_io_in_7 = fc1_io_out_7;
  assign bn1_io_in_8 = fc1_io_out_8;
  assign bn1_io_in_9 = fc1_io_out_9;
  assign bn1_io_in_10 = fc1_io_out_10;
  assign bn1_io_in_11 = fc1_io_out_11;
  assign bn1_io_in_12 = fc1_io_out_12;
  assign bn1_io_in_13 = fc1_io_out_13;
  assign bn1_io_in_14 = fc1_io_out_14;
  assign bn1_io_in_15 = fc1_io_out_15;
  assign bi1_io_in_0 = bn1_io_out_0;
  assign bi1_io_in_1 = bn1_io_out_1;
  assign bi1_io_in_2 = bn1_io_out_2;
  assign bi1_io_in_3 = bn1_io_out_3;
  assign bi1_io_in_4 = bn1_io_out_4;
  assign bi1_io_in_5 = bn1_io_out_5;
  assign bi1_io_in_6 = bn1_io_out_6;
  assign bi1_io_in_7 = bn1_io_out_7;
  assign bi1_io_in_8 = bn1_io_out_8;
  assign bi1_io_in_9 = bn1_io_out_9;
  assign bi1_io_in_10 = bn1_io_out_10;
  assign bi1_io_in_11 = bn1_io_out_11;
  assign bi1_io_in_12 = bn1_io_out_12;
  assign bi1_io_in_13 = bn1_io_out_13;
  assign bi1_io_in_14 = bn1_io_out_14;
  assign bi1_io_in_15 = bn1_io_out_15;
  assign fc2_io_in_0 = bi1_io_out_0;
  assign fc2_io_in_1 = bi1_io_out_1;
  assign fc2_io_in_2 = bi1_io_out_2;
  assign fc2_io_in_3 = bi1_io_out_3;
  assign fc2_io_in_4 = bi1_io_out_4;
  assign fc2_io_in_5 = bi1_io_out_5;
  assign fc2_io_in_6 = bi1_io_out_6;
  assign fc2_io_in_7 = bi1_io_out_7;
  assign fc2_io_in_8 = bi1_io_out_8;
  assign fc2_io_in_9 = bi1_io_out_9;
  assign fc2_io_in_10 = bi1_io_out_10;
  assign fc2_io_in_11 = bi1_io_out_11;
  assign fc2_io_in_12 = bi1_io_out_12;
  assign fc2_io_in_13 = bi1_io_out_13;
  assign fc2_io_in_14 = bi1_io_out_14;
  assign fc2_io_in_15 = bi1_io_out_15;
  assign bn2_io_in_0 = fc2_io_out_0;
  assign bn2_io_in_1 = fc2_io_out_1;
  assign bn2_io_in_2 = fc2_io_out_2;
  assign bn2_io_in_3 = fc2_io_out_3;
  assign bn2_io_in_4 = fc2_io_out_4;
  assign bn2_io_in_5 = fc2_io_out_5;
  assign bn2_io_in_6 = fc2_io_out_6;
  assign bn2_io_in_7 = fc2_io_out_7;
  assign bn2_io_in_8 = fc2_io_out_8;
  assign bn2_io_in_9 = fc2_io_out_9;
  assign bn2_io_in_10 = fc2_io_out_10;
  assign bn2_io_in_11 = fc2_io_out_11;
  assign bn2_io_in_12 = fc2_io_out_12;
  assign bn2_io_in_13 = fc2_io_out_13;
  assign bn2_io_in_14 = fc2_io_out_14;
  assign bn2_io_in_15 = fc2_io_out_15;
  assign bi2_io_in_0 = bn2_io_out_0;
  assign bi2_io_in_1 = bn2_io_out_1;
  assign bi2_io_in_2 = bn2_io_out_2;
  assign bi2_io_in_3 = bn2_io_out_3;
  assign bi2_io_in_4 = bn2_io_out_4;
  assign bi2_io_in_5 = bn2_io_out_5;
  assign bi2_io_in_6 = bn2_io_out_6;
  assign bi2_io_in_7 = bn2_io_out_7;
  assign bi2_io_in_8 = bn2_io_out_8;
  assign bi2_io_in_9 = bn2_io_out_9;
  assign bi2_io_in_10 = bn2_io_out_10;
  assign bi2_io_in_11 = bn2_io_out_11;
  assign bi2_io_in_12 = bn2_io_out_12;
  assign bi2_io_in_13 = bn2_io_out_13;
  assign bi2_io_in_14 = bn2_io_out_14;
  assign bi2_io_in_15 = bn2_io_out_15;
  assign fc3_io_in_0 = bi2_io_out_0;
  assign fc3_io_in_1 = bi2_io_out_1;
  assign fc3_io_in_2 = bi2_io_out_2;
  assign fc3_io_in_3 = bi2_io_out_3;
  assign fc3_io_in_4 = bi2_io_out_4;
  assign fc3_io_in_5 = bi2_io_out_5;
  assign fc3_io_in_6 = bi2_io_out_6;
  assign fc3_io_in_7 = bi2_io_out_7;
  assign fc3_io_in_8 = bi2_io_out_8;
  assign fc3_io_in_9 = bi2_io_out_9;
  assign fc3_io_in_10 = bi2_io_out_10;
  assign fc3_io_in_11 = bi2_io_out_11;
  assign fc3_io_in_12 = bi2_io_out_12;
  assign fc3_io_in_13 = bi2_io_out_13;
  assign fc3_io_in_14 = bi2_io_out_14;
  assign fc3_io_in_15 = bi2_io_out_15;
  assign bn3_io_in_0 = fc3_io_out_0;
  assign bn3_io_in_1 = fc3_io_out_1;
  assign bn3_io_in_2 = fc3_io_out_2;
  assign bn3_io_in_3 = fc3_io_out_3;
  assign bn3_io_in_4 = fc3_io_out_4;
  assign bn3_io_in_5 = fc3_io_out_5;
  assign bn3_io_in_6 = fc3_io_out_6;
  assign bn3_io_in_7 = fc3_io_out_7;
  assign bn3_io_in_8 = fc3_io_out_8;
  assign bn3_io_in_9 = fc3_io_out_9;
endmodule
